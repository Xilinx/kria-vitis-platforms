/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dD6sJjMckNM/hk590wWgo7QyLBP7qvuv1GnV/mfQB0w/i/pvS4BJcnppdBuizaQbHZTE85H6pboO
mTjEC8kS1yUyaRKX4KpOmRsaXVL7/iV6Mc+EyHoad/3cx2lAwTCRu6nptqi96Q/dtiPbQirlE0cr
bj2VslWvQXYp7agPImHpkldpbIx4OKKY49/lmZgzjQmz1uAl0Vpqn03TZsorFhKrWNa1NL2PWEvy
H6r6Q2NnxwJibsxIu7/DaDQZ9tx7P3Ox5rT/+t7OV/sWKJMNsqkendhSkyxMCR6Z1Ip9YxyEItGS
Bld1ucslP9zp60t9CzMGZcj/WZZ+ve1NzjV/uw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="NlHs8opBWv2KH1hFnLsdY2EH/Cy8LVzvJ0P9w8zUaYI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3008)
`pragma protect data_block
jOrE4515xgbASXSOIDgmJkXcXt7RETFe/mPq2BnvaRJwyPFDl1smas20v70GQpkf3qeD7bj7sIlp
z07fV96t9+2VpKfAOu6WpsTNkYx3HoKr5g4kzIMGPaao5qirLmlvZJPo13d3FcbazVTeHp1Kg68X
T+q9vHvyJkRGDfJbq6g7uWe9pDCEkA/lQhh7DDK/tHi9Sk/qUWjlH37meqgzDIn/cojxAD6A1NZ9
GtlKHIOSQibGw7ipVgbo49t/jMjgj9b6lsuu34icdAvJWYJVPLzXIIVdfRxZQc3Ys/7hw6/JJbC3
W0lBVlMrtGa4tWAmBxCs4XN2VnLI7j1mbhPAR33qw2mFUU7TPnGJGFirL3jGsSR767vMOYFYOpKt
IeRYghVIduSfGrKP38vmYdxP4X2G0zuGBGOg4EdNdMRLmBKTL5/EH0kKxeBmBduT+xeAu7MN2xzf
g45FohodAm8rLjNvgInZ7WV/dYDqOK408Kd7OK0OZFAu3fMISVzP9kr46Fg5GQFbRkXJHvdMBltH
4A43/GCP+mPq+OAqZ55Z9yXfrmLjtP4HAFyfFZ0k2Blj+ZUl2YISBdc2i8qSRkVl1fHlC7C1hjNd
jCLCV2Grfq9ARcflyU+jok8RFgnwgjD3M43Loi5tdoYKoymmJkMSkuc9D1tOIg3SgJ01UE028swv
EhTWV+LxrwHTH/XbkQf9R8wNOtm4PS2ZqNHwob3uWd9eavm5zNWaigTve5T9xds+9hIJZoY1isC0
WzoR0iduNXKKYXDZZpYwjliHfcOKu2rjSvRSSaFazGUammbMczhytVIwghtsUSMn2cXpJHGyaicJ
OAoWWUVFDqYMmg3vPAoPuX5Ii/4ISf5LILwlYImyIhnnurwEL8V05eXcRs0H9gVAXS9Bx9B2KoY+
V08LMq7unYvEfI+dLWiNIYPHhpbuD6T7idgqU0PCxsa46qzqLa6eYtXrNQ/QwlQwjQSdG9PXS682
s1mnHdF1N7roKihS3vMtWQqfbgr4N/RtFw3DzuX4Fbxr4FQtaVaXKGT/R1Mk8lVFZwV+QkjD0mTi
Ttv3KNWYq4yIAFgBVAYNea/64ZmwimBhJ9sFQom7GApoGn44OTDbLW3cQgDGQy9IcT19/crS0KgU
5vvoZRF+3FRa4jY3+5knJBLD38na4X9nbXSn65lzTdk4vlGolSs8hZ0qCI4dX1u8ZBAnXBTmSeX5
rXaKitOwZV2Ng9vHUfl+OUkyvPCGRQ21FpR8mcUg5G4npLZ5lIcmTryiQ6r8FCY8ypw9z0+1XElI
YhQoXvsaQ2GJqsZOpFNkUkbZj/SBDY/UZeGnPVBHrNeFausXuuTgw+nHdfguMedv/RlXvljYJuEr
+QLKPPKq/RtIzBlFlInNfIHXwaYsIdGb2O+RU9RwkM7Bdhm5uBmhBx6NRznDnnx/fEw7mOvL8azr
kK527xT1xOjPjHneQCF4miZBkXOIHo6U6/WThLppro+Br5qBN6jabxt4EtOKCkHf15nGdd5/KW/o
1wApFFVuXrc6SXAY8b8Gx/TSsJ5dV5xsOf3Y7/N6YyJp69RL5oh3z6ulQyJJORcEN8uMex47EfXp
8oZqnx/QiVW41w/SYN5nQPjaDEHrA1mnayQnx6W0dA2xrFo9wBf6oFyJisqix1C2XBXSMmKgqHC2
r3bWFz3i0K5D5VqAhjQ+8zH6R01GWmXekCREDAR5pNAqaZYDgOZxRAQ0CPftKtP0Fjh28G28kgSw
WJ1PUpwj4UakmFWwtmo7R+lhjc3qm4PRzbXvP8KtPSQrs4RGZTsTJTnHQQ1IupN3cXQee6ZCNDhI
KdUYEYKCbVHGUkP62mXbRb+XYEz+ByUHa3rEXwIPlLHkb9C/JvCHZ0CbHKcGWR0rTDThOjyye0eM
J8DghUuOlg52B3nk3rDaS2Ij1tP7bZ7W4IECDQTA9IP7tvUTvCp0qLK2X2jevsSZr0yHzlbB2uoG
EdisJ+ej1DJfdoQkFJH/FYyGx56R+HoZt8Xq8aI6anafXPlpm0NfTSMgsnvdHm9bxb9WcpHDV+Lq
UwOCp8EMzMTXh6YdrLpoWX3Z52LjdWGgswsRbh7JSe5bFUWopObguNWDQsIErjKvFfDSASyLhT2d
GuajVOOxDSRd0r+WU6d+H8qaxCeFh0QnMRscxMIohzRcDy2d4BAFmG8RGr48e5loVGKUMpCSOPr0
NOMIlV7ecbZPvHTy3zPvcuu433810J4RZfb4hoAda+hsZziI5l49mDAzgXKO3zZBTW+VBG7sFbzP
qnKHrgXZ0Z4Ben6MiQnpq2Ty5XRE2RuV5m9+T9phKEK2brKwWLFz9Ru7fv5pI+mg6Ca8ORwc0XEf
eviJ6RZ44jJVPNMVSGSCQDO/7JZmKHVTYD7fV3eY9c2GodyNzdKlnakE4IYp9BFCFeS2Ea5pDKmz
wwS9BxH4Iu4kePTckk7nkW3wEk3wiJFC9YBEvkytVxpa8bWUeAfrsuR9TFPXgj3LPuIACIYms3UD
uaEy9tWBlISKLcopViFzYrk2UbZW7Bp3VTj7zyIQt6AU4XOCmquq4cSGbJtUIx2LwtsRW7GFTHcZ
kvmTtR4BT+o+I9Ou6x/9dhrbc4xslGwgqhbtnKjZvqBRVtkGhJ9AsVmSmjMzNulYQdhaeOqdpuvX
OvGMMapZk0MvaZYx+rU2FD18bPZdMnygX5aYvyDelctS09O1vfNt6vWs5t4szcCCKZWKB2MnOAl/
CBOmhdIZcwAgSdw9hEk+OU2prDpiQxsd+80ksLiUvQokOr33tKO2BTq8Yikg9gdsWF2fMJGmR1fU
L4f2+5XYYPaPm7cMz/VxkAH9vzwdvpmsmfE8tsmCXmYq/dmzz5fp8mRP2XvIAnupRt8wJxrPZmtj
XCR1zivpQCQZPeOMqwCeSi2K6UZI2jkk3JZ1Yu5j+6o68b2bmuw3RJ9uFWtvowN552OgitlgT6Nr
q28LYnqod4rcDhXmWwjYmq7I72p3OogtKGqjD4vgZ5gEy71wJV+LNXGnX45ju+LPDw2WgXAqZvxS
tbSRSWdBfXU4QF0CeCDc+MvShK2JNRcZds9xuQxKE44KhuJu2sUWB4L9jAAFzZYpHepE+5TAfOsV
JnaEKul5Rqct5JLOKtUNoS/+wGKFSE1/sQZ+v7L/MqANfMQKdcbhqT2F5/Jrs0uH39yNg3WT44cN
ipSLb1QciLdYR8uzHknWoX7Iz+Sk6zSclxm76Mqe9JlunSpA0FSYW68wZY/tyR5ZbeVG1K06Zkfb
JuROrFTr7qD6b3e6st8tx42vbSjugB8LrblN+imxqveYsoNEXk9mhHtQjYT41/ARi8tj1WF9rX2W
ECakc6xQ5k3koDLxrbzdM2GVApV/aa/SD0nSA0lg16VYsAoTBrhQgDIyKYGUoIkDCveynrEgDBWp
U54E91j8i8OQxlpxgGmOnXMTA16M1zsQWSWPsTIk2aerzuiC5yKVEl/CQBHVGNG+OaNYCO/eQSRW
zhHMiobBPOR441MAsWrkI2P7a7F4VSVAzlmBXCynm+tPxtHJLYVfmJQF8evnfUujpRJdUP5euJOm
Cqe1onTGlNpQuqWEPmUgAixfB8zpqbA8IKt9cuWRYC/vH6NlXGGOkm7MWjPlNhX+vFpFOjLpdt0+
TZWaL/PFgqCwXzt/g19046fA0UnRbYFWP2MQCt+4IFI+KFUpAjhLL4pdMqnPZ+DFf8C2MoBT4tUw
CBmf1XGEbibEy/BCJuQzryvp4xqXK/EQhcJIsPXf8xja5KSyI8j9zyTZWHE1aViLjMYtyUGtCjfH
RsMWy2wy0XuBd6tPzvnZFYrKUdtnUJB58slwKErMZpN+CCUYms4AAMvc1m07dvU79wyDhPlrtkwF
x9uoERK9bLmSP6KagoZk1zm+OcE3c2qsmrjZfJc6uPuFWZYImTvbnsA3Gr5jB0Fp7Qd2NzeCDhvo
4iM/rlZJ5q3UQ0dmkqtTlJpt6nxsrHywPAcw1fAYwcQL3Hl+BJYiOZa6tfo=
`pragma protect end_protected

// 
