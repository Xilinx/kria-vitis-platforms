/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dD6sJjMckNM/hk590wWgo7QyLBP7qvuv1GnV/mfQB0w/i/pvS4BJcnppdBuizaQbHZTE85H6pboO
mTjEC8kS1yUyaRKX4KpOmRsaXVL7/iV6Mc+EyHoad/3cx2lAwTCRu6nptqi96Q/dtiPbQirlE0cr
bj2VslWvQXYp7agPImHpkldpbIx4OKKY49/lmZgzjQmz1uAl0Vpqn03TZsorFhKrWNa1NL2PWEvy
H6r6Q2NnxwJibsxIu7/DaDQZ9tx7P3Ox5rT/+t7OV/sWKJMNsqkendhSkyxMCR6Z1Ip9YxyEItGS
Bld1ucslP9zp60t9CzMGZcj/WZZ+ve1NzjV/uw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="NlHs8opBWv2KH1hFnLsdY2EH/Cy8LVzvJ0P9w8zUaYI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 880)
`pragma protect data_block
jOrE4515xgbASXSOIDgmJo0c8SZbBjVFRDwRcDqfwrXwP+X4O+KaIFDjVnzqixqB4+NQvRrsuEmM
3BrgcJ0atT95TM2iMx2RlpUwRuPcQ8Hd6CHKHPhmu3KuBjccJW4D1qUjw0LYD1htrvzXUnTPDQcI
yjjFa7stZeKqe/GBYQOeugyDMHvQZHUR0lhAHeRSt1c1Jg0ZO/gOETGQhlziIXRqBzTdWmyLVro3
j3k8aw5du19u31olCC1dm5NypNVYhrxPU1JkyAi2ikA9Kf7rpMnII+c19ufn2U0sPXkE1o+XICxr
oOaf0OSFGeTdeR07Ymf4m8bQec0vtNv+UCosOeO5Gof1XvUXlkKVL9BQb9ua3awmSOST5hTjyyZT
ZSBTVvxsZwLyb3f4O3z+Wk4vzrVUPNd1buRRVGcXD5LBzxtZJVwJKKhGCi/AJSa0grxodMFmHok/
fok1uCSuQCuJjgmHvkz0QrOakSM5uyv7v6nGaYkbAuqy8RWMehdA2O6yKzjS2+8E6oeDHP/3Eajm
z4ryzx0khr2w0VUnvvHXhqZDSUy0oXIVxkJ4vpTcOxuwJrLPQMZ22RlFOUFRcmB08hIVQ7C5x2wL
c0kmdRioe1R/0plMR8tSv1pmK1sG3cyuvWvhdOv5WZ6KHLAIF23WSYTLsBms80k79azM4Gw9l1OZ
MSqSwtU5zIOBZKr2PMOWNwAR9rxp+jaKn57oiolGcDqPfpo3xkn9wIocxYW8QJOJdfrdCGUC0xxY
MrgCW19jPQhplB6v1KykBRjjhCzh8BZ3dBEwDjOZaI8NiDMYh7xtjFUIJBqRPElsXprz1wyyi9jU
UGY3DrvTetUAhFIPlLLb9li99KhVup2ceNR2Ev0DYdbNZ8hkdjW81U+6DqZfCRmF0r+erQJXIFvV
nStBy7DfF5/vPwJ3gCGbhTazunBVcPhdsva8rYSb+CrFCKGBCQBG/c5/h3UUtfGcMGy4HfQivHD0
LjMnVAfQyUQ4MHR5ESoop2eYVsjTu7FTCI636JfKg8FqRXvFBV+pza+JTqYqO5hUkK9MXY5ZsruU
am0YGiXqHgKhnoMoCJ1N2OjMu+SVbpLm4S1AcdCIFKKhIYv31BOWUNOhWOXi1gSxCtSQJtSuF5Rf
eEO2cKb3NBDPHtlBmwVCKYW93WZStkEslg==
`pragma protect end_protected

// 
