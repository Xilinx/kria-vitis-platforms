/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
CaihNQWwu+qKJWjcmdIgzgKIXQ8l3vMImmWHnChjYqoa51yMcErBScyiE64YZSDih9WCUqsVfjEZ
HfdPZ9ljuyASaDAJWOBnJBbhrePBDPO5jKkFmPbv80QoBXSWaNMFc5sW0Ulg3lCiE5qq9SVr7IMd
vkFVewJkI9IJKPXIqEiYLMio527A7EkzJrjUXC11BQnTYghbA5n7/6q2WIDOwjQ+BdLZXxGdIUKi
ihIieqBZEgdd6vwETSGv3sSorIwnUPSueC94L800xEEoFQmghwgPGvLA3IEIqt1YNZfrY4rcuvTH
rxE5ve/ar6tMYP0QdSitAf/UOVre3EWtsP+Jcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="IxINXwVvXQ/n7KwTaYrPoEaEACBK27oPy3cRIdl/LOI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3696)
`pragma protect data_block
EiGu1ShDtOnFp1/lwt6Vhfsr9gFnEckKnswcEbLLSwr/iD5ZxXbGXzMqMrbRcIl1KhEa0QkQHY5S
A2RDc1xzHxQEDjuJ0miDGzuUabWBhHTQfh2QgP1ybq+SSibsaey/C7p5fGQHilHwaPoRTIN/bPnO
82yPdqTjx4lWKyr6Int9yGjPsA39B/8FKpxLkHNaaxmdknzSw+bgK/L8d22eWH+342T6D1XM8kkr
Y0sWWqxUfOmclElhHR13NfFSCP0KNK0OBuaj8G36aJq6g0g89NpWJS12EPPQDj4lDq/C62Xb42uN
6sCNiopBnPzzN1am8dOtZSv6y9PKkNivRkvOy5qtJkEw2HZzrSTmNWLXG233CcksD/YfmgPdzhac
ywUVs0OmUo6HaxxWgViRr6iwPUdXAe+4Xl1+Pc3CD2iwmHJvhSWi3egYurGiwzQDYM6uYOgJ+Pki
pv8L7iudRbQs/2tu+moPD5xjqcqNNNGbvD9tZo1Ix7vQytPySN+A9wno1rjsDpUbOJmJk6zdlfY9
Gm7ec2hSjZalkPGcwFy+ngv5D41ouz9aUBU3Vq9DzSDclvBXqJG75d2hgR+Ah9MRKY7pz0lLXhHy
h3sVKdrj/5LLVV+zx8QPXHDbaEJrYcOpW2NBp3LcOT9AYqRe8nsdzXPU8r0eE53+YarB7Wqxyh+h
xt8yu4U0aOXU81991lyGCK//Y2UFnCGz+1o/WZ9ZgVkczOqRadzxbWz5bIerIDtLvsqbNwgFxmWa
qRk/eqZ23EOnKIRBK/vcQWdRo9zxJpkv51njZOB+RNNJLOlzTdRjzofWIr6FXFn7E+mC0nsL5g4R
OvsMdTCPeyBntDO79Re7xNAR1Tmcqs45szObE/ji5eIogvrIYLU4sQwExapnEaw5EQhdHM9eFgsy
n5XjqU79SK9zfJWWyrKwzNBcW1vhDu5cNjaTM4JDk/PrfKLSV7K+ihfqSXsyHnkbjM89xFDkiOTa
x60SzItwVYeiPdKNW0vJ7c+1oEp0pVtJtbIuxbjVlDSfLCe6JHKc/s8QeDIF799tM86DGmdAp7yU
eTkXVCOkLysDspoNlsxEa05MpfeokUlTNjQmIIHh3+8vjKbtmm2z6/i9A5beEBfPvWgvnF0c5znZ
Ig4G+XzvyeXDavARspOpdj/bkorTA0Glma66dJYGul0wgimxzRwQMdUDrHLC0Sxto25YbYWHyadO
IR4hT6J1XB5BMl0wepRu5yqBvK77SxXClOsnO7XR+sGJQczVcKBntfBQbyu0z07PiHhMKECjYC33
7PkxNtovM9nUsVEEKybm0tnFWlXX3SmkuctnyxdkGA83kHZhk2N9+PLkTq8ySD7PssuurKJf3ODE
5Gk7eOHf8qgOuNKgzA7teLVMBdiwjsm7fTsdJ6jjjV2Sa3rrBV4cvtPA6F5Z/HWIOQomJKN+Fasq
86/NijWhU6us6zGCHKa/gcnBcMc12E5VZoJn/rhujbB9JNGedr25VXrrFU+ro/vVqmAMHDPQZO7z
P/EkjlVd+oNUTgNr6LoJLUze+7BPnZkYJjkj8FMQzqUu8ehevf1dw0zAbNvViTB09K8i1pyVWPWI
Vs0Fh12s0XWiopwoxO0iZJbEDc3XMeEgJPG/txOEcBcJ3l0kTmgk5QVbCxCO469ndPvCI0i0qk3W
ZOjBiSO8vyB3dpCPuAq4u2uDuPZPfFJSCL5xGjXkBE1M0CWQRvt1pfIRonxSvsDxpYNkRr5IjCBB
ljFlrS4Qqz1skRQAoE4zNOi5J/DaC6CeEiGDTRTcr9hkUGv2wxqtcHl/ykT38bRjV4ACZ0SApI0L
5I0AFYXNVy/HyDoq7bNP+Kn1k1myWeoMHrX+oebbPR2IDicF7RtkLjvocf6TlmtOOpYukyNd4rzS
qQXZFTvubLPMuWELsXT7kplux7DapZ1dzSQS8BqIwR379ho8nKrgcHsf5LiPIYj96Bh5Fmp5wj27
Qnk4+xlIzdRhKXITSEXmX6kR9c61VZxVEYatgEGmhvaqOKxme9vRPmHCjGhGqwwZkRz3aB33AuL/
Q+v7WZhLtWvnbxvRCFHtbJFYARw+m8hwhB5HmyHkq9po6fnLVSEplMBddiqtEOZq1cpr1BsRcyYz
9fIhcIXBMzYBB5VFLQdbcosUYWLGorncHTTc77916jED/9hnFFVd8g14+AzqqLmQYb8PcgMysK8p
8iJd0u8L6PrKMdXNY5kG7vGl8dNQfVwAhwFpN5Y5bBM93/Hio5MkQ3HLU0QiqxYlSolmN3/Od9AG
V+0Ty+zIdKtewdYzTUDPXNCB7mV9NtEUCXaKmNLzp1cZ1l+cHnyB2DYFVaiONygAQV8nkKggFZU3
trJhTg+gDMA8h3An35IpOX4xl6235PzFzXPNz+6Hb42BRdKwSeb0yixwl4tpSJ/WJ34A2gEcB0Ow
0v8j6bqGUNu0e4mcPbMqQ+w+IIVIDO6Cn4c0fVqEEo5iVEZ6zxiWxIWLEqD8Mk0ADWg2UmodDjlA
za3iJYHS4IaA0kj2bjQxIJa2wCdDJAsO6j+D3WPOXqy8WUggDFrwYnbiKX20Lsu7fG9Jt3uf1Wi3
bgLXsssYqCTjGFaIwAA0G7NhRq22fO815yH3x/yVLMZFkr5zqk+axJ88p/VmfuKn8U5z9YxNKo2+
kdX+UBFjwKWYUPNqlDMSroc1U61B3gnV8eKcXAKrRc55eNc9c1ed16sjZMdwhM1s6vZqwsaDf2Tt
NKiZOI/qSYSjxFAKNQy/Wvfo1wpnErhBdEYiwMgfO9CETQ7CI9Iv9qmXMo2fPbPS7lO929WFetUs
9+CrR4cIfciRePvw1EdmAkQ+JP6iKrbo7+KBfR3Cu2JTJpuddL+jkQ53s8asAjcx6L8jvG+mJ8/D
t/3W0fnHkrNRerP6OUnXu+xda9vIlOF4a2u99j6ArShcT4sMRk7jVnLC+hHeUpIcDj3sLYlIq4NS
Py0HmHc87HTEYEC1BXU/JFd4uf8Y2V7WBJthxu8C9l6kH+qx3aD0cYdXJC+dAG//cQ7+Y5nNzX6j
YoHIuS7pdSDA+QupcWrXLpGkoImwDnttZJTkqHlGHXlar5zw9QO2bxC9B3KYQHHxVzid1rs4YuS5
Z38J1kE5MkdyIHy+NW4vqixMWJV9lrT1ldhfYGtNPpM82LmTjcX5/jM69NfOL7OZzig04dQJbjgt
3q3OxMS9ANFdHBzsflpgll6qJwHcyl4jVdXaNbExM++U1FjamP/Xz+9Vi55YxQWbft2+qjcTfvrz
qHt8DMVnzBGTF6Oo/yvvLYKNFoyQ3Dp47dYeMSNCM8JLeNT0QdHFEz4GciOdkgaM+irZpdEDAwFI
+4yJ7wcJ5mWNfhVnVEMDnY2MbDcPbFPShjAK0PEcFepV5ndu987Xnl5fwy/CmSX+nycK1RoDP+5D
BQqdIdEyIe/WKTThKaWRBRW8LjUDfWvM42lOlBg8dT+gfnveXH7+uPVUq4baMp0HR14QL/Y9cjhz
7klVUftYK0ZX+Q8af+IR03K5inpFTGQx+3VEpR20G3bPH9lfi3IPf1/no0OjpX5xUqDmRs0R3Csj
QUfHYISDAFP1Ie5bo5BUVROCBPy9sNAs1zkION5Vi7Q4oCe2UNo20KIPDcpqhZtNExksj1I13BBn
hP4qTAPSva0P+/YsC+M+whEeT6Q+NgpMuETwzZyDFRPTv6KV4nVCZGXjwNWBytYQt7i97lfSAPh8
YocwYrC+vLcSqev7pVRFrFW/otmgCEVOtvP9ueRYKF8Rp4JVTFHehJqvPb+QbWNbrwrsQ9CDVyM/
Bmoqskx4R2bWTjV8ko+xiiTvWn3xoMOoWc4QfLKhT5P3aMLms8Xd08+Q8IKEfsl1KH/XWTZMf2rD
FQ1roNZvL5Xj+Ls1Qu+OkSpDJ6Vd6IMi7vAYv5O77CfT9BqbZsNlT39E8omhgFVWUaFvw4Qu4rNU
8GJPFRV6L/w76CgUCtVeuacrkjTgtoa79GDVcY2RfxE+kmCEynSagqylUSBorMJvKINMkCuZeF2y
XNCbSEJxM2nitvBWNCIv95Qc1DkxblraUJjB2UoyLABz1kBBMr1zOT3D7xHK8iNFqfE/pbwyHFC3
fWXvfyPYdGjaTdPRwgCbNbOclW4bHL7koEy0WJ0ZpRPtsGjyKT1UdubEueOVCesZ+4jxrT2zkqZs
mG/qoTCD0pl0/pZXJLQu87nVT2lTOqgIiit/TmZ8fAmN72fEvCjyXnPNhNVwWmM5DLaI2P9VK1/6
SwZJO6X+dDu/C+zZ2N/dTozjajSHh5gJOdq6qCvOw8i2vAhNEiioQhxomKd+vHyD36Rl7HwNIYA/
Wwl4Bsk7/9Kuz6/MNKadEeIo18ucTeSGEupb+Z4DKHTT0AVTGrlwrxp9S7JsftKi29oNs4FbmPiJ
SXzewZ1L8erqlAieG8wGPEMIrWF5D8v3xs8Ed0VMhESaY/Lme0nF1cokJs1sjuZCfMMNLaIrtP7L
gIlyb3sQfwGl7CEriSsYwpYtU+45tlsSRuVHxcv6VbJu5QdEuxJY+i0/VI1ph0/03VRiunlFqUFl
DwiSglFQVaUaiTZnLxh/vE2E4GM8DljwJdrvsSSgDq3ZPto//2kcqDQRmte5O+FU5AXhBV4m/UdH
9l7Xla4zlzidb4uni8/4OIsN0t03kMYTTQbSzHviK6H8U2nX9D0/tAflpG2ZunnXrccBiqPXngDT
G4eKNM5McYejDQI162GwAw/Vj97lbhLr/13Ei5qXEitATflT9lQJzvzDD8/5+0NptjOYroTCi5O5
1q4GOGbX85FkprsjgsRGnGWz/IT1xfc2PLi7WgIPZJi5H/uuCbmhD45INAT9yen7QrPZOI5GZrCW
Q60NnhyUzTIXNd6v6tlPbX+oQTu8wFhBnC2pOLNpyHvlHarGQtweQnH20ndwku/A
`pragma protect end_protected

// 
