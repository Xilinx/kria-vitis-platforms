/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dD6sJjMckNM/hk590wWgo7QyLBP7qvuv1GnV/mfQB0w/i/pvS4BJcnppdBuizaQbHZTE85H6pboO
mTjEC8kS1yUyaRKX4KpOmRsaXVL7/iV6Mc+EyHoad/3cx2lAwTCRu6nptqi96Q/dtiPbQirlE0cr
bj2VslWvQXYp7agPImHpkldpbIx4OKKY49/lmZgzjQmz1uAl0Vpqn03TZsorFhKrWNa1NL2PWEvy
H6r6Q2NnxwJibsxIu7/DaDQZ9tx7P3Ox5rT/+t7OV/sWKJMNsqkendhSkyxMCR6Z1Ip9YxyEItGS
Bld1ucslP9zp60t9CzMGZcj/WZZ+ve1NzjV/uw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="NlHs8opBWv2KH1hFnLsdY2EH/Cy8LVzvJ0P9w8zUaYI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1219024)
`pragma protect data_block
jOrE4515xgbASXSOIDgmJivH1BrgF1rw+6BJcQoBitrI+HvZq9gDrwocA86EquicOM5HsSBkzDZx
5BEJUjoBsfta2i4Bv8REqJYjs0A5nuVeRVtaD1ee8Qp+gKufqTZf3FNUI4d4palWbc/9+fF+Ok/F
cuHgim3m000SYp18ErFZOyZRUUg5X2brii3ZBagFgMRJaAbRtMjpsjjprJ5H10LBzgHjj6ElO+xL
TVI56cJmxdH/XyMTub4H2zPDcgeqNNvCkzfpj0LKgYzr3Fzznz2Igmfhmt72wRYhUoWtUMzkDiws
n/TaWHohzRRpOisFCmxo1ACvO67DkWEgR4ZrMwrmn+gCC1YQFAdTrh5yHthDeomcLUGqyD9SZwdp
0Ya4A5MSrxUHlBnhgIuhNjbGItepyKiWfbWfP0dv9TA86VvLu6DFfaGazlexRN+DfGEZxM1Q2MFs
Mcl+iU95bQTfyWBH3eO1YSSBFHMhhzoYdYY6twOEdwmnBo02gkkAeGULUJFZQgz8ykgx0Zhyvedp
8NdkJhc0izyvlCwdEn8Qzp8DXGsT8PDh28YBOahQbnKHNO/NY5/EW1NnoJzrqWW78lkTi5mzcZVn
9+Aqvv0DD4W7WYrAftHg0MVqJ40vrH0TOmQHYr4TNiVSOGWQP9ph4MvK03YzGhj/lvElPxK0diUp
iSOoaAY2WWyB3KYK282WS0Xs4dj96dOhOjuo4BIDxIA1ccmh3p1jfj3RKloPmQeIbNGUat6PqLzJ
C9GuSZOWoLKJ8A0ABuEzgeJX+Rvlaphd220pypU7KAhzy9A7JYgsEvdGYhqcBZgARQBLCUChqCQL
ZjQKkLZoSkES3rlHbac3Q6jro2V6FYSBUTgpwaSts4RLYbbs2tTPYQz/YzwEIEU/1pFSYPEKCeLO
rcaaAOrqMdBMPYfnHGxyP81itwQNHZeTmwYSa4ms7rrjjhxOH9fa/kHwIaE5xUPXtLscPrfTtDmI
IPE5Czi3tV6vQnqmhniZCh1Uu/3aozRbzUDru2X18GOYNe3OzVFwsUuFdo2HZ8tB9j+Eik+UmN9y
JZOZBfwM1PgRJZgBnBxVOXqTSkP0TtMHyCvArngyZze23LaysKdhaQQnWaNAOFfG8Z9QucZVUuT9
Eh3rNUGfFak9yAe7W/mQ3ME5B9WbtcRqe9J+WNeDhMuhGX1RP/wlyoMfhiyQXbLZ2CVq3DxeQ8Fc
69CqjwS8FhBBoIt+47iCodbdve2TkneZk7G2/4mOVydqfULHar/Xh163I1nVRdIt6e27XOIBfFBC
duVUq3INvZLS6KUVm+CZRhQln4gIS8+nlIQ20QGSv+wY3VYNXP66Ywlt2uUGlBTIKAkszY/il4I9
Q/+m77oBjW9Hd4IdMKIXq9tuL41EBbUwUO6lPpnQ+wRrZz5Z0+F9hQL8zmYjD92PcZpXENsY2pGm
QSWKIvMyBZ4e+n99PjNgKvXpzLtr1wEoYzWKNsKCXDa3qokMARP8UERranbGQKMScOW3E8T5wnTW
ygaOuEGG0TLPyjwezu1VQT6AJB5SNn38k2hnLNMlbbY4o5BYiGK+VDdzaJgcuETJ7LpjBh4G4nPV
CLpKKtS+PjnsJsHsUbz8pS+152EjW7oLr5/v43kXwg0R/1BqMEX5z+dZ10STwTr559X4x3tb5xVE
UUSXMi0fIgqKGkrE3NM9H/BH+vsB80PXresoblBMKI3ykGAZ0jckLd81QkwCCgXGyTeAmhlgQnrS
HqaXe1sN/6WGQrxItpYJZ5Ig3DXCOSn5pgplFol3ktRMwa0IqSWucyFn5nhuh8jufYxJaUkbehTL
yqWL7jX9/vtHoDjTRIQfZsjeqq0pyvjgKezQuxiv6CLoyzpes3hRZPq+qPSESV6JRS5GOdyYV/yY
Wv633YvHA3Y6kPLtDN4cHAiUOP6TjHybZmBRwkh/1o6x2sW+ZkaFIuwgeGZmyhzn14/wHYl6fyCm
NYjYYFbmzzfo6w/yRX8PBnJudPL+pkzoGkYcg3CL+2KovvOMqtfJs0UwjDjE1S3bf/W0NINaTzDZ
aA8eRl3U62Y89YqZeTv0e0d8xreDjAGZEA2iBTU7Z65674Civyw1Xl6lfMW5+GSk4B8d72yXcSHo
TGY6FUj5wRY025I+Ak27oou0BR+Df+Hi5RMfRkK/CvopUuRCfK52Wz82rub8NQxyaJ7j9u6LPlKL
i57f3fx8Xwc74Ta9YjfKghDb4sowm+eZQpmdOUoB02GGCXuxSm1uQkHcKpASBBZ2P1SVF3LcsA/y
pEiT5fTbwQAoYJgrnq9flIeMxskp6EEh4XfVxHoJu8onL/FgL9bIL+FtYLTmfwZ3rQtlOIQ/2nUP
G0xkQWklxxbtQKVnCIZs44+6K3sHqx8Z9czkdbaRuvzWWYGvu35pR9IeWvTQl2noaa7w116ViZMI
RF2GYjPgS7ArQ3o/jHMPi9bNTF1d25zARI5C/z3Ju02z166VQESIvFwOeuhkca7K1ZwSphOjq4p1
Wd5W59aUDoaEcmRPSVJNgWCLKAM32esLQ9fu7k+tjV9FQTEOtT9KkIojsyjG+LTGy+1Jq8pw6sbC
yay6CS5Sc0oHIXr5bKFtmCbExTHpEWCCTQY1xUY+L1yZ8GWW1yomSHufEYxd09J/K9sQ9tnC/EGV
rH9rLfF2UuQvpI1EijAQfp6uwBFKf7Ig5uFN7zba8N5QHI2FLH7InlOsNfc3+yOkKT7gliOtmlV0
j8hrLLEh0XbE9DkVtIZ0sbYJ7Bm8emJazQT4m3cRwgaSk0w7ShMwlnN3jAmv2ggGppyyGK244XiT
KEOGE9xkrMO67DEvl44/SscI3d6/7QU4Imr2l64rEtMQwu9PB8e8Xv3fdIpMAEBtW70S7LB+X2cD
TU1O+60cy+DzZwJZKN9J1B4rEMsv2grxf91cvJdQJNBWxT3dyq7TdAjUZ64VQQ4Hc6Jc6CPb2Tzn
5f1FNBkaTu0/scG3A+8Lu0L8fCzISI/6ubtiXX+HjDCtIXSaAQ1BGehedSvesK+zRWRia8owFZxb
tUcy65fVW/AmuCYdL671v/EGbgMQztW5zvuIUhZJrBQAHnyUuU5JeKIQhFQy+FGQ5P0HE469nan3
QDJA2vC2Gm0KF/YylO8ADkSeh0MKnsHoPGjiVCqtD0UxxnDkkZ7EoHs7GTbHQaECgXGtXoFwc+As
yllhMSzBrE7rMLu5EEGeIz/NQQQi9PChrLLJNLVbTyDXdgFE7a8fn5LLNBoyyLGNS8MVF3N6sIFk
hJQOyx/KN1zOuDLJU4xZH63bEMyf9LrOiAdyleqTYkGcQFSodTLpk8bGjIw1sU2M/miCEk+AUht2
+gCIzPKsVyuim78gJgfKktrEcFgLLlFZDLdQBSARLYKELhXb92hnfePEIITIT30fhQZdGlzocpyl
tYdboCvlH3dZcOzU3yybD3/nJ/PJ0NakEF2OM0eFf77uhVuC6vAjxWsHvhJhgeOxq7Wqyh3uwZXt
zQfoxu+CV74ElsSR5+iHWFW4KV3HBgoA/z+Ry1UlmJyR5f2UB3XXGU6w3XUpqr0uXqJwsFv31/mw
w25LUNH8aOXmUdLtmWtmfDm1jvnoTiaia8FWHO2d8K2k7saZBrvS7fB5p1EfbBZ39z2txFISTZ7C
yhz0OoMlEFfLaDuRZYJ3fmVyex/lHNj67CXdPvRZFKvi8adkmezY6d6VLIKvKjCA1FC9SahI8Ym+
AWGiUE+8CmXW6ATS7yN37CqApk28cxhFZoIwRRCk2RJge2Q3BJ6qcAFIW7k36z8vxrMNF0sQjY03
b8LMM5L+/WiC07fJyjH40nFqkXQaRD/crnCR8JwCqd4AQtRNKAyKQ+dXR7l4CgQ/6Jrw9ZOlxGW5
Znzo+RORJcW6saSdPRIXjniw5sokgKr7ObTWHP3dy/7iaqO4xt8Is1Uecg0Bd4kdmiK/CxjQn1ol
KpqlyJ1e8qAS4c62xyAnEGieiyZBAU48OFDxqOdkhkZi1QzHnD3iEuJfKEZ5y2rHudjpLZ05g3uR
OyvxvqSo0k3D9ddKgOeyF6ExlXKAj7qiI+aJsNZ0SQFjZbMXUx/szqZZNie8N/1aK7YLzmq/bzho
aOgJNQDJjSTvCbRH+I4gngrecShRMWuLZF54CmGuG7wPh9V+KUOnkzBJyvdS7SYLWwQjHzbeedow
fe0Aza5pFjTd5aHpQbqpRHOg9uhO7gPWqJEIP6UnMQfqbGkAbkACxh+Z0UUbkmmfAEsrnAIAFaOY
nd1dM6YZ6W3qEYOravN82Du4hb/amUDNMZlBExvnO+e5w1ImwajU6qSyLppx0gUaCW6U+MGHRkvq
MK5f73Mrph8s1W8sqc/007YynPjLvC2zT3fkXvaZU1IbO4pRQ3nzjQRJHWVWvlM6r12uJL/m5bwV
9xsXzumn0BRK3J4+D8OVOo2snMUPEzrmZ9IxglvM6yjqOpWoGKAEC0pnoYLOM3JQ67Zi2MvWq6jd
z4oRzhXC1zv3zjIEzibCmSeaGWLFiS68SUAySWlq6mnDIfqhqmT3MkGgRcgdQkECBTYGu6jhCPnT
qARH/i+g/OvIFwXhxPTALRHOeCpp9tNFZXoeReu7jUNgjnb8vilg+WDY31jnHqAkxAtK5OShNIfV
L1c0uPaaWqB485uB3X9ItZx3DYEdYYZnkA6VRg8s6JVDb6MAMUMhvLj8dpERp5hEETuW+AnVAWxp
7XdFwXkYTIsYaQG4G0RESH/9UScJXpkgPWe5gbkYd00/7+vOhujJMYTWO1yZ2SZHhoo0TnoYJQDP
QgFLBqxwvJiob0UoxAsdWeqKb2pa/DW9elkw5ATNzNq6diWafKrT4HjVFd3r+eHGIk8IXJAKPmu1
Xn1JICz8Om084PZPiCBu4Zl2SjVUlxlIplak7gKfWyeu3hVSb4lA6nz3BXuL+g+RH5xW6Klu/CqE
224JwrMfi6fiUUZ1HtEXI+2LuIcrIcIt1iy4ssLUtuX2bTgPP6zL7Dir5wkgQyf1stcPc6aeAO0C
02KfQoRVxa6/qtzA+qamKzQewPpqcK9YvtwX0pbIBrqfVVCy+l1EckwEv6O8CxqITxS8zctkIgOW
xmb4IxcLO3tRiKT3cU/qvM/jUOoNcpclttTKps4yInszPUT2VG0xg6YVfYrRJQ7tFD2/xx67PhhB
jXVrIdhbrR7sjIpgGQb+DGM+01E+jthVq9uFcG9kuGLPlGmTaFBDWTRWV2v958AQfiDYJmDGDvT1
CwqeE9RAxzezsyG+a2fkHH8ROWb5tHly57C0KJVQZLfAT/eUOp7z3ouLTnBQkFx1IT3ngrwU+edb
3Miv2Q118Qt9VaEQwb9n6GdYjPYShhXJt2e3Ct64seQCrFAKEtyQ9gQZjq0pKAb7dih8SZsqkwic
2KHVWm6JuDywxqHC6tJyyqwFuYzfmUkhpPuoA/5S2g9Yj5rMkkGRBQkWINWSZ5c4IQexbGqqOfZw
YR/H43m96smEpih9IeZQT4uSAsX33Du432sl9OPTFJ9IYhUsNHlzvMw/POBE8uYdaVhGpJsO9pWO
X/MrkdiVyT3r1xT/C2XhlIAOaxGveg3jS2ZxOXjuGxhScHHnnLwq6iJ6oqNs20+BUj0CPcgtTr3Q
1UKCCi8c6GErEEVARt0azIYKPct5zyYFxmEht1ite70hu8Rvsn8DPrziIFUvU0SFj32raOwCzV1E
GlcZtR5RfE7cfhhGSREmVQjC2Vt0CGhd1mELVTLnHTRSlDyOj0PRhs+dQazpDpfynkeaL4B+Ubl1
bzDtfb1EyVzkt/xtiYF7l5dUVGLMO+i7dZJoIB/QVBN/XGX/WmzkYwbvx1sOmfZaRxQ5qcYdXdYA
0D4uzS1eNHl5ATRc0MhhBqeak3CQAIi2egZwdVnRGZavM4AXwhoOzUse/dLzZfKCC9KW4jCwK4RN
ST8vcHTC/MJIO+6HKEDPn+65oXbZkdYkJMG+PCtUAKFYSs7vBeqzhrGNF9kjRck5vYsmhYjQ9LIS
L10teJCifbBG/WS9y8KO1ctSH7sApH+hLTacEWXUgeh8b1o64v7om/rotw7or7PM+EiR+A77HaSj
IqelO6O48gkQlp7PF0+jqiVX8n5qu52a2324BPkOnt8ta/U2tyJST28217rIWKNMnbM8keB7Qkg4
FC0H3NjTb/5ySLzDd4xoryrpJXe4E+idJi04rci3mlAxvhZSK/lLMVkhLnTZXU4Bcp0RsrHVIeBT
QtMC1q+/345dm6ef7fNr/Fvuv6dIHgS4OZuec6DHRMxBSgNVArnvU3rF6aV29A5Qc1FAe0JbMuVq
STgYca1yKry6OdFKtMOOq+9BoFpmdZ5QnebiXSm12X1GZJLALqBM2aFHpYuYYSe5GanHDlhbVIrz
lWwyWcSN3qtStajo1wGvN2vHl1rErl2zvQeOwI6dIR9DGniBpgZSXdT2pchzjFCqwsAMyFOIbSy4
uz2Nh8MOAfT7l6Vgn43EnD0QzslyswfR1ENs+DHJdWB/KX75KW9L4el+Mir6QD0/Vl9PRuerXT4Z
Yjzs8gRDwgbHFE04aNqJaKCoCZGp47X5nv98t16WiHHYgM/r1mfRtG6u4S7OB81ogvTjVmqEh4in
Ct8Ft1DlJj9Yhjoky4JFyMxnfEzatQL5VO/TBj2gsbMsS7zEoe+XPhWkW3EaC54Sl7IV5k/ytsNM
CyAKJ54IqiSpWoFAvaksmvm+j3JFBWHYKK35m6DpBfclg8pIZqe4BlSigLIfN2XpVjCkei9Fj6Fl
cGMHMIqs3fk8mwjhBNhtu/6EKA/gUzfuM4KommNrfRbJpbLS+LDjLyIOmsUSk25VTH6TtNlx20Ho
PCvoCLKtN1Vm4kzt+ss3pC19ppkUSJQZgKjYPzpaweiNa1XRFZQFYr8icqiqZtCMAwKZJlNjjwxL
XCqnR59VHxuoyO/uiNjv8Ze0kz8F1N3CWVhhhvp2jH41JwrrGAms185x48kO8y38haDRVYyJTljw
Ps5ivHVJwz1X5ioWMJLkU+qLDj/4KmBKfIrrCGtH+0C/rlKyUXF9qbyJKQujAKSb4xm6WJgy64FQ
wywxrOeum2FBoVLbIt0nAMep1JoYD876kPcubS/j9X6rG9xsOIVbQ90Bpn1c6yViqPv5NqtVPnfI
u+8vY5sUGWzf12q6Lwr54LZzC5/Q8pkXGHDb7DheMdvEiRVv0abA0aZPNCyn74/aXcBx2xky6Yjo
pskJYjW3Wqp92hDshaJenJli0MGviQ4b3yZ3c5l7qfLX8N2jzNS8Qpe1VUi0ncjjZElnPT1Dfe0x
EVJJqpeABS781rt7Djl9c2vefLKHGIhyqHRAgUTbwNFYxCl62Hi8yuaJCZ1TQEMNt/zqT21h4QtR
7cp52rL3FXX/miPTe2HATXkfZ0jQDpFu89d4UU8W6o7QbrOtHuMAlTyPnQMZW4M7YS5bZ43f0RUh
P3Tio0fwbZu8nJIDCrNaLkMGjYlYxLKOmLlF6TsCvWWCP+yZsot7IbDZ5/i4CdFHpsQn53KATp5G
zoQmc3DYEnnz78fRJ6m/Gx719OrK7gw4yqpcwoUHaiZBifAGgyKxmgL8QXAXSZJv99xWPIrFMX0s
Fm8BYh6fFs89ZNDleepONgHT92FdlMZsU2oZhY2ATeBZEpszQg1ulNteWIrYaJXUR59TvHh4GLkC
lGxuyx6Ch15JBO4QgY1xQfhyGJkcv47hnTC7lCOIrNm9i25DMBgB1loSVb6gYxoY0q6/DvY+ikmQ
KXhUE6TKYchQ42imrlAU+z56yTLU/7nD5Uc4Jn2+n8MvzJIQz7oNjDnnAwSkKAANtavdDhYwDTiD
6frpQyeGUGL2JAfGtgLAPi2+WF8Nn1X4tHrggJU4ACZ4IOWjafDDu/Q/qt6pNLKCJ/2mZ480m6Yq
xjFI6stM/mGH/qiIFrIIQc5TvoJx5gFuUWzDbu2qQdkwMYwheVZ0Y3RSvkvaWIoVxwg1YCf1YHSl
y14vhBa81V/K9+O21GaKDzCjw8rolt0cjpHppKdWgpL+rnNJsXW2pzOWXI2Y9VPUZ2fbUAvnVF4U
PQyNiPNUwAfDWyFFEKJbPQbXyJN5VOpj00jj+Ds/VnfDW3poNeQGqF0OOBHZQVYrabNxcx9ymErx
kTldNKoMHn/EHR/4QCEU4zHEvrDavD9UA8t12CbluJ9iKsKErNeXeVvYsp+LRKEZDhIFPisBEanZ
8FbCbuf8vtWmaFlqqL5ALRXCupl9ZW+OgI8pdtri6OzskhoUltdvbOcHtpVC/hzgWbTtecvaQvyA
PhKrtJDCHrpgnm/el/7QnkaCIHfLzRicjfYHPlq/4Jn0hU8NmILtFivMB6f2fDU/6W5TlP8AfAqO
FIn1cW6c41v+75myOyXth+1FR55IukUy7vGMCXiLyAyhwAvOYf3J5TkWpOvFTmkYcw/CPibEZcfC
Jnpsvftb040mgAen25d7lDLAc6PIbFaBbwME49av5zfMWRuzlwfYShLOlokfwNojVpfeT+6yn3+Z
BrnmEN0zhX46hK1Q5qp/PXC2LnqoHeuS0Dlyl5lm3ZlVd0EGqkVjPXYsUUKlK97C/TzI+mhZsSy/
KGNYT/RNyuPx987XwwWg7qhLCvwGJmBy+J363ERc/nbgiEEuC6DvnP5umwvlNuLBayqP/RRh8m5i
KQZcaLIR0bSgLlpTwK6hC8heEFtkvGS7eytK4yHRpV/P+S0Jal6k/6C/KCXqW2++4dnUV7al+wWB
/5SzKtYnwlSVbSHtSz3EP/fLV0ufBCN6t9+s9rqbiSAEQtkgenOpDRSKBUPw2qoSSwnbDLYzZCA0
T1IE3gu28vUZGQIVl3j4DwtkQTw4w3khSFsoI+jqwGuk1dCy8YJcDeKuJOQjPZDQJiAPo1S0mAZ6
xbQ8UoLMGsDC4wL8weeyT1wgfujdn5BmaQCOQoQ796GmUY5zMuNUpeC/77p7DHABiiGKmemWg/Ou
mnEtWnS8QQ4WbY7wz2HrPT2YaBfX4c/MWuHfegyqrJ49RkN5NP0zu8UQT1sgX0tNPvtsHdxQWh2R
UqtCWRip+DYveVm0r6TzelCdqbU8VhzdcoIBeO0SrrhdMwDq7IPK6+B1tAodNnwzhiugeEAPKZ7a
rPZFxNXTkcPKax+58pIQuIhUBHHYRQtsq0nel/afLz1PQoB6ZiwI+gAx0JQ8yKY1+y72LS+jl1Yj
c//FYvd8llu6NGTuktOdc/q3XrXQoS4qzxPptIZlqZJq8zBSHMKMciS+huUxsk3vMk9yy/lxJ4NR
4OnYfWu2iLj5M4FM320c7cvvdEPjyQE2X3fZqkfzd2eZCqt/9t0sD+O7ytUEo8xGqh0h+JEDSk9D
sqvYfUxrAdaUBEDN2Co0uFaLpzb52DEzY3CBUFuVDJ0JGzg/9RSGpOPN0cRPCizeOFrnvvAXtWb8
2fxSuLavKRyk3U1h8A/Sh+7tnk9vQTXi3m0HLtiiHO3shDLv9IWAlKrP8o5RXy3jnqQ47Z5TvWpC
cmo+TemL/5S2ob37dPZls6cTgtlYhg+4iOjov4Sdh8zTG9z6jmSt5NBx6nwYLV2O/9LcCOVg2hdd
6PRswc7H3d6Pyjc+hvauU/W7mUSf5o67Gxe9VLSFFqXp4aSptFwqv/CFRsEGQiTRXWWaaGk7HY3N
g+zSv0lKCrobqx7rWWc4ANR5kiMxQk7iOsgx3IQwHrsZX61FnlKnM2HN85tEEByAC0XM0Eiury3o
VoDvi3N+l8o7zO5Q9t9qzAJ76xrpKlbq7ofy/xVTsNehpIozo8eFhVdDLu7UglfJbAeuAtEdqt+x
9UODa9jlO3zxFMJ7HGhTlqC7mZWX3UvL3bhPuSrBj7YCzx2R6TRbSXbXl2SD6/SgK0+y2EbI9Kf8
kthz8r4nc+I8GhM1bp5T6UvbunUl+wcx0GVbXurL2O/tPvzmFRsOyV+XqrcFrWPp/qnP0eqD5KJP
9H/ZhISp52icqHeAjlYYOi3iwueikeVuKx9px5amROTHdErfPotr8JVnfJFqO05SHUyFZQKZtuYT
K7/BWiiU+7jyM92NjmNd8gfq+qWilsJbZb+9UDPe2cltcuO2t7np/zyOLXI90nuQKd+Ba9RY08r1
9CU8BR/oQcLS5CkeNvMKhVpATRPybF0XMn0+gAMdh8c7Xazw94yGNC/6OckFUlgjX/XpBXq/4WNX
vDKrsiW/pJEhmaFTsJ4Jp526yFNMuMTNiaN8+BlbiWIMpdGy9untBcKN2iFsdRuZoJsUQxUR+kLa
DYzKAE7HuBAdrwNfWlr9PcUOGY3XZKJBlgBfZshd0ocbpAclaQjk9+vIzfRPRP6U61AuOjzLAofl
xapRL3cw0Jr5XMniaWfqAQS3UwvgCrcNAebXz/6l51l4czp8wfhH5MEWBRCynTnbhANiXi9AzKNS
DltYrw0c+OveUuPKqkA+MhE/nM08+Qvtyu2UjbIBOX/f4wndxV2vBYUflRMTYGmBmjfujk8BRRB+
0PMldix5nOJ3NEHR+FE1H++/WV1CjV3s+o7j6qQfJVyRscEOuJNGt9kDQY4ZLqgZ3S1dVuhPWx+S
2EHtbg1E9SM+c9kDs9nKYV5GM5l40EwDtccUK2prpc4+cVF5dE/slrnggptShyD7QMGCpNvIhz5n
56ZxNYjdNhpQ1jIjRDIBfeJqZrJezcPjxAP9K/FgILNVbAhCEIG3ucZqk3z+gHpWnbwVNqooZlpv
Si7woLhqjRPdhZ2hLbwdj63Y+wmVEEKYcaiVucDwMH2Nb9xMhEHkPheKFKaNhLyqFOCxFDSQBatg
kwsTArnf7RKm8sAVQXrcliGXjSV4wtUhNtyOFPG6wkDcJa3ahJVZijQ1M5HZmlAakAu+AJkgCtWK
Rmc+yVlR/SgEAgprd3UWACQsOLHLAGO9fUhJlJFw5hsPV6xDM8uvbY8cNrhmoqbiNpDGp/iZSedV
f4U6FAUUMvRDKLHoDa/UTGoVfrVxpI0O+dbac0YHukisPTAYy14FzYc4UoG/pKiWGmlO+g0ZfssE
omDjIc6Sb/mLfwIf8ASyVpb2Qlyhd0Dn1ihxbSRL0hHfKzfoivpDCp6/7MCOu53owGKFDkGGM/cm
NvuCAQG2ObjKoQ4/yL7ohruteqHHAGnq33/cR6kRQOfJiIdmIdYuK+3buwIVY9q2uI9QPVNn8580
4EP1zZ1cpRRldYFRda2Q39B1XGZL+ZQkAvpZna4F43gRTpGHYM7UV7PHrtr9rjLPQ6LhVv6en71y
TQkOw/xj3pXUEZytEYYZ+dqkE32RtGWGOVqdXRkgMyP8mNpCdozXM0PNfO+53gEgBHiQdnUx43G/
3ZFtCCrWGGu4vMSctVKjOvSXe+P8czdwLh3ZBxftyLnjrzG4Pwq8sR55Ulv2C30aGE6cwFN2wm+O
GmGQc7rmv8gBLA+ctXU7eUgLlA8oKSUowp/m3X1+BJJiR92vkpTkBNuuDJL6PlPsRyGTbhWA4CcK
pvutvJMcDv0YAPDCa7qWj4OHGq3LwxzMF8LXV137Z4SeHyK0weZkS8HokeMg9YgHxFq9Ae7ka13V
i6TVUK9RS+i4iLkJfxYdhoh+m5RZDS3McdFiU1uI1kRIuddA9tJx9AA5bf2TLIheZ9cXmtfw29Bu
clQGWaIXapzuBNhRbpnC1kaWVQcxAOyrOjild5pZQbbsMcej2uaOQxHbfrxoJg4fgMHH1lml+Ecx
eUsWrE1qoJY0sEFnDCcJWE7szpAB49TZkxeSq2+MJSTP+4cUUh74CoYHEC1cD6sI/PjGri/lz/qw
9aIS3lsfH79pTZtsVeqjaJ7tLOplERHB9YkGLqN9SQga36mIJD67mhPDXvAuz/Cz8PYTuActSIKq
kBs4F2tKZx4gazqk65D+IaVcHTnUVJmm+d2d412ln5gJW4wKUwJ4s93lbR9H/nkJ4CMV5XelqSjz
lBKiHs1GjqRyhKwzb99VVyCVUSXGdyKRWn/4Ixx5B8ObbaaAYPoSaLKQPZ8L39DMbU3Vtz0TZ8c9
nNAXdDsD/UFYpNqJ2L13A6GoxpE4TltuaHcuKt1gpX1czQSPHYB0+zFWflrvSr/l6n3NH0aVjaf+
en29fyvKH8M2Ir08dRaiucWMtWZBniQ6V5cFgsMwLDQLLNt57MRFYBzb+mpTO9h0JZ3AzNTi+qMN
1sxxQidzKE2YzwTM47BfOxONh4bk02dM5SURS8SiDL9A458J/HghtBfDNpf6M+sSKO5jsSDlip3n
PP4B+8h6baA1vJcesedaqq0Sa9yf7KuEApph1GO8O98SZ9vJywoP7WcosNI3hGo1mwr+o7dArJjP
tmU8K+S8rdVRzbHN6Z9vrNkM2ZyvgOXYY0dhYYWAg88Icalr0vl66dRGvrhIY0TvIv+ja1L0Gc1O
K4T0pL4hKTEioEQbnCMAUE+k2sllA2nhNPcDeD9yonhYTcG4d7urX16A1EID5bbmuWHcgdidbBeC
ii/yectOZxfae+dAtUmwgiERnrcR4rjYdZGv1b5/xB0UCvKyGPKMOXn1nyv7qdUbOsFD6oKuPnJX
tq4zXlu2mUwupcW73SO96Jukx1SUFFT2Rr5exNtr3VMj43tYJpEvqAM92fYNPlupz4OubUngvNlv
jZ0jseFyuZfgQUFSSPNnMnMtQJg9YTvo+bKGqL+zm1XpZRnt1h3tn0L/lthl4VTNm4dJFUCRjDsU
nOG4Q2TZ3XAHj3GI9iihgzqplg6hRLHV/v1yjTA02gnpKUl/hbm0NjNsO8EaI8VeGSr/yB4CcZ8i
fEj8qJXHa//FM+PHfVuTZujaYQXzU4V2t6E69X2WB/7a0wq3ZlJ3YKmF2mOjUTORIaNkYVu/2YRC
lQ4bEiFdkAbw3pgOjsf5Tlk+JBk1ET1HtJEWqhWyPM53LAIrX7mBVtEVv9GEfV6aKTJc5Y54Q7K5
ACNenju1KCm6vr2DlTCdQSj+l+khH77NoJmIEcFzvqDLdtlHBDL/fXzwgecJkTIjAC+fb5SvTpKa
dNBuE8VBAiWcdMhQqzacODZ81L4nhTn3Y+wh1jdOISXV6uH9rlqlAc65dZBxkNwem+g6IRUqf2f/
U5YZ7RsK/yRrGKg2ZuM3o8/jIc4E6r2vzlDXWh21/8E1lh7ZQdy2jMAJEUtAagxqxex9MeLoockQ
D4XdL7q3VaYtX1WKBWFMrKhDkCc7sOVxl8uM+amwFDvN45zgHkqLW8req8yi1lCL/Q2jS8Vw2yVS
U6l1lZfkQC32RHeZ8tZrCxmpA5gjDc/AqMtyLpsawVIUVQsYs8J52g4x8GK3WeozWIyBu8Aq9AnD
VhVxE2JZkBxB5x+3Opdp0nVzlt91yi9e6B6pJZdZXvumCCNKaohsTKaKic8dDvz9C2cVHozc2rLI
2iuDic5tOXYmkqUQeEDB2YYaCyAcA4oQ0ZP18prRtRcYeYcHd/Aq5V88JTlUtTxcX3exPJGYEeGU
BdN5tzkkSTDg1RwAYIRVWxynuHtHYrILvxijJT2aO/674NPPYxYxMNDK85W7ATXiPvy139Tda61l
kUO3QCC8I9YQ2tigmZvAzHKVeOf9B4/FeR3T3XZKE5rKw/5MJNboQqKWZuJRYvRaY0QtznmAyEeC
Ei5lnKSp1FIr+I8tx5Yzp+FHobS2e871sd/dnRbdDaKOhlxB6W/Y2jJZmK6VF+NfqQZLOe6FlEgY
j5oP5L56zYbFDvYgf+YGRh5hYqNZWFi+lOYgv9CBJK0clLl5+Yu4mJ34R5Yu+78ZrDJf41NeHqgy
5OXkzUB27eKTSs7vuOCHOQzICaa+sGr5180T9/EPnr8tO0TNFgFXpGbhpZchm3CDNAf8t/j6gw4f
CktqiOpgoAXPAfhtW7J6sSzY2sWkOd60u3dkYh7RXQaBUcwsUjQxCfoA/k2mCD4YQecGfkq2nZij
YZeLj2c5/ii1zJa18v3/+NMjCkBr6gPXhguqg4F9KSvbuJnWjQfYvOm0ZNkMK2k0l5/4snnLStK4
7WuOHUOqUHCqHNo0tbXSi3Jt1cLiiDnmVxnvwR9QtxpO38hZZ4OOb140nSG6t5AlLsuhULWM2o7E
PJYRtgESjJOJjAuOKrObt+BXj4brYs2y/GgWNFEQke68BAU9R1UXUOEOMM/4wwO7JEdYqss5rh1W
7MXxrLUdlfzOJi2KmDvr/XzymeqIwmD+jwqmgAHhVe7O84VG+TeNkEDl0DKbx14xmdur0Gx0PjOC
v/BbTiiYAPujRyti00ZsYRc6zHpjjWA2dofwLlADSczGo1M0uJmioHOUGoUxF8ImcaO9w/qY2UGY
vdAFpYcLaeMl2GCXtcMshzKWRHyk3gUC4NM19hhPw8SPWP9RCSr1JJ1FvomfEOjDLjJl2P03vXBQ
uMY4lSFOtxzEsO8z3iPK6I+K7o9GUz6R2pdQIklmTQZwzqymQDZQws9zs4u+g9ZD8sVcMjMmjPX6
VffPpNB6FKD7d84iVsCA+q7N5C19VwpcgbsQgELpKrJexfSOWbqgxRlodM8S4fRuVIJR7PEmjQC+
OLCjZVzr5gq+TgQqQ+Mkgo2iUMFk4plf5nCwVST+MEhN4v9nRHh7Xwpaq4p8X+P00KQl64AAyay/
C4zPhBJ64H9H+KC/ZYH3K/e1VeQwNtX90YRSgmwSplQHjDa2z7zLA5CTOZfbJFdxJrUSNP2mQsL1
iu13ErkEdXi6PM3Wbhokoc2W8l4hfwTQeD3uEZR56LCOu0z/bg7kVwhjhfj6tqS14G/KXvZbE37A
s8TJ2YQP1G9LyhO70b/zMRaHqjinNR0+oUuk8z8uVcnnKlNfh8xcV50YoDups0RO03xwpySOdhMk
zyxKGDlLBJxBe7vMSd3M7LpzpafX9jBemDjftc+1aMXHvmw39WwpwaABx/InIt5x+6sEc844kQ67
NspxhvOfH1dimOEu1wIXKN/Kn9Nm2BViWOrKo7QGTr4XeQhGkJTESqndK8A46S/awbHggZH4utqN
eUM+FSiQXK1rAPE4yzLmR8q4aRYEA3aPJkpbBkyylWBAdLmfdJOf6mK6k8m0MEo9XG79xtXEB43H
2bn++UZTDp5HJ7Fn0rMIcvEK5YWcUE1WhpRDezaQH9NJAigwxKVPMpzyrQHhio3MYxbZYMwR8I35
YBHxYq72uUb2j1L4tvgwj1IAWQI7nrmHB7PqC+Vy4ADIg4X5b0PXOzU6fzzfgrsM08q+zezOYaOl
qU4aguSF30M3G5ZjGtgag3lEXgyEAutmWROSPOAPnpzBlvC0J+S1S8/ZeOgT0vE4XkAB3EsbVimx
CJzpQQ8c32x+oLp1Ym08AUcJBwEJT73rc2W4CPOqwI446S5qmDhqLWanmLP9MQXWHmIBCmb4O1xj
RMzrFsY6IQaOyBR6R01JVlEENFY6bVWhc6c3v+pu2oIUvo5vW6t6H/njj9c5nqdP+kmQY7sSBmqy
JGulf7TIm6YzcRs3Rr8aS19RnvMk8n9bN6YfzoyK1t+5KWccxCNRUmHwzWZR/TBT0nVkXBb7fgJA
c2c/VAGx4hN5jHx/g3qdVGsZ1ZHocC4tgK0jbigAFL6u5EIqDPxi8gHKdHYlxoiZOl7qPGiZwzyj
ASGCyZ9acV/jeZLqRGCLlQnLof7Yfyce3PHsqjNXA62mJ6MClNyr34VvGjEKXeQs91BIW/TuD24l
UvfbYIz/RlAl/8yK2Tsa+pV6uUEJECle6qQsBjWS6F7l//i1x3PmMwlh7YAs2k0tNsJO4n0ld73U
qJhIc27DGUhHLXmF0FOTAhWppnA5+k3JEzK18PXRQE/ER2Nvvixvmyd8hYK3gd7aKgKgE9YGr8eT
DfW0FLD68YX7jGh9LoQe0w+LmmPIxdqH+38aPnDcFzFzZjsGoV2TqCC2hmWv0RFnYuXgtvdlFZvM
AGFezHvEDilgEXoQgnW6SWrNDJslgq1+AXvWoCbTELf2cUEFK7yqvoiNp4CIEHEli5GAMpVubRE0
DB2YuTQmr8BP64w0+GTKEXp1hBAjznNI32+N9u+UOH6uo1lDSsTOORJk+SWd/LYfOiT418ljg1nq
GnVB9fM5nMW+XZPc26Vpt+lyE2j3JpEbzMJzINyxZdKJ8HBnR1YBSeTu15qKLxTe+QZKEParjcXP
+jP+Jc3NFShwbj1kNDoXHjNlcsRDeDT1B2C9bYizcdbiAl5dpscc+/PixgHyPYwKinl5oEODhEL4
dLWTii536sGjh7bDHrL8fvuO3qqPrRcwtl9i7qcEjK78BITeYVZ5I819p2wa9LNf+TksEUGHap+U
muEiR6dZX8DvDPyUWGPiGFC+vCyNTD4R4ke7Y14Hu7roHG+r2jJ5ErChbrA6+6Go/NzMFWMjsLum
d5VyP5OOr3MEbtGYCeaGixKUdLv/YUFTQZlQWdphje2lgRxZvLSl9Fmfc2VuL1DSb3d4Qc2ZQuUl
hQ+MtaGHSQVQW9wpQQpRUS/EyBbYV1l7z/XuNAX+6dId66Zk64bYYDP0y0VFldnIOCHkJ31WHoyo
nL+vWmgFy8lW154TZefyuDOeysDSVLxm+JRlli9uBahBvEycjIqKy/vCgLeDUdKsPke1dC44UphW
/GWUZBvd5O3quOs8RjEAIsdP/hKCcPGg89XSz8vPeVRHORXmDRY39lhEQK0mMu7fdHcyMvEsp60e
q+LZjvpK71ZbAfVao9CccCDBtKEI+yPMu1t9xM/3PEwzhnX2vWLdl/zaNpuOWzE0zkETpkVdFC+j
uvELp3F1U4B84EAbYiwbGz9V72dJ9oembGSVpy4ZlqwK2p4pmnCvqUkwqHVY7NsFDI8uhz/22QuC
7wOZzX/LDEWmAKuF5rRkUMmE2w8SCTLPlb4pzFJk6rZvswxCQXcST7s9QeMe0dVodmQeORf0eg4b
qde5EYMXKmthPD8YeH9LQv8kpiA4FX2fTytHsSpYGF3cYjtPF2KwskTZ20q5MMhJu9hmp/cnlHj/
8EmkwLNZ+pVg0o4kE7p67DjTQ43X0IlDQFwxyQ4FGQcoZvSyTr/rPKefRBRDDdn2gMJkNWLbyMT3
pRbO9jSVZrFfhaivLRKL2xyeaBqgLmxDyHHPVUl/KlpwwiN5CBfGWvfGrvnipwWHLYfxau5kFuI+
rDdFVSMt5EXnnFYnqk4C482Z7LLQaau6tUgEHj/YTs8jhMC6yr9YWGnBgvIXb4GeC9huCy+pv8uG
HXsE7xW4PtTxvbziCBhYrxlGWzIv+U9b0UznUx8QV4hqsUOL8F2sLI4IT7cozFQPnAgdpiTirxne
96ed0OyGrc3BZGvx11BH/PqOjOS1hHrilM2xMtdHpYIqfSDwfJBZXn/3ayoNuVXs6EZlsakl4aqA
hMgKj8bYIzVccPcvHbBwn8EifkGsWWPutDxwYpLpacI4duNk2F3k47TitNthQ2qRcdSNXLM8w1G9
ayFBwL7/8q4fl2hyZW2X+Gf/Yd8V7v1JPyuWhlcTFqlHNIatSj79ZLGFkJCWgvJvUn3lFL2NUDdu
TvdJp8QlxwceSm+yR87G0HDV8lehajdIwzjh3Y3Krt6xGHXBbfS61ZPl1MXZF+cXsSOI2SGoO7sy
jcryVOmRLq4jkn8Eut2i68zT5Slwl8Mv6JS3U1S5OnpHo0iFK4Ehq5cawo166ZoGDnLR1FE9WQxH
d3hSlpLKKub4J/c+14i5DY67H5qajAEsTRlrrVtpRHL4lwh+fTQ9zHEcm6FQy6OBapChfsU4zsgC
KJU2ODiLaU0JmLL3rmOYgANglNWRyAyGGeXzGgcosql2EzK4a9qLlFKg5hjhRKDQLDdl8cW6EaY4
KRgC/nyYygITCpKknlM7GsupB4YVZXw74CRezLIHqYZEsAZSTsnctkXcTkb9fpk/LwfReuFDLvwW
DEw1vkYIfehSdG7YYBJXjLpgqjjj65DSVZ5feXDIqMQDdytWuaPGpd+5pNy9rx5JwR4oKOD1m+8b
v6U7BoqxgEuqCpYemOFMpzAYOWzaEbCmonD+zbbcXyArRodJBYX0K4YHCqBPFdMTUd5cs5DkDYD8
5T0ha1k5yPWwhy9upWgvtjN7Lg/nH4ouPMaIx1PUoDzaN8mJ3fZZTKerPcC6EeDI8qCDDuPPIZ2K
jgDwfTx6S789kkShNCCn6c7cu/aCOlX1MIv7lXnB6LX5CMrpv9asgQ04XMEqhXpxqUh9Yo4Gx9DC
pdQakFkH+yhPAIksjRHtTohlqq1/r13CEjV0iBYbGEcSm4F02XD8mo2h+BHYxiFgXXZB9qs36F+W
KRy5a9XWp6/r7i72ayBeBuuPndjxoQ/EnQ0VglzogfbQpv2KwS2Cczju4Yz7lhibodpka9tBqjZS
oYJXl2OF5XzUg7UYc6T7ftNIKx+b5FIWVZHgOzGYyP7G4VlOZH2p4G4gzX7NqrElp2/gDyYuoe+Q
ZzktuMIT6KUm4fM7L6j51T9m3gHBUrXr2xoTY6D+n4JfpjMwGi9tS9HV8tm1fd71FVBTNkyT+Lvv
t60YjJ9HXWyXPmpYCS4PSCm87dMw4wfUM8H9nmZxkP2dhP/qbMxBTnUmXHeCe5DPK0AkIEaDwEJ5
qZ4f9CRvz+5wtwBfYXNo6M6PB4WVefnvm+A5MjjwpOJPMGTNmbE6A+xTVTSIiqrvDjhKnHLyyYl9
Qv6kH8xv4GrLKgQiA68iYSu3lVvhNB6vWjWTjBh3lZdePuMx4ODDvdNcVGVcll7DJ4SUG3Bmta+8
ta14pb+oQRov9pR+A9ciTSF3LrWDVMmYolGDUFnFHHJg0Rg+L0lcm3KEPcx1yB3LtoslYvztoKC+
0cMl0jLWTM5zIFrtIk9mvqdoCl/LnMx8nCwQqxe7FwxGxsN9Zug4V4DHz8cvZIjHXu0638KXxTIe
CnLCxhPbknr2+T6NAGIq0TmpHt+x2yxKGLpslNUboUj+QO1IraI6Twp8xBQk4OrF5GNSpnsf7NEO
j7iepoHHuU2M3U+4SvDn+I7NmxtTdTpPbu8BF4OWoRdY3sZ9xdJjovFHddysdH1fqmtFHWcSiuXK
yK4qczkIzWOQXyNujDVb5nYnE5N2kSJZYXzx4szsTt3KcS4IbHrH4/tqp58cY/BTn96RRQ+SHj+v
iYVOUAu3xchduMrCQhUbChEqD3ipObuw4fBCqKZq/ayzDDqpprU4EfuwAiO1gX4kKUmhSIi0EP3j
pV2e8UBRz0HLFQk3NFiDlPR6Yc19wM3oeWBGFx+NZcc0NM2udHYQCR8oFgSmBAU6Y3KZ7nUOaXAy
G0H0nvVRtrfajtVF1JBj76pgFp40IUKLNQEIJIE2sBaOGwBL9fj09UUf3OP3JUX5Znbz9cQzJJ+G
RKCc5RbTs4cybaUXV+QTBRxr3jr83Gqsp39LBdEKEDdt+pi8MYayyWHhPfm5JrB9vaQaMbBD1bkq
2wak/jLwFtL74obyjtxi4kuMRSky17CR3DU3VX2z1bUPCbSOWlt8QQwkXQl/zf01KCT3h4paFNgK
kh2WgCyB3D8Cv/b0x7TbGQG9aplhXNXPcpcJMRkov9GRPS7MDq/kO6/DH1Mbj29i6ZjTP7qZP2St
3CuEttqcE6LbEbHXz506ZYTVkZ8fTnhT6h6gxdGaBN6eFB7mXE6lyba6Rw7/vMbjhLlC/6UaI7XF
Z0++iB47OL24akKpRatiBu8CcazzvqMPF6Ny9p3c3FMdx4XP7chBLo8qtF5gr+SoTPwA56Znr5Pp
jnpIrZy43kJ3rjT0uh81dAdMfuDJ50h1JNkhWu/m22mFgYsrcluZ6wgo5hunlnqxnev1M3KoTkLp
aLQdBfxjD5gCDdVCc9nk8tpwqsRWOVmW4zGvFRL9Zex0yA+4dji4zSolRn5aYDR6LcANxTKrDiuN
5WzM3ZIiliZBQwKGoU3C+E878hZFzHv6McQCDSVjgMJGG5YBoJ0r2Ydg1kYkyCGIfTs4CzdHIupT
rDFXCLda9nK9Dc80jvwmtuXuIweqPNZaD5/gnweZXObSnst5KFfT5uylRd2Zs8aFXL4wXc9DNhHD
QkAJyCROEB9xMBFhcT3fYB/bdHBa+MHYf5sXQSlAvq4QXN7APRD8GW8F4ymurPoHrxaPMiWcC/V9
Pf7zbB8l0XkfzR5WYVu0a8FBUBCraU4g9itkkWDz0wMFtHVgsQOGEa2sg4LlS56dvfrp3p8d6Sbu
95WKBVNiEgw0nOgSjOtK4HLbAxJWsRggui/XP9pnuqxZ7TkuF1RaJMjVW7No81XCdk2sbDsNS4Lz
ZZrHvkz5G5ZNvW4TGbXbgAoYfpaQxDcgpMHUJ3gsVK5NiOWKT7c2mEp5p+PC38S86la1hwD6/ByE
fwVbXkpXu8tcT9fwOoYgM67xH80lZzTVK736+abG5LLlpYbdojgGV+9Jtl7wy0XktTtbqnIrBhlk
ZBbW+hYpiO5EJu916sGvyQvVk6bGqQcr9LRWQmfz0A86DbWqtxvVVQne9wsp90KPv/8VjEPs5rSw
Za76enuUtvW9RocT/RdzddC2ygQt9ScLbrQV+dJQLyZH82TKN8ML6J2j/ipRZ2yWXrxdRGPBcGmm
pQEfRmI/wy9rco2m/xRLwiOXGbB9qQq/ihVgQqAAL5xOuhEIj1UoAZd4LBsSPdQedzJcanJEU8gJ
hdt4LjOYZTtO9VZyKGXmDOpDBlHTDMOLMG64kOhrD6u6Hpd214w4m/qK7kV18t2btKwk+WHTDwdB
w6cpdtXyHqE9UkDhNnZWM1m13THKw3LRi2p81Qs4R8VqFWRhp9JWcqPaVUO2+wsfI/jeVLe5PgZ5
7T8rxS5qwR6aqiT2siy/ufVi64bh6HNhjPV3AGaH0mrlwv1UoVBs9/D17UXk0iE0jSwbLc+z9tP2
Q2mE5Bl8/UYkMVLxW0OVoXltMB0+8JCPHkwFr+f1HwTVrBMRbyaQgXGN2iRL5U4FYfuePkeNKZ1J
3OCBrkVJ80hMjsWKJq6BcP6N/d0pzZ5kEJN50XrNDW21FabQrgcLrDmz5JmK56jmVUUZYrsu0tEH
BGygkvM/mOAz88MitXy6FMe2yF/pcnYCqmJXAPEvXqcO1539wgvx5KqBnqDjsf9XEDbN6VRXn+4m
Fa5HfdwLoO5rTyQn6Gm2gA1C2tgCizE+GbYrERWlgcwcmp5lIRFQTbYx5TyB/C4WqMmGbKM6ORNP
p2NpE02edzqQ1vnm23VyGaFlul3q+fSc9mWJpgJ3ZCxaCCFHK/DhszgNmeq2OWtKyT2VUZt11RsO
eFEInNsl1zBeSXGyIT3Z+sG9R9/YJmkg07zj7Wd33BCB1gk49Z/S/4YZKuQwh0Df6x2sysmGDGL2
YtA1VjAvLfHmTPSVy51vorIvmiKn2u1YTOY9sKobGVh346PEBiQEl2co5pcuTk3CkK7hRt+wUgO7
8XNWA8cmlxNnCCIksn0gSWO2HBD2V53g+wbQQSoPbXOFV5tHt27YEhfq5R3R+hjb4uNc95UPL6u8
7BHtrVf5Ri0JIOylIeDuoAtZTjtRyEcG1yTgzCKl4y+mhbsIovnOAIqzDvvGX7A7YVne/6m9e0Ho
pA1/XUaGCPWS+oAaMHDc3kRd/V7HV6EWxs1+3Q/czmLzJcscoQBJkH22Cp/4upeRWIsN0ogoAQRK
yVHyxxud3bKzWBta5R1szp+3/v359H9uX3wrzmHrDJMMFZuNZ+cPe1ZWTuGvHhBz5KZZYfy9/G+9
yxEwHNefsG0oAQonlAI/7kmVVEzM84A9DICxB05nRbIliNjBsKjbiB0mVBlMGTclo9kDtDbBoGS0
0oHenBAlDTN1B4cePf4L2z454ZzV/+AXltDVN3/FN+cTeTeTttCiEjf5nSZohcgEk6UhlySBAbHS
qM9QxB2OaA44HTGv+bcGK9K5aRtP6Z5C2kXb8aue+ct1m1mGanM2tH+/U9VfPz/EM3Lvh6Nn9X7R
1OJWQAKgnVmYMT8UV9D3OIFwXvegmRl4o0Dzh+HLOcMe3LtuU8gDZjBEwmczhS2BEHWGjzKmzrMS
aYe/uycnZt0UeVB3S2Hd2DrLLJJ2VDa2H9y4zw82EX+VvQTmMYCCb6nwwQ7Ga9AU3hyhkeS68YRw
AUV9IARWuC3IeyXAoDK5DqGJzGqgOVYTQ+46vLST82ebsVNxGw93mV4zjHuIiuovSyFIzeVC8gKT
vr0LuRclAe7R4aTywA7v6mmg0uFG9OzFP9Z4cmPr15h2FZeYL9kVaDtvl9cjyHEiFr+x2anRwEl/
MS5ulLwzihe7oW3Bj2peoKLsAy9DeRW6rE12rpJnjgHDJpeeuWxor3UIjNZD1XJdFYdkDvxZc0iv
CdXgNBWgjx75H9J77s+DWqR0FB2ywNCOOPzNa7BW7N6CGUlokKuAxXLuTOed6SW28e3xSeKCgGjL
sUUHFpCC7TAbfuek2qsE8UwbcAXIRtrHinMCgKGuVyOWXDh8GYP+SXQfO2x5/uxY/V4ZwDAoHHBO
XX4IBYKBXmBizdygp+Ut+q+XwVAXX7o1tYN7HvumxEJYXED09SIRDvj2icV8jcl8dyti1JSlD/83
fN8XtQciCpkRBDImTWn1WWsl5m5sVlzQ+2Jr5DMaoRlz+FkcM1eH5q4YIQ1RePQVtywq6Tr2+1Aq
PJQRLf1Rj201b0M0/QYCXwFcnTQWu94ARwwG0bAMPzoxxONjUckFHlWPWH/zxxYzMEZ8q03JKTq8
ehWyby6SORtbMuhBsiNAR68yV9meee00A1+B8BiFXnvE61wBTpuTZ0fHQyfqNUgWtL4g+OYZ8xoO
uqXQzn9/6y7s5AkSkNoUuKzh37w8N9BiIvwi12YmPqI2HMM3BQzEn2TWiHZXJ9dDfskp+Lv0nCMG
AUJe27rsVChSSHloWePHodQVjNXjzHHIj0ZY9tjtcTvOjx3sKXsQF67jQ75U+UbQ7utrh561Vfnq
UYc5p41FJj017TP0k2anSQPOQwTfDlg9B6QIiJe/jdRo36UYyCYjzDrJoUBCCGO8FESvyoByzFVY
IB1o7EUnK1PgLJO/BxIOReJLrCj+Y3XhLzNBt2hYR7cmV9LTdasOO+rELJZtkIOjtlQKWsme1Gpa
iyuJe2Mf5Fi9iWSuMyHJylOnbln/9UpBUJ35+ENrgMcprOi1M6+wDMdwgKiPjikJ8Xp5TXUlCwRe
Pc7PKxPB/BpTYrhZ5JsRGye5ED1GrWe4mCqZe5Z5Iphe6Q4SStHp8knFfl7pL1wgnffryBKe2Jww
HOSe4tpK3I2UHO+aRvyeGac77bKxHMBLEd0xGN1oVHz7W6Zxrh+6niyVXFQcVwfSdbfXibVGmx0g
pdbPGuAsAZlC88r0wDlK4k9dOOf2a39sPOyuJEuSgFcysXJ4HZdtuUt9N+nddPl4ZsbSCtCBIb0h
0TeBkQCseMSaBdYcDy0uH5uTb1W9F3p08lok56HxSISo9xnO8V/CXLvxcYUBUH/oBvwoUAXcOC+u
/5ydx/5A3lllzmZzzUuG5PcYXBzlfGnA1+b8oT2lKg8quy8+OQPVTJIYCW28+sm1lJrh2NwKGFT1
HCcMi1xiqJU60iwfWJbe6Ly3hX6pEhLrdsnFwJ7wQVC9dkGxrBSPXQSUFMaJV0RhvyRxh6Gfvde3
lkyKpS//kjA7EJqyQVN8ZSxiZoFMtvHBG62kt6e5BN0FNnLkGorsMqgHe/1xS/4UvUtt4HXiOFhh
c/nmUZ1ZyQBTck7g3ZHA6cRpk77opuKJpMomF5o/lYl/c9y6ENlql8WDN+D5LzaHpTmxboBa1Gkc
y5+2GVvy4A5mkRGLuOq1GnZuCgfEZyynpL3j9+jLeXjxyWqS3oI2zwjUd73tvW0OtAf+U5zbSMg0
9XRPTA0JRel78pPNMCaKdmpuVEX6cMep7pY7pfCnR26hWVmPQXkES0heFybDXWCEd9KLA6f5cwZi
Qy+9rDqDSmMdx9ACDb0rRch8vPnV0YwIpDEYCgWbIk8a3WdQDd0NusnaQlZySHNui71wmivLtmAL
lGZmIE9iwBH2Rtvk6oCGhUwJUY1ZrVG/eMc0lAbM+/eVqAO0PsbDH580eTMhAnX/r/dCKtL/9nLP
iZa0z7LijJK9rCbdZDH7NgwQJKUe7VbevrF4OtubQqz6UNaCDjLxYjnlhUgUUkM11vo/QXyOki9+
cRGpY4hD0VVbekBLGd4HzBmthjnW4jOSCO1/kzCevvB6xHSQeYOI7fbupobRts492QvS5osy017J
w5vbWlwbFfHxDCLxUNrDQiOniGQDYg9l+gY5Flrn4utsyzW9sc0shcx2Idqr05k1RepAbsGkRQTV
LBoRpzetMkg5/1Tj+pMC6XkpqLrkZ5Po9CLVBDnqREUvzU+7kU5GYYeCs8Z4hzMGY6LO/SWcUHPk
H1buQcwSmDTcvJxLNgSNuuNWxYrAsuFWt090GTwEs3kYNrBW9TP0VFut5LxqCTR6VQZv6szbKLtv
IXCUQajjHPmnJcH6Vxf6iEG52XuZEv0tJu/QH+amfJOIoLtS8/2MNAcwxst+KRi45C7w+pHHuJC3
S7z1LMUplfYC1QNeJvqboglG8ERl8UIVOhuLClqdBA6axSSAAWsUDFo7VI7bSBOLwkSrJG2FsiM/
vSbMzWNPKHuYtXqGKvqPDK7yV1HJs/vkhczSAo8Cvaoj50WTp5b26cK0eLJy2OzD5FAMJUV3Kpf4
zPXtGrtNpZms+hBepdVBqDT2f9ki41QG2wKbMgx+0GSFrjJhGRThwgZ24mKqBiK8ut/XrynTIYaR
EmDgvPk7IEm9FVxuGwkPAMhY7/ivmgVSyU1gNwU7rfmqf3tsS8hcknRYTzIFj3C/Fhp3jaUl08MK
shwhlvHFeeLD/0dMv+jT0g4kFru6T1LQ/ic0b+FqZ0FStGGcgrgg/Xfge0cpCVt9ohkb4LjGQ5Ox
asMZPEFBXRQIqpjnmTeKDcOEethEo/r3Jt+wqbHPS0hr4HrghtadU8vsSssXmwnMafYm4Zax0hZl
0cHbuMqeN5g8ZQOzC7PrSB8a0EBxX0wkgj73ltU9d22OTkajeIo0rlp/NLZJ/FGuuvIzSHnflJh1
RzAWqYl+l2jPQAKzMrFN2L6q5qNie8+CATe/NouyMc7YpKWW6tDo3Kf/Jb+ISDiqj2HQ6OQ/Fucw
OZYSYxilB3/YYc1r5bgsav6bbFQsLcTGjWmmrV3kyYNETRdfWo4UJkMWlN9aj6rjj+x8Iv/bR2Is
BnKhoS2sVBX+HAI/2ox04upIAnqfrkUJ9ikbeMoKxvsbtO/XOgGzG9XJ3dVt1GSJucgixCOneeFc
lxgxggcHScuJ8TDJjNe4emCXmhBkS17tAmSum5Pss6zjaECdyw+h7MTTnhz5rM+erZqgSznxhdip
kAHG5M7S4KSx934jpGjU9dSmTQL9rCiwdOpOPUnx1W7FBJek313Ay4FcZQjVwRB/uM7BUNrkTG/B
UWtUJVcKXNHzoSclUL3QRbvng43IWClWK64JAKdguFCm3aZxSltg4yTFMtU1mbJFdmAfusJnrzJ9
xl2QkFu4nunh4RUMGsJqyZl7Z93qlWJUkBhEEfb/k8J78ZnaX2uzL/vtW8UbpL6vMGNaNrdepTzz
dAOj1RlOXTQLdYlFriZQ4vF4UrccoWidp5JKUhtayX9OcTh9mYcNUj0e45BYpzozTus+uurnuV8k
GXZhLSof1qgNxlTD8wBb+Yn0TftHLEhj2B0u6GkoVr1Lyiyv1CIE9xcKOiCR9DiY/c0GOpuQiCbO
O14xABqS2xTIVrH4/bPkWAxi+8GU4H0vqvi84Y1PWnpWBxtXmcucDTEpu//l/xAT1/gLHg37TqUF
zddrbJOMRGdDCG69r+doJPN1dSf2xPVxZsLSJOEW1afxkhNBcXFwlspAG800ZG+0PQRMNfROvCom
Gy40zuws1h99c6JxcFW2micIJ/XYslka+kYRTe5UuKLZrQ20dwEC986xnqgapS15KhofTkTGl9SA
LvsSSd9uj+uo3e/CeW+d+Mifgzo0lpSgEA+HBrbn69MU2rkKN/0l8+18/5yosSE/THqmbjy0TbhU
Ymb7Gd/dX2Mr4+To8szGKrriqijaQR6Y54klPlT45IsBAfg+uGJtUeb7qx0zwMrScwsIwIcXba8d
4WZcM+2ESfU3zWW/ngn8gteV+WwJAmLRe/GLMB5aQN8FDIqMKkC8847g4XfOUNjw3IDTcyh04QX2
TvjJO7sl+BwlJj9jojDYRk3QVHeiOUa9+zIvgR5MbHgwfBAAc0hxhNICEaeSt5aNm6Kf/0x1HnHS
0YksW9klw94XPFd6h8rV4ghRvbE2XooSDFxuJPKkOg3CwKBiL1gA197hzMbQ/R+g/m4JoeQfb94V
dne4uqzuALaBc2GDwPA/UVtYXYC5ozXkyluBqelfNsbDyTzjn2w8pBd235S5rIDka2CrUjt0OqgO
RVIm/WWLvEKfdpK+zTfeLhEWZyGE98N+8eK1Mg64VGKRgk1WNJxo+BbAtDq5v3kv4kYsmtoW+Rb4
NdLUKwYjziBoWn5g4xnDkLG8W07vS+Ptf2hwfaNMNqWIjeVA27GwH0Lqow8SijAXG2RE5DwN5JtR
DM+uRNYQSE4cqFuAsxV4fA8u8Lfg3+iB8zvoCO3MI74Wtz/hJxzHN0PDkRRmrGQTnrucBKwrRQjp
JgCRnKpVEYYJr0nCWa5hXuYdkT0vq+qfCV8JQtU4OZE1uZqHifgMJ4CKQ4qIf71tlqzH5/3w1n1o
N6plKgOxtc1214ds4G0aODtb+gtvQKyl89ylZHSs/GJj2E5slXDYchLo2lO0p4G62ryolLjM7q3N
fSftA+3+JCPtNcgSHHLemYEQDYMOY5ns5QD3fDe0wYtX14etvF/eF/0kM2mMtqp8WJjCeV9hjh1t
zHp8tmNPVdmZzdxrq8ZWYoS2vphI/1Lt5QMxYrTYeeLYx4f8kTeBdwF2IjMwUfrNK8FoPFz8l368
1yVU+jzH44NorsQad3t1+beLfZM1kU5/PKYzowMpc7TcYpXm17vA2WZBeGuZiuak7ehcAnlPGV+Z
7IuzPBuFG64hGL8TBEDYlBH0LZUOQ8QClJJS4nri6Qe57gxz4nsokSW0pIC5+ndmLAmDDMVWs1DN
2T2sbkYzGyEmFWkXSztDeXJHNZZw8od7Efv4+IBBQY8E2I1oBVxn36oNRk5w89UA9c+K2VR8cLG2
iMM5TE9ZMLj82MYVsZ5ik7Dme7wgHB4WkZ7D2qDbDkiOKlN58QSzDY4wigG9hnE5koex52rGTOQk
Wb6dj70E4ppVt36qfHTLlPtmPlWZUeBGw1DvTwj+9KPQoJOoxL1z+KzWw3f9Qgn52YDYp+1qHv6y
5kJlfHhUyublninIjUgZlMQlOENODT4C/d+YkIFhhL/xZwhnLO/ZFjCTZfMJk7AiRA7/dq6++WOv
U1h04+xsKALT1g0cZvlRuHSPkRepO1qDmdf9YPbROt4leC6ba/I+EusC3+1H5cHeMZJJlUcm5WHy
HJ506ELPfJjzBpQwVw040ycbz1qz37uDZJZhAlEOc61KjzC53Oj+ZxbxoT+OZHyNHBz2zv8cust9
4yHq8ptgKWzujh6sjuV+uM6C16z83N/oFUWKa7u5dDXWB6kQsDcAYSPz2GyOQvOrFclcM++t/pKd
BG8fczaktk629PLfLb9GIN3JXH6VDTFa4NUM/gngNv8yZUK7uHs5YNwK1zo9kzd6TDRNn4pUjbiz
LMKGvpY7yuAtEubvURQLon4MwdHnNCubWG6mZR+kOzXqUP8IX5sU7PahXUHv8xDzV3AiYxwWWrNq
RPXLkGpFoHD9AdhYfITNeAUS6Fmd2QNH/0oVVTeAEb+2hknhfB4IpFcbRmI+fnVUjA7WU1Tc8tlV
jW1HOn7A2ebwnkMJD2v0E0VTdWd2kt+0ilTO0g1BUOctgpKGe4Vkb/UMlDVcskDl8aCr2OkWM4ox
8rJVXLmGZdlLBbjxSskmRMJQNL3UZSe5yYMhwhp2dSsvFv3q7zsmK7pgvVLmciSe2ruNaLnIrP9H
y0NukFcmZxwnGJb7cvNgLQdfqFKdLu+fzgwln6reWCJ4VW49SnkeH/5EYDXbvxGOMwOWijSug/a4
mpW2zD9ZSLsOzCQbWl5peltDJpbMNYm0L5OVIiy28Purgxw0LUfrOP/IA2rq4RrMTBO6kbuac5OZ
8zGZ7Due3IPoOIv+m0tx9LXKKv1EFqyVpCwTVku4NgofTX5qJ6ACHsLGxZAwcCr+6CtvYW4yR9Mj
Tnx0MoMANei3b642b2Mmec7Yif6W8lfte4p5DTyMLvXd/j+0irBuTO14OVZcPlgZjpZzj7dQAdWv
EEALfqhUxrU78Sv5Ypu2cllxCclUc8OhWa/NxAM5cPga+vvv/jV4BbF7MkTClXlbeDtxR31iNz33
SciVMZSMaLKoAxLN/R74OVfp5SZ/2z9Y8rq1zxYVHoprEEJIlmALH16drbWQokBuxR1OtNy7X+66
X22FTkrDQkWT9fx8x+WyYj/pME0HUlTYQys1w0SNsGREW6VfFFPDexZ/YHx+e5byx4IFht95D+B1
iQ7xw3LC8Dh/mI+yt7c+uu/EuxtOrs//NNLBj5B6n4Ld5QY2tRqezmMs0+Im+k7Z0tZNxkuOZFtd
EzZKwBru8cK2a60KmDlMfNutLHBCtY6gSsUTZ4kKAnCB46p8YCtjmJT8pK451a4ChgA1Zd/U2f7i
UnCsjdxVjUC7HfZo1ixML1z1vpxwQLMbwOnIgpRNI8QNHvxnCCR2398GKqdXz+SMDGQEvMPE5S83
T4mu/w+8emB3gxM23FoUyJ7gTyJSs1LrS+/Tts3h6xRcTQsaGIiTGIiqEaiqJzUgzMEWnxwNESvW
AzSMtmRKcHKwfZOuJc45vl1OJTOY6pBs0RRPctWhIutd+3/lhYCtVBFSzQXqQIbVVRebpJQeAzDm
kVEIbH4O6DpSeTVh2cJZrv478MUwXQ4Mwa4911V9NJXWC8T2eiwtnCLgx8L4XK3x2grV5kJI347B
YuMkf5rv/yI8egdoW6wFM2qPIuoPVpEvyrZDb3zyd4AHBhFTHDO7dp6GqjXEZhs+avhat2vV1osE
mYhemmsGTPRWMea+m6vdnqzuRGd1vY6FUiqPvHMnpMXwqeSxTuJ6j6DAFVSaHpj7GYlXbwaAFUsz
GHONWJd1kwKro+/WN+Qfjs8C5ByS9ffJ6GgfuWgjICKASnul1RLMirSZ1VAZkW9s0xYXi0Cz96hg
0YLzjYuTHYDJtEjVOuHijyalpsRuNKuqjICJWgMucrRz98PITGrZ0AJG3VC2f2ewYJEU7tkN7JYE
XDrL7vhmiuQvk+zs1RV1tAnF2iF2eWmo3rJKF6SIrc2RWr+1P2v3O6Mhif7HXXtcfT1Fbb0rwzzV
6xT/eB7KWN4rXnlk/Zn6RvNoKZoc6EJGtsQrRNgUfkWOBazVuVeoKVYHv+Z9e8QpWcah5zY4R/SM
25o/MHhGbIMdt76uYLsmR7mQxHfaTkbyjgq6erkz68EgzagwMCiloJARokYmGaAIqCUaolPiD1ch
SUXbBx/t+ROjKjbtFmKjcmzPkJpZ2LpcbPVzpI7akoZnzBYynoQ803crw4IXuJbw7DgAoeUvQSju
VOQ9W1a2/PmjNfFwjMka8h/jk4rxesx/wrg7eEPbkOTymBK9h7I0B3kmN3ZKijWBfbGTVmDdIOML
M2+2U41Ixt57OyhpZ7jsVzu7CnW2hjvBFYxyNYO+0IEcspSqwDMIz6OEJDY7HPTv0NbgnB8irfnY
QG/eQlkf1Tsw1vJDmjckNyTS39QWvwsey5a+rX0S4xiIbz0EBkZe4DziJsJyW2zxokI1u+WWIn1o
dFs1wTTqSt2ZWzNN9pChHiz4eUCgwzx1uvdxr0WwK2nFnDXcQmOanWvaPJkJ5+J7DJ8yDXLVyHOR
UrHfivdufIIWPlFpZ1jTsg+iaP5LH3DiAaew3ZDe2jDOANISl2gDkcDjtOcWLSP9cr/vhUOVc1yw
Om9oS+DEvH40CC3ugOluDfn49ZdCI/lQwrojrFrz/7xQCPK55nQOSsTgD3WtC+jd19P8i5fqEb5W
2m1nOB+CpQpSBhWLZ57c0coUcnlYiidjNl5kQuLrvJGrNJ0f4AuFJAIl7XEMbG11iLIFobk/sJNe
yxpoVVNS+pwNiDcx0R8IYDp0TzajtkXJ9ibz+IWSGe4QU26nlAA4zSbJpnHh3EW9ogcbia1V681P
rQ+S4q9qtXMB7FzsjpJqEwQIKKzT9dhEYF4H0dNiCkEp3GaxR6mx2q26Y7n2N2ETU4fj/+Qi/LWg
jRVgY1nnfLpkUSqKhjdlOU6Gu83PIts6H+lSeDuKeaE2rVO+x2hRCaSVdRlw8xk4XHI9+bNpVhOi
pBdZEE7u6qkhNeYAEtY3ycasbcsuA0cXup8fmyYAJGbXUo6mIcFd3w39jwQYWwqqauAmPUbwX6h5
hJ2X+iy8WlLMNw99sGBToxUDPmpKY6BW7E+mOZ63w0na64fgcQyRt2e+kdOXxJv2fNgrN5cifRmT
N9UAaKZvVbi0SJTMStgV0rHg9kFlyC4dO3JT8TnAnGB/PiFf4YP5JbEnUJ4oJxTSrgMPEG5Peqgq
CCNYv3E1ltEfL2xy6BVK0IGb5NK7Uss/zB/QlpSasik89dJA8ux0/+WUKfCaTndzsEixcsJ9uUI1
UPmXPD354CgTg3gTwOraK4+4uWnd3sFNmHNpx19q8zNDk6UdHiqOtHqKcglAH/EeOk+cs4EhEJVt
Aa1vHZVxJ3aorj4p1cbf3eau6/3PqSaihDHClAw0Gac4goiTnLpHs0O97SnEgCEBIXb6V113gGZI
xUJTLzJDMlutHfry6RTAQMwvHKApS4dfeQ7qK31B0TSAgZBhCGLh8VbjATTlxQGH1qzzX8Um2a2W
fwUEX3skL7Lk6dmQPGbCA9YD6xWGQ7sJfk6chnDmv0rIjvofg9jYOzW0z0cXr6shtFVvmmcbHdpt
CxdU3jVWZqmuaN9qnacdlFaFnRhqiDbr+KqpvSsqcM2h4Csp1gdEuT7O2VV1LuVAqIsVKtq3fzEm
8zW6QXfldHhTvYaz1/Xy0m8Iq9xbyha+fIxTNALxwYecmXIm1EuNS+s/GKY7IwjlEeV3xS7K/1n7
w8lyI4YELi1G8wrpgbnR7ehzDDuP1D1JN9vBEdnBO7sMmaCAI+GwzxBI0pFnvxR+Zkk6w5xcxToA
x1fy+hJQRdNeJilu3dgFMofIrWC7Pd+tKel14ohnGcyo42+6X89qupfQVBzAI1AaLWpwB9+Gk9yV
sWcS4zpiXUVvBeIUTPP/1iuTzaCwOq2T48VMaos9Sx4Gtn5Y4+80lBh17MOqi2vHWLM4lXU8tNLD
CGAEHMYErjdLeE2Vf9W+T2msvNqzojNR5TYmw4EpC0mOJ6B3+bwo2IwpHEJBZV3Ka/N+7eX7cLgr
FPIQvXGdVrI+BaVBWZPygQopNJKheB7PxAcWmRgBIcNN83isR0qXfBGIBTI+04DTYuBSKAtFbuoD
DIID4NMjs+ViSqybMGAqFx973nGTxRA62JNRJqKOxoPrRqnpg8oT83400212jMiz3SOksXdHd3xy
Qtz65lQRCzr7WC7br88D8ZkpRMt0hbc6cEfIvocVEsoGjy/VBlNhGScoouPgYe4aCumbTjjQFPwG
Pz+WGRCjl5ZrWzpxet5DIZAAmR5isuO1jkWdtMiITkUHZIY07p4L/ryR/h7R9dr3Fd5lbmq0VEM6
DafRUSRFgq7kY2t6vEDx/LTQ4krZZUpRaKoqznvImzLGuz0t4OsnqSE2i4SHuJ4l8q4onvXKtnpg
+ouAn53stMjiv9Vfn133NWsi/rVUTddwgB+M0ORjLpcgxp7D67iulkr0Gy1hXFVQhwqSOv5QHvaL
J0j/QYnNWYQcNggcgAsSScLxzLJzC1nuyRIN/K8Y/vFf9Xy1/AtBI/YxPF3Abv9qqkG0Uqk1cAW/
rGAbdHHu6IZxgnwTj4w24yEdNDWrS19NOLe1zg1TS4ORlXOKs5hHuChjukCSeCQSCyVv3Pkkc2nN
SFRkiDkFSKhQNmaj+9TFWkpOgaKH3wbq5jV41Nyh/Zp7WE587Oe4qycVxb+EFHnzi24ujjlE0NEt
XYOg9H6XG4+6OeoiNRDcE6uuHMR5o4ClimDxk8PtP08//wayJcvNfKnYFj8ItBARwX2ex1QOKMmC
NmM478ymeJjmO/Jwk0UXLsf7Q7d62Mj6UuiyqybCsPKgg1ECihj1heZfdapaeZLwLziXA9ZswCoH
U4l+OTV9oLcnlfbkB2o9NJgGIv6HvYWGYoCjhYutOAJidOeGa0ygIQQTzgG0HrrshMLCIiHtbTmY
c6q6SCyAmadH0GeSKJeukoNDM07g9vW8AscMKT9XorVSU5FaHDvTAbGB4pPqlZCwowEbY3J+qP+r
gRZvjYSvxs2E2OjyizgZaT6kuf1dK5RU50y9EtAZ0RoCmeOBO46Z8ijCJsX51xO+/z1jXWLxfudK
VZJsmeamDv9ML+xKT0eHYT9i/iqypGwz0qJKuCtBKJCWNnfIfq1/C6708NaEEam7U1GCN8w0IOo2
iGdf4fBJka1JSVHNJtAVvJIl4gY6nnCe/HNIW+rrQ8f3YE8WsNOSE3/joV5SEsTXrm3WJsjd8f1Z
LYZW/upCYrqeq8i3ld4GHUWkrWOnNDuzJw4bgwwtEWvujGF2si/fRYcPkU9grIJJkQo4zmsMJUQM
DWBwkQz01IE4Rhv5UxtoXVSYB8CzOY2y8zCl5dULbfKG5t4XsUbAiCEoygfNhvWsNamY+wUD5bEs
+dpSBSi1Apfivuwru3uUCVwgO2w4BUAemXhMY2z5izsmOHtb+2BmXOULknlFDgUU7Icaw4gP/W/Q
q/1+N8SKwDp2CGEQIHuTLZpdKCvBQdiRJqT9Tr8qTGlH+e4L/Sk/iK54MzKpmT5q4qhyjm+hC+Jp
sck5MZQ2dXZP38IuO/8KgyQItWCVFqPTCZANwbCa5UWsantYW7phHk4YyqV0XucfvcpKEhd0sc1T
aIiSY+M341QY2RbBRQ3pulzRdUn/nwIzB+E1A2K3Vf7KmDF9jXJQKt9RzlFbmvGnQS2eLA1LfgOP
0ov+ev+LVgB1Epab36S25RE+kuakmX4vqM9N+FxFF509HWsccXh1pjkUCXrapjrFLon9Mx8K65sk
I07cts/wtLbi5f582vWEp29Uhq6pGcCNy0aSjbxjtkjiyI2ocHyl1ar4wfxmNDu7jG4ZAvA2vb4b
CR79lZnIt2fuPqT46KN8lncBv7LG7iIilw4INsOwG1K38eUzxYkONVvwqNCpRI7QhOploC9e1tWG
BXs04xYaJCK3tjsbCRp1vGSEm5OmfvUNVpvTukp1GShUnVaecYnutqETJZTWTh+zFrV2bAbe6K/6
27vgwV7Gaebvs3g78regakLO3NV5QBYPYrcOVHWwzZtr86R1JK2euc4ctbypHcpT0LVESzyGFN17
lFYEyjeBDTb51xn6MjN3xXjMD78xm0Iv30PUXEhZpBmymJBWcy7ghoml1uLed8BwJWhjQqPg2G8/
y+5+nimasLzxe7LfQFqPQS5hlVnOuz3296EZXRKmfsQqLclPcP2W4kVrHU6XsGjQuI1w/dETep7L
GdqfhRNa7u8jbl99QhL+qi7Gw4K5LVXyWjx6PdZHpWe65t/J1mggVqDpYsfN0zfX7g1v5raZsoIM
YKAeBe64N3tcC+u6RMEQokCFYEZBzjicAUTocnTuT/kLt1rEKwN99Dy7yBqkABq+j5fOZPMHTuCC
fQ44ordnKHVVlukdMRji/rKRlH8PgspsNE5BsIr+BHqP8veJqoxLSSSCU/9UtxRM6/yhm+r+QnY1
23yz4a1R6ITSmIQ+pyqynBtg2gVcckat/pp98v7bJy1P2LDfHyHzozG+cQw/SqBFjq4gHsL8VK9H
s7NAjUEkEO4EpxetcTJYv5L21UIouGPSaBoaa+S9ZHDwX9cAtHIc/mGg3a9jEBdV8bpgAG2FDX2M
0RQMcGwCGS32bnUUbUd+XqFF9VJoIdFH2WUARcM6BVWvP9wcHKeT8pP7Cwf8IFTgZqPLw0tIdxAu
rnSTwoqsLJsMxS47M9WEnYWpslh0ykzbBG1Ft/F763m73GyCCpAGCaAiDtFf2iirj9VCZVBxRta3
fe6rsuqzzYhsNY6c6Ffq+90BZIVyrazWpD6sdlc8pV7/avyS5tLHFDFIbTs13Ib3J0f0OLyniE9V
chEbWTRwDblomDfkWMEznt/rRa9qqa58UrJzO28T0VKlxgTmzFIPzGNz4bbU8fpdcgaPsFtNiTSH
ZL7WfKwvGkOYtCDE+xI4ua2Gr2o5Ih24aR5SE/E5SW6JSoJmAEm5hU/l6uwl2XFXfS/UZT2R9Mtq
YcDSK20L1fCLVtGUZKcuM1GkVqUyXNR6H1QHwZfixCzJ+C96kSbeegMTlPx3r/abFlXN4ywaCugl
McjgfnUu53xJ1xn+T+/tAdS52UDOYKmpgxAIjt9J3npV9JJgFd/9z1lQLRcUGbKISMEmhob2ANuV
RbRn6pIh1CbEV3lNpEumHrObeeL/zSQuMKCyEa/mQf3R4KP4/cZHYzpFRYmRnwkzdtKlAE1/9qED
g8oH2rlbhLI5GhmvcUDkdEc+3H++y4CABbE7c0OJ2f0q8NkKxBUGJ6ayEUZuSAB+QqpCQ0kdAdBt
agw0RkqGekgKzhTt4pjANeC6W234/9vOfpoLqN4Pof28kcyXeZbbd9FwrbjIh5DNPGb8DzxvLiHb
7CNuYMzpbRGSJLgURRHLTrn99efIDxjb7YeyC/rEzyz+awFTANv//kNYnA6YhrX+NDSnSg9PzzUY
vS1wxLThyI1bGQ76cCR0YRFrY1Smb9DGikxxe7c76MgLOnzE+5KUROQXXpd3aKjIs0gzTwB6rVLz
b29CvoWMnhJkt1fJqAVxXDf6xJcKdRYCTPWTWM+/SU7DQxTLApwE4624SVbWHKchT/3P2lvQ7U3g
nzBPmESaP8gdcWsGtWx6s5fVUI1VqRx/WQoE2I1TWUfN/rM+WdWU/NohZoHegJr6dcNxG32L6VhU
as4QKtZeFQ8I46qJjqd4FFGgdIcsWG1dD35NLLYsoh74a+hlRc6Fr9bhBGc6BIOvIbUPwEIoeppu
lIwIk6cA1dJHQQq28U45NanugQVmiWxmoMUGi8eE9l4EAwLkUT86fgJyInI9dfsGfklwsR48nDzh
zy2e+56bhrDbpHwgbyTtYHCUYqKjR11f7okehxtHzir8xkssjfY2a6evs5T6FqJiJCDceVzTkW+b
sqSF1k4T7BBW4N89VVunnv/dPcs3dTjGHtKXTWQhsrGM5wm1uueH9s7Yi9z9qoSzltk4XE9qgYGr
jm3HfkPkGyF85QP3sJOYE1Z/7kyUoLBo7Q9ey2Sef0cviJMv8JxrvFYAmObGT+x/o6d1WX8Macnw
AuIKC6WMcN9PSzdx+4WDpHDZIrl9kusPn4dR8JgYyf57Lnwnlc4FGYceEU0LRuL2nbH/RAH5VY5c
HiyCmNiGm0768nWVmgViIsdZ9Fu3iMmctDgnwPouvkijPnYiCqVlQ+cF3kV/7c3RW8DP52eAfeyl
iANhlHVGH4lIvny4h7w9FUjblpyx7cX+mVONKy7EO0pdrc4NuvAatOttQCT3rznrJiAMczluoxNm
uZuUzubzexP+QnYhTTYgqg/xAmoqOtVWLrxZ4XyoglJaC+Rr/ur7aE/YDX3eKRt2Ph32vvZfWdI2
e4SKFiILRcl4TvMfOruypjWlpUFTI3KSs7CUB8F2eK+8taJ2r46LRErAHgVl2QeBB1dZotb/mTAH
j1Im3deH4O5PqfsywpN0122R/trJlpZ1bV7WFyOntiLYerqxI033M0FrUnMaMWzSjYpL/RLPp+b4
FHGCY5/Khtd1Jl6htIAGFgN1j1n93g23vwy/XseGCIpBFLzHmjVE8CzDWuHOsKd+H6ieHII8/AKg
NOj/Mykok8FH0XFq+EsDcZEvqhuGT15NlU91TzgvCPhcuoaE2ckJspdbj9iKT2VtsS98Ib1FnB31
zz8VOQ3873jRSGwRASQnSPmIiWfohlRAJ1/8MpSotXUvWBVWtrY0uN8dsNO4365/pEHkH5ix/Biv
IfHPTCg/PIC/LgTK3bT9UJkjKw4dR4QkaRFEWCW5Hv+tUI3rOx+OtWUyBjTo+GonBXVL9HIDkuhB
brNba43i6k+GcqY/h4Q5oz6LOqgpQt5QONyHZBrCCUUSDng9zxGNwyIT29EbbiqBHsp1WG4U4wdG
d+GaUohL+ab98DtpoHG5bIYwbNeOtt6pDFiXz1P/mvOVE0v82+6swhgoUecUckBl7FBmlrk50u/d
WTxEWU2kYRPf7rrl22XgCV4Ka5rcnXuRk0l85J/G8bo4h2CgO7byxuA9W6xC22QiD7Tcy7Dh/alz
PqrHybcEwsKORx5jQeFLXCn8Mrc0+wDJ0ijcR9ylIbWIu984gQAv+rxQ0iFRYs84uEjgROwn8WcU
SKhtltl//BuftNA1ehCIedqBrf9p015kL7QcJHT8Zr51oggJismSH9BNdD+O8N8o1he6FjMwxflW
ZxttjbquJ9r0p8OWwm8O/1Vii9MGx42I1N/v3ooXjb+5Qe/keYQ1lwEmw1Q5RF4N+lfnJfxPgj5t
g8hOnhtU0tN1yzK1w5gne02b/TfyP9puGE+TEFlIZ2/Qt1dbI9al8HaN8i8Dxwg5OHW+zULrTiCk
xmOJ6irGUX1YbkQ6mXBBwQmzK1FyexZd6tlCPM8qr1YjUD5WQVNGnRf/M7b06GYOl/LgIf7JVapj
FKBguTrPF06Je2vn1QZ9RxJ85Uk8dvpwWoBPJ80nCHHoBVeYM0JW07kldW4P2JK3db2+q3/MJtw1
XCTU4YXu1xp2KeE1X/y+zyPYEPD+EKiYD2Fash87QbR9AFc6uU4dBeWwdzKwVLwkA9U+rssAITrh
27HLYJ4QbXbajllFk3ZFU3j/mXNJnhOuxn02SG6hnvKDP7WpshxmMkAYbnUWvFIPMpf/FLVj+Aed
tb6NmSscUuElzthVz4oh6SUSozOb1CSV4d7zfBpfCO8rPEnwz5PF3Xpzls8jKEpGYZnBYYINRWb+
IKFiFs2x9vyfBhC53RfiUNINmXdWTD0SPEY2i/nMY3/Z0DFOTAjZZzKjvES04Yr6kc4BnuiziEVh
W0mV8SeIPMZCJtdYJO1CdhDyP0NPXRGN1zUUzWNPBWiNp0MscIM75EN+Zg6lQYN8OsyKEJ5lxQVv
2p9k4tyfqkHCietBBZooqviviU76Mnn4UYKrTqpPTO6wJVSYu4f/w4OhhidoB2D5EeqBdM4Sk/jn
n1Zwjl0B5crHElZt0yx290fzTG2ryDf3iqi5h8A9EsB+qXncZPUWQ/A8F5FU8tiMxk9OServ5Qqb
NtWIWWS58knV0E1xZBAFG6QTJeshuF6jUUFL2KVEF8Db8WjEX0JqV1Est/ybCj/sWqqa9ARN55BZ
ejzMjlukXHUWs1fxJpFCOm0OWjrF6WayzxJr7MUnYb1ukTXhriy3nio+UZrCDKR5FO62Fc0bCjmo
ftAT0ORgvGDSw1DYS46RXLqXdYzArYFIR+85lhlV5g8Tq28gdhaY7+O0ShJQ2SvXO+nnlowH2uad
RUZ2O5H6926MQttgpQZllGQvlVun6r92QVjEh5haAagE1Ee/rskb9Pnsjt+AsAoTjeWns+KS86ST
69pOtslrdgYNVq4CK6/Ow6UQOBXAtqeF9tpIJBHpZ3MCDIP4g/VyEGXBbhK+aDUgnWj/y6VlLM2A
XWbOFF6JFW0CU//ZtROmuKWK4ivnYsRFu4LwNtPfLxn6JRq9IMGSgQM+8jtSxMTksTAuPRUWqfhh
vLtamPDD9D2iq9x+qfaEIBS22X2GDXdBpCF9H6Tm6DsQC7+eN/2OhCqGGN40cQjMoLAmHikmo4kj
pTghff7tpRqnHaZdiYKWba/jnviwqWOZIi+P6v16aHGWkHJQ3IdsCzEkQEIBX2W5yXvVtczacH9O
Z4Tt/AETXccscS7MPfCtYunoSfJagFQwEvoM6jiPG7/pg0vHxdqaEnDRZKfRUqEA6ObZMxdv4V34
p4xsYUEhjSpFP0MWfUN3LoZmc/46ITC1hscDSHbvd+CYwSsj+P9oo+omhBixQlvR7hBx7iCAbmKQ
2SpIKm0gAWGNYI1yrIzqNprf2c2CeQQc0x98YwolHzjFXr1dZTV0cAuPX3xrbD5GVRwU48RD+578
HnWi+VvGQPVyRBZ+h/LYltv497oQ6LpG7Zrbv1i8dnezYtnlbBFJ76X3bBYfflkGEP6DUTKZ2HD+
sjVoFC1mJPgSTqlRzb1FPUw/sxXbjmDPi4DCHZWcdtch9piAuKdM9G09fNGuovxYemUPBuOFeU4A
etdsoAgMZscW85yO0N/bu8lWLVxPBlRfcebMC8Lctfz3O3Mc1FZaYKOYyHyF8gCjXC/b/lnfK14n
Iy8d2bDjmWwe1BztWQCUuZrk+VAa/cnVqcYUg2U8F8JKEodaQlFf0wxQrCDji9aUZggIACkIXK/s
HXPiohlTdIyxQR94D5cPUUBJRiJP0RiEuxwEZ9oWC7JVOZC69rlp/5cv02qoVtIfv1dNNdUbH3vH
UJT7yB9cEDDED5ZcY8uBW3PerOItYvUsaOK2374x5L0jbcLdSGEyiUE33agLJghFOQrT/KZmw3aY
MVy8FnU5/PA2YeZW7VnImUqBssUVZ92jpPpP9w07DHW2wrzfgnJXpbTMZ6mcii/3Sd9NW/0g4boV
syHikVTtAQerjnDbuWu8M3cq/HVJF3tdSXCpRKH+5t4XsdJr8io5vjTsRySoYkNV7trdrUT3vaLN
6xSF2M+NRgn2V8GZ2pQxJXI/hApL4qv94NE3yjln9wMBHduee9IELzWiOpMglflYZcp11H0Ug/H3
Dh0IW6I59epeG1DiECuypuBP/kCmptxf4kg1tnyydg5f1/Ax97IT5DVpAAYOqMJjA3pL4wG26MVw
W+LRO7UcaO40eTqCS1cMhzfnseMkjQXCFHi/UqNgK7kfpevGjkYudnCbStOITJnM624uDNJQkYW+
RuT7uzdRh8Pv81z3YmZZoqVrp13fHjPjFu9kyg5YRfRAiO9qmqVH1nYs35G6iUEapCao088sSZty
erH7G9rNRPTLQrOgEJxdEDAGr3PLYFzxJC+BjPjoKKMsa3tAxO/X0M1WAgs9EZb9vA6joq3O+o6f
34ng8NAEPui3XwIi/XAy1B1AQKmoNqZ5tHiJO121FbcUWoL5jZKrI4R1sqUUohZzvEV4S2g49lgQ
a8bk+xXHCDfpfby0REKEZk1Vw9gEUpsBp5PZDyywF3mXKKPUqtPyc86xcvHW4JOMcLGLO2YLy4YB
RIgwEb0mRfeQGgeYB2na1SidAjL7tNc2Qo3q00jwexk6LfPMLGBNVs46gXvQ4BmA1PsEeAY52olx
W5kdDk/KVtDESM06HGN1Bs2B2ev/jv3aoHRpx3YIgCaQbkGYzTsZnk4gY1+fvH6Jdfy5HcMLysIS
3yJS5tt9tdedOxkyT3W+XUhoPhfdUFkGGphFWtuiaHTrxQvhWxHNhfyyTlKjv3pMyl/E/pe7XUlm
Ojpc5jTpEchIbq/w+2JxiY+xZo2BgMT4LgBgyLaELVSsIge8upcKqA31cNDbn2eeuj44amHukUDp
MUWfJEKjoMEKbFtppkYpBl0nIj0PlYr9aVDPbmKK1uPj3MOl89YCKoZcu6/i5ShuzWG0teZYVmm3
AuaYPBdis9u4jRSFhQTwewlk+oritDIaF2MMWtbJvIICV4TZtVKq4fNJfLUkQx2n00kQUK3oENBF
IrgMULnyWOLx7rBTb39h17WPtZmZL1827a0SmR2VzexkQX1bw5mBMDYcCBPV8fVBwtVy97Y9ShUD
SPbiEIW8T5/cnI6mF2yNZfJ8ncqpDkFIkDFkfFdnNBSNsQK2cWptzBCg4uJgXx8L4tFpijtP3QVW
kHaRRYCGyoMiGoAOR60AO+WhS9kC1ASzwNDB3/FFVduMt7NQizHunZ1Wic0GnXv9ty/n58vV2aiO
ICsROiAhe++BO3dkBElJR0zfCgVWUOO+31vjkcVaQ0sC4/2x+S/dmNB/BXBfEF+dAksGtEFCfiPl
IRgLdtCHCORG419L+6GKOyEAbIwND2MxQu0IR8YHgwmKFGQPHdYp3KZGpq+xtcbD7HtuNyFGyG9o
rAFh1pkY6bei23AAIXAynyMwOJQFTyEDvTbCflvgOEUY5bgSSEKvzbO+/XUUnat41VzliMq0ysF3
3LGkeSxlHRSCgOruHDu0kAOCFh+XoD7KIdCD5ASv+F2kDo8kQMIjPLPdX4PEyse5xT4PAa+1qNa9
ETY9OxBlFe3GFxqpTapToWmaLNOIYCYgenOjJcGFv+2LR3d5pekWJ+v4RdkJoSWAFIdJq2mjyt/g
h9v58sFduCS9L6qf8dOGa7pN+SaEiMlCH81YAa5rDuhGWgH08l+WEUf8HU3sfBwupxH56zre/B6Q
TYfoKjKHYD2KMufRK4cewwSZ/tIoW5m7nFLVzQdSRPeBBg1APgWtZqBT3vUN2Ofx+JNph8p1AjNd
L0TprFhjtR+JtEJCTrGClHzj/c5I26mieuhtz22XC87wcVwKipd6sKkJcdJNAkK4Bez7eXgwekJK
WdkM1o+svDz7O81bXs93VFuMfSvASxHGrqn3V1b7sclAG6RQVhlAiL27rnLcY+Pxks1RmV0bhumY
BAILfAM+uWZU+4ZI+o55X/+7CXlR8j65bTfXozL7CzrX19Rxms2Vfz0fNHQX7XrWsn2f2r0Z+xTX
piFRL9O7vAi89UiTBAdTXQoe0kKSovzXdzJ2wW233GkPM1ZU87BDzO5hVW4+5Q9P/5i/Jkni6DyO
Lw6UI3zyaA6Wy01EQgybzU3s1IFwzlD6ayt99iq0GQl9TM8Yvpmoqt9XidHRmoX6RPTik/V4ww5M
iFCWgeLfWEszOAuzKimNVyuZzN8XDYQpU4U/qLftFzCidxFB6yj8Wxb5TIQI5n0yIQZkABuECjlx
r9wwiiQABC8mAxZbNfv7l4RPyDg4jTan4IvmM4HLiEAjYs4NOsbp4xK0vJhcoIYGC2qQfOizdKAv
a73VIY654VbibHUCfsbEp58vY0rZDNzgWYQ31nh+xnSG+NW2NylZSz5bCdnYxWPUeMXApRGMjUwn
XcihiiqtOsxNk4VNAXhTTMEf14zA0Hd3kzVv3UoYbuy2ChZuj7SWpBSi2dwye0oUW4/cZmQIJ7oL
5Ds055Tf63XJvJS20Y4pzmTke0QV7i0uBCFyOMVtGaMaazu8YBHlhB3YXgp1sg5AXq8hd0SWKexq
0QixjqCSqbBxQKRkr+4mMXKAE6YGWHzAhHLWzHEDps4AN4DcKGNb9E7gM51hlT73Js+bE5LiGEDQ
t4xNO18DoB0AHO1lKlRCrXZjsvWy1J5hqfFQS0UsUKNHd4n2USlI2sUxsZGRJPyfnM2YRAdrLZpy
8ZXNfBZnqgvk75ZlNt7W7fPXnTYK0RqNvwPSBDL+vboSKbrVNsuKU8epr5m+8epn4fZJdlALxJqx
Pvj62Lz807yVAe6JGe24kPhZCld9yuRwDuauDvgtVgy6i6oxFG3PKa/4YlUb743SVRSQlO2aPPkB
HvPhd9xZajIK+kdJzJBbAIDOpkRnmwlFv6B2/FnAAOUKlboMiSX8MtM8qhSpib3Gg8Mscl7g1v05
LgeQd1VR0SzmLvwTIbIzyCb2D1fNmfLxYm4/HiJ187pKoTpSYPX6t3OlPbYRTdCQcMPaN0+yzRzn
UdoDT5f/A5ou57O9etgkFO3sgzxM6wxPsU/DzVtTWM0oaeRmMLu0w68rndZCdba7uiS2aQOHikBk
J/L06pV0OuPy+fgYPMROQmC59REEgLUfWZPly/4T5Tc8alA/uwEffihV0aMOWhArSEjCMN0RHq7K
kwoBaUaTdOXQ/NIxjQlzXjoPsUULxL4eLgS7Ejg8t2zK4Nagx04mN9LNrCFe6hNwvye1hCXHP7oZ
a41cF1/hmARg4Hsp0dZjSnIEhOYh6cdkoYOg44gK8m8yfgmpBVFxx1L2M5fR57Lzq+DdIImu0pQt
3DOpIpmzjJTje5VVh13qEowllU1bK3gR3NhZPPauAxijg/G0eBRMrjijoQbOQ6oIz4EyMB4pYXRQ
5pCDV38BXoLgnOBxti2rsy2aqDo2TjxkHFpPPF06ma3ZggBPKvGL+48WC4dhfp0muNQS8sZzdLXr
X2OOKRNiX7utpmM+aFR4R4ftURuFYsYa1AJtAx6JUG9T0AwC3mgpCyjewQP9E74Q4pGPlltxraBc
wR7+77B/RsaNkEWWKDK9q4xcZA2leOiyLvi+YBQfEe0pwyivJ4cXzjZsO2yPjfKgi80fTn+ZnXF9
p62tMPww3l92DK7XvOMBw2bS1LeB2YcJlLxFnC4mxNKEnKpETdhnMxhbQAkh6ncbc8DWd3/8FJag
moQWUc6U4Un4NkfCHV1tiGVBdgd6ptg6G88FSX7BUQpPBhcCqRePkKZvdi/Z92UbnEtun61hFLJx
vYwq9w0B/uKX3k16vvTY16RFE9Xlt5JDRGZf8qAs8a8zd59D1WIwZ+nsczrOtQHoenbd4ssmb5Mg
KLSBS6yzJMLeIJ49hieEXgJFPARidWn5yUarQNjniz+TvmZ/bd3OR22XWMancDWPVkzjCwtpTEOg
4/RNiMdq5NyTCcfQdkvJPfkRuiIn3UucEh0Hh7c615qimq65NtyRK3FLhgJZrL6rNPZkO+kscVhO
FvpqcxhNFoOHvLUzfkLszMBFs4CwsZfvZrYNX6FypxfyNN8uBEjT6+M5rbxkWc86V/u1+VMbanDd
Wbvssi+Gor6eV7qEWJ24/6O1ImCFxhBwEYg2D5DscNwCRM7Fndtrrqm+suuuv1TC5TaJxWYF/Mzt
M8zSeplwgC1TxmPKvlraaIVDhtjYHRHVhBaxjSW79aoxXebAhaubY2VIPAjOroi1rp2S23z4mtqN
Y4nRk7zjeLD6eV2enU7i+NxYFr06xZ1EB4sV0+cJTAO7rzUpKeWHDyCWctnnJ9hmZ+b7p8jlD1GR
z6+KwOyhgUc9pC6k5ggoRPfAWfH8mYJ6ckuOZmud7w7d6FGayKw5UEyycmZerOOrXFTR8ZEcC7D1
r8TjXS3HWKPsDUQkYFWFJe78hIc/xJDSWNpAF9dhp+vRy0PUrytDa8p2j8qMl5n/4/M2Sd+dUZKU
1IIPCPcvQKZz8DwiJRU+hqZMTggAdSkM/I6GPtPSMq3XO2V8UzcOI1ow0hDxuHXrSYNzzM+LJ9JV
poH4H1OwPLL+6atJ+ZXTkS0h5Yj8/+iYzFSo2al8K0j5yf+kjxnRylxTcAVXXet75jb+23qKkDU+
OoV3gsPcreRlT9WUK0SI86L3pceX9tt9L4yliSE8Dpo5UGRqTHs5DYaAzr1+nVT+WatM0qk7ZyJZ
ycUu8tP4gVOD2JMpZdg5CnoLMqzTUU7tTwjE+4mrqJbRmb2jxqdlDUMMAw9MCgLfyaJWQ2X2SYjm
/WgMHkkjEs+bIKPUaStZ/+n2KJAFtFHu9r8q9OYjthCw00rG5IhyvEoHgY96lmhMi2wmg6B4MzO1
NK2EXk9qXlG5SH+zb1sPVhhPJYwffYxDVf70USk2KeowuB3zu/ZBxLDuCMO0hZN2KpHqesqKJdwI
uOZxE+l69j0kxfEXGJkH3E/pfB+hMzrKBoRTJRLL7MjZ8nvWm9rOlmunQ4S1zdKB4caIOhIrFeqR
IJsT5ypf/Ltdud88YUlsH8gVfhTgzFBAoydacJP9DxnDaB+ro4zfRjuPHqY+H0tqj1FHZXfRKnpx
pZdctYKTL+AEsjWI9NOhXt1ahztgN7N2xySpiVtx6QDuavDJYy+PdAeyY0SSBsiaMpC5ginUOpxm
ZhMITs5I5hVqhulooMDVIWby/9Rl3EoTZuM+A/dVe8/p9pfp1YjCHXrDN0iZf4Ptxdz5x9tqCgnI
jmlroK9Z10eRzkZuPNyFQfa+4pOepk5xDu0rXqsspy4owcrO/RPP5Od4aUrS4nhqtlrBQg9fbW0z
gew6GkRopjfSyddnZ6zRLWBe/LYTLqCJlJOwTFONpJJcFog83oXxjUCcFe7OTftKC2esxXxAVzch
34uIiw4yKZN9I25hRY/lL7EFu9v0cG+RTsFWW0E+yA53Fka5Bt4TwtPMgp2KI7OiFFyTRyk6lVSB
hoZolC801eWSrT3f6zO2c2P9MZYDXRxlqIvFQpfPwwfWXH5kXnr9XSVfgjlSprgwxNDNLPQZhSM5
zC8PcsZm4wbRuzpU1I5GsdzrW7K17/4K/883EVkCVKuAgEQi2c1pocpXDvdREnDsbrVmXopUXt8N
tJVK/D1inueXBYu74IADoaBOI4TY0j6lhmxQpYBIBR66kHDmWbe8/7QvJviwRgLjEKyAukIs0Ule
4EnHvYaaEFZc7lhPRUeA2YJB6/PasSxZh4KGfFxVW4KOHrogqYf9bB/h4WagBA+FlUNw3Su8c9nr
nwTJh0Tw4o2N5a+a475Gst6pbcNx+k088gzw2sD64zwg6oWhWTpDXANnz4NQx36gc3I8cvl64Y+F
hJZKRK6vjNuNs3UK1v/H1xWeMbH14pJ0+L+RHsRYPrzD3F04lRg5ebHG6w42GYYrtoadRDY+Jw98
t4gtEbYd/24Vs6muFl5e0HaJxoUGpxo4SFuwPXSA4i9+r6KPTF27U/BBcT71bQ94CVL1/QPoGEbg
BhHhCi+eLzoCruODh2RUIUBznssl6MIh8H2hN17tLJhusco/vVtKtkJfQZ9IcLHXV3jX7RT/M2bi
w411w9yD6H4ZYFBG81LTgMaBNeLZlhvNftzfrKeShOX/tgQtgF+Cm6q3/toUhtPhIClZfo/OVqI8
J7w4gb/95VvDis5Tx6l6AYBG1UcVvomvmJIA/o79qy90ClmSIbgr/WiSX+fe5of4wjdu5K5SRfZ8
xCH4eNjDSvl7UQBXRBJA8MXb6XFaLX9Qi93XbRQ03sZoWbjOfu9IS2tpNc6DXR/OW4TV47BDrHIP
XINnD9IFKWIA7gR49/g1JJh6flxmbyj2tF7Nb0UbYFSY7XwKKgekcN+mCAVQ1jbOsiQfU7qff2hP
zQWQivoXJAiEM8dkZ0PenEwe5/nH0XMUYmw4YdiiBktkHSi8mvs1PdS5SCPsOXO0KBxO2Ae6noTr
na4/WH/Gk9v5Y0ksEXaS4ris/q/QBnEby1muIHfm/k9wAF7W/nGYL9xoHR1KrXy1bzRDE4mmrgVs
odkAUPUPr1Hk73sN8pw6QKaYXP/Z5P9UIbmzXfX/ZMdtoaNYtxrppezBoc+MAmY8tkdV7cwtHPIK
BtWaqOP0AS9a0jO9lHJJaqZoF9pWXdOPH02Sy1unxpzg4oUgxCzfoMWF6rP9HW/zaPZtld15RO1u
eqX0hZ9lIow0J+RvUdae7jGj9FS/RVHvdUirIi/+P0DfobzwsynueQwor/Zkv8AuraA4XAQplCXe
k4tiMcZri5tfk1UID5IDN9xmX6xJxThzaV3TKsm5rM+TtklZLdtZgPCrGAMR1WegFrYhmGe88dSc
wnn6NcDyd9Hnz6mz2MNIxHfZzsQxsMgJ0hAaAVKLHdYhB8C+81opoYcztawiCoCThdE9ey+qKR5M
iwcVN9VNQx4BJzCpbH6zAyrp991ISG+XuhnMROtHlbIvxYXphzLpq5dFig2JxYzOvZcRmGE356Qx
tsGH+gj/qbo2Ezf7WXjIr86WzSODbCUtGn4lPXfqt1hm3ZHjVFjPs+cqc+kL1+4sC3kpkON86vx6
XH1kxA5R+whFcWZFEq2D36nsO6Ii2SSZMOowuyYutMheDX03S1xbZSchf5kEJ8vWJgA29RkbLmGX
PXmzxe8rXeHiyaJHNRsEnwQ3O33NWNgM0hJyJHZuAwHiKu+IxmiXEaOhckF8WePg2cg87jEC4Wj+
wfMMYl4Vfk4Qfr+zl7THN5SckG9+DPSeZ+2CtX6qhZ9/XAWWm3c9uYMSYs42eNT2qXwVn49Jca1D
2ZGUwLRxPKGtoPUOH/IQzb+yjl0A8qZdDO3X7nDhJ0AYtEjDp1Ap1KyD7CWU4DK0OhcY1E9HgXNk
tW6hp2ypsSgki7K0fTYDwyHNvromj2eyP//+aveKzYJpwvxhVTrFI/0JY2HyAkym651o5URmTN0e
yo4u1NCJpAQii41Qd8L43wmt7mnoZFhUXeV+9BI9vXaygMlwMT7gAnwiVKPhiCYj64K32YeIww9j
UhUI54nO30TiX7fKjhvPeRky0jR/d84fSfMrZEuiyhj4UmcmCHs9xAiSnEPhSsw6trAyPk6UX5At
7f7GNgJvQohUmbRSqShL+LVUbikwxO0P4vmGh85i63+gs3kDZwCOA0DluAQKlpU9c0WVt6/aPy1Z
/91ntO14ajGs1NhXF7w4s3r5XTI8ply7MiaH6IWCb1ihpFqam97q9zH6B4gblxccBF9iyZMu4X7T
fD5t1KGYDz2sBsgoMrSWL9DAG/eFpfvpsFb1j84h7fQarDx0vpk8U5GGMBdfvIFp7mo3oen7nPFV
3bGL94pxQWzXShBMWkz4UdkAnPVuOJdSzxlacQ48U2b147Lg/2Fc1XmMEcQWQTl39jlBL/C12hcN
3tRkHi14zpBgSm1FcdbJUXKGqPvTPGqfPoO0cy/Y9zk6uGuTTOwm02FG4wte0DKmgy9hYACslnPG
ruYZej3Z1n0rCSBNM/72RII16+Txtn1APyKcyCuuDjFCKISYDVsl4TSKrn9DSAE/OYyWX+cFjRYj
/h4A0mzmaMcQk8AGnBl940zZAI2A+ntnJCjS6ocSD3KKpHOsfCBGaBvTbthoQJyoeIDt50/MPizp
8WFOhpKBn8EOa5G7hJKJkkDjVSUX7kLDxnYQEigH0100tdzD+gIbL3LtMqueLbgBtKI21Tm1Pdca
Inowz36A2QORwGKSXtYsmf3aT+Ve6JMM6+xIUEgXJG6JsAn98BbYHCIk2znSHoXzP0pxFEwYc0pk
RdDnTykqWY+B6MJyUUrX64qK2tbiEyNukobdYO+dWSW+jx1EYhuf2fLWL9Df8+r+f/ldMO86nm7G
BWRnfohlBSIUKTBv/8b6xcsKz77+uX5IZRDuw19MnJ+2IgncMgo+6FNPESjdaAC0BAnkFYNBPfTm
eXsp+Xbi7NEBZlsfQzK/0AmYOkmk/tQ8lcTjGRsYbxtuc7DIdWTldhT5U7Pw/i7fOO/GKSLNhsw2
FCRTl0YcZ0bjAqjWyqe+Zmh1bO40mMSGDg/lWbqRTkxxzqh81JOJaiG4wU05XjAuExXo9Ezkv0XX
dK4cCQP18ako6p+9NvTYc5GuxEmhtpotIf5R0mEMrcyZi492vG0OAUkjOTBIux5HE3FDmvvcPOdJ
SXYTEX83y18dgDCEbFtnHp6njuQwrHU0uJl9oLsnJHP5WWr1ltn2qyEsaMrJzUXbghLqwz8o5R0G
VE2hDZl0fpPhIBAVxK7XBwiNNDdd8zXa1yqdpXvhcm57Idxbxgt4F6K+JNKzxLTZK+MVpndMSr4e
g6jpt4/QM04dAKLeD8Z4wnxZgU6XRXOiQtuWMAO8B1SVwIS/54WX/KW4EBjs7PxlI3ptdLX1NZAr
BHU4/M6LNUjk8x1ooxe0lC2bS54HHzGW+w/9VqHMU8bdOaORdmQfhhdJ9f2eUUqAepi5jA1G7W2i
WXuUhTZ3oyNjjzY7C326Qqgrg1UjQkbtYq4oQUssJYEwjvm2oPLdzZ9KJYhoGxURvAt+tMlf1NUu
w2r0k9cSZ1DXQ30sFGeo4FKrM1AlM8iwQFsK+xOl4gkMVOC9AusRHbFOKzfDVrYltZs8JYbtlWfv
RU04qxMkRaSwhP0vExTaiuwlzq95vG6mw81/35li9kmBUQcCjHlfMy8BV52SHw3lEKkNsf0oBX3w
nSosWN4GpzHIATQ3mNst9oRoDNkKJDs1UvWkocMCym6B+LRyNIpb/VWTc0nDy1DFBzQBJPwqHwmK
L7Dz1+wKWU6IYiuAjrcsoiJx/ppTyZC72n5Fn5I/P/kb0GlTsM25K1CLvua+MHtyU6WatCT24h9R
wvgNxkanMWqXTwCk7HZ019H01oKLeYdNqsdfJ6QvgXeGP9i8dfuM5x4R2DRGM1Ink4iCPLr+6C6K
XLdujZzzEUC3548rxRy37ySo5XqjLm17HovCAf4Okd6IWYOuOA4YY/M2n8pTrIaDrxnFCVTvwAs3
CeN3+J2z+AP2/lfn0aG+qFzAdJARCfXVfGO9nRMMNkFzUVS46lr2VrvM44l+V09AU8LgOYwLeA+3
Q69qg0P4xUiWENhELynwEboatXiq05nvLYCmIN6mtxxzuh+NdcaPUPeOrm+pqTnPLSEslZz7eLd+
0dsnMakjf1WRsTylqaVSdKITyNQSQLRG3zcoxXSAN44bAJ2tgCE/XTTJVjjf2bMH5d14X+H0+k7d
sgar49Jh7+ATvRBvMuzqN9CTxzhnLpIsgT1hAjn7vxQryXqec8KDiivlXw4Z1Lbue8vizNL3P6Sf
dUv+vZ7xzXYJvL2PhCItbqLzbUoMcyuHH3gHBi9rWpFfVyggSufzExlE65n+RSWb/V+QZFp4MoxR
lmx9QNARs4aK8KJ2hkZNo0La6PpmHQGhv8ej8QzCx2S70DiN4no/KLxcgWKZXVTYAUTugpOFODVm
rIaDoqMoDPnBT9jciJNfPZaw4fkNWvUQUcUc+0It5AN7ev67bOWJZ4lBbQF8x8QPoSeI1QrNql55
lzK9iSgHSdz4vY+n+yt3oN4K5p91zXkEm2NiuBANmIoaoDn+uAvVs+wJ59/6TfOP6tvOascjUhQ8
Pk9MKG9V+GxjA4jZOyyRHU0bUkFdujQ494S3Len0FleGLbch8AqZNXQYNNZbANnwtO59CF1zYJ5p
hj9Mi03p/h2WmQplvmaPXHw41lckuq8z0Pik2lSLJaB57YBc2nhCEKxXNzqBxm73Z7xXNqaPlmbt
KaMeaTc0z1JjkPQgUjdYLJ9C9nU3s11kEaXboJXzXV9okx6+GbkoV2fnleTfOejq7gTWxDZ4twt1
yodKbYeRF/uxblsVKgBHetEhLXzD4CU5mnxhjCsQw9kJTF1q/wmNWVX6Q/8cdQJipx+qDCiDWkBS
LerJw603pse+QGmHF68RW/ASB/R676GFlIy/WiIeyEuRoeft+0qJwTiAM6iVRJF3YbfQJx/4KG6U
5Ng47B83jfxy6NTp1SeQDztUCIeNj8sdkytKlDfJXfwT+4dhTkXmv910yvkith/oXx8gHLTBaFjf
360Zf/pMYLiB3YqhvrdZX+ZxyTWKvzu1UTGlSeSihoCnujdVUDHbjUC2fjnT1+dXbk2veEEQx9mS
KD3Y6ebQ54LN5zuaWCPz+oOxA1qZFv2H+phOD4r1w1Nz3gk8nJLRJPr9yIjZEdIaD2WmzBM9MCeA
f/i4lXo4oduAWoDw24LSnpSMPFG5M/A2iW//5aAuIrxukLNubXGwOQC5ErNGq/qd5u4c9M0WfevA
vbP8fDlxrJGyrUg8jxQk3iZkNc/dyoF6XDNQiB9uaGAYVRDc99rPe1mZSnQH2c8FT/14IufTl1zA
30IiiT4ab81KDOPKMhRs4bZiziIdCABf6gj4TmnfjduBRMbTqhg68K/Er4+sltXv2IP/hLSaD1F9
/T6keR4hXUT7MXBHwtIW0233lNnIeWskrd5zM49e/LePLIVTPtLaiNLYQImAKEcv+m8g6zA3RENS
alpGvItitu87rx0ZOqKtawe4RFnnzoFUOdU3Q1LOjdFQ0hadsZZqkwXhycMHrP+FZp9c1U+PkWzl
H6B6YjdArloCFeDVx3yiYjunpVIoBp9waQ2quRrHg4QRwC2agRS5hi/upUzNyl337mmiDQ+MWf7j
COXFRUdOdbKjBIKYEfbVeCFinc9ExbQk7YqixwP65z/4XQm63I7AYEbCgrfNc5exkaY5H3osFLg6
EoG9hIBbEB4tUH3iwVz9U3Bh9QbfuS7Cn2M3VSs672VF3Q0y+j1TaVBv8sdS+EB8f3VewEYoLknf
p/2kTDisSNR24beP6RtWXIQ+x5mvvFhmVjSlq35wMsJiLOc4utzhMfYqzySinZhqUlndxw/R3sKj
TKCxULK4SYMBYHGLYGRPDbbUeMe6zgVWyyASGG3GW5PbH4QKILVyEs0+rSpQZerCNndP2D5wXSLw
Hve8XRQiYZ/xAcpUPlOAd4/zTHNhaRjvjEpxcL5/GZsHckyjckmRm6PS3XlpCO9TFE1o1mMwOemz
Ij1aynVafjSKyUfQ8e5HuesSpaNKVBpjs/89rAFr+l1CMCdqe9kJwqKF6j8xfkDHepzbarBfNFrA
FspEmxIfYqeVqqmBJxbr9PheYZEHVK0ynhVTRyKJcDw2/g9ZLVkmTnv35sWTQ66UNIbScP8L/cld
xAbaoo6bHDRZOReTm2k2kioXZuA+6ssCbEtXqvgBpr9R4Lvaml+TDtfG+A2hRuUCvrxMu4qheOUA
h7wjhfyGYQaduBob2rYc5zyST9MsEyLuDSJ2yqOup0bnPiptNCqz2QYl9BiMSJ9yrbzJJ8WLfQHw
wJ+GOW4Qv13ImzIhVuAANdzwHRpqcAJQuw2MmCerTqVtUjEQUltXugkriAaREMDOe6tcWXi5dwFz
K6Zz9qUvaKbhWCrZqk92tgslAMF8TzOGAeOumfV2wMEkJJbLV8JdM/vnfDtYrQbvzY3eSlkj8foG
IGu0sS5A83N+BmaIrua86YxOm6NuoDZZt3/6DwPvXoPyJ1hhQQA/UbXS2MMtfcZkQzFCIS0Utgqd
hKyfH1hCxgwKia65E5+bMi+a59xdCrG8lsuNpBMI0QTXlvOATFxvMaSOpRfMe9KrPP5t0Eh/FAZj
PNhPzVq54KeEgwRR69I2QmEIv0tNAFbz2zHFAmrJM2Q6BXYzZ3YLe4FUxizx3n1tA6OmVREknMK8
MoW461smU1F53NYdewV9GnZh7onmUfImxDb1kaL8CPgGB3JiAwB2toT/LKIlwi6bBOAdSa4zXKC2
spkJuULEnoOmJWcQxrDI3omId8tSmioCCAT+J6LlADvztB/jDGqxu2Oy5a341dbog2D7afK3CLaQ
o2Va15xFV+MNIaRCFMSQajJ1qc6WXYgUdphcwXBOIdL34DAAVuTYHHRpc3TuUXOpVplS6WT6PDic
PLhCPJu6x8+dmPSIk4DPaEwcUvb3u/Fklp/8siXs9eEOjXf4IXEnKrrmGzxihoZHmPWkSSNXUSOt
hTG74u4WBJFRYhFZH59dWohpjaBr2wp+sJRkjm6iG7IOyQGNeJBQFLfRPyXmToEGI7t6rLw+/uB5
mtvPnygf6EhtLUNna2DiG+YxS0f87+HvZR7ZBWkYRMiHWVVd/PZUy9VosJwZSNxvTQWsMTaK3/3K
nvbi2iU/a7Ad28lE+bSN2jD9gCk/Tz5QPbIBnomcHySQrFLU+iFEo/Qke+FBnBAeqmhkXaDNpZI2
ejuXtlCWtKDp9OX135Ry5vouOsbMeNbwnPdig12winME23/SmM0nQDK1bRDFg3IXqLHPz6MDZadO
lw3MWq95wNeVSobmkSxDBWgrfa0ojXXhRcocBHo/FwCc653Eck2iIXRuHDKrF+kHWn7wafoy+pXb
bNnOg3F4NcLe1UtGi8WCwsxOE1qhZ+58awDVt+INZ/kTxF2OU16xxx5ObBWljuBU62XSnF/jZdPX
74FhoM36z+HLtEWYD+tSm3YO9m7qh2/VaQ8B9dbYv4IryQ+eUcS/CtPZlzaQWms+dZZ8BWeGfjNg
q1+CSvMf/owOeSs2uma16s+wgokNwXEHpdB0mm7FnLRf4LxesAzmkuNQcm47mgyZhlBru0jyMXQu
mNCva9mXptboRKJKyGlHzsHRzpLSZffKJysjb2z4zh5j0dOuhuXWsZcwPjD+67avP0nwukoV+AFR
GJsbqIgw84WJ3o/Gncp7QY05ETBhOn6XwJMNwzYFKTZPBSV/IGmWjoGckR99MAmk0CbkQAQvWxsC
3dRqcjbqDHMHixNq+btYApPYi+LPjF73OD0JJ6E6MiSOcWauzmES3NatDqr0TkUy2cLpHOumb5Tj
PhLbTmpOXakX42WD9mrJxW/QeknQK+omc/LM1NbrFPMobBTTB6Y7Rd/GUkFZxAxOoSvJ0k9G5rAT
YqvwED6bvYhCa4L413RoC48Jv0IBeXcZUhSeXqCHj7OcQdBDjFR//VRlawA4xbu8WIdrwaPsb2g9
FZoeJPuxe2KMZU3pKEEhsEs0f0Z0uGEdC5DLjv1J3Fw04pMmTN8j1MAgKPTZ32/gaRrtwHgW4Qta
AslSYjyLwtq5ujuLYSljJwuO6DHH2Cvu/a/LNN1/f7Lnv3f4mx/VJOPNOSAFDamymNcUkhBsbP3F
1kADro+/WtA9Y0JEH4A9TNmlc7iCKVprU5cE6/cGdEXYrJAgn08kF2JSV+IsGSxaH37EB53V6xKk
vc6Fff1Ci8itIc89ZWE/4Vcni73XMSM7V+VPG1dGqdtnvpY8mNJeL55CHJLS4aLQ5ncp06xYpZIW
i7RpAZ5qb0JB/sQAckOoSRMgn0n/mM0Ehm7CjEs9qz95iutWeAeP13H5CnCPQknSdzsP/MSVEcNA
2bX86DuidqqfuviZQq+jE6TinTY6/LD49D1uK1oTVC3PAJj0GYqdCLeaWkmSMNbsREqABQR2KlwF
kZqb8Ab15fmA0HYo35INI83RhCrfrVBUVgQ3YxGMCm5q0q2pFkUJGpBUkPByRd5WRwonU+LMFKpq
dFzp2o0UC/bMzDAV4yv4u86KZ2GDmqUET7sIAZKK+LZtcpeaQltOy+3MzQASAGsQuW1zaNpPeLfI
x5j1uK28wcUlcvqgK73EsZcUXiYfeCA5qZZgRScH4w6LQGGwZi0bhgDWo77ymEhx8gvCCsMuo9Qr
HonR8i/uX5C0jKhBMvnP95m9Z1t5e/zgB5fSvO00BK3Wb2YYgehtccK5m+tjgNIG7N+COFT4TdAQ
dUKtr6rlmEgYpdfX1jws5r6BHOzud2va8mOQ9sVasa+DGhQmCLK0ndwi++rFkJBG+UqrVscs1RYP
TdIhr73/1npkyEEy2pC5tlstCUTL+7IDaw2W3H1IGigG1WSfOymc2PSA1ftQwJHLPljk7MTW6Oly
3JUqvoAjaMnwHQtKVklhE6qcvSpZt8nKAhnqhnr5Ft+Y6h9sANWGB4n0K3O8C+WPPF7Qf3Ukk8mH
jNSw2vOdLLFz57TQI1ibmYphygLbXss0rNa/a6DIcc0SrzxpLIVmf+2IQCCvh1YSPgEInH5OCZtI
lCJmaRbePAq9if59MDWVIABWTb9hJWihhF6r8IkFVPkStKNBx1z2pdzS7DJeSOJWkL9qiRIjpvFi
GwYCU/74aj21neavuZbjf/DjVdIfbQyx3k9A1xBRM8G5Iw7Hi0pfm8vfsu9g44ELEHKtogsjmPLL
udygHQotqW2phFGYJf+tLaL2ZjK1sWKTjU3rsxEsOqRtf0YuExQ2BS495nH8KGlFcYfqgH21X5GV
ZFs8kq7nh8gwWyF6nL1JRAm1t5YpKiIZtSsOgc2Gx1F4uNXnZdvzliOqb4BF5cQDrbD//7eEQOgL
vIDaEOy9lyKamFEDXd6LMSEPeCO5pMt1s/4E2Rc06sD6J77SesYt09B1BH/gOGMd5WG23Qy4ZEf/
7MXbgc3cK9WcZlSTso58XUFTlK/P7xXiVdQgBs7Uz+/EJVjQe0l32Ry4EfoJ6E0fUaIXH8MzybgJ
2K+M5rHyNiNLlpICxn4dXhftLyJL0zDerNxSLMHwLRTXImgGW88A5582af1ztLHwgKIe+z7oFYdM
hG+zZLsHSL5LcYd52A/aJu/WPTA33F9Gubr00BgUbxIDeVq/4n2SzwjhzZOOpo1luZfySJH8atbX
LKuWR9TTmgBRr081y/0OwmJO0sO3/gcF/dIsvTxVpuiTdnuz884kOJOdK+76gewf7God8gVPBgSL
G4n8aX9V3Cj7x+u8e5PNpebHLG/xNp5dQ66/V5TJt2yzmT/60e3Vdxan3xCknTzq7s2apPInf/5F
3IPoYcpudpPJVevWfQx8OGpDhOgVLUSNns5Ar+lL3wBDlCCZerl09KdnQzMg1G2x0/VI9v1GUbT8
tBWsCL41/Cqg8aiHSjLWMWhy1c40wp/aNe7K9+AyTkRL+2yY/K+InRYbPIhx/kEfYBj/vHsdBTzT
8CjvuStvlhilgEG4EG7b98CuNzrdmtX4nPkb1qzxsh9nPCwJrzpEjTD6aOlAzBhR9Q2X53qoCDrx
l3PNvty2P8v13+O14sPnPtoR/JehcC3nskr+mCRafcaW3huhf97kQwjdnZqtQPHpwJAFW9ELq75u
sLlmCqFleUVEQvV91Zv9Hzy/CPb3HF1OUGqKT2JgCcrC7mEu+3yc3MXTJ7imDKxSaYQ20JTTFU+8
Bo8xkrjFAKLqRiYfKn4825a1pyOwgvf2PuyXQt+FxF3OZ4G/wSO91kvcs43+5/G0cKzdwlJPHyxT
JuF1JmTfPVtBM+ct2WF7YT8kN15KTwq20NPNZJDWABB7AleD7f5h+ysqaHsNGMIyPuMmJOB0eYfz
jHfPaxhdIXFEQiiq33cX66UibouI+99pp+Vz+GSCoNETUWI9CWMJD7eWf4QTOaa1kvjPhzooyKf7
zrQNmV9ZbpLzmlOD+o8L2KkYkOo65vTj/FyIOUXiKsob6fhzEC+FKWU2zDwTor3r8zZWSMW+f37p
trI8Zgf32Y+0TjAAgKDFeUWhnVyIQVXdYsgiLQUeIJ00czgIhYwfyEwDLCHiyy1ZiIJo7Y9WWsfL
mXbRFODCpgfEpPlE6NLuH96Chq0YHBQ1+YLpe86AyMZFkdg7M7SUiM4Cpip0Cz6iH6QomXQe11Th
k65r2cwz51oFqvTVdmIP6xRunOUNoQoF187NOxoNCu/0THNHi0QyRtK2N2ot+S/L3yMKptdGNl5K
iMA4ZmJfTZLqR2zCIiBXHPUVXy1WbPnbMkz2sIs/0u/6v6j8+wpv7Is+aemuStF4yic7V6cPncdL
0sAUo1oC6MK/ByjQQ6uHth3AQ3WDA30xXfXXfiM6DjvFfnuu1S6ud5pxgqrqJ6B/6XaKQTZ2Gofb
75aRvrONxfUQeYi58cLfs5JRNyKFLUYGjeMesdLqiHJazRwqx2ALnQnklYk557vIGgyaCJ8Mjzjs
c72mOHLWF8rfJuI1jr1oDyN0+o0Y7TScQPLxJxzVi5gIY9zvIWNs0eE0FtynfwlnICiI8Th65rW+
XqR7MnGxsgsGy1T5Md6zBLjLaDd3nRjEFZFlvnCZmOvBOXauYi1ySoLDD8JfMOYqDexb3UPnogsC
vGZ3LYKWiC5iglMx64434YGj3oICzPtiGzbnY9lbnaiz6qg8msqkC5ldPGHuOJwiPnZVP4KEXqZU
6pabNEMB6EwVnHbR1Xx3QNsbJA3UCHzWmtZ+r9co63bl1c/4uGOcCarNga04Zc5odlVgfbB0T/uZ
fuA3DPSFR/1AVNeIVYX11+9X7ycSwgfMBTq+Kx8pjVcvjPINrNzse+j0aKZnmysWTaxGy/rV7bR6
X+gNXkITTr3l3MqTtu3Vd45CtLY+E3NbyLlGRdnNXtrTBV4Dl/Nn5bV9EWP40RSIFvmsvs1VnFKB
TNjslRs8wIZd58f6/Yve7PbZ5Sc846SO15Cnca9hVEivO8k4z5CmRe4sLyMmaQBYyD5Xfxafn6AT
S0858ueLvM7fuXK8sbvim1cjwLcZjqu/K2IeBh+fw0HbuQKhMrznVe6sPs5hxph+fEqmbJAe672K
ivuV4NhirsyhlBXtr9vbS6YHQJ5X5p3TIygphedLPuuwcY73CyCKbsZXWTJwUcgcyjYR7x/JQB/E
tBrMmpOj39uwHfwrwLAvnch5MCfDPeJpX8nw+BwifIvGswX1+iyeLJFPjAtQZrLkvh7/tnUvboRT
HUV7CdWf/WukL1xpJxnmsemwJbpG76qDdnJ//1QoAMlpmEaaZFyyWwQ10EAY0eDj+4jh+3PNN0E6
Zy4y416KfTgNhBLdhK/DCO0QfB3MpWOnlX+NuGCPy6/smAZ+d++sIEnHoZ4Lr1ykw77hblUiekZa
SqmcJgZgdJJbjsuEeBMBqB9NwdGf9Shb46YgCkFeZWK/zQDMAEyfnZWJmPIh2wZr29ebcHNQ+v3A
GKxbR9zzLDgYN/pmIZmkTFBNNyQ+0qQDgZdugGyBHxc8gL1q+GIYsa2DY+TAeAdd+YHd0pukbF/q
ZYO3YYugBrBGXGwEhwOiYPhN4WQkg526UQYVqbyAJk16WS+hdbfDx6qsw9MQurCQQA/2blS5UQr5
1/GmwOyUNR8Mc3+5IR6FCLdiBjGq30yECepnIFKhao1DSyVMKzwuHu5cdl8vvCD6R/TrLpFKLs1L
sBG4vdI7XaXDf/O5SLdBecHZCGGskW/D3+vULvQwjYT7/iuUL0jmcOPxgIkx/jUIPdMzv96S6jSY
8kyTGUJAl92qLBb2Hfe1c9IjpJjlPtwLTC3F324pyLv5NMoyaP5UtVK0yVdKlfKQd1oLhLAfv9Dh
cDSCJffgjCkgjrS2fDEtHWAlfeGjlwBSy96/KJJPiKQuBXItdIgoPxIbFe07jCAA/po8Wno+kASF
6MFSfAlKKzqCWFunFxFRHGc1RgJ1bLoLg17QBKgl9r9iBwxUGgKUENMAHHTVJsL9KmYkrnM9iwQO
FYwMBWeTnlRYVrUbbt3dlOD9ZwZYLK+K3swX0lvIhIUe+2OuZbxC+0hTsdF1Z5uFF+1kkZWut6XB
S+BAlr6E5zot3yZv51NLwoRyoKtWGsCvzYboRg5bwIbY3SbKnBFglYiqZaNnrVlnKGqXuFI6soTm
6m6U4NUDySTQ+YWN83pG2XGcZZbvBjC48I/gRSDuAG8eSUDyfjkdIRmnuZjGTzyXpu+8wel6deD8
vGFBwQz/BlroOJCVNOxzSwe7/jELtOTxzWgnEvmXylr2ggVx/2y9TGHpEKqgfaU4DIdv6hQFppM1
RVyhN9LjrGmIClQABD4YFClqmo0+AeLtpTsPLeEPy7+L3bZLY/tmTLtwK0Qepapd8y0x1KcuDVcY
0pH+wHDw3LgpR1+K7zE5qbUgJVs2wOzg/jkNrN6q7FYJcjRQU2nz0eoDL9MzE4hfHvhxNdb1XnbA
C8cWONJILC7jwdZfolDa8rU0stX6aknVxdkYu8DIot3zlTDszzr9NtbFzFGrYWIolIazHl58ByLi
egu4A2SO6iMrOc0p8OZW+qz48j4n9Wmid8uArD2NK4jTy/LzB8w7fbyD8XffSzwpBdMzkTvzxVwf
/cN1qF6799rgO4TZc9yf34DW3E0pRfjhKYbTq2908lH/4JXDVws5gspjh6FcOfwVUTOxGYrA0Ggi
KV7ObRhVUm3Lp2uwpKosaeUFf32BRr2fw5H9bTWyGOBIJOjHR/nVikd6ob/CjKIqCf45h7eYtUNy
dbDZyc4GFNyoYcLIFWrT+ZEmFvTBhOLe9PlGk2gddpREqneQRvVpqvICG1ESj0L4SsD5JXMpNC0F
DqtfAiG11Anhz1Jb1AW7ZPtsbukr7ZGjsWpZXSfWbm3KjwujnGjyN8VjtCdjERh72jO1ZIhAzmby
UjN+087xSWYtg6H/TY3mK0fQsQrMOS0gu89e8Zpjia+XYB4sFFhWBhK4pFlhphmI9AELjpl45R9I
9IPVs3/akvjRu4cbUQ7cm0QUEJGyc7kloIkedK58lL3QEhgA5tDjZX3CsDaRjB3dH5ga1oDDUXtc
CYDZVEKtXShtdTAU0UMnHV7tGfKHjsFAbLi05FCGvhAZlGluTpYh51whH+hAIkUiNjM3UHPgrnia
FCYiok0UywN1oqtwJpeL9OxjCM3ALJ7cEjFxjI3kLEPks4CzTYQv3Iimc6H1tYmQ8fEZy+91qBny
D7Zy/j9hKkl93l8Cj+LvcWSaHECHDZYGQrCifsdsNGCFHc6nZ83vzhcOl+TTjM1g5BCpmz0gUJ+2
J5j/1cy27h9UAncy1L0bo7W/+qs18NwyqnIvxhgNfLh+w0tqYPdUywo3HBNxTwNPfvzW6VHUdcQ4
3xBtnspuWbCMayZxr7uJvNjdzXkGVdYksdOVEsvBVzhO77UEWmjEJb174ag/LYGaPYembA2zkZyH
ZdmGmLGbnqcuHq/vcSVFh3nALzkq9xNq25U4MThme7cUu7bAGjZw9Z1DcOKcrykUSQTCUhptdlap
wdvdbKAmAFKJUvzEli8eOab/DXdFzeIiFiwsfJAHXNHdDFlSwMEG53erLhyd+QDVsYJLZ7CJgoti
WvZTbiA8A9Z8pmFvSvnRqX8P9rVeHyMN49wRPbm2nB+SRvzkyNIKKnvsCSTHSSoDyNtHL+1EaNJV
nr3z3HxCyRnoidAfcWX23Uf/Co1m7dea2RmK8fKs77sfefhuEKMFEc9jlr/IY23PdcUHsA0y/MQy
l3yxMnFsLAjWUpEOorhqjpjIzGKlipnJ+qPzCZiYpWAciNc8zmbYAKh0XOAOUO4miDrsDIikq0Ox
IrPKfFfjAghtlyVmMEem5TnBRe6kM24P98vj8n2Z/vXf08z/yiBmMl1Cp9ee4dalFjfPUuWZblg9
F9ni1PUztfvjubnbtv7wGYZwxwvWPw+th+K9vV1oA3lKMF0O2FBTr3IqIBwILDltV9TD6EaaTPdK
VsSlwnwbkumFDWD3NTI6rE8fJlJG1E6bvPyJ8GeEYwnwr4I+vED4mLEa7QDaEGFNNg4xlJl3+/tl
G+P8SqPX/bVbRRNpjZ4oU1dyfgfTQ2729V4nuSrT2nqS56w1J9kmm5wxinu+Umg+xGaZoi++Wn3Q
eZMePF0EtIiAhXNxHqkqXS5+nDeIwJ0gn99BIGUSow9CkhV2b+2w6ZsqwQKpKIvgIQzqMO2QuYBS
npdWOJvrQR2WmFhgnWtnvRHqvbq4GBeFQDaZZ7/xrzmAIJJVti2n3JwRMRSktCxiXHNQ3kkgzm3X
4bkTpr7CdYvbVwbeUpvRMlMkfu/yWgzy553URg4xXjJ6vdR8Tm7Zk1EEfhgtu0ybY0tRTujaiOh2
Lb5CJRKDZXVE/tKumrxdbvzzTKm+XOCOBOTs6/3ZPmTyuquSD7ZXA68WVgdfTgpamJIIVtQ2anXQ
P78L1VkO6j8YUiqv/AFKsof88AEb/bAUKvcE8XzIO5/OCY4FsyLL6vN/cA+s/H8Cd8Zbuc0K4YkQ
uenoVBfUU7iD1WMmbmwrc5BHrj2Xnd7ovjF3zV6BKIhMVRtdqsIHuoJzDmN4tQ+7IOlr86jyaF3P
i0v7GlnV1kQRmzbXPO8T6SrfkxbfKvIgAr3+GAzMfbSKGyCLGnJk67SsjeOHuE2DzSpL6om5x/i8
+Sz69wdNcL0KJUay7PZTG0G2y/+iL6KqBLLmJw59bf4UeefAGdxdTcp2gLNfHCnVw6k4CzT9I4PK
h+TfqUdyYNPgba3wp2YDVXu7+uqvaTWBo6iTiZHimIuJuioLXMprENna9qvJUf+EYmUu0pQV8gDO
HwwQi/5xQ6iqvdfvNk3dXKlsYLJJaXgu/zruid0CDCUYI7bouqwUjR9U+I6h+tUUpGvHt+Gkhl1V
ePa92MCxfO2BHE9z5K5ipe7ymO9m14JraKQ4Dt8DXC3pWon3TBmgHDG4u9HC5D9d6iAryONwdMlb
D5iPgFEHEXQ316xjH10Bie0b8XNVXUfAGD2um4KQho5f8oHNTfZepqTWdcw/FNWcZbK6u8P93djr
/VDcLPX8vil1g3UvIwia27ELImTa/X9vyt67wG+sNDGYm9AwKU7v7uqFhhyQjpvBiuz5Hx6/RTT2
qxo5vR/Wgx/p+vTbZuaEnDr57kablG0BCEVzQ8Webk3PBK50V0kvqau/kUvOnpYz6ttqemOvea8w
wVGAUcphe+kBvJiNAa625UwP0dfzvEPK9GX9ENxQYfRsa030Kwj7RWe846P1R5X3sGzw7gF0Txt+
SupG8ovxYCKbpdxImygWJtW8JVG/FMVHDQy4YHxO5rwOYjLBhkaKcZXb8k/6enw8814AIlGBoZA2
mtJ4BNYIWSngtQvCtnOJ4AcfXVqWg/G99NbTFmFGgOh8mInleCC6oq0OEsfck0LoZKizlY1gShLi
l5pHAdsNetFhhhTeS4xAX4/1xBY8DQtBERpVx1Mm697xCat4lkyWKYzS+77jDv/yAr2lBivUwAZQ
vzEiELtsSfld0B9brC3NcAgNSrNFJ4yMKoo9ezkL7T/E6+WS9FWLE8fYOQ/suXlJMbSv93cLZt6c
JfJe5/Gs2alXnEiqxCQxuyXbktkaFCtj4FdRvRzeGHoTGDqUvNI3RR7n5jTkPg690rABL5QKj7Ug
hJzz5Tdua0YNjKejso5w09vdHXVa2aTJ/9ZjscPuD7+mu7fpGXBrngdxprVMuxWxtufgCD28T3B6
jJ8frXCxK0QNd8+rhAULNK19VCxqZmQfDQoNqxqnDUJWdjrnrMMldCzTHsGABpcLCJFarGa+DNnI
O/XhahY/U9XCO9oJ6T3aJHNd87tutpkGrq0c/n3htZSNV8VhMbFIB3nagAKvl06wnaBA1vmMQrAQ
fNuIe9lODV4yUqwLZIioN4jo1hcMweeeFj0JHVwWOdKZUzJRkd4ZxW+8eqHS9WvNcara3nA7PBZf
jIgOLl7CZy4zpUZ6OOmsGG/Ro75XVgbojcKQ/9nAoxSEqNHLDDt/UbAJk9UodOMRyZ4OiOldWkSY
aUimal+zUFDauBqN2ulrudnq/F3PLst24uv55y0RBZcwWP5wVASx39UbzeViFXK/VVs+VyADSx8h
h9TgUprAl7cVpRv7p9V+TeGTRFk4eV95eDhx1d7EYJ69YO3RNoJyunzpfULNMqNxk2/o5tHECf2Z
PNRsHJ7qfLMEAgThV4mZ8uvqS1xSTYZDtynZPd3LG2HYpTcr1U6s+m6B/I4x2jWWrIVJzQNdqYG3
r2DUg8unKhcuXHxM4KT9wos+aHtNOd3xFhbAJAocSQWoS1JduG3YowQ6V0pwKaXWYprIHQHzAGN5
HfyNCAbzKqfTH5p1bucwPjMS5djZafH2f3GAzL+ka09vNAVSmQuTwjeUU868HSXdhetX0iWo890l
5hmuTUYhdcosLD1qPtq9yOkRJat0BbjSEMsmmdGtz+OxzzucSfJMdpcNlUwlzDm4JpiC4eG5aSC6
mFEB6J1hXztC4t1g0mOYT1FJJ5hgNU/hDVIr0S17xddZBPgMnLvGJlzizTRKA71MBcByxsgZaG5h
f23gjTYqNlC0WtA6sosJmvaWh6ltwMdLe5LThbC23tzC1atVJbQTCVzo6SJLd2I9sKaBfECIk/ZJ
DqgS1tSlXw+lt5BdW6M8GtDfVr9Qx0IHNdfWrgy85/NRM43xnT3nt46dxGdw5zxua2B7mWMigqj8
+m21iQF2RQ8al8LZsfHu6FPueb+biojVCYLIN8vndTSNX3asZNpCFgr7m2UvMUqWYckylAV30E/5
QznNHaaheHo+sPzQEJ4TGSYqWGSdHTTdtWnu8kZ4CPyezp5UgOp/ZI/TCExu0q9vEB1UUdG2YKJ0
OmHUM5sgg9U8Yk5Po0K5nq6b+UKggDQgQqT5GAbirlanUnkMBE469xvkXK/L93HA0LrfbqHD5oB0
fvBiK2B53/3shlu9hzHb8oXwVYvJaLsImZAj1l5JIKIFOKcBuVdItyaJXZ9BwpzT17OBQeEqt5KM
iw8/KnJDIbcbJjYzNW7dghKwtjI0161PFvlgKDpGDFAnmdgQB/k77v+kTuhxtqGVxPFd1A6XK7en
7hyNkf21vk/RzvOD06ZszVL4L6BfcNdTi8Vrq33Lsq8uAOpqVD6hYsd/8mYyscQohE5g0FbbtdWS
wbNSCaAeaOCh+MRkb06209oZY46JCQsdOYF6BriFXxaOb2xfRrmIE7CJJk1AOqjnHVN9S55ch4x6
VQdeUiktbbaKfeqLmp1aPnnG35E2c5skmp4OhiHd0VcFg/1Bxk2UH2tE64r8rSNmY6ozdVKuu0yF
gxynEMViz7U4qoowbbVhFqPD8a9VIaMnu0PN8QxLDyXDI8L730lIFksUgzl9y2oU5Q/qd0tXy7fT
MXbLGuB9Ggc6iSdg30Vq3fv3S/qCM5jp8gvESE2ag/1HPp00BEQCC007OUOZR3YZxeDNMtXnPTM0
1MswMZjpTRyh7tZzDbYl46WC0iaIqsTZF5fBEqQyBr8QpLIinLN0HOaZ7gopZW/eutvc+Ho0+O/L
dH5vMOj0I4BXiA0iaEUp7wpSi9Dewp9gCBTdxukCjOtgY4TFwqOYfHx4A6A+Rc+2bSLkzGvSv7rb
5QqFL2bq7eNy7KCgnPVlS9QnFofDb8Qburrfp+zerZylbti9PPXAX7zse0zMX+xaKH8DSNz1zPth
is73My4XUPnkpd3hCPo7liM3d04rvkgXPQX6uaMwy8ufAhtLFO2lLQ7aN8VUdUsYLKX+/zfL/A4Z
pUPtSGCb/4IzlE94ehQ4k2W7SG4MmH1To3FYyArDxREFmA+amuLll1h+FBxtnS6mfQEymW0Y8DNh
bYHc/ATx3JI5ghGeJ9zgpC80fr1Fzyei2v2aVlvB+WZzCp+J7mtTkGq3N8EI4Mrdm1Z7clG5g5rJ
QOeD4LV0DED+eOeAhss+rE+QoxhHzhq+EpCYY+epCIfKFTMRA5QMh8knbTBuxDd++tfhwkh36Hnu
y1DAWXTGJ4/dKguMK+C034iI455MuY1c1YsvNJKq6uCLrnhjd0reTJ8CBrHhBnmaiKZ2/MNr1pWF
xPVZpGiOvO8g8aEkKVrWUW6yk12gU/yrnzIpWi7hCEPjhGWyOkgYlgwJJ5j+G/yPIbleL4xZvi5W
Gvbf/3wGSA3SPFAB58/C3YmlFW34XOTf9Ktv/ddVOa5vV8JSwKJQXHA7khPBclXlS/p3DllZn3Pf
ph3gmQe1JDKNs8XjZ0BbhYdvtTLbG4VItYfYqhFOSbwQoMQjZlss7/nEYeyNiFF25QUVPE7+4/OX
Mjyq/Mp+jUXXEopjpWZvWs/S/1+hfMX1u9SPuF4GGFPz6nCaIWrmnjwZo6vyActvvJM1UYAgqg0K
XB4m/jG10YRNVZtU9h1KikMrq++UngsUK0jWfcGjMzSZo1uzfLzIke/8Kuhda4j2FQN5bOnAjSHW
3ixnYQL3wMcEWNplJ4umDBHo+g3ediw/SHV9vqUNdNX6CtBBxcs9aMzjJhxvFZ9nmLmV+Is7fQHp
OoNDIxP1GoDNwd2KPu/ClemyMBhrefR1804RU/pqLbK0exGJSIRR4lA4EgOMO1f/zq5phGT9uQay
80xjjrGycCDaIPzxhGgCtoWF/EEzNMGZCFGnkutZmlxnF7NtNzRXq2KqobdXAchPxz5/JrtSsM9A
CqxAdbEKd94ybBl2NUSfEPQ/pNw1ncka5aLPn+z7yCciXwGWDVZ0tlkfKFvEkFvLwPL3GNf4j5IM
B766nz+k/epYnyJedU1u6O3NrDQ2zY36rtiH8UT09QWWUMXXYQu5ZbaRMJ2GnrIKOcAYgUDy9pCA
VzXASSNOfTzlCdX1P6gf5U6iP/sPP5j1KLz+kTI3OibUMPP4lNMwSestWlWvkuDEjmIcTVXi7ero
9jMqHyVWSdRh5vBfLhrpvDM5PSSHKFp6xKwYc6MLrk0NC8VyTrCrm1hXPeDwfW4NneGqGEKh2qlw
itBOlGj0vIF5ecRlTgtbBQb5Sv6EaKsoD8xQzRWfiTF+d1ITnntu3dX2GyZJO83qBwMThSomTtQi
9u7DqF2lfhBSqW3lsULMlv9NZsi3hylO6iOVdi/YfhIOCeiWG++UQkCgJxvOZsnZf8qD3EyE2K8i
AA6l/k6cAQ29cAdoHuTiXR5ONFQ0BgzVPUYaIW1EDaBgdMNJ1kUViHttbFW9ahXip723CWrI/57j
aifzLbB57AoLhpSjm+n5usuNfcduKBjPNc+a2vi+wBGf1HPrmPJhtNLPOJE92ZB2wrl2Nmh8YfTm
Wlwjfq7VZAc4pJZhW4CvR/vXVmpaGIkcTDBStFX6n55dG3AK5/G5xRnIgUP29GTqKR88BVnHV/cV
zDQSdqLPJ/Oj5xn+zSAsT6w+35I2+jl0TPHimsBE5ieaadj1JrlLKGwBYaJJMrXZ8OoG35FQjXdY
Nc+ljiVxqmKebqcE8hpFpB4+VgHGM42ehWKW7KbJPodq1Hdp1wOQK5nap1Dh2quDN4CQDPcOt6Qg
sy74bWw3LuEEtH6o267bVAGm0xWQ0e+j8DhxIoWQ4jqSp5grrLwmKG1lC3AYpNsoknf8HgsVLeLM
7njZH4VV0DRY5VO+dOfMVFBnNZOr4Vb3Sc2qSNgrdlE4tjHVWAYlJDyEbWNXbmHNbp+GX0Asenkg
bykW12k1aEguazp3NrHlo5UR9zkSlAsfDBaGTyRu9HaCTOBvJ3HoLcRVrEutD9xFFEBDQmA6HYLp
h5J9QgWcJGs40IOJvEJO5D6h/buLbK6OtZxAt4BjRbvLv5ICPmIZHDLA93jFoi+ymsK8c5TYiLSt
n1S6I1Jb6jjhGjzs4rXT6eR3GZprF9wAGIgRq8liLxg7HsQtnavJpk3JTdJl6/u1jMOImdKdizQX
xLGqmyr2b/N8nSrRzMBBgxf1Dkn3DgQbay0MPOqVk1pzv3m0Epni6Wz+HugWSOj3+HAUcBoYbKvs
dt3SWX7hG0TyZxgfVZ18lCTnaIVVRk1wAErc2faTXx/XFCZ5Pal3V8KkHepf36kAzpoW9QS8+xgC
FhYrRpGxK54Pq3796tKd7eKq7J+aYVqmI6+vfPUvvBUqhdfJfIp0ry7ur6Z7Rp0fOY/4GM86MZUx
2lPWgevuZ4ceQnVO+NTZeva5Fai1AIjX0L4wCctBwSTkeTyb7BtpaTLmO9mBsI5ZknUfvv6PiL4+
hIwj9etaCyNKKsd0gY/+XBEi5Q1U1BjVf2x8TmkF5VYPN5v4yPsGutrIpTaRR9Ox52V/cF+RB4du
9Zn+twxWu7WLScENGGVz6cXXjRoYMXw0M11QTehMHOCmI24sH4lXoylxvZiuZluMniWCUbzfKLNx
Jvq6B0gg8r3BZDYZCEBYjjiPsPmdkIF5kfi7RZN0ZeKrEjjxaL/M/8qzv50ryydULzmEe9zJdwef
nAdv4u/6QiZ8EHul+A7uu35J8WXSC/8o3XlvNgOBehUsiYB1cd6TzalJkmhdrRtw3wJ3LbXHGbAV
oPj4GoAcaTBxFJQ8YxYgz6CVwPwF3Gje17TcdAfCarwVur9PTd6BtEJh2kkCUEhNvwcfpU2JFZqU
XG1PbjqYpK9UCHsBDqK/0Uxg7WtPm8/w5d+rP/+mIoFBkA67sQ/NQNtinC6hnld7noiPdWy8P0LK
y/x5fS4jX651g/7iq7HRUT4mdwEUmg7lLDh2TDabtOxQxgaxP6LmJXhoOLWgpQBGchoXVdA52en9
Lm4wrn/7IJsNTmmNQ3TC8mjyPH/7VounuyQ2VT78VNTqcwA7U88OKvu1Zr/yZdgz3HgV8TfG3sYK
Gp3BKiVgujdvPJwivE51tuAyjV7slkNT1OZfDOH92ZFX7mTo8H+tWKpIcYyzTh0Pt23ZxQ06rfDG
CLpVAK0huB4CZJGuWRvdAsni58+2qViwkDYtwytPVqM0609zY/Y2KDethrsZNcowYu5p141HAV2l
wR6ER6YN9Kj5d8p14y0htVH5OMT1oLt1g6xR8IASnXBt/J+h4y1UnUoBthaIdiIE64i3mf7RFZYd
MwCMPega2fxzqgcS/qSLs6fdWKk6JG2SVFGOpgk23rBENgyWt1C2GRvcwsnXGHAmS1VLDEJp2Y1W
8xLiN9lBuGd7/4A1m8pdgT8IIWJPgFPDRK+uUiYHyQaY45yFHfAq6A4Fu5Itr8eVcAlbag1R3iqO
LUM4F3TOUtW/xzqi1Rb+FiNkVzvIOrABTg1KG5bGywlN78WVfFviHjDa5oypIIpjyJHoMGqP6tRg
nG5HYzb1rJgtsyJBN64jrNgX3EfvcD/vZX58A5b5j6Ukw1229w2IC14JdXAoK21vSZpjMtsH82SQ
R5JddOTdBdQU0bJ4ZFXr13RHNXvCeZ3Bm1wnDxWsFmIqYdrxPUIlOQf6roKOZHJg8OULgNVNHmJl
6QJnuVuj3ftKgRiWp3gYrjkT0qi8L/FGqrfpDcwWlNs2RwMI5VEZH/+LPq1QExdCNV2yhVgl5EeQ
3Ed0fJmxjo5oL0eiIdD4zJ6EkkRXDg6uvimEc1PW91vmHPheZ3Hwovrd7K5ziVBan9pO3YFlbhen
4CVQAM9DhUrZyefc6r5+f3f9ekfjN7nFieNn4tK6VTltCQpXK8O5XEJI31lY0eE591FnCuLS8chX
ENJgtqlkjX/RAzHUz/aKDm1al0H75oS5nqAEdN7WrkhYvP5HB18wm4+ckSwcx9fXzLD8Ehf7qij7
ECzLu4qeJgi0BB7X+qChcmlx+4x2QyPzkRm8H78dEex4SvzWUOywRPrTwUNtsHyOv2bDSgok1k5S
sHq2wvuHPck5NP+zlL4hJmNyzzMP4wtTMJ8eO7ilGyH8NUOVjFfCtyMr7GKth791x8McEwHHfh/b
J7b0dGuG30vC+G3/DnWvrCHIYUsFeWiwavZzfuC4/wsqAqP8ZURtnnPhzxClo3C85MTMO4G61RJ+
B2lCdSnJqG8LYKHA6t7XU8mvy1NHf+8MF+BHBJhPV204sFEkIAbNGlJCVCvudbvcl8htND8jcvbt
9v127YReqeEodDjV1Zckp4X6PYf9VTOuvg7dlpraExkcupVIl7DIpwifL1XG4jvxnkkM76YiPUWJ
f2s5DTHb5T5XkbA5IQGW9r8Y/VWUYt/vtDB7yMRLCAuNTYtl5n2BSUF3s7JJT1ZycLb10YyuMjhY
oK9WPRraRu6J8ibd0nyXEs9mu0YzT/4TBq1BifNCsGH8FMRBfeOjjEky+e6uo47lQMD0tImml+R6
qAhy7xZwrfBSX+Wxrt15icF2UEJFi+LfZRpYInXq0oMAK4WejihqGYr238Cv6j+ISkQYbYzt9vxi
7KAy2CTgVgf63eWSH1aofOJ2DOz7/rOU2YukC1kH8SCZGjfrepbPljQUWcyp31Joo2d+fh+OxdE6
uhHsESmK9a6uVwaEIhX3j9tAVC4zcX97jHAXN3Lff3TPvYA4MRDcSuXqmt8Ix/RweVeKRpmOGUA6
3h3qCvp5TJqd3zDpS7nK3m9E9k3FgtzvGPyJoe9Zy21G9CUYntP4o6UJPcdnPslQglJVc1bXZ/t4
i0ppYLahXLliixEHIfkm8Na5RBZaViw8cHXYbBMc6IxS6w3Lm8EMrYfuFnexuV208uMLGV7pURJi
d7YwUcwQM00aY6OXw3I108vaPU46WcP0Y1ZIaR+eZVcAsGGonGQCG0XOwmeIJPdIbtUQQoqCErq4
3CwkJYVIgDcC0K4J4eb+OHGt6PEwEwM82UUJvPoC868Yj+Yf10J7J6MoacqnCJRFTjNcrA2AO4bO
uEiz2q8bPHJuVjFV47aHirWrys5he9sA+7N+HeuNb0qwkF3IJY6KqFa2vkilgz/NDqeHL/XghEeh
x5OwpZSBT5Je+sCRcoyd25T11dIznMYyUsCy+GSwR+qAs8v7ZQWa6q90IcaO4Q9wY7GQJVJUVXs8
d+mWZeMZTF3MRuAAu3ir8ucplLPpVyC8AzxYnxKO7iu8Z0b5y/IpZ4y5LvN0K0oWYV3RWQk/R6+M
8PD4hM727nCt8sZ2EWpEUxtNqRouaE+OK31wOO3KnfSfezMpuMr3bDjH/yh954Bnz6NK+sMJchgI
uifBkda+SNpCh+flS40/hl+GZU9lBScC6V6toEgQ9tnSw0JBA6N3HbYuM2wjWM4MAq3NnuGT0kDa
spKGIM07E0NY9+FRjoIVJzI68VId/B3j6nCDJo8vk5/Jp2ZuLnmeo7DlB09Ym6pJOvG81oPkkP/W
vX3hpTvMHwuYnxRQnlQHSkwXuk75Tpy0q+ydwwVykICtKL6CdBsrpizc4CYv7oSrFSn73ug/MgOh
XpD4Odm4ua3dTfCYKFsQKNRDY/EbOPp9FOYOiciuA1ohm8Izc5dw46RRBTlqdA+hekNHTdYjyPja
MUq6k8pFdij3MDqJ2QMho44stuDTgIfgeUWOuh0fvTKXBypHjvrOYEIkBXrzpHLyZqElW4IB8bOk
aFQIL6yY66q775AeWd7e1X//wgFDeYJ4jS9vEUbb12P4qR71Lh5yeURH6DvNJ8TLA6vgAyU77QCw
e2zRfiQyETjf6Nra0pGBdYwy6rQ6pQ7QnfIp2iyTD2y+9ZS1RVuccEAOH1lsoWwov3yNy9dwaPV3
cx8Uoqcl0RJntk0At5K2H6y/c+sMbrWC1FeOUOS1NUzV1XKYcSUfp7CSUHNWjpBdzrxyVJJv4ano
vMYHVLj607I6uB5DHMNee65bC0Q4dhyoe81oTAOXMgryh2YadIeDO5NKl0ruTNlQ4DJbW/5y2Csb
fmeNa8tm4nwca8RLu3dbgRurku+t8uVLxabz9NP03LnvD0R8v5wBm/Sx/j+CnvJavaJaXYx5nbNX
cWl9pHaNnCr4UDh6xbuGITg3o3/S66V2Dkwhz8Lb8XZHi8WKK8hTL9dgd+ruHzdyQ9YOREy8K1Rf
qCCwxBLzs9UwnbORNwIu+SeN0hOOiDLeUJz7FJ4x/RWV0u7kL5iHDgJEpWJ1ldxZyeLUzswzCFEw
5aTTgxdsKECvfN29AI76nBSVbEqO4JFyQg0KgwdyEHgB+bgz4UCVbyHyT5tggJWOhBhTZB0nqiWl
YK85z/lmrWurRb6qZYsQcrh0MDlRV68ertorI2iySmPnWze+UsHs7CE48dAViGAYsDVbOqoEkDwK
wEW107XtD379kblJX/tLsYWK2WB78yMApwJVpfU02C+CPJA4TV2HUCc/mntIhYfNkgaWveN2QCZ5
LboZrvMs5tLobPYoielnih+JE90Fh4GgvVUQlQaSWkuVAqR3WR8ZE8I2SB12EgozRlx+nPRKA8S/
t5kZtvLTClfVu/5O/aHzJTA1qIAVPQPDBVNo0cJyj88xWA/Bb/JvLyBns4L8U9iRxeWeFT1CjCyW
hVdg8cXKBezo8WeZHN0SvuVXdJ+tjpTiwBuam2ynjJ0SiAZlTdbp4nWDZSJpGwnfQcH3EBRd8Meb
Z1iGYHwWKfhwSfbhQQ3DFtBZlNzc1OE5PqlSfYLYTYSuCovpxBB/Xap6dqZgDONvgKNkv35Zjorf
l5UMJtLbDaHLRIDcxXUBk4qWqVYAtNjLKlJPCDTBV021sNI6VhrPnKCwa4BfnGKa1oJSVnfwF5s0
etvxbJrhEu875ZxigF6IucK8u2dUPmWipzKEUQYKiESwpr5OQeKOKM3SCreY6rSzx41F1NMdBWJ1
tyeLf113bZql2Hr5S3y+vg+Cl8B6Qxsfk232kDnnBsW2Nw+pem7c/x2bgl18/ftMmaG5jtuCMQks
J0k2f0yP5lTKXXykG6waSmjx+c6gOykWHKk0DHifd3CIr49/yDtrws+2j9uVb0sUC2Qv8Gh1i4A4
1pxWpEB6DX2CXZ33S/S0WPNL3h4V8AXdOJig/pPews/okydlzvYdSWorL/UcBo7x4tBiXxF8JAdA
olptj0fuqcq+fdxV7gvZaAP3zbSco7ojhD0SzRr1KJW4jhN2gkU6RPSPGFAX01DIVFRnHM+vDE2/
mCsaK1PT4rfEEAtOBwvaegkzpWkFaVmep9dRxLDGkHVcAheUvYrzDxFkAo9y2xGcDRGf3vvBWXKB
9hWacPhN55VKrrBpd2jxePflVY/5QqPV1HDSxb/aXlY6xFfu2zOwyrqAlknbi4fXnxToRq0DTXaH
uKivNw/po5Xj8gNqkIQTIVOGp+wP7qYUAj3uyG439wTBysdPgJkf+7SmX+QiutsSK80yVXW3ex3c
yCgGUYtirFtF3+g2xlg2AQVmhO6c1Waq2Fik/yqRm2rtKTqSJVyqXUs8RB5txvl4PX1cgEzwcen2
Dbp47Z/4pvph4DWpI30/cEk9PvtAYdz/3qlaXSBzVyt9pLJfqU4vNCgHhNb8xiU7YNm6x3I4M6hi
ydJHrlABbmc1L1mukzXU/cX4iX2nv49qrhTsuUSArp+gkaZiyg5XwbAz6IgoupAko3czzGAmv8NA
6RSJ1QiCkHyMn+azE7D8ORMDgvkUWSL/IpprW7lpP6JtsIb+y0LEfaoYjOs5QtIlKswr6w+yi/Dk
uVPZxX+/VIw6zs2/mF8R9oq2LI/WRtqOVWcjeCZedUXIpJ96Nk7CX4TsPvrERr0i/bN7EprA9+m0
AfX65D3M0ZibjwFQudnSbiY6ohJ2gWGJmw4G8A4wcFEuV8lBERmdzT5GuGSsBuZNknWGGEIt4Z+P
QB94G6+oQc/V5S+qHeTgxERjyLwI6Rj2CPsKkRD+sER3nHTzM/oALIP3gfSp3ZPRHVVvLicD42S2
ifqrK/NiVovLCn9VLYx5bTa5oHb3s37YlIe+LVZS3RROgQDYFeD8d1bVOX9Strhi5qVjHPPQHbvO
ZLyphw62e0Qz2pwItMGRfdq5p9X2hu3CKGBD7evGYOX64qs6vYOckO0iOlNLmqVus86iRJGf7pG0
CcnrQux406uuOdosozfqJpumkRwqS3yARDNqSONXsjXFVV6Vo2H8j8ru4tRNFTZgPoabB57+s8D0
aa5iUkyurMwV1f6XW1a86louXCkoE5xU5YjTSmNNVvvHTDLSiXGYKPq4rvDRFGNFdwoW20GYv7Br
eyjXNtpkG2ynFSFee/1CCf0wAZUgAiG97sbzj6t3xO1y+sOnSJHJHRMl++nw+1krQNvpu1JktmEs
IMceRG4/GlrsjrpWxeC32dSIwwbAQdixABXeGLs//shO2kySaRb3PUtk1jd+qNps1D6d8jv+fvKC
4EDIRDbxBlKM88Oc8h3CzDYy2kokJ8+DjfJXeV30q5Hgw6hzGEjvn7Squ4maBNbtyGMSkcFRxwpK
Es7DWWHlR4CoFH97xseUyZV5KFIblynEP/3Y71PuiBYVB7U41/unAXTrG3xcH0fMOQ2T7O3HkgeK
kYtLr2RhjFebdW/eEiyncQvBSTBM4hs5K9gfLgfW9bin8vMorofNmnSd70XdQuPHvmGkbjMdyGTE
9GdBu9hcMn9oJeHOW1jOF3oc3JgfulmSLZI6q7P/DRLk50rWaKSsgm+P4v33KQGcvaQI28uaiKK7
4eJdM/SYp0DKW1/fJ+N4wzsx1G2IPB1BeUCXNNSnnEhxTn8MTYqZ2a/jcBt5dx5V7afhHXETO1Vj
JQ3E3xom/OIifaWZlS16oc7bAnypjZw2dK8hsRLCHSbG/UfjushRopggyaekGMRJtvL6YQAz3Gwh
hkGbtqVLBBGkA2IAv4f8S1Evj6AwBRA0XRaJiH5LkdCf30+/UItIJaJf7hn/CIx9pgEAx48kriXe
OSdHWsZRqM5AoiHmqfpECYHpSApO/UEvRWgmFDBoAu9uSyOGHSh5oT3ewqis+xJJjmH5y3qNrSpr
R5oOOM/S/dhI/lV+BoeWvh3dS6dET4lxyxGOWoft/Tlyt9hCcNJV8KwoRHzJPXelyM6JKYkuu2Wg
nUGT7iDtO6h5a94MFkmMu+FG4P2fWIhrNL8G9HcTUZLeLx2RHhPhnw7PE6KI0ZpFnG9dhE5UwhYJ
NhUGtQb1B3m8tivMItiF6XjtTUH2xIK3iKOk/eavnmEVKQ6wfEs5HouehnE+099oj1iQN2g7fP2G
4w1JCG6SizYAaYSOdTbf3Te7QxMj5c66+o872ElXkxeRgp427mdJ+QGG3Z2XJCrIwS/x8oD5BJ6o
Yc2tkso4oEzsIvJw0vUhDnk3Ut/1cOBWwSn+8z+5UvGU3aGB5XxLO556KcCq9VVZtUZvtdjH//Lc
nqX0Rd8qRRJG40lN5YFGBTwl5DHzNEaPEcmfRqWGyGJ6ziDvlxQ4cVIlK5XJXp4/+5FdZWcaiFtr
qfkXnytKCTz71exYm8NH8rsPRB8XfXH8SOXs+O7TlvXynajrWunzSSr+0j8iEb0CnNS9uAEw0Aer
8bQtk3n2ru63uts2m8Tk7lNVeTBOfxMZJdNRh0ul2Z+/tj5eVGQTQwsQ8HQLs3dFpimz1l2ls1kw
sA16BKrGGEoyzRCaC2ywOJuW3N86hWkgm0VgBJEjPhrlfAbw7rXhXPeibC/rpglyhBqsZ+Qcyb/O
96109guWzYzyo2AfCPPFSxMkl8nP7cuVVRPL6t64itVFK1v8g/8L4+u2Z10Tz9XoFVv6fEFm3YPm
rKnTLgEFzqPBLO33/Aj2OGN/wepyz/Kd3VCoeuzeT43DTakGswi1rGOJU+OVnfqgES1P3CJAC1py
OOL2hIK2Oz5s8/d7vbsNKttQKYK8bbVuCPOR7TO/jWboMAHteccMTsceweeRvgBPNzT79nnVREUx
bsAtKZBBXNHI5AgmyWvdGt5n76gcmq2GODeCxAnqZpRLpvIV/9BfjRl38bbJw4h4+an/TU5hvwNl
qz740xWz6lSBvbu/H6DVDSoAAY1bJyyoq1JidJuYYRXhnS1iPXavg7TI0ATZyjUyTcD+t88w1wK2
clB0W9SyuzHEGn63leVhlhsNAlA2lePCLTyH/R8FZyWomX2PEJ/ioh8VFvIUrrbfzyQVYwVv+L1u
fbSWPOZ5hHooB/l4eDL5LqoyijGPnKRQsnpx0V6/zpT03WZly/HgUanxGclkwt/DOqgAM2fYfSOr
BbgWFgmTlSGgLZm3TcuRUtwdkK7jdINkPxFi7DR+W+X6Q31UMIBtofWgKZ+lRqmuBjOH4X9/KQnN
O6BAIGPhnHX9bMcDGaE4zaR/f0wg/8QWdmkvJpuyr5s6oQI+/CwwPKrew1P2o2egUpamb7rfGuv8
O+UlQG4znnEHYVw+xx3haq7jDkco2AK5t2NEt5btereyEVUEsqS/+R8iuveu3X/j0AWL8CpBWn9c
xhmWuMISa0FM++ef2whf/PY4eAl+FSJxTCq6w8oCnhb67eADtjer8geVc0wbn5v/XhrQEGMT2LZe
Mz+zSlEBrCTMtlvIIizg9eBWx+gkwxfcbbhUIxGPbsAMvTXSy0DOGKKN/TyCMD2LEramLI08/Fmc
xrdiBFitG9HyVg4265T1Qv47YV9YVH4j3J0A9vpYzpaNZji8eEGwetxycIET/2n2DJyAOPxbzC/5
focQihfFgE2BjUhatIiTdtxFLIr3ljRAO3w0t4k95G+zBL2Twa3ruy/j/15eQwNyDF6ZcmK/3qvv
RQa+/tWi9Ts+8yhOenGm1obK5leNE0/ocGpwK5HbfDg5QQXEt4EHBHUoL1qFTNysnsPHFKFED+XS
SK9LhDGVki19WuRBtsIaMmVVxbRuLHwscuR7Dvo3SG0FzUe+6Ewshv4Qe6mvqeLZB0tjVCk7Wroo
DqAMJcVL6ycioRIigD4Xb/WkDB0YV2W116pDNwfOfjwZ3hpv35QhwPSFVe8cy9VWbrCSpFdQzgwO
vd1QW5IHAftJ/0bDnUTZv/dOBo7I2W1iawiavOWsyeKvk8PqjdKLBDGyv5qbujSrIGr71YszN5tH
n3u2a1EJJn2iTWa8coFQn0M0ST1XX9i363Gh2cmojmi/2Bqs2eIhapsl+9bj/MJdQ58a6160Unpo
9LqpAbcicKJvkDy51fFVRegU2EAQh9a/V4T6xkwKpNwhfNH3q10YkVTj13RNfQBF/ztp/dogHIKB
toeQalOhpwMruNvLVqaxACvkbaJLLtvScOQ7mX54ssYHX/vLD684o9u/4+NUTrbo5d6/ODFu9z0y
shNZumAgGPNKwx/3gB6Qfi4jsQC8jp4xUZxCuNAFGS4c330AgrCAGkyEGtXnuPJTXpaZDa9R1PT1
36almOAo+plNHsJBjrl2afcP87UZ7DL2VVCLMlpuUlZ+pp2fb0rQpLBknWY+wsxekBqGoeoKwIub
seiq318T294vhUJcgoABQ2SBhitrc3PaqkPia1/vgFeb6ZYjIpFaHvJ05DZvsVYot0LiblaCWKIr
EAbI3ZsIaZTykBHrIOGJjJk3414RgGRkwrTge90Y9kvS6XFBsompvbT25U1sz3pHf+EvMZMGG6+E
O9WT94Zaa4CLZX7wvM3LhRVGdblOLnAfSxBJwOp11O9Pc3pi4yUTI2sdHoSk94QHZ2uPMIR9oWa/
MF9flZSVurv+Po88Fnnt/n/7pCF7sVZOMkPesyzsb2YvKk9ry9P7Z0yZJWTys9ZBhlpqtzso+gR0
ATBotHVuGPjRtuOATq3nwYBu4z5wtrAjkAlOxmSzF6RYYrEzOItHhWBqCPzNYEVVmzn+ayEsVPEJ
nRKterAHnt2jV9Rmk/PhuI03khmIZCkevv22flqnspQgt6TTEQ9h4tHql5XoCPzkvhJAp3f7cIpn
Zqi8IE45noPARIobEoe2NgIMPt3Jy3mcbGzeJc7crjIVWxD7/ZVWbZp2w81zsTh/JdFJPmIb+mAt
/WYuGsMtTv5SRTiKxm3KOe6Bo/LoR4R00rJbx7woD61xqKJQdfbXMzdAJDUhBxZKN7zRVnjr1/fN
8DuK3T3vsOGKotjfK8+lahkpieMo7A609Wk52hIoqaknI7pQexX9hr+eIBKt5993XHlr74pgl6lU
CILomkEhgwwwMgcNoCt+CsZKO73SIhriQW5BaFuShrtMmhaSS2QSclFWRnxRYBlSrIHlBcGcEcHC
Zrk0tZSynFSTzxLaxosk4IEIQJ0rdHmNr07mau4pv+GP5fjchAhTQwY+EXr8vxOSX09w6Wt9zgkE
3AWoTbGYJ6kL35qIUTdjpKA0DxIYFLMEsQ22+9wVsfY6MaVuY7ewlgarhK6FNF/J/g0qu6bWMuNo
ONjHSTIuQRBEQB5keoVsGCQCPWB4B0K4j26duIS+zKRNPfWtTl4606Kv0rpEn7RWYFeV6BTVbEzA
mQo0P3/2ED7I+GcWgrYvBdKqdJux6t3cC+Q8OL+QYsM23SpdmC/rmttYFAyiQow9CTDQOylsQyxj
RsHQi703w+BGPf6ym/oMaC8sybi3+NtrR44HUu61BgB4AVSDq9qrIKuXfA9DruqkFmM/VCSZ+Q05
HiQJe40auvRPQ86Xhn9hZYJC2ARXC2UDMiRVnXQR7DqnDkgSWwiRAeT+eJQfCAoRGR/xWGMf4GgX
1hHyIjjjrLtczzyYDspmWxdeOP/Io1yQ3IhSCqsryhcBPaA3Ae8JIAjcu6XcGZz/2e9p3ka2m/lz
BdsYyzyGL6KLw3i1Q4/qGsh6DE1DuQnZoEkVNmmdAtFGvw05aCPtEj7EmlvuZ/DFfZ4FCfjGfKjF
4Qko1edbgoBVVid98RMmWKY8maFSzWSZ2tqjCVAKsap57/ng3g5gcV6RjIj+dWDDWdWW3gFZ+oW2
KLN4DUYCfHljw4M+d63udhaAr/ZJpRjk/xCKyyLcmDhRn20c5YRHvP0yce7b5P0cnNf53crIG0w9
EGOVtwbChM6JHDAlXlXd2vW55BXriX0/7xkFJ7LGGG8wpW1GHfx03mfn4MsTy/3jsjJPFAEHS2VT
jjDIYTqLfc3/y+KJRLDegyN1eiA4tnANPKmzUPMa3yk8tNCJjL0NZ9oJyiT9zyokPbr/YvLS0/BT
o0y1kSWua4Nq3x3iXzfW7bV7ghSuai7ujBvIHc/otLZTesGvbfHwxon7TF+oYLPKLCCCyJJce3ry
divrC0GhLT8p6qZvxC4nOyemoApYZLE33VSh/NrRYItqmLXvwtbWbNGkxCCkfmxrvuc3hWnjDj+7
Jrr7n0mCT1P/EbcXeY1R5vkFumXujLCIhT0ceW41H9b5rzh8x63PBbGAi6E2/I9m0a/nFeOYXg+d
xzg3FN5bi9AmrPKVIRXLcV5M+pnCtjkdGYSJqEkrioe8MCLU1+6DZmuHbLvReRv8VqDpGzBt0oSL
zTUZ4+KTovz7T5h76+aN/i+Y3jtJF1vIphSxKBDP2vv6zU4tSqY5X7YbcyIWvNKmvri27l9AhWcx
wqzvQffAaAl5yET+FGChRUnY4iK5X/3VGV5p1t8kVjZmCuzrAWfCwj4VTpOCnls6DQHdOJ1f3uIM
6+G8UFlhPSjHtYc+DnWkVdRguq3N2ao+Uf0eq0Q5ewNn4yb50+tyHLqaKZDVxVFY3AEJxLboWzB9
xVyW8rIuC5rCj48XM16dZ95tKf9RsPSsfHXebRyp3ydBsHzdRgZ/s41AGoDN66Rsp1Kj/ff2GCV0
ri9xEOV3pjb5tpf3Gv6NsJn+gAP651EwyIU2lDBqDdEv9JL1S10qsj065ruTPaVRKDlVso3qP3AU
Sl+2AFmN5Babc+Uz/9JwSGvOkXGD3JD2Ehjrjll8Jq6jziUq2kayHHma0X/6Dw+cesrjDDXPbG75
hCODZNkBMdhD3HmlKNOp03BBANNFwvRnRour3I+SE6FZZw6BWQjxViXhtyLRHB5yd+Jn4CSDqPDU
DthOC5wrZ7tNg1m1NEIglYUI+SMD77pM9d6XDNbuCRlEVF+I6DsGfChPWN/1gIm3o9h+TgSKTX07
gEk5p4RyzLips6wxLOL1Q/4iRQhLqeCoFN4l5IThV2JuZZgIh5IuaNo1HBYsZU6d2jjPC0l4jwpY
IKLx+sm88VmX0z6QcjwA3kVcYdi3Hv25VNBHlYtl/1+F7UkZVATNkdNfv7Vl8/GMOZc9a7AQcYPY
BwTV9gc/NEila0TW5T5KVjBs6PSXRBHtI4wLFZQfGkS2bppOWKJpxazloHHNH52jUvEuDZu/mUBm
7VSvcVbLR6o/JhrjEjlysKBQHbuJpFvtr9ONXaD9CWWBcCMwJ21QvaTwwREaeUEJ22iMkKQnI9Zx
L+S0fzPd0tPHZMc0DQpaKu4r8DhVtdU6FFlGND8HYgkI6GOZI20NJYYBYmp6h8os0vP+Psmdm2hb
TylDDYV2zqCu4EnXcAadQN5ud9EKl/tMfQSdov7fWNQkzp7BcPzY/iVFsqZUcEhhkecnBMvbz4Fb
uDY1C2PdaQ6iUnPFdwup6oQbE4tq1qtHFcrY66J59vRBiyxSwN+M8ZyuXW52Zusay/9LREwmXgDt
WjlwraKKG/Edg0lxnpUSGejAILcNtzbjE59FmXIIJGYbGYit5hAo+nqvspnEXBxjIBQWlhAQo4xN
38j1E47OLJ7HBxNho8zK+45sT4dQ9jM7d+D6fXPE+3EGReJa4EW0FGEtv/E04wkiiSl1Y/kDqt5I
J8OqNbJ2h0uwAtDI4YqPtvxloOsOTyYFDb4LI+aMPxjsh1IZQQNVBoBFaz8XxgH1tqllAbKVp5UO
vTJZBiK9GpnvVuDf5K2S/xOQtS7RY/8DipxtNQ973W7wlOBmv2lbgWWxA/8E98ky88BXM9xq2P6B
/p/fwM2KLK6xtyrUeb+DPyKPmCFd4Hj2gCdNibZum2KKOUNX54o79oaPUI8RSt+LJOGDTe1sz+a+
iSyevTV2UF31SPxPY48az9BOKVmcMoPB5UfkCNvVeU47qWzU+koV2AcbBPl8RdfR1BnQqNvTYhia
9NFFTSutnYM2Akp2hmfsFtAcfqKTd9lhdLip8gN41ZVKZIQxWwll5DMVwfooMJghR5qMjZay1WVn
NPjbDC2rVJVH4i0jqfLlYCltCTycv3dq6eERo6qG2SlNkxWGpOrkeRseWPUZG6iOrXDp4Gz87Hc7
aKHUaSale0w9FQGBB1SqjG32F4ZVklA7OFybpyovkTpmwUfMav2Ry1QQuXDb0dmIpyV/qEfx8foN
576qd8U/1hbZXsSVnCSOTgdtMck3kF7P1trtNGLSkLa+wbWyYLB/lsQGdDy2sJZgu74KrZ+Y8jD5
Cf5XNSQ/HOHPYWV6UTQx+2LcS8nEw0OQGV0K3V6linTBSH5VPdHbuq+1TvKBu3lRnExz1pTPzqpU
OV2Djq98E1WFoQg/ETtGpmz0vymEASiz0AjwR+l7zahOsxZeUADnE3qSUPf6nmUACLy/sImJ2Rzv
3kc/T8vmi2cBQnpjtBrO9ow+fM9q5fLzcyYbfHTPwFZG74MvwXYWpCy9BUCo/AQmxsg8SLgkBR1j
PtRJf53URufaKfsQKRh8DCqSg+W61rZ0+Lxa6orzQW8yhcnlX1TEqTRWOnPCchGY6+2ii815s4Tx
F0v/REx8pzW0DffYttx2pBUby/Z5qNe7mpdTbFcQVxYsWJTgeRkZYdnO5ZdudQQQVNkIaJgdFVgI
DuC4shBt1hX7AxOmseRwVI4KJTC7BO6+f/UXJjtYNZ9fX9TkzXlqU2XsDBRoUb8gAd3V/SFveLrs
ULhpzBSakSIeBp9TjJLZKqX/dUfzHd96TDZWMKN02w5tCCCU8ug9iOjDNghKbNgiLrwFWvXMnEnK
l+HzheD/j+S6Q+PQceFMbIlrWNF1YyKjk3lQs5ZOtreAinpY8bPmhytoGzF6mn5PvvikBjEgBzNu
+F+nXg8qeTmNFVT31dcbEYcYrLQrVU3zTh74DNoHiX3M0XuS+i8ADjsP+gbkOdd5YhyxismNbkzB
O7BGMs4hjfcNF5bcPToXlUAQRgSdIY9odKHj1DbwUFXqVHT1mIN3c3DVlpdrWUM9shc2YDWuSPF6
D6VRpT+4EvcQRfxqRmWKsXXMC85sIF5zC1GBaFUiCG3/id46MxMRfP025m1XqTVR3Yjx2mtVvhge
zi7+iHm2JZAZDeW7ngRYXhMqvvKllPvZBWroX80QuN3+MHZZ5eIC+satILjyeFq5lgnrypg+TRh/
mRoXbwqEokcvqSZOhfN7aPsbjiBr2zEMkPiJ82WzXtbhKpiuR0VhgMhSQgH4nxd54/zJbSrD/pBg
iTAUNYCjB4qc0rJZPJ4hv2uhrYTfFkyntmytlT2V3OYvsGW9sxK2J94hcmi2T937RXJBFafsYii8
QiTc8V1/fNfYkDSw3o6dn2WYBBCXudhiuuchhMgcDi4ekA+gRn2rOzlZhQrv30itWRbo6HUNpFIr
EIvfIe7R98iI/SpH1H00xTKQLBk1g4ua+0/OZm7/GFUAi8/rnaluUJRHzf5hs2255pDiRonucBkH
HAzBfib0M0w0XEo6u9N4IQDIcV60GiYYRkBMBU8WVlsy9qW4qwgL6I5KtFyF1db2xkSUbxU/+MF1
QM+gqGl5MTwhp1wTq9OlG8tM3DhqvRhmh3sCkMcbx4aKY5sJGtLCRz49uVfVdedGMR9HXgLXP3UO
YOe1P5x4oysFFbw+is2SEZkapijnvQ+6b7OnQnTisatBJRKbsLLmtMajzOmA2TGcxqbtKwMtzQir
ge1E+ubBQEbjtCYA/QhFtp4HIK2NAW+8ECXhIrdXtSN7T6wUhj7IND/nrr33qyCLwqG/5hlMswro
tjrBIBI95M1uRNCpoH3GMF885oFmXvz7gkRVIdySrIBiYErxHfZg6fSM0hTDGhv0ehERB6P/M3Cu
D0TppwGXtQuQ9M3qa1iLSrGtRzlahQMKWTG0+USpm6tt7GtZ3EpJN6Webha9VzppyWDNhOjGo2NY
LtKUInsoNVZGlAKfW1L+PpYWoDVAonZjwviSOUdlRC4xCnXYmykVwhY/RXZACfMAnMxn+O5UJ5k7
uWSEKsItbDTLwDpKBFDAPFqeib0Shp7HxDmpCTXGnVj10yRSxbsr8XeWrCWnrlz1zRwSo+wvMfl0
zlVDFAgwTLD9O6Rll0kmPDQ//y/DnLegJOJwVp6VKtr+aVRooAnIBFa6MJsMDRmqqA2zsotiLyo0
u7R1NVrztQP+i9Nb/3r/YDUP4f126JdILl5HdwcoZx8OFetEs/sQba5N65wbqo1ECawWYgmpXjBZ
bama1acOcnogxAFVLIY81DSBt7/Z6ZfkM8Wm1mz8wL14DbKwlDkwtj4JoF85Ekdvw4AJXvpq999L
NoqH/HLHOOlkol3RExOb9rBF30pIj7tvw8REJMPJuGD0Ol4RwZuS/RmAVPc2ylYxoz+MOCeBC2da
bo9CCcJnb3uQFcj7IkQn4JaRczD65FB9jDGeg5UMPflRb3TVZK1EVUU/ZMGTZ8HCiNFKSisxphDV
1wC9UIupqm9tvRTIM6QkyFqmmhHoC3sO2A55m9toNG3dz7Sbn3NXd3XRbVn+7dvHGf/XpThptSu+
ylWFhJJMJHeClZovuu/2WsvBhOHgKeaj250Yml922ShpAXpdChUpArOgjlZh69uMDyIHU2jkiwvX
cWVMsKREx1aMPPlEKNYofExBvxyAuOBalR5SMT6+etVuIWwv6kAKiT5dSMp0gUgLsr3dtRB9mCrl
KrHs0uMJ8/YyGrIv9Gx6dktyRrtvef8rRoSasXXkLj8tYM2RbLDl8BX2RCUyRINfDMQvQHLMnwGQ
q0SYDWR9sgt2KkyW+sN1TteBymdn5K7D1zGh/S4kFedQ/1yvKyw8tchZAp/1Ngo8QC0A1MPzmk0B
ZC9exCFEEUNv9e347Eoiz0YhzMpzwsoYCiT6d9wfdA7MLdUnoioA5s/BvwV9sRRvQnmHwpj1kNVL
E3B/V5m+LR7bEiAXaSw1uV+SSzylw+gkfRG0CKycFK3Xm1dyXvLtyGM7C+0uWzpM6M65wC0c72Ct
v29UH/+fEuNuz7kdL9NUl5fEf1sE2nbVLU5ORAjWk+HnsUj9CaL99sogZHSxE0xI1y+eo8BudlYR
ZAKibekaRIrRPD6WleSJSZQthkTUFNLN0p042iec5uPTLbk7gxpJWQvfzWkzhfUtuOE6NxG8sFaT
ITfVoZpasoF8iWs5kq0nWdDUT3r05nk7WdqqmoWK9WQkWOjO/Wixmq6rjtJQ2kBGxsNUQBRsnK3L
cscM9u9hJbSQdOzzYolGGlsSv8BJ/9KJxc+5UAGHxjDDAAUzaCrG8cI4zWcOMj/MsZcRK7+osn3Y
jStetZfoYDV1VsohQm7kLmEntbGJkwk8HaRqVtKFzvWGwd+ptIhVvpSJugpcjemxLHMg/kei0ryc
fMksTxlgiZi7loywxmTop46S5K6HZNOONPeE8enzEdqBFGJNaUZ26HE/E/d6tHpHLP4ymxuxWh5h
jOyhfBNhD9Mb8sdpxvNtP8SStkKrceDL99rc3SITLecgDSvoaB6ZvAFSzYul6e+VuUEwTFS4xtZ1
snHOa/JvKgjGKDdfd6Zj2xKJ/l4qr29wCVV8wV/rkJZ0HFOMR2F5HUglTGRU6oUSO8OVwiRLUOR0
q9YtgcYS4G5H94VnDCGPB+LKJo3ohm7rFStmkgmOZT6ou493wl2H78iB1YWJvxmL7rAMFUJpFN8u
03HkM4JgoW/qpUHtM9K3gpBpJqrqkROdMmlFESxz5+ojw/M7Bbsz8Y7hNN8NjZzux4jCAAGNXoeD
btJxqofTIz++N6KeXykORJ0HqjTWL1LwqoL6abzHRF15FV5dCnUbRB65r9OwQ+M1fRn9DTi2QXlV
kYtzg4zc/73SbwIsotiIzPQ3L/S55qDsH99SyZDI6TpS4OWHi6b4w0RDYesHXcZmsW07Wj8UAMBH
NoohOhEdYmAKPzPeUDAFDmhCR2GaYuPs16HGbR32fTus9PokRY2bwe+giCTAPFcEW0ewBqaY7xeN
ofo3soF+NS2ca5Mnoi8HrZXUAWLj8tNq6v8aHStZTjeRI297gWqcJz5orQ/GdK7FHJNIf3NtdkAU
jA/9dBaYDcPnlpiSC28vOQptW9LUFmX9YXuXb96lJY7qEdqhi17gMeDjEBuVzbjUEE0rIu3sVKui
uXCWSL5iCJTrSxlzwPnTZQJA/g75mTjk/GpoliQUfFTWapa43KczBQ0mqd2NvwRJk/rsYIuJ569x
Ha/pQDyfKbm8GT4YwxOhR/VPLXsTF1sFGjFyAFdexvWzICFv0UXgO/cd/vqdXTS4g2kagI02p09f
P5ahMS3orDFLQKmMm4AArxV4LYLdnr4tmcLiIz4Ez9+IPcdIppWx8xwV47nxwzH6A2GgqUtYlUqp
HhVR+xVSpvK3iczwP+dS6YfFOwmP1UXbK0O2TfEp/C30hwssb62754i+uwdWKCDswmKcrB01fPB3
T60bPx3fiHGMmtErYs0JvH2Uxp2vQ6t2WYt+7Qo8vQaw3PX4MWeP4G5XImpn4y8LSDiBDgiLQTS3
LPd3LU+e25GBcUTuuhhMdwLgo2zDUsiEYyF80W4JJN8tq7cw941u9XOGKBQeyZv2at1xkso4F8Sv
iYWYoxTGSxj5CcXPB9ayTjPo4OjnAMIEgF8mPmnp8nC4zqoUEk1CLpTrsWTzSENukhI0sK/p5aFC
xLsdV7+58U+vSQ0K3yrGUsr/u2XGJFLlYQuBqS0zoE7IKoD+M51iySnT1VdHnIq1FX5qpSJQEYyl
jTi6Gic029F2kIA79yIAvCY/zuwii3VMuj4QZuj73vTZXQLjxeMEmnNj8shq/umiMXBwHnQK9wMk
FuQ2YY7VvW9mr3uaS2LtYRKxe4Vlg1R0QCRTGoBUuhvwV7XCwV4OugOW37/PHL0JNWJ968jQq/hq
D802iFE4Eh0aeU6ijquKPGO7XdSXXYD2D41VNxQkC+vVU7m7rWwOTu5VSBaYgnTorPKDQJD3JEk8
1qS//yDcMnG5LxONFIUD2XCI9rtA58I8SEHIUegJV80y6e6Mja5c735EGDvFJBgNU/9SEyTAHLNz
zvjgmv024IrNcP1IGwoeObCB7v8aVGc9P9hJeJKxQR8AjTxqJ+bLDBzSKK5DEzrMk6BMm1nZrt+z
M6WI0uvfWDuAPzaRn85sZnqIDrMftNBkOvLc7trvlR1TxPQm5rayDdfL/+qEUl6KhFM1MN5asqVi
AnQtFpHjycLYJVasSgNuxDbb5Umg/11g6CSJKXhybaxhcApJ0z1L8hxa4LZGvsJ1hn11fUTByAim
Nf21CAQKnzFGIPXNOSwOVD2vphrszKNJw71UeyfvEQGFSYMX5yiRV7So3B92aCAeor8YOj0QtJzh
phj0qxAcLTKrP95Fp/8swXriaGbLW+LdtvJmfyVLD8ryRuXQev+heKtFcqtR49KnUOdgAba33l1d
9G93/oYKVEf6TjXIpOkKpO5RzWbHxVnFs8yQRFaUHfapHZC4K5cnoI25U+fZ0Tn0c3arNYnfCxjn
PVi6v8xpiWPpazkuGvnt/lmKNMCZ3EHFNPuIT3Wv1IQc8V3XXqzfLaS4kQp9eTvmw2WZLSJCx2hz
SKs78uYDWGbSbuCgY6JQI/LKPzY1vXjshd1WKvxySIWwVsnnF9XpvfZROa4Is2/XQfR4spivRR1G
LIi5K3RzuUz5eskCQNrvckQpTUipm0QnaXlv57Bil3iARXVaTOIvem65aLCL8ziHaipUOgJs79di
basg8/YDaHd3WhxlzMivTV7h2E6rkegloHq056QGgiv67MyUdJ+9Bz9cYbXPGkZcrJQlj9fXfPHP
Ejz2ROGXLYqbt9m35q7fbDrGeLzgylVbtUPw1Oc2yVYojp1pgwpTwPGqRazxhnB5HQZwqppzpkzP
ceaZTq4OmMPIiG6BDXMVlMSp5QipS+ixrSwESRioPtqB0Ssilmx5tmb7I2hbTsi5YagC154rgr80
7KiwLT6Y3Due/1dP5K5sU+UeLfv8Fx3guIlelB/7ubxOxKW0Jrx6Mi4ZG0KPiBMN8wNVvweai58e
3GwYOjC+3JzDqrT4b/y/TrFV5W0nsWkYkXMcHF/ePpsXRw/oY0kpFucG5Rw9j2TgdsQOB/KihIgx
TYAIcZBr+PWBTvyMl2Q9NAW6Kmz3SuWy319NYjE+TbQEwcMPR2OtKacMoomnXfolpB+T1tpI/go+
6iKOtgHRBGvA4cI1X4WX2d4iU2OUBRCypZ83f45FVZpm5iBc30rPIINKFEHGDidTL8asyGC3TFnz
CI50bOHirC3gZXNMrOpiTk1sL1wFwer435T09M2qbimJwKodF5NrFT+wwD7R/r5FtY+Bd9MHOvHg
dWUDr3vBmbHBT+uDoMaS0rtEa5sOKml5ZFNMY/9ts0R+VEhzvHhZdszvOXj3uWoQ8Ffw9Bwb+qMq
sd7WfNs1g9E9bGznXHfgWS388XorjA7aWYwFXn7JLYvF62bFXh/icH+UmU0qN79zWwLpxdlrPHBC
MPPBnScNf6PyoJY+/Hei5iFBMXOeBfsJL9yuMyNQ8kPtC4aOoxvAEIpC/8I+ehhzzrIckTXqejS1
4x5S6WVBs/8zNWDVydhHWNfxguCNUQJAlg06h6mN8A936QHgIJAmucJBIwBJX4dXrmwFXKegbgDn
2329Cxs9YgK7pwEyvEfvf8E/buyVInmkGj66L/hflprAPiBS/t3K5qtXUOZQY0YK+qy4s06QH2Y0
AU9NXTbjKwS8rJ0SHixiiXQtvygJerSj464ktscELgoxkCAKQNPJn3QeFxfod2xEPZbGKvvbUrSX
FFRd0PgK0R79XX6EeIIBDM7mJpr0PEsaIvF1fVtjUDtbQspa/IhXsE1pa9WRSlj+f/7jHZ4Vc1SN
0awkyWxpLgDKayZFBhQy0TZX3UwNkxZ5Jz2zSD0nzzK3/GIq342nydpQPZbbmvGppuG/Zr93T1rk
kaHaXbavuP1PS47enj97wRkaamZnJeMIMeS/F7omLFVEqh+bYw0BrAFi17BTjN8+KVbVu2/h/whi
xWuca6ScKkKW7J413C0GwipnlkEExAMkODmijD3wD11iOvn1MfvHbN9O5A7PKKOTaboADcTyy9Ga
hO3SgFyrZ5oIvmgXmNlVxFqywylwHNTCjwighjJ1LPWXZ/ly6HARafIIGvWWvll1T9Eodbe11IO1
pH4PMsiKko7kjHXY5yoAeWdONN1Eol561Mt4wiU1yCzKtMBvt6qUUAI97ddR4tZHCut0LQLB8Pee
DRV0WDP8Jn4Junwku8Pv6oGZOAsi+pfD/h7Bw9ciDFsiFQtxyxn5wJlHSdgxbPmBV+LIgDqaZ4pE
DiAhjHcyoRi+Y77Ogsh76MZHwuWIg/n5t9ZTcdvoGm06OQ4OhnAGVqivCwrOEMAVjnCJUMyFZqwC
D4efsu+9u41acTOSgJUMSMrPnasGey5z+xa5LFJxqO56kbdJk3pUPBQqZ7hLb1qPZKfV3JRblgcj
oxH8HDUYc135RYYGmCumnHYk+QVl2SNQoekwdxYVAvYjSMPPlryixf63RrXAR03U7tDma5UgBtmc
nm7UbsGMP7zPLg3+qiro1ITO0AtS6lks/FBiTC//UsiUebYrznkAAMe2UNMJLauIfxeMuUN/1t1j
bPjPYKq1PJobXJel/CsvH3AShelOP3c1J7PEbWVZIsqRfZE++lyFctxoefWXZsXBSunf9qLm2Lgq
dstGqftftLl2mQB9frQlwj2gXyGSVVaiRU2+5JxwzPe6bcC1UAKilmzzTzBKAfYVxHba9V+1ZP2x
hGL85T7yrGvq0hNmpjggH8dRPi7NGT85MRY5IxrzB3Bj8xGvc9J73JeUhDPD9CuF8jttB0q65ooq
IyOXloxlbWoOpsrkYMuf3RRY9vnBlrGJZTFzbfqKm4tMG97liby9D1h83t7tJy5ff4Dz+Vfnz8gy
9+r380BEW9ybfwJ6r6UUbjZ2qfDpQKamKeVRTNsGJH0mcf+B4hxIHlSvEFLzImlb+Vtr39fUFMS5
btf2IiztZtyJzt4ukEdp30AFsAszjjmEUMT6mOcWysW9Qt3cyELyKa7s6ipnn3F0GrrzzjsHSnXj
TgAGhWFs1++zdjqn1yAHDPmsGtiAlMkn/BFoioultHPEmdyeS8flPUchYKXpDQj4fHdIVhJ2gY0q
Cqtypbcltk+sYeiFskPsgZ2ZySIl4j45Tdc5epjcPON22BAhKPkxh8uHRMtAQiBmJWSvOgywLrn4
LwjCklk/xVzSA73M+QMBewwCtlgjPmtTA2sLyRIYAHNQbyYetKtO0+27LIyi+HDnZcWG9T5QQqY4
JpSgXXU+R9Tr5JR+6qLw7+u5BxdTM7Vz2iuH1XMemVqLR+ICVjd1mHMEX4W3tYuzALaLQAyQ1ez0
FshUOytHbesMj3W4ytoa1tk2b1LB2sEHvwN0QuzXNu0lZAWr5/k4jiP4xjQNZgA4s5FyVUG48QY1
zdyn0QQmx809udb3u+NYUPIWmjGQU/YO11xabrA4z2E/u9pGG9y0xlXevJzrwdOQTcZcKLhxzerh
w2wWqCT2XRSxV+gMD6hNbxdSZDSi5gdAuipHmgnjQl3JW+n37rCrCFD9ZORXcu7NNm2BoshiLr2v
7EOusXHmcSOHCfwBYqSUI4dFArDSu3mgOEoN0EMVIDxTfR7h/bNtL/YQFjQ71UsinlNEUAP1Aace
qBWJqoS4Ksd35HSZKm16aO6M3ftIJkoKFbw/6obI8tC4qQWGgvoJuXFaV4tvgoVpL8q+1tc9kNtQ
LPJmSwN0Zwuv/Gx+H6LqQSpBJ3RheqdsjciIfX+WmZNr242TNFMrRjpYkC1yxWiOFb6leQfAayO+
HKgc8pVp2uM1R0QfX1agUPQ5Sz4TDAKmR2YDJEKVgjwpjNQQjGcFAOYb0BYAUPzhobugz4xm9oSU
jxuTDh4HeK4o3UFQ3aoQmLi3CFqSM5wtlwfCw9OYp2ERGSf0xIHbPBos1h5nlNMZ/5CDkx0A1rXQ
ieIRTQbXmukinmFhu8iFC3LRklR5JbjbyhkgLgdk9g5YG7mUYjnnMoO9RdLYFHnPW6o87G+r+uyQ
vPb2Q0ETlKTxGKK2kMcp6pTSmYF3BdHh+AWocPRcQ00GpS7E+XrGQJdTWzIz09irIPVhPlZBcf6/
+GGmn7Dq3jd+Z4O+81JGS4p0hmYisBqH9uyJF3g+0kh41go4xBJQ4nvyUaRszn7lWLjIAdlgqJpo
v3a1itZmu8CFHkjwZU4YsGhLOj5+a4ngauMomPw4P7MnCZhsjtcTM06ArbWgUdZM2S50WwGFanXK
kBK1I5c4TeKAPtb2K6PdHO4jTuiudwN6X0a9oZqa/fwZ3PmXxlTBiCAtjb6lk5FGSnghBC2PNI5m
PsRjTxR1njmcMN3dRkWgoYrdAgFwUEc3PO/g/xwQ6YHnEcUH9bW/Tbkhy5LnNSgIbUGUgl4OPBzo
SbNTPXwPvSvLnAWjL6NyyMaa7iKdS8NrLXGgJot/uQ0yLk6L8GXGVbobUR58wn1fSVT0myeCGsXL
FG/u16VmIUMAcGxjaOKjh7Iruw57/nk4OODdHLa2uZBe0msIGnm+dqjMk4cq+/dPgAtv5Fy2R/uG
wQt96Jwj/cLZPMNZoWgOkSmFk5KGZR4hro7KglS0obWu1kyhTl9AKxvSLKfnfRvgqdbXsyGcoW7o
Gty2/yXo5XR1SoAI3G0tYbvfAnemsqyaApLqORIe3Pxgvk+WsdQJOdU7WY8HXNQRvCo/u05S1dl+
HUsFg0baL/MXh2q4CBcfTJsLLOijfJLANypSCz0cvN1z6vcjvd5UjQPJ6ToDHwMuu5mBDHBduJOa
9rIc0NHF0iQZlyE515c1A9/77Ajx7JSwNbA960jc1O7e7WqslLYdFFE2tu/uPWTHbu9cVYHXN1ym
MsbegoTM83GmzBxMMIGymQ8MnR3cEDdhj3fJpKEeSYUWAgi877hO4G3AGyEWCsbbZRKA0maQnP4b
hR0yqfNR+NU+kNlSIR0Fl5lFIox0BRVAYfRMsE6eNXIjyDvy4fh/teHgbvYsnrIV+34CSlwWfFUA
Vya/zUbcvx3lWYWyNrfSONAkUoSZ+yMB425xN4WAht+bV+HcF9pJMKetJk5LlZEiA0gnqmEsDqz6
uRuSHFke4Bzo8CXFzZH3loJVEzwcjD0QStr+FfyIrLK/XOU/pyFuu/eNIOfgB3Vxg+T6UQluTaXs
pOf3hE/Lv7Q4igV4ljGBzZPaSFxlk7A1J8XTyf6rFhxug2zTrZkXJeJOBxcH5K7gdCvhDduCQHRn
nWkhinuCJ4GcePQWogXXxiC/nxqvZmG9XN2KG29XXobjnwEk/zFqm4KFP/LJowIHLsqWs7oG+RvZ
UPtLz4BS+oCXAzejSiZuvzOh8NaODsgZiGy+ROfpsg5FCrrX3TZ9Hn4EjGf11xU/Pz0WecjN5SUL
q7agiNuSGJcUWyXIvBgOLR1QFnU0NlzAqMsyKew7BXvPD2MfDGGMnfENnP3xzR3CtZieYzJMZ0aH
5O/RPCpeME4jtq/Bsr309gtXisIfTUoLsSQSHcJo/NP9fPuepjnwxQ49pNRX0hWg5n4IlZDuifZC
qHR3HYAvuFATTjxgbj0aJYsxbDpZF/wUDpTsGBW5rAmDCW/99VBW4qK7KVwEcd0smn411QtYnwIf
tdK6v7TakKJZDgHao2eLCPfIdwVxidNFt272qCB+t8zJNtM+SWfyl/L0HYFEGVFncYE4rf94xxZO
gLWYu06PwsKpLQ4o868vVGqQsD7S47nEojMf40bmQOquDIgHtoDkUfx3eDZ5NOFGi+1O1GaHz/QX
QGYDo6YHWys+lP4aynv1pCzpqoKdPMvwZXkQIWDy5ZIU08t3Ms4n052MvK6cOo0mp0yubHNgV20U
PKNxwYERZfBhv2fopu3puivZbOYBn19L06B49dwy86j/bj8bCEujKqkuOWNXHsVKNj7HbrnqoydL
PDVC9ybGrwwokQ3Al4blbZVHhZ/B2NU/Mv57K/I2myUIqY7MzWrqraLP2O0NaYSg1FKtPXPVq1e2
ec+y30HRDTJnEQ9bMwBBFjnQv2Wc/Ts0hm7lOS+/pdpT+uhGgi4/nPhg2d69gdXjj9nmZMxR+mSh
lKnEk6/E28V0id+/JOZzWDVK/FMFVc7DtGyRESUI8wM5O7SL0QOTtNZwfpbJwpglaB2OLMzm42N7
mKJJAa9X/i9D9/+VEagOyJBJBjq2AxXSuNwzto0KSkEFp+e/APUcgfXwOBgL9Du63ssP1OEbfRsU
Ze7e5lQFhBxxozpV1RXLCeamVYBgfzGxELrqbjav6RJZj36IfjfIkJDUKckfsDQaDFBqCPYPmHL/
EoxSnIEN1SZs7CAb5iFHAjD6EbNo1k5xhNF0WNlnYSALUux/i1mOZLD7J7spIBwPt6X5vwpCa0xn
HMn1/cSO2i02S1BJqvNzmgtwf8zGMOfuA6YysDI41Yx+ZR9g3+uGXHjVdu+UPdpUsf7qvd1zmsXN
nfvUgF5973cwjByjluJV1940kkWfngEwfR+TVZgYFk+sBlCJqRyP2SE14ce+GxMPwLbnHBybECC6
vJ0QxyaIGxZ9D/zASdhH/RaMQr3PO4qt43kmmMulspsAnvY/5dV30aja/6QcBxmcopes4A4YaYl/
qPlC4T1rqNYf8lt5N96ltSdf8TkjAnhYsZhvVWBXrjlQc9edRhfoJ2uaaydc4Yeyo34pw6MBJcaE
0ggUv0rm9gZshPUBCg+vNGlRTdlHMCFCkaDo9aB74QT7z24GIezWAG7fk0yhtdhHLzGe6s5EA6Hj
elmEjXg2aAwtJua16j7wdAaVksZhttNSFBKkHZBcb2M+pzPQdB0LTXrMiDNUJwU/Q9j6hQssxXIE
wBQuzJQ5uXGByjYN6LWo8ealehJFMDdJdvfQiBg9N01+Y3jYbIZeoGUVvuYxocQs0rbvMVpEYk+B
tug9VU0fvP54U5vQ0cKfbZsLEKsYtyNxvG0c0elospUfJYSpJBzPdYxmI6nIxz7gSFSbpUUsFWZe
emMvi/3d3bmA/UJDoWQQWU3L4nil6cE4pPTr+hgbYcSffRl2A5VHoBj0+kxjB7eK4sXr7DIEG0kD
A4HrFOMAZ5kNGktc+RxQlcaEqI/YXY5+ljxgg3BbD1VpAFhN2p+Vk7fwoxNgBxxdNFgOhnepDfHJ
nakOdx7/O0W64bt/Ok0peUOPYYp9YM1Klu/dSmOOpT9l4eQ7PQsq4eEHTu+35ljr4xIzkvBaYYm+
ZYAVPg4IfGUTnE1ZTIqzp6H5KHzY9TPZegkB/7nOlxbZvN0wwmX51SD4dGTiJq8JTYSnnyGNs0mR
nFtWY+/frlaw6xqfDuVTWLdxOwwN0Gd00Z0jkgs8hiRSmrKid7PPIzQFm1Hk9sjCWhmMo5B0Hg+w
5sGcKAZ4YPSUwLReOIWptK5ATQXmZHOcUQXZE/oDajUZxPko6bJS6vYV46VvrD9pVKdvUBZLSjO2
zHRNdnpviI2bK4NY1f/RMNdfU3CW8e0gmVYjLiTr7lMScicyQnwlMmf2MjkQVCyN58SZrUFrcpgx
dK8D0qygB90Qy49pUBIQ2XQwBs0nGi6xkjHyNWntxQ/eFY+qmQT1w1RMvZSMVXbTcFbko5FVWrUS
Epi+MYNM2dCRL2uIp+LxinTrNweQ6+10PvkFz9HsdYOcGwYOJwFu8XM6ykYHrCa2y6Pi7xZ0kICG
gHIDdCWa7MsF2CzARRtrQ+X+VJCkp22K/GxNK9j9xcF6inV7mMeUCW+Bq7zLC0O+GXHoM6JLZH95
NeUOZQoWzUZa34A3IsnmKF/C37qxVIgPHrQf7948MYng9hjKZdWLLRcIo5TZ49BlOWoMFLeObPH8
PYRgwL80S1ZdeOxS4fJXehU2wF7ytsjY44oD4PHcqXv3+JvOlFclxjYcZyAWKeGg8IPMrIfn8pRZ
wK2TGH94bLpEGMfPSyhc3Dp4O99c0aRgWhnRhNfV6c7UAmRDLnR1g6Xwkf8HdL11VzO9Sfmzn23w
FGgkczow62FDT0UZ8tIphZc030LIZzPLie67PP7BY6N4JU7Y79vexxXrnA+d1G8A1C14LdGzXfDv
xWiLKitzt/rs+yv08iqq6jK7BmqYMxEbOKCfSwhx2gbMOdXbWFDD33Txeh5mQ/8K1EB7ULjE4rxs
9H+KzovMEvGbDrxY0fX/qsMawU7gyv7nn5hFEHuctNGImkOWeo1OwGY/GNaiWMRkj+R3iLbpabkJ
y3dmHo5BuWy/9BO069n6EHKYTuDw9wC38oEqf+mhjeljyU7JUrddL+kOWgBokVLpJ84Cpei8wl/0
jEeJYFBiJzW4tinY5J1IdE4U4bqMuwwiifeOy55S32KaiLnrlHW8ZRZT7H794Dp5n/wnZPPOioei
seBN6qpKXW+0lUrdsckJCjA1LlryQZ0Q9KF37YzWFTbMUWEzSnlIlYJFqk15JblhAP3tbTZuvN6x
ZRO0w+EhJJuAtgm2/0oTFL61XPf8Q5IaBhwuUlkpp2RpSpy8c4xMtREPbwOB/slpjgshGde0yGPB
duZqMO4ixz3+vHQ8iQLi00V9hYIyWwBcM0biUjtWzpb07G2rzEtsi1KU54qQpaHmzBA4M3pX9id/
sJVElU8Dha/X7caDPFvdcyq6NJjHu4Q8Y8m/xnTw8o0L7mGbU77ydB3gAXhlLM9Ihf+cCd1mllZS
3D1nTBMt7BG5DixRb7El3rr84kAXVdAP+DjBw01VTCTmYW6QJKanl34HCsT8dBznAv8/ogshX590
ZGYcnPzFpUix07Iglws24X33DGZslY8+i+DaQVZPcxgQ5X9J9uK7zl12bfBUXNdGLxHeiMlDCumE
fEO/p5qBjsNsy8YVhhuxNKssSw5fROE+SVlaNm8wUGvf4gIDFaOjR4pI2KwJ9kMRVOTzXOcYEkWG
/5NPTLixRuh97h4YkT9imp+Vdn2bDFWEHbU2/ljW4uWYY8pU1iJPCKo3swb2kkerbap54QOEvklT
PuMWmxjG5uwdr1GwWDlUMlHSOfflL4hJotAJ340kiowpLV8fGGyZJMsVBVX+sQagFVdPqKsdbXx2
1khPtg9T+XWHolRMlMVFTDpp1PVayQAtw9VxXyTBEHr5bq1Tf2H0ifAgXlgtQgXhnOe8Ml21TIca
/zwxxYSoyzazm/bOSoAbHjCbnL+kBcPKlzATfEGvAF+sjG4AGVRhjeFe45MxuWz7F9r+8rl4jXyK
kCYzexH8dP0rgigAKHwvjAj0QKFF3nVqoXNf5u0s8dxz38JxXVpTNdzWq/ytIeI6DKN24P8CWbMe
FSW/IqF0auUqL+QUQUtFgEvPc+QQWKFTi3A/HFJa4hrrhVOHBUEWzYwtw2uD/c04mPppuA1UBovO
kaebUKMRTtmhZoAd9MnLsK96WDfV2WeJZTV04EhlZnMm6dpvMN3BReYSuSRoXvt6AKjNLMO5jBkJ
kWmSz8y5k06w2Vx1bqcCOwaJCph8EhglxfMnAse9APhcuROc+NhSMizCZE8E7xnuvKh01q5MMw4N
JjP69wtWkcNgihv9BEzdOsSjq1jWRr7BcqVwbdDAcnTSMzTx8uvWEI1EWAq3puR7yM6rGP4oyfwD
w+ecbJZTIKeQSRWMD2PLqw4bH50LDd3v/601nShY69ZQU118EX7e5EyADeETZaSw0ODOK2fn3RBm
DsLE94qCIWt2ZeH/Gn7Fe2c4+dBrD6WgI4usbtwTQMVjerkbgQsbROxrTGcjJqzMMh2s2PaV0tkW
F5yoJakc8Y/NxFCV5B6w+xWHK6stX1LFEZhNQRv9fclmGrVc0Sdb8XvS0ilnEfqygvHH/zavY4lg
w0DzVly4eucWXotpJ7ihrNcNxUO7Qczd57Qq1jLkPMhqLI3nhvymeUM7PGO2k4LNeuz2np78IHwz
O2UiK7f+mj2TgvB2VAPNaQCEKp5+1RjvWsZUx2ncicxgmLzEZbRTILA03gq4eH8xEP32csokT9zp
ewumS7ipE7TDYawSNrH6UCRejJpVYICouZt1y1gRXmcCMSInG00VwQB/1Jivbiobko0P7IeJI8lQ
rr3yuTZBSv4QSPgwOCy6LTi42p1/qRgTWKNrXAvgvnyPSVdlh/qCk/Fs4EJMciEWrtgDGMARu2Pc
JBDHYCDG01GAfZmsKHRp04KxyyFFw4gC/4BJNQvxEQG7xmpMLwE13Yd6r8aU/9/5zdVKWJagmyB7
Qe1XV5b+w154vNhj9itXRl/84pc6+V+lXxcVCqK0srCymgbQtdmT8VlYFRQzE3CoKk1FnoNm6szq
cJCaRh7BU/tC4qb/FTUofCKhh7iqR2HC501ChSzwF5VtShjn87KvjsGsec2w2wPXLCsAJC4MdJAe
EXIMyIsaDeSMvL82afkexEMh6182PYxChZxSRG57Ox3axgJg6tXIxi9abeyHieH60g9rRkj8iomM
y6LFEF0Pt77Dhojl95R9K4oN25lUI3MRPbsUz6Mz+Svxld/mO16COcgpin8QKskv3V0Q++0rxbRg
G6NdMoGA+KU5YoGXJDmOEw3i6NvWsd78HS1EE40X1WqcxVQwFywYjelEgE0GHc36Fwc0WyE4ofqF
EUfYhnd0+T9qLcCKCS/ySfDlgwKwxgX7IfSY2C+Z8uhqrEuUMDdWRBncyUvF/BjEZlGXqjEXX/0y
5MfgyJAUVJQTdNuQRzMSwbzmJriuWjwMInJsaJymkXyu+a8OBTra7N5CbSqTdfzw5P/TzRn31ohV
Mz6Mboj4GgGjaaDQ+qYnSwfWbGxjW+pp7fE/hmoGRD8d6L1BLGntGkPb9ha0wah52LCrcj4BQNOA
bWyYtj/v06Ig4I6O3MJDA9yw41r75fdYrhL/PsXwvYe+Lc/Upain2F6BpiEhgnj4dfSfY6JtfaiR
7ddCEov0aL1iENHifqqYDXN16nPNJOT3tCLC2ENUuupeRkzwvJjOj8TvloQzrc4cAaNsQPtXaK4h
2xRuipHPQtAU/frtgyd/GOrGWFCHd1gG33no3qRUPbIRny6D5khq11+Z+EDS0QnEjoVGbDRHUcy6
njoO2Eu4BIvksX54F5YlrNaZLR3kGTJ0nykzp+qo1LOf6w6CSGzyRE/kEfMeB9DNTZMQkOPN+/qn
AsxMDqNpk70LZtFj6dEoepABLbV63A4xGF8GzhZVA4/PEFHBmbbH9pho2iLJFft+Vsx+LDVSdiGO
8boPERcbxZdT9ndoltRnyjXwfkq0FzPL0xJP4MeIdyHXogwJaZM9/K0Vu2SnZ+i5ZLE0oZfjHzA+
dKDQjXXD0nuofYCZMf2X6aLyxQ8co/R/IVavaGliOIYezMTL1DqUyOswX9LNv440rdxvk6C7zBFx
xD4CevSU67sWzceX8m58AEFC+uLnHNM57j0aAgVHITiXxWbyMvou+fYnTMRhQTXV1Ly11wZDPd8Y
gsQVyHd+sKVlnYO2ql9+Nt7dHr3n8UlMed0YDoKvc1RXGJqkHI+deJUZRshQFqvByAtN+pqDN/yH
EHkkbPDBaHtx8KYPmP2dPDxYToh9ZvXqW0Ela+RquFwjt67ufR2Sis71KlyAvhylM5R+dsH4S5A2
KW+rEkI/w2RcP2iRgsF2PG8JcTfwhsnAsgzLkTzuNl15YVR3pYPcE+WxqBzzU/ZBkVcoomrLWdVL
QO4UfWm6dWkUqlWej7I8XaoZUVQzWdSkRmUBtw4GeYwZYWzyXpy9T14GxtxNA401hC8sV7XcRoYS
uy6QmDCEAmLHFfabNg0VWs5EIDlsUOlzvGAWRCJu9JTPverx5l05hKpBQc6Z4oYj53iMnbwB/vxF
5mGH3oHLFh6OeNsEPhUS1uxuX6TxKsz0O7+BrW6yFKUXwk2M+P5iy9UBfcx8Zu+UaCCsEZKjxBf8
aBwHQQ3U0CNOMusoAtHjdN/Z3Zhy1NnqAS/RRZYD47Qerk6IlvHf12xk/02Ksts/YQF23miqocCE
X1E8eRsYjt4o7d6BJmfBfLoYPA9EweeYpugSwIxnJhHZnBfRXE12AdN59kNCciqwW1a2yw2Nl59e
M/QLPrrHBHI4gYkiiwCvfsaXsVo4RRLi4vuNsYaeUNrFMvs+0y63rrPR7UAcaoeLcRcFisRFtc1m
ZF2VmQMn+3u+yDvW0K45YcbB/Hf5m3lVV4brNYo0rzboYWn/Ga43QCSm6BeX/mVEciL4r5EfRhf4
Nbyu7+4bkxG0dMjSU9q8YJgwj2PuqgE4+wA3tSGlISaLDBPLNPPpb7kFl+g1yUlq0Z2msMjHiqHo
BHkUkuR2ZGbSseWKJwqZ5S2hQLPdRBPD2FB8LS1cUbdP8peFdFWxe1DJJrRRA1Q9ICufg/kUHYQP
kjZQaGLIiFBPCUli4RZu/ApXWixm3vQLDSctKUkJgwsNRJKlnQvcnfJUA5n4BE9/yst15i31RUX1
l2Fqn3cwci3ZSdzdSqISywmbNGUbRwrxxQozbpVxo9mjXk6ZvNe8BXB+3DrnYFvWyHS3i0w8lA72
v/2bfl1+yJihnfsamI0A1X6dDnmUzY/vHIREMf2Xg0MpjzzBYUqsb1OlMNtLcQzMdgIhkGLqXQzg
F11lh2qQGLRrWIbyGBI1gpODlWHixh2qhT72ZW6FU0YBY1HY+EZd+TqP/rrWSRN7tl/MP53SbJ97
R7MPOACfPBI/bvrbewICwKXkJ+yDjTUB31Gi4NFrit8SysO/aVaKOgt4qz6D6WZrMQfzEn3T/kxN
YBDs3Y69lpZ7c5Fsk8UiyS4LFlkES5YP6Eo5+oFPqABzJfjT++zTYn/txgO+AT/T88IDNCeofA3r
QTRVOFNzoCoyMJjRY5X9GboLWwgoGK786lrBJhp84ECSJyDeUCGg2HZox7uh+M6JvcSAlvAKII2n
Ce2/KWwhthpJDiGjpbkYYG55TsQrzDw2QcADliZY3E6nLhRHjwL9TTCQWrN0kAx8GdJrXM7VSDDc
zUOaLuTZtmdY5t7q8AoKJmHY5EH8nw0lnATyVYeYAq0nTxEHSVFr8c7PAeCAledXvWL5mUWHmk6Y
gGhWtsvZTrrNPNHQ7A1jIXGPYTI0tkMy9TZ0hsblcO8K1YC1jQIR6MNyuAp+bweC1iL5J4hD4FmH
AGzEyjtT7LctREiLRl+Wu9iWtP2SMl35ShtYX1aMJykvUjka1zAnXeV5DSkkWBNQRAypyIC64iNU
O3V/AowKc2Np6nVHHx4XrF/c4y0PxyaW/nDXX09JN8ZXKZfzjGPmcBHkZTNX3pebRPj4w8Gvp5N+
qUkSly57jjT7wedQr8ios270EmdOxo1XjMdY7zMRQVXgK1MDpf0XFSCilRjR8Ctz8OdAdgd3f4r4
AMY66TDo2EPFsY0sy4k4GwuY1lIC/WT5utvBKRM94YyZFg1ta6kJqwva3Jk+bUsUzvdmw7XfIo4O
jcxTz6vtRcNumLJeuFEFFwk5Txa6iI2D3eX0gy3xhQcwmLiKY3ptadL7QQYkEhY1p0ydOH+CE6+n
oFrwY0VD5HV/MrDdYQfmQQEEPcJ3N3rYgzyglvBxkTP5tJpo1VXJaczfHRtPllCb2c+54nkiqlUl
QJdTA56DuKDuMdJMo5GWZNDz3Q64J6pXp5v/EdpbdJ/6hX14GUAsKyuFjLeZIaWHBZRJoC2LsE2k
ChHTV95/KIz3QnhU8YLfmcJlx58vbuHO4n9QacRqDUBVo6VFYwAwXx+AybmbV+kBUqprdhPGO4z2
v53M0OCQjL84yU5Ar27P3pE9TQPSCzXHv1E2vIJn/9FzKO6ETT1uT8TPn9InujAn/GbWkiL7aKuJ
9mMzSzN2ByQuUeA3JnZFqs10d1Y661OEUGmEDZ5tXRSA9kf6FmXPpQLTonz4lpfWNb3hCwj03GwT
E1nPCyDtuCjM5CBWAvgftU2F35z/UYupRDmsKlBSny9dnYYJ/zOIcOcyK4BllbVhP1K+BtiVuoG6
1lTNTon7bAC6+zy7o/DsSQ1UZMH1dxqWdcXSBqK0mIS6v9A5hZCsDCsS1cMnCm4mgs5BFmzZetBP
u1v9JCrY06xpfDX3Z+XNFJGqzerekWH6ZfP/8Zs4STR1MT54325LdxfyhZvysiYr1RPPnHTOBVBI
kPbVwfO8I1N2BLfpdgnRFp4YlQ5+RxN14EVDdMwo2P3Eph/GRpHY+VbaDMfteQ9cGmidz9x1ZEfp
WQKJQppAYw2aEe4sINi6U2+QutNPH/cgn4i6BsS7XlgfTy0GXhpufNk0dDBDus54d/w0Rsu/q0dt
AJGoXTg0sYqnP7TCH/TGlSNZqdWeZV56d5bQPqsyYZvi3N77inq45qZrbyhQMEYnOJxcoYEbXakM
w1WJ34tiF/DboIqIbofKxiP5IHYLrlnpAY2tRZ8Pw/cPmQOrpR/6/D+x+568hH90qL2utPoIjX9U
9d2k5JxJIf5fEPrWEAbquLjkOGMSvDs8oGyDWBaqh5Dl7aJfpiwH2eB7WKG3HrfAOTfaApI30U0x
MyuaKbEtoWiH3vp07PnpavtVignmD7h3Llq19ajodt1OkiXDQ28QMV5wT/B2dcdbjYuwVFlPSTTi
G2QXGxmx3+NzMUv0BOuDW5ynaSeBNBCCq48Ewt+DM89OIjqIeRUnYGwWQYm58vDLjEHY7hEPgIcZ
nZUXyq0XFg7dBYsveDB72gFlgk41c+LRDYHZByKfjGLDZZUdJOkk/sGddKGMpXZZ1rDaTETsNXh1
MhJqR115CM4r+252wwdyGcafwoWyZtcHGB040BM1zoIT6fAYP15Vf5vroI66O2GDpkSz2NiFctnf
iQRx/LYDIp90vsP3sa7AHzxa/GuWpvqle1vXu1qjWuGmi4OjPwSKpuJb0njfTipG0SiQ4KvuHlPV
c18RSOKv0Ms6ggOwo9h4zQ0lW4gu4acfpDONJYLCyQvs3uSX6GLVRU8nVU3RDToYizADE9DGdKDu
fj4tL28ahMn2rPvF+IBXjZdp9cZRJQYB0ul788F+1SQAWoY9JcMNG+9k8Pe3eGGj2WiaIeJ//00p
FmZbkJv3CqXa0c+0txlGdcxV2Aaq+PDzhng7aE3nCqa7WVO71LbB8QgVLrOelDmhTo8lCcE84bA3
0CqSMvBvt4k3JYZDs/yIMoAnz0yLSBAw6yG483bdNuuXdJoqrh69aBDVfRBjxABL0/saehauzkLs
WOvqb00Qy6J146Xy45zzV1pFCrMeFgRlbnHECz/Yo45YxdSnlFJkqgQiREFha5BC9Jhv3IU1x9aj
PHCYbvE6A2kzGcGpdDZasISTPkEuw3L8j0PDL1vVQU5Qyq1ZrQL+fxeeiw6lZ7RkzW28+GtJRagX
3WVIM0oeltOifykGl1qW+dcQc/PSV+wYLm45sbgCPd995HsFJUpskgptcWKOzIAIvPISax8bx24U
WpHEWBaNhbnaYthC2OX578wYQhgNxxiCeMpVL2be8QewfM6ROa5MXUY5UE3GiiSRkHIdhmlyejET
45ZSG4DGPNtUV6QUzdawahB7fkxxcmOLQ5hLlXd4z8NfsXbXy8Bnul5UGJ81AF55syBN9TKyoooB
LeBeF7yKf1lvg2dm3ca6vHQJ9wjkJxx6Kf/SLweiev1FohPPCpbnOifJCyFxomrlJ/1AvdI6oDoj
JD1yieNUY3kz3pVaNK9I5OIIAgI+hvdd0eXMlZcJSh/Jw4zjRYlwFRHhH51XgJyBREVHM1OI0E1A
XqgpOqV8ktu2RO0PjPXj8UnDS1VSXroCaZ9l6ZJbEkIrVf91pyoCaQ1Qqi0+mnjh95om1VRuEunU
+RKAsDFLPqd+B6AXVZuXI2+Y8QULJNj8e3P7vMV8gRDSteBBtA/cP6LsOL6lSVNsGneSAflL5m7G
bjTCslYH+rB5HGSr7wPirIeSnqXZE8buJYY/d0JE1ICk0llMqQK3pmFLx3VIOLdZAbj4/0tUy2Zh
QIKZIkGr9E3pMAj9Ixb62LxcNN6lMckO8eyXKpvOefaghdyTk8Z0G93SjcR3qlYn4oYOTVzE1Wvx
0r2P8pckDtVtMTJs+gjRnj54ROZYxxU7WnlGPTVAGH/vwnawTMNdLiYuZZvGI9I75kQsTEYgGczf
SWvRjaDqoV5HXnUKNKkj+fA9uvHEe8omqoSKCI9bcaqd0T9KO5V9z8qLWnf92ongTNyaiQGiGMed
rj5txJxC2ZlDlJCnhElaVkQ6K0cU6xSQWU8QJwBZ3VZRYdMiybC1mZxCRKG9sk3lT/rq7CiqmJj1
ngumvk0o+jH/qi6CKm2LmXO0W1IDSZpR+Ss2K5Fx9DE9PxHo9jIOGokER1WFCrb2e1ShPnVpU2zv
Y/TEFkNSBxL6lxA0GPukZme4AWWSCZqSab+q45xfsb8JdRMhbt2WpNVJXVTLbw4hF42mvH/8uYZb
gZBtHucPwBsDkfhU32qY7UpfjHOb/ZjnS9gIAc1VPVFDytpChdRpXg8iMoKgm67VODbPDBZZgC8c
NYZQnAnZANC5ywWlGV5hypzCzlUVy/qBt3OHKvwmEpMyNZFz/AQkwR7ZsW2z5DCciyWM8VGZtBBq
A+rs4sjKbuDvE09FBUAEJc0OXwjf3IS31FnDZOIiGiAJZBNYUVTIK4T1Cl7jxh/9+1Le24M2Rglg
/c+S28/TVXXbXXyAKfZYt9uZj5a5YMYUYjwvrBDwL0LJQUwYe9xChQv68Ize+Bs9+i2lOkn/7gjr
Zv5aZT60NMVZZ0BizL67WoLkGKnKC8I7Lvt/7N1ZShdR21NeWifK6PF2Ii/TpQtUN1c5y/cGXEF5
5pZTEzLHhNcs/37J80F+qtVvHjHF3R1IcBFP26NSlFHgw14ZCz02vz9EZWPUUo7Nbq6iOUL6RHiP
FFv12hGpWdG8Ke7YBt6zJoVezNR+oulCUIPULXAYEUm/Wab1vSFuEiaWxWqixDUGTzDJDTRvdUP4
/MFRm69vggpf+uNM04GO8Q0hDJDRoj8kt26OXL0jeFGwLXKb4Sx5ZayZNk8IjOArLpUeyLG340NA
/9h0IOuazcT+4pkStMzGnTJVDQbYLPAz16Gb05uXx3xRKLT4ud/0w4oMPNm5+A3rSjsbBoFAPQiX
iGTmz1qEqahD1o5PY1QEa8BTf0fbUKVEhZpa/5H5J1lkUiitfug3D/yNpQcFi2c2uyvv3o9h8THW
OCdj1Ew8WznUgD3uZprhCugdKzhYr6Pisb5SSMD2eER4YxhDrnSHUt/Woady6H/sDYiJ2R2Sn6Yl
va/AfUEYDHTWlBmYr0UtMjJBYukjBWEW9P0O4PBVMv7BtkBfMiIlcx87hESwPVByL7mZmkMlSz+h
sOMHnUR19tLG3/WUw3tcyyRI3TcvfTLeyqzkvrtnScvG0dAGtmLzpaN02oY2FnA1429fjlev6bnp
6GBSTjheyY17qQvGoJzt23AwO94NwZHgXvDOISGB4Yv5FEQ8Qw3mwYcqPEVQaiXiFzoQotOkPn5t
6KFPSJKTpjamVSzCM72D4L30bhmlzYGrl9RfQvYMWOQm7UORD1hhth++c7H5sw1dU507YvjZsdPf
h3M9tyOcJhhWuWdi/ML63Sn5lBZLGx1GMNb2dV6UdIZ9FRfagsAoUdlCVh+AP6eWjlo73jAXhbCW
nZicO7SEyGpDSZjHTykvHwmDVxFBfpxG2vvhSunIM0XOHvA0PhPdR+TJB6PyLEvHx+6hblK7USNA
aZFG3qmMjeFLm+5joaZhXJhgQw7WOELJEkzOHPBILTfoa/xfWhf0Vc9ajuxoy65h3/4GjuZpo+Fs
EXRWLzz5B/cbGVkzjhqrXkbPEhMrkNoS9Fwa3MnZKuT+GX8X4kbMsFHLeDLYO38SY1NB1Xz4ktul
tGkNFL94t8ZJme3Cz8Jh8Wtpic8P7ACCxtsTC1fUxrI0cym5L4jWB4JD/i5JvRXHZ99X1Mx/ipaF
Ej8OTdi1T2WRQ4QeQWEJolqPrItWtjm2FBLkgQxtit54Ve0RHwy5Ypa12fneSyYd9zjVgo+9NJMm
9Tzzi7nN1OjRRh0qpUxIZZEBTRxOiAHsxUCfCGGuleoWwLavMnZZNuNOQ2MRJ+UjxxbEfojOEb/e
eEJlW5/BbmiHZIoHwI5ALp+g1eXJM3Q7aCV+k6ljoXcrNUtAk3QXm1WCNIU9tXwpx3oc3GwFeaKE
nqujBzZHcnlCuPMgwLjwcvuHoL73d2gUZ7mWU+ucI8t4zs/rmFRFvd3YXB0qSn0z3mLFly6HhWiR
VkFvd39z61+dMJiw3LDlqizOO5sH8HYSaAkar+/w+fvckBRjOh7yYQ4TEaHgOHWZzLXK/ZzvCC/q
f1TEqFTN+nWHHmI/C7E3q7UG9HK30rXoCeGyaM53OhZPs78iZdjWiZAz5TBJwmaD8acsYzzRRLNH
hHobaL2awuX6wgvvoyMcviTZOBjlpLcn3xCPRc59EhH3wPMVjz8olrnrJXvbQT+qXHq0QxqG31q6
Ii3jf/M5cYsMQsszFvg4cEkhEj7HQxwgPei4do9PdrC3I+VmaBwL5sUSDoCx2TlWEggvyz+ONiyb
91gxHr/ccPPpmQM92Xv86tbFzx3FlZ6UvfuSYJMdAHvRpFb949Xi/DZY+QTfYp2NMavP0C3DCBZy
2pSqNmgthvXyBxYx/NfFvEeYBmVkSWsSSkbh9Y8fwSJ3qt9dJjfYWSY+wgzpFWxN5jtI1cwCg3Zc
ogrhCgXE4jW6zVqsz83uIL8FKi36RLvPdP7c9RIPwpzt3KQk/0XXc379H3wzR8Z7z2PvQsZ//DFI
vCL8DIAgcFN+d8e5EJ9A9ZmvOdXLr+Ja+3twZP6eK0353o00ARMfVGky3MrpDY4p3UDhi+//mKd9
DZ2VMaFCY2ra6sfMwShzUo6GnVvMEQC871M47T7CDCOkyXDvA96+ZsnCxA76ZzWAZ5meCW7AvFyZ
aoIZoYnruIbFwpDtuikMytOxGqClVdZqJHnepkgGy8JJR2dt6XLbV7MdgqDiQlhSXFQ/lmzEWstd
WDjTTxufbMX7StKST88lwqE+uLFQiwy7xCxg7U8UXNmRswXOxCNQ8mH+xp0CwFycA51uF3nJEgI+
h47dxXaWg+hTihCGakJa8JXxvzItGfsxK0DB/JmGxyiFqlxT5jEPKMxbS1Esr7TVKYnCDz73KUXu
lNcmV6xKKAEVPCu4G+v1FTUS/RSkpksNNtxBiwpe7S0xy7bnCgarTMN/yI/Z1OvXMnXR7vxtsU7h
uWnG80ai4g9QVexgYwrnAZHYftdqKVAKR/6CstgaWlEEDf6Usi/7yV5Cezo8K/tkUuO5etGYcB8N
Fy/gy8yZAw3VpvB390eLsjGNqkVi7kcDMtvagTi+mYUAUtKhphlbj+EyDc1vWtDt1wAp6SaaRvbG
n14yvy+y2z/y/zk2F3RRxkSCZLWARdJU8iUdwXUDeb+rhzjAYAyXy0K1stGagrGCEdstAb2Gmn7K
/K3NW6ErQ9/yz1chli5zTwUfmg4Hw+/pKzWKvF8wTpxsB4BAmDlkvIXsziZfsdPYqXaue2iADDH8
U69x9FUz5eEiRbPYeMD/QhJGrA8/nR5ZhN7TaTnwOAR6eIc4jEJCnJ9v4w11C3/KeklZOuK/wCU2
e6miwD/+/XJMNaDSzAmh1p5wtL3STfCCpkxa9ZvQgg99G/SAyY30JC4bwRcrxLVVdsc38SAHrKAx
dpXGQVp5+dV4wJ1dtiwRZOsSqYJa1BRzRkW5J60yhX1nMYsROweRvWVEPqaAKsWo4o+1iwoAWHKq
fGMfe+oFHi+SeATrk/JRgys9suUn7RrmYhjf9WmMMO7gAPNxkuUREJGANuQkHqcxr5Ojm4y2f7ek
VUEqmHOPhxZDzA40PoE6urFIrjgXKIK81zE5KMHE+PzSPEZ4wV4cjR9sYSyDUvHHwcL1mU1I5Ymm
Vyezxe6n80V3+YICqeTG3B61l1UOoqZaW3Qmirrga75RcgwGtmKk4KXL2F2NESNJo2diwtTf2rZh
TaRYnRlCLN2swr3g2fB74MpOIHPJDg7t33IyoTpNvJYCANUtxOLwKa7L7js1/q57JFOsXFskIOfG
Nbrmty2Lbfwn+ZvK2IDk5APKXETKTjt158g/PVLdfN9uiCAGbnk6ylIgh073aQthfdlNQYnx+728
FfWGOt6QQZBBLZH/DIAAaQgqrikUrQACXnlWJP/6+YsTfeHsguBNjojmnWhQsuFr/CF7zsI3LSwl
rITQFZiGt5Bh9b4p8RjmncXnk6mVUeR65mn/dCOd54TGC3mVg5N+/a4cx/RAjHcSdelZzykONy4i
xUuVbbO+9ZW7nL7EeH6r5aZa7CzkfCYix6LLR38CFMYbcvu8dRphEYNkmDGvrdXqgmh1Wb+UrP/J
qrq6iezBWpHPCOUITFINzMNs/WwyPGkdw+mtmHuu+LteN5nd4x42AgdwaabJMkNxzKtwcYFXNQEK
CleUJCCNdT/7fjER6sGb/VCfX25d+bFqFOKSsI4rMvQWfhOAaBopytWcn/UWvwgXdt1su15hZK0O
jPqFLL7uXwbXYHQlIiVw3KV5sBn35jDxSVynsV0e/kQjpKMC09u/BXv/PjOIk0qz/v2nSWfHZ5PE
Esi/VOjeZLGFatOWISfD0XhkHgIC1M2DJnt8F46J2t6r2wBFbr7Dq0jzqTZCUvFFktaaH1Mwl6ei
AEepeNyX/Sqk3Df517qoiHKG0v+iLkXferbFmD/vXGjtod0yrar+666gDArT+T4YgYO7/sSDm6fX
p8avK96RxeWIBAvJbZK91mebT3DcbM65icG+R3uqFxVNR5oH+ZQ6vS6dQGUSxTBslRLxxayuXc8p
Kp9CxOhs6ekz9U8Cp5KiUo2HatPQ4LKlMarlRUd7VTRwaIN7PyPA0YD8T9Bq/zvs9/KNbWEQTDaw
uFM72F7ScEhhmiswWSzPVCQb6CIPMrLc3d12PjT0GeCGoX+Zs8tpLyeyanePxRVLy43CHl9onsu4
NrY/gbL3zeMyJaGpow0fSU8HWOOq8zwZFytWDE67NSnXQCACE5ySvQAwZnWzYKYHUMU2AhFXb0TX
lF2oPdV9tfcqM4YNA/AznBXWiiVT1BF8uHaJKpGvw5IfbImO6FYAKMIM2yzzEG0F8XzY6qSPPgkp
99ISqQOaEXOgXFzfQu0qMCCvmDQca36/yxZRBlyGd5solhYg3/VHIs1xwb4n8dltGrvqnqS90aLY
9tkS5jefk1/ZRF6OvsT7CfSGfvz9EFyxOVWDSYjrhBrV71InPiPpXWYpoonKlpVeqThVk8yzriWi
ZQqWrZCaP72GDSsAyLA5rfBOts0Vy7pfXmYYmXa2DLHPoY2Q3/6JewzZ2jFsdHf+xGRTzPyB3hWI
okevy2gJbUfxn4/farxZAArVgeoAf7PIS1jyblEuBxZgQln0p9Pv2yi6vSMCjRpQi9C9KuMGYO8y
lCpd1+ZcVlKh8IA7qNz+QeLssgv5q4PiXZF1gREa1BpzFbxdN5Y97FnSxtuKpJ/ajK7J59yeKWr1
NG1KEr8X+a9rxUacEWmVRPeQmvC6XQsQ5BI/eX6epGjV809NHtIi6SS00qynTPO/5ysNWZKXJLOs
Z3QsZ1GTbNZ49Z8nC0wWHmlOmk857sDFYSGgZNS+06rZUM3zU6vRcxWphIm31eQLgqxa4z9FXeJW
dZOmcp3AIhFdJ4P1kA58U7NSNPigAn5N/REM302H+6KdkY15wxHdjwwyUI4W9bZeT2w7Qh23+YFI
Y+Gs0xZ5jTD1/Eyjr2nIYsobyhkmMdw1SFQZJVszUJ0BSsc5nIiL2uH26b/8MkTeu91t47Cnw4Vt
70fRbeBP4QcACaxLofEYS2ygFwwxfu3bUvZUeDpfAqJA1l8p9cbBk7FR3CoQdM8VQ5ADI0ShTzxz
pC3MSOPt+7E6YYsw0tRW60WuwM1gjZsuSpMbZTUSnb5ys9f9RYsIB2ztla5oGuSRt98U8zyoGpMr
r+cz2q0VXyZojpV6JDueeRdlgQrj8IRkBgzbamOPx3WVe6AAohrsEvxDMaI0y29SvFke5fbM/8YL
3GCs42NbXx9IDW4zXoEFStluBaSVEseIs/imLsOUwdT1vpKw++80E+SFtZcGUV+dM2oHjXs1ypqs
ZB6hTq5mDvUmz+VFx2ouQpGb1YRSVqG3amp5XKZ6+iAffRPziCt+ARUG/N1K0nxWmkZXDeD1FU/S
KErokKpeLsSW0/4JJqDTHuIpsG+9/tobJKbAmuWtyShNnPHTorjFZOV94y2h4kzEJ8dd6JiTxFI+
9qJbxhqE/4H7GCGng66LpANFTqvK+RIVMkqePrwDRBYf1OD5ct2/hqPw8eDwnN+AQYlT5wdanW0R
KkzoIDw1SxvUc78P+Z3ukHaQk3S0hVehwhaAKzUOAD/URu4CmFiKEA8po3HVngEzuodRltLY7YPz
DipNQHTfRudl/4PfON0HGo20NuIeCmTWyHHIyw1S5k47koS1jdnLU6Ssre2dBSEk8mRpIaE2iVYi
vVPZCq2NZEfud7x87tem9/SSiNdsLofpQJgAWqje+4jjkoCBkPbddUAyNu/N6UaVhmMWvJD2Yckx
IWHY5CIXggbyHXffBZZzp8D8EiPDeuvy64yit1AhkpXUAn49ACXFQg5XuQ+huBf39DtnHta3f4Hy
yQkEzeOHnZEWUtSVoOHgtlfuCDerkxKPcENvMOeWoGL9oyP8RUve2S4guzVEheaa8JbEEHaJqWQU
5BFl7gwEASnq/Iu8QjNpQz+KJO9KsSigErPf7ScvDkuCzP1FwKDKp85rn2CB+UaawZ3CZQpyT5BQ
0E/3MQ8EFnTBzQMUROsYP6x/wjoMaE8rqPt9joPHyXF4ytnl5D0r7yNIePGQrUObArZAHVniJ6T0
7n8mDlpiJUAKpEhBdPnxCKBr9e7uLn1gvMWZYkWNob7uBiFnO5UdBW/lWr17gvxgfiG120jExzhZ
cCrgGYqxkCXhXWRCfU9MvnlApG2HEVGLsMxo1tayNh4usW5EhbBN2bp7D/OS+oulhQgWeTjkDu1z
PPsNk/D6KEZWt/yn44slTOFiNdDlD0JjcV6DZKaFFf0IN4YUNcPGrAJTNJUqwDIo81SU07detJQI
aDM99lZx6jiGZ0NlvIbQ5+uaWHlEDDtpgJ7OYFlkBxc3bzEum/fvvQnJM/gDhSF5i+8UiWnfOJH2
craCUGRiz55c2CYnoHf1PP9aP1p6UiMM4aqqb2/Z0rKn4hneLktAApk/g9fPFTTx8WqqIcK946Mi
zju/UNBKwyM461pMTxTEC5i3COmiTKeSOT4diEFrpArxDiLvIsLxp+hPhHxKQLGy2ARJIrd0zTfU
R7v1RIPpR3adoJc5r46T5y1z6+wcCaE6d1zRkT60pFgQlcvzyNdSHk7MZfcI8yTaF6V0gkMNRUB5
1N+2YgqMJXFkZm8K0ZHGXU4NGEg7XLecBwcj/wUhIZEdPgNGDWuHLwhlwyA7MGj40xL6VuVWzmD0
eIfQ3rA05ipCCWd4uVArbAne6QKAB3lmlNwALGdfF3IBTJPFfo+bAD3qD4VqdH35tgJs9yT0JOyT
34TgtshkTRwB1oPSunl+VoP5ZB4ZXYYWWv+tLeUGyhoT5y25CZQ1imNkyPqPJSkn3dmlIb9N9rlA
Gp4qq0svlbHBUl2UdhJzx3+YEgltB89RtVpjHGmzwWDW4QtU9S2m0rEiIBKRbI1cdno2ZlLvYFgc
GVPqcqJlRSMChdYSsysVTYAf1CCw6aNxEIn7SBl13bazVQjtNNHZLeQ/P4JoopaZjtXraHrEph5i
3NwTxAqdUrxUrwHOv2OJc8V4eDMRnQuiiDCJs9+OPm+c79TPoecYep1hZYb8k0E2A9umxr3r3VOH
KLKWPlKyJJD7UZ8xDm0TyO3Iguvtz57maOCmXfA9l3Xyigz3GrvHr6tgqXRkNmJnZNeOmqZhja6y
VOkjwijOJAkAdIQVldbCukPY2EvgFPSDTEq/eQa8XaLBXuepdwu2XaroFCBn3Bku2F4tKHpY5EHV
egVucGqbilQ7qj6hazo2AyTP7eil5jsKwCTA7/vyT13ImsrgTk0JSPmFguWQnUH8FjfEQb4C/Hoi
3BM0zEiQomY0gCZryOysZ6ePeF5BoL4yeXteXhKQJxAiVnkYq2T5FvPR2fnCAQnAr4QWhKe/2uWA
1rtfnxqRmMfgGOBNnXEuPSxIb8YZz1cZi0827smOusAt8MvNWQ1tKIFlinyOE5vCMVGjmrJTaqEU
VgppZTMltu1lNjkP3q+PB4pYF3+9DEzEyLGR8rzl0vodg5TgA3/DUdsI0QOCSpH6lKB2AbC7uuFu
xXsJqHBpwiBS978GQuCZbkPvWJI1M5G44l5yeLrBVFMBXws1ULwvPn2mta7/HpHR0JF3OmumoNp7
72cbt/TCFe0f7vRO7BS2rI6nJAIk8d4I+c3nPhJESKCIq68onrUo1j831fHetIEmhvT8lO8uLfeJ
LUImGsZJF8K3AW6IqsxhQzoQSRV5stXIobH2kNer2Jlu3n908P67vD75N59FHGU1XjqsBhmLjoIq
4GJ0UrqnsFwdaXJhvUooSn4MyJwHWC1oRdBQhXNwlLmQOGGtkfAdKSlvkeTdzB7Oor3/7LrMfXO+
Un7lhEmSz+NC8xWXDJkq6PKCpS602Tu5xELScPfYuvud15og2yRa5yYlkS2evaIAUJ8u6udrxH4I
kE8YmQsrPdgcxh7BSO4nlMqnKAevutk8DmvVVhus0snEsEi31QMr0m3lQGZ+l+IzyNXw3ucK5a8M
6s2kKNIHtIcQrtYQCVJNmwgkeeDFyJeROYfUt07NT0rLD3zpX6RdTuBX0L1QD9FQSSwZUYYNLZzQ
9WC3RPa9Q5YHE1xoFue3RaJMNX4dy3RD24gnnkWvvT2xRjIhe13drCNFF5F4Q6wmE7Sj5g3nMclE
1UhCAZ2FhkzsLzKrBzh97B3i/ojtr6rp4wf5pdKafLF/E6iAFBWxpZBfSPa1lHbDTF4gjaowX/El
w08N9HOcY1gBLECrs9lI54qs/n3r8XHvPJXng2OE2L/2rnP/RyVj/QvS4bnSscXFksFaY7552WTB
+ejBVPQRM+i0Z74gdrhdcH7krUbFR4kWdxIjXSJcQR/o8AZ+9zKlyJLFscnr1MtBEoJu0sHjnz4V
eLyr4JK8BcvX6ToN7+Nhox/zv08nkernwqxo/sKGc/yT5pLcfqFFY2vocg2cbWpM81n1aabhgjNX
P3KJret/1iGU12Py/F+05Yp4SzuFbVkdm1bqX0MnC69R2Ids9tj11nMbV3rH4nT97wfi6fUI0olW
wPKVW3Zqd9q4PUqt4dDOE7w/LbPzSQEd6xzbvWKNwn+UoVRUTPPPzwbgMJT+cbSDGFnI1yUlCuNr
ttt0jGdVXM7MOOGaeSUiSb8gGGDgHe9QGTBeAzVoBGUTgOPPRr7Ijq2m/AF6OZPFdNUhMvPfPuDN
MhPxKKYonoZxfgXBk+07LP4Cg+pLFlsXBA3I3t4vRn/Avpl7PWlxMdQ+iKf3EwQiPaOvKgHxLvMH
ig32fSCn0AS5+Vm3Hep4W2DKRHWKYb8WUuT7vp1z9pbP/qFwLSN+erys5N90AzbMCCjEojAqo0V0
9rEMqL7T3n3oqbzQCMARAw/Coem5tYFEq+vjXshrEK/qG/505cu7/k0WTmV2rdAMMTcqVWaFJrUn
SLsD30/60ocvZRmzQfT0ClISUR3hdYbCFbxbLNecK8Xr1QMHSb+juC7ZSyT4TUEyneMDlNUluPTJ
QNtBpU3aODRR/KuQXqKOeVtg6obg/pvQbdANC0aq4z+/pU3EylbF2ncLdmIBU5h8lb5AJVTsOR4S
8yeMEcz2ZhU6nvCP3zfp+HfqUgP6O4LcAlZt94LtiGCbIXUkRy3KkpA5Hb5zo0WFRY+LcB2O+wn4
/SoYOrowybKfwJWk27DKVkf2H6FwmTvLA/cUTc83odqVlUupvSfMyA43gnKksrmuRsjNrz50Dm16
Q3+Uk/b9Lc+6oswETHiCIoUO23QcigwTFfwJrM8UY/MHv6bd/0nGlDWfGQrrPXmRl2XGkwtM+MHr
WTSaComQjMDz923wi87RbAYMoFsnvQPA4e02JkisYLIvLJfaT0wk+oLgq08I1UrzTA7ZlXbS41GG
Uh8HW+zpkOnv0eFRz4C2V14Ej9x8IgaSLFI0N25Bx4ZH1b2tPKt0+8b5JjlWMQDwZrwuWN9jwQ9V
HywRwFiLtlljJNKyfMnzrm4JpUYdzI/rx8UegCf17CxXGNGTvSsKX8uBhsnW+TtwPiDCx3aHS2SQ
8ADkpaMlDVj1A52Z/NUmK61zdKro2Rr+EODNNKOF0E9yaR9cTymUsgh/8vbLm4fHZJGfl4P5qp28
p95hlW5Vcpz4q1+stLF9TnnTmuaSiCjjMj4KZkoh3fwf+pTl0zcrpJneTN5TlOzgUTYNUgzGk/BI
RiAfe7N1rC0qFa1mJBcWzErVen2nLVoSxf0WfKBhpnJ+eitOHZd8Bqz3hUdpLTflrY7JtLLP1TWQ
ePNxhRAWGLY5bUAwZOFcx+st+TQJYwhfPtIGDtfMaL4AQzj/eQ5cxGNE+D8HnmG5HWYgQbyX2Hu+
zoHUn16z+NXBXtYaV2zTPz3RR9AqP46FfSI3Nansx5ZjHJtVnWBPhnHReLNezlPMYl/8QDK5qAcZ
dDhz6+rm+Hc8cTum5rlnrDCPvlp+X8Kj5lUhvyVNDhJWQaa9xtAelyn1TKVzi39YHU3Ncvko0VeR
QZatSTVHNjjcsp/RT9KD4i6zwzF9HAtHSAIUF8FAH8DNK93xgs1n5o5WKL/Km8ZrOSL1xiN/2DiE
GTmr19Wz5Is8Vtsxw6Fjf0MlKRvHogMpK/EpMAkdI3qfcqVR009Np0834lXdKIhW/wmaozUoT+4V
VZnrv6ALbnZQIpEK2XGl7y5aXuqzd7oiShM6TEFnTVz/GNQih1dYdFLzdbrir+O1l62rmAxdzRdM
wRItbgBXqMs6KVl93j/BwRHo5M8oU49CNfXGTZ6HmHw3nwbmcPKCatBpnqmT23zF1xtYpgS9ocqM
VX8/UfCgqmLsl1UOUyUgBEQ3LBCjH4WPbCWwDhnjFMDCfN+/UcKJWWR/y2tKmiY0dNLFveWJ+uYF
JgnQzs5uunLyYZQLQLQs8mu4t/y16IzxWU33NhgmKmqeJNAUGb9SQkZXkR3iETlxaXTlm+GtWv9f
INbFaua2eAOc2n2/dWMqofkAPHaPCgpyhIoPrROlV6Ntzr4yYmVNSxYLM+evSYNhJaNewC2B9LBP
25bS2oHTyB3cNW+zxEqRL4RmquJ9CxhvxC6pkrLluNNQz3WSC736yeYXLSkXlr899Jsqe1ah4Qqj
Rg9pemti6OECcJ5fc3Xq5Ty4PynkSMpRJKUR6e7OZ0x4KdHG0kUsYckscmoCufutewJnozi7J2Ky
9wM4ibMIMaL/d/0iKVyk7SQz865ySzrKVDiKWtpWFH1zWtvVF2PvyMo3Tg/yLhb1di+Ky96JvMon
ZFAL0rAPDQaquHOi/E+Frrxhex6e6jmUeeu6Qw1kCxARMybmxALFSHimO2BVpf3RnF7x+qeaa89Z
zwzQiZR1AbKyV2gcTfZEw1oEBU2rnQj4B+f2DmoTjK5sMXDQubCAVHXB+1wlP/zeAPN3Nn2z1kfY
zUoxk4swFljJrOv4YQkm3ftnvyb55uPh4F1u0M0+wXnkYqyNPE2+ab1nAqpCp7usgwj304FhD4BE
pIrWHcfuYrp2nUycpr8sjXGW9Zm+I0YWjX1wa+TPzfWGDBjqblVxcb+4QK4b1OB3/XKYMRNnQ695
8TcGYFRvxQuC0QdQ4DOwu2YipCER3aDVVRhN8ILErSz5U3QstYaDUFx44aDqWh+KR2mXU84yK7Ca
8po05b5C54Ylfu3l0U3di8DTyRPFcCKuwF5eLfEHuwqPdV37/mrausondOzreT9hhCKSOKm/xAXD
GGzvb8H5tfGqvK7avmBowsaOERp+iwVi1f92w6dHC40wKFAr+OBiJ3jQROWX3DpXvAmILho+xTrm
W5uVqwRQ1KrstZ5o3hK9gqpMKB4I2E4DSl8T36rFX9tDQuzK1WgnPWRfcf50fyfttf8k6QzGk9r0
FVY40JGiU90qPCHL5e3+7Maa7Y52wvMzeQeHa0eSS4fxvfVt4nE7bgRZtE1KAxcV+e33LA/1aPBO
kZKsImyX7AVnlttibHI9spdYZbqmal6+2wel/i7UdKgpvBLB9K6ftD9d0qnMHzsoLL4NW9HjnY7u
h+olheUSXGW7GDQ+ZtVroRXUCf+H1a43bhMgAp/+iNrVf6tkMQVRsg2rrVVGS57XY4tyk32vAdN3
LHeyu3luZ/n9YdPWyIp7LbLNwX+ogFBEwx7S1srZaE6uIQjac6+T5upYX1TSaQvFx31e9RZ2QmMT
JC+bQmdVMM+UFE2SJfxXDTa2an47UZvydhF1+9529KZruVTHgBzPGfDfvOWyAH75Rqmd2PRu1Dza
lpm9AG1yPBce+B5tUNPwrntPOsad1F//Qas3euS5YfqK7W7RNTYQETx8reeLzSJSssvMKrS6pMrA
hbbt8dbGb08u1zEp65tUBtP5/CRwvyehTa67+ZBIBtmzWsWSw3ii+GagaN88pINuELkFY7XEWtId
WI23VY6iLHyvif6jtrLY+M/cDM2UjhmnbvIsQWx6WjtAWEl/dLC1h5CHCc8z5ydErYUxssGQeTw3
YipCWUji7wCKmewTEsP2kRriSf65GPgO3pYyc3kOD/UWlY7hWl6gP9Hv68viotgf2eKH7m0+ita3
pBh1TVHq3MNr7HfR0zGDVFgk5jp5rmU8W1clFoBD+J13BKGNPTT96LZc4BCui01GPx530m33QMJr
9BxAZbFcwlU8hjqX3bH2oMhy5llR0LEI5FIAs/tmcZdJC2+k3ZLmEbNFtfHahq7fCwfLbt76nvWx
g+kqbldZg0iR1DW/LQtEiKGmziWtMwP5sNdUpiOaRMm4KIOvSufJVFpK+S47WI8zLtTRpnfgzlpX
lfFhdO1MyMZtG2hBFT1h3ULtR5z1XBGBijzN0nJmKrwvuts9kDpaKVGkTWOF93IoJH5IzOVXincC
f6arlndse+b+jo120WFVk747Eh4LcIDBTGc4s0jbNwtyqQJphGENbQimYmyzAqr3n+/aly4vLbk0
91mR6ItFjpI7fVJjSdjXGbvJT0boavBBvIG81swDkc8b2HsA9mKdtinPHcY3hPW/EX1Cs1KUr+cN
GohcGvPsP5tZR80ESSjYJWWQyyOWuI0jF7kSX7h9s8D/m1ro3v64beDkGGq9HAZ4HAnQzIUjB7Ci
DqY5WbxnDiqv0gp4kA8jZqDOggKPVlUmm+8bU4Xh1gxhstfamaFODWu6d94l36m4AMkTyF49mLkS
Z1M+QDo4e0GqaIzY7BC1LrwbCDx/Dnq12Thujxks6kuQIrEjWFQwDqIPNsR7x6JspHPDfBZAAjqb
dyQ5MURUhqx9LOSt28VEoMSjCxsiA9cGAqfDf1NdF6zwWUrgrqlPIwjcw1bI92dNnrZotL2vG2Ma
2Kw3lWTctbOSsq7JN0aRrbcTFAf6CHUaZqprrEjRI+rx7Bi3h8PW1R/IlvST0RveqvF4ukR5+Equ
wAib4vEIuKOwZ3LZgA7/6waENph/48c7bCehIQGuW1G7qj8Z8aJEby9vuVm5Hgmv6P1S8L1cSfi0
d7m07y5AXBwBjIjHueeO1oC7VPLPp83a/l1To/hFhdzPD/ARhG8Sn+9HnJrTvjAiwmP2xsxzH0Gy
X/21uE5gU497KZL1478Fe9E7ufQJXSOhxGNvYpW56wgE5H2Pby7b+NtzTA4ug+no/nHty4LJzmb1
zB4OGBjEjFDcYNpJ2rqSjZRoiBsef4SPDMvfpILO3uO9I352TBtSPmd74UPwVgoHtp+JLizCOi+s
qxjdINA1zeTyjnhe8sft4uZUvbiv8QvPeCfTo2fard+8Om0fp5YpTj42VvHz4nlD3gv5QmaYSJhM
c+/dOpz7f35e924KQO8oXgay4XlTmVM5cNCWU3xJ5DGXoyWMq2Gw9wT93pNKBDsTrKaVeyqLorv2
Di3TlTBRLxhy0g4to2/0BWr3kz2sYiEoP1wdVN9HD3pcA6F2W3fJfxJAlwFBN1TiVdgAVlAQnaN2
m/ynN9lYPSoo9h4+4kcAL1bYi2lb2H6dabPoY0H/ji/SHk++ExdKzWzpA67OL720Lnytr5CQr+pB
pUWXndzld+arqVogPK9NpbTCB2INM+P3kJBVPTwflOeVhSJkhXVDiVt3b7ABbjDNls1Qgq/qDOih
K/bcaLlRCqddFlNVJyKAWEMdAC9UrDN8/nnAMNLqt+x2w6MAVc75WhnfI5e6vW/31xkN1OF79DtU
QKhHHo3h9Pvo3cz6jqw7wI5fPdC/dhaXuGxC54TzLpYNYZvqrmxQ3ckwSRyqqXoWeV+7YT1sKsnU
nn99Zp/wZTLAJ8yUBl/DrVnxgvV0jqn6tpuNpMuHkMq00w64f8LNYylEM844y4qhe5LQdox9MPvX
VE4fU4INLDbXAYpMnja7ckbdkV9Vn78/4dUKL9n4+lSkPmEoEkg+f+LqJComXMoSHXwu9prG5Qn0
1PJCOCg12r6R7/0/UHgkIf1eIpDIrp0kC+67Z+K3Tyxaxpl1UhvFR4wFlbDZsS6c8l0TGL1WvIZw
TDfq7Jl4VexxgVIq/lFzuqV6O5wGy1dVCmHlOJrtaj+p4q8rUkPLxzPmQDHDYsOqZlZ3SbNtmgWL
GYc/B/lQiweBj+XZsReFG0bxbkLowVWCPt3rW26lu5FHTHCknjo+3PXUI38xmwjTTaYo56hGBMOI
ycNSACHq9YkBCfjVCfTJsD88ZKRdLFxOh72Bqz5dJi8HUcvvn8UiApOfB66MviefdoeI6fU+pSwv
q0DRgq4n2zsjTc3PK8agWl/wFJo3ABN18qScOZdCZLuD+YTcMF/9CFmYVE2/ndYwOgyq4Irg9hmm
dgo2Jd0SmNgVfM/L3sz/sA+AR/Lgb0XnXqhikumokPUs5tWQDRMHjd5rRxF6DrLrBBZyP68A3RVv
1bClDPVYAFJ9JYaU/tWVhG4xAkodJ9JlGSiC6lLXasNEBZuW8kIldznlmwyIdrednDhupw1zW4H1
7luU4DFw5xC2yAnCrzFteOtqn769ZuknStZwqbn25jTaB+Uy2OVyQ3ntzQ/6IsMv+RFHQmWcgIrN
GQpbtb3F208RmyikHZe39vtxhUmPNiKYmwcQOPrwwAQXVtjIs9EtUEUz/VpprubRdtqNRYGOnLN+
Igs9ySyUfZJC1yA1V8r2GunLHJjB1tS3JRggfwZtjgnNKsoxDcWxbkkaSdRxIjsOn1Ea8BK7ZOc+
kmlxewWS7mTVkQXsY3h5z1qinKP+T2ODh7MqQhpppkw6KbFlFiXqwbiyCYOp5tvb443gbn7pSHLx
QmsJhQX6JLt0Z9iAWwUZj/I7R+/ws2dnVdO2UQglbLhttZ22cZSniU1pWIqo6AGA7Es/9AEC2iLn
SPtX8Aj6fBrmyZa9paoyjqZAmoGqlJykH+MWzDESML1RGK9N1X76kzKI9DGcnUekm9/4gbsnI5OT
565uNtzMElt8jK12MMoGHSQ/nKIudWTFr5ZU9HyKFWXBXGyuFXyiuGZY37oHo+PGkQrx1m6CSx+C
2QW45WsO97QHLolYpbVoTOam4GQ9w+3Tu0j3v6Aoo7WtqBaKFSx2CrTNFM0QyZ/iw2fWAM8wA7N7
k1M4Syu4MROkO3Slnuwa5QL7pi0w6hRLJscJTDARydm03STUIyEeALDruVESOOS1VIu7NEdVYe6H
aCf8pxoCUTNEm2f0chYIb/MaY6ttdu4dOqsWPl5Qr6MxdbFyinLn6d84TV5h1rj4mi/1fPy7Pa3m
icitkNVLBMrOuRixqrOzTt9EdmdfvN+kJvi71rzGat4eOSrZjNoV9pleH4CZUmLECRk7U3/l7vdW
5YT7REXpXV/Rw+6FIp0qmiAy+2Ny/TQXGp2GkM5mgmLLXJV7+XPIVPI42mZlMVcTFW2xXrDIVXWn
g9aBsXr2pURSh/BwIGJyW3pNH2jyxEw6C2ktzSvr97yLfnYoEXfFqYDZL320k8NuqLvsIjSv51wf
bla4vqBOACjnOq7TIWME5Gq1Ez8s2sOzD+zUKFbDBBrHo0/3f63KCSCtP1YJm4DMj/uHjCqEAxdx
L63Zx7oV4LAdJg0OiH28lMt2OuqmgTZUvyHIRMLHpnfL0fmilc/njZT7091HQad/w/AJQIpNpArt
yp6og4xeWDPmS8i+S8KOuuUH6XTNDph2+F27wsANmWdYtI7lmP4nGwGsF4lVIlKaN7Mwu9h7WVX2
WCUPk+vaQJU8qIXfIBvTLFD5+ZcryAVSapokM8iOwmjj/CThsLc393nu2ICUQP7B8fGUwf5clxc0
Xy+iGYdrMItpW3MDRPdXtl/tkc7ZrK3sPv7Z3hEue/qB0FFFOz0uoIJ7a/HbC/0H3oKQlxj5AQ9t
nnIkyQbLfewwRvP2F+ht8JmQVToTx9Aq0TBIAKmn80GlDPrIgb5YD+ZJd9Ry5EZGMoLUvJKPHrp0
9tlszP6Z22AKoQH+VZ8pcodAdBAtrGk/sN3jWpu/cxjv1vCK0mxYJ79XkxCCSoer9Sh+q695lDzJ
9DXFlUlq/KXxlAUfmx/FO/W0DH1Mw66UrN/2mN5umamfTc9nQ2LXebNzpFSfgCdw6aPn3Gv50NBG
J2SaiBBKiH1oy4qeSX9CSYfAKHjpnIctXOyVenyENM+CbXLysriSjJsHAwPmhQguPA/4iifzfcmk
Rgr9/Dzk2VC2hmg1tsIMcEUJMGL6Ut8aCaUZaQQNpN5GEInxyIDQvDg/eH+U9KjoqHelIqDaqJqG
h1rEEyNlH7AP5swnDYJcY7ZGw6/neftX0oI865k6lMHNaL46FU8oKXKaoATZM2gmMnNTIp9dMdxP
8zxyCKl/VsALdBGlZu8ZFa8Xwa/8rrddn8gPWIm+nZLDNTmWENHxwx4a9Ljuse7uuOg+Ecbp+6Gs
zoywWnTJdJFJA4NJj1K1cS7QAvXoTrhZTo2czVMIInuPLwWw9BkXGj76/5XNvKjRCFMd3JDAW/Ef
fdMdcvdUT7Estq04LwXaa3Mzu+/wx7uYzU3Xrn8/8iPyo3c83Q+CAUL1G2j3HRdqLqt1qvlbXQ/v
8Sx/FFZtBOZmfj5lXJfQHQcJO7DbpnXLLeJwyHaNqALTiq7/tv4QtyeEAxRVHXgfeqYUjTQ6l683
I6FLZTPJwH8eTJTVZg0WdFKOvnd+WZ1aLxVkTqrvarnR2w/MPdRXbIJ6LAMOU2hJxAO3EhAVG1Yq
smPBtIuDvPdod2OTPTh++q8UNp41BqP6KQs9QxAeNP36FA2GMqJJa8JRtv1MZjnD78sg+lRKZBCr
1ZhopE0tmOUF6LguGjGv30wlnAx+dmU1ld8fpqzSh7zVAfebuDot/1qGfRfC4ymiHbih0LPxL4UZ
bTTI48iXRf+llrgWSge8tjRZaCguOIXBW5Q8D7wSAWNmRFCwsROQ8yZZDB+fXb0tOSGV6FVyMbzM
srSsuf2lAiJFw8DLcJMuEiFQX2CkT0HZGr33KKbmmk+sJrNlFw8bchhfAnleCVX75/EJMziRc+gf
KsqLCFaElztf5+1hU1K+9YhkOcme/Y/UK4HruUJTPgg4u+th1mtStKrP1RstbYw1Y4IUEudP47Dq
WUh1LDJL7S7kgkZc8p+XV5Sii+sz/6Gc7jGSXuCvfnNLlQL3ufS144dvnOgWnfbI1xXAbUAuIsdZ
W4jn4H+hSXX+q5EImnle1NB9HAmzFWFR6dTBe+EnfMkk2pTFdGCJh3kN5ITk+lBkzHELaCTLfgWJ
oJlBo+LsYmOcMibVicMxRwJWTCJwyTFymqmweLMnvuT6E7eUYEUYDWoDpkMoyMDrcLAXNHpGgxdz
JoQigTewWcC3phwPGljFx2/7hnBZSpNotDYaWGHzr3BEOXL+SvxY2z4Xh/07QCUWYwS9hUI3aCcm
VwRtTMmYdbOIFzn3Ns/m2/L6qGmO8VMxW5T181xc/mMnC57D68yqqu577utpkPGr9ohGAaHiSP95
Dy+rg4xVvqnCfsgXRHduM6TGseqUZO0iKrthQD69lwtcBMkmr4Jm2ogh8qEN5J6pCfzxfUgZK3CK
Hge0aAWrpaEAj+4eWwQxB10q+umTu0pen4cFOjs+G6CTNNudf+2m+u3o5E/1DipjxruJMuNCy9d2
Ezmw54O3/qbKWkSJ6N5XK+c6BIZhzX6SjwUGIe0C9V2BEOwbTh7kZW2TavuigWWAt3gKTmLOnn3u
oaNmfNH26h3IQxfRayomlqpxaMEtKuI5qAql7B/273Kg6bNvvkd1cgb77WnqaL0IYPWwcHzNs+P8
Qx2nPEYCESG8ruVx/h3aFS9UQElrJ1Zn/OEFltQJ/IxsCtMj42xLZUhJcA5z9b6shyYDqkbuYMSq
1k4Bu5rXaIge7JvAyT3fS5Wv/JtMA9kjWGVSS2eTSgYrRUxO28O1L8z3Pwnucj0V7JwYSp217JJv
3rmgAFt9xjmft70QZTERjaRYFcuWCtYXjtCkUx0bjEPx+l+DYC3ztU5ZppAAqeXcnjs2iir9Bng1
IsDT1ZWrGtZxGRofIbQY333gVfuvMR1eAiwhm+jH0REO0hVXwHS+bofjRHiTQ9Q6HjuH2xi3gtmo
E3oYaup3Rv5BRwYnSMrfcdcMRitM3tibqUad0EDSLpR3wQQn8itNZ0/rLS4QG7S6eQUnzJ3ZC1iX
9334uCDLIhxmUc971hSNOTcfNuCcF0i+0olMrjUydl2Uj8akSAYsSseY3AWL8nHL4kI44sic27I7
c6F/G7+71qr+JHKtKL37cmL6iR7NqjfTusgc1mdGNtcKggNZJMplHW6XlHczpXcufBM05CWxTCtN
jBhY53+iWC33mlTVpQEZGNCnAKvDXyo4iBpl88oyGXuvOmkNiQwS1ZtRI3nzSFtd3O6MqRP030+1
QgcqlbLd9UYndqT2fQfADe0K01KM0XcVnZcQb3W9ik5L5gKuMmY+sXBNCs8yNCGLtRvvkRS/rEoC
JkcMLXFSIVBqoO0XtoArAPU2ksw4A9TuIaN0hBVr9jXdQyjBCie6Kn5/FsdvBqWVMSyXHNpVebqv
fYdV3Fiy4XKuoR84EOLM4AZfxpCYxlzBrfnbXUEtI7DqLKEi5Yf0+WfaSU/KDmDJ47N+Uw3jYpFN
D5Z2oTlC8GF/KqQvL8wND2OqLns0NDk2o/m58iWC/1LMYCTfdZjvItd0EZohtAvTrn/2Ic4hKZpW
DWCaQhl+0gWSHcuugBDaK7YT19M8tzD1eVoUOAr0KTGGOW9ud1wWz+v+leyd1DRNdmI6hsMTUPzx
E/b7HZxGzRd8on+ZsPy9TNgFlqTcEKX2J9SD97ZNQnVTaJy8a29a2UYTjo109+bm+4sP5VKxsB1x
9queigDZcc9A0l6gnRIqgNM0IIrEd0btLElc52UwiOXSX6zcE9WCJcmLBwt/U/LnLy6gyDjy1O+t
TD0THaS0Iok1DuNpz6RfZsTu954s0GMhJY4qn7ROERaKTly6ypwsq4P9eE73X/jHapac4Sx9n6Hl
7MXyFZoOL3RUmqEzZUgVC5yMbHnRLeweYRyHsgxo1b01hQlaL08JWs05nVXin103l9qmtsbbSEJ6
D3b3bVWN4TPDBAF4S8NC7Df3eKIruInj2S9U01v9n6ySGkZrNRz5n4QNmp82PXSA1Z+Hd4fFjOFj
PGVy502GQq+G1bCKmYGxpaJeGl0ri7uAzI2r0ciWeF/R2Eko5qDS0DJo3p9HnSl08c1Q8JCKnVpv
c+hIKLDWx4xq/5TQDFYAdhoAp0pkWZ0gFQX0qtCdZTuZOUXZeNd7sdVhtmWOef1msveb4VrV2J6/
X8qjCcbcuvtAaMXGtvBpo1GyoAxAUxVj7j0LsFVhuZJOcYtI0BVsWmo8kiB0LLshiIdzYe5UoiF6
hQVLQ045QI/ZMHSrk5tpfWjR1t2deBpD7yY4alSA9y0Xr1izA7Xe6LSVZudnSyGDRvlDvUEMY8Y2
XaobUaWBLuWKc0ZQASJ9oJjO7QiIwUEZZr/W08cqExoenC+uTBiTEsczbsb9Ar3RPpVNgxNeqCxn
1ZV4kzYAZJn5iDc8obiV/NYujyDkedzLlPaaJce0HHywdcLDLO2ZuGDzRAEm02FO9C8Di6jWj+qq
hOqUvc8LqtDpotb6spnSKZ3TKIFwLEiRdRz9Ydum7gzUuKX9ikUyq/7hvr/C2CBgiFDRwWreavyb
pj3KUV4NeUA4KRjl2Ict4xflngxgWjUqZgsX+8d4rkcQiYbf5fvPEnQNzjOHhtU6W9c0xJqmpJyH
oqHfOyU6DUCH/l21pmaONrp71eEd4qJvQ7FM/r0fgO9kzbiRTJrsBlcQAazI/3azu8noe2g+DCWH
CyKHoyChhqmpWFpN1R4P2ZvBsGmm7g82c79AOY6yPF8HNMhQO7laYCVIanK4cdrERzZByVOk9HKl
3eS82Y1LKloRAqni5ZhDD/gn/NUqRsxuHdPbLvDs4Y5G47te6TvYsF3M17LOx2pCRbeedCMnqeee
TFMqMuKpTvk+8Z4anvEWWzb4ASIRj4eX+tO1XkBmIv0kjKZc2GSLYBybzB5ylAslrExEuJMBHLOg
ddbvKjk4ys2JGzrrr5Gdy0Ocgrwn2ZP58BFg26kRJF6ZbIvhJ6zLjYPA2DZKPp3it/avMibHK1/L
O4w1MqTJcvr604UuSsvEtPyE1UO9LQ7oXMNu/n9Ti6NAf2SEeQjKa2mg+BvEx4nEJGQR9WIRnYYO
B7a1j0lHnMgZbpOyy4hay6S5cuTozj4BSZaaMxtlBBy9ygrTyuf/6Mlxkauwn0Wg7P06ETs9oUKo
iMMocnAfDqVpwc2hgYc6iIeaE9IsJJWyk8OmDrKxTtv80cU7PI/i+boHnhvHl9JnUcUXkM3yGZMj
KgYTtRvK4LfMDnDrca8RLKSifa1B0vFuuw/qrCWsLEzmE5LmuDiziL+IcAtNiyyp5Fe5+QateGdF
9afxof98kkFsndWurxE+nGDZaOrERmmch4T8SxFFyk/59xrXUVgRFkuFvJa8YTOl0c4IgVQG7KDn
LD90E06Jawa20TnAQ81KNqQFlLx6l8qacAKENkKaRsvT0OnEXNICiaoHxuo2yXutd71MXQlXk60s
t9MrrTu0b+cnxV9N4kSsm/2SfFvcOZjCZ5SVrEEFjo2hPwDPozkf5qvmbiZgLAzvkqOaJepEF9yJ
rFToCLquZHp6I8k0b9slUlh5Z3ZixfOB0SXKrgMKUlJmb/9n5KczS25hBXo82OHxBvxvqPXg5Zzq
/mKvspOsajwua7uYEYZ5hgujo1GCyjALir9MmwRH53a3yDi5il3fWdT8H3N2ksHVgNK+XEqMjB2i
oL9jV+Mg5JrFpipUBCSt2ImVdTnVCXVUzk2KIq1MB57OsZTCYswcnuFZaJYXVu2s6mOPk6Hl4OAH
mvRfw1eIRW1CaSOb8rborRfZCzZBnkuJX9TMcAYv4w4eB9YYsmSfrPE48UQoCyEU21VOm2hP9rAw
BKaWE4gZmvkfrhwtAM/zGoGbcmt8nr6tRNakUUMo5UYb7eOn3Z6xpyCfTtbP5XKVc33+Z6as1IJt
PHtd7rvhIqvj4LzNHJDPjLrenKKJu7qPVogxI/uk9TBmZRKrrIQkNSb9a+u9vxJ8vku93jxU77Iq
CMjij9F5naqaN4Ni+rasrWG2K/JJ7CHk8b5FRzLlWFTYLaKu9FhgfAWLehbKN8ZwNvZ0WmadjCTR
+SJu97v4rjo3+nUitmAUi+nQzdhNsJiTjrKbWy4giLXg1dEbB3Q91W/QXYJp/J9mL2bGUfJ5r2Pd
Hs2011A6FN+Me8sfYh7TS81OR/pyLunFlUoskRDuNQ4RchO1QmMZJKtUwKFbS04B4jbTqHmtboWl
4Lpop2kLdjbTI/Vyn00Ruo3Cfq9EQTwwtWUCvPKZuVMNpLbL3/zkqOnke4XM7XMnMUYu8bceMaMG
jeZKeaVcWjKd4Ymzjhi1c/nPOScdSWvB3PhUjRepxDGtq3PHUweX7qTEa1yEoFnY9CYpWRBNarX5
58HdgL1koQN9jF+bG52LTPUEQ9aLLHAih263CJ5iDdiYdZBft+leNWQUBi2tGiH8rKaB+4+v77O7
mz5erKejW1F/2Gy/UL4iVVZlzjyjOBSjw6aKa/ajuXkUsXOFezjmuFaUqPBwx01YwnomT4GfSOf4
v1oGADcGru1xRSSuEpl3YLlPDCTmPGdPT9SQNHcC/7UKC9cfzSSxAgyDqqVTvJamHcib3qvTO5C4
9/VQ5mRcPnEOaGCjpoukPzcz6JpMafXyJe23c7DvGqIOulZ1zdKif7Fj4JP0x6XqAkw8X5V2YLTI
7ImWdiilGPYvL4D5yekSSoASh1KXJxTIIczsp0PmLUjkdSaKnVguJoAyckmzXckcmuNuYht8QcUE
R1nEcMAOhJEISDWg+jt1ECrSLPFTw5fVP2X3TXQhlBxM7Eka7dU3HEF250PFNYIWycl+5HQ/DQLW
Sq6BPZTbMX9+2IwlhAQf5QtYzIBcJ/ejh2cjon/xBl85ePaxd3qTaXzr+Ek+qEGdh+431SSsY0tM
eYILSZYQH8zrHyPofJBCK5cleLlxrhveVCFyn4cH585k4ZKbQtFQRBCt2LPOYqJVv3iGP6DiTcaB
KHGiSu2jWQqa2FGGUfpY+te+ridZKr5b66qkMMtuXC/7g2w66a0nHiW/2KV1DPpF2NhitR4+BOyF
fyE8Nmd/gBLFiu9buUFLB6SqWRjPvp0OZW9/qhkUBoh/jn8LM2Uk4rTC8l50/mpr+pMH9Bclrp5I
THiTmStZwlC4VIX4eHljw2p5slAsvUfylVXMWQu7GFhoIU6yRp91hVj6xjKgGGcQ3Zh9M3MCxjHw
oaDIXTTmvFVgxgzC1luziF4OPDCGUEDbSOyklqJzGIt76nbHrb7Hn8/1JS8aylVHikYzB2EbEkhA
89mJ3AicBe/LHgp+ZRgVxAS193wiTPveiLQTf8VEDy69PQyY/gzRmte2/TQeSNsoE4I9rUJEPDGR
UC83SSfzTwlDsytHNIxqWpPtaTGadL85dE/xotWfEI9aA9EQJGXupPXbLhIhruyNbDlGugGMzXHT
6qLtvB/9vHP/rBzh7PGb10/qZIw0JNtE632boOrjWmUDr1Z7KCDMjXsBtf0ILFl92B4ROGNf917n
H6Emni4s7+maSNFg67rQPBKSPW01lInpWmhLrErTOwAr4Pvgn815IYCBn4wtvu/KKb3PNHjYUmxj
FIOhv6HltWkZNDJmCtgQ069kycziQTfDTe89wWRzCaDzHqqgSrXY5/zfux16E8YKsVYso3i4qpZD
bp5rMW0tvQ3YdFukjkCqbn9fCsmYdog6vn3HNN/gMeajEauDZ0QSH6YyPDZk9MPYJDTV0vW9Oq4A
sIkQ275iWuHZAGMo7TovJ5bVoAFq1sAVPKOQy9u/eklVgAjPWCCd6ZzakdfYtpJmVN2Rq+pApdfE
XUylP1HllBIjdGqB4WLpfltkcxY756bQ9ZQi5rGDR8+hPOLUIdzVOb1kRv9EkiEBOPlVvAq4Ctg+
x3F+7V84UFuursGM22uSRNUIzleTx46YK44IGpXd5mKmMlcLQG7liG5kxGmyXmlEhZXhcfxyJIf8
XTqXxsrst1SrrPlYp4mnVYTFxiDy9f7QjZ8mOzbSdj5/J072GN8BHs6io+xaGTFlcAgYt3gPThYg
3hoT0IyY5lEcZihKNhqMKNGW4JOO/tQrehFwZS/A5yKaWmipz5rVZjYE7wW8uAi41QFdAc/lrwma
n/JQ4XoC7o1+SpIViubhdp600J+pKgty4Ei3RSs5/wNJCe1zV176FRgZ8ZYxP84q6hhCqFDcDE0a
sYyB6d1kXIKWrCY+6bKBzeKX3RUG8Jx6ZmTmxMzSZEWbR4MNOqtEJ5BN8v7LDdPnklf71qOg48de
nW3fzkV8B5mffaG9GbptVV1SsoZm9wqiV3OIIf4Rgqwnoxvj5UcW2s7qnspIFY/fPRBOPBFXdJGf
fvstR8hjn2ernrpBIM/s3280rHYrq0x25BmD0w9PIVRO8RTcxWT8BgYiQ2U8w07ZX4XR7P0fnIfq
oowrZREAvw95UoKEBCEw2/+A9ixa47an2bjlxAwXDSsF/phjj3T1JychVDUNaV5y2MIAt8OCd7QX
ayLv6MSl5orUm7/42SXh7NLX8kjYF5qnZFa1I1zY7IYMVe5cjfcvlHuZLQGNPZ2cZwZfeD2SFp7c
hNgc6t8fQSfQYjv0AUAlfkNqGldab7emmR4/ZZA6ngGZlvzTb5iXDE+ypNXpHk2vzc3eZFvuaPn8
bqKF/m6qL7jtQbHR8P7AE+3Wk+KW56ecP2nQwffdcSRa75AV6m1SnAN/tDuHs5Ahiih+Ya9IdWbH
s8DUd2LxNToAEK0VjFhYjc6iHLFALlzO67K+WFTUj7XzptXZwqEN1wM6F5uk7/nAEdThQC2rpJvW
9WwbakkrctuODB4OMj1Qp5Gs8db+WN8gA/tzf70UQeh4NHoaJAUjkB9JRrJO9UNgxg7bOQ/2rpUj
YWiXz6VEJDAUu+QWrbiqyP997OpFomdWYspHUqIlHYOESyvpyfksAYbEBeruv/tDqx4ESO9Ha8kk
b317wZuCUVmyANlXVq5l35zjjZ4qKxt2x9w1ipr7m7i/TbkrMU+z7qc6N0XH8ryAllXJ77lJMLeW
DdkakfXD5nfJUGymbfYua5w+B1+pBRa4KGdi2KwNFTdeNrzIy6XReTg+pnENFPRIQCmyvZ1xyawG
FrRGPxMnCIqZVR9aK3XLU4bbZLNGrGqxbwD+gKxOn7huPm7DhoCb4OjaIZjFEf9qAn4K6OloFGiD
AL39c3cjUKRoSXkGyvD4oE4eg6GfxNJeI64nvdPrErU8esH2Jy1UEGWuJSwVCqcEIiQXYx7DPyqi
eJnzllO7FcCQ65Jvt7x4KCEbP1uklHG8e3k06xhCdTgdQlGUi/Gh9l9Wwp1nVE+F9VW4OCiGRKtQ
reELVuM/0rZDcyCFhIHSx51W/Wy2VJms7tVQIXoF6aB0s4qwf9BI2Q25JiiX9WMH9zTzk2qZmhYA
PRgH4GqrnFMfvQdl/DgxbE1el46qU19UsZaxwLe4edJ3mBKKaVHcxmFJnnJ1bI9GrIrzlZs8hg6r
i/0L/m1L5b5TGukvnXgcKGuZil5fAAjMjRf8eQi/1lkwQsgGMlhQ8sPWrGg1xwa41SUKXfyAnx+T
mjCpDEcEzox5mhspYJPQ1pO/OUIXt/va+JLsVDt7jCxLhU/IgZqpQoH5t+oOon3nWtDtN2KFfKvS
O5gAV0Fsk+y/uzrfnMl2bCpPTP1ryPtIoR26KMhkQ5v2CYa4m5rn+XT+kAJm1bIpDerv9i64GnH6
r3wMs74Y4M+LIDBGc95XOU8JaFo8NdAFBIPZRBoieiuD6ZG6X+bcMjmUps2RoaOWSTjx0RrhwGQQ
pYfyX/iohfyVq4ER12ZaWM+mwj+5u/HGWJKEr8GwIjR8HVNgLtx6i9IRUYmfeU5j3Bh2EBj1Emel
YtnMy7EMofnTfXGI8nCkUpTAs0H0+jLTlI/vI17JPEuFJ9IzBh7R67BFA4NazsE06hZyQt0/Mu3i
wmUt/rO7EnEEUZ5zcsU/Du1TJazJN+eLgUmvWImZ3tGpt2Yh9jyWuRexQ//0jiRqKax0UInn4m7H
ew1lfW4yhLaDT9fgoWPGWOuQT6SMK0UH4TVSrh6CSyMyaiD65JtKOzdP3F1WCuZat0ynGz1KZ9h4
pK2oVTwioAEYlicGc4lGl60p7cpM4chLIZwR7XNakCjCwqXiTc80VayoEZ7fekzFcCWIU5/dOeVp
oo4slHtmMwFHaMv/zOG947fYdXDc+XlyMu3bhFVNOqzs4b8gAh3nAGOpc+smQaIh4Jg+6diR6ie/
iwkwNuVqM7mdkoFw4KyJaYMlXCusihSHvdgnRG10fcsAMzW9fOpHDuKeWtbpjm/zSSdIfhyWs405
jctWMh7GZ50nSYBjrFKkwHXvj9ifhxEiP+nKro+F7ni2HHnKIOPozVOWADbU3imogAeMmMVOh6FP
OyYmsvgEHNCbcaZoPjrmZMl+/2GpKalPaMzo2wmmFOahF51uLBfotCX4ElHwwGPihtILY5RINiaf
jUh74NleNHPNoR2hvFIG9Q4Ei8+WOqXHqcPkvv8SJXo6MQaTtm600poGwi8qiCim+LnmjRIXVhkM
XQlQJYrtGt1Srs3F4eud56zzr++1rhVoj4YtPsi5m1zHQuIuAOs08VQDchcvyD8rr3OjCwXxg9zA
CK/FhyL+Ja2LIPvtheo+DfxxGrNeci4d5Loh7A8ErqEokz/xUnD1cSVbaDzE0Q7ChCDWGWKigsCz
qhDQikbJdxam3EygqCCWhpLgTSkLCa8Eoyw6STkDIWQrLu1R0iX790QbXahhiYAqm9R8mCe6gdos
PmUdG5nvpZ7XGJE712PtXpwGtywk3g8t4Hoxj8atkNWOtEdZzQv6LXYAc6IoCgy5UtOAkVvW+Yt7
kKL45R1cb8x3UmKkl9hkhLNANobWlUzOCzKWOgWiavLIJLye76cNKEuJfHP+ZrN0UXAU2rrP9a/8
ajAMiNgdaCR0F+KijmubYxUB1o5e0TWTBRLz5g6wCiraEPIUfoDwODcN1YgeRnyd6lyOcM4oS4B7
GC4jnTaxIYHKwOPT6dTwv/DQc8gdxOs1nOJhf/+OU9T/hvpsMNkCqCtj1H7KzaMkcfbfMwfzqpCx
uFknrWjvSBb//16836huJebvaq2NpAqKoXPP9nCG79xkLbtA8I3BlgQRnxi8ODWs4aWDT5GvYao8
WhrKPvJ4If9Au5FDfwDqo2CK+WmlXspbfZScsaXTbdriX2cC6i+nEqyfhaOGwgcvQEHwAoE+7FqY
PcVUNP5GA74hcCSOCCwD59il/dcuxP8bs7k1jxMcVkksVuFL6lTnyBawKANyQq3q3ffJULOJd44/
i9LCai+dWl9eaZsDjjswTv5plrDxvDZ2lQJmialobiu8s9B5tPfUflaJhfU1eVm6WFJFm4jOhv+c
Zx75l19RiLzAXemREcObVrcRAjjwvKOsvCvCyJAqNUDTZG1SsXCdAZ0+up4E+TskvH7GOsRFb2SA
HZzR3baGJ1bp2zkx86uLFMGmYRLSatjqv7D6rDA8uObM5q3+U99bnypELPviNKcCU1g6h4SsycLv
2AHrvt1ROhpPa7zinre4yja5OlMqR9pqpiTBFLgie8gz5g3NzAlFBn7g27AI9zhaSBAhqIQMoiGt
RPsN6sq9kAEqNmyiJTW9G8JQcXOnO0Mv9657rKFiJHfRVLP8FovDCyCo7okTyDDmQyy/W0D1G3ey
XIUnZtol2obPHk72UvW2WeR7KXRWuNhuwzMe8t/jYa4AF2SEcJPl6dIxhsiCIHYdKQxcyTSxFdE2
RFkvF6Bt942HwSjNd6PJA3X9wMoTLCuY0nS6WlaV/Eg30WqJVvWQGhmyiH8sNDcNi7yJHKNMmoLc
SrxoTk5JknLIG5X26rvZOTxHAOBIFDg8tW0Co8zFpuqX8bXQHNMHy15WbIoN1JBWkKrdTnsAnGA4
uJlVkOYq0UTHccCUfX8zRXTgGzERpgp03yfYoFOYgOZFdV5pgUY9x5CqMEg4OY1RUSsBqccRhB/b
Kk5lcXykRDfRVrAlWimwRzkLBTcLLLuOEBRAdegonF39c2bRN4wkn37X5E7g0O4IjLP5YQF9pEbH
GwuqMracYT+iN/i9Jfowa3LJgow0cPi20b6d8ggk7YcHPce27QWqhKaPmw3Evz0GbtNEHX3HO9Md
ZAdeMNZADmc+8YHmDrfZOLp1Nu+MWzkl5NRW99naj7oaZNxGYYyYcDLVT2Kf/p6vBZYO4FmXWkvO
t00++6VazJvlbPq6Y6RfWbRHrJdkFxpM1tIXhHcpRth+xEw7mVPn5CXehbk6pUeA58wfvOwuEMhj
d1RO+PZCXE9UnCHH8MQV05aW9zZq4YROFkpHdJDyP3CyjksIaUFWR6gLBQjQJz8PNM+FNtL1x2Qy
sp4nRVHtYToRKY8cKPwdGHhXz8HfNCwGQzJw/TDeyiKLE6ksKW2RhT120KgVJb3pelTCjbaDcGom
Icy38WOJRogTZ41hz3M0OulKsGRVIFBo3vD70Qunv3+M1Bb56Gy86kKjIvhDrO2wn5FC3SyIUx5k
Xm72OgNkBfYNoESdMFRettm03C7mUCJb4mA89ilBZ6JgciHL1UNFbox5/KcZOc/zUdPsupYE6JKj
IIddnffoqZeytaGkhERgSoOoyIQko9VngS4cHeRHaO3vHU5G5K+2taDNnLOJ4GzUVWy2eTGnbiwK
J7C4I9qYQTucOJI/yXF78khOY5+kYQPsiwXJg6ApxmyZP3xwpYk5HLEPF7I4sYwK1twN27QDAxZc
zjKujxnfB5sn0cpplKMTREKmY3Lt73vHo7f2riaJv30AzN6gTh6RULHta7ViDHa64g91DlrcFUBh
e9Y+M0MjdlucOVhAPu+++D4nSlqTs+zhpNiq1rZpdnnTfDv7B9tLd566xr+gBlS6VwrpdXh73hkO
AuC6e4e0LJuRHRZhzKY0p64CN+W6nKP3ijZzWf+yb+fA366W+MA2KmBU5d7y1RuMpM4a7h62qUTt
VTMIkImiCHU2uraEKGv000ESF+qukLqOR9Gv78an/XuAEechjTGxuNTkwzXBOeWC/22e5T/hJF2/
O5HjV0Te+lJryOpvAaV46IYKy+E3FIB/wRNMm1u0DoWrhbfHuOPCWv8au+ZnvxejZHSM8fuzle9E
u4zPPgJiBCZ44CbT+NhrWp6fB4kEa6fvpFHQTx3n3QbYwl50DexwQQ8OzlmHsyfvmYf4Y1D2XjUL
8BCn2EdVZFqkxjy+rzDfHeehul4kJr+7a3h+0Y5I2C5RJMRXY+M/hlUPzCveQd58ZMuNuvYOR28f
DJPFgyD8HaQwckyZSl0Mu2vyqy7X/70VPQ0lgnneFX6r0u5LmyJ85z9Ty8wDiICUEsAlWsOT1JJ/
XySDhrqErUR+fsn7GTbw3kO1BlYt83JGt4YfS0q573oXyuW2sfh3Iz34s1UAXl1ElUt572m8kMoR
gP8SnEnnEzMuGI4Du0aGhANBy20cb2jFpp7/nezeSKwBcoR1rM/sH5b1Zxiz9YJndpe6ccas0EaR
GQkMeQ0c/Csd3IOSh9ecHJMR1wYMy89CusK7rhrqccaq/cesVMBCqTanPFweumg6/bsBNRrcSL1l
ooVjxALdkg9x9uXtxMHPNHaiiw6ZC3hnkpBKHy24A47O1mUz63I7cubrrLNc+I14F8GuJqXEXvcv
ON2d8FdJqVjQwMZqIe09uh5mWzjZ8loY57PgVhSy79bsDT/TDd/B39wbzp7XfyW+0AbNiW45VMQw
aukUQRJXxrFPRzmN3peEblI+iaG2BzpmATjYIFUjwfrYmHV44EY3nDPbrJZtbND3rkBZmpJNCKmA
een2jbpTybgTETaVPMIpdCahLlubWkUluH8/IqXs5tHSurQne3+ehmZr1dMnBXwFm35z55OD+/iS
kPR14HpSLy+xMbMb5mGK4GemV0H/uCmfpz7do5oaPkfW+2LSAGTCi+49SCohjAAX4Ed7K2YbFLDp
jinbKJypfWumeIx0mwcx9uKJEVdPOfISBaMQO6OX/Y3gno2q9CeHzRBjucdxiuNtY0zjOW+BKBLn
3MZhWug5aZoenGIXPYff22jaCxj9YdMrItPKtw+0ZJV/5bQcAMT4sglVFUhZWxoj0fa2a5mDQc7j
4cuTbnztLKGuXyGT0Kowoa33FRk/4Qkk9cWy3hbazCxLVlTxrHJmyhttbhE67VpKT5hWDefCuNoo
T+RP/NXD5Z50DKW9OKIeW/EQmczD4vgOVVAu+R5G7kt47I7tTlK+it6EO+NvKUC/nd39r3vRpC2R
YeBKMyTzeolgRshjQWh0hK+5hRgdjt1AIuqCqjMuiBrd0xyyXztZ023pmtUZHur39UT4M6YRuNfd
BUgSUx8al4S6CrTFXGkodBZDEKjKG8y77eNmBe4Rtyo6Od5ElYr3N3rlnyOu+YQSePBJkjkNEx8A
mYKo0v4PynEsal8bMocII/V572tSChPVgbV0CcD54EHTpbfOiLC1Z6rz6RUCuxDtuKeKSTpSzZD/
JRsrwguC8Ke0J7DqqIT5SteC2N/BdVck1G85v4DFEuCZAJ+enQuWNNAxG3FQBnCJAFika8NPH2FS
U7LUpCCghXJ6Y3yKKx80Ax96trcOuwBMReVuVeJ4a1Nl9VGK4E23URmPTyGqCuNf23X0BjL3BI0y
vSK14VR5tJaiychcjOHI8RVm33ABzredcnr7vgY0lUGOz3JuyjDiSUBnqHU4od6WR6YXXoUAXv3U
OBnpWyFQB59vCXq2IiT5gbUSW5N3UqWVqaF9wXRO5F9X3J4UJblgNfmiwDpuSE42kc92ngnoF9M/
C7KWvZTcOu3RVq7C2WKrVcS972RRF6O3lR6hRIPOaFbPRsrSeIVqMnod3hNra9sI85ZhJV9BY3OC
BZzu61Sy//WXJPOCJBOJSBBIiFVkLCEStRtEjw65iNLQ439PAbxSuFjILI/3yvtSEfz9OUlZqwtI
8TH8WDAR0TnzoFynBpNQ98D4o39FSl05py6/u/mgjRVyoZkINgLxPqyd/sP5JrCegNNLSc/nhEnc
jdYtez2PRrs6WOFf0l6PyUUFhQrTDWRei2j4uufPpyWy1NHV584gjOp2DXtu9uH6O3OS9UTlOSuJ
dYP0XVJ7D8eIF0uGVRk0l1Pd7PQvRcAdjNx/jSpT5cvkZtsXwDTXrvHYSFyaKT1bBsbTuIWpeb0F
si17mUBHkGkrew0aQJVB8lFLOEXDDUAVIqbIJ273wQn6OS+PQnUiTSEVU9FMwXR9eiUGu2mVyD9S
+DT591Sr1BEqXwvAsQCsdsFco8iDuYEfxdiNmUJ3I6T2DFaEP36Lewhw8a7zzXpDa3YeF1uu0glo
HHpAiTfxaAAWDS9m+9g1dHOqASYLbtYOjMj63+Ll/jVePVfwD8/JY2be6B4UfgLjwHqQT92mjzcf
Jf+Y5yZkx7uMsms0RRqZe1g+dMVcAUhUAh5cMs9rxmlBidCYTQshnUXA/iLWinmzRGhekkFyvTWA
7eGHSOkvP5jz0jazZSz1ZmCMswfc8TmeUTeZrCnP2WKchLWdsKSjMEsUnW8CE9D4DjVWIQIJ6KF8
OQPY+PLsjkfwjaFaoRkGJqWwtN+XxzROqPXOvsZN44XSeyJIpHJ6N1UZD/Pz557gSWFTjTDg+jAw
3hzHsOAjBsRCR6eVNH/tt2Z7nyf8a0ZttD9/lDLwsEPspnbhVGiLjATYPew8BwPcNid5z2fQ5YQh
MhSjoB7LA02i8QEi7WyAKjiY9fN4Cv+Pt4QEv40JZlcctINuGK+ZyX/O5Tokv4ZqX5K1Vod1rgB7
RyzCMkZ3BFJ7hC5OpSVB4qNXFDs6dRKGjBKHlXwLw/v/3iLGT7WqM9aSCSu88LivAzq6m1gHfByo
mWv1p2vNJ/aIydmvvXUB1pQzAVXnALN7mq6GhrV1o4A0jghm9jyy2XSalQLhxpemBIBP4oF/76tE
AJgUN+nQPCB6cVR3CcC67izG3SK3tr0LtUkcmIkdKMlnXRCPjpdl1R04C9dO66068nZwYfVDxHnl
MVXkN682hdDU8ydsMtk9JgrEpTIGPJQFf4Z04qH+4x78ZTHNxaRoXVJZlh/MAbEeutG0uTYvv/vY
nuhRQGO2wV69Kiuwn90X9IT478Oh4LYICIqmIwh8YKRwfiFz5kre8B6/n0Ohdetq73z7KsPmNC/L
yq3MNuSiNPqgwo4p3LFz4roVzuwfW8PYQS8pXhkx6aD0keZu3/TnVjjKGc0pnz/J5cw333RJdlYP
O8EliKAmORHGU7Ya2jfRK64cKu23Ccnyw67GYIlD+fgP/eWYr7XLE35c2usDG6y+BruaAsYITaNi
sbVas9enX64EMwjEpamAPtnQzGN8c/Pv5P1rQdZPt6R8XF0BFJshWOCM2pCY4hQiKzNNCgwy2wtF
9y4ZrJXCdgaNoMpdrtCREJLEdrx9bMdSkVXP265HmyXVN337Nq+uMk1y+WhUjYKRJ1LbjQMxaZ9O
6NDUSudQb5MfaAOQw/fSIi1aBTFfurRwsOkMQ2uwzQpEEaKMpVPbaR9wTvjv/VSg9EvxTtnSmsRB
rGwDf/Nhk92iMwHO7uppiLBBCG9YxmhIfp0L55hDw+k+FtnL9GAxkNnVsOR3DUWjemk/nkoTv7U4
H7kCp2TS8BJgd6Jn9u2iWIW1j6Krsc06bCqlZHbqPumckCzNovH9q4/Bvnx5Rh9uupT5+XZ5xBPP
UWjq3s9ITf5WYZieoendhoX93rllfyvnVMYgLRDI2TCoKVmz5rSpVHS7QtVZvUNULaR10zMncOCI
WXzVTEi73Y1kpBj/aBIZWCx/9WQmdH7RGMclkuxv0vzoN3Ae1W7h323WqkrBdPyomXr4ES+oDaR2
f+8+msygXUvJLi9ZGjCCHQoEHA7McZQGp0rU4tyA9OcRR1Pmok40Wcx+2mWK2YF/xp4R7c9Jw+Td
L8i59U/5BEVAlNPfrx2PtEb31ZGU23KIovd4XZ+wodVweaSPXqR8EniBy5rBAzh0+nTXhdcjc3fj
8jnp9yOBPDazHg550i/Sni1xjRFABjtcve5EFXDa4xiwuqPQqnyaDq1yQfEwRBEdM+cItXB+F3RF
ZS4JA52aIatOQbmcZy0Tt+fj/rDrBMJDUoWQfPWCDFjW8S5WUxogicGjn68pQTbHbozebWM7pxvV
y7exouZ5xyr6hIgEaTDXQgOPY/1nBwheXiQoYZ3GIkysjpLxa81RA22Fg7vxejg8EApNbPfX7SF2
qaQJzQ483B63ItiEl52eG/nXoic8VEb4ax9066EXntIxmn2E3jbMS4oRlQ0XD9CGIZ3ifo+FwU27
BwCT42+xAT9MeznqbjnokKElAZwQFdUxMYk9HskSjKHEpv4189TuDoAye9FJi3gO2BkSpAHH3I0S
azm3uj0WWpaZXAZ5B1Lk5oCNQQMrSW9kQP6ETMdkudnGMGKgUQ0gF2PUn68m3TTaev+pBnHJUcDi
J/PSBSYdHGUlciEXHh+OuvXiBJP9TSVzKuDe0PPb6ZcfxDlku1HZn5SytXzgBKxKooNFLPzR9+zf
fFlwtXBWpykQyF/XG8ALdYH58trAxHmkL9GnktFCYVyTm7rbqbUiNokoDAdRxZMZaXw/VE3kjeOJ
ubmj3LRvfLXvp25ZPepNl3G1DGFTHU8eVaAzWELsr8qkszxhJb4IPgPjgnpNHEIL4sH/8+PQKxxC
eVNx58A19pPZE76h4EeVYXSTwobllkDkV5zrMf2MyDLA2fDVMoKVigmjXM3CHqxk5UHAzw/Suv8G
2vaYVg20UXVFfQOxyUmdOnhqdTT7QF+1FY0D84NnnNQxQjbCqs+ualR3hzuK0r1WnTCSsIgRVKWM
7NHdd3hVBlNltTzIex7hddJv6f+o3biEvigaXi23o1Q9kMmoM9cEFJFYwXy5NN0OGrbU7dVAxgbj
PQin46P2Yj4zolwar8NEGYwxiU92auQ+EATanniO0qp3E0mO6IOlyrP9qbk4YsKaoCSGm73fHP7G
p2zcEyanVieNMy8OW9CRCbzh7ofYntgj+hUYC6Xa3AGbzMPB6rF9GcLwFa66kUHoo4UWLhLGKlZp
/PM5XQQ7qowHmRRdC+Gu9Vx1caBCpU518+Cu+SLqkJwwK6EuLBupKEcAxlm+P32/Q1rJL0D2itHs
Xqm6hMZ/jfYE55mxQ02QgQOhsCMJs4d0RI6ORBb4c16xO88SAyi6KassurOlbIxu4xqyWi4YoYs3
hVm8EP15Kf3iHfF2dCTyOLjHlNDN6dY5LVlJ9y7qci3pe7/bZIzXoco5m2D4Y7g9bR8ydlb6uCtp
uwT2vZh688TDG7GpRIRpD/ilY5cMKI6V4rqQm49x9SgoAFc9livsIrGrYuuadjsEriJ3Zw8oQtDZ
xcgYlbZ/bwbo4aCOWcM25ML1BW9TTGYW/yJHkhBkUw+4szLwpb1UNy4oo7ZkDAr1/jaK4nBYaw62
xHa8XeAtAZZpd5T1gTPDvycatzMiXxfBKryVV2r4EZD8nzZZJEbZyo7ErGc9IHaez42xLIyb1+RS
AiOyAdnDLgyyNSYrxx24K0FhC7rw7GbAgaiantaGqpFx7qwVFdDyYQSjEEG0rH3E1A5hUrjoKJY2
WGjXyYMHM+amFZBlcMwpALx6u4f3lKBjmzpgf4QfqNCMh/CktofsXREXRTBPn7WhzVARZA//aN+E
ahoJLQpL2tPdj7IWFWZvwN2c1K0y60+9AwNj+cD7oaCtqJQypY1XJtuG7N4pNLhjCyf6ah4NbmMK
pkZvab+mgIYBTy46c9//+moho64mRZyYXJFhbbH889yDaT/0ScHcjflsK6xKAWQXB6+OOY3bjZjx
pA2ZEETVHKht3FrL+GfiUcxXy2nW7wz9/pVJQTlGL+oVlSpGw5Q9FzcNeVZtZEiJl9Hi7soiibss
dahfKgkbSdViLXl9l0F4tXQLPpUTzPEQt64RPYtwfSH4vY1llkTbpy4f7iSU1n88RuzaaGCDcCb+
4AYBu6sZFST4G47IqhkBFWYuKvmQB0jdLgD/I/tYQpoLSuFNBXQEZskwaF9LhEiLz1Qh52cL5fZz
tTlbVTC2tRDnqaLO7u89V3HvMp4qiYdYTXBoDp/4h0ev2qAyTdHGD3qaeV0Qca14LfwlNrQN7VaZ
BlrwYtLIMysQW5VIXyY/Jc2bnZKeZr2KLREqCUjRL9b6ba6XgA3FoZ0aa3TKCDmFIIOxkQYE1dwj
JBBEG2/WkmmkjBTEhHaVylrxmmSyWd4hdsMVfhFW8jqMPtOCZ7nRAkFGbHZL8cIafJI7MmdJWXVJ
b6eGrTGQALHhClVEjczMYBHZAX0fyuxoKhyCLACw5HknegnzcDisPT+bbSpUY+N/4664dzt4FLy1
WUeJTKbUZjX3VLxfpx0/0dT+5xFDqCE8WTyrGTBOvI6H9jJcWu817li3ItkLPaDz8tYmsdAZtgWT
Va+jvurIBDCza7NT9gg5Qr2k6mdwIgqUMo1LL2/m6R5I3nMkwvMHvmgBAmuLERBcYWvUItbhYnMh
/HJUJD/6SLg0OZJZZfJgQ9Sv5fvv3fpm+EX3qY+36RWt6e24mRYQXBX6InHmsShY5rEJ0gDy4JOx
3EWiNxd/ZKwAjAXVt/jQW3f+LPT/bptT1v8SRloD4p833/UdfgmyyRr5ryBeZNzC5/k0QYUP54Kl
wLbcuzuHLkaSeNXFL+ngHDp/cUVu9ccqVBCcx8acAOZW3MS9uX1s+3yZ7YfZbR9BpxRmao8vF/2H
+++w38+HALfz7kp4lII2eTEY/aRkaBJF4Rhia3ajKcbjPr1tVYp2tPtCnthexeyAsbNuaJAizpun
+ufi5Pu3AAFdubuXegz9tHlhRlOR9jV5uupcrCMzdiHg53MwwwlSsJW+H6PFKz0x4m7wQXdXZENJ
NJXbnoL+UDUOHxP4tSpst0GOD3j1VYH5md+GhFnMFVRxNdI4hMO7ng6gKl0vDVAKTGt+hGhTm9vI
GktlQUzQPtjjPGtooawVM3pmDI0E4M7qbOmLC3AxpsPZQeqlqDL+orwkx1Zvy2LQsR54WALMHvgR
1+qvfPmdtL/vXJXdLfkkmu5GemcJnFHsbBstVZxJHULtIUeJFpg7+YrFcxAQSWv6KwH2uA6SMFZN
CCVrH+QV1mMUoO4idPA+G6H4hd2mn3aoeKZzastuX4pAvGl59PwaT4w6fIB4F9fnjNox9PXw7WTA
AzcjDeIff28xqpZgW7VW85H6GLge/8AxUrSaMs6PUoBsUpu9qc9rbrpK1lhT9+jlAE5WvROUIS7Z
OhJ3yIIzyJaxwUYwCED408uQ/GgJYifrV7rtjeiCZeOfu0PCSyXXg/NwdrUHe1E3GpmY3QCcvnQ9
zVj1JkKXid/kSStkiRnup/DsygyT+eDVNtCqVia9IpfNsy6lSFSgmRbEHd5QRMZ6kTcn/dttE1R8
HoasP76oURhEyJJmhopOQrfa3G5kuTsxwQDXTGvwBcOpGzaLUQwJip8jYxQfIBDtfCaSaSBvneSO
A4EZlV1dFtgb/2lpy+u3prl6Syd+cMh5n0txbtlUPev46pN+Z21uBTV4zJE71Srj6g6CTUVcU5F8
fI5eOwTr2YLCKkuOFVNXJsKWzvAyfqSluPkKnzjXrM0zY7VNlBZCrxxfi/sV3N8M7SQ7gaKp6SLF
DLb2lK1CCP7ydkRifNGkEcR39J2LIdUesvbFfPO9/iTxDsBMvGpuKUsOej5qWiw8rcYo8+vckI2D
VneV1NQxNZo/YhihHLBEguruFXYESklLIFUr+xuKafM7N/4RdFcWBBmejtWaD2bFmHxJU4ijH9sl
MF+WtwPEuJA66pan1yJa82kLTmEepucyP/BTD/X2AddbubtdktaxXFUm9gZxAruRCbiWhDX/gW/+
rm6TUN7urA4RV4mIozrZoFM3SCKDQU8w4aopcnWzSgSfAyqhM2GWdepPHgjPFRsnjN2u7BwjIChw
vy7AK8YAViC7Knd81+AwA/kZg3LKPplZhGHPt1h+R/0K+FCiMeOTRs0vV/wEKING+uYbPL2Nekst
/Z163YrQ3fnLVfCps4m8+yCxHd5yguzIq9dwBuBPgUnxehduksOtAdZcOY3b3R6CDTR7uSaTLn7F
bda64Ftzr/oXLFDaq8CKYKM3sB/5DMx4riO+qWX6ic3gpZBcBLZxoMnVef7dd8XzUzRzG3GrLC0Z
IC+53IcXLL6J8k31TUFfQmIHlBpyX4uSH+Eoc2Sk4aukjRVJW48UycxiHzRbjGBPCOLxOci5ztEE
CLGhM/BEqCzpfiCyUllF7E0K3DStQvAnAzUAoZ6Wq43japJ8U+hfBcwFDaDswdzWEpmCJkUcZvtH
TjNn35ECKzg8EVD0PCl+RUXeNFNkN7OHJDMpu99yduJdMEher5EwRwmragtpSrY0dPgJpPkUXTic
iAE5IH8vhNUcUL+TUmIu+Wo3/myQfyDW7UykbJVrID5sPTi6BGqTPZ+VoZZAWFFRsfQk4D0MBFvK
rRVaVh1ohGBQ4bYg/stQhEe/Qnhno+xFXsQAlctv9Jx8BagvGmiiozCnzvEcOlhfBJ3pYAs9krrm
16yPa3cI1/ko4MdTODul6Rcv7IxkQSiM1Q3ihSQWZ/aYisovZl9Kpy0E7vJnfDM1WlyundPVYrV/
DOcGyaSgnP7w+BudddnEUYiLCvOC9mnB9OEgJ9ScFOfDFMZpVWVb5t67D2h2LdJx2dDBOeoXAr9t
qJpuPdBEUZEfQzODuyQ5otUneYQYrHbAs0aQoqqeQTC8Od0ppD/ttQEWjIyvj51fWr4JvhBnm2/h
sx+lts/2a3zeYfoM5hRdU4I7pfg5RCS4GZPRLZO0yltlZDvPDu1nOxzn9dkg2JG9qToxY52Ub0iM
6HVmgJjwQkSJSUaaEkxNUbjt1S/uA8oXfvNQgQQ8ffg/ViAhocpHPh/x7VuWr8mkBTjyg5j2bCC1
+BPjsEls0eXW0PfgafYdVfSl+99YTUWUfFqEf7yHxwEH+UKmtI2SaRkizjvGjG5Qfm5g/Ti9s0r6
BCTuq5qmWXw+MRHDZy1WxBjREO3HqupiVQdogZR0DEueljmG3nrHr1wytvAS5XqX54HZpWg3mAbR
2fPhy5lsB2uwYsZMSJQlw+xzCxqugW4O6gQFUM18iV5wlR0cHOiDAPZcPlamD5FXxuYnxk7/K0J6
6TWJfCYDwCyR/DumJEb1fx6axKVWKumrWl3A7wzbfClvTH6z9XjylMOr0E8bNPANcqI74rlx8KB9
z7kKZH1LZ18/3pHH1hzxbTUyJRjH+Kziz1NGlfTvMDj9Cu7XTqDrYo/UOuF7Ss5n3jhA5TX1Ofc9
XWhMFb2wYP4WJHtgWpqJdgp0Ex5rErCXrDboBZo+EhAeMGmpApSm3RIcOuRKbV0Kq13k098SG9E0
n2fPF6kXFILgJ/8GOJP7e6g9UByriHgzlk7q3mnLhvNZ47YzR+C7/kOLMlcIzUcp18t7/LQz+xgQ
wQmTQchy5dkMPGgO9xb7W71m+OQq2Yz9qQaVEVZ+flf/h8sy22atd9oPLN58KIMjpAXUauo6SPTr
UY1nVMUGmF3JogxhXZsabZpV/VqpL1+2KGc6aFphqsiWUxQ8pXbQylSX1h2EdS/CqKXvpEmSPSgW
X/YFbKb8+SUd857XuxTRFBsE9UOvsU84qgP/MNkYKj4nkz0hF9Or/f+/Nx5v2u6OQaJOFgjU00sI
Rbtr7H4odcfAYUW+UDyDcOAcq0k/XCy0zkf1CS+co9vWWD1Jg7vudprvJk3HdONLDSwPSam2mwdy
3P5baeDMzirBO16WBErIocUDNmkvg3/T3rlMZZptu7mjHRzDl2OtC+mpYISVt+2SY7r+ws3tKSb/
rOwbQf5JX/RiK8O9+0CPAzITF7W6a1J+poXp8cEa6HnndHkQ5YfyyQdpPolw3G9R2OODsoMtUYsP
XmfUa6nxov5jTHpbG84C2upESBwGcd8fBpa2n72gGW6z9qb6mYYt8NOlf6+GhxV2iiZKwVT1hEYR
62WsnPMDmOnZh7RUAAdP6BXWOPzNhA/XjhPDsG2a71rSNniYrcqjTyd7PDHVNCOie+N/ZmiILOlD
HY75zVjHn3lmQE6Fk+wdQmhg5CP9HZ4xMn849w5Aaoqdm2b4r4QuhuWl2K8koX8LKFwyv7r0KHsH
9TUSO/uA/LzlVEFfV7+Mocd7JuXoOekMOOXjaKkZG9RKlm3JUuP18iJEzbZCoPba8Tp6s4RaDWjv
0UgOcFdwS8ZSXEt0c1BvfH/YCqT+vZt++3SJDyZjCgjfhvJEX/D1C787v4e3n7QMNAhfwaWnWVhC
XDpH2gD/z+VF/2LO2tQAmmy5X/Zpje4sR9/VO1nkc8lHaOiZ919GrT0qKufUp0l6oqIvSAJRkcpl
wq5ZXIjJJfB4/hAE0cawTgQ1aCDO7XtWnFA6+LaizZ7YY43e26L/MgyGfoMHN7uLGymL/fOXUswF
ztT83WUSUEoTtKYP1k316svNvG0nl7/RugfuMD19fVKQ6RQ5sP9nQwCWFQiC8W/Sv/at406DcFde
6UYDhsuKL9mfAETBpZQZpDE5B1wjfDJJFxP19I9Tmhe3LIl6iwC+2hxMGU//yIWwb7qqOJ+2kDy1
QPyQPh1bKuR+TQUXtQzcu6/5n0N53fCQ8m05txxjP/0z6Pi3dpzEhEjmfd5trZrff8VT6cky19Ba
xtjM4Pb9begjeS0FeKGnUSN1rlQZ8WVZxZHKx5SRxvzG7ipSOBq1mqrWYu0qJgkndI8rnP1JLhxB
Gnxh3yyWuBgJk7esCRJoH+f9A+36iZ8euN/7Kcd4D5H1xd2lWlxv6RtbYzSzwbL3UYPJpVliN7Sf
yoUkJFE/pZBUzxu+yypIk6RFHQOtVL1nmAh4+d7l4fWPFXmt024nNBzedns0EuWYLGpflsLB/w2e
ke634JOQfwERrJQHILl5MN+ya6obiNSkfyU9tj+Qml3kTwyVcrRSsEM+fNLjtgKKvAxrBwoY9qoV
/4Uh28BT1MOA5NJSPmdYWAc2Y7GAdN8LCUx0j2TUfFwZ08z5BJ9Mg6bSvxmwI7FuDHfFibNvs+bH
FyNBpDRMgZUx3LxFzLkpRoUhtw1o9nColg36LsYjorCGMTBA8U1+kdAZsY64JFH9ZXa85Y2TQEsi
Q7oT7KJyhY6kwdd1yNL+yQVVL+38/g+ssNnpOIFNo6qVSsy9e0Khz8vBW01CblSAkIojxfVsmnv/
/ekL9dLBH85+R0fsp6lwejLltYRQF1ou0hZQmf2Ll4FdjV2CJwDRaFdBnZt3NssynsMCNlCUseHG
oL29JmkFBPDPkuwaWXrbsyTgvfZpYtgC1gy+gR+ficoj6mglIOyeoZuvgmFo+B/uNJ3ysccM9uA3
v4uFNb0+Fv/9GpVoYrtMnmls2XNbXnRIydQdaxGgBn6htKliFDOgTpcnMq8tz0HzuknJf3+KKXPc
DNnHnLWfgrNGTxlCComznLgnvRP8PpjkXZj+YWuC6sclodxzTNZOoQR7frt/URZs/pa71A/N3HxG
lK0M5rPibH3IBxhT5kJxtvAhZHLEGNmaURWGPovnl2XIHP/mMvxDYOtVRv2in1ierFYy3D/+v8KU
KZVf0NXmmT+gWYStdVWZIWgfOmp2nYBTM1WG4B6e5dHELyd2L89q0nk6sBRMLFJJIPIyirIhmRuE
ZBNatg9hVg7rHaQ8TO4A8ysZhbxOP2JZxmF9zfWNbvFl9ObV7vP0eqwZylAiz7Wp2/iIcV95zv6o
6YptE8vWZEXY3+gLxrd+JpVYIIIAqinowbGdDafBn7Gk2tq1r5xDQygoNldKcDk+d4O3vArL60mi
tMx/I+eazTq8LPNi+tbSQBaX2L5ZWCHdxfyifPGeFg1TN0h33tgyyTgkMUipR/RPcHQuYkPMW3TV
QN/dw6mO5/RInsvkny75v6XaeBpg6jWisAcclZzCA1unKAbwIrLAjNU8VdK8Fj5/9P07iIxGgQOw
MV/8Zsw/iNeRJjs4j4tlvUe8HyOCXCrzkOdCIosLdYaMiVMpnmW+HquZSmx76EWfUT6KSyhK/FGe
xNHvk7B7kTg3iMxNgs4TOTy8YfDXJS8WWkutl3/2EiLSKnT+f9f50I58Tmz4YoZYC2juWylEhhVo
lQmX70Thh7EA0NXkn42hWOIvHWyzJMpBKZ1iewtbpjL6aQt5tNFntKRd7OM48HsfTsot4/O/Llk6
+LZeHWaheTS9rt9b/d91qrAgI86g3cFajA10YN7h4cT1fJYqYIUubFpbIfcwEPJeluNSZzJyWAlm
qe7N2Yisf3pFTKHBrwVVGdOYyU32DHCnVRUlD8Ow39lckiEdbE+FPcUKdmUcs0yssFmvBvgtfZGr
o4To3mjuuXqnBzRP64cGCXxQUSdbrMOIEs5iFBVIRKG+M6EKWSI6P7lC46A1FaWTRHdThONjoSGc
8sQwUVh7Om+8YTBCaglZQA2UM0SmcRUp6hyXnwhuFkTN6qAQrZwh+yQ/Dt9/2futnYH8ZLd+n5EE
1IZEcK40XHzkPcFpkjW2GGJa7478rTuE6U1ActQ6hJ7wHJIdaNdq6o1EvgGCerBGKRZ33kHdUWuI
d4pHXnmSQ6IHIVFGuYUg6DC3otZkPCGTQPS03pvtfgcFSybEy3HDeEtCwVXqy2VL5/Rd4NFDwdEQ
cy9+ZvlYanwFHlWan06TiYOKYn938dcEtThrIRcoOlNJI6bqmZ9hmOvMsXntn0r1bb0aFKv7qjdT
N6Lnt4dVfMX8oDX29DOCnsdWDt0c5/KZQzJp9dOFmubvY0Z4lGedqq6wCLKYvyYuL0TPiuKZAbSV
+58G2Yb1jJZ0YY6mXFO6JywRzmTLCHGid/0eoo2obJ88vjJk17igE3fbX8L7nr/ulHJUVGJIAdeE
mw7Aqw7j03V8eVYi9dfCYiqxIbyxA6XmGkvu3gAo+Whzfq27Dcw90+2HZQrga8tyzYoHCG+TXs+Z
0glkD2+vBS72rALxfy6Bj7Y7iAQsAGlTMEMGJ1ImRru7QJxkx88323zvN2iIGeLfwG0QTJEq8KAg
lJv+8NfdezmwyR38O7PaACVh4/QX9uWXZgAL4rp8ymB7rkH4WuqwYtAUXGRFYBCoTt61ZRsssnlB
e0/wB/Mwui7aUN9DjsomPStoniBqOpPXDgLg/eNIUbZU/SYCTqS04eb/ctjXBqGcLfy/0hUaSh/8
x3PpxpKtg3wizlPi47aoN/rp4bC1+PBkt4mux7weti8u3Fnwk0Oc8YWzyjhkGEMn1jQzFm4DKwnq
0pTijUtaRwzdIwKUe/RrXmfbH1Ml1zBZwJ3yL3eZiM+2/kZVNT/XCmrWBrr4k5DuIkOFGn0nuCzz
rJ9HNXw8nlA+Ayq40Br8LIkg0qaHbooj5rSAUe7nv6xVIZgGvlKvpssmUnhfbTDm0cy6ZAMqC/TZ
IexNAgw5080ftTre9zOtIwpxF/n/lFv/Dboayl2b2IaWGsMDOKNbdFIBNFO9VQyOKzT6VJOQ6ym5
wLv396avQ7rUaUUM3e4+C/aE3A4qucL8AxyUbakIv1Cvf+B4Mc40235RSUmthWVGTlP6MeVM0Hrf
5kLVrEHZbtHD4CpMDp0t4qAXHYM9ndd73sYEJcKk7r+MuPEZ/xDxFjFhG7yo0doDScZ6Np2tSL51
FpXdwDL/D9+lU2zefw2WVJV/sPOliHDZ63uNeMK8Q3Z2E7hLCoplO16WqhNy7//DVyhGbTKTDr0P
DAMTEmb1apt3SLb12ImyicExevhvSLBLJn57/jbxACR5+KF8GXSeI0euE38GJQh8EOtuqzyOOBl4
FG1qYKZa7xOOdem5fV1zIEvgi97xCNlcYRT7+epqilXEjL3RGJivq8jT7azKoS6FjzUo9qkNp1wg
P38M3BRZqq3D98Qi0ZuWFu8hrDQ4fW+d4G5vCmS65yvNOJJvFNW1UhKFjhW5UsylhDDgaOb/k8R/
V2vxkuEh4W2S9n6wUFsr/1QhsuaJSRhTB/y7RUV33ai8BRCTioRlEIuDuqBPx/p6FPhms8AzY/1g
ct4QzYTckFsS+nxTN4YmvHVAQMvTGhG7eTNvwHTWc031C8WSHpBSAl574B25XE0kBLZy3MDX0Fqf
RCh5Lf0tpLUqm7lZy2ZkxnlL/CkqeXee74O8uqOk2tIzxnoJ/WdjfASWpTZuWIKyDuwNf6ORcQBJ
T0NpcvwCaddHrCxaaR7IVT3ia9JQ/0U6edaoFwqBkkctUCe8PvEmDlA89bRyi9EzBlUhEcwYOh7O
QEo2sVFw4MlzvYZH55doa5SRWaqT9MVGuQYAHcHm5xDbchXh6s73kWbdnSbCYoKE4VsQ6Rw/8xyP
HxYjFS3MVQXbNpVv7G2iCsfCqHwLD/YLAIvaHscfVlFvdPcpkxaWS1y8X95UJ62rX/XGGtVO64K0
R0G19r2bnyvZdp2Zsmquv4Alw/s3IPd9mq5pf/giTvXl8166f9lc8GY9lof3vNLyuhYkPb1kLjGw
txa7I5X/NjukRJeDtV4w58wl+IpoMyWmrRMcVhDnPGzkR4sO8FTnIe5x06wezaf0K/DXKi85akDA
Hn3kt63OrB12/2s3caE4wpBje9EfcHw6ACGlUba0Iq1DUt15+lkaNdCyuZO0hLKiPTkUvaMM6dQ1
VhphR6jvbr/zkd2FkKncoayrqUsXEOl1vDYveovOl2qJgbvqU/+HSj8Cv5+0Q2nA15p7C3VLdSss
SBkDbBsqPFaVDtJlQezd8kNuyJ87ZPEFw/6mdjO+VnGljDv/RTp4blQCd+hHqIeCPXdlsJAVY9cQ
SeTscpeVVrybaIvBkVpT7BMLNtAAXk72YOsf+fo+upGTU0+VFzavxMJRuo1TfhPAIQ2QJ0rU/6Mw
LZmJmqJWbz3MyuJS8TRWpRbQ/Q91ipDW0ox+kAg3TSllLTDpFsNPIr+Hd5zEygAkiLSLOKonbzm0
4yCcxeB/nsoiCvtpE9/VgDNc6JwCcjvCZcTtFJXv2r17QEUe7wPfNGLHUP3+5wcepksB45VxJ/1W
Y/q8EsFLRqzg1YjO1Lh4qPl9qom0mD30GCkDgruFml0n7IOiBWFD0Bx9nFIAloCumYLCJ65k1hqu
O6lTcr+kbMahJa7BIMovxMoBGTH6E1O4DSCXRX+rZRNwYNfLSlyL6a4DhRLNfdSm/jc0U4h+jF6Z
keq0sJnLemWfyFH73VD3NIkqLB1Y4w9lqj5PToAn940PgcG+/ldErw1sdddqryXuSUXhgCxH4hZ7
xqj2iudUDpZN2mvX9DOsb+MNJ7MHlRJw8ust/zr1lw1Z47RHTIDNkWL9sIIExMlieP+w/vWtjEfX
pL+vHQ0xVN2mXp59TFKXdYMw31NU7mif/dDBPrq53JM6jtu1ioJzOwRET5iJ09wxiiWHSjiHZtyP
9fPtC2IBw3U2hGwJ+UL84gSiReMcoeejKxI7HXiWIYDRghv2LQriummsgVHOFix2jaysPMPHrG+/
la27e5MSsBJC5MS/P/xz2iLPFi/joAet1k8KHT09RJFR8qprrOs1ZFrQ5JQlr+92xcA9YeGEXCtz
t8emB1pohROOZkeNRPfHn6eFarG0z9r/vsgeWSRmAKSzZLlVsHcE7sQK3+68P/WgMjuqz7bmwyy4
cw8EN6ozuDa2OR1Jdw/qEdaIlTCOK6RMqJxAb4qMA9bjwFhEs/C/NYPEEpaosN5HZOSU35Lza/y/
VnzZQ6NajQEnLd7DYls4ZwphjMzAs4lrXN4GRNqK4IytACEHNQmQFQ19rM44FpiTRZgsnEUQSJm0
tj0ie1rw6Fw/r1irJpjV+QNwcwxMJpaLzsw4wacZCMjUtHZ9MI2q8zDPaBX0sJZJTO1nuV9eagWj
PAvwssI91AW5O08xNSVEtTKPVyCwXmFe7Ii4QLSPzNeqMYm+Mk3h2QaSKFuvsvjMx5bIVRdFIGbk
K4w57H8f4F+afwdC9Fmnq2CUxZC0GaFzA6KlTAt+2j+SoLaf+BBYG4P+LC9QFIe4+rgBmXJ9ucQY
ha+6OcpTDBH23Cdk0Eb9RrrsonPw0eBtxumS3n4R6ygxhYhwElextFl/sF4Ey7Fq6I3xvpAsHdWa
etxQThry/qSIgmU3/pUZNL2EYuJhOclXa7+5G3Z5saj7xVhC38JN/utLmkEQuMNN8ji+4fnNLclE
GW8nz+gvX3JCFNx7f0Z4I9bpDDZx3awwmWJRvr/sOGVqs0kfms4zTwHHOT/l/dyjV0lRxM5jpX54
Xs1ZrNnnsK4wFj8idkC5pxKT8R4EnvuzKzQ7kPXZlouwPi8qt3GpJTSwnad8g/g9tYZquj7K8FxC
ilOI5SCCRiPDgEfpFwwKG9ao71tvmQfzBVAZtNnGN6pJqtY73e5wOPWDqFqaxwfg3mVT7cB/TkKj
v1MBWzxNnjiezt5GpcqtoVvDsDX1PNyGRnb3Q0ugUnxGQVjXFTGkA7AEPLP81FuZsqnPQRZHHAFR
3GJM5t81c5vWKcj4ia1alPhiRtOeMSFeGOIU6wsH/oAayB9kD2/BLjD4gh82Gf/9fipIn0wI37f1
kbQRuCMU31guZkByxrfay1zgRGgfZXjZh5KisjNw69socUEaqPJTefI99yt9YhLj1gXqfhUP/rzt
Yr3Ui6oVnLQuRLrTLavjJ8WHZqptybbhDJcYOURKztmAiVJ146MBpCrF05It2hMyFA0yIlzWK45A
NkHC3oH8F+FfmQR2JJDKkbwMogcUMueDHM99x5Mu5R/Uiiz4Fpfn+fOrs9Se/TtIQkB7a7z5YI7R
zBqF5qwJmnUgEMr7BQ27He7waJr06rPtEyntfKlg3OZwWWvMR8qDyYjhF1fPqwqzAC6tCRhiKGQH
RWDVgR85TlnHTpkIIACHUcd86E3JQrLEkVNmaKd+KmA6Po5NPu3vOvhszw0OLMpwMfmeqsVLJywo
D3NEhjUJ4g3IjRWvfEQCAbhOXpENhhPqDoJgndu3hZ2SmLj0RFNr/WzM66205oFBjTN/Ke4gKC5p
LUnOPqlDvu1sdzTvlnx08RI6kf4r8+quVycwiNJEiWPzDCsCB9n6g+Hn0GuMoZ2SFTkACyPCu8sD
JT43kdiZ/c8ZHs1QtzbFWMAaU8mdZnDX+hN2HEc2GSNZEt7OeF8enKD5RKncDU2XabUJxvOGnvl7
9KshRVHB2cXLooxpcHG8SwxYTZIym8MtocYMpafMNxyDEjUsTj/XQRbd2RyJBqUmmKyXVNcBLJaD
XWobLpZ1NNFGomcVPfi1W0TSQWw8d5k7ssCvboMf9smfiD7RdzGEuDozaiXNd/vVAj6RQdTpa/Va
SIAUr3x6B4+jj8/b8XH9pr8SU2MLCHqF0BZSjfyrZM4xO/7pYm11WWvNDE74NYRXPplCOIYIQa8N
J1x0bb8g7Rsj9U7B/IhGSf5zKKKVK2q0ed3KSUX65O/2q8pvfyy3shMENgwpXL/w3V4x/iy5UYer
6uJgWFARzrgoKqTdsqaZstpHp+Ya6fp80HSld6w79pzPNYkMkt1bVnGC777qZMkBfMAqmXX8zbXp
b6GD9Ot129QpRKwTogdDdl8FRq5/ZXQRJWNjVl0dozDvquCpPgdZRwW4eyTnMNCXf1bimEZCmJ5D
MGcgl8kK7FTZP8Z8H3GzXJY0PF8b8s07UuubgG1RCnZ2eUlqPbUKdnoPQG1P5oBUgq2ZOHS2jMYz
J7ygH8PyqcQBxs+pOdO4HbcZJKQijLjhlwIR/3gRmfsuY4gX+EMZuXxbgtuz+v7c7oo/m0iZyfMA
mCaozaNt1Z4Pav2x9KRWKnJ/SmQwLdF0kjn/YXkn8pVEsFMU+k1Wbp9oylu01HD35zbd1hVFCz78
92KtPRf0XkMTbwBbQ+QbhLxwXFhJn4vnA7DWBPwm72eV01OJhMAKlWzQEfiuCAYUmbrToAnC8sJ5
DGT4gdwLqpabu/T2kLBToXOb5nsAAQg+ird5C//KmZ+vDCYwBguo22FfwhY7CeOXAfb83yqC7j6S
+MpNDHhurFfLUk2qjoUSvOxEOqQ1rpg8yzCg50WIAIWiDrfMUq2NVja+XK2TcIEd6xw5kq76F9Wk
Wp+2ClGzhOdKlrzg5uNma3/LN7qvN1v3Bo6hs6vFs9GYs4DRdpB45uosg48kDyA2IJojkvqqiFh3
JNjEXpJHbXjY2mfszhZPL/HkvNPzXfWSaAR4an5HHCtpOZKnSQnJ2kuxLraZ+yN2hGgEP0OXJ6Fj
22Y+QFCqcIDfBoI/arfIMNQjNKKlbWQesXt+G7v77za3nBKYVP/99+HQdTH0gV9kxvNuHvvZSbc+
XOH8N1BVJzhXQA4V6PFW9cNHut+BuKg2yUxrbqR597cbPoo4A533CXSKofDupUN9TSNZ1JWkknar
G/yetZfDuMG2f3yivGjbq9LjDRyDMO75OFL95naaOt+F1HwhqodFdIqJiPvmxXL8zSsK/fgRjS7L
TxKsWrFe+8m97EKk1sP6UrIHQ8+Rzdj4V9FjVRwtaQa716VREcLEHpYj5JoijkTgpKaxA3kt0Tbn
2MiydjHogdyOes+Rz16goe/IN7tTT2mdTK8IB9VlVMzhW+1YLJY6jafcMeHQM1ES7C/QDZxT1cMs
WDV2dd37UmntdbiR+/TbdikGq3XQI8dd+Gm5OZ3WZ8BEFQCmldh5+bcpmK1FjOrNTFv0xhx0v+5T
u0VearD0ORS+bNH6/rQjPBY3WRcJg3nlYKxHetcyfBamyFJG4KbW7FcHWwk4EgMv/hwXxCdPxTmi
82b54eiZ4ynp7SBN1ncyiEQgzmJwF7u3vZu1oOC4sy4NhjVVLh0oHJdm2iyuRm+OBfHhciL/Q3J5
NAf6l1VHWheu9xdHxwnyI4GfXqGPlFI/VGtX6HLVgJ+Cvs4158R1nC7+nG0gP8hzoXvtnr8+VXhO
u7XoJf0Lbd87463t3WOESbeMq6lT+a5T7CG5IxLDeQRtBlqGkHQFqevBCiTAi0R2Qs4/VcPs7WI3
VzxEROgONG5eKa6lx36ooIXout1ee3YSCl3vWAKvgj82Di+k0ogoP+OeYzJa9G7cS7xsOcb8psgc
f4xlbK/hZQZ4+6MCbEF3u1xOGrkzgj3E0+k/8OsOarSSL+cfR5SHhD3K+tZPJbOsHKrARAzJNHkc
lTtCj6G1hIo4EDPmS4NEivPOQoNBzc5p1m9dBjRgAJ0GCbuhK+2Oy6Y6BRocbcxuTlXjyOexbhej
irnvoY02cAppuQAT1r+G0qqptDoMEa7a4dUyQpeFx9swzQi3vj3uokCT8/z2aKLpPbviujDJHXOv
HYXpiCMrLuvsFQ4d7EWYOkJQpYW5oWTEplAJcn2JLGx+NZkdFnl8VFvD13GhfhFy+kiFLVKwtxA6
701Op5ViaIgXR1wvXDjhOVtHjFPTJ5kQ51UZZxe/aAfdnOpZytTkdt9LuOwhr/c1zx//96uBR0r5
y98oaAdbw1T/UNIoNI2eLa9+yaaN/eXaiKIrjwUbt89AAuGzaR1xTZvoLyX7qOwLrpfo2Ngv6JSZ
GMoYXMO3u4SSSPo/Z3biniMULc0xuWON/j4HQBgko6je96/E+J/fd//hzKftZMEl1gINp/lLyul1
dQgAUNHBlow2a7FLVXJdFiyIwjhwqK7AoNhwHXq9m7HstJ+cymywBg/OdYU+F2+UY5DO2HOHPLqK
7hJ3xonLFw+SIbVjBATjMdXczhwwryJv6Azv45UM0BvHYI24oIZKl/Jegn3IgBJKTQgLv2kkKZXo
oTSMaIwggeU8cTA53vQNtmqPki4gYee5QyLZRDDdNWnUV/dScCD4fhBIr/c48UM+Vxfoh/ChqDAY
mbSFpg6dSnuN6RE3bRHXVsiIUlKv/7ANz7MAlq0X/BEswyu51Bicga0o5wxKKuEyNGuzHZZtWSzB
ABELHRyC3Wo8OEWR2XKcJtP3FCxayfSI/TdFR9FbSElMUv2tfFKuXTbtlR39DSzHefwiQom2i0LC
lwPHwntXtCWvdnHZ3u/irYpPeAwhMT5B/D6vzuqN21RTo+hNp4EJIq1sepzxPB1G+kwzix5apzol
XRnqO9A4LyRIbZtaSQ5jWAm8LlNnKRxc3gjPO4ZFLjQqrjdqNa46ertFo+XQGc8ukb4sv3oXZs+v
s+zCF81E+/xN9l+80tYAl5DQAftdWG422ydny77Q8TdEFsf/AxTamgupWLqnjeNSeLAZnCVpSvIM
1UihW0qhnihEZjkqTPh/kuAnIWn3H5rK90gQW+enkzc3Zvturjnicnnfn3CVuwzlGxRyRqFp4SUo
6Slvycjrn5+4a7UOm3fLVbFLQ/eKVuakh2BK0VrpnyOeQbtZrVYWl+ChHtLw6QYX+727uSTCXL0R
KjaVp2mrf02plPOxwH3Vv0WVxacGzLSLnGoUypeHDIYLbfOKm303h053qvOzwOA+rvEoLkqYPXSw
2Tb5gQ9hWb/gmUDXVNSkVxNbUPDK5HtRwHTlA5Gv+slh7Ib2heVpxEDZn4cpeEh1o9ICwYC7btn0
YEQGFpe9tNeIJWdvyjllbTPEi3qRKY3UFsCpFXMvA5NdF6KnH/CBWsKH+4YcnVeV0QU5cUPpfhar
ha+3FaVqcCH8D6LWYzbtqHE2lttuRWC0+wbIACse8YK4ZG16ZQRpIG5nxitOts2oILo0yEJcpRZO
Skr3k3CZK6LFC4tIKebJwtevT6y8PZwGoGCtbGMGWd7cf2WgwrIgPi25f22B5vlXjLyI21PvaPB/
QmS2GayYUOgwjsj83mEDM6pSd/6l3z/CGtnLTCz10iFyLd9BHgr2ZqWTcd0RRGt9i6fQBvv/17Ac
NAEKZ/KuHPxS1/q7Brl7uLc1T8CBSwCldnCmLYcCn481qi6Yuys3XYe+dAXKViznMHyxJVAmRNur
98cfAJTXMg1aibqe2amcqhe7AvsHPMT/rabIQNK4nJ9/xaGPoUy4BZ4uQpSiYGfYm0f7L8kCIyPH
10fa96NM4MbdZAXrTrtfknax0C8du+b3TE7IbFy0wUsyUn/g9iG5wgiIL0pjQxVLmlBwnH9/wLku
9cujovOWEUgspLGBy/FcK8LsEFgYeKibebikvwsfWAjeBr3h1jg2T2J9Ncm8jPXYVNnil84yxOmO
3ApNjozZyvWwre3g1xbVuERV3/azghHv9Hd7VtXCN4GeiszIqj4poMlGz2pwaomvD0C1vYCPKlU0
NsIkFl0EcUP3A7VO4WZv5lYEboPrs01OuCpsVv+j46TiJMm3vLor0l/awhvRCQgYAx5i5K8hFey0
x6qM9rAjxrHCUe87QRx31JWj3ygtYEK8L8AUycP98t720KUIM5MobFSOC3hrKgJwkC/+5mbLtHkx
mLh/BBQ3EmsH/1iilzzZCadH7jtCozZ/ZI0BcTTMIGudd2ThfB1PRA2cSfmG4G8U64via6Ws/om2
/HjXYyRr/O0F91JJRJOW9Zd9genV7/I5RBNysbD5xSWK3oKUBEIjXGfSOuXs3WH1mmpr2p+pxZal
2N2Yny344Y7ffM9iCpOO/xRx65ZXX4ktpwfq3Ie8JebXUqKG1ElqQZGBN04t7guaO2r0wiyiUKgA
6NSnd4uu9ips0U/E3vMvmfeS8VNnqzRgww9nolLZjmVKCvOM49ORJqpZ6gVppcDhexdd15DTCyf4
GEzBswwuL9npGDQyNmYl7id+XKJRIdejDeAmwjwphPq4Is0jmOKm8TachEKnbSVMZgJFSx7JK5/o
Fp3cwOALhHz4f+Iic9eXnx2aeBIlOH090ZhHCgZ6EY+/ewgjxt8atDbqyvMkW4qgKrMJL35XvgFw
hMNy/N7CZJjQtqNNANG0+I78H/imRAm/SAlhrPZ+PZ8ZUsr53ySNxXcn2bAVj43L8vQryAJiopHU
LeJoK0V8VlBFolrGWwJFz+JfeQRmUYMiLvIbCia5qm0AerJEJ92vIhEer7yeeFAzpd2W2CmW246U
bLuHigPeHtho2fMXAC6Y40jo79FSsaU0f6r7qTJoOQxMrYKXcNdBe/eAPQxyh6/LDZLUVGSZO1Om
bd/j/l3r4ipM2+DjHsuJryaPSN9l9nWEslyJRzUHp8quirY1I4bKb9thL3MkEBjk2LOF4sljwUuF
EMxRAjttNEK8u4lAzBdDiuwFXbs5o16LRecFgZVynBh6S7yf52eSywchVXYhR4DIC5AXK8uaH9SU
rKVw0XhOTaPus9RE21elfV+PRqBtxe+DS5ZAU2M/K6gazhWOg0q2WDT5k+4zBI366GeBJtTit3rT
koE9lEKscoEo6p/FcQxskMQERFe4+ZJ768EPI4bZDgdMHak+iQiZYQqlPoAmtZt4Y2CwQ5x5OjTF
83aaT4PvBYTSOuWxBFaIqkPuzXmAOZaBsudmNsuI/60cGdnb0kalqoC8NfwTUug8IYgKTrFE7ske
6IlD+4NId+ppdyC55atu5VQdwMdCC9aDZGguqrLmbQCq+fTJsqj1x47ttrayySE3OsMJAWOpo3OF
5rcLojZSigGXEV4lUbax59Rw2hgzjOXLLlafx5oX4ro/c6rTA5Yc6msTq5ZEX7eToxWflK8fKtpb
/wHfnqIf5E3/xJrDWnu7AtLLS2oNw9ULdURQsvWcLFFjYME23SclMCkALaeYk5Up9/wgP5H3oLgT
526N+Su0n9dPXzAHng6axY1vaXLjXD2esrjnshHhmpJ5jP0aI+8cMPgqCX0+5ZCWEkLzjNyJcIE7
EPO9P5xGgIPysUFEEBb3D4Q6zerx/58+fwJ/iBeXI/Bi1mS7zAOOtoHZfWDv0Qdr7ehYo0o6e+QF
Z4BZkpXJaHH30sjZixc4SurT7/FHDGrj5Kje8R6gaV1m5wdnYTLdRdYhv1cZ4kII5OedAKa5SVGl
o92onGdIZR7pMgT41Ee39nhb76U1+cALKB3QQwC/eW0eil44331qeTOM42PsFSi198q6e+Y3d46v
Hqggiozdk4FB9kw/5hQMNhPcZ7TrbabhjXkakBrLQ9kah1la9KEoIrck3EM/ABDteajL4Qz9Ilm6
HCaTS4Hw/8Wb1xlpXgLbkC9i6VvhGq48z1Sj+aXVmeBALQHgPtgriAvErbC0aqS/3pgae8uw6xxo
ed5lsKi6DsaBSUhJ1zGpQO2laAN7Xj5+GMgno+M2HKdrYe5GzBI07NvGQ1MFVAv+KY+1qZ4SO9br
9uVrkeJ4iZICt+DuOwv7CSHXi/FwvCn141FT26MGPVNnE4T23jfBgfq+xIW1dNTJe56hUF0/hf0e
pMcBNzxR09nvJHNRGcoLSrknrOE4ReVHxhfML5WbGXdAelY9X4VSYKrsifm7M/PTq3oCIMmwVBZk
lEkjUZUi5BwjfKTCCeo2+AholdW/Eq9Ttz9tTmLLInhnL27QFTNmjdTSpl7u8g0nqGT9QvQj0BrN
c2sQIEj6fEbnSlMWgWDpiVv0C/qdNzoSiKTIiePm/NyGTWeXRAxh9/Ja3w9E0mTYAcMnLpENwS65
C7ARXEHFt2vxdq5FTEezidzwtwTwPDZ0+svY+ues8ct087itR93jMi7mmYDd4rg+chjdJwhAlq2X
ONze9PzPOrXCpuQL+xbzCjmv5SlGzupS+2NTo83naY2kUkDaoryUL+H3YHpaB0XhtMWvrWLmZvrR
vFBET3tmJYoMWjtKUR+rSh9AjcQBiDDIoBAm1345YpQZ9K+zv3N25bYAS8zu6PnsUxb/3h1gqijF
eF0jTd9CsG1RB2d/So6Hr7vn+MIAvpQHJviA/Pebcxwn/yRgwRk7/5/JesWnoNWGlydSPz9zGJGY
PoTvHYt5naDCCMjjARuU4EmeS2GXRuS3yMi3Zd65bdBesgvz3+M6/tCQ1S+qWJeZ6FgM8IVl0JkQ
ELC4WcbqoWZS0ncKR9rfYTyUqFpudiXWGddqhb//ouKFC5Jek1KYqN6VAarGmyd6aPgWkYwgufaX
XSxtHq1nR9hTiz1LFY/B8ddgJsgvWqWJ7UtcWUw3iDOkUW8jaCX0rIR9ZDSPJ3Y3//XOR76bbXgn
tEpnpcitS4guaLbqPWNnKyyFnZlMgMscwhumaceHAMzcoCvb431eUDRuKdenaADb3MBWIE74mIF9
8MVu0o+a3jQgmXDqRUPBPzMFcsA9cmPNalRV7TOJJGI4m1yVpaSC+WIl5W5GyiOOZ4GQTH4wj2Nc
FtPULs0l6cvMlcAAT53HfXQtM8nRA4C7yiWvR9pzvDm37Eb4ck2qF3yscUAKx8pOhS/jhjv8KgET
AtQZQiTtmOZDAQUmVs+N9zSZ0aSkcWhwnTyH75EwR9+uuj6N/cTvhypTfrV/Dhr4JvJ2hEBBFutq
8b01LYMRL5I+gtuvlyggDuAJn1h0IUMyrwWVEHyHxrv+YIfVN32AIMy1aLIY4j8xc9/P4TSqron/
J2NYZ7nuHrt3lQn63nuQcRH5NOUxnUcPHQ6I3+4mEnu8ZdiBmVhB3cDWuMQy519thfXm3bRA+aaT
h5k3UebLQ4DoOpcabyrVcFHav/QF5BX5KC8HT01rQGu41mggyahvGahjd97j8Q7tkaz2mVUftoTW
iZNWBsKDdz2PLXUI8f8Zn1OVVJ6zmhb1x/PRzXVBM73MwNGizKobUrE0BLrdIqo8xdtaCVEXkH0n
Dz1TsOTQyyTNfCtklj0yZtdaR6vfhX+jTOK6HnqLiqeEHD9n18UUB2wusqqviyTR4SA9eaXmkQYi
xvYmtgVWgH0CoGIojvLDyEZ0Ugmq+a6S0fDOlIsvrFBzEZfzzd+Gn5dobn4hgf4gkbxeRvk8ummc
36/vIJLHP1LRl6eFNCqqEp5chCvmAqVVJxTgu4TfPTHN7B+848DHRubQ3M3hzmCXsjA65O07iEJv
dWTJvc61TusLuy+DPQe+HLWmbACEq/PC7EE4iELvyIrvz5iPGZaTuTOwl9vblz+K7w1Bccud4Lpa
lp3GfKp+Hkz1GrJQX0AnXxeG1OGI2T4NRfN/o/yndADNcQA/nqdlVmyKxcbUWO/zlj9kb+Zk+YAR
++hu93UWg6RJKEZyoSZstXvgI17Fm6amkQiZF4qXcSag+IoivoSddsqLM5B1nJTK+tq1+wjxC8C1
jtcRtEhzy3JuJinqUidG4jFY293KBHxW3s46Z5Btai7DeNxEYoIeHHf+FVqwuJmZBLPVx5pvcxIN
0PQOcGICRivpC0lEDo8rrrnl2wE2pn8OhX2ovZzRgdNMnInrCRuUGlBFf5R/HRqicS6ZS9tuC+Us
kGGoj+eJG6TPUlXIqHVi1fmktr2p1PKC2DgKj9ZWsfnZiZVIQ6hx+SygF0xyHJPT640K4C2Lqet6
PjERVdSwzxdiq/L98Hevi93z1Myh3B1AMwYDfY5gH+ZfSPp38oRDUTsG1/GilLMSeXKUv/Ri/0wS
LZylLvEUmII/FXCF8MM2b5Kt7UQbIY4xTrq8FsGLCWfr3vcvH90Gf2XzxR4dbDQS7AUxrOXou/pv
T/CTiUH+2AjGxrV8pV+6PrHsqoiTF7woXQUNErBIuPQn8Kqc/GdsdiCEl+6n/sviTJx6v3p3Ihe5
UpojcUsmptY1X2hu5YmD8jxZ3KAiJ/LvYte7MEIXw/nYZiCuJ+9osYZDY3QjPMIfDsF+KjUeLpsg
yaTl9hYHU5x1V0BQsnYjkB+PrjKtiZZyVGlw7lbLFVUsDkoHEElloDDv3EiM22p8K5nEQtsn2vB3
juBAXZqjaZM7cUw6mq1nL9N1tdBTHt6TMKzxQi2JzTMgs+fcSws68xCBaHT69lQBVrGENtnwXMDS
4UpLH9AegRg90QJN3JgKR7OgpZidU/M0Leu9JJiinT8blFECavgnbp/N2X5wf6jOIOk7baJAdw2I
9Ty9OdGKAJ8XlkGj7EOseXGu1Yc6bUx7yiYiGAsJAigdrc7wCg0PuFGz5TAXgqCNYZrAZwykrrZ4
QE2AnrAwmt1zBUvwGxPsU0xAYzFHURRjIjVLLUbT6mvvB+wXxu7x1xm9vii+bdcCYB7aPL6og6Yd
/eGxdLLZPkX6Og02SYywN+rkZjH6hkxGFgdUz668MA/9fzbKAjGbxY1LTayWidT2kijT0UdvGJnA
HnVD2XINUPdSxfyj0BwSDYixxxk/aooxQNXIm0g6umuGIn38tJOkKHbtjKumG7yl7NmRwgN42n5W
DmpoiGVeKPAglGHXaHPiX1aZPCkDPxFDF4w8pCHCMXvQZZa0NRKOT8PFg0UCBQ+7yAE8cDPTP2nE
JNNNOH7frdRgFjhG9R8P2unSw+1kSSwSeNbqH/yYpJ0EwjjU8gGtOCJgCeOa+yz0Ew6ILNMjykLy
rbE9fZvw5zx9WwZh3cm2xUtG4EE2aRJyLFfdaQek6ij1NiCPlQA7E67ObfNaODD6/mKqxVojxxp6
rQY+tdGX96p4MFnJotDlUzql63p+pMShfkuL5aMkVkmAwO2w+cTCe9WKShV3B25xfjdzwS7p0Tcn
2KcNaIMX/qfPm8ejAg6YErCrV0NtwOp9HRUufG/kCyil7yp7fpqlRXPz5ioHw4SbQuhEkHtXPhAP
UKaccmxOXcBU7ilotPbLKXH+8nwpaYTVlYmgiHwxu7BkwMAgVhj6dL9rn6bUcuJ+fSgPHoJZYlk7
nJJfvZuGPmWZzQpeozNDU37VGMlh1xVJul+JRfWWUGPldNutZtXi51AfuHqR/fsBEBxD/xQthoVm
7WHRAtKdms989bF+W4F7CNwlT5ZvjNunC1jZDNdLz9IpVZ5/hpvxzx9jpIe0ZllDEq2DjFkFuRZP
Fw5Tf5IVZWUDrh6lURfzGsKfZBczUiWpz5O29k0pAJFVng9G7rrpEQD4DHa+4vcNZ454VaiSIny0
r6F2IjCyU9VHOOtkZ5SOy3I9z+X4YtRm6vyt4pE85nt4SgAO9BOrwtGQX1JT3j6zTdfJJNvUMepk
eWWbdpNhnJhIz11Gr9/hqXw52i9W7YRwxWMc0WdA383TuzO6XOF2V7ICxXqta1OCnCdt+11UDegy
ZfE0sLWBJUALPVg2rMeLhOKEu8DTYUnZiyFEpB+7U2IrIrTwTJthF/FATJY0PKaC+Uddpv6FHRyK
cH//NoHOidvBQFC//ZvViTesN07TS8D+pweGoJtECQbqbyZLn0pB4R7anLXsNitniFVTnozdzYdl
CUVA43881E/ZiPqIttnccN5Von19koLjytHOt/DKu318ysMxhew71+vAJC61WDtQyS/h0GUXOysr
GFuSr5UIF5yEIctU1xqxnBYVIgR7aeOsBmTBx1t9SWl9Ap7McE466WNyLTNBQWz2Wxug5Wapkh3Y
/ULlth45Q4S6vhHWWmRXuyQ9FmciMJa2fJZ/qJz47MLO3VzS8sGSDXeV9iu8Jww0sNtTyddsAaiB
+ZL1OD1WsCphMeCydhPchqxNXmb0KdqncPz/WQQT0rkJOjf+dK20SMD4vUu6L4GDXvMlA18RUP3h
bCCb5IgGFTLkNb4QQTl2DL0ql4Nr4lHVkCGaCtk4D7EN5k1QQF7P6cZqwxFrYZUJKBuu0hK2QZGb
MHjcb8RulEQOExZKl4rxurSf3ZRIVR3iD6gjEcVaEmFuMJGx4T/VCijP6Ys5v/19Qn/nvoSkg4rD
Vgl3k0eFo8mn9lplBkEElw+5W2pZuohICFGNg+qSm1jfnFWDZdstN3NWzdHhBMONqQhukiHLbF4d
7OSktkdPz7FKgKJy7HBNd12KzAqoJ1LZ7hLB7LAtWDfO5AJOzCI6GARO0VdbIyg7qlYkbfzVA+Uc
dILhVAl0ZmJNxcYXVdu9xeX/qJvoR4+cGDILSorwAWzryNzHf3t4RiFSJl1ChIMOo01hnnHBEfIJ
/HAxn8vwm2cgw7jjU9nOvr8dlQfqC2V7P+RDm7cNkbEAYzMirtZBi3trkqnMLdGvT199mH/ccB8B
poKtUiDk1j33XPXrntGD9aUporG0qiiI/w2Val06jZvImNnW4AhJGn/aoD2owrq1hOhREaQ3+yUs
EtUP8f7Z3H7XSgXFh115PIHjkPUNO8en5tbvbBRM4pDbasVP628bOSMAGmAS7Hyiw6YI3kBfXfEG
GJTLHskhSV6Z4rEPBBu6TIgUYEornEKJYhIarqnv48uPveZ1lq/Ic/dv45bcGOhkUSDS+z/FWI8i
5ynxDhoKHTLyMNdp1pwhvBNYULq94C8agQl4NghYbgvoJanoB2L0rOa3mjsrCuHUfxa1wk5MAiRG
KD6/w0ZNlVbBeS0w4ZPmTdynWR1nnPfIBOa2TJe2gS5Umt4lnONcF/SG7/H8dvN57od9FlgHMVOl
Bf6NzfNIDmEcY8iE3D2rlKvIbJ1fU6eST8RUqQ61Ow5lan8w2o7wtMb/iMYf7YTHzrAkqv+/k/Ot
n12dtdwXqO9hQ/BxmGexioGHXTBH/OgsKhpW57UdSERYIU39+x4d2pYmvbl1Y4zDb56Ar6hK1d4i
LqMy1VaL1SEyGc3DM0CxmG/ImGyYLcEmihRvgI6RZB/6ZJtFvr2GES/+R/qEegU47qFX2a0UuNwg
aDxsV986teuQDnBwOZU2kGDvrJNRmPOSZlviPUr/S6KqKtiSZeylg0Vran0Pwce4BMgUbkdUDkUy
ifALd9eZdpQftqyGxjYOu4SZv8YtW0JItFeSQQzMGhZH8lA4Y/YGkd2GCBU8zRvDNb6/lrjbLH84
3ZLz+B761omLvLgBhK0sqav0txp9uC//VXQwgD34olPj6IUkNKOEwDXW4hu+pjcBwl793WH5bYLW
BOkry0UwOmG8jfMgittFiu//yDoTUlgM3yEO1r3GC4dr4riBvLflP/3yo4RD7QCsL3pb9+F8VVdq
donEL/McrvQmCGKux72ET+5mAEU7fAzZH4KQVPPj9gtZ8fh6lXTq0b0J/ug2G2lHhFRCVDSIBpLL
i/cJbOtN2fEizM4e3ST+b3GLfiqqoelvxOGrC2v1C9DJUmPJyuD/NTkVxag5tKpEbVLVA2zF/Fhx
M65cdg6hduCXsCW8ElPdnxDEajNaS3iCQMugkM8NzjBzdqbnDDRUcoYC8dZumpygQ7ApwCCVrOLM
kYLSzuw2vzylCgyHnWJkkEE0H3UQtM94w9xJbULyqxlnbGK4heVJ4EGZbMctAzKuYYWIP4u1PMwn
51BJCU57M/adMrPxPvrcslgWSpFhyj1Y1ACzGG0/0TwR0DO2s2usFWtOGknpf6alwb8HChdiuX/4
LdJZXcYsW/VrlCGwu9BmElQ/kTOoA/q6PLl9LuJvVJ4H0MUIKieni4MIDrqb/KZfKdWVtnCbrZBV
rkMxYUody0fGwE129/qJAZNWxqcldtGVV07lvcGgNT46L8p8FTEc8RuKU0fvb/va+3H5e9jt/Qna
DUI0EnxRAluyEhBxfeP3Sf6mmU5AGDcG1bJKnieIol8gBfzfpgbPSGkV3Nx44OJXlWo+0s7rD3h5
eMlRR5at6yAyV1AgeH6SExTpc13ry7EStZnYPwGXo7CFaxDIBak4t7G8OvqKZkdHRl+QP7PeQRtH
U7BipCHxj2rHfOiMj90jA0ADHZYB6iRdp2dymGUoRmk7C0328K/fhXJeF10pPSTeMOpCN+p69GDn
I3XEcmc9IBsCyB71sRJbCski/5Szpi6fS/V3fMzPVfHZng1+OD32/Pk3bsI9mYfkb3WAvPdxV7be
zXAvmkJW9vxwsqq2U5mll8MBT4eKbCiN2BZj8gn+zeVTxas+FcV1Pfvj+FBgEvU2bPFvCi3e2p9z
3pDt+jtgUKSrw5F6v3bRP8aMGiDDV/e+kOkmFU1ypM4J9GAv2ZONAb0+4iI1jbXGORaHd0C9jzMV
InLAOrtpI3kCarUQqRBfHQ8C2Wj9yuwfOlpW3KZwRtBfM71hMtpfuTRLHsGVzCUTwnOxptYf+pjH
4o3yndiBMf5Vf0Jv0l+Sou2QIZA1YqtGkeRm7AyD4P6AQuEKvlSwzXORK5rm97DkpkS6QF/sORXr
HQH/GAnxmcf+raFwkoy/8ADG4sng2EnPcQoCOyogKfyDKm8r6WgV2uJe3Z1zIgdFonVJV+xFa+oc
Rfi3LpZcdXQbu3847XLv8NeSiemp6cI87h16Ls/d/hqiFm/727HDy0aWwVC6V0xxog1FqXIwU2Ek
yjDG61ijUBRXQ9Jhe+ELns0a0LXiS22HhU0pETJXhEXN7oP8MJ2fTBUxg8S27wOXUEQej33dsZXn
BPWEnmnGgT8pg7kLxgMNPqb5js0BC+W/GTq3qPfjKc/Yy2vJ5+WnGsWlMYvuihDj3bC2BkCeUsHu
xeHK23ZultpMNMjr/AbM7XYg7LBPo83TtS7CZ5DBKycmISvTJnGlQriJhRff/WNWDmM8sJjBW/gY
0A+YlHGkvcthvVxbx56rfKjclHoa16JRSo7GkBPKPp6z2RM1r0mpJxAOdAVxjfX3oHXiqIckR62N
CmO9V4dL1hcP6MadGeDfIX8//zujsBV4URnB7UG+kAWa//CkQaw5TNREOkmaLLEZkHAdckDCXlLn
5cFcjxGF1+3d0RCEOr57DbCaVT6kvymfMA7VOVGp+mkLioKOCOCBY8/v4HOPGy4NSdE1jB9HeRxZ
zNJfi7IbCuxiufSLHa1fKruJsbwqJRAZdJcmqfLk47ANnKmg3mcDcGGV1/CsKEqa74y65K1b9tNo
6B/aMwUzgUYwwt7HjNvCY6WaIx4LU9gVPG+yyAFPNxy4Y2yKrhprfY3Oe/8Yyw71LFXWUZd+rldm
s0qNRLSsoAcYYiSdd8tUVuB36wd+IrdTG9cJqlW3eZzdexABXkGGrFtiJUSsaRXi0W37qRvkTKmR
3Y9eFgv7np+Kk/VKCExVJf2KDdYNkkzAw7PxpArPBS1KTn6i8jQY0qelL9g+1XaaXu/qpaEcRbsJ
DzFQtZpss6IQ0pmAAw6NGN546bOJMR8lW9cKVxpvpPWsDupSNghbTUUPZmzAUkLUji0o/wSs51HH
XkqnxMCXeqWA3K36Y2vcIFHbUQIRCiRNNxS2XnhWbDeg3Kdq8bPUFvc3N5Q9kCs9CGApVH9EMzZc
I1bA6ttBZhwe6mMze6zTg4K7o2fzu9sX83mPPaHvMEaKy4lp43B573Dbmve+UYapGcpsKkct7yjW
ORPxMOkvYWFpTe20SYz1/F1jmkQizUXCjqpag9jrHJC+qhFfnj3AvH0MJGk0xe18x3ESxVloyaz6
1EiOVrsyYjH9U7gX5uZOtByq37ZRoq9wFh6X1EMFgFKvwUnMIL8DwRMCcN+VD7SJW5cfk3VOUVm7
f9tfZagUpcT5VgBBA+NcboQH95yh8iQhmvh48PA6az9UwcT2PoRvpQilLmJp2v2a19PIVb9YyWdm
MRGcj1jQTUyyRj/50yNZfFeqAtIP9M+oXPe7KieMKDNKTdq6KJ2Eti0cB4MuzpMolSlRejh1eenv
QV92YrTiWcw/oTVeWUf9s0MEeHTbn9R3ZJ2g2iMjYRjK8k3aAkMY81YpIAxYX1QafvRgWlB7rq+0
NHRUxlhQIRFnWSYlTd//EaXhVrwxjn2XrB/e19QVDWs5hSX9wUg4brtxWb1orm6Zey5Ecee3zt+w
KQs613C9Ap/ByAANMryvXjzlHco9kQYRZOaqPag0WQXW+dEEQaOyNm5zm/vkNqQBTCSyGQNHTdrd
I0CiunjCGYq80o5LvtVk+XkLXo9Y76QvV4zkG8uEHL9WCx+GCfncXdS5sGlfWiS+ImUrvvcByiPH
Ejuxhiy4TXXSnMf8b8sJM/L5Js3oJEPDfATPE48MZ15f/5LB+rjOBE/68z7igdC683LXCpuLZwO4
KpI+CV8DoaZox8KSWl9RivF/Mr7eAg6jMEGcGgIfijW6Yz/Mt2dZftFIVn5XdkFEqRBlwp54wosb
JLMmL0hTZComwYn9NNOQfpoCUP6pXguARe0mgziVmyHJYwbw5ScQkKyYZ3KpSlKtDcUwZL7jrJFK
C+rLFKOv8hk2OZrdfDTMULGGeDC0Zs15dAYHzrAdM1YyIHbyXlXOW2xjyEPHguyB4QSkapwjyEQk
77HobzhgU8/ZuS0P5jrKyleIOWG+X31jN/u+X1MK7oUKo5DRqRIXttd7lMpmn9g/knx5rn6gsPJs
UsZuihuhNolGszD9kcXyaVdb3TpXi7NfCzB3E9Oldcj1+ivRdgcRI5PebMcFG7O6k6D0jXCrnLF8
haqRorB+Mj1rlBtB5dqFx7D2VJCEdHpoefyf+ZsmJUeTl9b1UKoMf4QprPttIf1v4f2+0RH4OkxC
6+tG+FjF/oxc31TJJulEc4YnVuJtVj2rZsoERGs4QeUXF3aImq7GwZcDMwfV3JAtSGsluX7eg5TA
RSkgekhA4/N9oESQuhQI1vHSmpMK5gWCCXgY4ZHrj0bEI49uCMDu8mRzem7YvL9PWJm2SrjktlNe
t+YxxwuUtNvfxp2/cdryloju1Lx9OiziDSCnATQmfLD+QwCUDaRq6h1EPCr15iq1AOJcKxMXkied
D+/8ZJ+NfZDUG5nTS2JXOkKLGTUoGzagXCKodvaejjpl8Hmp9UlaojQP7uPKgQc3IbcoU+HzOD5g
k6IjSiuCYEq9RVfaBionztx4/cuX8YMqvtPY0AHbVwt/fh3/hUZUchtfVA2FzTmA5CEqdOlcHdEO
XZ32Sj4vchTTTziDVWcU/J9WGm4PeqgqQiI6oLv5YL4q9fxw8edw11CHJQopu+2StDLBvwGa901v
ZTkbTfo4kTk1Z5lXf8WxgnAiXpHeIWCG5RgDOnPt6APemphKz4i0UtFA8rLyWvMj+YCPs508ZHdo
XsS2jwtkGCfsbdktaH+dEXdFqSDotqXNnkI9qI+K4lC1qw0uABGOv/yGdsEVhiOZeMRs3OnpI5DH
ObUSuf8wls8Bv8TNW8RsTNyFc1VQxp9DOAyNHuk3v8VwQtW6Y9bR1eoUym/fg38B20Q5rCUrjDC/
UGyHBibVEjMk7X3lQ5wxx96BYEoMkWEaaC8VijcllfZvOL8tPp83+g6zevRr7D6YJo+sDt6/H1Fv
yNnnH8WQvhoj2uFYVwRFFKUq2OTpJlksjr8ylUWrTbpsqsxQliRzGLjPA2Logyx1OVHH/yNFKlK8
vHG52jocuu7bSzrOHRLuHXym0vUjn9SxIBZaPIRSAqs26XHsibURGMYiSiuj2FekyP+rSoe0wlB4
h2dw+wrGz4/idlpn++MU+Fn4U/lCe1p9rSGBkEEXNctC4TSokaNow8AYWg+082ahG/5siQ0rwf/m
L7BB9InJnqGQZkveDmgXGeZKnaQ2Qows4gbl6KNm3wkScddQ29n3jZumUEbNmoku+jl286nbmHfE
b4W/Mat937DdmGJgHsQxAA09pjo6rC39eJD6mAknA9SAzwAySatJp00eFLaMQOigyjbp55LcfrDE
ATIb8hJIvkrM3k3xQ0w7opiGq79bCMLOeADO/ulqPScgCuRfb7oFCr+yhflw7ejuFLYQb8b69nQq
oCx9OSF4R9q0xFgapiGXLSURM/Tb467HJ83iemn2Rh+wJLmauuhWw3Mw6VLyrMPaOSyrp+akUzhl
/QPxOof4JqKQlhmO3nVpOGK7bL3gfKOtn40stc9T7+BhlNwVMVRnD4VcLFv2KtfPC1mmCd9hYs5g
gbNu+K7zIDtJbi4/mREkdKnHRKNhvThA4yfxq9s8XGu8I860ldekYUllP+5enHkGTZPaXBNP1GKt
Cw/a9XKD0XhcIVJVbbOVlsRGXBpajrI891eQcGkM8RCAldRcyGUzR4vhAhYx2gefb+dw65oGS1sY
0HSnkMmWeUOMilT5KTwXh+3Wn1ZSIEcgCHPBC43HIzC3aRtXtCkLG3cDRzF5o3TedVKQlBJEn3Nt
y60ycxzM0+79rBBJ9GDrrv2jII7vhFrx6QCa3WvJ+pV/c/ApXR5b46o5D13IhQPQvLs1SqfQGMjt
65Tw6S+OthZzGPQNpyy6oOe5wh0RKCwrknQyJVkDYcqpuDp1VM7UY9KEP3AJsvUF5GIeaac2Q+DF
HM39ZbItY2xYLoKk29gBL/yvOrszjHyZ/iNQ2wXG9k/Qx955mlWBdbd6Lf5v8yhaERmNSWVZVv5D
iiWUNYX6B3Q7eV1Oqko+z48j8cvpecTkMOjVwM65IqKyEyKvI6hILQOeQ6pEr2GOx9sSx4zZB6X4
mwI2ClZZcExm97XTimozzwhnwvguqISL01i+p5q7NJfmlz4J1Jkj6zAXg9wF5UTSXVXCjKTo+8U0
NLYTY+gSd3NF3H4vSvYcYEcRjyh6HyIpv9nNQywYg6N3KtpUh10Owk0B1udTy47AZqvUf0KnUeJp
WSkRG1baG49LtNYAarAl2JwwDQAqggysl38N1p0VoL93Jo6IxkEg0QQLYRC+Mm/CgieDLD+lvT/Y
oxAhPyvJ8ScfTWVOfhZGRE9Y94pmYcAVCRV5Etup5IRxg5HkWC6Te4i1vQ1myUuN/HIWBpf3YSru
hBQFkkbQu3M27I8+HILyIiBekH4PQfPXCSunx7GVXEWhorONHsBhdhEQhShZBc9QgsCq6HmP1t0M
9RC3eQlFCD8Jau1Iqt72BgCF2MKO6TO6Gp3AGpNIucv+Crld2WlX8jLOEBJyujGRL9sqMCi84Qpj
xBqFJh0LKAMYMOWrjfIWxpS3XsUkIEFh1MwG7M2WBDqjIAZ7oGmQ/FOl9xYb/cMUlNxn76z7jwf+
X1cvo4/jmA1Iygvp+pX+9Oc2KMwqs1L/LaKciv0FSQ1/8/xuoGKtfOEEZr6BNM9R7wfPDduLSj1e
zE3uJNdREfs+vQ2GcHz7YcxUqE2G0ZU0fPXuJXbxIQKCGQI0kdfdFuXZkNZEpvU5VIr0gnzg6iEL
6vx8Lkl/HI0gMbxFfFbgPOnQLB5qGAJY7y7zdqDhlnCaUGmCVcR3plThmkQFM9CQ7Co4j834/6ld
9OKAlXRcSa2u6hs1Rq+VZXxu/fGvheIxZkqLDH69p7x/iRO7M9B0o48Vt3azO0JvBahy7l1wa6nc
qIMCnFKFN1OluLb3BeB4rAo3na8tQsZmFQrG3+6SWf763KZDQkVzP3VdjPqSOC1Pw8UL8U1zIj5q
xXzjRM0N/zTl5dw0YdJRiQleKnCi5oyDvAwrfk4gxko5XrQXys++VQ2XLYNuCxKdF7hy0FyQ7FzL
lTUK4bYQ6GSVDmJlz6wEHr1ntimnxKMIGCFlPDj+bwARsyW7LYF6rNsQ3rVMdFscRdlfutPkixry
t4vpiG15mbzzc7lEjLObu+6cDAnetHpFWo82it1qSDWxcMwmGqaX8Ij0ZFf2AtYZAM2Dk0ouTa4i
GoEx1plTD/RfqQYhW1rySNXTHvav2vIYoEmk7SB3e7AidHPWLhxQ/OEFNzzKqIxvHmIxamudWhL+
nU4wSHHAtmcwPgn6AciEV9l569/JTiolOUuL5RM+ZOs0pWuSM0Ayy6QGW7EmIxKqtZrry+rqTwj9
FdUX/znzAPmB4QKeeWLUZn9BVT56xrB4hAmO1lbaOEqmyDC/0w/rYq2ReiqkT+CBvUfQMQT52Ep9
hclih7+iqYcFqpnCflbUXGc5C6I7tzidHB03qGy99B/TGdQ8ME23q73GySWCD4BFIipTbpG7iEyw
QlVKGEnJsUhUtLZGtQIssD+HBhy2o8cyEyB5b+Ksr9IYQM5OOQZXqCQpgpBTp7Y31hVTYpOPoT6e
nLiMokhvY+AZoN3IRKUt0aop1+tDmKKA7X6tnrN9R4/Ooza+bGM14QzLMqCbpz5yOSnkVPPjva9W
/YRtpyRflJcOdQzDQTWtgXojjU04gtNIHZpvnYrGw//VcCyjMr6Rq1qbvErTMIvAWSeInptv7695
sDkuIJXHd3BJPC8jxGCWFoenBoE2DYpdu2ZUyBwDc7DHFZcgG0JNC0V7hwEXmUXlFIhE2WTXj5pi
ijw9nUNYNp53ncPcwA1cs+wezvNhBpxY8hy8UCx1mjMKa7SE4qn6LjDtxWPyQAZxYX4Hb+48MEpf
bB1F2pPE5h8JRxeOh9PNzh1+hvHtmbKav9z/JlPSINNue2asSt+kiN0FGp2X+fHACvCpA+T8DAW4
RRyG1/YDXcjjAi2f4o2lC727wudADLq+8upNpuJTwRIxvf0lYVOHjkOGhZdwIZAvjREjJZMRParu
HDQSCfbgMUrJ2XUxkkW5ANHGhlwp3mYDT9sA+ogc6iAmWUHVTEyWf2HvJAfkjJb/2Hsivy2hOO4t
t/6CUXaIKsL6LCJCUcHDsUh2Zp1rkF++LbKwH2R4hlHp/0Vbx+DpVkYrujR8j9Bolf3kL4vt4g03
Zf6yreu3+TRDW+9GRIVztCl09YvH4x9aIe7rGNDLq4gf9HeRMGprq9mW2ijYS8gVlU4h8lQV23KW
s0vUUABYNT9BGJnXWbVenggJGlh3vwONh2FKfCwofFvhIdVBOUaW+E8IAJrFd/uiEGBsIL6ygqg0
oaVnDDSMWCRiaSz5FwKMmgolEvvkp5tWnHAGLVeoNRAvLXVgIth0WPepIUDwsfQA0viNNjbWyrat
xb7d/BKYkuRfdvGsF3pL9tAOVnTtEevtZnsrp2nwz/VLmOkK/7oitjpBOcPV70hr7Tu7mFQh/1WA
fe8sQVzLjBIvnqR7fYMcondYaSTRH4/MPNfYRaqgCW8MN3AC3xmxTUOGfN0kF6QGSmdZwNyovx9o
ELiSecPoLpuH/uSpATFLC48ZpwUDD5pLK1p9Qpq4URAn85N5EYHXpePxu9jVpQI3H4U11hggA/ZF
NU6hJYo5AS7qCEvTgLQmTaRt6M0ZrnG8xcvEbflPO6KRqXnHz2/2ACMAVlcAFFGCGPgyAJIg5z4W
qHTp1z7sls+QutFerBDAb7uwF7wkgPhgWgMzPqVGh+2JlivKLHW3XuL1A0tRFywUBq2brMssqdLm
GdhEhd7sStLADWdBWOuJx9e/ufpJQrgo6pZSX3TOjELlEtnaLnECvcMgqA6dnHM9M1d0rMqniUmw
8P8k7wFb8YZ/jKYJviqUNUqR0j6znwIsxALU+wa0PMVBjyslIz1hM7h9RGqubY+6cXhXnRrHDUDI
nWWMY0Actzba/d+JAw5hp/HYycLSPOu95Sui7sjnqghA3Sql65dB24lM16n41Bg/DGzMsmDeVS0w
1BTqYdTuERE7T9iG/qgFGi7ObXAAKc9vFVYOn/R2qpBvvYNC83alsC2LyS5B6HF1h15vSvcX+Kj+
1ZjRx3clW8szaO5CGQDQv5znxDMrH5ef4pzMnApAfHJzyiiRz/81i9S96MFY7fiGM+H+Qa+1LVbU
59IqSf2k0W57sjxZ9PBoO9YLgv1V96HrPKKwErEO0AcxC6h3IRXyRwsqdZUzv8wuRy8ufs3w1xoe
xRXv5GQOfkN4L8UAaanq3G7JXOHsIPjDB+ORpzSv5+AkQBR2ICjkdy6Q6olrwXylv2FkqAT2l5u/
/76NEHzEi0lHf0S/TEIJW2/TZOLpVZhZtL6LhNYkHFqfZNhRugVH/AAQ/vuoXZomiUkfb1koaGg/
gUTzwiIeuxlxofqFJ9+HhisWVUJfuQXEtVDQBcQ/cAak8cB5TN4/xKJPOG0XhAlAvlYNV9cZ5vBS
bEMdKzC7cwbpdOBtweE86QxiHqAOh7UlmKUHxdTFNIj0Fdii9NHwxwW6RGqGAGIl6dE0sRil6JiG
DgMPpR5UnIUU8SES0aOPJ2qwqIAM0TjQsaBQMKwNFB2U86XmTDEI3N+8/Y0DeCpMEyaw+5WSPIwe
SpAQ904dEQfKFGS8aXz1Dio7/0PSLd5yHhr96kKYtCY/g4iYOYqTonrIWdSXNLOb1aQBqsn+b4hp
goWnihcyLnK0eoOJ3nt/u17Hqu62Oq3zr62KsHSSIcU6s0pmn3LkxeORmzmzDfVUGyKADu7JcZsY
JDgMN77MpvJwhgqT1piPqkcik2CQoAlS7QVq01jLbp2E/X1cu2Eg7Ynzduzew0X/fOa76qhnqO1g
Y2wZntCYheu1t0zn8vL6iZR0OhXCfysVZnIacmJeVuBgT9s3bLRcIFd3aCSUe8Za14zPeomay996
NUMozj4g963zygVuSSDpVsQMmIhD85t0BbGigQ5N6K0h1ZZKv/Y4yEIqpUUsSfbu1Zhbqbrn7ll4
FfleW5nKw6Um0pcFTXRiHY5SrhiJMfoc04SMplzLbfoZoN2sw5wZJW+GsiNBInKO42ESwvBsTIRC
Emnrw5Q3ftUjVYdwllDHaEFpRkV5f/vlqa+Md7yk+pyqpKm1Zw3acXIthguOYC0a2mC9ch2fm8Cs
j0WhzUchlANuP/JEDvpTlO46VsaaN7+mRNqN9qoPM/OXVGf8/UVp4O82Y1JjYMJLJXOF2tAFlIht
x9izQzKhhfaDBNaIXhuhLb0tkslo86q9jvsHq7H9k02TSN/6da5iZ0kuRMY2hMnLp6gOonsnzjAn
VYBVW0uxAYOxNj3UqYgsEhnukgWIdCsJLfh1K+46rrM+FLICeSli7PmDXRIXV+LF5QlRvTlHp+iQ
0GBSYVnTkBsB+7bDFMHA3zFlzHpGPHr0c/dqDb7IYLL0/z4mrhNNdMlDfSpGO/UdYltCFwc6CDZx
M7xdoIgvcdPam95INiCRQyRUFW+pSUGQV0wVOF1V0NcAMwPzmS5S8j8trKPBGPByHJ1+vTYPyuyz
9OUUJoVaTjRVRe/6cFCbmlKJRAsUtYPZ8Htt/k4uofve+omIMnyE8O0t2xWQqzt4zjPiIt8Q9NRu
nLLzqw4+Ui0NehkJXiAxdyWECxkOFCTS3H29vRCe0Ka8Rn452SzZr3fkvb5JyTKup+kBhXPyyd+V
Z/XPzQRnIpKQr+3NfKuB0eFw0jPz75lLim2z1OCuU4a4JMhtW/aqLqZ1n3jkW0FmkIXyNIY93pGC
isbXwxmmXKpsInzg6ofRCHWaD0cnlcogCRedkYD9WPW4Ojrb1sUEXQWUWPQ7eglg4dZp62t/LeeW
ENQvRb85vLhs0TybcwtJaE2CReKrqSXMHX3Kj9y35nuOhagIam737Kr+gj9cZnzYrv7l87HjT/pO
tgEE8do1luAvymjIwO8nmo97YpV9oK2sbGPSQFt7EGGEnpiGV+IV3Wlms2VFQ8OeipWOJgEYuXhx
NLMfmyAXBjMndBMl9Rq+L+Kk3y98mGXi2hfd3kY074dFFklZ2JqXH8o4YGBnABWoFHjWhwqazzG/
Ji+aXQ9uZJ2CyIYmRe5Nxnx3FacNF2k8GPpkorkPZtadmbWkTieGZJBOEengY1ypWySk/gzZUOZ9
hvYyTpiH2v0V1ol+BHqbqDd+a/wzk+pmSI6Ppcl0Mh8buaEj6izlR14V1JJ5sVL4Q4d9se7M3cll
7jWwiwwy6HLfZuF3pFJqnhkGo4XD/dvgHaM6ilioGdVd1dUsc5R21DkILXb6qWGAY01F9KPWmBpO
fV0/7+vLAWn95YOXAF12Hv1s8AQDaed8fD0NivTACAyAy+ugwt9zvGB0k9yVBltfpsPDI/2d3pT8
MKG7iMH90A9z6WJL0qMWRZHsm5U9v7KxOprIDKkHUqzPJ7P0V+kXdpD0DVzkdmcGupbn+ItbeXX1
jx0M90CSH0lMml5WkMdqChpJpVyUYAGGG0mrpRdlkEu+wUDSguhece0QVYYWBPwi+QZU4koQmnRR
v/MxFVMiilfGR/vcWTjEVLUyCnhUziAZ5YU1K1Cuvt6i1LPu432Q03DXNPLBJpGbwfRdiRNqZykD
+ifD5dd2IsRksAmlpIX9NTAJYJFe7SY1h6EqIggUpsWQemZr7mJs8DMhiDVWC581AO6Jg/DY/wqO
35OF0M/b/EzoqXEHLenoqs/UctPIX7hPN/43w65IVG6pQw6UfwlhZVsMcpZiCj2HGaMpSysDIUoB
mAHw1m9aBKj1L5F3AkV0M7wJ0PVfilV7Vy3FXm0yaj91UYCUuYozS03RvcSjODzKUZBmaMmf3f+p
Un/aBsqbrk2xAtEq4SMyapjVmSzxm18ttZJIG5161OrVtflxIibY3kbGpsCyLUA4eE42Qq6Sy3od
okAyXyTCWLP9E1lgukUjhXHZXSqGQadXRk47pRjTOSxvQW3OXzxGcKEOWf4MibfoaL0KqtGPVenO
gvqQ8TPRYWIc89FlSQL78GboTw2FSbV31uzQrzw7Knil4mheLNUDtSSlGAAem0CtxR/1sJ3aaHX0
5kzfrd5JKVHHxIObOUq0ti5STe7cGjwOt2FOV002hypqL2tf738l++I8vPikelZN7Qo1qLDjAIAv
1dHjQpZtltSDyMLwrnDFYjMyXYgcMVVBVnUjcv3Vqj1J1sjWEKGfhVOKolKWY3Uoy86po44Lq5m0
EuS7y+21u+NORnJubAI3EhEJ4gzL13kJu/tlRQAk6cOAMkbAuNG4UPc1xucyydSoS45yhx+/k5N+
xH0Ty02GjtECG/wbB2bGVUVayJWnKNAIrFhhGkCyHy+TEl8mKaXD0nCNNaP9sggHQnq7HdDVVhCm
jvs7lsYScONVRpBuMGD1yPbcwRpgcDeWr1stpFRwkKX7uH0xwbfzdAskSuMUPqToLgxwJuomYuch
BRcjllsV8zpnr4VGXIbt/krbev5aIrZ2AoMRa3hFW/GSQ6FRuZ2ADPRATySJEFmIa1KQZoNngPtH
0AiAqML5B5lzXDMAzU2f9izKTaaVLu/zb+u5U5uamwkUAHYB2Y9oSJxOZ6XkF09AZLmfDVaca1QW
wCAWLVM/il0wK8BLyC6pCYBqeFsmnOAtIZIR7/MTb4bZbIQ8lmCtMqPB4vR54lWNOrS/8Jy9VV3h
XG5rSF0pqBeaS4IeVnt/Z3TFC436qNsZEYuS3xEHLrCJDiOUyZzTiJd2VdpBl7WqyOMfyN+7xDbA
bRw9DeZYcgyhRwtvxamlVxmyNBBjxnzYw6vAR32m0q3ItdhJ+HhGDreY/pfOeMSF/DHHtxRVZsLG
ala8Wh160W3gy3JP5Wlv3UAJc/vztm4i6FblfOG22RH66kdwkCcxpdR2nkW95ZmBYlHiC8AAVmBD
AS16A67UuqwTVAsAuyPeUrRVula5fgKb+ubucAyKRJnWfKBJW0StNPufEXiW31SJ5JLeIbMWz+0N
Rk+B7StiIun29m0pNxCIpyA+2+rbcVcH7hqv7aHPpc+SMofERfK2OT3IAxMrxflVKjYzo7VoEZ/n
JFZqAU8bB6a9J8M7i0LQ15Qv+ICdvb5vgpaSuzEjwSTaoU/sfkT51u1xf2Zl6h30X9OPyY9ZX/Ya
QMhECQB1TKUPgLhwwJinm/yeHJhw+nT1eUfW2+k5G41ecx49i2Wd6wVCD10N8gHLSBP8wxRwCEKy
6TX3/8Fm7gLecqcm/sog4CcdkwJ95zfcZg6Yc0E4jHPi0o7J+d5AhVu0exTkaysnL7wDjRuPr4Ra
gCXnVKC35szlyVwOyBKMB48dV2K4g9h1TFjt69ShIGpOYLef5NojcYBJ95tSWlbkKr0FdugPzKc8
1Ixp+bQ+cKHbWNf0uwY9yb3xAZUM8dW+SPOQvYg0YFGBPOZTp+0KJuTA5cw8jYWKNVaJBBgTQ+Gl
6eutb2oVAgmNIng6pAro7yRmrzlwUdwzLpDczS3xWG69uoUuV5ZoLJnqDXwG/aza/pgNBA05jP/r
4KX9JAAgwTuEVgO3sM3uKODDgEj3yeI/pt2o/sceSMX9G3ua0yXvZQys/eU1cXKXiq75zCw6dFVZ
9ewa86IfjbNmZcEJSI62yfqmWGq7+mt3r0SvhcKL9sS3PZGC0d4BRO/eOeRK6/CrDht1ZhTcwWF8
AtZ5+UXBqs6zWn2PNw3uBhdikzYg/hzrRmtn93xyykEIPMMxpb1dCdKjhbiAiUcPaSRAjgQJUNoR
KQzuRQ+Q6Qe3TMKRtAyIgsBCtHj78Ghc3uyrCFIs1rlPJRSfm5yd1jmUOaNJMBj/h+Y6hsw4LmFs
kMgM3Dcn9CrvuyKv57edCN+TO89b3DIvyGQn/CefJGEyxrKQXGPyvIRx/lTw91G4M+3HyFZWIUCy
YU5N7As8xBPl2qV2g3EF9C09krF7xhUPP6qRNfiuytn9Wdnmkj6xMC+oS2v9iXRxst+L87AfGKVe
BWJxPsSv+df5BATskVpsN3LgXFQlD+7XN9UPO4MqIMyzcjpNi84bTLhEF+KHZlH/uvrxSQv0a5w8
XKgWwLFmYbuIlkf1f+K7LoDNIF9hwxzIwLQ8ByC94afeqsBnHtkcOM/k9E9MZIZ5JojaHUM0LtDu
6mR9fmFlLwoj7lgPEqkVpkUa6HcDe1fuacC///B7vax+qd14P8UKBS7WclSBMXyuK35giXbgRzuD
iJnl/hWMyxETxJOABIYTwnKgydXHwYP2Ze1CYwoXgQbKIX1yMMOwh48H/seF9d1aDN/z4ksF7OqZ
f7p0ZtMOO/xXOMZ9stXNxpHa5XoA6x1Mkwh2dqsDqY/pcpSia+84CpGINl+jRy66oxSamrrpN19R
I4wgYkP5xNq5DAr9ruwpIbSC6M0KdPUusYWE8b5TS7334K1OAuQ1RcNzBz13I2xQ/QSkllc0AI3w
U/A2BhKAk0WQx35GLSkzuOMEAvs+jBrHRHb/iOzMH2Czl37gWTtquW9LBm6ovZMl4xECYeZZWIBj
xpPl6gVrZYc0Ilf7YKCt3f3f1Rn/iykKLk476RlnDroxBzNV77MGU6h6TL4/zC4suPw4VUA5G3pO
n+FgJFqdCKdTWyqU1E2VVUSkr3wzNwsflEqw7Ya9wlDlOpjhpd1+7VfnHmrGPn2nZJ4tgjiTM2G2
jZ4Ebz9uu5tVTV2vEDAH5bxmprRaOIwihf0cYyzv1t2fowBTGuyaWZaZy1qQeRb6GTIEtjK+CMeM
kQspyDZYYLvIm99F/2nua+7M9T3HwFFsm0E2KEgCIzBmQyoOh65RGfNdB761N2+06RfHiLZpArEb
HFdN+83WH4tGhMEQDuCR8EFyur8rqYZqVX8q+0FvjqT/K7N7g+b40+rNVR22Fhjo7zDjDCeSxAWK
7KDu0iguY9Eq3UZh4X92kobB2lBAXZmF4d8JzggPsCWj3i/fMSpUwNUoiWPgzcoOFzwZ4zBmDUpH
+DxPu9A/ViPYus874uhpvVdrfXYNWeUsCgKhjE+0iZ8Vdw2uXewmooq1mRQyWUAtubQAGYFdzCbX
DRygclf8L/RYsp9ql6HUJWo6JlNOoMNNRQV6Ri3zXBcm+xlk/TGhB6T1b4/8/OGA0gTPR//+tiyE
7SKn5ehhcgbM6rZbHTQkz3fvGJDYlG34H9zppFY935tgLgzRcIHwW+SIPuY6NwKA7HKN7FIEqdhM
eb3u4e/nEEQ5VYgZE8zC+Fx5FtrMtM23etPBUW0KNRPVYvlevFw20Y+5EIHjfEJaSzF7RkjZJR4l
K6jP8lP1RzYvmfTWsTqg3WVhlA3hQdASJe38KWJ6YGKsOdEpXNeEDz+iRmDtpqQrc3BSjA5QlEon
5AX+QVAfDTPx63WxYKN1upUQ2sSAwTMK4rk79W+Xx0IyNwJT9J18E2lv4mOcC09VZHfZkwU1hBME
2juoc+X08e4xGE4eLCWjju/iWFbJt1sKDewe1eIYsRRjJoTu1Jl96bX1BUUKxvTwDxie68c9N9dd
7XwWjmJMHeN2ywT8/zLJJrM/eRPX3VeQz9k7Ya+oNy0Z8Y8pOY94xTdU+Uw2JtQb/NCHeFtjNPm8
11nbwtRbN90hcBVVnrp8+C5FZqjHpMM7nkDBD0imEITc+0xx3jfNYfIwHoBTezT2YGMzd+4Pgz6Y
CY+ROJ7RWV4gZ3KlaEZ87a9rAGTX9DFEAw7KFUEbMUvZfgTUn8ecy/UxKiuTuTf7ebd4ncokWhLL
RPBrTLlZ+ukBbehxY8nunvrTdnHkUP025e/OhFz03L9TTvC3pySZncsmC+83Iz4cufHwJvIo8Izi
HguCZv+7litG1EmXrrMpyorPWCKtxR1GDhyaNQ8oZeCVUJIIl0IaqKf951fYuagTu3opw19M4mrt
YhWwXYyK0A6I1U/GsElquvLrAb35c3uXlXFrTlE4RIO0CIgFseDbgm73Ms0KoNWlN35AKupDeatx
5cdIf7exkLKidYTEUN0tPA3moE+us4Bu6aFqgEXbKDq9lRIgQSCO38pSPFGgyT/U66vQfcOy9VUb
FqAh+xm2/n2IKnwJWQwfE65UeMtKFtgBEKYpoZUxYVOKP2qSb1uA0c38U7SK7CCWUYj5uThE+jEA
72WiTq5xlk+M+CGh4tlCpjJmLaRDpGQy96hGXuy+mdmoJo2E/UXFtWfojHh6PjVz8l4r2nApo7Vz
SXmGZZ+Zzj4OBjKRr853xYGijD8nGCHvQqO0vN0OjjLKTd8gBIdvH5FE2OG5fpWwNS68PlkuhXXE
ao2YqXCGpg1U+RKB5r5me9kdEvjJSQlLZqzTGwJRz4OlAcRqZsBnMd+sWcYwRrkkqIAWcxVsdeT0
9R3xN8PH0jsXeJUml4B3SubiNuzyVJEI5zlh5m1I/pHUFPR0GUB6F6f0FMAHLycYgdbqutVZTejR
EF3MmtbC7lRFvqKsFgr7XytJ5eMHbnekvqJ4i2LiTiU3AFaSSxojl8GwooyfIx2VMlavd24B1C8p
3icNwIXuxWA8JmHmm59sVS/6R/0pXcua2U4mEX81ihZRj2PB8NbYBs4hcK8OPqkSxjY6wULjk1zh
/1L0yXkBE+gitjM8Nwesl510SvUEJGht+nnCItXtpto1f/mlDj0Yuf/v7ZHEvYV7zlVJVA08LCjO
IN3cEGxK1mwgyivXcD9HDi0gpgzJvl4kFt4ckStMDqckxacmR29kOYKNCj6HEzhVo1Cmla9XKQxJ
z8bhm4q1XAdej09yEWhUuap9vgi9AuZpu+iZNJeeHmZDVWe9/FJkzE7fNJHS4L0lvTdaK7bsc2aD
U/W6mgJLjCTQ0wUt2hzmX3/2olLcJeKvQ1hPoR+VPJSfmXU1lFtRC/pRBAeqx7KLLCxELyUnPeg6
C5V+PULklBAww8iBmwzH9ZKQ8gN5deEDp7WuUaR3N7daMuJ6XBP+mQfNze9a7p+aNGgNbjY9p6ov
3itBQHAG+CziRcy4WdmWs098eZnq6CrHES0RK6eXQfsg6EVM6f+ljeLvqOxbD6pln0p5LxFPcGbW
1mYSDC/UyTq8xMD6As5zecsbIT/+IYTybcprUOSdV2eLfHI3tt524dKYVz7Pg7yjclya146611cd
JQZTbOfqP54g3HoJ54+6kEkNSWagoKQURVIICg5zt/NZIOW6gtV8g//OJoRy50mJnbGvH/c6FXGz
5YTvxEII+xIjKjC/Zy64JduHUcFkJ4ESq6X1xGbpwxRXEN2sBbG0+5mt+xLXur/JRiXUMisfCxCT
9ZUysJ/CptZe6VQtnfM6o6Pz4lqJuiUcQVZY/TZgQtogPZVw+DB5Dr1QKL2C/92kjVPwlFAmT5v0
XB/Fmva247NpRTDmwaWFpy865v/m3WVterx+ad+Z2jgijt50vAdYIzyQseMcmAU+FEvUVDkerlpL
NsfsKYwVJ1VWJ6T735LKDIBfheDifHeiUNoC095HmHedSDbWZSKOwny69s023LoyBOQOkwkst6qN
79HbtceNC+yie/9igwhLXf3T+mguPmWck96ce+SsRyXEQeWTVHB3om3Jed91FjOTXvHJubpHTAf8
Fx51j3viBSUuWr6zSem6ow44RCcshL1dm1DbDbGC371Jx4PgCv9jwvCd3ca4y9ELy6Las6zSiBWG
niWpmrln4tVWlezZR9VUQtEZE9RDgvsk6+pvwMBM/HjA6tmBEFts9xK1twbBI8gvCMZEvyd27n3r
2a8kg+8DLy6cwnrKgaFE6TIMmv7OiqxFj8+XjSsbb+KjB70UUGnKgeqP7LVsJyZUZWIQfhEuSs3f
hkQI8KdvtoXr1arBNachDl7PIrQURvfqjVAIZVAf1Aa4cHqesc35fwXLgqH+b842p/5Gbv0shiNg
z73fxEddjoy5N+mQAIkPETVeK2XC1PIpnxAYQQkjAlbo3nc6M7gXJj+GituCW7/0GeAqqhwFVxdQ
NATY/k/C7q9OUnCaZYxnhw0B3S05Jwkv/Y3QQe6kVq+76LjVbyJltbdbNt43P3aeqke5dnUxDGW8
Ew4KhnIGWKmfDDmLlMWBSZEwctiTJhzSZsMsi9NVV2T47y/CUrFNr6hWQnv0c0CvgsU24QRPV6F9
ySIBGsQjnwgDap7LQF7tZeGffi5ZubdzrQRFV1swz6kliltdmT3hTWNEckzwrmFrF7eVELrwcuFS
p3nAbO+nR1iVZ+SOiHDWW36t9JOpwIpWcuaew3ZFKbUk4qtdXp3vcUZqqheHsgrlMFKcL3vWi1MA
UyMVzWQu49iKYbA2IObXY8KWYXqe6wgX/1OLrWdDqVHL3IamkF+NYrFw9KCMSXdJEc0rI8XRGltP
Ezjrl6fEEm7BBnqaTO/zuGNMthT9yBxYEOjSgrAGpXxjJyJUCMM2eGYxDtQKBJ2T7FkCbRMJjS9X
fng/Gu2OvcdXMHioitDJs3GA6IDRMEFb5kYaUV0e4LEAuqGnn3LXze2OzWXH/f6KZbPvYfK4aMwL
QwYod/ePgK6tDbAZjgrYibCWZ3k6gQrHgbqDuL69Z6Krqpf36H9LMPWq3S9BcAviGAaFYd/mEH76
q6/J4/PLATKxUZLCFMVn8wRTZA52zNVjuDwrwes1Q0WSFRr6/QBH58U8immyOkJ3vantCqtJczHN
uDJrylWTj6fnCLaOdtflrZbEsF05H7XLJYh+E8GnxLjmZXM8ZUt8k/3vxDsjmq7RY1w/xRvVNqjH
ke6PHE3pnWJRZo0I7BHmqHa52fz+Wd8oJofkqpnhKBc0vP5vzrJy8uqlLpF/LF7UCa56S7ZcSfVf
yqFjU3+AOqqehUVlyJepRskY3sMsMnKCSuQcJ/XtZntsT/POfW1SQ+/pzOpKpNS9vwneL7gU/kXs
W3o3YmR6i8PWpKhtsPSMOb9Gm3bFQWVSncJ2Iy3C0mG77b2UPc0OMe3k1M0s4oWP2wdvcXQgrTQy
Yrp3eFwrW7bLKrYYP/pH1fvJyuUUxty5h49vGzE0uAtNLclcx95apYSDK+KnY6RLpJZCzS4BFSCG
rSp3gk3+czqtfvrpeLi5wyYHMvWW9/l1xN/P66fROs1TuqcUQwHqJTCr9r4LH94bIzyl7VrOoehq
amx/EPPB1vqimUqjGCjD4LsvXqCFALZ5b+u8QdITX5qvahoa/Rvqz3/UhHl5LxMt7Sf9r8PzWgEC
eoHrJ7eBQRLrOl/o+/LeoLGaZ7vdKesL2PiG11WtkWXnU4egZbx/PTWX9g0Hyb4o8WzU5RcW6vn/
z2NXi4awwVDqFKz3kJ3mHJfs9RqfhZsG0SIRO/fRvNIQKV+1EMUekiYyGxs9FLvb3KoicPclORUp
IXco9DlkuGNyG2oRAoPtkfz+PLJc/npwKG99AzsWe5dicaEIgHN6QPwi+cXKf2ltpWbquuiBQjWI
we5SRooaB0w5hRSx+tvI/ysQF9tOspNu0TJ402sQNcTO1t+2y/cp0wPSPc/O1FgoCiVc8hj//yBD
iPolQPxfnz+o1Ayu4VJLWO7fmi/rYakTqjKvgZviT/kXQAnvKkk7+pJiURE6K74y+YThnZTWas6t
hkXkVNg4/m5HzSEerYrQ7YS8hCtB1+NlECnjRHe0rh/+lYO2mkH80546UI1SGtgFZlONYQMOAcn8
Pqy5xA/pFkeWV9nmfcrXhsWEv8QoJ/zViwnzEAOdCpM/ZyE/fLu41kRedIfoRKGaAyMu0kZXZJ59
ryGpNv2vHHnWYBkzkp5XDddSzwkotB+hNYZ06Bs7u+CJq+pmgzj3ozAsR+OFQ3iRPRfhYsJbP0Ko
kNy/yahX6aHHF+SUKAdh4NTanw8EXLF1JrKm64q133+MXr5y3RdT2Q/IWFnxmgCNN264kVTeEw0b
t2fB3muHzq9rvWe7k7gWnazns3suXEJvRo167OPwS5zrt2c6jzyj6tEkJG5kzLGR5qczvgWNiTNN
ufbOwom8VHFDwuHsRdK2k8bvcDgrlwrJP9VI2Mtg17Kq9b+vIbmsq07/HxUVaE0BgkFz/57MwZm/
DNT6kNbeBZmSbbDtDu1JQp/xDGQ5/3BTcxUiITHFEgF2WMaixlc8km0FVHRfzvTcmLuEP0ZkLm5l
P0y04KVIn7sLov6ZxrANL1PT0OmkNt/bo6cxcMOMC18wn/+bA+MbjcMiCHyxb+DH+ig+kgBp8IQz
ZDaF5fSMuRn836okoNuONhVhKtHuYsDI0IlhWV6tez18WNQlxDWJiED2X2UIvhcIU+1sqkR6TGww
x5I0qr4n9pzqxtdzlg0MCdeqyP44TTMEDKy+wcfbyyru/hqxKhMOCCbQj8IBKe0pam+NfVU7s3kI
/8jH8yguxAK45s1ellWdWaLRfF60SZVAvtt0rP3mW/8VXs8iICe/5QrtvK9ddtCi/JxzNl83fgBD
2wmbqNjqSGG/K0Kp070K/39QJp/yQbRTD+vKMGd+rSAmoSCPRHztrW0Bpx5MvPFLEZM2ok6bAyOW
3WVsivFY3VVs+SsQcPxITP9ctL/9JNpElRoo8wSCGgpAo+nEZhIK5onnLItgO+iP0HkfitkdOJAY
trVFAnmEIMp77yM9LR4ezGTcTKHMPku0Q2MTmzXYe/Z8pOKCtHt9Q/852hTlXHtozKhUkvtfdqyX
p2W45UxZnWcwoD4Kb0YaXI18y+WM/bsUw8UsMtlXuIOwGJ+5TwHKURjyYZV1GvtWh0MWKIfigzPT
V1KPw+ZeixORTzp7tZaH5AJ6VZDQKCKyxgmjuu4sYuKCnsT6ZDiKDPaTo0OGOMeF4uhltM9YEvH6
cof3WW0SRx+PPy3Z5C33tQGJ6UBxf8pDqba+X/6fgWgrYRUCRa1HkTMGIieo62uRdfgSsQXAj+el
4qzQJOp2Azap3LwRjqiROWP4Ksxa1YurZVriHYD0+Kyt3IssT1iB4dywmJY49r3nDgMawhfN4kOO
PQIBBLo20z5GahMlj6N2HpxMJ0VHDfYKdhRvLlY88TrA2NBs6DWHdb+fcg4KD+HFikNq5DgF+Z+t
R0u2gzkEiBsCzJj+oPigCgbYtB98l4y9GZdHxpTn+jbY5aheug7EVlwn5IAwdKqlIDCt01p9hyU5
xZpOjlNe9kp8R8Fqq+9tUbvij8R370/DmlUGmkqmPPpf37/OMqTuLXyKeGS989a86SZGynwWBcJF
aJxPbHgnAIkgle2nqnTACHUAz8Xst84yQDYaFkjMm+ezg5awaDJPzLmTPQyU0nCpuydErAskXmnW
eUZKiMPHomAIgAZDa+ai62ODGYy4KiNNPdnfuYq5kYG5Ysg4Yks9NWDgi9BxWrzRRvsvxlfO9A7N
SsPBTZVObdxKpp79xOoKAO9/PMm3x68Gg/xUxYuUnkjCQjs8RZvJTf61WEC2c2qtrd61flSE0bXg
veu1oOzSsypMZWyZNOMyFj5BIUZRL3vPPwE1FyISQ3e8m+JLco6/n2XRYRfJQxlQo1RfuqdbIvlC
nxPuUMN8OzBn3IPkTyD4P0pKELTLLIAApSbAFyfWjs7hJIfwZbr7P6/q390MI0bGJ5uuAWoNinY7
MoaE46pDQEIAL9VMBn8uve451tRQkJjJEDboK2T8UZJrsAwZhImSKwaMPX9BWdm8Kv4HugeGQgjw
deHYe4+sVg63Epm40Pht1JsW05im0c0bT4Dq17Mryvk4Dk2GGcQXGi/3jT8mM2Fpjjg9x+VpYYJ5
B3EAMS9/oUhXi8Veh4XpHEKzpbMlNIz/BvIenv4QnrjfTlC+OpQKXXGG8E+m6Px+7GTJ1jRMXoRH
Kd2PvJkcWK4SQGjHK+mRUpj7LuMDBwKO1ZoXQM77ahA//2IpZkb7Pndm67JcqlpeIJo3PDkW72FH
A9AQbibOzeEf3U7rRkla/FvGQT4fYZgAyNhkR9SAMoBOpEunOYYni4O/iPPvoRHo8J/8gNfl6VT6
gylJfceMSFbQoMCWLj9QMxQrgiYB7hcYQ8gH4MTmvkWdXPyDTJy7DvnWGmbGuJ5S+lyuKfgZoUIy
bN0Y0dCLKMr90wg+shESkJsZGLYAgLV60hg8GmgSr62WxUm6ajFLTpO0seI7MsbiiI6YRN0sGLMg
A/WPgcHVOVzpEF8UwYMTXJS5dt4qNZv2Q+Qb+/7R7uUid+i11X4l0ZUVx8s1w7i+SCbOTeS+iE34
M6qmMuc5fO2gsnnQrCuwj/VUp1AcO7sif4tAYt1rqKB70gsyl5X/av6v1qHOgjyxsD+3+dAn8tbu
gKH9G/ODt1TWYOpV0E+76WZQQ205BAMRZqTNmEzYWmK2PKoFzlxh33HethfUvxSlNKUDPhz8sqKD
i4TbhBIlfwpN6oxTMvripR2WNip4vCGdTe1Uu3tMVw/N3ZgLzX7fdm0+MiszQwV1k0gJ653p8beo
Ev5QKx9DO9KzcvaAs2VPZWJzjhPFkSVWvDzxusnpko1Cjy+1oyNd/AX9HFOIH97zR/72W4soR3s+
Lf+euHm8pDQhfVO1wEmzLtj2ObB70OUxoAugj+h5pO/GTuG4TbiR/2VoCWSNRkD+/GvKRKi3z++S
e/HcoeQ4OieBwSXXuP+q51tKa+wYO42SDs3hFx8W0wAPBttPkfd+D1ItOaRV5rQ0Hr8OU9mejeO+
ercvStDtXs1QCbFm+w0GGBkqu1j7wcqD8+CADk3dDtEyV/8fyEv3IOaUkWlSdPLPsfXRG9jpo7uT
JP1FRBrPXwgAD4uHqhYOvPofddvHHrSVqPCBqhjI/JrmgbQs5hRKIr+O4HsqzHpQIWVVuswgFm3Q
xsox5Zlo+HROzS+/sBCtcQqIucoVZSKTAeSmXoNChIPsEptKTU7TLpqvgokgd3VGUxomiIkFHxEZ
mDsgcZosjnMxqyx3gjGLgyPHOUenRQRnJN6YLTdlQN2l0KkL/n+NPzGc7DfqEWuiXs5nN0VbGtqA
uVbrp37h5IGs3i5l56GcU5r4rpheJxZXdMhxV6wbfA4hqRg+1RMx5xcm41o+EdR2Tg1sTiUSpnJQ
2YvgjtWM3Eys3dFoGmkvetACJA++0mUzPR2CTQ77d0iFF3oJqAEtX3/ibAlozrioFN9sppr8wArq
Fooc0Uh/nDg6k/oPhyjr2u91AmnWF5e7bvmQbo1dFlKuvZ5mj2WvIyPbq45f70tIlQSBqDcYuYza
935ksUFY4DEIeTr/aSD/UorR7F5wcSGon4ebXXoMit9m9in9NFbIXGdajdsnQKoCeLeMiwKLKc2x
eyQHxL1wQItyc0oQ3+FpGWBU2jrc/WiTl97iW7n+NgQPGue2oLxuhZiVi90PbHm+lnJDh/AcbxQO
kgXypMRlAA3j9TYlKjePvXRKiCF12i8yjDyzzcF5QDsFCL0pXoh/WkP53KrKDqjBkjcu24z2hMn+
livL8zEOeuB2GnNPXe7VNwZBTYFi2U4o4oPud2xWNT63RA/oc/2wywI6BtFJV3RNyibNexFArgQn
pifyZAcUCnAwoYWTYVFQDnZ40zV8H5Nz8NHLElNf6y3vL+pIwrjcrEsOmkbsjxVZu0x5GH3hGbLF
dljsX0va2J6D1F50XazOrViwG5B/tlOesD5wlj7LRwYlLuKZD0OFRquUjNXZDzWku9F/2lQguWTK
8sfcQRR0LrwZfhtw5tlxZfnWLbm3mi2hAmRXEeJTVwFSZ9kGkRHo6JKpoVfuMc+RYu3bEOoN2q2y
3VWeoqIfT9QfjySOPxStjj/S1nH085KDsKPDrqgzCL2tmwcLkTFxVXfjdKxxqMYAAGfFw2ve5gVe
aOK/ewJohCSQOGmThcCHMwyZF1qgVHoqS2H3f+vAjy3dWE7Qt5N7AHBVytFtqkKCxVjM1FSzAnJi
cPRssJW8OW2WOjT0JpxjaGXkauLUYnImW5dO9LTvZqIA+24oNSFmIQq43WchcN+hE6gN7ilVdfQs
tHtifuPNUprqhSUpsFwmuqVm8x22keCh8vKwmt1k1/M7MdKDW60+ET1DRb4OjygVpR5MMIJoF6Go
knegWh8bVjrKI45A2GnhpIgQEWf76nQysnZ30CqLLuzHQmW8RIldWFC4CkrvZc7VB6YigOimMv54
EbS34+lCj+KV+w6awMityLNVr5rqfgCdXoW2V7kjIKRqIBi6+ZVndmARyddMK5fRRzhcY4Z6hM5k
yM9nA1ffTPvxxSQk6eWqDTGzg6eNvkwDYSYYcezBPBCAR/KDyJ6ete8h5+qAzyXZxZHYW9uDybwO
4lGrBV+sL6jQb7G/zHW3dbR+7GU6R+qcGm1WbQtmUztOvY+xKmp/zl8LixveReMNzOmFJj34Uj4m
aonLlqQDtjKcB7F9Dmlbm5uvPYznDJHDNlljIh0QfFSmE24bMAFUGuz2HDya1sVogOd9ij5NS1Tg
lXzuPDiYHBLq01NZIyrL8Rcyjvjd3xUAODFSwovB4AO59BI3QmpBIisrn8sA8ONnoOYNFgU3bJq+
HOMao6G5gj7eSrxZQTiZMLuSlA/l9iGgPPtIeUqNoHCDPT+r3UNNWgE9b5J4RAM0j3mTw9jrlHER
p8No28PUou2bHHeoC3QsmIGPaAwQoBkJxLjnPmZWik5B9aSbsCeIfagrV+mUdOeAhpZncclIVg1R
1l00UM+f4iTF6hhX0NWLF83OR2OGl+OvkDqc35030xkBtRujFAqPWC8X8eXsvjqgjNxAuc7T3sqm
FKs2ncl2p1nmqLWlVBeyp5eLn55MCU4nqQCEKNaD7/4NlMY8zLhlKkeJzCDlj/1qCXPMBskFjDbA
IAuh5pxrcBI8CCxb+WppEoCsvV5gPE7PM5ngp+T11GfVDTsDlUa/W8G0PVfwRvVIdFtES9pObMTA
hcBIA8eSDg6PBAmnltNyUPZJ0lu7EyquiPFcprzb/+hj4rHGTxHANMENgrOG8ac/NKhpdZZZMSlF
w72Hwe68hiOZ64GOQ+bFjtONgUUq9cdyeGEYRr6E4R618Tj+QvfLDrDLS2WZ5RKp0UAI72WQ6kgu
xDdVagFWoabALmt0nM5XmqigjsZvbMSAjevzVtDMqaYidBS8WtJyQK6j0ci6RYa6T564ayDN7t3X
QWWRG9M1qNZdG+BiSHivZmXs8tEjsVHRvFTlXC7fr5VUv0gcQoTUsKxFGsSUpCnzp3DhaLT4pMNi
aV/AmFkXl37SeFHC3YU9eyYBBxfuR7ATl2w19HWKm/C8ecMpnb98+98eWieM+SXFgVlCHE1Tup6h
+pREMOL2wY+7zLKUv7qS74x/Kz49ajYDqBU+EGMXH2/mBD4fKfxxQHfPFe3jdKoe9+OWL2GfnTzm
jHWyscrINTzBGw3cRxi9yfx1b38kXKnXkTfypqwn07SqZ17Uuarh5KaXMggj5zG/DALccC6vxuYG
Avj6fuaTAbS5YDzAYUYhYR4TzQ350HG3BiZ6fCk5UyHqhlTSnYOStM7xe9X+mY7KSCxLNJdt4CT7
RlDwKAqIbd7Xb6uAgpLF+ZGCogMFkT7bJEP4u7N8+eILgZ/EbQUk0UoqlRuet4EUE4ydafmbiJfG
uDCvyzCEAJsS2fdKZilUE9pA4mXbH4escAui6CJ43k35rdmUfwXI6VBLC16PUGOi7/mROeaB0PQZ
hzkbXW1iyUXn4yq9n1i1UfsHHZNqHQaBCwGc1zxKR1Pl4jufZhoxKViBwnS9dM9+YHOAfyBG2rFY
t6gZxGT0lJ8u7d5nFKjhQSkJkBi266va4mE2eTMCjLCV9thL7PxBJEpYihphdoWBkvNVHHAN51WC
Q8ruWm2ATLxj0294kgqBLdbnoGbi+dhI8lNMStkkHWWoHYnZooeSljkyvJWlAym6DjKGGzo0AXFe
Ew3RJSHGPqnJCL/5qqPSAJZbxbEIX1lDLgA4JFv2fcEAYH30Pe+sXl15FaNeb4Wg9QQ0SGjVpby+
djcQNyJv0/knBu0xgTDuZEijP38MPv/FSlQAsQmAGnOowQu0hEz9JcCtEFJr+soiportq8Xx3OEV
murRoxwI+kyvrE3wiTUl4v++MRRJgMseUC8S3NucjdjDEaIoybSKhc2V0X1jsDCOkqNPReH6JHwI
/Dpy59Rm++tzG8tQO+27yVyz3VYZTm3U+bHzgWhVCgU4txb2kR1vANxYJor/0GQYeVkb0aHgUS7o
EQd1iH8ehzxk4ouZ0Ag970CbDKbiR7TCoGYiV9p71zAuMloQ3reAmCIdGCSGw926NER69NP0giJE
D9JsCr5sB+RmKtmuDVsUoYzWXysWMCSAwQYzjxlabIMgMDea9DOS+LZ3s80YNmajcuaPbHnCeA3g
pUNZrAstYAqEg0aFBEIqmR2mV2OVBUt6MRFkTiRSldacGKGuGbSJOESb7ZYVCRg89pts9JAci3bE
+Ku3x0GvzrHd65mkQW19ws4z2v6bgQ8/NQPyZKai/FoSd+cz87S12656fE7U/XC2q3TQzc8ukssf
6VgDnp+lYQC9NaQVOccvRqoZcMz4M9oH07K1fPSQrP1RmI0DBBHtpbXXoA0kPo1iyYPevM2Q/56n
AwhOqAUuok5smUvB+Nv2fO4P3owOJuWVFZaObCiQgHEJRGahI+U+mtKMruqImin9MukiOgU8dcgj
/QT7YSQNIDhFe5jpnTmVdNVyf/fcnOO8BvGjhtQFsLqbGueS57LAYKU5WFp2ftoXzToJKDgPuGMl
Rx9+D1Vzfljydu28DWoeNIw6iCDL3v2MrCONiyQneVbITwfr1QZiuT93mmGeE1q3M8zxKlrRMlwD
AiNfpz0IBK/PXDrLGrxIwmutsxuSG9dNbVt+61tdEmc7D66owVJ/d9rX/3BrolYx8AJKe82ua4GS
+bMvIoLe2nYZHQsrQvUTETYOwCd00y669PItb7aTjUidJkd6y0ciugm6NkM8aKDahBcCGPlv/1DP
3j4EUIyHmVVTwyYmsrwKtHj+JFm92UnyRkxYBNADOl82OkdrQjxPOFTdPHWNcWYmh0T0MCwnaT3j
+UCclsMEEuuPcpp6AaLj81XP3jcw8bUeosKSuemjDmniqPslvhspIqdWD9e/b+liMiCdu25takUj
nk+N0tlopqFsScCKnJRCkGQSd+Z6i5TDzs6PHnS3YJmbTA2UusJtzxtlwI2b2ytwrNQusxgogjgI
8MFqjKrJa+ds8kXK6X9/fkOA8nH8O517DDFfwEFa4wPUSYUPsiKpgbI3JqhI20gpDBwUq6kXq7Hn
0mPHexBxWVFFkrOzZEby19FoFzI3W1tSMOKaReNIcDGHob1oJCLL1kJSxRBncgrGzzJZhtZAj3cY
TfivXVyvsz+hiVy4hNLy7+BuIwkTy1eVyVxh2cxt3yBrOvgLMiFA5R59LMt8HxRr3ELYhiLEGddi
PHeE//aR8tvqHDDQfrz7F/Yrn4D6r3HRAEdgEBT2YgdFGBePtynLfjox+7CHuld1YIF6cNA7ej5d
ZUhUKvSpsEs1rrunloECLKobr4g5ihD+aR7xksFovass4V8wybE/sj54Ur6RhCPUxp1uG8Lp1lX+
F/YT9vHRnFNmFZclISWQ+TapSq2MHjyLo160klpP0YR5evda3l8iwMb5pbIJV5Pzk9IIvWqbADV6
vJMThMMTwwW1CvH3Vl9Ns7zir4SFqaaOx6JoUtu68yDgswENMzHsUQOgURkx6qDiABRKmI658x1I
NJmYi4f3DS1QywQtmDEIS6QIv//4Mti2SGJR7021ZVUEBOG0EQIQP5T+CYgn53c/f3H2oLdIS9lD
696N5u+rRCLmC88J6dFZKbQMWI5fYMoho6adTKl0x6fzD7flXMRwjAXsFh0FbDWr1ub0N/7sY9+l
qLC9cOqi3nJlR7eM7AJ+Yji6M0KBD/DqK4qDpz7hkKiz0U5FZCULpyT4AscFtiRWE6GIhzoQ0zcg
WA81pN8YQMvwhT7VquCGBvDAofbNlHnR6jK0v4GHLmq7WZOrSN0tHrcyFPk8tIlAtscaJF8Zxvp1
Bh8WhcdlcW6AUOsrELBT6IIewxuVhu7rOdoXPy1GerdniizHQ2lwOQuSNP6uxq1PwJtbgSJ1HIW4
w5ur8n+071YseWtg2srcTwL28ew/+buof6Rk+2PTowzPdoiaR0zfgMcHWpuudsiYPhM4x/CUZD3+
7VZWhnxlUyRgyUzfoFIPTP6GWmTVXAZdhIIqNny48Mu/+rMXM4imXMpHRR5LH7DAjFXTVCvR52o7
L8oi+DdxxlNnO5bUkeQgKtklv0YPT5YDNZC7Bdva4QprssHiP9emU1K3EC6nC4e2MrYqNAIEjMJk
43cF8b4poWfNT17kqy0rnFoOfEucNKylOCGEcJaxzqktSq0I2WY8H5lu1l36AW81Ik/yivpfjlD3
QZ4H5LiahKBnmWfJFKHq+Llg1Y7P9ygcAj4TE2ImQcGnTjhrPwzp8U4rXwLmSSgNIVeqObXbl74v
SEXfdCVix400TiGc7RLQ+32i7u6kwlGeOlf/luh5Wu2RB/Kn8RdmJLn+84xui3veUeRlukE4FA7a
CrFduGOzKFVgqV1THK2k1U0uI4MEvdVNAnm6lpSZTLBHqsaSkN1Csr+XSgYmXOFB4hz4gKEJN9/E
OK2vgoWMG3cp3z3D1MhmB7Yd6rjLi3Wc9GTsVHKHTiYnLatu7LcAWiteM7VvE2It3xtW83G7GHky
EGRpQMU3eHUp5lR2e+Uz2SNTAPAR38BFCx0wv6wfFnBRzsvcsymeF1deI03FnYWKD7q43pe+Jh6j
wtKXY3+D+Yl09ijk5f/p4WfoWiflHdS2V5HEJa95JeLavDExmTuSmu1U8ASyfbbwM5n8nDbFL55m
8HYfXMg+XbFKG4ION3NDJMnRsoyC8V3DP1P+L5wLdGpG9DMKDAzAGxQiEEClx8a6VVi9SvQPfq7F
aBxo9H4s34pC2bXJh7Zfou+1YOvVpUgakyJdPj8Z+xIfV7My4RC5DnwCgswvvAOUlchDy5u3sEHr
eViPGEVEgVTRUCJPg682aZWD4fVgObREuTo7NyiPfQFFKw1Dxcy/jbRPMbKq/KnK5Xmm0B73NMcA
ji8xP/4nKHyDsoCA96YzOfmuaarc4+hDJqPO/FBbVd4Jgkcxx0GJYP5A4lLVOR9ghQ2GYNtqK88V
8zr0DBf+f3xWHOJ4uZVMWO1W8cXSYXjksn2GFt712jzDFt/TsaAHZzsq53thgrW9ACEehRcxAWaO
QZTT55YhRbpelRuD5q0QhJ3YNSHhkimDHdYjWK+34TXDlFt0ckD6p9QhJRqgRAmm//IckJdCyRNn
UvHITwoQmXJgoA301+fB8egmkMPGBacV5NuK3wcow3WLE7L50fC1Iv1HJg0vMAi7QtqAMtbLM7EG
aHkzALRqpjoUq0+Y0+0BzCp3t+DA+fJrVIfpPX/qW2zH8wWZzdvKZuxrwNCcaE/53U7joMbelQ48
HTLSNBDShNC0sQ9yN4ChLPCArXbOjXnA03r3y4ZeBOENl+y14fNxox9S9BLSoQllo6KyGPvuPf46
bEHknCp3ApY6hsdD4wwnArxPlLKSqBwi6cpwIBeCI3z/hzXV8evBHBnYYq/pBc/3MkEI8q9YNqnT
QrPFSXEoWes6SSi/B8vNazc68xbh3YkHbcYn0mSIOa6LiKAPyzXdRRGJUYwacwpDr504+LWDPGXC
p4wIlqrK8rTRInQyU54bPrnXD9EqT4d9oommmemLagqp9mcn+pEMtKMbUAcsb9o9GF3EXemEGQUw
ZRU5h3MTySw/G39F8hQozjkIcB3T0B+hzVkmO/glS2sOCCDQfvBO4TI1bC/CqNjmvYlYNKfX+u14
KvvXEdK7dHmH21q+T00XzC13FqUZ54J2fcHgjw0GX8Uh7U39agMHsJu90z51PAvk9d/Z2AFb7aqw
mMqr5bckUC12c8q30abVnbyPd7+zjU+LtVqliUpXPBsb8RkFY4XSO/mv8ls4gZLPvLwpQk+TXqxu
CSVScoCecmzmhA4mZZl9E/+w1HLoL4Qq9MXI475wd0pJy6EXaMTAw43AUXwQl9N4+uhTTmlRarxo
7H9EnjTTqUwaFTOZB7oKPKLhNxQ2YpLmQ5FFtpoBdIdnyKbv1jgcG78GDk/0ycErMp5luMLh3dyw
Qj+6u5uuFna+1zGKISZDlPKOT5+7Zrt+eTYkAbHkqhhUhQki6sJtSULf9qc4St6W3pLyFUClR98F
r/FbPxpT0JaIZJFITtXxWkLB8dLT4MiKiBeZphbpfnHGa4w1IVdk6+tynYoaaHn0pS7hQK06nqkt
Vbr8W7SOQQI8t0cAAnwkKAUNUQU49ZNK3P+lDY1/2Z77NCFj5jAlDpF1OWCbMjsya8+TdQ0MlPIx
9FGT2bauxoJnw0ZXbgaNWy4OJh07jn4wTBUW8EgcxvdnYJL8yO2hlw00001AgOGmaP8KOSTrGAAy
7ROyvuode5yMdiqjSHWpqC4e+MTyuEUPQBcJ1dihVcfv6ZwOIdZoBXPGrhyqMVG7E5rLYEjYruco
rEliZdlGR6w5B0xRmMrQ/Kic6vgdY1/W+P+su965ZcasiyGQpwyJmpmlE1DIwnOsI/EpDGseuS7d
QtzDWEGxTOfRrwdokTeOjrBdxtIrIFSqufyB4BpMz9drjwxW5Q/JlEjF4SfxQf3k/dqmm5AQ3Yow
cZ+zWonALx1UrclyyBuZF8/6FURtyCkvPcSqdL9t1sHobLkdSKD4/63IcJqWXy+X1U8xurNaMqTl
61zB2pFPT9SejWr9aODZRW0/FUDoLb45BOpfEmpo9DKy+kzjscUH097JbFbJ+fngGSeJcNHgDRej
dnbC6tf5fsoe6vaCp0+2J/xCn2fGwFTaOYACMzeUtpTSHhhUaNWXTl6ELwdfUw4eZUNxVL3H3WR8
tzp53/rmHu8a+sb6beCQSp90bW/rct4joIqCoqtaZSJcz14M5QAIqZHADZ6OsX1Lm7mGBQ8DgjSs
NzpZVF01mqkosOR4HrdQMweSjOB1yybA6DDs6DAzFBtngioJHvFLTRQ9hmRhCJhwjeLVxP4PRPi6
bBa+nMl8GnCSQajk+gk4sCmuU8YsrJ6jbKj8VijRYRSXm2iBq2VG7TwLy445h26fFqFVe1ibbXp4
S8Z8XvOvqoAE21vM0XBJMHYsYFrp15MzWOqD/bDJvR0YHDPQABLb3aS5K/IuNrYpY3uM6i+aoM95
QCvzmT9ZyV2L8TN7r4eB+fVAJw7K3E8Z5p1IhoqLrqxw6lKrBxo6Vf9VeRGvTtOgprbN0IRo8sm3
k78yFwns2/BH0Z3FeZP8losbHliO+eiAdf/2YUwdGwoyT5IjtISLLM4Dif6dVL/Du/873x/ii/KT
0hBHaKYmHwVD90h0B2n58KsDkeIn+aDST9KexRGrNyojDaLrSNz9RqlJ7ms8Y3tK/5KOx/3KVadh
acnTCL9fW3+4VxCe8i11xcAG4/+l26Xam0RzreLWh+Wu/DiW5ZZm9WGnag54GQyauAWHFQl2IsH7
YAV03XBxzS5LJX9JucfFGfF9HSTrmMvdyhxdVEAS8krEXTiNIp/dJglN4Wdd9K3rdNXY0g5amU9S
96SmtlqVT3HjPvyaxWjVCSKvlQE2FcpbwUHEAuotKpiaJCiNuRnjSwFYmwHXo6S2lqAKBC5WRlC/
jC58JnuR5JQ8YuCxUDcaYWzh5CDE6B+d2aleDrVfW3pncVZN6iZimyK/PSDcRGdieVSXVKuvbKWM
TqwaUfujzkLDL+liOqKlCDbYdsEtRTlugQLMT2Wmx39eXe21yYTDC73w+WQm3KaEp6Y8rw1xlJc8
TyG3cHym4iykzidrZEUA0jZcW5vfSMLnXNWRAJx+uHIT5TVS2AYKciji2SqH60grZYc6S+yRbOBu
5RHP0u1uSavW1D1EOydG7zPIE5eWHfEEhDstL+pkp6cPIdngkAfuxW+I+E64YP1Q3q4EtoCEf5kx
YmXPuoiv/QE7dBtfquDduIw/Ojo1+tlrQ22z/P6arUKp8fVj3OHQd/YsvD4b2O8soNPitVRKr4gY
IPgQ+ghqL1O8cbaG24tXNEp4+Bh803nSbd3TMKzELeyp1KfcbVHyYS+YLTSPVORZM8eji6quBrpS
nFSWooMkB4QFyfeVTXXYpOBOt79+YMoJzFT1FlM2dySujWjqienCk0ik77QN4Lt78p8eUHaazsMW
MiEuWeCYhNaJwI/EvGqILmCUSU7D4WfkBscZ9/BZeiUNscZnyTqZNLgAZJbjTTU+A4cpuwWpN9SD
m8YJK7dd3C67ZwmH4aQTnWvCbo1OTHxvPLn7qB4cELXy8PNETErq42aMO3NNj84iiToHZ87W1EBu
J4wKMiPgNAQNok57DnFQAufB/4fZ1cI2JtVinVJmWvnpAZm1452KIqbZnms9i+uwOmrpCFtEH6Ip
DOotahJoU7tfJjFCXZZ7Ilqi1Ucr3R8nAYVdv4T6ZA6++H9ggsY+RtL0ed3AcOp0KDQDfQm5WOFz
zc8Ntf33cvTrarfKhyDqFwIWeSt/rBk+A1aMN/5nO2HSXaB7wfIdN0CVAHmtN0yMJvr3yJW9mPE+
bj4AOBl17SCojlft6euKFXDhMNmNs02JO1BE2hWiBAFY2misu+OcfJemhAW8V1SLGwcqDrWxYpob
xPUxEqFfp7kQbZk/ElzZnwnnFv4pXOo5xgvPwDmCFs+evArNgEXmhSMmO/sUz6uUi5wCSe+d1KQk
rTkVYpQbqa8Ar4Je0p5BtlkPW2Xk6JcM9pJlrvBn1iHltXal/UXgh8DumQZjVrEfWLF22QZbnLHC
VOxwbIdY//mMpQ/fQxmDco8IeAHCdGiOhe5DgX3Y6NVdZeapSnpvyZ9mLBKZdIcTONuWfEFOboDH
QWetJVq/QmdxEtvY9xXBRGDQe7vU324mCxK/7yhIoOFBBTe0OxrccO+b1AIrlxs6XXntaMFJjBZ7
JZ4bk5rE8B2/mryKdy32XcIDPcmIntmJFJB4fmWcc/ZWUvraja3q7qgSed+KKl7AMKI4tyEprsSI
yopn7wtfBbj6UPeZOxObvTf46p/0sZxyQH0gys+gqbvCAhYwpDJ3BOLcLNp38zPmQkY/2qO/rNkV
nHKFzqstkRb8WKpGEVFQ3Zi6ZTZCTBX3cD8nWh7qr8s03uQbgy7zBzyFjVpi3RKz080dSarPklyP
Xygzzgga0b4QrAC2qUdLs6BqQUVwWuRSWIShIWSLfklvPkrR4b/Gc3/R+N4gZ54P/5ppl8M2f+H8
SI8csIspUCvtwyO+IJT5sBjlhv3wfurKb2WTRmSZ/G3D7QPIkrE0IG9aY8eaoRBu78MDy9AnorIN
4z2xBMh7pM5biL5g1doWGvkxxD8mmal705QVGLXOCkqGVHu1xFhJUGKHfVWIO4Jde4Th1rSETjzZ
UnJ3pOeOd5j5FLJZTWopxFsGJPwFX3bvjSTp0WS6taq+gL36XUJDvMn8xofg8INE0p2jV/3QOWHP
8aBdmEIvYKes66B0IVVXRSyVUpiu/Ce88uZBCmoBsw7fcSltCkF++Lr3hL8jSdEW6lAJxpS7I52i
VHbG8JiOjSoM2JT47t0rHFQUEZ63P6dIjHA+fQQK8t7sYWpWSwkQLZFKpFxRUfEx+soZrTzaaKhc
HjSpIESJmvpg1McmH6/ytbyuyVBKMppN+N+CtvaBKs3YPIN9lbfxhsxSaiw+6vLReMlXmRLO6RzY
Yvg061In0plum3mreiLnIetBapJaQLkzc5cFPm2Jm5YPgakX0mmT2IKNvfOsXKM5UtkX2qkpa7Bn
eyDvEyVC31y1ZJjKDjymseRn0zkqcae/emRi0vOJYtcEdsOteJXWkrrN6X4+0O6P4UcE6KjHY6O7
u7eVu0pD2aFwRfe+Ts88QeJTsLDMVZgYmJOjLc7kEtiPj4eOdVA/+YYkapO/MowYYUkKjIY4F3mB
F+k6Z5EU8Xa7on54ca+6o0J4f5IJMSntEBj71Z/ySqK/v7ayyF66yB1QNq1UngkqJo4T9K8b3cIz
a/AqjrbOvwM3QR3MXQb7kiiNlmx8vijzm88BN6kAFYgCGIWp4ddqrodbijIufAOzxxfxawsZHybS
mJFDm0E/rc2MDTpXEtswuoSYNV9IXWckgeinKtdbLkXqkgfwLVM/cDKRknhcKAjZoeJ0QtJdkWEh
njmW0//qNLO5Ffj2jyIl6reEDVKSsH8OdEbgkJbDhyM6T3N6MTndFYfFynv5IBy+Wk4IhSx6ub4l
7QFontYSBTnXqsTmssbMH5pKXiHPZft95ftvoLnmDmRAscOTMVDeUHqFvAglfBB5ZXNBqqkEujcv
nYxOQpzyUeSe2y0NpNBa6B5NUnorOO/BZqKfASNonx8U5JjOmahQPiQJaTXDiMQHLm32fJz+2xXr
a4kK8x6wSBb/DKC2OeLD/kAYoMhvsh/T0WWBcEKeqmHDU75NQA4nErgf5W536ws+1ncLhGQCFwt9
md1g6XPdXj8cPd10X8iJoB+GYdwfR0PJYPnN+OZkl235CBDigGkWRLq2z5Hrdcaqpt7J9iFSqpsu
QVtkYTmS27QkkN1OVZB0vbh6YjPJnDZE9Pgg2TwlpxxYkNFfjhMC0ZD4FvbSiNNptiloEzBdHm+7
QZXfKwtkb5XSoMLo9IGeTTl51qRb3xNk//oF+kuU5WQRqCzPJPk9C5eIiOWU40yPqG2wArBb4b6p
zC1lWY3qgnMyjw/KQlJX9NvFFxyqVIU2wwjTJbfN8pVJifRGdmM2x5qi2dDsFs9hTN9X5Ob1jImL
Y+m+8KffVeHlq5NPjNjoocDAMtDR8LZXdn9SQBtTyrSsr8de9aO0WnbgLt3qZkysx7T5c8Jzc6WR
WiljMFGx2vEtJYkW6hyMWkCsytTeNS/EXB9OZaMNOeMZai88QwW0LHJDiYJGfPO/nsQSPwYWNvtJ
0KcHytAdGCQg4IHOcvcC6LiQMo8/EqHujKf45Kw7duNW2/sRDTzbE45PKJb9Ok1fS1lwSXEm7t3t
bn5ubc64c2ys53k7U/dOczpn+0ZgiBOZCsIeb9v1BDbe1N50KPXvJKiwl5EHqkQOjuhjBTcBhw3L
uY7duIEWZQjeQx9NI8SEukGkVJbRWXVn1eCUuuxoGwwDphX6K/H0Rh5CtbhxY1JcsCB5YnEtJaIJ
49lWGctRFKQuBd22tw6/R2BbfoFMiAavevBq/s/mbEXxkMRHc20gZUB0GKxI63LbEUSclcJSdWIT
CZsb4EMF4jr19oDn3P4G8uomBqxqh7EMrijKuwO/P/m+z2EMyAmJbUo3Fi5rW41RWbNIe8D8EpfG
uUKP/55/3gCZCS4yhOX2kFwHBZijliMitS61nuW5oIpi4NmWo3HzfU/W5hKmmuck3S/dx4woQe+j
lJiKN/gunQdc/H2XK6jtuuFCcwV6oXDyIoJP+IxRxngpf26Ht5f15pziR4O6rn/ybHBScYmuRVfq
w3zb9g7bx7FKyEudgQLtKXaC306yB6CoDkwLjVUq8hnwpIpLADNnAAHvcd5Ow7fHxPhX5YUDOTrh
fWwRgmDRDcMNFD90aD3/8q/Gi1p8eRVvurFsStdASflDwM79JkvlbJMuOPpA9zc4a4E9Da7ZEnFz
tBo4LD4sCKDZzH7hNPr8vYecKYCcryOoavxu0NlZoDc8wIl8y8m7leYD8Y6tJzyBWkWRl2yKJsBg
OXvO0JJwrLd0w32CA1qfwWL3/TOsZ8uD1jr9TYaObIYEhRQVaeFjuQgAFmRUxA5rKLy8fVDh5xzw
49rx6z8fdzI0+JKWyfp1M1eggjZ3/MIJECxTYI35ZKM9i3tCb2tMG1yeVo5lv0xy3oSYoXvUGQSb
H7W1hFh8AxNDgHBHzqAuA6kb1Dai7I6UvEEZsnfuRGwn2Q7bc74G3H/KXa4uYLPK2r7GnpCKZBiw
zZI/wYDW2BPYz2ou1qH9vsBMw2C0pG+AO+l4Cw/IPkSro0mfQG1zfeBt4bw+8I2MANtKIfeT+czv
h+bqvFIkFjYkoKZJXfZbOoPovSJNZFpVpgUX0JqcXIz4pnYEQCDQQ7lrwelBS4FoFNiVeYAuczu6
BLXkHRBhwoRRPEYZXiB24r7pvC+nUIhyVeWNNs6MdtXWabS7+JwOQ/YaO7n+3EW6QasUB5Z9Ug5d
5KSl6JBvCU7YlHiuGgE3zh1+JqOXFMfBinYtVQRjFeZMZFEtHcYu/xrKFZIyKJn01YWeQYMcBIHw
YW2tGDmKLpNKs9aboX6LPsKHW5mzedCbv0dCGkVgH/OOqeaXjYtNitNunQL+xAO3TzAooWag7+Qx
ptzFRbC35b/Z5dEKOh23HJPeaqJ8K2wMx97Dc+9XSxTbgLx5OV+zk44dgu51n9gY+fOTE9tZURmJ
RLoyrHasOcdNzvujDlcuG5CVhOks4fHPmAfAbK+b7BA0zijX07nFsbEvu+AjH8mVrqhNUPl3zkVY
wBuxDflwe78kuRPYKrydyRD915ZUbGAcZQ+m6weQpWDkF2IyndNkrDERzP7Ehtl6Wr+Atx0qayrC
sswBaYwp2Miv3XIMLlj7v3UxlYVubf3od10jNxjK7hLGYM7+htRnbug4ieXnM7GIeJyUGQhrSmmf
k6ocPmYJSiDFcUUnbFibGhj4hgEvJLJCObmJ+7jNJSs5iaa9bU7FgbgAwgtv9Qs7AiG74VQtWNu9
24CDWNz0cMrOcJbKIWF/u/CCG2Zdt9266oH82qN0Fdhps1o9qkzs1EZO8LeNDg/93Hf7QAdN7sFP
YGrdC/YD/Z8HPtR71O7/LpfiT6WpI1/g1wUL7LYftFwVy1h2Tg4iSiP43r6BtRkgxPSPsXus1+HL
ZShAwyRoKHVOt7qwz5S/14TAmcH22x9sT3QP+VZkELTYcqWveojY8KLbIgEEr8yIJ3ERX2V67NRm
H0HY23FZLTJ9C685LNHdk21g82vaEYIG0NzSvsiUmWdru44OEk40WdjwZVfWPdxIwdOwY29Ivsau
616oO4X7qn8g/4IjJRRgzMmkQfFJ53SUoLSBWDHQAYoN6nY3++DsX5H1pj/CAUsmLMJV15JZWGIR
gCyA/k7dwrP1fpDwk4Vm6IX5rGpolj7TsXhe3IYMVz+gSSkZRhmLvV4GLgGlzPhm6DwDJQJym5CE
UP8l5xtOGajCqbLxxjPSyjk+Ept3f9CTsAfo3y+/M3EqW22jHfdySyNWw1ugl8Nr7YxSdsAyVRbw
1HXhwu4vCPcjjUTdHhe1bW0B7xJZq0I9lLeFiy/z9Kwxe2XDVRL9IMH+/NNyKwqXK6/0mLLYEYEm
2EBdrt/XhjZXkiviq4h5TGLijK9uHdz0xFMdAdJzmquIF0Y9qOvLDj2cJBmV9sTcvg+7+zYsFUGT
nIudEhc6iniZgCgVkkxKSObx4b4vG+hCqBPLiaNFSELv8qMn5mA+gf/fGqB8ahUYJ/OiX0ba+2/9
AuhtUkB8I04vxYLBCxf0NhBjnTHp3UWF3+r9vyYf147/toUQK7ENwjd4AZB1pAKvzjFQqLAVh+Aa
HYbHtdon4THEzSHXazYoBQC7Iy9Bbf8/mvFPOj6V+8sF09XWKI0mMhE5CFp/O3Z1qh4A3vO6s/yZ
H1z7YEJL+dz88Y2F81cLbizwAKJs9AsX3hy9KqbeN1F7MD/U8FglEyCNyZ1B2x/nylce+BlBYTah
5TsbbPtPSW0jOr8cjqgRxe3BWd2qwrhyXcupkAzXDP3nFwxJg71NzTDc6TQ2G49q2KGdjlIsxFNN
70L+xZfXoowyb+79slWV7OB13rXtzLhqFJpJe3XjoNYuPMLIhJab3KwZ05QcMrFzV8DBCNyaKTl4
CwLK3KZn3GCJKfC2oG8zCt32+K2fO/C6LCI13so65pymEy95ZVG7GLDw1yQ6TTafxTbUdGL/0bra
p//QZOzMXygyP3kalGVzibqaJqRLx7IBb+g+f/doxWTqMgsieTZbz3WUiRiLMaTzwsPPUJlkpHVe
WcKW2+HVOTSNsHaSxOnm+8JRYv76sc2WsK7hTzYruP8eoRunPrd1O/OiMl0w1QAUcteLYzeZquIi
FUY6Vr8WVjU/fIdxJQNQeE7BzJtgyK4cylj0xIU0jB2a6mSILFN/KP1yJ8zGWt9sbAdmK+VMrvuG
k9vcKgzSMZozNfhlu6bZDAkcezuC+qvy2bMKTgp4KKCADwt80BYBM761dZNfuEQPA0G5hVF47SSZ
LTsNw4AeIKsL1oiGu0/i+2Rvuq7hxfJf7odj2n+coLUmKM7tFwFPTZicQ3NgMFo9LYRv2DtemIVQ
/o/WaPGZbylw7+xkHK/njqPs+qCltZkSv2WfvDduONDZZyqWuJ8nSo2UbZyTTrad3P158NJwNRwo
sKYE5FyuApKfqceFNUKNYd21DhPu/OO3L1M0H+x2Ov9PP42AODhdQL5xGpSi21L/iNJHaYWxm0d4
jgle8PIb0Fr+LF5fIgLSXtTs5qQrVmGnVU+YGiTnAp4NQe1HaXi9fIta3xvPPrQeYpzIBc0nU9gT
14+DLq1X9zkJnZ0kzSggwvNMCQg4ClMh3vRh2kYg7IX3h8RzVbhYGKx/R1hY4p75b9Mz6Ev29yjQ
zawlJ1dwublApHNMaIfjgGKQoWhXd2HT4Kbr08/pFvMzms+A/isKjuxNjHVoUUq+FTrWHmpTU+8B
PyernJRJMXe/cUZZUt34m0PDZ7LByHD6WyY++RuCRbVaqNzPe3vMOAflO4+v4V95P9lep0ru9tgX
OP8XWhMwA8sT4WMlRn8dHR9fLHLWSoh1BksglCzKVq/dGuVUEhUIREMxu0DG74GJNYcMG4zYoiEA
44wnzp8x+sUhJvxyZLwKUHrHhSuA78SmoUwHLifiC8BHMDvhH1/ihHnL/tYIMyYZID1j8VWo5b5L
ucVObCQc2kAEc/7P9XResO2A6PKfLZNi1TA1gke3frMI3wpci5Dx+LapfWjKyBOrsRAqoT2j+pXY
c0MwPAezDXw5tJhliy8ysTu+uVG5nr7cPrTBge5cjsCSffaqdxtLQaEAGoNoGEw9uc9axM2EBRIl
ondWMQVVtpgW3CzLDHNo2zuKyYrR77q+Z9qyapncmzlitJsw8QKtmkSOfcrwuZXbnzVN/bntwTg3
SfiWoXh5dKJv2/H7s7AKt2ocSowEKp2ezVvoTyjA4OGhKosjNyih2XSZAMG4+6aI+ij/Ua6OaOf/
K9rBRF+HOJLCRZhQPdNb1b40785pI9IqqI0euyyAvJR4TkLFFBp3CJmUE2zG8GDTVt6Hqw3ASo0z
ZYXlqOx9dIwLi1WOBLMMkhQUkkGZ0OhY3A3wzp7sdtMvZabc69IgD9LHH97jjfUuHafnGtG2VHpj
SO8TvXvbRQwaGWoMeLODdvZmSHd48C1uPPM8WbzJyGut/nPdhVArDB7+pH3zx6MR35BxccpBobVa
x2X7IMW4wgDFjke3RwJNSTb7jIOPf5u5xqmw9tNZF/gGqErKxRLHDGYuwG6+OgHVrOSTb5JHxutT
8Mhb0OIezmoYm1OsIwnYSQnt0sQAx2x3srYk39U0Q9BTGgYjw92Kwijd/E/y0tM8GBx/6x1OWHes
7fa0k8acthZ1mJ+PrzIDDgzfKO2QPENMmLZFY+IOivIGvBjFLyznNjay5BTmCUs/KIojcuQGyX2n
RqyP4D2OKoU9qYVZuqoPtD0HvDvozGVGHXR8HPdxuhDCQkDHWVH5wamvejeJWly3Ja+Zds6d1rMw
QwQmOyJbUDcxm45yZE+2NUoEImkVkMOR34Wm3U6GMNLSDNaQRgcw/5AKRc+Nzie4vAyZmmOdhBgB
nvzZPKWPs0Wezy6LKBCPsoch4zAwGpujul/wpYAUwz+DoT0bF6UjcTlZbgdD4EyIHK/duczOwvzc
SZu8Yk+Yoq2yUBIomcop4JBZr5u79zZRHIha+q9iOZkzk+8ssfTsSHvNATnJ3/d/d31mwlQxM5z4
kigW8K7Tbq8UjOIFagr4mHo/YorEsWfsBLRwQ/4W9eW/JiQW9xTr+kQNz9y/pCGBn6bY1xP1qB1o
5txNu7EKYJLBed+iam+DwSlP49YVfuSPZNQ/XyyAf4zLQPoEmQ+PQvfc1Fsu0jAU/I5uIzd/uk3S
mvt3bPQA+VnqGClSok4UJOvVG9d32vK8lzftZqbpktcEWxT0H6t8NDoms66vAKrxFNRqjM9LxiG4
fPYdw1z+qGzBC+iNN9e9vOvaI1OFv/i6a4Gr4N6PD/tO1wRBMvach/9QirEqe9XrjmiF1O8ghGR0
haB1IeUREfxL1Me75h2mV9wsfai+qYNFPjWzF8ElEPiwkvvNs1fcZlohHqlJ97RA8VXv3GCAV78+
M2UBwCNIRW7M9WUm7LHHOSwlVSRBWGTv23OAs4t2yKYVTVAXVlvt9LDJ2BcvPrlD+frGLlYXjtZ+
OME0nFgXjQYa6s+y2bGtKgwdChUexgkej/g4G9nkPwC18/pLdW8VINgjTXwoozT5iLL7vZGeR4p6
NgeBsyNWoynfY54V1dsLPx1pJ1sfCpW6y0Lf+kucrvNMLL0gR8zPM8jSVGe/PtK43hodlfc/jK/g
rxJjRnvp8LMX5cy35qeXJjwiBZND6WP3fzTWbkTYYSVmOphgphjbFQkDsYC+zIT4kLJJX+bvcO04
umr6c3EJfx4B4UxQpkUiJy/h41GV97kDP1JfxLBsIsYgMnn6hFXJ0P6TetRBARvE9/lmubUdaPW4
swN86IJJwdWcAqWZc0OvKwvbLqthO8OuVE2Dl48rM9ozToNubwkx4my8LmrzY5vhb17Mdb3+wEe8
DVScmDeftibRaZS1VPn3QfLxeO02Vv9KQbKJO8ohM0GCs4Uw1OUwbKMatS3DaKzSj4M1I3e0YWfi
46cCg+Q0zEJgmvmaaxQwoYdG09mSRgCSo1GDGXZrc0mJcmOb6uCFTTTXYQPGwR1/HGYw8CP9YgpD
0Z2tDkAal5gmprX7dUi7zjj1YZwD3bsLQLhjpIc2jmRD0srKHNExmkJOMD9G7Iz1poZKmztA3n4B
746Fv2kxaZL7m21Kzfc+ARU+1yxttWIePBLhz8Sus70s+Zfxiydw76fRMKS5lG5ffZBBAguotX1j
aQPYGKqf8JH9jJ6PUvJHWOD4IxwBOIz+sHj5OIIw0zdpHLnAoTkkLeM3d5XYyrYzaNJsaxUuOY8N
zU6zAWk/Jr9WPCpt6Xif3FPkN6FicrqKyPggni4FZn2zCoQl83XhiX4I0d0vo/Ztxq710LBKdvQ5
h62Qr7UNSVl7wSllf4BizT5mJjeQ+EnoBYg8+4S4UQ+B8rV+OsDiLvdbu2D27YF7VsRE4hXfoj+B
qYDCrpGplgWfvSFLCIfmJS09iBkRGK8srXDKljinLONn0XNEXukOADOn767H1BYuk4fwM1XorZwJ
ttkpL1S1wATrvKM8wvgtGDun1HUpMvZnER6Vrf2tFprORO+CPrxoKRoY5SQhPk6rp+EhJpB6G7a2
pxoZX32TsCy1C6eCO0b5zFIe7dKBhQuGtZvfIqm4LuDh3yfmGZ2LfjYXKJflO8Mu+va9YqoldUcr
AlYYdnOsM6jpM+vqlh2BHtRSitM188Wr1c/crbhXASX/XbQnBUnbdcMnkI3lUm7CKsLFMGfcnLpj
vVLbIkOemQWmOUyVGHwe/65DkJyZ2p6cYT5WZtS0fFZbDTZB1HXtHRVabf3mcR00lnjXLsu/8CzY
cfUXSTA3E8I6tT3H7cUibaOZyQjgghvfny1KbxMFZOiJ594DsURwqycTJfO0/iHnyvR+GRldHMxi
UAGnbiG5ljh44osJncfBSpQ2pfZHZ/FXu2IxyQJwnWO51Rpg81BT4gggJ4GX+KoP5i/0ZJievpU/
9HW3/t2yYZcgKE9luhFWIS33J1nkaM+KzqN+ile4/tJyUR5lBrtidENkHUMpWJt8gZmEfEIM1Ra0
bTN4qavABI/nbbaIjki8t0deCMM96VLfSqKfwg2jHnxaTfqZavcmxmAu1CHquaJBR1pXFoIK0ZcS
vqlH9AkTWbnOz/GGqVQKZwYJTOinYrVButS3rB7gMg+2GFuN29VTRMFJn75WlpPg6mJWq99gEwsZ
NEkHP/3Ezg59BQDV0FU/hXYhuA0IF2K9RICnV+BiBGZVP9heAQjH3s/eUepFuQoNIgYob9XfiQ92
55RU/UC9qr+idCLVyI4fOuO281y6L3K9sPVrTQafJIaeddsRWn8PzttN8d1KzTlse3dmBBojloPZ
zQ5CnrVQkTWUD8HbRVusGrGN8r2DApZaoO7wrY5MbnTFTe/NX8pb/JAjCuGPLXkazEfiY2olckN4
UMcEd0G8qVj7pXoyAsgfk2iHoKESho8+vMhD6fz1dez0i/OqggjZmwkC6XAXxUpnXbDDdFEguUg0
VmVwJp2Z4Y9r6NUH0DZn1QR26hdhvwyHUC2dRedIQzO2HYtn/Th7MjtSEesmQVBw8IiUOv7n8cxi
oU2GarTuwWpsvlcJL7tMZtugqqBfigxOcstpdHaIFM3PDEz7Xkdv8NLzwBlVVnHBGmjw0N2G5ZNd
j1iZKz5SieBOBBe9XQdsTDoW7OwiJq45l/X2JA1DcEFLdZty5ndjKiFH5zJR1IstfiTc4vByeMz9
08MFt5P2tfieSIJ+biaeoJxG/sCFm/I/bim8JZ7V0/dONQ1EEQEV7UcIjUhaV9yk7Q+itrGcV0Y3
Yoy+bFo72nlCKZcNqLFZl4oMFg28EqhMEQxXEHwIpf5aKDobv6QhYMjYESJQQfSMFSh+620WQsNx
v83HdFjEbFRM7WZHrHQUBxC0yR9MlT7+/BTcq2ft5Q5rowVYBdGyI+YJlkBZpoj5977rq30N5+J+
U76qwEC+zgGkckmrwNLgcz1bX83aaZoeGhhEw3GYzJYAHJbGrtv+EWeajbLUG7fG8gUwxpo2JzXo
nS/SWGa1ZNkCviHvoZ5urqPdxGXHvzaX47kNjRQQ5REggV72wF9YmRwVrGgNya9wXI25bmhc1WI6
w4xXp8YzEdh6yTeBoJnp2ce7Xje1Yi4JUpV7Wdxrs8XwVXmUuQBVsgQjv/IuKGD7EIp61jsGnXPa
+jF7FgxHt3n19b9IKWZ5d6WSaeuNjDCSrMducFzJMtWXgJM14qcxKeRbk3UER/UfQfEdIELoykAu
xzoy39DBHHR+Izb2HEM/VCnooxclZGQc0t/MKQi31mTfSgWqSixrIAnkBY2UyQWZInGr5qXYMCWR
AkWPrrzjGMEOOXyg72BcVbzna9u/+FpTjDBJb8lGAInuc9sHCH0ayjnggI2e75+duvBUaMgAjEFA
ZXmS+KA/XNIsyMa60qKHxmrb7t+rV5lD65A7690H/KV7ILTGtZSOqEukjJlRx1bQxV8KIUJWod35
SQyu1BFRjLmfS/iQMtXGR3iQXsdeKJFZKltNum+wTZo2d7aL9AWGztnqOb2EtVocrWoYoMScMHRW
wl4j9SrYXsJQi3qWT0LTZd6CT1PWW/KJ2YVm4Awh/dgamAZFR3dkQqh9M6trAycIDSGDBX1TyQTX
nZMaKhbPBB2yG3Outyc2u0Sj+jgvdR5UpYHPncBjfP9TuSWOJyVxCwWgRpcjQ4HL8h9wKytJojg7
Ccdsq6VvOk+KME9T7sGaNq/azHHDg9XMkVF8nQh6uTMB4eFdpdIZ//QSJCsjQKUg45cCEhUF+Cbk
N2Yz7YNYATtHj37/GfpkJoM/cucX2AEmVUslDz4kbpPeTEiDNKdf5f4oryUQ4iRH42Hm5rhkEO/z
0i+TUFYgNFWe892TAHUPHtStgkOpbPY5+KhJqtoDoiTnaSC4NXI9o9c6zqQBygoTN68UP7+kuI6T
F+6/TZ+yvOdQVdcQ3YaDvTDhx0dsm1xFBoDNUxIx2CI4OR6pNjUy4VPbcW+tqH74xLrYnXX7VaGO
R8KNIQAUuTb0arzkdRGh3xDOCBmiAEbcQ0SPodUQkGPrQTLiegW7Lptx2YxggM9bkECG8ch4gMK7
kJNvZS32cXoNuL0hGd3HOv5jat2CYT13Zfedn2Je1ePr2EZhbEWR3xUSXaj4HNelaQkoX56NaX+b
YHl0TgBMgR5+T0yNYy5K0OCAfhbE368P2ucB+hFnvXT1njB0vZtEdZFD56pWK67DQOT4LW/pECGc
vonmiTRTu0aXBm6EC8+C8Ku+2KYXujsR13Pg/23HOksnr5CNqaNzdeLStTVjSARSgcQ0HL2Q0wjB
mcA1NCN6RWc7eO9Yb8Nk9GUKr5Eo7TBejfRIdtm0Ph65SlTDzlR8YLXBEuZL0ro+96ObtOk0hAwj
Rhm2mZ5EzidrxKsFDyZdXOJRdwkNUAfjOx7//FcRUB31XZ/AdEgI1THwEsAB3GnHpiVDCAv7kxwd
7RnorbrDC2VhveNLADi48g6L0nQI7MdxtSltTb2a/RToqqp+OprqK5tombK+NXPBKgVPy0D0qrgr
dUJrmDAxzQRs5XLMduRdmW3LMjwd8DbqM5z75IUgpVnG2AgkT93IOC9DDfZLiRPO4QcyiDn8abeX
LUZDpeHOJ89KHaCclROPGXSqe7eBEwN0Yvb96KHoUpCqPFxT+C+SWz2DjRJRWk4/Kj6LtQ1+Y9+F
AV4cdCG6icpKVXImn6r3a1MkoSkiIktul2ZOdHzqRcqE8urNLQfgARkgIOdpgYVWy8VIJFNxtEI6
M6CR6oN2oQWlAhl4+ZysX55d92diFav3BQyScZLTtDyjiIHneJ7+KUTcds+6kHBpThBXCmkamDPo
0XLp3qZaJ+Xy1gQa8Spl9Plunu2t0DZHipzuwN7ro6oM267RpR4gpLI6IRwWAPUvKRMCiUAO5KhR
O5rkOLA/jqaT/wRs2kkoZtsxqlj1ZeGsb31S74iEoDZfVHbvozQPXCqEf0nV5T9tAc7fnBLZWkOA
Ny7fCVYiO04R+JPSvXQjvfo4s5Cb1Nh3JoDDEi3r+WNVGvCnZ0RHzAqAEIp8mMstMI3ybf0bkLFr
KMKNdGn2cGN6hWboaHQnNXcGoaRUkyUgcTLeOrOp8W0+YWfubmHmzsBUBcZkgUTZwQwFOlrZZ4rI
gKsoJVBxbj0ZYJH2IgXnB/7BBt/fYCKRYceVw10d21RyufZmvsao4YyKZa04Y6DZtToBjgfO3f1x
TKjn/Dw1J2R9T+0lRviBPOIQrEKA1y26kJcnI8pfLjWDivWhQ7aH+qqcXIgzCe2r99GNX3fmUySz
G6o2Jb8vXhJEcC1y1xh7xc7UtGTG8UfgF41coTE9Nx7PPI02rPrUd8ZVBQiS971IQLISrghh4OoV
drd5mZTPlIdnGYNJ8lMRhcR5wa6l4Yyzc4EL28fPcoWnzbwM1S2snRkBGB11OBDNjJgbZU9RrsVp
GMdeSHhhW6rulIXcFJhjF1h59nUyWBauciRGMjMgmbFMli+OyJucIzXl+OHETCL2DL63IPR0L3WM
Usw+Sy6NV27LuyhM3jq85pLW5hNgKKhe2TTiLN85sNJpFTYyr5DTZVpLPMfZbwKoHjQUdtURWfzQ
vuIw7rE00moeqhfJV+lkTRvbyNKOBVWKXxIRGslNGCopRavZOldCBU/ZOiJE0LhGeMwdUWYpjLJi
NwUfiXtHO6lyvs8CrxDB7pXmIlCZk0cdkiOvN+giO/oKR+Ohj3I/TEqieSSwywmmE8JWg+wbQDnt
OsSyqH17+Sqly3uVMpI9ecFDQGNrsgLJJXEs/Yx19kHTLmVevRt8c4FhwldEwdzWg+OJ7uRpC0hf
KFQfJSzmGbat4QpiMp8jhSPU+2Ia8P+/U3einW8ES75pF1A+ucNq+Bc0f/sacAq/ICAi+EkgPPJE
enwnlTruehSWovW3oxe/JT1kD543aLW3smKfeTqfKOQ+VSmQo8M5EbPeQ9bzz9WLO7wThhFqwG0N
F49uOp2HAyZC2m46VB5WWCq3LBVzppgmftFekceQBapZOyME1EnbjcDOjjXj9NwnFx5saNrl7TFl
UZjyT9u4tJD7Cc4BWJEEk2Bbdm7uNgKmiIvppofehENaDApqEURi8DG/L+2VmAYbv6b7Mr5ZSQeL
UJXuK7hAcUCXLW0Yrm2/ObzjscUxbeCZnr74l/5U+/tfIiMtUbN8PJ29JTn1ypcrOeaZruutiWf/
/Bb2uEZkxk984aSMSwCC/kns94DkjlTnhyRE8QBfbIF/9ZaBmZGQFkUahkzWNx7nG5EejTmWnINC
9frY49zBJGgp0LZaK3WOpDmmlqn8ny4Q7sd4dZ3koipW+j8ixWU3jekmp4ecAYnWNsXfIaua/sfj
IT/j4yrzn5+r8WYk6WHdsWkOlOPbVtvDVTc/v76CV9ymUnKah3hBR9SUs17mGz/UU2+GUbmGLYEw
h7oia/0ckzH8C3MgNC/Y+8wAQiO61OliSdIzS22Gxmq6bOS2jecELNtsTkdlcx5PW5JTwjcCbHU9
HGygQHPRzb6E5MnaRPpp9FSSEW0sUKV4T20PP7NmO/ltbmAUDBEIzQoPlg4geW4VtGQoVUfcpjxB
4AGKl8ee3+lkHiAec7PHBxfB9/K57J8W0Eg6O8iCyPVSppvP48wTtFv6IrNDwqwMU2LcfPKEfLI/
l7CkI8DDy9NX9MtnQxE+suxag+bq73nyffE1RUFcPPEZsGi6WOSraURVSK+TpauY54DbRH7QcY96
nuO2TXRNfXJXgZYfI6BVAPVD7V4OH2Y0wTkynOkJkyrCXtJ0nOHEtcuyZBU8AzNgkdtm2VOli9YA
DnWBSSalybWlpGLYt8+jHdKC4tSM0tHr1CRPOWguyMSzHWQQcS9ogw7G6NoHuCycJRuTNTPOfCzI
N1sZksXdjQnbjIuGtXgEH9OTNf/vm8ZRzBpIUrLcimyhEFnh6u+5W5QtnkAXgydRuFcOPMWDxKzY
02wmat6gEZS1vR1ozVCRwxUzROxq5V57mFTHp5WUyHtglJVZoUvUgEdiamc8bD+kNtrBPTGv946c
U7jEJBa3rFbZOKHeNr7+AJfk5Mxa0DFYYndsUkbycUaMjx0NHrRQlJQKbXBJhM85cNJ6kgYssoPp
mNk2BeOziULsxjO2wUi2HMEr6tOI2AhFxQYWAY3dhq+fNPjX1dhw+L55E1Vc4pXJsLuH8SdDPCVm
gnrR9v/+z6OQdRpFgUMdxcNcNUIv/dLhnm7XZ6Ibekk7HPwOO/aN+gL5QTa1E29yL2APElc1WBFN
BoyPh/M90CumRQFabbrGV6eIZBtzJsf2Tkw8tEnrT3J6ylWn7qCp5OhNlTeQy+3T+ZPsFkmL1SFx
EMNGBqN0cdfFHUe4fHtCyWFTx0X8nHgEFx2OD+b9tLOtjPSRNeZuNb08pzhicctmkpSWlFKkP/XE
or5DtHO/EISlkeu4u7PplnCf2PylqKFSAgW7iCZuy8iP8/q4lbfCT1wkZV0WMSsrtL8qqjvjYftm
GxM/4TNcM8ZL8PF17xMdvo9GzwMrWk1yPTUSUre1E1xVFu0WLF2EeCcl+8fZ0Do10LZ/QEmLuxqR
C4RUdEZjYcyRXvDLgZLY7VrmYNByHq1o5Cm3HOfsHCE3g8TzqT0dpLOCfAfl4NBtqU8AA6TisJfC
qsV7IQwJNGyTwMJvcOPLlE0lCnuN+LsvFtl0cH1B0CuMLWikBRw8IEhG7f4BNCm4O6Md1ZC+pDEH
e8kz85J4bOS+OB0LydVOGoDmuuP2m70mJc7TbevcKVNyCwLcRD6C9ci5rItjZgJ24UlHGuLTuw4Y
p9hm80gtJ53890ygGDqjv3eivO/SJNBApCAPxY63nBFDwKpxW5rfMkCLetEBiu+hVmXHHUe5gEpJ
Ge/7WQ9+PP+65jMMBlnq1AbhvkuCh0HYgM5LtE1I1/JJD581P9a/cpttoL72iC9bTjtvGL01oRIr
pSQBEXHB8Br+9SmGI8a7tAjmbIsjlETXRX+t/WjbhXqAa/+IPjO8lhUZ6iudclDJNrtp7YaGsABN
CCAnoOBxNdygOub7D9dBsrzJkFvN3lmcLwFgfE8IRj6cTBLuNYDHrDzPcJQzI0vxCbZw6akUMrBA
pK1PZmiWDKC1l5WojLBNR/BCdOAF49kN35KUsgQuGFv3e6BPqQecOvMNqAPAOuNe6AgmBJtToX95
fYhD2UDfZaslNcsFOJK/fab4t+x+loLyELozfRMMt2c3KTuZfwppUZhUcw3REr17vwdJHZbkv9a4
iTmV8lQw//QfDuoJr10+koNAQ6URDjdaomxu7o54aEr4dQo7lnUwuqrwJIAQROPK+/kW8fg6/VVi
ctnw5MW5WW3PTGpUf7Cr2yX9Ap6rcAzfZn7jaQtrkIzQsH73EB8l76JyAYlXj/UIYE8WLTzNwhoo
io8INQiGseiwDZoOyJqy/c3adPTK40tM+rnGYNM8IjuJ7QAUFq3eKcqhPQD+dHfdJ/SI+Sz2BrfA
EKOLrrm44TCjvzMm7A8VdrT5rul6Q6w8X2j6Vjmtu60+Ni920x/1d0lH4JkjEcd/0x8sbn56U7xt
2pRNwBKAsT4enbe/Unp+E5Lz+AfpRk7v7e4ZEwjXZRihlck5nAS4wJQ+paLThSFTewf/3d5iYHtJ
LoNz31V5ZBux5nUyzcwP731mTeEDEEthPgKhQdtsx/h+8u1+nN5VmaCTCr9ZXeMxHz8icrLc7Cu3
wskhxWc0rGx+m8Sb/jcF0x2/G2czUkW4JiAYq47iEDto73JzAhLpdjia8EUEVN4LoZiVQ3qDXCk0
Zgfz8cGlMnOTwcp1T9jQ823WHCK/8pNzDI1pvivJbL50VXcXGsbFyVwoR3P8jJPth2w1w0bLLZ4G
2M1O0Tp2qR/jOR/4i8QkIX3iFVMpnE6IhuFShZXMaGxsVlrvAtAOuuJ9ssDdbym7h7ByB9kU2BbE
03TuKqm2aSnbCu+jFUTVyLDkKQr/nKVcD2Jtyw6DB1qKHa4B5YNRdyZ3lcVJVSnLXe6PsX7vv7Bo
56B4HB5yTNEP3BP0E+k7hfBVRYoL+/PCDVa3pYBwggS30YeGgwCT3roOPI12pms+uZ1+EkQoOcHd
9o9ZrYeB+WbTQzYvr3pCC1nizoPjTen/zktep+VEzhU/MnrPX936ncChWIy4C5P4xzBV2PTCnOfZ
bwaAEnh2tXXW0G5jXF++OjOVtWbc+qSDNjj+kEsihP9E8ykzPsq4dMY1dwDYkI/5fYps7V64RpS6
CLqE6NQSknx6uVEJYAtkWUfu3azn8Aenbyb28yvEkhQGGZcs7WeZpXVm911wXHXgGfgOWXAtxkcO
EiVYMoFRZouXxueSCv8+3wjCbYgOeWxy/Hi5vuqzWBA7oar5mmmRgfhISPmseppcKEQLnaBBgSYq
rHPL9k6ctGZy00SzHi3Dk/hfeGWL7Cepi0bZFy2x6wiE8WaiuOnshLuuTsDigxNOo8RawUfz7PMB
84+uzFn+gLpbNX6Jz/yaKqMvbP0/vELbH4e+PD+esF9mJTGAJRTmeZxTjLbi5M7aVX8BkKtlE0yl
NOc9q5A5R80Kr3aPN15Adcrd/svFKDbe0MqYXfhGiAUkedWKhNRJiGtGdfZ0Hbayibf6NaURbt5o
4t/ww5F3+OKi17bghDmXftTOb6lkFxF/G2HnsUI44meSxmjELLmhvZPb3ex8Fa+QXXQFxg7PYP6g
ts7IkRB5LDMaXmADQ5rJXhs4yJDwJESIQdPxz+llcGrcQnKGdkRjvy6XzSWXhc8Vut+lwA0BaO4U
4E3gTNVOQ5ye15B8hw1vVhPqJeynUVs+dKXjWnsz0UbVj8S0vL/hEt779wgktyCaYrqQI05GfjKB
jcIgcj2Ijqn0VPISJ8+ZCNV6bjOxqMYJRwRykON9YQBEEGBj9IvmAFA5x6XnjRThBnkXUGDzIn4j
Wsi5n0VcCFeagNts+AnKUVJ6dkyZ9jTTwL2SwDwMCdy6JfTemif8dqYyWrSf8800jVQS5Cx/LeR+
dh0GwU2U7iF6QOl93iyJbXaU9sgKY13Dp6AlZGpAebOSnIE+vLvv52jw2IwdtIg54/+fPDDDpYPr
jZBFDIs++Ky5Aw/JIbQfztKOdMhj5etOyERrRT82AxNLABMGngvTxpygEL0Fg3HwVblwxz66h9s+
SYx9wd5PDzmknN0IEZhVZw5HybzoAa76J4o6KwN3YBl6DwFjmz9ZqvcSg1Wasvbb80fdXplncaMD
ELFPUD6hf4ZBKFYoAGXLvS2JtMa0/WIcgZbYkfh8pMzb1h4H9p5lYaADz6uv7ftWvePuoq6FOMC4
8s93HoOwBjL0iyw0TppETVfKlE/l77+yfCWxSpsjs1JH9SFTeHi6TvRjGPwevzwI8jnCwM4OJLge
R7T+rMhjZRPvPEMpUQvVIX01nqFy7HDesgkZAq35Yhnwgjtscnxui77Mt5Zmde5DHlbSbg+uVPgV
S23gqd6ScOypvvD+YXkiuxvTmhAP6HsFFeF6oYnRjO/O/Brby9Gr34hS0cEK9+L+QmrJR02rpoJe
Hg7lZCNvFhGugumUk2kiUi4ZSElltEz0z9nqG+JQxhEZWNJ25hMqvYQ+LP7r8wULDQ21/0nOBNRd
nLUl0lyUkX3zzdUE6l5jFsxd5FyorAgxex87ZYjYjDpwwLIueCuGqfSZTn4vPmQG+eoJFqFFPcMW
I94RNXiPzmQSKpmY6w3qLojtqh8HnnE4Uakc3vhBmZPXtq6pDOAlbDsS288UGTaVXtsg1kPzk0e9
YnwV/eg8/+adnEbW4ScXFZW+Zuho7b6IA8GKyoF9QXScET1Ftuj01/np8NQL4rFyLuye50/VGSUw
VOhosNczhLfEUX7N4zqpaL8Fe9y1/icXJqwg7ncsfMMjDfp4ut7ll5+vKPVR1AbYbwM7M7l7umne
Cc0F3I9z/g1P6u9Aa9bcjJIqibOTUwo09Wg6434Yyem/jJ2q/jr36yqbcLL2GiD/NNkuHKA2aDgu
gU2UTjETOSUAcu6pb/bkGn+TwOnxTM+lfGI6DR/t7Dr7R3iwnlPvcGmLwedwXRdWBPfVgAthMWNN
Rxoq7uP8ay/H8LMlZX8UvCQK7uw3ehcnwsY/Ny0tJfyGQYH5qT51zxwAWXd/vZjA2S6eUTl0oO7j
7magt4SVT+/BeGmBzi69/DRiDGHilAxNxL80ryWVMId+7ryB6qUP3lOvMHMEj8ApzjnPSYWr3tjA
dxPrZB5rnh57MDldGcOVikYnRrNBr/cu3ZWnSfI0UBWX2vrO/3/1d8IuzD+r9y2zObRMcCVz4/iq
64ZroW3N5CmIBNjEDKsVQMvy5/lqktukk4dP+dwsTEabNslWuw7br+6sl9ukVzM66rMmIrxRmddH
QdHdiXZzxUtZ2aslBmTiDxIN5NSNBCX24bC2/jpNmwxie09E84u08IOrM4YphhQRCCukGM2W/WuF
cF90R3UkumHTmw1tMghw1ZxESTmHl5mHkRbE+6eV2F5UBGXALYYdZisTOXnthw221nhKKPwOkvG/
MW+/M2bfgvRigeBk8RSDpam7S+AzrKK1LrBb9HaEN1PjtWYVSLZwsXWjop4me2LAvnc/SuIeR3+A
GKDC8aItHWclV+V5/gbRlyXYksdvZnQgCY5e8IEL4qJnd2A7jX4GDL64O7hm1j8zvrSB0fBaF7dr
bpX5iCUqtmXDSs27jAGR2Y6hghm+Q3FzlPhFZCkvkKtUewHPQEmjd+U4zzs+atW5TVXf9Uzqccgp
1F3txBGph4o5Wr26LLidDSKuH0WdVHSt8Lw8Oae37fISgsy/kRK1OgPNEYbOgSd9g576gFzPrLJS
xoYfBIs5lHujR+uAbzuTjHX74HETguN48ddNY4AoAt1Ta8qyzL4sQdvckB7QXRMjbpae6SUcwwoJ
4IXf5PUunkrA4MVEWeMjoRgBRVIKtRmd5l746BUPCiIlSeyJliq1hfhP+qlUx/uWab3ZIddcMQuk
CZxMU+826BVNAstLlpMsgn7MFt87gs+oeB1GpW/YBYVfe0Z2a4bY+ba1RFVsl3qRXqMuXyKC7Jeq
7NvCYChuRtU8lSK9dUBGc0M8tYLLXpzwvVhIHnAJ9eln8HnZ2DGJwCA/LNy/dMcjezRi6A5n/KT6
albUP0y8++L8SrqG4jztfOlgVhkmQOZNSKXoR7qT5StHTruNUNka2DVdxzYYq1bZqDcd+GXPxlnw
OBP4DmrZIYtKRMAOG0qp/fur36h3NnsxuRmWpzMDCGtv/HTDHLOINfRbW2nBkUP5tCOtBvgtqY+G
nkUdAmbvrrSnq1ClNLyAO1L07oT6pl7hPd8Eu4CUcpZKGVzPrOlp1eSeOrfjivNZby3guMo3zWRs
QylBemMzBBfukKxvGfUcNW8x1PMkhmtUrgXW9qInsJ6LA+3x+dmo7r3+diHv4V059YrEKFVMI2OV
+LgFSSATHwxUZ6Eos2d+b7R+bcun0pzYZHw7AtLuka28Vhx2cYAjIBUZTurqriyhoBQIMAtySfu0
aH8HzhmruUw6Rd07WP/4ZwCILfjHsCxNcjCT9KyzYngjBXNRoXnGUj0eri7/GYIZ00PGn369kCSt
J/Pu2ye/n6mUONuNeeQb5ZQGrHoSA7gLSQWw/+ZMmjM8DNxwzlOoPBtuZo1KO42wdmBX+pPfys+d
kKeutA2bQdIGC8XYqqySYbE7yJrDpQUt7qQRhUAOWtn3/+DzugdOVzQddkkpGXS4Biy0ZnOoSK3a
hMPpluWXSKYd7KtNNcurhZgZf2031F9ExhPibLkAcSN8X2t51tuQovO1cO/tdW6BpAOvYKJE75hy
QlYQE4C5B7IA/xRCr1wYPvTG1kpZ7canGAvpkBW2fZM49uF0k4wp3zAaboBe4zFi0x9erZeXcNYp
3bwUHZH508KZQWAJq1BL69/A7MOMh3y3u9L85UWuiAg9RJf0s/094dMVgdfZcyBoRZMgOgLo+91l
PLBJPNylt7xGrhqZ/kdwFlR+bxf1sBmmzxHflgSiI4N2lffzCjoxn7dSV1P1OfRA4JvtXVPr0VCK
WY8OWEgJzv6LOMHJYW7QzIYx2RozjBGGBp/C8T0j4zWveIXXuf3iK2Yr3lkTJVFVEOOq+0eTl6OZ
XnIvulvB8F4uW8KfImpEmB8KfZJjKqov2+zLUMhVTnlbHNvbveyEw43jigNDPUbNe9RgfMoM0Gei
Ls0ixCG0RN7NDOmoRtaYupQ4UR+nKUfRcLe4wEtLimy5YoGv6sxuel2kDRq9vSUN8kJvFU0VoIxl
oLP09boa32IpO5Ik6C+x5oaRdWai0lW2he9aPfmcUyINtHzxm72xJRCnYkTIH5y8JHhyRqOItxUm
HX1ZPY06y2W31yIvb93IEm0AslR1doWf5K4AXGTAVDX7+32Gm9obN3qhUjO7trJN8p7TO5KWORT0
u0rBMh3aZIXbntTwLxAkOyrdAlMSfvWfHZfQoZU6R0Zjtj+sUaJHIU2ZyMow6obSnK1RePlWCzLo
yTq/JKL9apYqTy4kixXmiQNwqQWtUjV1bUJn0EHHt8/e4WKpHjrff/bPj4Kv4g85w+LqVi+ZPFUd
dBeQgqwQ/xMWsBGDJDilTfdBF4AcwiN4uZSWu5lLdwivoqISqATE8nGaVABpZvLGqTLNharov9lx
bHEtW+QVvX12dI7/KjD267kTmtKvqvlWvQmwqAM669JRgb0mF5xMoVPJVVohwjPgpARu10f0cBJc
02LSTbURr0Oc8afBbEm8l9Nsgb7QlitYsUNTJvFbbYn6E+lOWvJZTIhrDgz/Iy94yGUvOJRvyFu1
ihhwWPsq9OgvVKxRVLGhEojWPidgsl1SbTGvcYWgorM+K/MaD+6wJj3pKVooG9Zslg665VxMnkXT
50ii69X27e1rsAgmw6VfjXXk+rh0S0SK9uSBg8JaPxJV9nHld4egqd53BOd3W+rAxkYqRTgntnXH
qUN32WSx57xDj9HtHk5QWweLfVtvLYussbVM+kPFAbDIZvt1keWz/X1vWfL07kZzouxUXa+jAp/e
eu7znyh+cIMFV2HE5575ontoNcihU1n2Yd5RDyUn2v27vZbvLEFsZIFJiG5ABQA8wIJ1Rh6dkTXg
qJLF9mDAC7O1i1qBQZHUyqkqOc8PEdWOd2qes3PnL80NZT0CXlYZeh/su8Axrt3RLYljbXYEBY5M
YHfDtQnyyXNy299osxiwUZ7Y5M4Ejy2liFw71I5FJ9hlxhp+bSFIJlxo7TgARocxHKuL2QzNKJAi
gj4epEuUyUxo+tCycWdsMx3VISrhFABnt6WQwheKKijAfzutR83GaExbE6+FjORA8fTG7Bt8UHaS
TduK3lPlIBuQm8A3qwRQopglQoUiNE+tprRZdBp364OkqVjpGCNrXRc/SueCmTNUULvg5gt0xlxT
x6l58ivnAazeGq7aWin/q+5CxEWFR7MFNsmEl4erpY9jzSm/iknUSEjqY+wzni8cy4xXOv06tW91
dtUOmmnn3zPjvKMUd+WEHom91dbGcg7MZ9GEzj3p3dQgMYgkFJ+3b/M+Rhmwb6BxSHL6QN5qVFQL
jemrfzNPlw7rvUAPBg0MGKnIlF7J/tgxdHQp7kFb/DHIJCtDUDp8JerALDwmefUiHFBcTQ6fItGr
cgvlb2nuFERpUutWSNrfzQWY9UcTyBvCX0RZCbcCKDh3gqY5BXXvHp5XurnUe1/Nqfn36Ws+lvA9
GfjjMJ3r/lZUn7BqlUGPdGGiGRnkKsvrxkH0S/KioLoQ1ampQN7kJZOsnNJL6GVor+1b+swOT+2V
OsZBlhmFrp0wwpNnRWtVKq3PuJT0VeV1huZBGzCi7/Nrh3ef99mZIf8OEZU1GG+Js+HpEh12z7pE
4rnmrfjUBl5U/325kZyZU9VqpyZeijLg899Ji4B3QkDFb+8wWN0JasGZ7FaAdffyzw96UCyyrH/o
W0GA4Anb5B16o20AkMQ6gxRVjMg3J/xJaUeec+IcYZ4+FUD0asL85W3SJKhTUnnpAE3EBKO47uIL
pvXS9JiqAkm/Ww35UYt9AXgeTyPrHN+axXlTEYzoZs2RteDo0EryR3o7W0SQTneTOyRUgt6PrGO+
roYKx4KsShbO07PtnNpt4sp/SDX/vgSSC7bsqWNRSn+H+6OGh2qKCHANpjrqz+SsqiVygF9qcQUk
w2hMOALkPtDyst4qstV9fhrR+TPbuAfJy74dWJ9s8M2kcqLD4xn7y88klXFCa4J05lyHWI2wlGBe
BWWLgzEdnYbWfQcsvq7EfxxRw5VryLc/t/+/5gH7XO/U4/zRZeBxUAfcz3lwWmiE2UdgWjTzSLJ9
rsdCPQQJV9egI9trE2plUXqlRPim6a4mKefqYElGtzz6vM8Ru+y21q3T4YOHfi0R3qK/JAAf0Lre
GeqHXxqcaf1PMp+ajAPhDo2vgeX1Ln9+0tT7CWO/RgbxHvlkzoI2exaYZfJ49x/LEcOh8tGgcgo4
LcrjOZTIL3khTqb3bm9ydPImiXBmzxuRh66SmBxWiLAbVUtSyudfFgmwIg7E3isw9S/SCdhHOdPd
tvyhygIv4SeV4ZfNXXSpEGxueFBb8mQuwRigKWZ0ju6+GwIu+sqhfqJnvUk5lfmwjLm0isudwkse
nYLcnd1Vm2IoRNxNuiTH8i2l7deMxiy0MlkRvuq0Gs4vJ3XVJgT806BsE/Yiq4CzoZimEvlcBCit
RsXH/Y6YbFCAxxCt4tt+L0+XsgJ/k6XyuVnUCyS/Jw92V2v+VUfap8HZWx3MBDVWgprfb/64g9qC
8gVeRWS4DDsgLCfdVeLst45eE1C5ILLzBDBi4J/T9jsn2fAyy1A3Uz0mapWkFbe3EI2vp6Guvdb+
FnX65o8UZnEDujZoszRjER2oLV0kJx/6jzt2+Mvfm8DKu5XcU3IN9PGAuZm9yAMTFLW6KNHihB3b
LWUdGhfzK//bT4pSSo7Cf5o7wlMhRLv5aKFXE2kzkoMl7jwosph7ICeczHejIGOZfW/KKcppGs21
+cRjBiAVXyPM3Y93YaYw+DD/OM8vKvNpTmhdchVgwaqAYOf8UxW9C4D9CjhyFxX4xdhlTH60NUp7
TBmjVyJKD3PAbsJTGxfPYStu8V4E5TlYvnUrjm/cqbn37NN2FK3fHzagVsB1z8I+fmkniys5mJdv
zzMQdCVpVrPegABjYn9uKkmryCmiK980/jBY/zgIpNzKlcvCcqlDVmoQvriRhB3RKpxdpBDKGSRC
EFjBJHyCctrkDJuyfs5mbBqREjmtSjeSBjMg5iSQbZt5W26tlsgcqxSSTZHdeXpa+7Bbpe6tpqSd
sf+P8yqE2KpFoTbosDmYx3JBpuqWuUuf9e4vV2c1rOrAoWDgT3G9lR3pC2PweUAY9eQhYcmaqalP
2hOEJBpSFzr3Ldm5GyneEsRrKsYrxicDddGu0XMo+61I6D0s+nCpYe44XEEwigHztRQFQxR1CWpB
wdgMeJZDhj+8SvlbvqhSTAdZOmC/YsUrOqKYxzyZsmAnsiHpIzPwaKcZDSXGgoBVPtlWMctZvOPt
Ic02a2+951exbOSdAIHWY6V/1J9+wXvV/K3xYyN8XWtfkYdcZueQpsqL6X+Qcn3+H1Rh4+V69bJC
qUxRJZ+hypKMZ/9EOGPdTE1IOwkndvKRrxkQ2UslED3x7glfEFfFX5SnWfG+ZaIWOd9yABVpWdjP
LQVELw7EWylRZqSkiZ40A4nyHAmMrj+dBpIYiOzOxTRQg4vUZV5AtjXK9zjXzcdKsVphMvBF/eT3
XzsjS/ZogU/ibpf5CttBalt18SdAIRnusEnLDYvgE0ynHM7P9B+8Kw06mzokTAuRjL3ijP8GZNGO
azkKN/IDfdFtKxKItScNU8t463LLhbOBUFt9m6bz9tHXKm3ih4FYe7Fpjc6nKvm6ekLX0SKosVkP
rMy8HIX3IhAiNjB3R+KIippKKH1ZhFGSgBQWpUf3RorqYkyUI7d+diHd3IqCg0ZsCqlMjE9IdUUK
0QtTgrfpdoyjExwhFFr9h29SD9tWdCLDMS9IaKt0eojIu2gKwFhzbZC3BajK/RRkNz0ZkEcUMC40
12jI9dwv9JGX86yUh9eSdsHtATi4Jp99bzToAsFyPlNgNQSxsKY8XbRpbC9mOy0TjJkIOX31CIei
vy2pxKnoTsIgJFTZBD7/9tdVpsAYKah51KE9NsrKs1RaMdPw14/Ue1iNSRCeCpJsZigkEdHxfQkx
f/PoD+e4SH4iBCUU1w1WiVI6cipKZH97OQJqw+fWJZMrzbqzRYx0GnOwDf7e2aZbv7gh0CuUpR6D
El6QA0HphYIYxiWNu2UtLfJvJhgHzopvFpWuYx5vhQQrgAxslVdEh7fliZb9XWC8n+aHBTlgyUy7
q13Jew1QJ52Acp+mdqigsmiFeaeIOeqSNniLgU5pLPQWFWHDIt+o+Shy97AR23PXSRPPAkd5TOYs
bPNTGGXGvelxaXxv9rhaIkVVBxyYDLNMQInCTkUFydthjGmtrHZqN9tSDo9EjoOZUvXLaxNinG7h
W19npkAOtoI6jQZGCpFfWm5NDcDQC8YNk14UPhGBU7UIWSrmLC4fUr7iNht9J24yJ3OJb+t7qv+W
RiqWXBQ8VCIQVx2LHf/OOKxEtamSiSkmxRjykP5X9u0lHuys5+BdrKiaF7s2zKxcMbs6u3N3HkB0
LddEsLLCf8Ae5xQTSVNCzHAO1JbWM0mivuuOrrd4gGnR9qNCs4uzjTSIFVDpFY0CJ7imbUkWQF0L
C5ZLFEvByoLaWYa4kQKnp3+AhcZR9GZiTp3fpIvVQXg0nC9XVRVZeCJ45YZipFfYBMq9Q3Ve79gF
aIq8MIxd4YlnvaUQiJ2TsaVaiMyzvIjZ6ymlGTQ6XH392tMjbUVHyU7T0I8qwoeaHSNvhLv5ztlo
Du3f7qev+gueFZSY/KBaTOFtnuz+yqcsbYpCMDxk9Q87uXBNyLI7QjJqvBTZQlOn0HKtWfCOqIY5
XzisXhSdNudG+KjmGLjxiLO4ajNneOYm4fvly64gXDVdQdZ3W3NiztmJIDct0HoDnmG0q2z2miP7
j7OEg2OpBDI+0Bv3WR80XCoyuHat4DZcEcBibYYAFc0HNiBSohDoaDWztzrSgm/JG5rx/xbI1UQj
ZoVgkx00pMW5xclKX9PMS6FTiGb4PTuA7lopQucnKHPmsEKKyDoBfzVQZo8B66DcTowLKQdl26e+
xbGr4d9/HYleHTxg1g+HEZ/F7G7o2MtS7GqWWw5hePJco2YiaUVbmM3nzbHkUeh5g6TkNX3NSOqK
5ggDYXd/wqMlU0QX1VzEbwEAsrg+WseR00e9QVsZoJ9X/SQCxFHaApfrHM0N7gyAlcjzXnPg5qj1
YOql3foeJ0570pHdZ8nIpjheREqlGv7ZxWCwa02Xtq5lG29zENO29pOJyMuJc/Xgpi2wbpRRMmv5
/koQrbdO6ADPLZifjPtFx8WfL23+WQkYzPcAxuWtrbsR3X9SBVhLfYvQgwLFVyDGmwq8ABxGGcBh
+eWAd/TOzLo8cWfNxzdEcZHLojZoAI2EbNAm3mAXUZsrG020hgCXHp3vwu7SH/ZTIFMS2EyjcK11
o1KQNaAZVaSDJXpLeDky/rPCt9+RCyqxrBkmxCvjWOxnjcn4yWVOSvWgXv00SIsrJOax9yW9hHnF
AN499Sg/RfmTpd4aKWGMejRwilHORKDqB+OcuzXQjuu1pQdQwHZD8xLu6s4h0BfPTspk4E9tM4d8
2g3GaDWJAIk5a7rEjipzPsb+BgoYsGgu/7LqCdTpmBqjIpnI9kIZVh0NoC3VsXsI6VVz9YptviZ1
UgeNBQNWdhr77NrDc9X6GxLQ2sAC1+yE13CUC9iuEhMqlcKQ2LS8exaRhp5BVkgHWHe5CjWYQDV5
GNQBeW3/reTSMXEoGyaKQz2/IA5P9TIOvNASU6QwDoRRhcYElAQv/+DPdNjY+16gqOrtXXVNS4Bn
4s7WNllcgkUiRY951KaX8pCZf2pUeGiFlcGhxOSKDlNvJEDLNbdo6sMsrIlKCUvtu26aOxdZfAVd
ugk+ULSnXabzzvK9xx82rt1MKMRf/bLrE630AY1j6o3SytN2Zp1GrIIi6RRHNyixVU+2rK3MmlAx
FmJ9WkoDYpdqudR/hwlSeLiW3k6UR7jhCUii8gIfHBdqN5IGVB/G/mfHcV4pWCeQN/DzdrDComx5
ellxPR+ew8ZsuHjHIah6O8LavBBWiNcYBeOEqMsvlHDMRXIMtub7XW47n9tQpVApIQP0aUkDDTaz
UrxbkF2FLP915S5f3P0RnpbBKtRNSxJUYPlFgon5IKbp/oxqoVVAg6mw1PNnzZxrPQvAA73mmteC
C/ubzB9kb4Tw5pKnS0Jnc0lXbfit/utIXg+xnOfsXKdhr3+d50t3xCHqsIZEXcqaJmbd/lu98nom
ylJ4pbDYxI9pHhqPzz59C0h5xJEyHkYl0cIMaOVqUtsEcnK00x9M6vLT1XEF8BHwFALtUa6lK3lj
/QZNTkITgryuSqrYlaBy3ukzPqJJJk2U1fiBis0Ak3y6HAiQ8PVUDitXoBWe40LTWMlEVVd8gGc0
2Kyys3Jl6boMhg1gRycZl5QAbPOmA/euIH+6fDOz6r/cEHK/WauuULw9Btgapj/kepzdkwo9KHSt
LCtQdg7pYWrKfsbDZ3uJprx7QJLPNircGX0g7wXgf9hni49OyIGt1iz4vm8RZYvvd8Ma6mhV81lC
0NC6vAP0bFpuUMTMF0qMlkpf7GK+hd+5PVJ6xNgxM2A57Cke5E5N68gUyJUSnUVs2ggIu/X22d9A
VEC47wN0ykTl0W0E5gmTFiMY8oJkb4Le9W0Jejzdj3y9J2QqT7T1Vkgp1zCIPxrZpRioIFlMZQ3K
rKzHrMataa9JLpHC2q6l60lZTvU1ukWcTpyz1Jup8WLp3m4nH4flIBkFbvTO0YWuzbQ/DIRL5aIk
+9L/lYjKqC0bW6nIkN6T5l9SUXgCxe9k2YA4nyfC+Xh4SglDJorZflS3HMr3BMLZJsJtA6CrDQea
vp6cJnDCNB30jjC9quwqN7bRJGJdJAoHnyHGbJRY6gm3Ct0OGVMgcJePHvlCGvfwBaRxiglJHPs8
HfmsexfW8Gi+0C/npgkJGtIvWdh0SPeAPL125ulx94jklBR6Xd76B+Np6sTlCKyst8xKz7t0xWIx
6odvMqSLEctMggNOD9PUjekX9H4PthFpDgirtCHfr7I0gzgiaRWBzFO2HGjlwqf4HLMPQHSOALVc
X/e561Wz/P+iqMQgCscXrEILQo3/gMkf2Btj22kob7l9wpgHHBirq1Zg3x0Uo4fhddBf//pnKouB
bzFqlUtB2M0UVPVr5/oS7sxAwZMIiJYpYBjEDLoXYc9mRQymYjh6VM7YnA8M5v1r/+W6mzjaXshc
pPZMOuALqfU12REdpYaAQ8pJDSP4B+nFulIYPcL/GEelwPst3YD7X4gUNLif/SrOeMk4vjlthb/X
Y5FFsHXdwozq1PgRJfdR9xhcxSlIPS2IX+CH1zDf0UwjqSCZOxXWP1RKIBeHBoIa8YDJQGliwNTu
dOzuLEjpVxJNNuMv2qfbGJBAG8yfPgx51VsRvFssescXhbVjRgESjmb8D3PJU8fhLlSMDp1f9asH
Gx7spWVtrMU0dQvQ+OLm5Q61SDBGFvn6BcOFar7R9RPrqU5Se/kmGhnr56W2a70GxZE+vEZ3Yd01
y2Rtpj1c/he6iJwWM5w8F95iWp/HTcM+8eGWKQJWpfvOfAVUUpsrY3Y1s+bX9uERaIgePdeWxvA5
4BIUkmXGcRgXKaTzeYyS8BSgznhesbSmVADm7rS5hAJMOqYNnbuo8jgiCctyqd0HzGAI9LE0PR80
Nt+B63T14KXzjt5tMZhGY1jMW4mDVAPpb+Xly5gTC2ed98AtIGMYpbbv4QXawUz0TLCjZOBNmm/L
unj3QQ6M9hYVGa0TGCJQVM29lVNjj+BGwW82bJHGhg1lu6N47VIJ2kfyf1ERT2FL+46nsGM3MOpb
7GrqdY75wXnuJysSKCr+QYk9vU3Wvwn37JQ7EzKi6EvrB0WvwUG5Ul8vvx4LnhNHWB7W2oeVdAyK
oq4+tw4BxDZIS6a0AxQTYwfowpwIUwktbgzrWDnXpuwFSglarlCJdsLfiWFBtGcH525WSbbFyku3
hFzwjNMyhc/+aUPzqvBb6i1kAEc7eK38Jkyw5xnrXSodgjo1s+ROxNv2EZXNmCibqC/hyPjijs+/
+mKCNg8Q6P8f6+PIEoVc+4i0efLZqBZI4J6M73H/2d7WJ9NYVX+e5p0d9w6toONDf2K9ulURu+SZ
RHFKnL1nUFsPn6p2RunUn58B8bEkMHM3UpQwE0JL56hNNLRUJUFNOVnJmbeZCORmaQUbHyZRjLwQ
vxaACJ/Br+Z9IWaLivsX72s6P9l9LleV3chqkPttVtmaJkw9aVniJej4yXRpBUw+r8vllat/OGcE
zwKxBM0XLohk2XwlmS22yQwX/i1BJlX33SlrkzySJj+qITQZQvBhtfZCOUOEssq1inX8EXfShVEu
ZzG8bod0aKRN8eLzpeovQaUjmWrB+TTwgjdy8ioJJn57PZr2e/X6cLvzySiCyEbhmbqT2li97yWo
X2G33/uzFBWIJvaXeOGCiSQoFr6MsvWhPjNb7nil+1nlrdNtAQRn2U2fgBEoltIWVs5ktbiaOz87
FLKWI2HnyK3j/KM+MrVS4h/jz8N5TPE/Pb8ZulTY8lIK1O3+Dy1HEB1kcdAmrWNOb+i3A8ISBRTR
NqNWeL6o8V5/QQtJLHF4+89qTZs1iDHkH9Ou/pKGY9JieA0YIC/rKi64HScV11LI4vRGifSYH2Bz
nLCaNzGHzzfWR+8DrO4KYuy+Mqw6omyjrEsAnOx4hzwq4TbW+mI4L73GtiwlXtGD9jczyBK+OAxN
xM0VJoBEqDHsCP+QqAZy0QmKhEM981nk4PBsJuNcMHGNWbgljJixWOaeuJQUfbHxIEiVnPFBqOmU
gtY6/vA/v4mvxMcj56td8AUZTOdGBEHzY6khy4QHmJuwC3NmFs80hEY5mAH0eWAoAMJ/uLIRY6qA
1HCvzOx3iFumsTzbw9Bf9gYgKi2btKPyrQQJYumavgMdeLwcW7h+s0B3RA4JrWY0ZAKPvXpRuty5
BwBBSqnFVv0MXKZUzNFNfB5QLGB58d8xJiiOMs+8JbpBoXvfkedN4UoVyFmgcVXgw1Rvji2RKwSz
0UxLPL98KS5W3fpzCBLBIPB0agd4Ju927NYOwweLGwY6TsZn4iYlWrbkv5jvhKyRObe4pLGTOmd+
0xQcoh2zMkTSkDywqsm8N8HfJpRYukmKusZk0COK/4DhGll6+uf8m3oviz5OAGkgEPmbyiaHCFzE
UujFLuZalV4UYu+kJ2E/Rr4DRJSuDYmVl9ytqmVlnW3WNgy791PlJmjOYR7va5ouLlWdVxTsZi+S
UzR9JknzOOg5nDdGxWpaAGjKJ/RRYA3ehFBMTEGVv1oQg6igoA8Z1cjIbOQNY9nhle0on4tMw5Ml
bdJD0N3gPElkCRBZVD28pz/HEEbY8XBrLWiklzwqsH7Z815+BLVX03a41Kh5vvrpidKjI+e4Umfw
zahvIq8wGXYPgWpImMy4oT7tjjUqrRFmTH1QHQOrnknZUwaLB6zII+KFEKJ5fwhcOVIE8EgfGLyJ
51rx8VwJia6M8iXLWPePtcENP9CwK0zsTrfXhVlUObdMYQknoSEgFCacoL9FcoWW+g/6uV36ocYy
5FBJdg43Nc50YN8HUfYCpsxzIIaUb34e5f33G4HUiD26jdgP/K4FkBOR++d71ouJx5g3izxqX4r/
ctFnDgngqz5TvPPohZQAJ2GkIUVJe2fsF/7hZvUgPJ4wVHQ5zv5lQwl/f+WFyoAhRWIFd+7glGEu
+pjxJeG+fjDIpvlgt34OOovTOmZpZew+thWOQ5CyiP3ESBPwqG7rC6cd9BQ19BKppH8lcsn1P+K1
bjP1DuoUiGD3OaGvFUK74LtEDCCiJF086j3NZyEZWhr4DH3zXDJox9DNtQugSQj2FQCZWpvs2AQa
maOjXLxUC/e9vx0Nshh8M4mZ2mF7RlN+nhvtSANNz8ZaFvraUWGf6xfp2c6wlAL0mhaXJH4RbWCq
aXmCLmEe4fnfWGZ0lRL3zwH0jrQAxENwveDL8KBjwjunTBlC/FvbL6DPgNyPZjBFy/I5W3ZfVBkZ
H35w04D0c1ug6p+kqSj5XR9IC2ZsPK4xKA2CQiGcq2RSgisBAtnm67ARY62+5o6wdK1JatA5yXbr
4zj4Na7jLUgGKphBm61gLUxwdNOYXjph3BXihzLjKRnM6ftU8LX9RWWcZJBXYTDuZjTLarWJBbUq
v1+eQBltJI7xPep51yO/EzoKp3zZyq61qWuzA5JljxZutCkVKWhDAbcT2nq3QQfncKNdi/qTUh7f
uuE+NEmOxV3heVxxCwpD6Vl6xfNqfkgIIJmzEHUQ3w+N37gRxxmBr0nsTV5J+DUuAvVzD1jkwWAu
JTNJ2LJw0a6AQuct9urtJDKRwb0drF7nvQTNE2bleowyfAUm5JTeFtVj5o9O9aWeXcjk0EYFwdIO
WAQTCNWRKsCXW5b8G1+O33TrnLDjdJvWYN/MxmB4Qza2x96s7j1AxXCf4fMycDLwjXJwb5jgsVS+
NuoAPxMy+XREJBoyHkB9/4v/dWGfWpcOCzgSgtqFrbHE8WftosjpgTjJrolspBH2/l9NoDUjA/Ys
hFRUckma24THNjqkaQGaIwip1q0Aitpg288yX1gyZSSRzwRP8BYV4YjGumwnLN7L6a3NpHN1SJep
ImbtPgJ4j8F9b5m4O5/Lrkrb1ZasEnzh/5bevZUnrOdyAZAeK43OD48T3SATJg13gEi7HA7n8dBN
debGrny5Jzs8K40GWsh19zbVzuBf7XLLoY1TJLOZOnVPH3njkn8O8M0onK0RTN4vozSVsRKBWlcF
JLzNsNYL7qTs0JUUQRDaKdoOXyl6PYW62NygujcC3ESNAXr+QU0uvr0pmJvgGk1A8LfXux8vwJyA
0tQoIpVZuevxaClMR0SClxx3lNH9R3nREAfJt/Ui27xRipXVf/FE1QoAdycU68kemIpx8firWxmV
dJ39w7um/8hQ7ADnYjVeZLTic01lNg2/ummn6nQ+6zjP2e/svYDwE4a1a261P6XK89BwdXSlRc1R
034RNyHn6An7VDP9Zah45Ty7nyXwOxqKKn5lXmbIscNTxdC9HKnZ5vgqI01AGs+kEr59MJDodla1
Mgo0PYyESBqzN2iQovRh6DDnxDVjYQtbmM0Jt8YUixv1argrmrwRTbXh1JnA332ioKrk3cvQb139
UZnM/N6dIbVKlRGNRD9mS7uFESqmBn4K8KneAV4oNRlerjEgkVYE4lwNJUxLu5x7GJxM1IKJpB+p
XTZfHlVtKExogADLwhFq8Wn/XqYvyC+m9EgWhK5CDzxOPRAnd/3O40+83LM9Jv0bXR7mGLJC3aoV
+/DvaxxaR2VZYYUoVS3Pwibakl+z5w4Ssdk9a4oEkiZeIlJx9bX6MnRHNbagVT5NXP5Nfc3JCPX6
b/bk5rc6w6l1mVB6xSYIA6WLa90XAj100mz7ZbVnDJsTTAOJzc9z2bsoQRTSXOvuoyHefUYKX6K2
GtRsV0u9VZx93viZUPoayhS7Qr6631TDFqZYHP6N1XLhvV3KBJs8ktbZ/JJSD8cD3hpJEr0WrdgR
24e2dI4umiFg8RCf4B4M3YKmxlItyfVGsiAo3BprJWq2cIk2zCL3Gcr6lCQTNvQ1QnuJcRJY5jkv
EDiMcp4kMpQVr+rXAx8wOw76qHTIc/1guBCvfUUQuyDBJvt4c1pjX1dzf4max3RFFK57U9vUPZfc
83H1PSABQlUwESBTYS/qrcNL6OKapH4pZfTS5R5KzOzTanAXTPC7X0pozwWf2UPwhYOBnHWEJgbg
yTiqglzt7uPiq5Bwm+4V6S3H71ubiuIWGSa+laElh3Kz//dNXdGqH1gJ4vug8LI4ChNdypQ4Gxtb
NDIDTHrbdw/7FfSvTcFSlCi+EkRw96YmADfZgNz1SxqK5w1pHcBkePUB/0UoS2lV1W+aw9+8sPf+
QPqGz1UYtS2l+JLNTA1R81imCXCikWhn+hUtEc3qz4kNPiYnOlaQ/KCLF0YmYqtCjH1eOf9XeL9h
yV680eB+grT7gwF0lTB3DtDQvXFBH1IPuxZrgdmNZamyxxnLP01YYvaHPALqy4JfPSjqIURIxV/k
gZBXyLptXe0arAOl8pbXjRRUiFX1Mxl5jEydxye2osXeQv7cCPM5iVD48aaTLf16c2BucTJ0jixH
spdeedbGSsC+fO2jwKzPenUxPZXTQ8yXkr1NDMjowHMyvykBW2k9l7nZukwFCtD/goXJAPt+R5ff
VbIwaUlzfPZOYWDy5ZomJesd/jyC7aDr3/x/HnQw12fhWhnAv4ygCdT36OcB0EusiQKcRO5PQ3MS
kMB4n+ABKjaAdRaZrq/BCkbc8nyeU77vPTLDp9ZOguE0ClKzUrdwy812siubwWhAmuDtBDrXEdhC
cAWMD8rIm3s9LUt7vOujizTOBgwq5orA2dfRl5x2lPgZtK8ze21zA9v/KgSDxOSf+XTy9dvVAXJt
iz4IMxHw3ymv/fv4qp7ohACzdPGvnLLO7MpDsxHwtV+CETGEhK0+msv0QzIb5WqSbBF6yT0YZUZG
BZQcVqBAzNR/gkCj0FXDTPCNtm5rfXdPHzUK3FMCgK5uR3dOcl4tGb4Igddbn8ny7esBGGt/13Zr
T/jDo+6vA5WYlMA6aYnZUb9XSYpP+dwj9KBrKshWDi5IUWf40kKohaCdNJVBXhOpnc2lG1OjEx5y
aSMZecDkhl9BHkFOAcIIm4AaDlOJwLMskJ1FAIXxYKd3BgN1TRCuykB8NSpGnef61cvBPJwBdkq9
c10yXwnlTOFY8EiATvTLagLgjWyge8Gd6ztd7UrouIe+fe1b8p8SI9e3zXan6+q+VgHgDuaCk74E
7gSpCnx2jFp8xOwiSU/N1N+/xxv6g29PCG0esTXo2FDT5MAvJ7abQ5tIN5+zIMl00miYQoRF3wif
P/0D930HwGbyQZFMSwarVQpir22E/29N4F20VeELZJ/KWCwuYMQTGUoBWug8u89l55zugIIkxigA
TiDhczoac7MdGphLy8s3DZXKT4vkX2t790CJY4/ODh2pKa92165EiqKndSm4m/BkM3+c4umdiTzf
1OLzn8+REVkagkoin9l2FLDch+xpyhPupDu+LXfVUrqEQToe+EkBCeYmfVjiOEezaes0lV0W9QKJ
AV6g0NUfgsvaaXbVKHPr8SKpsom1dLGZaHdW7tk0jU7ON0v0v6iaTagZT7/je9/YoAqIWoQsvkET
b/9Me8pReZVK3E2qkem7/BDI0wNXIaojGV24+B/ormLZD1hcwHwsgi/EJ5AGHecUcqCMfCFBH/X6
CSU4WNk9oKd9HOCHD6gmBrsE5b4kHeDyGW5WKPF1Nz0ChpHTvsgMMdu+j78hrtj3XkqKchpC6nL5
cAO52gEdxg+09wYcLiNk6YaxgFcfgHKlWbVi953jYltwrNq6Thgw3cofDdOrZ9NMXbxXtokfoR2w
8zfRupp28raEoao/KOEvT2v0IaA6OgBUQDIeUynVjpaffqKH0SEYxI3+wKV/umeeAR6pUuLKTj2w
yJ+3JknEBR1GGyuXCYygWxIxyIbj42FLsm0HvJax6piIFhKROZJ0FkG6vjPO8btwZlsJOk3nrESU
l2kPbQnFcJFaV8LCaNlyN2dd4SbUUshadh30HOIibu5vzfXFhQ6KFKMrL7x1bHzv74jVvI7ZMFxv
TB1AlRPHqDYyE8390cIfANaFrWsUSqFz1LtrslE8/S888Ju27lvEooApMrzPocc6GeQVC05iJapV
6CqQ5zAduaf3FfoyEUFubsePoWxzTrxZOgNlSohsmZfk2luf8jy9fFj1zlQqdueaKg1TvKbmbSh5
51TMmR6JhruJvI1+Q7E5IIaH+B3Z+CU4xjoI2RL3gxJnJ1vO50v9GVVKzOjb+ktz9FCOnBasj1oM
Wd8sQE7lBMqu+KDqDwlkKyq4KGJNLe99L1PySniLXKaKl5ijFRkHubJmlvLAgv3jkIRmy3EJf7O+
S2n/W9BHszyzWrdYHxzRH5gJOxjCK6pPhFPcUlbpO4tSILXPdOroLIz0MctMewf8ORz1/bKHcI3c
1ozL6efETt01Mz3WEdCnVhqgvlXvC3sGWVPVApahCGaldwbsD7LjOq/zDTvUiEv6xTnBtXXgPphK
WSjUcgb6hRs9/j/q58WKqh4/BRflNqkN7oYSJo6P+aLmvsuGlZDZjaw+JzMCAGi53nCO9562UOO9
X1d2cjqPeE04QfnzNyTYqjXY2QVgjHSgOZ+kb+3tV7l750OswFh4QL8UL/qDy8h0efEHA1Gx7/Ol
XSL3im54IiuPd9UD3NlvNtSYRH9/FFDrTt9O+Ia6T/g4h22iXHHdX74JphxSgw0GB3vBd/2drdTt
0epi1HFM6JcR6HA9/81zzwrdc8ccsLDywE7HxZ5IulbHD/MP77GH/M2mE7a+zxrkfyh76PlUx6d1
+GzNzI7lUpajKCvZKJKuOtMEsayR2clcc+f9gQlWe+7yuutxoBSmGNmkAK5gFxPbeFX1RAjci3pJ
g/lIcqzkLOw3DdD88p1a+OICS3tikzL0ksNy1+DV5EaWyyoPZ4EH5SNiaY8u8ji5I0vBAD43uBNu
Wj7WeIEiMfpMZtHD6gCpvraaqnvLvMnTSZNA84qRopJdtxrrf2mm2V2x6uUeAeVuov9gpQ4kXphk
eqMVnbnzli+czDsonKnD2ZsPbJZSrPFUbX0h79y9LUjOS5yHVpf5Vf4CMt4pmnwUgJtGARhpask/
zWZ38LB46OSY5ZvVIwhlUSWRHJ5ZhWFiIQnzgunp69VQDAuw2XM51cJIe9gMnuCcBGLp4Tmv94yj
RifUqSLVW3yEQuezXxGI0vfc+4NzIyUx2SVa0GgDLy5Uk7KhFSBZv270+mQ8NEJB22og9knONdk8
Vs0cHavWcXezBD9dMgyjC4SOiNV323QKEQWUwq4onQjTKyGkx4j/v8cH6+Rx99Dep7OrvX/FGps8
AyFNjJfQTBZS2Sy2Yq5dqC9vgw+Oso+l3uWLkVd8Ru5wm0fScukU2GRC5L466w+d1Xw0Zau1AcTo
uVjl+Tl6EFsgabZm6O2O8BGzRDwU/uTnYhE+HFdnzffo+CV72TDF/uY8dflgGuWiQ62eL/j3SnIe
NHL+EPredqXsrpx0UeD3gNK/rD3qnlXjNydqO9uGpz2dQXnpmXHU/fJvP1XBSufWc9wW2azWPxOC
yaY6+7kbVEcsEKQJOPEgbNDim0055/b/3UD6lrXIGRt91yvd2zV9MqDCJCHFh0XAMVvwcp49TVKQ
ayyfsMKcUysqPY50DMPvU2kpY8DwHWd9Tp/1dM6yK1J07JKip2ENQ3WRoRixaJtAAwN/KLjbOsCW
nAbsYfqYKfVuVJHnKC4uAouAB1AJNpJaNAw6GXcnBdLs4QK811vjGApN6Bwrsi/BWWa4t6Sl3G+t
HrMGYZxqxmVORbBt8qrB/nQHsKXd98HPMYtYSDMOo3lQ1Jt1CuV0UTBYXH92gfmYDdARJqFmE3b4
PJXqHDxCZ1XvuzghfPLaznEEr1On6IykIWlg3+SN6i7AH1uCci0+2FrbfCVF/ABI4zsPts4NLuLv
fVUULOtpShYxTd4sRF7eE6Q/ypA9LW9t1Ehe+jxzfIRLmimKcg3YSMBGu8QOVPGhzz2sBwvcrn9g
G+QoxQHwCsW5VE8UYBV5I5czlRpH9+kLJ19GdFRsVjwl6xnAEfYBLjE2dhiU8qQBcVBeHQlDuf5I
MsofvtsR8gFgw5LAuG/Y8iozQSisjPKDKrpTCOxxEmZWlQqqYqCwHPO6DSzkmEQWgZbPruHqbuxm
B+Vbitl4HZOHOm1vvB5wHf9CDqC5I5w2CX28nnBHkhX7qTPd5mT578h2p0herln6B7yaQwU5o88r
FilkoSR8/4W6Hi9WfYvBL5THUZSPCJjYRVmcHwab/2iO9m2DB8smech0FDBdUMVXTabSLSVwNubg
6CXhGS3cQzUjjCsgN10Zyu40VLcAUF4y+LI1tduLUTfAxIA3BEqmSZjG5f9NAFcwB9c7vk2Rrmz7
ej2n5Eug13OgGuQsMhb8L3Avxwd0eUXEng2527l9r/nc5CXsEBwvMpIzDx5RYsu8cs56hPDGMWnG
XTl8GBveqQbra/9jmLmZDNu2G+wWha97f6DSXN1W7GeWW9cGWLQGyj0YCJxD32z22c7DyM22K5lx
sPXPjg7SmHAt68YWQcWw6nI6TQJHsLuy3bCWBszDJRoHwh22KaAmHZEJ6K5cx1bp3F+bc3wonWBY
EWBlsv5BbfMD/9O8NnzscH3qyz5SoWok8/f7f7XFP/38strd5yl9jw5EzrtPOQPGI1Z6+KO2xJpL
TTeaNQs5lSTpswyi/2TxeFEwl4ktbGlK+OEZ7ifyiyZDwISfgGCPOSLM21lWKqav5r7TmQ0dGiRb
usIOjPwP3XAHl5SFP+lgUIpT9iOnkq7Nz/SwzOfQgB9XApB4u7GoNGeIlv9kTlCAJnBXWpz/4lf1
2mHfsW+DNu5MoK4mnTw1XcnvkxqtXYyoshQk59wVmNHnt2IgVJISCs7e5eUxAF09/0PmAPPvc5Ky
pJ3znu9rK7wSN0MQpMfx2sQC+ewmQRmYVBUP3Ge7fC/75snR69OiQv7XrjMvTPIsrKLOOeluEdfZ
WhEXq8REo2r/IRqsEVwx36pg82mKgOomN1hLbUnQR42EYjUraMol/jlJ5pk5VVrrdMNJgYlHKT51
HAgk9zo2E+414DteGQ5EfExpB8oh9TbZE759byEt1VS6UBcQ56ddvWAJyYYAyqW3v+7wUCHVZ1U3
2bqaomfrzyLBEodHBXlcDFZsnM3o7iocT56k2aIu2Uyf6EAEOV4y+IxfBKX5plV2TX/i093QeSSV
0/2JgAA0uY3SavdT/bAK2myIMgpud5IaCagt6dMX21LR6ZUb4UPqOCPOH/fAOLgEZz+NgRWu/GTR
Bstqz9oCWtx0ZlwYJDjdYNz6ccrrp6RAKeCSL3mqQIq2fJdtGf4M8roj6N5TqvFXMxQibM+n0Dd8
hOXjnMgOOWxXYfaX9caQUzfAHSaD+tAUahBNOu+JlaPFgk1py0cNYytGwu3X8y130c52/RQqWb7G
l1m36scS4tgye9VqDLlxdrTiYeh4/giwX/wIVNJ8jIQ3PAsCauBJkbkcX7qONzibSzpxrBPqZSYW
U3pli/iTQUps5GC+c8d7A8q6GsWBYOJA2dxR9jnnqwlAF5zPhLSJVeJ/KIxuFyrSRtvfOEk9fMeK
R4E6sLDusAbtF938euh/MtY1mtObEoiHp7JVAFu4crUKob/AchNUD219tNlqSQcVzw8GazcsEsEa
dqVzEWpfKnneqG73NwKO59hNh15PtyZafszaGXT0P9AbJeH6N+q3p+k6A4iMOrkYORD14Kgy/1kf
86v16XsLd19+83l3blSHN3+Ez8TTXlvDvvfEuyjmM1jdMR5+5qyDbbN/WQHtrBH5+FBbciaoD4Ye
VHO+KXO3wsS12iXx+ioQ7rca+Azg/9peaIzpqHwFnZDOcqXbQBfTGnBzFw1z1X20E1cxZZ80Bs/O
9KIDo3HJrixA7S8Ms0djI0Hcu5J5KOGSwiLR4ekFiF+8LCh66iT8FVz4CahvZ67vgdlwvRvMXKVu
jHcB9XH946eCMtSykCq0hJfLusr8AQ2izWnVin86J1mKPOVdOmJ9sqkhcOqvGtcJoRNgAKkZM490
OH4V1qniPkuMRwt6wiOReM5TLn3PrntGpvwDIL25RGcpGeb72jSG0CKrEjWlR16wNk572Adf2+yH
/vuUG0lJiV5GDV9JobEG48RP9E26F/YGq/hmUSQ+bfwt2f741HzPs+UQHbOfc9rr/JR0M2E/RTQG
4mw1jOvJBejI+XGx94KE30CiMGlTKzjOR5kzAqiM9m73LSzgrGroqB+dN2ZPMprePNxo6kGbdbtY
Ih4JPb86Jv6zB+h2CPbRQK8vRrSsp8lTe/ro90rKKGKDVEMeItG4+Lp+nMzVqH2isyFu13hcTvzy
FcGLPg1bpt8PBv2Gk64hBGEdW/2Puyz3UfIJ6OHBa7gWtGxsYP2GQtz1fGtlQ1O3DcX9Jszql6f8
A0f2ceAqWaRUvRAU4TjU2oPAQWCI+ptK7VBkX0HUOwXcL3hM7CaEhNEDIG54byVpoS/DVYKvzyKI
H10rMPIWsUBEV9iL9ew9gqKvE/srSNw93mJTAnBfozHpto3kwAQU/saDduhYAxm/LCMMw9HzQksU
ealUqqL5IpCchNe7AHp6ybhPpR5XB93w7cGDHQW2ySPQZskHQveoiJtH+IbjxUYa+L3J/LvQeElZ
MT9M0pAgPXWa8D8vRFTHph2EKtt2PVT0XTSfkP0/5QFynlTTgrcOFlqcg88NOdn7qGdmf0eQDaHY
e7TwDvLw5rYg/kj+4R4YoETuFKxH0NXoEUbX/dluydEcsQKpEBKs3lLjl4Oh9Yq7KHH9hJ3l2vD9
ATDLHtpdHDDTyAE2PrdSiOVGQIz4wc69rodSui8pPikFQnu1sBGsks1dph7noqhvh89AXuf83c2m
DdwHY2lS+2ybmb9u9o9LG0KoH/a9D999xX8c7ajAwObq4WR62HRFYOvewZFooejmSfJcNXBnJOq7
RMvO3PVqMdChZ4lztwXVsC9iYQ8UDAt02AzcVhfU/wABQ0C5lMOP1U7ioSwxUcpIZYXo2va2muk7
xv/ZlujMzn9N8+OBuW3u5H+15obFQ9h770+zotlwwzq1rZmSP88mDmNS/GfAlvMFFcYUeVaxoqSA
Z/xhEoPFpDYPGCgTN+iJDEuNtEmJSNF0iqBbjDaDujYATfQMFSHqflh3kqjmpDovUo+rhlXEqLBU
3XRpUVCSgNZMIiDhcXngaenwKppHurM8Al6sAPnc2ZRZKn8dxwxivDVZjT085vyWmNLjYQH/wINK
BenSHWWkrqu9i9BQy1yLjQb0qH+gqekiApXFMMbx4dAOZHK7w4EM24zYEzyUvctcPRBxIu5dITvA
FYQKb2y6UdxunE5jF3wGEu0eJLrC4FWVk/dvQuHcz+i9g/CuZQkPd/ScBGFU1k3yTpO349ATUhXN
++673oSgxRoiEiLDcxxRxf3MlKj6CfXtRDw+0dvpoN7LOqy28hgGH+lfCsjG2LGn1b5eUakAP/N2
hBbpBaq9/9oPPCWNcmRYZM+sFUGMyqQL9tx3qC3T1F88DJrLiCLgdQapzw/c4vazNtf/wFxdCmjR
SKlKuWD35PlRxRr7IX8xiAUJkL/Jv3eLSGNbcyoykKcIkCRbXrAGmwmEpg5+IzpeNDBlHfF+DtM5
zTRnUqoXUqyGr+YGv2H5sWZxOxcWS5GOWTvv1xonJT2uOkxWMdvlAX6BVF0g/nMxZEJ92DkXbxpH
t3SAMd/CVPgZfhkGdkkkoxiBbFbKQrZmfudH1z6Y6KiTYcQ12tHhh9moOQI3EHQj3/IDITvdg95m
c1qnnLx+41s/Avvbr7+CgdbJKNR4GWfwI+vbwZFxFy33OYGn/5jC8Q3ChfIce/1Y2ITkS/0whhv7
tnt/OQlUOtOYuYJswVT0Usku+M/dWgbs6Lwf3up8FmwL+GSW/T6BDMGzZW9lhIuUYJvO3ks2RaQe
Vl2ikMtXmxMt9p7f8rjE3LBSiKlxiIpXmWHUakPK5/JBK32PsFPcI7552KIIr6u3apHPCG0IM13D
naM34DyD2+qXri4tZOqFuaSZh6BB6dASd63L3RoLxMwF0BTfJbtM6qbNhOWj+Ku+KiC0EhwbF8+z
/dO4kzmU7HjPbyuRIy6kfSost0/RnR4f4A+KvGlULHpVuZHNlukQeYvAtNpV31l9hwI3mGyew9Iv
jNeRon1yvO1SUCafXqdolBp/V3MGpvP0Fse22x9kmqmu1m1OZO+7A5urXTBSDV3uKAiFquIKV7P+
rLrcIW/foFq4GtE+caROHMZiO0HOrjgsb0EU1v7BpKGXFZ6ggf+iKJzWxHYhiG2ZuyK3ol8SuFBB
Bkyzfd1IgAMTElm60KaNb/km7a3OJjRSXGbXEzhz914knvydVSir7kKCQ3Gp+Hg8ARou1hXxr9AK
8dbBGQDHhmU7gVv0B5xO1e87023FYnduCjaZXreZmUDVKPu8iHXMcNDkKrXXXUZzAQYhyUYSWTUp
R3HqRyR6l5J41i6PsOxARd7m+xOt78I0mAzloNqVUO04LX4Vq/fVMUnli94ig2LAE8mNppJ3JNOj
B3d3nxsxGegTCAtvHy12x+oKY8SGwmY7orjLTUI0h7B4JAsWRj6UxoCSxN28ztZxv294SNeIFMCm
jtQYPdkc6S3Pet3YaFBnfni4DB0Vnw2XXGU2VQMb3tEKzadzr8U0inVRpZJVneIi76rHLZD4tvn3
yIMnsn51IWyWeYOY4DeSZUujf2jWTR6KIfl0324jW+DHxZaNwfkrIXjpJ4oZ9zu0eIjHMKuGbFlw
zPUA82ndjacQ8MF7nvpTQZH9KDKe/mDTTwHZkaquuJ8SyfG3ck3j+hixCDbsBtA/Y/BYIKzwh3xc
Ie/MxviL1Xo9jsu/rFSf6o7+RMvA9Y3bWxXAg2pnJpQf5UWGuonfzsC9MOwjX0JYa7YAe5WI6Vjf
4pxQ/qchBq13XC+6ZthNfUH2SHUZRLRRR9VwGQwYOJoBn8MWFrloDZycicd1wNHji0HfMHk0yu/Q
5ddndLovrG+jkXHbk/3PkElhELe6hBxWYItJZsQYZeBsQb8uFUcbufiuSk7mOv4XXVi8/Tpu1RPm
bxuGjdGQ9+ZqwRqI0lpR5KZogLGi3fOcFpFBhwpeZJZKlJjQ+OPw2ZPbjf2pIIumfHEXi/HE6BMF
ItwCaPLQHx94wStrkujYhcpCKRG//LbS/DAcjj2dGRK2Juu8B1nLpOTq82i2mspyeKE+8OEcLm19
RN4IpvJIvqlu2NI7oSHYlYJotFZ6m53K8jVkA4/5J7+spJEAIvnzA4GLhqWuFisQr/IsSu7dU+0G
fhj/LGn4VxRzCOtESqufzdzkL6XXM3Z//Uah7f0TXmXfDAy6ArnbHUixlQLcg4rUgnTSY5MkEZOB
3vpRWkQC6RviSbL64GMAYCUUVSB8UPDHQlrK92mtZS77XVONnMkeJtR7pgxvWz5LWcIFJo3KVN7X
pQ95twMQf9FWXzSWhyMR5JSUbn05oeMEfpkp6ha6x3qf3o5wVxT5F7LAbNXO93+ry8pgBXXmEZti
w96p+bT+0x+ZUqWCVi6HfPSm4vJV0/PXChHsUbH5dWw2CYpQ9W6+SlQTo78qNSJGw1KUMfvh6fCm
61WUHG4QaXkuxV8mzZXwXMd6JPtFLcWs2/X+aau1fUpqWWTqUk1x1WgJhIQ/xEUCIxQj7knjNbEu
J506OKvxKjyIpCD9U8cp1FofuoeZdmGYb5cRMaNcXbvucmeKzsxleayKijvsZ/Bw+HBuqF6hMFhy
1fbGzMmAKafNsneO/ipJVwEzO48aydGTKDw/W0MVMglAGOHjIHX6Ad0DgmkIVzXFVedVQfgnfUfv
etihM4lOfOJkdgoj13JBvBtMMPMN9zLzmWJ4Hsc1oDu1LjWiVvx+nd4LTN4XeE4nBeJ6zc15q7uu
DD2pef8fnodQrqeF17kPaPhkzHUOZpxtqAHboGc9YtfMNO4YiYB8Ju+kybyvpA+TR8O4HTdRg/M/
Vtsogei0qEAmgfEfbrpK972tZcyADGJdZPo0sh5cUYynKvf4VMDtiuTl6vCv2CKH5GoRc4O41L6J
fpfK2baOygKxY6r7rqYX9IWP/dZyekxCb2ZwwiizRnEVWHkvjRqPDOXYGeAyL1sZPyEeYSnjwAi9
U79Vqn77ierYWrEavgsJ6JyiCvC5BgxkaGICaqueSUWfCSI2drEboriMoes5XbgO+wcI9V8auIAw
HQ5FXIooR2TL6izPN5Lbbj4vrVknHB2xSmnXUzUXvjG8HAzBKsJg76l7RbK68NshztzJ+oD1CBKa
C5DIW9C9AKbYaQRUQ2sl+g68+9gVpbpKdj7HmZhmn2Ka5JZITsdjo8xqJpwfymrLZKneTHZsiAFP
WaPMmcEe50r2YiQqnULaY55KhwchQ5M77D4MZlC5E7z1mn2OXjBIxeB+0gQvGtI9OM0YvMxYagPK
PS7HNrx60Yd6drzeN267hiWDkHyJKy4E9P6JiFdYXzJ6260vRi8GjhbgrnBbqd6VCVIgcWm9f1kA
5jFnrHnHEEcr9sd/Be55H0sELR5Ic1ENRoOgV4+WJED/OYGzIzBKPl3FDrQGvnfAb6x4V2qHKDu+
a1GJ4rkfwPYPgcCzTVOoBpPnWs+6L0UcS1Z0l0/4l57JOtrAaSgXM/IgVWuOpL1MnHchD7rq12eI
KHIg66fx1lT15Y0XblzR7SzlgkZK/eUvxRNplcgRfiMbgciMjgO1u4khpBwdkFJqR+qc7dEfvgMM
1/tZWUPPMSt/P9Vzjk6KnL1gN0PF6rw025tm7nUAqA+VfKAWhZhKrx2T5ZIXJbu1MRHI4EauYJQm
SlGrWk6771eU2ggbMbDVXQttTO7SKo0jXUfWubArLme1p0lqZczxrPhOPHGoA8MvXp8tvxFj9/Q4
Svc/kofMKkTRucfsYpZSc8CGt9dRJUHkXU6QQsq3+0QmRk0b7/dbL8FoT6BVx69O6JfWHwrxF6sa
5jNc7pcPgsBBSqnvduLoOfAXdbzJQntPzpgfi4Z4NT9wkO9zY1zooE9EqV1b0yD0YJmwxiR3zz+W
Wr/5Xu+lzqnk/+oZJ+Mrsc9lqkYy3v61X8B5laEoAazuoJCmvkS7jck1Vh8MFOVyx/NAmLZRTj0Y
6veWwwKSr3zEvKr8mupNNF2sVxbSEnU7YUp8WQr7CwQ8U+AnZR7Vbel+mteHClMk6KruYG7jizca
9iqbnKLQcgYhX/PrKKk92WWSIpUN/HeP1B6mv4c4eUn8E3F9BS0BK0GB3zos7++ibWymerPGp/8Y
2Z+6mX/i4iec/7S2arGv7PoCjE7wvB9QPzPKN2H3d2FKDZ6DC+kUnXfzbQJozAwCXtuHOKEeeEek
tS1o/GL+t4uWj+wjfXmi5jYbNkh1Q+MXK1hr9fUVPAO5WPxqpI25GOKWkq06G1N56y/wRjGfYQF7
ItTulpFzXlxuGiYdU+6lWpPRa0QbcDVv6yFLW8RsEwfID8Gbhy3s5OXrI8+19mG9M/b4UKGE0cxg
RIZVXyMf6jAPGfRGXlU+sQ7V5NcBcKmk6xAyRL2ig5/7JsNTtUx4+qgkkTPPCVBqbw8+h9XU7ePz
2xQ6qZRAimkrRHLXdcTWX9XplJ78bAkPMd45FCvjhgb3TqfxiGl/0FOg8Gw+meQPdSbGla6bviRW
uls+xPDzwxtELjIf9162p1gFG52L6H0wNgQyO6yiwKptO//dM1Aozmz2OgaQphdXnDNfMdGGlt6F
BDz1PRf8uUN/O1mEARkF8uU1N2LGmAOYogVtfI+e3iSu91vtpEY56jjYMvjiBiTxk1wU+uEpHk5u
PGKEA1culS0rBTpYcrWsyfCadECiZh7Bqwrjs2+VmJ7G6BKVkAVb7AqLzESHQcTrz2eYqWYc6u24
MgkuRg64on288lvGkTlZjaUhB7ozPlxTk6OzlEeC4V346d5Etf204sOhk+vPlqqhnYjinhCYl4S0
Dvcssl6ocny7fLdiT1E/Jj/B6CKlOD6nUJOHf0lC/olQbRXmfL7T3aEeTiuibuh9axgkkSCOn763
GoatjeaDiF6vFRsfPKomA1uOXJ2LqWbP/ayIylT9ffbnFEtOmx0ibwx+PLjHln3TomfPu5e5YgpP
Scp4L3KlRo/eulaosquwZQM8FdT+J2DnBsVU9TETgsALi228hIMNADeufSiI5X+u0tUwAKUbjjF1
ZfMu/Q5/4KLv/Ea8kpSntMO2ukp1aGA/to/BSAo6HnxXv+donfy/0Zni8mp8CevK+KhMYY+hdTAX
LWi+LCJyXZklEJLTGfxbT+HoiExPy6tIXwq7zjDVUSV7zAy/rSFAUVDpR9TyOrPGFHNP01SVUhl8
ake5jjJAdXvQlpMc3l23I8Ib5xGj9ZaKqHn7aQOmUprS85LqELsPM867vIIhN0HkRI31vxnoXEuW
SjG2aMNEIYLL4J4iIpfU5g8YuO0kkHWqvRrjRewhb8lMBmU9ih+/qA2pLGOZtdr4OTwHrtH0l1nh
EQvwXCcCQn3BSMer6eD5FSZstFZorYGQnPDhnbCLVQQJFNtVQsd+7iBwtzQ1h3KI50MYrG/CWkpG
dXCZnMw7a++xivWFCja7qZHTVCidevXkZNntEL2JI/l4St/FefCtQt5nuJ8sd1CvdR0QTMAuRpcB
dcMdpflBQcC1wa2VgrB1Wm1qpOQ5Nsqrrii+XIa6o10q6rmzwquZ45+hvacYp+nTDozrwHFLPtom
1Rak8KoRoZloy1vDB4IgJz22HsE1ra18zNXPLbgeNKNv/gzW6GA6gT7MkptcXleFOwDRIHpZeuOJ
A0jomkIhOJS2xObumG/LPy7vLRSZ3Kk02TTCMKQ/ZITeDEw3M0BO1wsGnLRyj8Xd/UsB5/wdKckP
8jutUouRcbk/rsY/3fePy7XkvAWj8F2IanraETyBBzO9HwuTAzyBA9A2O0Vdy/6ac3ijDMHkD59L
D2A8fp3AZbWf6GtBOWeDnFW9IazwX83SZXeSgrr5SwNeZ+Q8DE+qOh+L0FtiEGBmdQ5LG2JWjtKc
SkK4PDeCidnWfmi7MqdQfSAKLkAugf+smII4/HGNoWrQOPEDW3Sc1RMvGDC3IFG5jRDaxrr+WEYT
frceAsOWqhtYBUT3I9Ci5dlzc2noudV79ERAoALobCY/EGuQF+z+KfD44ks0SZuGuzqbotBUfZEv
/x3Dtyczr08Pdh0EFVLbIC26vyAFg2SjVzi5BB6BKcCS/v5YnKiWyrhJxJT97pzkLr17+ju3kHxq
3CHgSL1zt/dsO3IdFFlav78nLxd1X4woU/yqfN3HhELCDmBcLIzQODc88YcQXLkqrqWa8lHY2ILk
V1+mrVqesfQ4VdZjIKcFwmmU+MtNM9H2oyB3ZkODWUPmNItIgODRbHCb6xooII65VrBIYQx6/n6d
7mb7sshs16EF+Anjp2l26yhVGtg+IfWzV4xyVZKuXpOvPZhadnHFSKnJUrP8S/bTjY+0ILLbvagf
3pwNKM/LKzFNuiVJMuUHxlzlClHc0sblHKhjK3LRdcAD9Vcpl9WGLmDRlGHamkQPJ4AhPBbx2ITY
yx45A1g03HcWgv+IqoTO2AJP22WCd4HocK4CEwH/tRIqrbljJUJlEbDXPvWwCRsg0kSocTN/lIap
z7f39S3rR9IxkuK8cUcbx2XQwks7npfcsgitSfl2PDTV77BYWvgl8ybXA2i/D6Dt71EJ4C5wGDqT
k5QQFVbn6FYEfbCl5cZ+gn0driFlpEIccM0Y2uHxwHx2iN1nHE9C3smkquSIKipTM/ImwU40au3v
WOdKo/Kuz0Duqt9mjOeXpLHSqQ4qLheYNN3Q3B5lrESkBjD2R3xPGOViRXo68TB+J1gbNrNw+Fem
s+NZB0I8m2gWALzMyWycU5VNovaXG1xlWJqqNdnnDscMaHiSJiL7oIqM21f39i1nWntpS6r/LM5B
s4ClG3pmS5xsARdxCF+e/fhqMZZ9MGNQbByY8/jEx8wN33V7dfx8Cn0aTH8UR5n4VaBHySX//pv3
N/wKqiXX4t0eA9CjR+FB8gGnbKRiU5GgWS/ei4toY1qlM5YlVf2gV2n2q5bNEaJeHpY7FQ6k0waB
hOtMNE8y3BaiQoxCc8RHTV+6xRroIgLUBqKag2SQfCmIyQoHsJuQOhJdMvVIzBG2rr07HFTQYOTC
HSthDKlqFdQmL+sS8JhzuYdEZAvAQvsPrESgKD1N84HiXEuBiW04An/Vm+LFaivqAaYvSkowraY0
Muz4l9320f5BF9UT9qNS8566vLP/jV9rmLw1rK0G4GpkFAkEB3IrWIdK7Wb1qaqaGYpprbsfo9wg
U1RwcXkp8sIEVlsAhJMdvZDsXPM581iD3LVGcW4VKssbAmm4gMhpkTGKl5wMyUv7fkhNgjMQhM1S
k+Ve/v+wEL+FdLEjYq8qDzgcycNf79AlN6UmrEtKIr/mP5swH2N+pv3gTL32wHV0i+S9xII4pbqF
RFPOLYZkKQXA/i+ONc7R5htuYlZiNoO10qGf29PFkdbGZamqMnfeopDmSMORUHBTsqThlVzRA+Mu
OsdjSP3xR9hUUFJmBkjXmDDDeu2lq+ueVBCdOouCWh8OS1gpNvRvZlAQC6EnNpl+rQr0g5AvC6cz
wdhN5ixuCMx0SuW4BYT6ZekSfU/p1jcVA5TybXYbr3seumWG9EXLkjTsv75B3GzmnKwwThVN63F6
oF3IfU9eSzJOtoCpwi+vWcaeCKdxYOTdOi6YKGU9oefhq8FHujwwJ3wPtRc59qg3hEU4DrBGUjjb
tZXXsPEuz/47XbD6mxgL6F37ke/sLXr5vf6AWYcmjFE7Xm7T+M8P+zz/wCUirB7lnRw71y/vxnbo
KHGXJQjIIrxUiXqFrdz/utouOMDxKLk2+VTxFJN5MiSB1PojcLFgPhRCXjWf1rWvDQM2W86GblIj
couNgH1/1S4vVyZnjlauDShU/x2bufUh10I6L5lCkm/uv3Z9uSyFYIY3Yxsyt+o4UmCkabzSucLG
oQaHU0viZ0++LZMlSpSDGE6u7blIeTcZnlWMpVPLwhvh+/DBfb7hp1fc7opefd7fhKmB036q7Im6
XKVivARCkODGg9/t0401k1ieCXNCuJHG8AV/uMWwOfAPWy0D1oIFEtuw/NpBOcyHAVHNjJzj1NaF
9oSi8lBDnEKUOkYJdeVDITRV5YMOBKh/QxxeM0dlorUkaexO8gUU8H6/auOMCQ/0Q2Bosi72roC0
PgA9jftgkFS1biMoacHxMhptehCPXGpYIUIZO/AmFYfMPBxloWt3fwPKefyoG+4cu2osU+at3d+y
qgbA+08d03meq4BMK44aVob22q5IfsaSaJLZpTdMsUD3Kpcrid+KtJmIQvnVbZ9BQ7cYX2LFVOuQ
gZyw7L4tmMcpyQpH8MacjEPWo9E7xK3gjhVejXTPg1nRTvIL5fOxRqeNOve3HTh9vc9Le+LsZat3
/DkuP71pYEs39E5zfWJIFvGoIIewvOg9zwDlBB59q8d03tZtQ7Qq6gdiBYhcFf2c2jpBdFzjJ/Rr
qTF8KJ2qvzJNsPbZvEyA27moaV71P0/qDNMdIy+VbrMMyIw3RGTMIjmxERc5yH6U18aE0Splul1p
GDZgNUUJANi/GOU+/ahG925I3YPUDr51OMgrH9FP4vBWjSP0OcbHdT6PbY3ne0ZcxPyv0j/OLpgM
ms+nIFGmsHisAyDZS/049D0LVEl5IhgoyUpTXBjATCjhguqCfti57vuOP5p//9fXjW2lRWasZdy7
EHPwC8KgJvHtSw9yPBpSOWkmBii8ROA5vhTLkHAs9aOP34zMPf6RC5PKrUWlfLINpM3JAg5RJcVo
Vdw/aR9NOwSTebbsiDAWDavAItUffND6NlBLFH2tV84IZ2XOeeeNa8m7G5SeAZOqz4Qa7c9BZlub
FZ8OHd7eGrJ0DR3Ihpks0rZQo8xk5lhYCruH59RiVaDr/lLnIAnt/KDTM/qUno6OHT0XVurUisB8
8PEWLytUji+EDS5HSa642LPEBhNbAVghLPMLPWvp/n0YIj2wZprNS7YSCeRH61YS+AlP7lBMyWTV
Y2lo4Xv3VRHSG/0N4xFY6TSdIelbqoQ1S5Den86ifrjBa6GYHO/g6a5oE9GROlWzPDV+vUs4FERJ
PIfc86sQ9jNF9EfMB/imCsE/vju5hj3GbxCIHNKXcacbwaxL8vnk70QRP5kWVXU1JCxj8zhmWnQT
AGP81nI5dfLoNaDX/eTkFSH+sp0ywsQ4KJvsVAKjnw9YooAWGdvwlhzrnx/nhFep79xox7IqeMGl
GPCV0g9ys0YtFdyh0WHstCzyQsBMA1sV1X+WVhnhMlwwa/lnACqoC4yi0/5RqTVs37r+oSHrySiW
R4mt8BgfiL9DmVfBSPnjBMEvyii6xh2fxLbwjiLnNhSfC+sVF9ECkubrWkSQkkGd1exfod4cpPFk
KTSV8p7UVHoSk6KMr03DSkZKhHlDixXniG/MjKmoW4WK2bzTuw0xIinzkv3ksbBcZAISDOxzJqmm
cvbI7dueUiNjD/Ygl97UiqzLq9hftPiM77kgYOJHWbVOswbmYkDM8OODwGns0MANoWqwEAMCBbcG
z7Ml6Az/WuUOMZG3ESh7jFI9lmt0s4MmpqJMWL7on4XAG+yDEVpQko9j2c4Ul7DUClaJQ4/JPmcq
kZKfYmBz5SaLgcxdrDIz+pOiafldPDYFd59jo5FhwW2+g3rJ7+ExmDfUcKcube+XMR6yIRs8BX8I
J9GEGTNsQ+qZQ8PfJo6saZ8VwPv79ovYICQwWfvcKE4pAF3WnPVSD9IJ7b404pAKBlhZjhP89juq
dudU85A2m/hzrdyV3ck0y34zShtm2uIVkMmAlDMyCu+JlmAdE8fwzIn5aHyOzsh6B9Be2dZXahxw
LkFJiOJ4H+kis6YVCBbc0hiqFCq9j5fujPH605o3rhidufa68ANfxrod4FSWacbgLzs1jnRBAiGc
dRSYMw/WV13ozbgGB3dINLU7BJU2CKcx1981qijacrKSQbBZpLLl3547X3Z6tPiXMX3A4YwIh68E
7Xg17m2bmGdq8nuQAyOqM7dP9/BgjYWCH+KjWzGEjtHcpTRBNWIxsl5NW9ZNaehdxCuciAg+eLY6
ainOAVNZJAlnppL27k+eVCDLj2ck7uOLKShkhexNLtoI3Epx69aqheCNZ8OIJ0wNsYPDgD+xWuUS
X2MynUGAFbbyHgs4ilvlh5aYLEteKyLDvbuOspWAOBs5zUZCopfjIRpnk0X+ylFxw3ABqMYkqnmj
1up4iyEfcUJ0LmRfRH3JhYewWmVjZit/bJ2X5siSqlOMEpmMUrlyw2p53KWzXYUGRuBkbsQyq85P
XQP26vsNmuRVE5g+zepRh8Uj4Gjc14t3sEAqPttu0UoyaZmuG4lWVt4ZjdAlxpyBGeAWm3agsQK2
F/ZTnlQm8JZy9lslhv200HC5Y9ksYJciLgfi5Yu08L0qShx0Qkm5Z0LO7d4PiwtCF++tbYFIjY6M
AKlp9F7sKvn6akUL5BeNJsZTMhV/Y5KJbcjnwJHVF4SzTzCkDefyfDi8uq8JOMlOIVIAbhQQLJNT
f58P7OepAEq+m/U5CFolSbzzppV4QbIu5ETLClew7sgAMLVVf3OwjKcpP6xgVLWLdQqO/r03RVR6
GRHG7FDXGmYQWSfXTlIP/U/hZTEG+SnaDwU5p5RnTEckSBoE8efGbj7vjRS0Lh2OqSu6l9tsdvV3
4/iLN0/NioNkIPLKPZqyp8p/7YrBFX2Wys4u2VQMhGhb6oouH4IS48qvnbShlM267yCXxr5ab3zB
bVScLJPa5QIhLt0KUtGzBWWT0gfAspQ3F0TV3Dri4JuNGBhN7HDD2laWYQJoDCeln41T56//Nc8u
ieeorwntUdNajbzvPPBkpPoSFiLystyJ3CcFSvjMZolE4YXAoyJxMeX6cHtaXYue4OiAbSKVIOQ4
Qq/x3NDHyq/fix3+9P1DhC3WFrXFHTiozVCIH4IRm6W2+jGyZ4VDZmSZDhWD/RJJr8VnaS3ZbGux
IN8AXZ9BK1EI+CD2KAwS/tVKZHWG64J8agAMmG9zAgoq+N9QT4NVAOzqSfqoizG0V1Q6gYV7QtED
04f+CKJ3N2x7SNAVeehN0vdxmkG8/FdD3JYlo9ozyk0NHaSz01q7ran/4A7I8brHGxLcSJhe6vS9
YiBJG3KqU9RM3VoMmAZ3E2VwqM/T3jm5JjvCPscwyZpVdsUYgc6qWkFQx55gwiHITJZchVRiz2u2
UD/uaHDN/XMmqTysozGnsn5aBwuaSi3tGT3NViSvWjBrr/pzPanx2RHVQJHDVCkK5u3XHM9+9m3a
qt5WL6BG2GUfsDrolJ2TJnUwH/Ssa+bY7eJ0TViFcRdh1tyUDriOxc/DwQ5VQrNW2FNG/hbw1mM3
YfOoTK4IImJvZQMDcSizQhjcFsvoXMGXv8ps9WX/qCSibSa7RmgroHH/WDgn/A/6HggGz6IVK0kM
QdegiSlvv8WRr5aHmOJyxs9PkI7P/0lEQ623CFfEDWQ5SEirRkksdIyAJZZP4ufYBLEcA6X3dXq5
aDZ9yBWXG6j2liTRB644OhKYiICpNempRDPESdq9QT69CxTLrfUJEvGPbIT7HzLaADLZ2HGeSMgs
XMHdwTMvjYs1KlUG5Jfkm+KBRQrPtAJh3XrC2wzRPinNY2DO4XYjKnx+yaiink9yWN6+0S6KMJiJ
UuI7hexAX3U8vab/6f6JMnil7330kqNTkaILU7qmvZYOsz4TnheYwmI5N8n0FEkQ7+xVUDNxvmDW
w+KSZjcU8EAbFTIgZr/M7b4i7q4KQPLU2beFpWyLYbL8NxjG5Jtr4gb2qgvSvF3KpA/tdB/SGin6
mE55K1GALaJe8ACcSXq5B4PjKfi5/p/AS3fAkjJbv8/wwr13ODgWm/bmXAiijYGoIravk5v0oajV
wNNzwnwumYLjJwd5+/aEnjN3Cv5cM/b/MtsEjtjToo3wEWkfoA0G9CWhZPnqwmPzpCqyXzkaY+99
RNY6hPqgYAmy16Nq3HsOEpUFY2dyhxkPNvzPG4gm7iKTXL0G5mQr42qp/9370qSMMIuE0MWTRCxA
8q3iHvTNbSl20F0Z6LIqkd8oreUTWyP1H27QgROfCJVYDe049CFoKampbiAjpCE5r2ko0USAus3w
WzvFAIDMOHqPTzd5wPnQcz1CfJKPTEP+9Ahwymk6fkZnFkpOplSog4sbS5PujU6HxOKC9LlwGI48
wvZHMn499AOGprCNH6x/YHb2pvsbPspkm3v2ghwdaG9L/6DTSrX7SOMrPdQxZbORgUuyWnCoABDn
kPu8RlB3LGJcsbE2Jx9gFMea1PQhCkqUD8j/t2biIyBz99a+A6tjV1+6vCVJ+BA1nZi3EOJne+Mc
3d9MQjeZDWYHwtgnyFdcLnKfWQIC47kNUjlN/u0lyHXfJd6UgqwJnOFrRAvTUhBd79Acuwj42KXE
t0M80ruwTjHiNLnjSr0KV8Clsfh9ggxYXwCHI+PBMB+i56vE47go2Gf9EZVeomPdUyzHcb1Q64oN
iQk2JT6qYfNnjPLqV1d4uoUTlu1/1bqCZq80HYVQx3ggScqswbC3AdfG+CeaMueVspkNfbIuJbPP
A924D+QNUAyBzD6xP1NYpoNQ/mokKHP3GIS2NHLYkeu9dNf7tVdzmYdWQJl5GnIX44aeW6J/Z+d6
KlI+KNVjZO5s6jJmWULiCPXs3FJXIWLI2Sj5q4nMTav0cbE/7S6psRBTwvHGJ+57k8ugkG17McUV
DSsEIoUCVnx/nx/mDkzqAOP7n5RARvdA21VVFrwS1aiu0ShO+2Gqdbyx/VZkJ5TcvyUDA0NWFi1o
zxfkB6dswSZk0+3SNw9xbtyRO09dd8mD0PJ+/EuhSv/ic1mTDAbl9YyL26YIzyHZNS6E5biESBQu
SyVfAilaaa6qf635nEtHM9eChlJFTVvC6Zi806P1yCMdqyNDyTs/ly8/g91R2tQ2sk1nY5/MLHvg
4/SDMQVDRsXJGsN/yduNS4eBs9ta3G7Rf7RdH40YvlR4LTCpJTSzadPY4caX+CDSV2mq8rpy/Xdb
5mZ3zGy8Z/jW0SbLjkfJ2Y+hUqgfOy/naoNpKl2qIQdp2+CNX/EP7HyUgfYGgH/exOFWA7FTZBqV
EavcHQ0PfFWF+ZFWHtEQZurNyRWNrZqCcRoL/95uiv0jq2KTO1vGeWLJlwkjGc4FmyyKK8joYqvD
aXMA/WeC4lUy/5wlnmJlRs16fJOf9cwMGsouR3sScly3P0msFu2V5Vo7eS8o6x4V7G0fPPOY97xT
13heLKqtFSlL76Wv77pjtE84lcVHeOkMb2wmFEZBoJFkYCDEwLgFM4GAp/+AMVq4x7EwjuEvtV+D
QYF0gcU3zGHAGrzhPmzhKbWI6wFfwLSOimrq/0/SuSgVbaNPMuqYVJbpWg1KhjIvDCpVAS/klMY+
FSYW9WrOgcXSl9e1M0q4jLUkyXCOCby5jvtcEn/wZ+BJiLYnHfjBrk2EfOfSKHtUvKQuAqU8Gl6L
d/V8Ei2YF2rQ7Z+Y5CSYWp//+94Vlaq3+T2GpWeNl8WVrZRze4Ctb+1mfQ9ZHv2DHbzjVuslb3m1
uyA21jAoalaJ0wHOoTeHgNhg9FykB8FGP9FOTheswKqFTs9J0by6+oy4KYRbFL3UfYGMR8aDpJ8J
L97DWZ0k+0s3XS5zIV37p/tKUAbBSxIJfMIuTuHV0P5NlG5PV+Vl2SKh238ehHu/8ncQtS4c3Piw
kVrWUukTsfaUEM9l09PPj/+fFAoCt0YTvbGGogxka3ziHqTvoZQmPvziZaMNeb9glX2bUrodwSfX
eAvhuW4oLXElMhkybKcy2cwuC8AUtFENy0NYpIWgGeGXzhb6lnAxr1ZxlL9U0QmXXjGWAA+qL/EZ
FpAXhGlh/Duq1JPOTi0m3IIJnjRFSyCn6wzPLZpR+L9Tyf2KV0+2GiEt2unzAIkCDraIgbo07la7
vfIPbcRLU15zFHQIjyOFXql6s/uMVZ/uzuZcgkvg/sszwQEPKISTUq80Newkht3GsM0XxmcLxS7c
X5EkK4yvW3IIFrTSSy/odN2vqHwmsT1TgL9g1pWKOjX1NQFdFrOgrtpuJ3DrX5TgRpMNiY/MtTvW
xdGnNZ3CStO0FlLD5cvUw0PisOy9ajfwhI1uV8/akoujo3X/oHQN4DeqkbHrSgaQCfg3YgYBrrCG
N1kTrF01CUoQKa16V5evKyCL/w4Y7i8HiQqnCVsdMFn/WBUrSz9/krjsPWIGX69Ubp33az96+owH
5Tj1GRXPCTN5n5IaoKp/6aGClrUt9dFhhpgPNaYJVqbieapoJiqjMRBTrJiTnIuW50yTwHSk/OT6
TxlZatHO9aWEAmv+8XszW5JpUAL9oTwOaUV8jrhmj+kWlgB9PEg13WPuLn70zLVSYdtRuSKIlJtA
ROSiLf602WWw6X3BbnFqpiVA44qEv0vE72vVqO4yeGnrcsN/YJdKQK8e3MNewABRDXwAyL8FTOKD
PAaAhrhTHH88K2DhvX0csZxqd4ydu4k3DCJ+6laRw0ulFSwLPCUt3YTHZyFqyXjAA34p0EswcFm7
5ZfXUVOjlQuiOp4zqeOZGvmUcQc7qoKjsdGohtOLG+goWhWROzqO2KpgrofaEmfPSEXgckpo0i2g
vmmnSAW16ebVbx9A/mempKHAgBq8ReAKCx3bkIiamoIDlojgfea6Ipig5wD0mDZjTiaMuPwNAe9x
ljbI89f1ErKy8m3cqesNxzLhGBGdnr3F/AIjuPXD1ZUKMfj6Jb7ZjtuGmjNYDnszfn8CvHauslRB
v/mG1t+kpTbD8vqh2Ew8iLaNs5ROExOvrBZBjW5PDn9K285PYslPCmainF9RYhJizP8ALaJQ49Gv
5Y3mcLA+5EXMNoknfGmnU0UEC4kzwjwe32NMwkT9zQQmBl+a9K5nus/rpEFK9EqNIZwRZv7WtV73
nLq5j9xTlCgur72hrIXxYjkzPDksmXbUff10Hz1K4MjIkAlcNO0O/9YN1u1d6auAmxPHoPUxpryo
X2yjHVb3X3EFj7mhDLrfyhqnDwPAouXxpPgTuVT7Qr4kCTanSHsUTRuKsE2+AOPdEcdWyAJlW4HA
hUe3X76OnDyU0yg9cPwmb50MGId+ohX0L62KH0sgabKrylZ/kZqaweuOWHbgY8FhJcqXvFjgZLC/
TXKXGd/P4UNGTVNKiKmq2q9yiviUVFgfSv5Y+uTbJmEck6VLOSeG6ZQyLsz1XucKIKdeyVlmGiUc
hsM9vkNDkcG5Vb2mSWiE7XF2kAmI7iZiFV6+ugrFe/IAtwOpz/z+srNoox4H0X3kkeOd2M+l1I9i
TXSkA931cIKmr6lQGrvyRd6jsyXhAfRZ18LRVg4o83HiP+ra3V0PTUq7Vw88qZtoRbitBG5/VRfV
hJhpwXn50HheBaAIwp511rDyGrHPjTt1rGVoUmm2FVEYY1oYlrHowOY9Or5L8cEYZnBAqkzNBbol
7+oxHtVAmYzGAoTgvTA+erxufZJz8BQ5N/mHx/v21vc0Ou5u+xBzBV28MK62b/31t/QM7PlzEAS6
LQOuMu3eJrajVb43moP+W0y5jCDywdboHYBt+6Q090939VLObdE17Br8IpniKh8SWpNcbb1l611+
c78d8kyy9tVA4XZba0axSlf7Du+fiMe9Wy/y7Er7S8gBQABYqD1/BOPRyUtcjX8uEJc9sSuCuwQY
VUKOmyXFfB28DPebdD/XYqaDVhtj9c0IJssLXtTqPpqZok/1lFwL5JUJIy/W0WFr8FXy7MA7u69p
nOzvwtwhVs+ruP9fCwLa97b78Y2AT9LnKjwATdqK07TZXRSf1xQsVAIOawiAmGrzxK3A0NWlFnKc
yIjZ7ggtsuk+v+lk25hCMbDVpn16jKIF7JafxE43MLOvXVRRvlnWx5q3bm0LOvvFD7DAk/F3WJUQ
QPZR8Rg5cj3BIZyElsoJNRRYoKpDwEjkgLpj9nN+AMk0BpVnQtJcRKQjO7m+vXSq+CwoW1h9QbGL
Vvr182p9VApuvzcD2wT6piGm/hpNAdhhQ53o78RwmOvBVWEoyBPIrwt2N2ob9MoohyCNZPlzWLXK
MNBZgStQiqq1ABf5v788d4ob1fVl25fhKW8iuQUA2hmc0lXQK8RIQ2ZI1VqQ9SK/wOxMWpLb0eKy
b/ZVU2l0cWhBYM1ojk1Y76nuvypx8jfnC1q2+hKsFTPaPXsB72Sx0Whd5rnm6NADRqWtE3KESi1+
WL86w+C0hnK4PICFgcxV21YW/e6rNXjFZMxXw8QPZFBivO3AxFFQ1zyWAaMlvVJ564wS0j/B8a4q
+/WX2ZhMSSu1D9z7peZ1EcNKFFCtMTpTbLSy+BqYngFvcXtHLSahtrn/Sxt8ONLXNAi+6z1DjxU5
43oxmJActLrUZIw6ljYXScre7QEmIAofz27L8PGx2wEggVB/5VPPvh1RlscUSBr3SB5JrMJG3eSq
FS5FQ3T2qTY8a0kX0MG5K4D9FOOEdv0x7KNbvFgHMgCASaf4Sde7uksNlFNbRW3ClNA9t79P1M2D
QRXxUROR0qZLlWqXG95QsYXtAOTvfeiqxOK2Svs55XGP4uXkuFRGfQuBs0Fkd/LjgsDqDbUFR6Tx
FnItsGjYK9xaSmExT5MlspK+zwYIE7JL1AT3NgVVhJ/h2yGf9dPsyh1wOntMqW5NwlnT3TBJ4dnv
+R/OpVULYUUrFRA3pckTn54rFHLywa2SF/x5sCKR5qIIBbyb53hXZIR7c1DN0w8yFfeB8n2CV8b8
D7dWvh/O/V2GUcPZ23tI13KoglgqLuVh0+gJfwk99OpRWnGNXfc2ic47FSZbzJ56qEPjaIVsp+uS
U+onUH+XSWDEo8NErHvfgLDvs3Ecv7cesh7gmZHD1j6IBFNb+bzJZWqlQ8zQIjUttAZTDq36I1ec
lhm4G9tFY2G52pEHjp6FM0P90M1kjtWV+oHPcagXnAHRRG1AEOhMEyuHAazdGl85KvkHtlQFia9V
MyRoqnRmnI9GwJus/W5XrIyWeh/++c+Y14koJHDBpKka5z6V040YcmFEs2+sD+NnqS8tDKeMZ28G
gU4iGYzsRUunfmdBzHf3Gx+WnKccGYuDARMgzTm3x3XVv/vJoQIomX18kfw+gWqdzQ4CHdi2+Uoh
z5MVBKcSLsD1KMhG7pCYTvMoaF3q/xy/7NJNhR2dyDdqf785ErDp3XKpwidg82ykiAwVHIWFniKn
qAaF/+DExcva/JSyCOYkDELpEqs73t1S1w3dhiWrmejamOqXx3RfYRbkN9pR7EdOLVxRrMjFMP4/
/vuYjOcW5UoSpW7uSlq0GA1SZT69N2qqeq7ie8+2fFrPHyD891G/2FAUvcLiCTqpfJDoZQT6oJHp
lZrzJiEQEGfP6GDUgMRuQTxVLe8nRTROeqvao3npouDhnNxeo6pFmHhAT7qbZxxNLZznUsp8VPpO
FV3zJtDPv+NB2zPl005pjvd2G7I3zQ1ovlDOYEbNAwygLRnSsr545aBhPbKn9N9DEPyl++tlXT72
ob11cPRhX5Oj/JMSFd8aXOS4ejhj17psi/1KRKgE3RhY/orZqF//zclal7Q773m5K4smPi/2Tpm1
zsVE2IK1+sDVIjrMtPGD7dzGJU+PYBqioy0Md9IhDPO++b6dgWC3IFxr7IKVvJlMRdSQAQf/Kzlm
2jT/RBti4lyYHksa7JSuQXLp+kqNdF3FIiOfcYRvV6MUJOCUFrl3gkHTaKizVLOQUiMSjmWzBxO7
bPhNwzdMsOwDxt9PItHxRdJHSGsJpjDuSIzV7HWWeVeELFWCWUTmT7t4CeyJr+6XBLIGzCwfiKVm
Fn15ozz6rccyJ94Df5Ct4i6lABjTOimTbTQ8JeVplVC+yZawphr4Ir8U+DmkpZGPM+tlgSdLOt5V
hXUgtwo11oX7H+tVfQhCOzI0dMIeIQVTbi4zh8KUgphDuxmMZ2Cn1ZtTw6CrM0BmkO7yKIvK08h2
L6l2jL5nTdq6IuWs4q7ZRoLJkKqiej0SbFCe/oZCK7gRDLVB6FnywK6Ny+YEZ2Dv+lvdJVDw8gJz
nhsQ8GLMd2aHlSLdT4yE63hJza/8BhKqf0QUIkUnRRSpuo/FMT9T4xIK4Wi6RfCc4or/AIIRV47d
JEHSYQiFku+ZBYb/Nt052Ui4eUnyzhoDKp+/6mfa47AoM0BAPWoGK1nBDhFpx3y+qMd2XWUT1666
ZHftL+xD4U21uYj6kwkBPRd7Qjllgg7cw/A5ka3/2EBHzBRacZSRWzDUGyc56Fvm7gALe2bxVAUL
BOU3NMyVGXjZUxQx2zFDZGqie9W6GNUPihCprlsBt60U6Ale1LO5BIGL8lChbGbfGQnK3io/4JQG
KoSfkgc6rv0UrGjNifUhjXWY2fKFLADGR1UDZce+BlMlc1ZcZ3gM6kC+BEtg1Gd3FjlDQ8cut7Qm
45uFZo3vtPMjW0SfwzbvCJiWiWQv+8Q1pKTxI8warjBRTyqerX/CHrC9FQ3gKPCW4TKJem7/MO2e
PaJWir/0PvmCOIkKdr1j+lxW/ebQVnWmLkR/GXdsQeUp3qxOw6SCwcsi8W184nAofv1eKaRzd9eq
p3lDzuTIRet15oVr2yYolfyjTcoaWEtN8+M5eq1K5zuAiecJwu/+Gjh9NeKZPDbHJP3qx1YzTZ/y
DQxJd+zl4ACtccYI6YQN44mlgu263mqIWmGRe80Vp2/u6pAIWt6/ft+CCCawBotCJYSZXCgwv2ea
m9nfGLqAhl7qGvB/mMt1WF3mvCmHOaJVkpsvDiRwySJgLbeSGj2auwi7PNSwk5AlJ6Koo+JMISnj
OeD0wSvXQtTEHBxeHhDIzcj4U+AaBllsoyxrRT/xf4WSf4m0iBoNVqQ2CNrb7EiU4wvwevdkeiVw
+8vCphaXy6neGjMszAoxH/PjY98PLuoxN9keeI1ymjdVsiyw5FC+GLcBoRmImosX9aHfVG+BWDAx
B17HhQMtR/0xqyVE/krDV4n2TTEPNnsNNUWcm9SaPJ4rcqI89al6ltX8ehaFCvMk9JhXG3ZT9nkG
h3qQOXxYrPeQdIyFV8RZV2J3iNY9MCCy8YKqJlpos+l9Ok/aWHqPLaREeyLLL2HfAAKCA8UTL5BC
Xp7sM9DZqVJXnA5rFZRcoMm2UQaixkJAzJzXe6maQjohLvxCfxvFGPJtS9XADVcm31uxY68Ym8NK
7oMDm2Ir5NKnAipCq1TE9w0F77wD1GcUb/SiqjyzhYluIvV4UyW3F7ELDqQhtCpKu+R+5ReXPU5A
Q7jtkXjm5MK7dtUqoboOSMPXFWq5pebbqdnmR17P3vzH0aDXRrkpJQZdWwoDgT/vu7gdNe2At+Hl
r5+EesOsafew8nij1r8vDX1BJbzFwtPZwRQAsMa70vp1v8P/G9p3UfZDTCq7CQsVdlSiZN5Bluts
W9FQ3LEh/Q5ryZv2zM7BGULbhxM7/P55oF5NkcX+dwg20bYzzsfIXz19rk1cA8LIBHCTTv3uJHAm
5KpU5OTKiRJT4AH5slVfQNTR+MOS2STi2vs2kWeXr6jj/exnn6E5zIxol8depFVqsZ2S2+r+bluh
i3v7k4iyFYUTh7vVxHAeqyVhntBFMOlsgkBRjq5FWkaQfdKHmGAQkTOL7S6X1UqwuLnXNZykQ4IL
pUnAz5h8Po6G3/LwaXahUKE1EFn/VCR7IecPnQuxdfp5tfj+tLdmBO84cNllgETxoq9YaofIfstO
ut8rTBFhsKs6VKWJTmsIJP2oZjhWT9KjsbVVpdN/l/PEQzdeKSMFNSU4BNrGirCOTPNeqhLSIwui
r/9u3DzMCQWCNPy92sU+Znz5JMlDBPXRY/8KIkISk+EBgZlQh2F3uTQO7iWctVUHuAO/AyWHwZwS
VKyFTTLG8pQOEIHz70gqYwE8GiEweyUG1I5bEXjP1WnJbvBBQ1InOvq9kfJMcsPRIAye/XR+Q9Zw
UGDfHalGbT7W7v+6wigqQYox5b0IvY2xjGcZwAi4dSKySSKgVIcIVJDQebFlHjE2VOGDGjqJ5n2O
ODmyOvaJLsYpc3NGJFBLI9pNehp+aXRanAqubWu2yw4DB8wpU2oUS5PU4v/SDp1hrnn7wfrf5xU6
Fg4XgjiQWgDOxbfftrJQdlftiPppKXwoqQ0GH3n+1laoz1imr8B+l3qXi283+R5262GCkRvA2H8W
ldRJ66GDWSaOgt5O4PdMPiFdjpnsfkOXWSs+XQwfiAH6oBuPGg75RjWjeVJbknw5nezSqwPktlov
uEgt6Ry6af6puebRLGJ/rXpkErIC3vxZlweoHHfGW6yMzM/MPMix91jmN7UXIVWMBbfaYtbmbBsw
hwk7khP+lqaDE2Af1jV2HZJfl01Wf72rci8Ungx+4sTH1ROWB4Va93alYAEcPQagDkG7yY9bm466
IM5PEOh7ABoMIrw58i9BqyCp3XN8szMdzowOYnlHL6MceipfdYCMbtDXOiBORlnVv/Dc/xHSNlPC
dzwY/PWc/KIBlZAebmQ2FleDgFp4CoIYh1z6oq2lKzDWiYGetTuK9HK2chVJd9bXFy+uW+jws4cg
6pgdDYZqfcV2Jep1LFryY9LvadswA5w3PtvqkUDHz8lcGDT9ux+6p46emSg8ugsDp/nRNZLDZZIO
IBq3W5Mb3Yuep8HJ5NpvEGObo/mTQWS+VMHcj2xW80FqLq3LJOy5FzkGebd/TSMTdTM0RbGUHTON
oBvDXMU5Wrk6kBVkw+jDlFfmllAj4QCR0AmVfsPkH2fM6tsFeHbiLt9iGOd01FFbvoUYII0DoKiq
K1ZLHmkGT0Ui8k5+F0wLqH2opK1QDAOoXkR9G7GnoSG90kNOXDVyaWlIFqPF4MV6hA+iOlSoF0CO
HVd9LPsNC/5PZcs/JOLXSno21lM+5lEdc+XvBFBxF/Y0jT5jUM72rIxTps7jDpXRneE+RZZ+ksRX
FP9/NllwaIFi/S88aWD4ClWHHjqkx7IjQnPCYal7t96KAGlO3p+q19y4rbPFr/CVzxpX9Zu1DQwO
6Xu+tpCBAnqc9JZxlpSJbOT+88++xrS3wNRdw10Qva/gvjG2UlmEp6e44+2TZT9wEphPbYVGkIAn
0Nugy25T+JOcJ8/N9rMUCzcnrqt1mrkM3R0p04VOngoFa29rLsp69A0M/O3eVRIdowdIxo6QkQw5
EMKUrWleLBa0V5rPZKsDPx1zzd+Kf1yMqnb+WjYPtj+pXf8yHIAAPT+ILoz9vXmd+pWA4rvh1f9K
QNQUjjiRGbI5SRZpBmlawCjH36i0nUJ0TKvkTq9ZCAdWs1WydwnxjkPB+a+C137enMi6VNMuxDzR
U9VSi3lBdKbsIMrfhMi+9zcvWlXqBS9Dqox5pzA/hEga5p03DNdlyNIGfyhX6puBYaEWPr/r+RS5
/zXkM5f06DcFu8zkwtJnrxrbFx0mp1AbpiER7IEww5jYlqGyMdWAXrclI6/lbql03wbbzHyrX10d
8Xw1UBGOKk9RbyDIMDh9yXHV5rtRNjpo8IYaHi1yn0TOxwHaykQOtB4KkRt4MbA04yHDMVYITiTU
tEHAaCRFWW9X43PseY5baNDMSEfDk4YdsHdhCCo7bQYJEhK1zZwq4iP89vs1RYPWhviAjCc6ZftC
DumOPp09ndP1pAmmINjQ4dYtQJqy8gVM1ZSSK2+7497C3wHogmDLuF3LGg9/Uc/1OaKCG6k6Inhu
u6K1vUoOlXOMxjLfqTiZwqQbU+HS6/gz0s4oQlJ2d0yW79GJHy1Z/irNPCf3NoJ54/+nYfWhs7gV
PBC+xSV9gJ9gTvN4TuPA3VqGiEisQIidTwdpW7bNTsE+4XQgBOpAGH2ja0aYdvewAM1KbZ9dIlBq
SZ+2+G9ctmmYqTrbKQfPaNcF4hnyvJh6VXUuTmmpjIr3sC9NJ4+mUytiYHHM9go5K4+oirXNiFJe
T+JnVH90lCkzxacw4+OTZbkvYGzqvc9rGWIZiwlTZrJobyGlzsSO6RpRRDSYRLT5RddkNigqdFBp
VkEntkb3oxHfoqJ7j9wePNUMzaC4CJNL0nl9ORGLNoeQgknLL6qcZRgZpRwPpqzs4KpW13oYDxOC
Do4sLMGCMxrX2WPDSsK+jv2Uz+O2ivqdJi5nY8Rjh/hsvKyKAoMDk7Z3I2P+cTbcvKNdN+KBaqjb
56YZwBMfJ6x3118Wt1CuEv6GDmqbTizn4XXWgi7w59tNEYLfB6toXZ/YlV7dWrom0f1Sg+4/TU60
3pBruhh4S7Im2KfMQ+WpIyvNpGZXUlTQJdDbLNIM/a3w3PySM14MRl0qs9A6GVq6kIG19+xBoiFB
umL65HJu2UALhfiv+A4lF/Yz7EYMx3ERVC1BvguKhxaNzZXQioh5ya5MRdGhdYmO1XF8QdVd7DB4
r6mCLLs4P3OTANvvnA7tw+23fzQi9JeldIGNWuj2mgM1X/PcU2iECEpqUAQkwVhC51AJGv44ByOR
0AiWzz0cWYCgY3HxczOUwIVJRmIlpizX7AmdQAFCoQ6UegMYlr9+ta3MIWNVjncnniaeoOKeiV9m
daEaHA6t0/PLXkBwL3MOfmjzy9zqSwu45eQTfvov4dGTM27fbP97c1kgxvfBXOchXThsZZ3ejs8j
1o9PWuOVxWmVFqaF/0g3en0YmvLYFykTvtygR7+1aa1UC+05Bv2z93pAWYAqGk4TrBEzrq3FgcGL
7kKiIcz/7LH/mzQm3Tx5mBraX74MNfIgdGclt9YjyrbfNpPYxn3FHPxPNWl/k2anLdiiSyOS9FrC
mzlLuS6LdIG51/tFzq4heVXQ/1LbkFxiREAuy7ab0nqQ8yb6WAkEfb9CYuXUgSWT+aYR7YvYlQT9
qxA6uoWlXFshkMRwbJi3HlFFhjkZlTNmXOhckeesfurq2ryKK4GAn6IP/hc7h05ZzncnDImy3nXO
SQcMvASYRYCHOnbBxqEyOkTUVG43ZQhLwyDlBpmjelnuLspVS3gx5/FgnSiYQ72pD9zLLTLU1zAY
zZSKmATRIWTV3yUMX1Q6mXGbm9gz3/aGC1CcfytVMco5DFG8rVqQEWPP9qQ9c8y1swtAXawn/o5o
CqsndCyXrzRM6whnHTi5lHBA93+JdNxdCiUAnRpNfa7tXNuGzcbSqES86lgp5lIdX16JXp5Z6fVg
hc6C/VfH6FeiuTRr2+G7m6M3dmDQVYeHchO9dDVOktXrMH4JzRKbNfyKipI295vI01Jeqadt+YMh
TEK22P1Ra7Hj9gNzeE81Cr1NAfqd0zO+5mBp80+aVzF32MS3TrDchIoRETsSb4C22MSAgDENA7TD
ObOlMYN/majwNfg8OX2WkEoxmVEYFfQDYxdydJDZQ/dckihMf1wQ+3M3TdolpeuyVZhO/wBWxrVu
rNuND7HCIFNix5lBpBO8w9vBIIJL+R3wIbgsWBOkqt2AbNTmSfpsNva1au6vIq91BxtNw7MQV8uZ
vamnos2NU+crGZ/vGhu/dZotASsx0/oPLQXO5hEASXIoFPhYCBOF60SiKH/EJrzJSjvyH8Ok9Xmj
MiEKO4WJxnqMfVMIYpBudwpqNLnnEwyX0zU8UjIA5FTsBOwlusAVooje3w7elG/qPTD4uhCuSj7s
o3PG8RZG6Oq9sVuuvn1vOhxbX5PXQNu9BBYFGpgpMoBe2SPiCPDKV0k+YMYxLB2ua7fWK0gJ1z4G
51d6ZtDde2bJVtpaJlAX03vKdAIqRnb2rZbM8rVaI/RUMd/bb7kNNlB/DaLEHyiwAmFc1Ydb3WDn
zcWrB6GFVo4EJF/8w2duxlDV8+nwRfgPDmPYEoa848gcYljs+N8EXt5e9AKTmJVXXvJaLesbheDj
0KPC698zrx4qUtlWKFNuU5x88HZFTCWfo3pt1FJ+WfKFis2f682ERSSUOHYj+r5Ln34Fv2pmNP6p
bExQdG088H1GaBh0rxD1eGf13qNFffTCmbPW8Fu+OOSBjTOBdQBQ35zOUTMpSErcvAFyRhP/PLmF
9Vlb0m5peu3SMBDySq1ZiXtST7eJGqvjDnACPajcxj0Spl6mAOMeZO5eDusW2TKSgUs6TI00PJri
M1tACKbBlsaXDwSRzN6512u0sS21zqrNJbEqRKyU37h24W7/Jk8AA1O23cEgX/a9ieIyei0xb7LY
061NomtVHCxvONstNtJXMu7R9rCiM/0RBftBW4N4dE/9E82q5fjv3C1HmyTIdcYLR7JumfB63LwP
alneZR70JAnT1eh0rvtQ5VNSoamIUqmYDNwtPA0Sqp61HQNb2gYh8NU7AwJ8F977VjIHLq6wpYd9
z0LzMNeDhQIxoGzkbNX/D1RWRZMISK7r8HsIDa1GEMOWoAgruRN7nklfRpk8wyDWKbT49V+iqRXE
PSrp8HWCUSmGT66ej9iHPMMZSXHUT05riI8551T0obruEl9Oas+sj3MTMOX0zxRCdtNlFTyAzQg0
Xh0uZ4COO+Bdm4c+ikheml2hVkGDNZqiRLaXq9T1h4wUmplhQmT7iBVLRMfr2Hc7F1/O4rHe53MV
3el0Pme4Q5fo0hQ+C3s4DeyQH4/Pgl1oZp1qpz+TqgRrIq5JZOEjbNStZU+GM41LaPFdOd6Hmknc
Gkw7WLSe3lBxEym6scP43usEie2mTDC407HpUjelMYNjRBRcKDapScSOpS7PX+ckUaaElJYkMMMV
zAXmTt+LaFj0VgctcoMv85c9jYu4CNMA3BYhq3RR7Ht3I4sLloo6brpndG7laztdkPbt4XOE6/j0
fzxosR/cO4DreiquVF0A31rpmDKwC/sKvPGfGbacyF11F1VScrOoun8TYerEoXsYWidUyblgy1w7
F+KehW+/i9HnUWpsmuQFyrLdJpL6eAklP2W/7pKI2kU/ptDBTTMk6P5bY1IZuMcIu/Z8lqWKLAYC
/KKUVl6zlMtc9JkJGYIIVT/284rH9WeAjyZdb0Jya2d3YQ8D0tE0sJfPxXqOvNZZPCQJ883ITGH/
H7RIF8/yJFgmsVj1+vbTg+s6xac+Li2QXij47HwFOTRT9mdQa6HqBHsLGpr3YFUZo0uQhLd6ivEs
P8mkiIYADw7uQm31QMpN2Bql5xtfaetZSMeumLcN9fcOMPeWalNgt5WwpWcz9+AM3aDZDy+lXTRa
nm3jMkC5wcXGlAg/UWi3LcyyLKSRuxSeNhFi72Rg5rdYGRD880mTQF26PwD7TWqm4kxu8BI1X7u5
0RV55QBY6hjfLkVFKu0rKtRrF5WtQA1MNZHRa1Rv0w+j5QBeyqOVAkWS1y8lGs5ZIkVIyoGRI3kL
pIc7ce+XDcGpFQSnpg+NfBjF+suQJrCUDAp2cf1ifs56LT8wxxf38uFk9SLVJv4s9Ay8au4eEOin
8wRt01+jk0O+RWBMjNYPOH7S3sfRUN4PxGSEKQ/FU1vtpILgnStkx7V9+SAJr4KnSdTPyROkMWJQ
V4mYVrae1IkwhpIe0GyYdgG54cCK2i5OFnXjErfz7avnm2eWe0oenjlkhZRk27aQOrIjdK7/8K01
UIBaARoRnpCTQvS5WtIsutAKm4hlpVyw5PuQgNOByd6OX6obuhwXfhbiqmlgBsWCxfPOSxz8LTxu
hVoM02GNcXLhp6LnEgDkmJgEj40RJSOjBui89kJgPSBqaF5hg9E3CoP4Fp5TZjIaEQw2GAbuGGkl
zYFjlGa+XZX7X9CQSuHUgsZ4enBt4T2AO4h/3dp1S0mYktW77VBvyrnuTTBBVp7lOUCuNTFmftNP
zlQxHjeFc55LgIzDhUJN/WPjrlr2xSTQAItI8mSmx8ANd7GP7jdPWHNE67H4CGgE5MoNc7vh/zmy
6rl/b86WDqBYoIEmXA6IhdsSxA7laOiNF3cpRDAcT8f5qDeuQef0YtJmK0AGsjxBCSkqZtx9ILsW
+weZQDvArefRnNkyi9bJi8QC5e5aeOB1hq59tAezrNdELMeOXYNQoKDtvrqtUZPz4jQoDL1v9ndi
1qYIdBLHDF0/zOKbRhi+2LA4Id3HSZcp4X39rotTO9vqX/3L7wl2IHDZPWRQRSZ1fSr+nudcGrkV
UsopGOYUJC2Ih5YNndta8y2dAlu++XEa/lzxU3x+dad4mQOXcIAzCpvDJFgd1/i4dx5ZtmEW/jnf
tXnGv3RYNd8lv0hskKK44J1P2LjP5NqntFYB+sNC+HG4rfZuBPavFwm0AM6dTDGZ4lXScjrR1i4D
QubRzqyhdlXDDus5MtE9Go15ig4WyzQq2PBAalnyO7TFzfFHZd7ITd5j6VQV3sAAfzHCLywZfdbH
GSmkTwvSnwaEC9gG8FHuLxHOMGHI11A1nXeYvQE1DtGq2p9N7inViFoQOV7lMQm2l6vlWoE8jNyM
G0uwVCTof82BbDCRPYK3D0lRAx2TjaqWMsQvCFH1ZhpILsDu2j7Xlsw/m/AoLM3w6ob1mGylLIL9
vRZIUdvH3e6FFeSZYE3lOK58hy/ZmFp7ZlDSPmuM6Eier8MeFobRUSruyRfQAOgK1D356k64abs4
h5/TlChADkTPV3V9Zv9aCW1xn7vRQIfbvXaJVFNBLJN5sMouF9G0N31t05ynO0j0L9z4XEbM6KGD
LKXkT/hh25aa8jqT+9gINFWUsTfarcB+vB75697pzGjbadacE6a2e8UT7/Do/x+MG8ssFx1sCg57
xeY2+E3om+xLcjJmWQAVzqxTq4mpX8vf4KKvlfP9IPFlYOMsL0y3soY34hIqmU7a3UJTDtwiHVCS
V5BbFBZz4QxILwwaTNPFuR1WY8hE6U0vDcoh5UMyP7HD2tZ1MElX7Xm5MpJEqe8PKRVnDXNGaAVW
8M6Lww9u+KLSaNXJmKrgr6UgfBSpS7EO46s6NyNeV6qLWH1qLq4HQ1qSw/HZEurUzPb2JUg2S3mp
IddOu1LoSqtcpONu4HxhDxY15JCfSPYoHlZSFhacUDPMhhWuRYfaLxU2xEceaCrjT46AmjPFCHiN
ToQdYzy9kwgRzf0dFkIiKGg98dbP7AtZwFeAalmF+Vzqkikz69dkLymNIvW1PO4p0+J5hcs7ci2P
CM6o1bxglkCPqknyOypFwJsrGV1r+pB0oYfVTXO/SwxZXCMFZBwOd9AuM6Y1WQo5IU1DcqR2wHnE
q/AvTpCRa//UErBpMUtSah4IwVfo8eMlJ81lTD6dZYMLkoHjq3yBGtQwLjqRLD3buU6CNqC8UnQk
X2H3r5ZlQ+xjp6x2OqT3w5NUNC1Zi77DEWPluIenE10bZDOkr7iULUTjDynHLxy174fIXuODFRK+
0US/uaR1sJNP6dT7oxnIcXlxyn8f3UthzKAxX7MEqU12nU8qzmFQAo7Kit04/EeT/tyiUxlzQul4
IXyZy+HuPaVMphB0SxMBy2W9ue+elTOSX37veu86NgrRxZrsdZ1/tiLB3uW/p91Z3R9s1yLbet4y
fiVUi2Yf7U2OiVnKf+IV2tbzYZn8genT+wGhVgRZUk4ipiPEsTvnS4ReG87hHIc4cm9u+xIAbdFL
VesEp2Rld/nHdWHtDxndauCJXj8K7abP0/eRrh4EwF5h9ge7Y3Pq3AVMHctnmPnhoTfOCjeuG/n7
KrBlgF9JA2n8N53idMLSU5zB+SwdSU9m+9zFD7iYqVcYKLO+WuqVr5W3OEi6wQmij+Vrtxt1Tmqy
36mMJVwP9ghQnwNyxFVF60d5rou2K4WgJwq/N2DCzyoB3WLfH5ZpXSt3TBTtyOpOjvWysYI0atrM
vWw6bijqhnPG4rEO24tDVKVTOese5zhH3duCkBDcCRhojG3/BVzpJoMy3uTudlDK9mkRxQxDfYPN
fUIbl+XpzoeyniX0yFleOS4UW4e8ViquHs/+u4WP9fRW847TzBzoepohoNFp9xrEz8eZOzAOOmAd
Z2zBKEyA8vqetAgSkYiarz6nHLNZXj97n8lt9YdDjXoiA/AyJRVyCky+aK0+mfOfRg4CYcgXxuj2
xRdicxAPqHfvSzr3D94T7Nz1OJtqsDfAD+JFeLKkzusY7tuOS7umS3w01QHti34zW40bIEmPPk2n
QI9RQRKHXNOQCKgiJ7lFvJfhTmOD9fSHscP+Ty3gvxUL9TONmXYNKtrhh8MG1X3qG2YB9SCis6Om
lNZnfBHt1bry41IpUEJfTd0JbdY5NouCR2mZmKHqvBvsH8waTi44iD14o4TNyoINQ9YfJZUlv55D
aEW8Io3uobbbJlx8HneDe4ZfPl/uPPO1gPhlaNIZdmqixD8mKj7jZbeHBLpIASXtdvieFwQ+28p9
VZORy1oIzS+wLkfYe+mB78RtQT5GvgQ3cTzZ7hOx6vc/dqQZkRW/zxVd9sfw50+20j+gyuQSVtXg
PVZuy8HZ7xjNcv+3tM9ViSyuCckT9/s0JAz4t/v6J3zd8w58zr3n2p6BafC/XltqSs6HLuhl38Z7
um8DPQuHqjBsr/MNl0TeQoHh/4+4d0Vh3kYriFWPJ75+aSF1ayEbvz9dI+C+G747IyHkgz92PQK3
SKxPldSAhK++HIXPXBW4gAlOleTRbhPHO6Jb9Daasy3+QtD15x+D1g5h8JFRTKvGYXJXZgF7aGah
3hG/wEbHH0FOb1xbwA1XQPoPU37jwYlrpB77a1WaegtZEeNrEsNzUiMZvMi4G2XWkXGa+LLk0lPz
xmsMQlE5qFgCXrAkoZ4P3MCC/3SMhTRFwxJrA6Me+seRUd7EKlqS+GrZ69ozfWQAtUaHaKlc18A3
phlnYno7KCBotFw/n1JauRAHCWEYRR6poJG61796hNEMZMFc6wg4YlUmyITb2QY7+36kIAEs2RSx
E7bgjAhMyAW6LGOIq8uOTPG4c7q/BBWYMWji8/qS5WsyQ91/xJAYrq441xsmTdrrwVbBOGxDUayy
tvRyqWz+X65SDH211Qj3PWy2Dkdnu0rTZaGDpdYNhMxZXa8jj+Rwuf92LP+wI+XnasoySC7A8DwC
zyIoOAvKVyfrJWqg0YgWXGtjhFTDAdLsJox+TdouHEcNYh0rTbUqDTqWyFuBgU5a+43tZrKx2LrF
8g5uaDP17af6+Ivj7z6BU2VwF9Z9p2ZN/Tbj0wksAHNhaP1x6Cer3tBgn1Er0XbytTKb9EVxQ4wG
2PQloKUAIAceunXfw6hE1h/SQvZirjqEkKIqfMZjdZON1nTzaKMRA0BkR2rw0nrkFXJYIH594+AO
vZJTkTzzBR6thVIzLW1/hcipRXLYkTbmEGKRoYr9oTg6bU0z/Qm52Zcd+QhhnwlHEw8z+Oc3xelj
m7Lo/KYNjtWmxywLrxf27XQwwmdwteLmbDuQWviPxGdOEaIFSezLooINQ3fNELHCqK8NwLkiVM2/
I82+5LHepWeKsrR2zOYjlHx5Phfp5uE97HL56gfZ0yEFAKEc5NgF4khGOpH7Hs0WTAnQbn2Rmr1i
HP2PZhRC0qd7Q+yNBcdygOifTn2OdZbFFFtfCUeY01QU/++pi5fsnAQFZ1k9Yc28gQQ2F7nndVMg
bqQZOLFmnNg1BJYtERbCORqtAl5t5r9yok5YS4k33O8lrpwJhIktiBYnomCWUdkcJhEdWYl2Hv4l
cb7yVuNWum1lkit6HdCSuRibf4Pqw2TxGz9hHYZZcjBCgAVEFi6vwBFDyDb2yR7rAqFQOvqqMe2d
wkw9jSruJj4RTMBfWVTcOXRHfMryT3dmYcqiEiu6tGy/X+s441Y2XFDbiao309BSp4mlsZTTFcy2
OUDIowyB4CVzUqMCC2NAyA98mx63Bbvtmi8UUFF/2sniYKEBRxsGeC7raodVZCjm6orfuP1x7hE/
Je+6fcJ6qjB3RwsqllrLrTfwYoT1UWNKCGu6nDljBKlhEjG7CTng4XlONAxmfLn1DckLW8nM1GxP
9HAro9U6lzPgrt+Lmppc2P95Y0KfPapj2Sda9JDvHRVGzDBxFR89BbNq5Ex2ZPY4nzYcEPFGDf94
x1D7bbXczQlOL8I7NVoZ7kYylgRR8R+Q3B/MKwFL+HljZbtkC0qB+NjJQ6EUNtcJFZQTGqXESIop
WQz6Bczj52qlrxn/R6ajnlMd3mXkfgbcHnkqa86pKDplEbBEJ140yqB4F3/p4MMkEJ+rvydmPm++
hVvHyZRHS85ZpSiisDStWlme4MWNuA1MW7nh9EgSO5EruaxYATqoIiHmS0XV7ZeF0ZzLAkMuc5RC
uveVPzqej7JSZZGM8wUZb8YVhu5O784u4Ks3fjQrwwKXlmgNNHbCUo3L3M0W/JqQaUcc5cEAU61c
H079UdeEB8HfhAd8+qnPGi9oeKAw/TBc62ZT2J749LT3jo+sgDT9LN2cBci85X5uZV8/5vvvxfdj
1GRV1SIHuoLsGODncohExHKmPCCxOdW/L2Bi9HlUKAeD4YdTFvnhKdvJbmYLxHWaJh/iL4nukvu0
8sG8ajVxzq/pQgJvgXfg7/n1EIU2qMl5ubio0vj8bQeC6wULqzdalm/c1CQWI+U09zfPLrzjyqKj
2cMWFQcmI6sqJCanQtbz0nr83O8iEiXsKSku6SZ2Ll4G3BGuT8WYB3wehGCOZjfqf79lYVqe/Ho/
sDzhJjR3idxZAApDwiXgyfkawQCo4ynHN3paB6NSUk/LOpPPEbdacDaux+IzYCNWMdKJIf6U+Vun
NhoHNhIC2lPskjVhkKS4d+qOhk9zbSqRC4grxYhQwgtH8rCWB8oyPOx6oTDtrTT33jtBo95F2UgG
5ZVK1mLoAu16m5JUpwd0QajaEAW54aL4uE2gqntPeZsuFEesMmv7LvNloudNQATsJiHUI+aocHlH
E/jAjHVlsbOUSNTsYhvOeBxffWcgFsBqyuP/2zckDa0E86/tLnebxDi2enNxniGLqRehpIlCFKDH
Tk82YNH8heZD5Rc7eX5sqSmulf83Eqw5ZA2qrst/iPtKEFXDPM5psfij91l17tqTiwcOGGKq/Mw1
12AMwiM9lkvqzviPZMt6/NQrBmI66Oxi50JBUuwgnUcExUsJmxcJ15Hw9hJR7dryHJY70pN7kcUI
JWS+91ZXzVqd0v2kYArJoM6K8PmpkD+vm7Hv97tW7Bv9VqIjWRKALOGzxlJ3qkYdHRtZ8ho8PGGr
Z/iaMniDOpr7+FpQUgFjnBwPMmAvEbG7rmFH8n2m0ZKrvUNsaijT9jgBdKGY4/DEcOwQfcPelOSo
wI6u3q7BfB/bVGSRgO3OK9PvL0IJKN4nJopRzfTBJxU0nNZL0ihGDyKxAnQl/6ZDIZCv+q3XnUvB
GIan/yEHAv9j/gA6r0GKp6fX1WK4JzYE8pENCQnrO5Nfwg1p5fTF6vOy3SaSp2TTBT3/jVMo9AlL
L39+pDi3ZnzdFwFM32DDSNIBNjsOV4emJs5kdUij3sN0HQKwNRXfV1ne8WwLjotIR9BUNvdv9tCb
qimOvn0Td4juOG4PxIeCILjAgAIwu6Kwif0meH3Q6NAGaeA9DA2Zbm0trymTU6N7kk22NAKUnPRJ
CBPsqXqsi5p7YT3rxOIEXP/p1J3kQfxm91o+MrtAQ212LlsGhT30HT4yIgo4Br2pzPcC1ZGNdL1B
wECxXHRTmFzBfl/tuHq6deAbR25VE4QFizU67U4mZD0lj8mgwbKBr8lKx521Bl3vbtsgL8gMp4Z6
jbr0FGukBhm5/27Xeq2nrRlG4pFgnBXa5qRf9/wYUHLGTyffU/XSnlj1KV+5Qd/0E/xjAV1Q3Csc
/ut/4oxWByGTbFPmWuPLNLr35KSn+1SMo6ADft0usxPAeU3WCXuIL+jFDP5zoWpkV17qn1x14PJZ
h+Oz8xGoZiBhGJ266j4MfP0+l0XZr105J7fHuH57QZyfgA9ENk+WNAc54dX9oHjYQbX6mObGEInt
tKPXOFiYpnFJPNXviDulXZ+iVtDyWwk0GnwURhheLyeM9/bWxGrfnFqETHx13SILM7Be5u+OVYB6
3KP2kyPZCgANTiJ84GbI29AKGzyDycPuwtjWH7EjgbupfY6tfeEL6U9n86LGjqjgN235OFatK28z
d6wEx2APeCqihO+che62XVk1ZdRXntKa3G3eb9fx6R4QuJakdgnVDsaFQfj4h976tXn6NK8Tb6BE
e7ZzcLxpvj82xU54PYzH6bK96nyxryiLAsT/QSpNLXugonuy3asFsG/JwQI+xiNTGCVBGVdEoDyM
ICQc5PiE7i0eA1RAGBoCjcQjfKPHuw/qXMID+ZZyKBrfet/gp9Af03EqGG7cqoo3ff8pqVKjig1t
ghTPLtCmSz0I+Og265/axwQWc96PANrxDeWZ304UNCTbWiKELGOasFb/65Z7cDW0D4SkhJms1BK6
9d2QbUpBF5GumBFcYf/7aB+3ZU1t4G7YBFV+Z771K7beTyeW7rFmekNCvAfGuHRrOnd+jUQNBRNj
5BxLXzDUGqUJKBFHU5bHN3t4Kg8WkhG6ZzCSTyo1KfXUY2lnZmJXzJIOZcj2AZUkTUNZ4EyjOAWZ
XMWh1dwNSthE6EPAeorNTY8HptZbVFqsac0ol+IAT/bRKapKREwk8A7ftewuqtrlFwT8xJYM7Eyt
T2IogiJm6u9x3iLdGYs32TM4g72mPX1wWhJCo5sWiCeXaw0Jkjo/XC66kYvAPJDhfrI0TlfxjRgz
1rNXOAsSDrbYv227vJxOfuF/Dd+cLJFHZ2TdQ2vMpTTzIHOGTQr7ZUpd2FCUqm2CiaoPYF1b/DEQ
2e3Vm8Durb/DDVTTRw5vCAIjRheAf2zqHYV58jJP2FjnaT0/1o84diMPky4ArOVXO59h2+3Jgsp1
dKRucfjxkyUi9u3Tc4cSQK0uVF7V6jRopaPe/u25sTE/O30D/n86Aw0WOwiMSgy+LIxxN9OtmUty
SPbDYq+wI2ENv+TKlxklyesrBoJvJgHIKOnqEy6n75uyK0fUy3XY2RiWkMVMrfcc7j4sO54JrZMV
4MJpFA5XTeqeYSoV+BqX78EXHGv5H0urJMW04otq8c1K0cWTt0/CSgyimKRuMgcuPTnNwJeft6Li
ghWkScqYcSVWoT55RedjvBs0ucEqNa8c3lzDtotRLP0r3DNhzNJ2bpx3AOxKE3wfjALoF6ZW/HCH
I4E9oVldxuf9k4RkE5GlGVSixJX9LEOM8o9OMls8wfRC/rOkMb9mlztJ5HgOH+W1bvAp8bIHQ0z7
4zj06/vUQni3V6zDVarm4sHvDUEnL0TKZB1Dy627MFAVsxdum1GmkfOrSbZWQ+UJReM93URLPCxd
K1t7iretfPMdAfqR3M42SVR8KBpg2zsGFn0OctNY7RvWqfVG38yo6CLdCGig/cF1ONSaMeI6JE/t
fDBkTX2DHtXHtEG3lmeQ+vYyiGmpnufZt6PLVppYoihjli/laaQDZWZMtDlE5uBWSlDeDb46nbLg
Ndg2ZSSrjrJJLvCYKqrYH0W2cVDjGINNghlt8s0gJjA1bb94cTrCJFv8K7oeJoxjoBlVS+yZs17p
T29YBv9ymq/yF1y55kaf+SfX16/yWmA20OZujnBMIZ/uVbsTRsASmuoyldjxnxQ/8orySqirskC7
61Q3vSOfTgeyTXX5OoQ6JMIsW4m9X/LROjVdbZdkZc1Ko9Ls2EdoUA56PHePuQQ/pu3aAVMsbkqV
Jyv0hzfRCxv14I56dsQvs5O5u6XdSz9+p4SGB0f/WPSINHkAtSPr/N4M2vNnAVVdJV10ql2U30Wh
TTyqSUtCFnqz6+HPyQed6ES3omygQzYgttC8Kvh0OqN47Gz8YP7OCyW/eRjuH0RhAl3RWJ6DQKcp
gfJA4xwH4DQKW/v8sVFUHe9vp9TvJ3I4NaJKl6zK4mzIG/6VVug38IKlnN2vQIN29YF77+/NiRoj
biUBeU4JncVuSx5MT5cstFQ18pgKyd7wfy7OExAsPZvwWwuQEtFK3W1FuiSKRubJMiWwzJoYkR7Q
uIaLkVWgDVNfENHIuuKRLw6eQcIWT9QB5xHiEN/Ig/QUMwcPSRXteTiblv6J5syfLXHTNTnyxDBa
FZ4EAOgXmAZg0f745SOTq6siszv7c4mdzMfzenmztuqTWzZ7l+FDnibhMf3xBQe2GJUK2HqRwAJM
K7MCgeLBgVUHW0VavZQSOWiMdLg7dDHcyitg7QKCEyhCRDg/b29S+9kfZrvaBLyGiXoF+WvflDMG
87bwNTOyorLB81JptslB7D8U2FNthOOhgrAPfhKDDKwv5ahy17akFdKJCI5aOQUzrnng/3valpsJ
2pzhwvVTtjbJ6d/iRkuG8LHQHQOZBZ9O/MzvM5ZVHrRtO1kseKjRdBow/SXoCCbkclyesp10ss5i
EDrDd7zYAKoI7AQr/mfCGbqtyHTmJ7/zEmFQj5sQXkMZjsDgv/T4CKFU65jUyuhn2p6/npJ8dKjI
hOvORti5Iy6DgnI99HPeY09NiCykHfe2MCMiKQ105KsACQ+1d5JoZIY1ruuuO/5D4WrHAIda8PaH
O1qPZWZ+GU99ZCOsAAbpWC7YmxDH8VqFWz5H8TwyGxdjXMtJDjw/E3H6y4m9I65DwxA7DgnA3ZjV
ko8uAF7fOBAj5ty9s0ijGxbhcSDpVk1YHYYLj98oGvjk/rfQIEGu4+LHcrL8Ac6Abphj9isUok3X
z4Gh9quvbN8ikc6vLRY5Tybe64Zs6IxnjchBQ6DD0oU640v/9Ad7mufnJxz9f6y2ny2tx8u35DcK
QDotkw7XyJy+lF7S6w1Vn4DuNX9vrjldJ9O9HiTCv9ttFzN+hsDue87n3rMp4ueGdZfFPTjKId/1
G80x71vll3bYCSXjl9QLFzJ0jF1mxNTHyWrKoyBPltlkjppseFbh8H/lqlqB6RFj7H6OqmaqJXX7
TQgP6Q67V1aGKfcm3y+lIaxaSObaGpngKMPX2JbJ6EhkfeauP4C+cNj6f2/J06pazOBPWMavzGPC
BkhpJcIRZtmGNxyzJ6scF5L1F0+zn43okJQm0N3P4nUAgYnxXrepXhMWBUugGNRGzN1sLnpEfSzE
tSUDqIWFgqVfNxfiEp3kfpmS5LwXO+lfai/wGsYEFkm++BJTjkSUVxDV0h24itIDN68yARnRVfsY
6/KaoIW7+IqQGbAH5tw5IcGk+zfos0uzFYFpE0f6gAutw8zKP0KixyI5uI33PAkZZQulBNl7K3j/
tNtFtam6L3GSo8Y0L+X2NubJHIdQb8CDwLigt1Fz/PIBMKRguZes9yZBpxtfCs03XNA+00vTUTzs
AYcNQVevNJuQ4AaEwojKjSde0CgMP/yiy3UQ3TOSYsBeodMAVjck22u5LWC2JcWGxRfDdlOE5WYa
Urz8ybpuRGFuqZ2sTlhtOGOM+7yH4fU8iMjdC33U9erdbo8h2r8LnO+JdzgAeo1TcddZ8+bV7lgH
M7O6ptx/uJi6V5n+i4MXE44aJ0ME3LsmKKY3ttxiLU0AETIoYarx7oBKKmMWsNL/NSqvUX2xB259
pqNb5mdCjqZVQPJ4IIiyPTescEgqll6xtlXWXd42av6m01eWNqqZRV72SSdMynN5HzujkdAmErsM
WkYqh2qvq9kjLT0t6HE1ls7q7aU3Hwmrkfdnp3YNh3HJxXK2TdetibrJHn6ww9s/xjRN1H8BRwgH
0uQhEtMoJfNAJRIRPpjvFAukOEppuC3mkG6SJlGDuYBOM1DhdXcwt8fcZCSPVN6mOCA6Gp5ZhM9/
NB46CBXNm5c/wUcYM8kAk0udnvsxc9fv/1VUL4ezNOZPcTGIV6MVmvSXbR5CUdQrWm5V5T1t6f7p
sO7oaq0wMXpQO/AMstGF/3Dir5amatwZ0NgcywhAUEAu5x0HUJ9zBMr5/xoAF9SnvYHbXm/uJprt
xLs1YmI11y4sSNej40KusN6GuavLwcNhAUrRTn8ACIxQ1+iwnWxUjOx3bEQCwcEFE3eInQDw6te9
UAfUnirxij64N3QHy08uvbv0HctaRbBFCugcDnP0l7M59uddbSPeTjrhgZAAPW9ZXEqZ5omSf7ue
qZYKjOumjVOXtSjWsuppP/R6ZGUZhMysY/+5XLywFcW0r89jW+nU0shqRGALujyZ4yWY0HDG3vUg
zQJw3Yq734MEhBqwhtqnFCM+IspHFQN/pE08L3eTf8zwq+QVlHDqnQPcrdOlK8vMyUf576KkaBZd
NbkYRpYFTIVogMt8SGBa3Blw+HXfxtZuOeQaZCEqLqjLAM/T7kB96k0O/o7OAhcdXVngFqHU50p0
uXeN+++IcuZkVFDVLgRXbntF9LgAp1IiVuEf4Xpbx0q+s6oPnZzeq1ojuYyRqg+wt8y82bArdWh3
7fWfhDHMqvXtCkD4J1WDyzsX0dhCL3opK1Crji7Q0ITTQPW7+6FK03aJSEaRuB36sTTsaNYiNBcP
R8vGie7YcSzEIbnJ+zdyycF7CpseK7r+HK6euhy+9lk1zuarjnKqaKQkoG3A4397gYqfwl3c+AiE
j5DMWXq1zaKilqTo3Xd+oF6DBS57B0H/6sHAPSBzb3z+aK+35bONiiCkvU01XWpftL17mcCb3KA9
mkvZS+Yoy5EpfL+b4OmhMQFU/iIXfh62dfIuv8n/W9Jkt9mVT1twkKIept699FBnNWb8ZDmR1MeN
wWeY1iXQgUdC/L0t8Kt9bdscJTH9UY8/HXZXthUS5e/bP4s5VT7/hojEY5XxJJ6kr4lkpurpPwrM
sd2YtOVX9/wbNDUdjeHM7/WQ0spA6YiReiPXA7geqOg6uQAh1vwiImqM/IFun7vVYRYOyxTWsNNo
dhnm0b9D+TaYU/2CIK5WQKUaEO9VMm7ZMjlw5YhD3UQVw225jSCyhcKnRluclaZsCF2UBdnruPk0
v1js907Zv65Ni9C2t6wqvti4Zcy/Sr/f9SpZsSxw0j3SXOyhfz9k9/Hwyfw7eBvetZenXyVaKmqX
XZNTCLml83Ii9sVYPJZGsHu69XAo0rKOywnmVD2ZS2IhXjePWwB/bQzMD+sDqfMZgD8t4sId7ykC
yNvRGj2/eapMBYhvYKdK+SYY0iadjGhqdIKpVLg/kc7occxn7Yc+BweY+HgYzRRUWMb8z9tcB0NP
rXHwyqYy+oewW/M0BBdbj8Ta87wdxf+u6Ar8wsQiJ36xUK3Ri0MFZxJMbruOZlMpvpow32yX7a3V
m2U1zO9sehFpZVF+siBRXBn7UBy9KVkidsy0jglDJM2yZYmEAB35YLdI88OQ785XQ40Qs1Dqm7hj
+LDJH4QrHRCiYmU8eAQ8lhj84V6tYnQf91rV4TX7WZnNZTgs+UyDUIey5MF4uj9A+SimlJgJdE1i
nViAAf9jfDq0Uv9OhfgNMCu5s8jAYlUGrW8XAQpOZm5fU2019SqcIGBM5crN4v8b+20iME2J70Hj
0+BbDtf9g1FVs/nQbzecAb4MykW7Eyggl4oFCnQS393S/CZBY7v7YEgjCrDa/X+3Ky+dq41sjeXz
q9gjryaXy5QlxN9nQew1Ipgzf67yPfyFFvX3twx3jM4rJyLFVw0g4QcjbXjL2NiuH4l0GISWO5wF
feBthELh3DEzpwnbHEzXzfSjRtZ97QzuGTezEO/QORlEA+y+I+jbpTELntQ+ndFYil/qkIgb/67E
IXJO6hOHjDOmKqolWTFCcbBv7XHW+vwk3EC95QxCkG1eL3+HYXuKAMmAnnrW3rjFOjvMYSIQdfSS
jJJqBVvXeKCu1RB9NaDdIs2sfdaJBz2j+G/VAh5jz7W39kDATsB3VzvRL1Vqi5U7Abrr4nfyVRiG
uf+B4zlv3zsm5JRZMZNyQhEYFpDtfXTIGNXns19S9qPrJlHOqxkIYdrwwtqMVuZSBMVBhcg7zxCN
t+gLZR+yIP7NmZojJJvlm8kJWbGV2zOgSJzwSJ098yCSfLceQgiqKgu9qjhufUV9uYhwYWUn2QWr
zBMRt2xM0TTqrYcHKFi8NTNUZziYNew1WzKzJILeTPoZ/vfC3hKdmWhDP5um9UxxO1Xmt1cX0zpS
GCnJA0tBBg0hawOxFvKP052/2cLwqnxgzQKJZ51ZoQRFojMYyVpnfbpsfJllcyBdvH/nFlquHLLy
RssZrUZXPpfAe8dOreJjwRUhcRe2J2O1X1r0Sopymp1VonCVXLw1nDW1Lxk169SYVRYXaymzvKYZ
0LRYkVKDt/UFPZcOzhWcasUZQ2BLiX/snfIQ2IXRAL7esEt/za6WaRBfTajhPk5RGWw/If3oowWX
ivndf9J+AaAaPfIJkZ8hDe/XemAY6gJYchM+ArBACfgtlS1UUR9g/0AuBkvy7I8vRXxnGckqfyYT
/JBbCNt9GvvQPie7763Iwep5BZFeI6/vRoBcuLOdJAzWB6Ew4IyguT6U5lKCr9TfobrvLk9a2bTk
dOWHQHbIv0Tc1gU5hpclNDEuIv++y0x2qsG4dvMoCooRZGDG3TTCzioxtF6S/6qznkfKp6QeL6aW
jqZA/NWOZx+M1Xh76U4a66x9ovcsFwQPySLrM2cXge2YCYr8r3wS8ZdyNMWML5KhFVf8WppYVUTQ
fBb1/e3/UJ2k5eiY5KQm9hmM/TeZ23KWILfywWn7kiJNLkSHp7jPWMWdDHy6TI56qdJkNnnffYg+
38m7RlCtL1yVlS/7XXzN9nFV3o5sJentQXYXdOZLKiItNY8t0b5z2jZTZb5LN+gMXxjKbooJHoic
gHONXDdhVIh3B+PwSLy98jp2dhsMxRf4Zl+MMDZK6ZFC7G25tLR69q7OXTfq9JNBeZK3CkwgTtvi
JUp3FsUXpQ/WSNmxVguY1zXD13QJTYuHapkIjOkPItHdLS+Oh61p79vsaSo3Plv2pKDtn9DnPcZ8
lPxlZHCiOsJRyaT4mo3WxsNqlLQvkxbXuScNUKtZAn+Ln/iODsdMiXUfUiPfrIpUq74x1Q58fq57
mrq09Z6or6SfalR12mIYRPv/ttn+jxANfZwbxnlJbFtqF0CmWmWIZ6dBMsSIWrpurVZCWDv+C8gL
1ggAb+Tw/KxUtAhGaBmFGQR8NGqh0j/vN/LpynttG0gmLJtE2f66rEhRfSELbgENB7W611dKwepo
uzyo4sZKD6cbjq/7zIRS0GswmJtOSCRJ5pZW7AFt/4/G8dVf9zx0VKU0C+AtsC3Lf8n9FOxOwdcI
gbM/m30IcZxLqezTiEqqSAgM0x5n5Ym1oyhRLhDs4uGhA3bXEJbbhlUNTrepJGCP7oPAW6kKXPt5
llE+qQOCxqlA+DDUVRTL7rWsNwJgWRhT7T14tOD0LbNhKfZmfq9fr7F/ESwO2zDOKKy+b1m/xLfS
Xq96lTK93zMNTkmBc2WMT+BokYy6Ri1mcx/6CT/9ujB5TPX71tU9mfKuwouJuXMRjs9QdE2vjh4V
gfFRyN1xYxsPLB9l3aDVFKVm7mRQE7gLcPq8l4C97u+uGVt8zQJrpdbPxkmTBR2s3urbB1X2lsjR
RxQcug6eHtHe3wJFVbtI3NMus04xTGB8GU4pYSHtERr8KsMlu7Q8yMst3IFFqEG7379xSxGtta4o
mCMYnvFapR9cqLI+uqIXyZ7mIqT6C1IFZ8pjVHMYZ8UI+0pkh+mIaPiizLfFy71RhzWdIzzAhgz8
zogLVGLUV4OLznVecptJJS6BiCQz9KouE309XnvB3x/3cIxaPzRR7MdjEp/d+UvhOo99da8mS6MV
acMsiNqdqmqJnuxltUcvT1BiXLWalccQkRgs38xa0P124DlpNOyjDu/Se1j+R6TBpRKPdpc3dQAJ
UO/vKIyYTNv3e/HaC0cAiMH2dfDXs1UJ1VvdXTrPU0WQYeAVYmWfyLysRqDLUFloj8QRajHxDhCs
hARqkKIO37U5hJnVQ0r3HN615KP7+RfBbnGajza9ttPR474bAZUtxLwUOFc0RCj1KS9v4VeTfOLb
5o2/GQRdJolmhHjqoCKnlInBuUs66tUFxOFjzHgZZHsc+g45AbG5pSdqJU9LxcerzfjLvJn8td8a
+JsQ2zfvG8Kgi++Sw4Xhqw9xZ9UAC637ofjXdYAbSFMuZds+7JL9TsZ/FDhtbH/xRTL9hyC+tbGb
UacIrkzlsiHH9CBjk0xZcS265H04GD62opF4TUfMsohD+QKZu7BnS7r5RaBdwlbVDg0r0RaM58Gj
hQLac7ul90TdRSSWOGdTOtJEs55mJTgphdDp3q5EPT16cq01YoNJ2eDyX/WvdYkFPrI2uxcUYSXO
LUyM0XC25UOxaYbA8XcTaWhNUS6J8Ao4GY4+8A3hGxz5jBgAQn330zdmiYsN9HaPRoTaziODAEeN
uAJrlX4kF4UkWudOBtuSegg+dCot+vlIm6e507OjCE7aphVosCpnqaUgfayU32/btUSrMcBMl+NE
Rkj4anG5Akb9dwScGDJr6KjluPuJHYjZj6mcS+HDShp0ddKdpQxVcmUq92iSNItYCaBmyvDctD8t
5/EvD1hMZsjlHUqDqfWMl2HyZLujqY6yj9TkoMW/DFZEjUEoDaZLlLIHYEgR6VGG/BuvTwsu4ID3
yP6DwI+nM/7svX6Lvm+4EW6GhLTaABhKuZknfaKxxk0QN0EgB2OhgND+snzQeJPrraps540sAcAs
SK7cd4BNWEdgxWpCzsWJ/MBQy9juWFiJ2XceCVRBFk5hvB9EfEQVSCYcbF88yKzcQ6xuNhewS01x
n7Iub42sRgJ7/VgHwKBybD5geXfalCGrjY2YEL5p25xYVBomzKBzgDkzp8MntY8dv83B3Y3QOeSL
soPTxFFfHJlVv7/JO7R6P4K4f/1dNRRiKFhfGpmkXF/xy95rfKj01AHpj3i4NXx9Rlvv3YVabv58
3KO8oIXjeMDtRgMbFPg83UDTv3fu5T/MoDTfjWw7KquOr7r4mDL1TpUxW/ORR6ZZ+oOPN2BQPIJJ
n4gHieEA50xMp+TkDxBpCQGYSU824hNd6mIzU70R0zd7Lc0yZJ/Xo/Q1hLXmnmRZ/3fFadVhHLuq
NEaFHlOEm2YrSly0zfvQxfh1m221JyGlknYkPjtK2L/a7Zj40XXrjq7/7oC1o0CCSj8Fe4zxAIEZ
394/B6KmSQjOOVuUPbd1caSoNEc0cq7JlgqC8lC3FqmkQKYo+yqcyIyCCyQI750WSs3WxS36YHWk
N3tzKJnK7ONhhI4PrLMrrPUF+kL0iYZjpMBYo8zjF5fY712/3HP8njLzLepPn1U7TC3G2uSi/oia
gl6X/Kv7Ft/oWkDXHfBrD+wvErntSjm40L54FHiRIpGY2YtlAKy7CDD3zFe1YgubzxfGjxSJeIBE
R0yGAhMQ2fcO956HKHvwZ9gwh1Pj+17E9G+HnpgSjQCKZtXcu+oAeCSOJQZb5q2Tu74Q7dsm934Z
HWdNdP1YTUnresul6wImTIAq2RnHTP55efPP7GBwxgfe5lORRs0MD33tp1dUX6OfOX+s6Ga6Ocy0
BL9fjBt4wDxaPEuA1kTfqgVtAe2AfARwCU9XvrzOFtE7SbCXVF1zlF9IKImbkQ738kee7Ybnjoqx
nh1VYN4h1BR30ejzt4P9Uz+WDp3QX9Xt41v4g4eQDzHG07HnNHwfqEb6yz3EqOX1ITJlI2x5qzGC
a29yWkKLGKpVkm5HiGdoTXfqQziRUhCnxtkYpVhN/BWQNEogKs6uvyc04TCHOElPuLe8e3FZNHVo
LiDjjVzikSkBXNIhyLvyQ3EVMl/BjL5nJvw6e+QeQaRETi31kLLiXTZKDlfAG3fdJvS5l7rYH0v4
7J+3aB+c9NGVnRhL/hKjw7hyDMMxtvE2am909H/H9GgLvQ0YF7apVOe/dSX7idduklJ3gx/+R6xB
Fa/FqV8Lo+JBzztwJanfoH8vfZoYAveGO/s6JVEbSufVUNbeG4QMtnDAfnVtZT3ZWzWmuBXg8qIl
sCLiU/4m+Khq1D7XpRJmBaK4brw6DLT6besnsShUGEwpxdFvuMwzYzqxgP2OQ1QtGdFAKkMer9ox
0SE80wvvxUobnmjTAUnJJuNvfgyCVWT6iFfqdM35otA1b+m6Qa0kaHeauAhu8MaGXYNi7CZaTW5a
0iK88YGZ5fgibm/y7Ta0dr6m7QTtOn/Oxc3Tfuhxje6NeKP7jrU8dSyalbB6PoLf2SaeEx+d1qGs
0UslPWxyUNLDEU28bqBXPa9Z5r/OsaVWLHGRN4NS2OVSgQuDCTIs8gmQ6LIyTr6mXiR+2jV7Swvo
6fk97Mmc8CWSBnKMzHi1eia0pwSiQwoqEWBTaHcu+R6hIfDkg/9Yrfxhi9Xt4VSVhrsImK7eRHA6
wwSQNrO0+0+1/4dL6nD0uK9XLzHBexdKQv6tN3VA7wonFUh5duBzH7wiWwkG8zhbB8enILSkdQwb
MUlr3W23U2/MYB6/Cb2lbgeNObmpSKmLFWGj+RkOM2qIwP9M/iyiRNQMl1gY9mAZwIWl7Lhp1B4N
V81N09GAVczGICCwgkX3wQ4pLRDnEYhTHWSvNBpzrhl/ahTorlJPdAfu4NXlqXIVepZmxIjDVFHV
QbKrEnvJBinF4zmXqBSqJHk4v7S67LfyZNBGL1ElZdMgW+9xTfV1bqJeo5FyP/ZHGYBJLq6NWCTO
rhcYELI6HI5ix4/uYzSqJXP2gqtS6pyd3Jd+bTHwpM55GAov6z9A3q3boqGwjv26HCtboi4jMJWA
FbFSPwDwm+BvfDWKQvxxTWmmuLw11Ebd2P/8gH46mcDSg/tf+Oiovkl1WGzx48Jlv97boX2adWDR
CBF1W51KkqUk7vSsWekJxkvKkbBpFQWce+bmpDvN1Zh8BUZ08fhL1w6U+wWGH7BntNXRviCUpNuy
c9JYv5eHMBjVgbXCgTrg1TGjJrriiV0tViuWhh5NCmhZQOFVD9qB2W8H4+Gpt3kh2pFbazl2WqLz
q9YrZfzJApWyhncx1H3Ji6zwcUpvSwukBc+0apyPgM6QHfXZFxTRxsTcBPAImw+Q1YIDE2oGJs+x
rzCjRb8R1u9cvw4nmH19PcYuU9j66o9uYyrGpRXGkGfX+7ff/WfddIfvIjmcSP3PKtwjQhgJnsi7
hwkcFmPv8mVZA08UikbDh1lu8xe1LWbjvBfuETgDpql54BQlpuC0KIRkkp6PKEBTQI3LD4WbIb3F
SN3loiNNeaprCD4ATSYqeWGh5pTwdmk82Mab87RhJthbJugA3Kds7eyJfdY/WdT9pOUTBd+Y5xZJ
G9q+K6gQuEyqCxIff2LRJ75ukAagnse1eW8Am8z0P3nfqNRI+j+/7S84anwPUHB8qciwG7MOP8bQ
yO2gQ7U7cW0LCQOKp1duhNk9GSXRXejAKgs1n43kbWBk56c9YBK4U7/NngkTmB5+AEncK0XY88Wh
S/ofzwXMbNk8uG3YA7CYE98ln+84+9OaNyhTCJPip/YfVAIQZZTZ/ktkv4LBA5kejn+gOGre+I2Z
bVHKyWpNi9mmeggJ9Ze/LwST06gRzZfdOa6d8DW4cn14N/lsUHwJF264P/dpDe7M8mU34i5tFWxW
xBcKri3kjc5WHbc7yUIGEg+RkMxlWLGjATdSEKv2snXBWy0GIVY/4Nez7/HS6skRUpenUto7nPy7
OKio5MRjpLNLDf702ZjQ5MbxjPilW3uWhBaiJMbqWZ6VmM9U1XJ4ZFz41/6Dv1jwvsY5fpHdqEHS
YtUYs/cT7EfoO3/vVx7I49ExQUxrqvQqD7V0AkduKvtkVYH+aSA6VeT/i3yJM5N0FqDaIy0EfM67
ZkuKL9L4bGhOzVcQbktZIvtqCIfCkRxDhgFqC0IHQ8rEMhdGc9+8CA7VCFTyLmLGyxjR7Bc3kWNR
emNysEKUg3HaaJtgjVC70F09LtAHxa9BhvWeWOQBhl2Ovo1TREWag2nlGAc/b7q8L0NKnHQmrim9
DQ15VGNgPCvzwR+AxW/fIe72Cb8c4SCLsUzIDoDklluJgzMaBn6hvWxUUmly8Vby/i7Yrbhc2bmv
DeRmvTRcIVomLxi38uZNd7Tngmcb5fkaqMlRnKVU9l0z5hSJVkz2stVz3Fq+IUPMdUp58W496O+C
JoGVewedUHr+6ruO7w+nhrik072zffp2ELRfCEia8d5QgnUwCx0s01Pa59CL0qYNwvZQZnBlvJPl
M7B5Zpacl/yiONFzACZG/l2vcnK/Js1cxR+BltvkqjLhaiT93ERpjUvPUgq+ClN/8hdXzx9ELzQ/
F4wpo5FR1/WaX3Kn6FXJBFLFkvpbprA4kG42vdX+UZ02aZ95pc9Q5nUnBKH1N/9MCmzuckYzOQr0
mSbUPIOtOHcs6ZctcXO1Bxy0XhnOQy6qnophYgsoPVmP/0nfBlWk8F7BglCKUJyYpMdA20Xzoc1N
inJUeGgVs2f+wTcSwyqe7A7iI1bYJx40FBXhyU2OioDrwsJHxAiGY4rl6eTtqtWEvSZXvFXiD9f4
HsbZwwOO0Uzb1aaBbIElq3nwjK7MoRwWjF1V66OKxV3DPCqISVWKzLCKkLGXWUgv0jDirfaSte39
mQ5gfHwFk7n8hf3OO+OOj0g9ZCKsEduHxC3FB4pUxyjDw7+VxZHiK+8FHCSd0m/ePRsHERDCK1+H
cYKW2VVqvAc52GKWzg28k9XDNhoqyYEIv4W7jG6AR/sjbh7iogEyIlxnNev35sqRsViODbuVjdxZ
UlpevgAHlPEyiNUp7UL/lkAV35QCLTaO+ZmDAVdxPYtwKfJoMLHvno50tvds6WJaBdU5cmwJrEUP
CIQOnzTQG4AYFt1GBIWSJIfrv7logudoe87HJ0LtPskX2dYNDXGsJS0dx1Yo+iJOs7+C+d/11iMI
buLfP5MjYBhJNZSEMvshKa8IbgIKcSMSdGhVQYr8f5RKnqEI13kTqEB706bLF/oOS/iIKijGW8PK
cuvfc2RevGnKQ8HXiOI2FT327HDFQJwwCQIaFSavczrmZBPVlOJgBCMOkfmf0Oy9AWB+C7e4dObw
80isYKJOn9G66XnScQFIL6eKrsww+Dhht0kSoG4tZfWXQgpy7q3K/IFY+nkGj58t+iIxhIn55Err
1rjycxtV0TQ7PkNbz8ZpBy6FC45AFWJd7AN+RV6lbfgVizLW9JrdZVNil8ZSyd3oIaQbZGhGsvVx
OYopKjWAHaKLJ7Mgo4sQgAjz3i6WqGbZ9Qxsfg00VBGBsxPwt9Xrb7qvnSRaA9tLyHkoyCxRSqmt
Xfm4zrYOXkMiCvHM7CI5GitOPGI7tWHC42S1LNrNwwFtHC7Yx7AnSdVi/3wPOkC4HxvaPwGgceT8
1Hz4XSihOUKriQmmeHLMA9uT5l2oF5Vdrbw81mxrojdMFBDflvZrXMGEtgn5UM68/ZU/vkrupHkP
S1LRMPGAMEocFmgu2DE6Y0T53KRDW0tYGIBNBU3LweEbJDBBblk8t2kkk6Pqh9dkvLqynfifVx7D
ZGJhgHUz3rUn5xZc0Rto0dg85i8q1uH+/KdRGOcxxrZKD0PiXMMFlpMT2LQ/35xng+0NKL/jC64s
r89982jTQ3YT04b7+HB6vpZzAg71h1rxyMy2titTqAImA3kVw6izk24sXwWFKH3VVrmnbo5ywYZI
suqZEMh8OOiFZIlUG1O3jiybwHXjEGkwOMuwNT9f+1U/FwHHr6qYB3c7LfxQEYA49IO1F8ASBhaM
Q6kHzdxwC8iRkqN0W6J3N5kyGUe8VApu+SgS/4rBDaadoV5oQEKVUkbw5tW4Cec/tFm7JQiLEiZK
OXuNTluKI05QbCOLySKFqlSaeyJoiIboQd/9Cl9DN3+Cv26ED8oHILif3NGKplZzea/6vmIRhgm3
IFM5aMzn3Q4DdYsfWOmRtPZMNq/8ONQ4LASqkphdwYO/SX4xc7pn8HbG6g8Rzlt+5n7pVKpKRkWX
6CqFgsWyqpvDsXMpv/W9lMzIGodH3BnRClxdLkBZapWpk4ccBp071evCECw1RDIBS47zDcr2Bjao
SV8tjwa3MY8oDv6O4suYknKGjg0hHOjRUIptPzJrvEvaesOYNM3hS3OZWXYF6J5Sk3LjXAi3iQ/T
9Lv/Sw0xuDWf3Co0bCLu5Sm4s1aTS/ux0dsvj7BkMTy/d424tL0bTVV7BIOGcELFUJjiLnDpYh1h
3KLMr4tIIxQijCskp7lYgvoaiFhz64nNApTT6CZoZHqK5FAHe23LZbORph0WrtPhDFdr9xmTcirl
8kRlpmGRtMPNKgS+qIeVuMtVuucTaQ2fMhOoXS9xDGm3VDdl+8ZWnOjbMC7iGK5hdMy4Zxpb/is5
Et5uuqy6Oo9hmC+izju97NJVoO9i4AdjKFEK0qzsEZVr8fKOza5TznKeMu8hdFlhTyzsl75424U9
q+YRc22jyXhGnmdVUvMQ8dX2JY4f0x8hCVxD0oBaVR0q6FA1Ovz9FiwjguDmakSKtEagzLRG1q2j
vzZu1C0kFdxhjMnAD3T72U9Z0VXqrepfa65/XjE5/IOH+y3+mUxXJfJh4+ogC6Evb8PNRxkUJKjf
KZ9WM/5SHDNVQvFdMoDJf0BB68vZvZBBUXIA3J2sLbOXte3yetCYzhBOqHw2Wk+UUn61sl4sgAd5
BchtFMaDle2WOcnC0pKod2FKcrr6dXh+hfI/SX93WiUDLBAPFdmd72DrGdUqDHEV0OU0k2dceO3h
G7NWSW+hzaFf5o3VYPCQ2OEP3EjA8XJce4LgBFJGdLoJo1ZQjXs/eo4mlTsmCF/sI36WyUDJQt2F
mrF0IsNzAodMxuulj439xDVYrKNwgL0y00OoY+6p78GElGoEw1WPedF1zjcidP0jHWnUJdbvYzmy
RV7aX+UyMwuSltKVR54x9Kuje7L35tVjzesbs6FxcaIx7VaN3Q4lU7vdZH3C0uC81v2tWdNZ0I4I
L4DU0U7j0XVlwOrr8+hT9UkMdLq0VUU/M8T2NUoY+rUv747qrQ/AxEn0POvXoh1zviThGu+wBxCF
OxwRbkMZ4bW0zVO64UD/3+DKSeJacMIfQ4F7pbq/v1epXoWZbISAJVa4rQB1oWxh7oYXGidSoQVn
0hJTzYuIwy7+7oLabZaVUqU4sck6oDsGywJfib0GgUHhUGvIWYMTimJ4s4TRrL2ghRGxgYn4MwN9
t9XhBO+wHcrhXnFQq/Tpi172A93bYPB2CU1iLYHvx+lU4qqWghzlQb8moGpRZmcO0rqu8rSC/hHG
4gpgBks7qntkpfGNrWGQGMUNFfCBU+0qnEv2mkQ6wH98jspOLc+o4ssSkCfsX/INKWDVSepOnsve
EOL3VlG1v6VCPRvMalRkS84wB8zJbq/FGk57hIy7o36ubtMlpDFkIaQa3Slcdnu2YDrVALA6vnwz
+Vl0h/UNNsIl6Ybx032JlLJvZ7ShtrG/pPvbuUMJhKNBGieChjhdxiT/Bdn2UBGIknnfOfqgWw7r
eOSWKg8aPKnk3+wGigIGbU3DMfTA7Mk1/PsKGHC+cQT3D8hgTiePtHZU0pwAl6gANFVnFoTXdZS1
9MgQNppjDMJRWNh2/GC4nz6tgo94Hhdh/wFKgleGOSZslpEBgYyDS0gmRFuON1YVGKROzyWus0HG
CLyEiPEDeHQRbQLeDyrM6R8KyxcK7RkSsnZWO4A6jtxsJcMl9fghVp+vO7/1J02E+3mdIP+/Hme0
UggEYhV7kYizUqNxc9fypaYpVjEcd7mwl62gZ3dPmKPPAg+rhloohRJIcfjBz60Z4eHx/zR5x23T
MojCS53sqFtIe1wgJkh4XSeN+H3Gk7mzuFE3l5qmgFLY3c6FnarS86oAq8ByEM+ABBKF5RfF0edN
iNQkw9HA2Lweb5jKuEemmZzUCIOuQodK9xUil147AV2NusR04pd/rJYMdU/u+NeV05f+P73qPjSg
jjT/uf4LzZf0HPkA/0JGlLnprqtt6zf6xPbmayMxOwHFnBRWjgqJ6eQ2Utr2obJWKZ+T6+u+9Vod
N9J/Hf8u29CCRiprNcDiJfELs+yQOFBp5MaiGepak8XF+SrSW/h+tgW6YRrcf79/U8WFMgn60ao6
QpGjIlJW1RTA1yzMKL0KvMHTtqU3sGwthbmvD3C0MTuszq8+b31e+ftONXogVPlMcmbWBLPujKZz
rSrYNRs6lk0jfxsDDP+yRO9CTrHZW1fe93GcyTPLdKO3qmXVjZZsuIXYXU5Vyy/cb7xR6fX/o/Vt
meF7IPg78Dr3upKj8bKthipLPbTqIJnoHIpVjMa1uS+YuPgtCogqNnGyce6GLXUj9MXXkliMyLdD
KuohBvzjP1kCZSKzLhrGkdQ0YkShvUumOGw5YMIG2ERiiQOTZTgkFmJolVgYA0mTH1zxMQpWP8Cl
E63xaIf0dNn1ORkjGW2beMoloSAkXNX+EfmG+rt4TErL//KPHMc3dLj1MJ0LzAeMO24ryZpipxGY
AmQrZq1SodHo287PIFnyzoDpOka9WtYK8sANLdbGOs7sZ5K0osG/dJO05JYAIKxhrAetpQYo80iy
+k1r3wjEJBXDBdrvYUy/9H7xwHzeFhEtKP6FyvnsDDyETojMllT8TeaXELYDnlmt/oVwsAIIMdMH
yXL0vwVg8RgcVnEU11eihTLWLXDOJiBorQKWieroVx0eKL4BD3RSvZmX3CaHo3pcKbeRhvpIBxId
4TjhQc9uiYhBv0qvqSaKKA0h4iUan+8mRnK0lfFUzMwRGDxGsTN9fHcXcvry9PO5uY6S+/TCmSp4
ObhoWsizEjwmHXBuDMF4dKYdRdsSB5uvO3jHy0tCe9E8To2+2qrlRSTpyxmkKa5jzyMhJ0UQCukX
OwlYcnq67j3KbIjgpOpO7Or7rE0K99ic39oRQZ+LxhGQ/sXkNjuicdzdjqVZpPIM7r2e6hUdI9/J
RhGJ0pgUL/enDGiDXEMTf7uy9SaU4mgt7lxMvTW4JYmwYYNJh0SHMYJFEyPFywA5PH+WgUhFB5eg
lcQuyVApKScWcuOOGxsDUoTdzn85Ia5k5ELphbNgXD77FGuz5xOdY0vrtDKk0dWtiNJnBOSQPbaQ
NYsdYL51tNgFeiFWR1uDgWR/hW34lrSF0PotUjuW5J9ka5745jRbW2cwIKkAHI0/Y1rY8ho5e6oQ
JQGSXAGrh77WFnIR6XQEZO9RAOaAeRPpA9RLSofN34/2ROXIWpmWi+2Ka19hk9ONuMxZcSvtK7Wk
ce8/dSOr2RxZZjhiL8c5OaIFouVwJpjmK75gwNSQ+XQEjvGSa2t3jOFvzcNCrlaKXXUJeNNtxPMO
AY/TD67ivvSpu/r/gYYE6Sj/yZVzkf0yr4PoEOerdcao5Ta6KQExOZ5IIu2jbwaFYRbNQ4YDwS+m
g72hwokJquc2UzBsOEb9xYuLgauk7U+HbEu7h+vQnzismYglUMmBKkN8e42Mbx8dduCAGREdoQz5
EODl2mx6c2rJCU0Otk/ZS6f/Rbb7Y932zwKF0JPnqjKXBq4ztmLTOFkwU1ViPIGwkbTWq84AZ4G6
DCls8aHCCHpUq/2EZYc6JwBxnaT4sBWtc+91svufs2IfrXrAp0ick5/Uvrnrovi/fxWWEQTIw6yv
vnDWAg1DSO7pSz7yTwHLtLzooOpSHDk6luU/P0BYfc1nv+DTb5lCcIRzHOZ0LSV0Yi53/0P4I+Ii
MNB+9GW/N8bRm43XoX7qkXRHnCHxFiJsQEEj5sbASh68iLNmW8+xHwxwRegd2XGw1BVRFRkC6X/8
M34cPsvg0/kyH7mnbSkf3jjsd3tAhffoeeoSSecKmDoXuDciKej1L030+hROvSEcWnUu84UH8G+8
kmNDV49PKkNnrP1kZcR7OdjVtnPfGFADjh/71Wfkpo3ECMQutX1M+65G+nJeKYGAuPzbwA7jhUTw
gt6/HpORhAYexfrlkB5/dC4dBdhDc6ObBxf55oYOj9mVLUYDLUhJAxqjdIXA1dJ0NcPK5RFVfWTk
XiBW50H7ILS02gz9hh20FwYXNgefXqT1Z5xbExzDnWisai9C9lbD0bQuW16T4/2xGRiJXa8tC1do
aozfHdMAVtNb6ufY2LoYQClnsCOzvOytIfm/jRdvmlMz22DccRM+FihsFSQgZAUvYvZXmqzKbFSm
t6Xcu9nF0jSezjUpC9pNP3eNPZHXatFhH2eDL60cnACJydKbOYQ2rQeqXK2May3cUevEZaV8/qV5
vXtyeIsY58QHrozXcMCJ1RL9yl9/BZ8yB8qB4uGcAW8riIJDgIMdVNqPC9IytM8iRbNT/eesTqLh
ezb+i5YJl962a4Rn/zHGpWHw68yAcBxYkcTOT3eeJLN7P2+37CGDihS3Wetnyw9lVdEjyjEFKV/S
+X7EoEyOxyZ8O30gQxf8etbKkTmuqPkECTwz6uKZ8FGpRxEEkqRsgZuTr+z+2EXNp4iCmQOiRcUW
5yebap4c0RS0EtDI3DSNWM60wK8dGF1Rwxkr42f/GLpXBbyKwcEbTodj5CZmaQ4q6XLbEQa46xWn
diM/nr3DqxgX64VBMQ5rTF2ZjsIZ/6WTD7qwv3XrIrTFQ8/aoAOSpPOfN6euOVyyGWqhGiei5Vum
ij+3kEp6/agcWUnfh8LuJHHPaT9tlXiDIcc0oZS24EFgqBkpQul8DQZ/Eo/aryCmJTWBkwOiUlR5
6wzh3OmW0JLRGUhR1JCEMFPsShBWTqMI7zqaLLN3X2jRPX1piyJV84phclYVoScWrgTCe1efBGks
+N4Lt4mddEjmPHRkb3fGl8hlYQdxOHvwWZQm1p2xdSeXShcdAOqLHMtIf16qFCvGYt7iunzrHICa
FIDI9tBD8wH4X8DZ6birjS4s2x1biY2QRnPlQWGbW5BBZX2cpPL5EHKJ9nRkws9fgTDoIIXXEo1M
I+RTbq+YKO1ZuZ8V+i40gb9ASU/VZMzOhoCOQtdRGMku3kURfd9fnrm0ALSJLfNf6wml4rcB7peC
OFsT78Qai2S/P9DKd+MkQ3lP1dD3QXqp7ttQSppao01mH1kv8MkOsAbWofS71NIRN0PksPJ3DSEu
fSzbFvCiSRGu2j68YHDJhuyD6nH6PVvvfPM9v2c8+GQ+sInChWFxfQBaXPxJbQ4sPg7Wi8LBB3Oy
JdQQnbOzynnkm3a5OAl+qd5CBmHirwjZ8IvYpJWk9G/oK0Ca/Y2ErHA0yJj5yyXd4zO7BSZF2uxT
1DL0v9eBGWtzXYhWByfr05m4yeLUNdFgFDZXmqP1PFL2b7FyRLr5fRv8QGb1bIRqzvYglO8PFE4m
t/BUjOTYw0s+Dt6fKJcfQJrq+Z0vT5LTzd6wwIHO5Z69nJ1fwTSdBfN4RQA3S4ShCd+tklIRqJ5p
YwiKhaNdbsYWsU2+2WljAr7y4RLDByP3mzKjPBquC4dR74lVWEoNSJ5jmpL4kdo30FnYT5/JkAL+
YUidjOKpcodu0hVXXKGPEha4cagJzDXcOoyRB/TlXwb8Ob+NAyW5fmajeT+g1GZivLwe9H5W8UT3
+mKleTIn31bdjYpfioeXffqmRg9+9LxTH75aE3FMVQk95PazZ+wYF6agkjTXr//wqBufntVGhQLa
HZmm6D9EbM2CNQE/gkxhCi8HJmq2okbZ331IOVkI/4+/45bCNau4hJsbHpvxTDRYWtjSWj7utp4s
3pk7V5nUszttvzoEKND+1z5imUA0e72ZuMZkCmDC3A8QntoCqxVzMud1oHn5Yr65RK9T/BiVW45X
BhJF6+euZ/7puuJdS5B42guNsZRs96SwfEOidkFqR9wKf9soCDFT38YzOQPa57a0pjt4G6XgeqYo
B5BIythY3nzC8588LAxuS908HD+8lRGbg5Qyzh4J2hD7BTQ2Mbi1TCogx2PIsoYBp4dSd++EkQOo
CWtHKBDubFcHbFOa6RsZihTJOk2FO8gTIOfZtJeVimiORk+G5qidrGJyNqaL7PFEX0RTAaeGGdNQ
S232rMDt4vTRpYYwJqlDQaR+ghpN8QzS7zRqt4auJdZJ0ulMN2i6p1y19aSrJikheWu9pknGxzlP
Mj4sfTMGLCYgVXVU5+ANP3PeRpPzNHD6pfX+SFAUN2ZmUTJTIJOSJ5PZqxPggxdWj4b2ZXmAMVb8
mdMdAvYRNR8VL55nqFFcUNaC54z3KwmNt3TKcEDvJzK8R/06OuwLj5asIVpqRs0Goj8wgIJHqISN
FaG7ccJiQTLjk9jmfrO3lYIjS2iD6LJtH+gYMEp3sEXbW2dVnTyDmAIojJzMHpEYTAtedQyyNfL9
l7gle98R4zLIbgXrR9PMItitt8XYCvWKJRldkav3GEsKzALSrUh6RjfJ/pQli4hlS0HKqoMnPRhe
fePjZ9SELHkM3hoMtxKJdkdNZUAd7BZ3Q0tYddMZbbcYzzcPqVpkRwCUDcgUEJsHNtquY2NXRrMO
sZ7bRGROfBCFjLC4k4h+BTibB6lQHllC9RV/iZoBn/jiItv0w8o7J0JmLwBcyz7t9vtcyAt+fumy
VFrIsT9v3cI9XizDZIM9Vt8vGWVlXAeL1IO9zFe8f2BvAAAFrVpyzPlKbwUO4KOCHWst7lsmvtl4
qQRzXLayqs2g/1vS96O47qVYMWwy0SHIx3XvDQrkLC1kwTVhC0rBRdwkQpHsx0Rba5GJez+2Oha6
naAvVeX3TVSOim18HEgmwZ8QMWQ+D1RjVA32f5jsZeHOCSmcq4dfIBqTDXf8XY+jhf63gDTVPJyi
3ol3eylcrViWBK0X8XKbg3XjpGyPdFHlhsyx6gMIeg+YLtgZ25QZS1D5J1M1ksQxMPE+K8CYgaa6
kKsQfNVH5L1ssprscKPyrTnaM85HcfiVJkAcHOVIMcgqQd4u6i6VIFkRPHQ88n/3ty59cGKnOgHS
5H24o2C5TFORp9QIsGJk3OkHH0j0lMFyarPEMK5Oa9CArYqsGY5rO686XYyYBpxGEM6X2U5yfqBW
RCHAlhiCZ+iCXmApsK0M4mrrAAjNwWEC/tC2O6UZ+NWg/7kHHNya+ibylEyGgdTLOHkn3NpnF3z8
U2lk4fTGOeW4D3mamBtLMnwB4Qi+LJ25hQLANuKNAyU0c/D1kzM8M4gxw3kYEGlmzP6Ypjw52oio
2+Qtg20VWtfE2BcpkJoY4wC94oGYp7DDmBWnVuKiI3Ek/MrzT5wDOkkgGnROIJ4cXkLAqHwbiEMT
aMfLXuIEBJ3F5stKIOB28HQkDi8uBbyp0qT5BtYD43HFVxZq3kFPow48gSSjCH5nq7yZBeqxLm2g
FOvFTYr2QTsTevxxqP/1jnHLAdPiEB+g9MPQUmmDHIa1j6/W5hWHoi6O+PQ4QFRnEB4jqfrI8R0k
A1QZiM59vUR1L4c2xCfMI2l9t+/7q1VJrEFc44YZZE7Dn2q/bshzdYUWxDWqKCM1rXRksEXUeCg6
BtF9jKZXbF9CBrFYfXMsBoPwrNo8pXcrO2wExnDGzuvCjfk5Xk6w2r1ZdZ2y6+pskmrZQ8cuWlZl
RYq0RDxSfg3EKG9xRmpeDd1c7s9KumMmK2q5hSTHQrSTU4idjwDwadWiTtMM1l5BLakqgLdCMsJt
4TZUgSvPxVOjjhPo7jsvUYGeq+LkQlAT3xneCcR7AMA/z1qddpC4zkz0nWCA660YIb7KFv0Oqd59
jDIDW4+xbwiDCBoidUNs2gUxtbHsakP0k4e29zlfZT8pBWVqBooBK82HWqsI/JZL+ki96Gkrz9M3
+Vt5uRZJ89vxDNAkBc3i1wcWiVBsnURGVH2pZul4iYixXaANThNLNKZ6LwGecgoiqGHCV8EPtxRJ
PZwRHnCPjfTVBI1kcR/56sWeh0aZzJrOQPvXGOfAG1AceaT9H6/TdMwlbKilhqS/mvR18R0oj5Q5
NHbqePvcGn3ycRszibD8kuh9atxuGXyfHYIz0IjxIj+Strd+g1Z2jzbmTNnC/CzTGaxwFNsODQp5
fMF337AUsUcAheRlCZLCysSaObzpGYerbH7CPQSzUeSuiy3YqLpu54mXAxSCgZ8p4rajo13uYXde
aC99nOQvljw+nU4+YdF7GwhaaQsQAs2MvdXgsguqIXmg/fw56rPq5WHo5Hyr5YQPJCOJ+ETqQM0w
oNyBNx04Cz1gYA5sWD2SoaKS1pu7LhjyXu3zYZC6eCepnmZOLzDDq7AltT58wYqgs/5d2/Asb4Ki
VDe3QmOpod9NGfOVFueHBDmvKZu5Qp932pq1hOWqWKTVyMHLWt6009t5k2NdImTI8qp90H5u/UMw
5o8xsoW5mKv6t7u2rnrRl95amzD8TuUXdGVh4BAvDlODShb/UIHLhIPJObVZkRjaIRhAQT5BcN/U
xlFxZczWlIKgR2z05KGuM7yIKQ9Zut+o9P+AY7Hrj2REP0bj58TVdcfR80D4ZZjsg8T39tkRnpZ0
UNBOW7LbbzarC6yajgM9plpVhQk6wHgylO5n6G9qTsUAkxYmbWYM8RNzs+EgA3xyDh3BI5/G1WlE
RhN1TaQQOIW44xu4pFM2YfnFp5pdpdJYiHS1tCci1Cr2xtBChcFG+rkWsf00zhkE7dMwdTg2dsIv
anyL7czlcfhNyGRBZ2FKYnlK/LAPJ2qgcTLq3aVK2eJ/Etf1Tekxlju/lT6L1VXN/Yd7F1EjLHlm
+H45rOoprCgOPNDUtXijpG7d73AOQbYkL/Z+26R4TJUzrD+DFrzmD+uA/NbMm+W1NkR/ZrmyGx8Q
vUsBlpFEQg6n/dxrX9/VFOPbJb/t+CEO1fUQCnQYOYnSefgTJs5OR9QdIddWutIaVZCJ4nQIpoEb
JpTwg4CYkZ2SdhgOdS7a0GxR7w1WchsZce/6nyLTHc82iMp5d4qYxn0tJhSRoJrpnCSRwRrI7Pzz
QDDK6/D2K7536kdWAhiDEUVmMWcCUVrU9y2ysqjITrcJ3YdR/rXY7qmtvgc4xEPkyUO+AOeR6PtG
lXPHLm9BautM6IJq2Hfz7X5EsUMznZ6apJCm3wRSC63L0H5lYukpGK6kKvC3TaKq1p+v6wm7zeOt
pj7CsJga6zNPzDSdLT36iTYNq03DFPZwe2HDdL1OZPh8G/r19kyVa8elIce0apH5AI1QND/olwbI
zJEiuL9H9APOMuuqseAwrzfKQbNM6M62sVCFF76rHSEwsbezWJC4h7yNC30FaiM9/soIq1stc6id
aKGiefDjLF1AmIytu4kCCYiqas403gSqk2ZRSx1rxD+DD6zaAw1fr9csQGPomAQtR1cR1mSz4inv
IPXbh9E32XMEfQakLoNxzvsBEOPTSWoAfmJVC5KcxBpxh3jeml1nehEZu7tnxBDJ9xZ4fMWOnzIj
+8njxaZKLnr3dm9qWeVk4iegNFheToRUqSxeIh5gpr0kozr3h5ZRxaE7hoZNWDsntNtVQK+J7i1K
KL7aaKqzGUTd8G0abnxRdefpMHc+rR2hTXVidIW0HmROu5DDyUgdumoNS2F3NsB/1E4lDsgZl0hh
y4pshWFHnNGgsauGwERaQGroPN6TOLCr0kCTZNoxX2KsJVYssRhWjjTLgNDUSjTLt9i2AopIznyK
2sfC8WpR/XYL2EG77Th2zW2qaAUz9Zt4VmpjRdZBU/CVIS1vX+cNAW50is2d4ls8FXgvP6cded0T
wXXPlUA+KLt9fsyi/7ZrEN+RDz1xUdbZ1+dnHJ4SHaO1PvMtjYG+fneXBKQnS163zpOtLqJQjUos
qQuIohNEIazS8ksLLdOr2YoeUbTCd1IuOGUwzSTRTTG7fSMqyOrRUyuEA9z5xKFEkUUWmfjNVIb9
5y4v/w+13ER3ZPe3U13LWGaQ1fVd2cWXXsMhTnlCppHDNAxBc8njUdpNC0K9Fg5QS4soJmVojoP5
3EDdmUjFAQu/vH4PNYex3phR/9Vst0C4XASQ6VqjKM7DHyLQDAuDIoeqpwxJZfmrDnn+xNjANraa
7aPua46pkWmV0A+Uae5QApuUgiEfck2icWQJuwV9MJ5t9uyTZwXvQdOyO9qVSgtdAaNGxyEJMXko
mxNSajPcAaZCMZB7wQxtH7bLZbGzEa21W80GcmsFGydUYv7nk+h1tm4rXxaqpAjisXiMXG5Ye5zd
QfwpNnobbg2hqe8yqZgOeMpDRRyw3n15IImIKVr4M9sSqo4vQsLC7aNpyeeMli+bdm0/yJNY60Ik
sYGNUSd5mY3Z7tr5tvKF35tiBO/C22RilkGSfAEaauh47gIqXM1FwT/xw06KcMsfRnU0vFc8fmRQ
64y5ix5/9sslg35dL24JJ5x9tj3CGzUmWXumIRDId89cvwqec/9s4oTh6RDUABC1j6mjZZyGWjw2
hTyuAkXkT4diNOvI+W8zONbzs5UhQjTEPB03ZqFDP4Ycrj/Uda5j1pD3EofPmeTJc6KEfiFz6UHk
5OP5lurTsEiE0UvqL7AWymoCUgmrGZf/M+al5WAW7adH00xUFvaMsBfeNwQ7htVOAoLb8bXC8Rht
GwWTZwXznCZvi6DhSBnSPSKycfjSM61HwcQLj6qXGHGJ9Tr4aflmDnLX6S0aSoIty4SxXhY6wjxf
5CS4ppTboKZdDhqXUIlzlpEQLppJmy+EzwFL2+1Beq9RmkVAX4sKOJUPQNjLDo6+W84ixD7uB7K1
PinygRKe7vUxhZeLlA2PZUkbtAVCFa9pfTSVxUzFgCHKY1UX9ghvnZTmA56XqBNAm6aRoedlNjph
WPbUohh5leHo7VCY0iXqmjb3Roi6/ZKkAw3fZ1Zdnee/wedxF2nWh+Zz7Hjhgs21I8BkoY41kUmu
3DJNbNCdM+VLioGHyGinAqfkyu5WNbVEgbkn8q7Stfha+6Pv7LjmVZE1Y/AJLQaAIhQkKQ/LPuMD
iN6G9zPq+WS9PBS1tnAmVSA63elVKD6EOPIzVMDC5uBphNBjkQgWN6anW/3scXTyAmxDViOkHqXP
ryxb/OSeIHQF/Pnp9VeSqFX1Y6L53SQpEvacfT8ejw2s8XSg+dBTLUcwgp1KbemqCCLiVnwTg+Nk
PUaPfcbte5uYvq61veIN4iDE0WZAepHOKYEvZ5JhhkOA++LOUT4Bz8MJpKbcdjQoCe0+l/frWBhK
Tv/IaYft2+6Wvl1mqeYE96FCurYLvSkZKLCwewRt8T3jJRnGzw1e7LhclXAiw+VqQLzykY8wPz7N
+Eq9Qjcb3AyKJb+uDY6RobIKj8O9coX0TOS2wlkH+JwS2m/JZsg4QMcz97XBnd0jGxgZwlp+WS0N
v7AZjo6RGeh50Q+1KPntRn+04reA8BYAHgw8baeQXdomhn8Gt14lJE8aL44GjDSJ0b0HsOWUm4jr
qUucKYtQaQRGCyT64z5xQyDMVqiCSUoE2FdA9zTBdzUUSwC9NyBHlox1nfllcySRSjeAHjZwH8ij
A5DD4DUpjQ887Q+d9UN3Ov2z6HMmgsOhjcljj0gXgaR7bgWtXHLvupgUMt5fTHD/6XAuC4ADGSEV
75JM+EhfIyiKN3YyCoqkJioZ8R8o3yDpnEil+FbKy4Cdy75ubh+i9GKNiwcoRRYW6RifVskE6XRz
/GNkp/w3NVgY14qqhXRYph7l5OD7DbzJ3UrKQPkXucAV5Njt/7VlEE4oX0nDdKCm6yk9Y/jJ3kl6
mackURlGOhkl6C7xPIhnAV58PywFEWFVVFqzHtYag+heJorUhsSvzgHtqwKIBO9wslmKtWM5oeo0
rISKbPfvIgmfcoZt5LTlVuSRCPKsyy3ZF7uK0wW0AlAl3nDPRTgsVJk2KwtK+0CF7vsW1zfg/BtJ
BqhudLvZCWrdLbjRBxmV7pYVO6YfSjDu7knoXD/nF2HUfKyoHpfMmxVKFUw2ZFz2yy3p0DP2UbS9
LR3FXcSuCG/lNkT6p0ITg5X+/l0RrPNyAdOpchQQgjfR6t33nw0k15o9/a0wdokjZFXiMCUhJfpW
HM7fFiUAgt26USFQ58cpJUVoY++02ShD4B0uhz9h/DliCIPHLQDNZM86CbPFl3Jgjt0U6pMjFm3B
uCu5C94vwqnjgt5gvXIz2qFWoDbP8xbfWFnqykOSHP32rgbEwL0/X5vtlejwF4L/bbjLF6ggnVt+
Hh1AQ5PjPB0plMvMlxUHzGF8MJkapTeo2NhL5CDWWsFp+nHTjNCI+Z/tMzoI3faLf8VBnSkfC08x
dWH+yYOd+vhGwwWDCCRXy+l3Z1s6WHX6byHLk39AAtk+z1xs6EtGNuIQYc0LaxXeF+qHeIuNpjJl
vALeLiuzwoH5cgPDTLtmSfHg9mB0K9DBleqzyO5IsUwESkwKi8aTRSABHaxoyiGVDbnaAWCqXBwj
Sd/pTLBu/A87kou5NFSlkQYNJvd2t+9yj7fi6LaurqPOtMhS7/7NG8xUTaho+2+eyCrqZROO//L/
5sXckJ95GunM2G5SMDkNBK0cWU0ItyjgStQ0OUYZi9e+RFvUfSPFqpRDNLOxxrCmxum7Ve9lT3hH
OY0w5ZfTZI+R9wuvfi82UDSCX4lqQkCWPMS/+kBejFz00A5vZdPzXODADOTcXwSw/II3E5fEj4ly
21MQeuMoDKOwgK5JGAdLIVaeNTnfivw+AFJaHzTc9XsqWMvEsPvO1lPKV0vTEz9I7Obk2p8uL+dk
2afHUiyivAHodD27TSCcnXn/FLtRH9o04ttnAZM9rQdJxbjszQwO/p2wRrGumnXr+dFk8OvyO8Is
RrW1Ct/R0kjIc0I4JnF3DiyBKF2lLCqpDxB3Wb3sy+AIL03OAhZCeQ/vhhn7erR6Xmqt4I9rUfco
Acv+L4fXq8N7YelA7FGY78+bXISN0+V8QBbY+BEa8jQr3Omy3z/2QeUJ9lI/7GITCnuwEH717EV6
ZLDeIpqyjycm8ylBlnpZRbdlc2FAoa1CB3mtEA1hE/7hTIfoUOz1tpz1yT+At1/yM+A1m71nxNCG
DMPn9bUbG25EgB17nG7sNQc5l0Ob7mZG6Y7b9aDKC2geYsTOZ8QLYeyf5fFOPU0nvl0plBzljU/T
QjN690W5TtNMIWERa0I9ELYWXFvuumOkPyZ69Zn4VjF9AIWLZbYuNak5YklNikdTBEbWABcAaEar
kBep/qugWZtbRqEltT3j4rW8Z7abWtEBsjl0M0a/KTFqmsT43+91Rz0siq7vwvcAyssCVpNjiv8j
ScKOq9rJS7QVqNomnVfOXkXxBwrDFYARLgcGNzGSXSB/4SrsAzzmD3qT5GQhcSkGMlNF7wjbFIYm
66mj3U1wCQMI5+RDIuBNigfccyWyFvX5v219dl6Uqr2EYjag+8dQGOjByxn++TqeWze8thLfU1tL
ci1FZc90eF4LowGp1rPqfpGE1dLeMiRXq7PLvTHSdj/3aKPMr7i9J1fTqpWeL6qe/DkqADVCpLes
fgjT5cdKH4lU+bpw0aHd4owZNuLo9OoAPPyvpJVhnx+BjuMz89dIImagHtcwpZln81pGjc+cRyqN
VsbJHDJNotearuix18CMh6SVINTsqFyCJ5xzDPCYiCpRbyqXnnradXI5Dko4/ZrfOYTRNviAYtrn
1XjQiyFjq4RF0FmNwKpmSda2KOv0QaomCaIV7VvYIgr5udVQUyutmPANH//1RYExthQNHHGXtWRG
64i6nAwUCDR1KpKitW6lxlgPOU5mgbXGkYYrX6QqwzRWmUlqouLjLXc59xLJW2m8wQFVsVgUgkFf
AE4ejm1TmGR7dfQnIE0xXJbx57jPwLeg1eGj8Mwma+/d3TNLEX6MTxM5OoQpzshelm57BnS4xM2F
zjbb8ymNB/KbCgODvhh/tXPQBVRkrrEzZd6gMNr6xWjtNI9BTbVEejX28QDJMI0uqr2dfAJ35rFT
q1WOxd9+DzeWV9Kk7/SxdklNjmaiZJ11pRHRmkMFY/LsgkZKW9ewd4uKxaztJyJR7d48ag3jLwSj
tsAYCd6ChfpaNaWqaqVF+2QaioOjLusjsM0WYmlBBOSBLcrOiKINLvFoBrKWJuEQo3j+tYg/Mc1E
8kIkHnmuhtjVwFZlngLuVx9QF6pCwddxG0a1d24XDLwQ4TbnlFvN1CX2mmnc7YlbQyy6gNK67qqy
Jqnwu+FuUyXEoqMeeMxfcz/7Q5PKQBXRcBFGD4lk9j/52bSLkEq9vfBv3L51YpSpSkg0A2Ez2Ytx
kNl/pYmbl2fBBaqpraRkOp4Xan6ce2GVbW46Bw4N+0T1BSSSnKuvoAjoVNNOcimoEHOWB3+TC3qh
XLsU4m0CnCADRPPk6JmTHlWb17HX1t2LG/WGwP3+j37H4vFTZw5RQbb6X7GeF066MZIBoiejyzAj
0gQ+yQw7iRBxRLQ2iu6IhrZEMh5KbKB7JUIiwveKRVAQcVcmlXs770hXOGLCf0N8ILM7TB8eEnj5
D95pPSXnHuUbzG9cofbWVGtXWdLNS73j++cQ+Wan6s2e4XuWpNrriFJzoiRfkYdvlxpyGBirpPXS
TJkpD296b2a2QVtnCW1pwylcOEfWPoNIRrXCovUEONNvcFvougGUETTHydGBJOdqkmK5a9IfB1ME
Ovs2wK4ibEMRSvhZYaZEj7KGA6TUQo8yvCFk4wIMHzJ2hMozK76DXDngLpi26pTzK6B0oF90I0mt
JLjada1BqvYYfPxx2gATAVPhBLH6EJI7w6RaiTfYnw7NrzfNxKsP5BTLXkvYofF/sm6wxZk5sF84
ePlQ/Z36PWHjE5fmy7SrqATnY5radreqAfxkol0OBitKf+SaLRXq/oAsbR46rGPzkP46QL5w7E3Q
j5o3BgjkC1gbR/tj30XKCbkOsvShj7eYYGMSVId+8eZQTl23bUQ50xYUJVbTj/Ef/PE/jwAX6Ief
Hyy9YoQ+EbHaDtT44TFYnYTYLozgRykXs0KowtTEEgcUwa/+YqEV5BiDHX0Pt+v2yk/0Bz0AcvRH
WqkG3S1f9r+3Ui0XVPAmaTckic689x+zOhwewRrw7WiTw5ysI81nw0XrzVANpL1oWLi0fPvHNUhs
1BrWnjRdbuwUBcngeB9UxEJaLTah8fr75YMck86wkLFBulLlyS6ky8GLhiZYdQ67axW1Wo32IQcm
FTGeXDK7c1WeUwbqHHfaHUoVOOUP7aDyTrwKw4dWJl1lKoFhceyJMJsi2K1RKBLTD+1mamT3PjEf
YlcMjQNreZ59b8Rz/X4H9biZ1hgnUwFcrGieuQhExkeCmqrA+l12z0/n9RwiFeu4PPC1bguxmF9+
WokkB7VeBNrh2C56yGUhLbXMQvXMwqIDaitFCr3/KwiBZs2jXdCkrHou3BTCsDttsE7OAG2wXjox
6ZWJeaCf7ytT1X3KqFmZrwFziAYIrpQwFJZtrqAlc+uxUpTq35HxYes+PEkpwxVwy0sx2YAn84PN
/K1gA9lzXbajUjKht0GJqcBT3E3nCfreLExhy2jR2at4WhSDCIppT6vEkueqwPDCqN26+O2em33o
ED4sR28s/P5avrsTiYmLAucHmyWlBLvvjNJ/XkPQj+4st/FHlED+Vd1VXMhGCDUkYs0BNl658Kue
elJYvgioQ+/3VgHtQCnIO6vCQ350yrVfuDLkyS9xOhLXkAJUNaDLWSEVOFXa+ExDWWryv31l3+3c
LSfI5Z5Kjp3nDBDW9J0zS412ZDFvDbMob0lPCu/Xjipj09JIc9IT8E8vjHg0el4+GvtViLNIFz0/
2En0nZPluRtL3RtPSnxDcfS2jmm7L+rqzxK5yio6FVrAWRSECpWKyfTunVuY6dxShnbZaYNwZr7I
YYCOsd45Wn2DSd0fw7HRi3lgugNg6a0BWklX1NVFODC9eBk3zei9NfK2SUZA5NGQYO+BS6kLQqyl
35tjyRNgVjYiTtEajrEsTsn7xtnsCweZLAQg/efW7bmj4Y4IS/9bj8PdcLEEh+NtOkCx5kr3lJoZ
2Z1heJrJBNWIrUZjFELyROlkAkGhyslbl6guvaiJIrJUqTytkdX0r//d9mMGDPvzMiGBPKw43K5a
VLRVLIrpkJPZmUKZtZz735GdJ2JKMRmUsdmq0cZ0zBe6BX8PsdkH1TfEQtUJMaFJiuZj9Arx/zus
pKyplUTjvdioNJY5mY6ki7NVq5r31se/zt4KhXRTJsO9V53gkYFSM7NkmQ3vsTp3Lz3qz6hWFkl8
+VRY0kYE5f2e1OrLtA2K4LHuZDepPKGlsHgMx+DnVAh3tju2+Dadc0aBWnSBn04O2kLR4WnZUu2z
l4gmg+Pb8pLKk7N67zUIoVEaXFUyQBkHgRK0UbUElJ0fHKmApFQd1GJfp7IgB/OoDC+A59lW+kE4
udvUqKE5C9FN5EdwBTiLTXnfB7zLR8pnTxBRUbzJ9Uxy79T+G+JTFbe1nzPBz83tD+xRj7d+nvCA
URE6QiSeYggCycGyF5zw26iCC1LJbhL63ewnogwzHKUIl0wgF5nbWMInrvr+wNia7Ddny5ZH/c5L
50zdyGBkQIk1ZgrmzfF0MM/tJKpHfQuHNhIuI9p75++R26INd5kgf3lzW09AzD+s1V0eoYQ7ZvLA
u00RPklakIO5EEOIf9gepnFjRER4IeDZY/U5Eh45MyPE42PKWx/SZqZVMaRZpnsKQktE84IXqrLU
AXU4bTYk6U/8GreSGQ7bblq0SyBMJLaniAg9H7Md3/WRXiYRyUxLB8SWrkq9ZyhZLxw4cHo1DxaO
5wq6ymqeeOQk+4SolgUTpeSQHkcRqvH1Tf1F0FiJ39FT7aYz63zprdt03yRDJxV3Gx+qhSAWVW1X
m2ttnN3YIQmZ/Wu7cDy58H9bamjfzID/YX65GCetcbM3oDXbcKcPB5gxswWc4iwy3i33mHTI+FOz
gLiqeTI5d7AjzfqOI4G7M5Iq8p/YGwZGofKVI/C6SMsTEj3M9ZyHhZfbSx/KV/in7kRlcH+IR9V9
7YBEopHnn7Xro8BjLmCUSQgVNiNev0XP389U9YYG2isWC1jDVqvM9puY8lZ/ZgDBEeBYeyn9vBzs
ueQR3IWTjOuzShh+6ptpd2LQpYWrGBoLpLa3kg/Cgw4U10kVhx8VtlliHmD0sLZ25NnFnijj/u1t
zdG+NsNWLut1B25IrmQxwghgslVHiYe8WbVPuj13cs38Vndh/z7XncpUA1LrOSDQh6b233e8LofV
P5UY/p8RJ8BoeFDUNEKsFHhMMAox/ycgKTAYD3Xq5F7W3RwTqy0yXRr0h5wtVU6elEUh77UdlyrI
LcMaMPsDP/kossOpOC0/h7+nbEyub+wH0NwFRQgAbii0VWbt4tGL0qrVDb7anNoIWUeClhjUpdoO
0b/GfCZdB8Xmx1WngcbcRSstoiB4wtUXvZHv7Ou/KGk1WViNdNyQWlZiJEbxdL7Of3N/Li8VUxdZ
77y6191Rg96jQ+S9uAkaaE+wZqTE4CYGs/5ZheNwoGka6AvllkKLP9vE5NxRG2PwhxIlcSnGK4jU
fqTR6hquhnLuHLcd44IcLmDVntVUf51XB7rbRpAV8NOBgUgm3sj/Qu+FCOdC66yOA3rnWVRQhmGQ
iiHcSTwvVy31XOC5/+yOqiaVI/AX6NajB0MzqAXHKwye3Zb6z6zZOX2qXVLNiSM/VcZhOydXTPfn
IrpzXDarvwvvDVBraJKSOZnh4u5nTkMsKM88q62KjMBfuHhQwQZ9Ag/2uwqhBGbff+1srFuEGZdU
IoGvJ/RRvkKoUOAb8kXlI5OU+ecN+9O1l4tswysvbOHTEAZpGX8d6Y2cYzdKCyUekRbBl4RjoNLM
QyBFXL1w0MP5QbpepPp6j6tq4yejuFQG6XxZJsh9N2VUAUARrXwlUidmweIzqKpITl+zivAkJ41n
QkmCF9fdvyR4qvUqo77St1K7iKS0JyY5CquJrk8NzSSj6eHrhOAu9yABg5L0FqEW2iAvkOFpmJl9
Pst6cGdC+gvl/xWfbd58qxK6GZj7s680jDgEGpefrmrhmMcjW1IsQu7v956tT6EndiY0Bw/RQTrX
WB1ssjx0I8G2yop+047OpCuANIXxqx2AnRUE234Eg15d1f0hn18bQ8efodIKEKaybElsSylHsYPO
/hgjYd21BzgDYIkxlyARRz2pPgZJ1ta6ZEYKc4N/GD+O2qhYDJ08bjw21jDweVoxC6GjvD36fDCs
FyiWB8YRZ3JI52Vv0SUq0L6KWy9LnK6dGPb5dniZMym2AKfctCKJuD3tyU3HJN/44F4ChWdBx8a9
UeYpubvaMtZ2ukP4SRMofnPFX+S7+KFs5C819ERGxeiOdIIhuSQ3EiMDCjUuFFcme0coP9WllZ4i
lNLGk6RRJvMoMSfvi2Tcoh5V6ipuZFDihI5aQn6UN3QOv8y18XSiXW6HKkDEDZfXK0sMdJ/bQa9N
9ayXWGp4xAI8jaS2I40Pk8juvELfIhV3XYm8Vu2oRh9upd3VBsmccaESfWRKdqZ7dIsHRrO0BBiX
92ycwb/ISqYgHk1Q4+U/Tc18qrEjW1aR5wQgNnz1nzbaMNF57X8UrdFCIFlMXQFjvMSoLOhlab0f
0vNtG62b+Lt2CwxyqBxeLH+jc5CQ9XCTDDcKeTdQoAstEQntcBr0pMUhReT5/i3TSYvSb6xDnT+I
MRrfdni2h36e5a+TvfWYzESmfMbBDd4xqe4J0KyPYwrMHJ0LT1V4z5Q61x6vBzhDXKz58cw4tyQc
nPHEEDSrch5m9JHOh00+K+fHdJXoNhrRcwvQu3+7oHF466ZJ4ZmuXy+B/Q8W/eJ1ZIcOo+XJNx2E
m5gGaNUb5zmeqnM/fTD/8fx45B0YNrA9WZ8NbrI3lXaXmFQdPxL3ewg+5bGSth9rjW2xODF4Zx8k
kigR9Rq4iK+tZ0nmeIDTTbdBsTSS813t742mY43UOwACuOvCb4Bz/6qXFcuMm+QsC37Gzm6gxUSY
GOg2msf9CprD+qsLPZsa53yB2m7FJAj/TdyHkcWI4eKIkW/SV1vObaAVW+2GrttYT+BGHl7q9g94
E2q7k8mSMVpNtDdQJqdmphg9ygQ79QvMEtnMbx7eWIi99p2/6v4k1qrigNwHsiW6bt7+gC0Fgbn+
lDb6a/8vufgvu083AfW7PPSRnZfWx4nr5ZaIpXbxfg1zSTmaHvK5qX1oa9vXunbWGP47Mww5NeB7
niCVoph9PkEncrErwEJJDEGferFNuaXACdHttZxwa3cPlrM+Vu/YdVmPIMFBkIV50MAe/0SU8A3L
abdTP/qUA46OlT2hEJFWu4BVqE+kcfZNHjBruNPVdhMjZqXxqJCaCm6cMXuhINB/CoA0SVLuEeg9
AL/+Knl9WXx66wh7MGzQf7IZT2Chlh7Lu3rDLEJlklApzlFOnFKUJdzc7DIawgSKvZQcFJdOgt6w
uGQ41J5PoQGs4DPa+sql+llddoDUWRwBxycLfzynfY/dXILd8OaGbrQnGGPTPS0dpkqM61A6nTlt
TiNApzpbkasb+QRiW5TTyPYTpmlXg3ry1cWu9jPzF+nScDLZlxKk4xq+mX4/rHE0Cgy0PWxviEEi
tKENwm1B6CAQ6uWqpyr8Wgbffq47r2Nr4bhD+CydrzdY1GlZtkE303C13i5bFbQbZUlTtN2gFmKc
+pkoLOMj//ww1jSqYqj13UVaaWp8+P1lNm+YO3+iMgFONH+aLAGBL9Z9f6qHwAALVh9B0EZdKLPY
RketcloOBoKGctjtEOJTLQu206Olgkv0OGTc/YKijz3REeVBBqIogFAhRFuwEEM4+glJ00Az8h4Y
MiHD+hWBxLKUxmnpI4xYt7yC1/oRwyfP2bPamqROekmeQDtAOW9jJrcoNtkVvoRmIv7YYn5Bv9RX
BJlqKYZGRDNFuqKwHqzAHnrxhTHAXI/rpc0YXEOP3/w+ek3RAz9tFOeMI+RXflmsvPLj8ZVUspCh
7vLW8cZ9uy/f7IKJIhNSH89aoAdub4umm6vU5OfSZpbHA+6gMNJmAfd29mCDxod9WqfbgRvc2/1P
6EKWcPBIMdABdCRjF3ptXQ/cU9oHM8/OV7yyBjDWS4218kewhmDaxwd91tE0gW03K8lvjW5F7fDh
xxy020hlKCwckZj8WLnPKv8utPdSFPphZMLFkhKkvrPfabsNr9Zb63M360ue6J2mXvb1y/m+pNpJ
B2aVO0qgyw528cN2+aiwI5h+sta299bmGU5Uwk/TpZ8uZgiu3sGqMl45EFGe9+uGBPVX1qsOvar1
kKzFqRRcYUCPZVkuKEu//ofIzgOqJympoULrHy0l4PTMleKPaJ0llCZ7N4G/PuS/1/QftJxZMht4
aCMrmM9udnw0LZN0qg51UXTFiIZZPlJh4qImagBrp3gSklB9sOGp/MHCR9O3HJAm29E2R1qkgf6Z
RbKP5FTG7WFXXB7frmQocSHkpVNQYa2z/yNjr3ZDDfr8eOaEO7Htj/Yoib/Q91iVar8mR7h30tjK
NaGCYQnc8uquMMVdivM3qTosB10RzAdwKWOKsNEmHXeg2E1P7V5rHthmQlzKkrTyIWlWitc+Lwtj
4P96b+z4SZX5+03eWxhk529sPtnHnyrITpcfg/3ecj8tYkfdVsn//sXINbSZiiSS3TrkEP9SRN8Q
EV8FoUGOSuX/m9bzpM+VVELEThnB6jPPsGP+eQMKCL4pVJ40dQ0OLQVzYD/mUSoNwn60jJYYPG9h
nr38ZVDuk/GbzDW4+W67GV1C55pSPpK7YD+rd55yw/3PmcU0iwG+lkAbuWeEY+dwB6qx+3gxh8Rq
DT5AuwD9KgF6e7a25kKtz61bTiZmtpMUrvPb4Pny6HBhy+8DRYCfA8UZRfikfnb7ThjzS2FZX4f2
Wopc5hpWDZI7ngU5NiYjq5E7IB06RxUD1OC8I1S/DFnJ20Qt1RjHxAR5vMmq/+yLVBrK8UPv/127
LRJ3Q2iPvlEtZBO8+MClB08YbyJInjc4XGCPtseydJVVRqW7hO7ml67/pjKlBHSFgbGNHlP5EFRY
TDRbec8M+BPAir8suv9rQ3PohAHwEGvhxDSrxkLdtfNKGBm8vIeA4jyJgdwpim/Nw75dWTcwPQnA
4zd+pT/f0ux1/bvfhvFo8LAKIMpRV7/eaX7kl45HnoaCBouTHc8bV3g++vt4asW/PwU/bo+vJXBd
vdlrTAczworDV5hgZaGQjxd9/PH0b1rnDDJ9EUpLV7pUBBzpBgNknP1JLjCR2NUeyqmX/ggxewof
mFFLiOHKQcD/Eca3o8aheJfFBQWyRPOErQ3coQ8yQ+RToVLj+nvfrP24kAy0WLl8QByhEbOorrRt
9h/wGvbpSaoCKAmpW+Y3PAKW5YaETNYZlc/Q8R6o63kWxmqmaU51H1ZVia0J43HPumW4/ZRSL5o3
gO+d+YT6H9iXELo8SuYuPzyWW/dAshjsGE/A9W8tH3o5A5R5h00AmJk8yUr1OOBfys+5WHKj10P7
ElbDVups543diOVF+IUZrSp4SHVGwICJrMSaQGbF35Q3/u8x6CbP2BZ0diT/DGF1/ii5L1xOcshV
LctrgO0iicbNsv5AGr68vo+V4N5oGg3uBYYcJMCqSO5b8gEVtKZLve+nXon4YlgiFlu57jIO3AEj
azJepryUXxmq6w11hGhw0rCWjJecwyC3QIbuELnxhWcH+UgnCtldKcXeLWgHKXi0k1ANjfpVRmVx
kQCT0j4+eFTHmHtjutJ7Ym9jKZZrFYi2JENSenFfRWJImhZ1SFrwbVTh4eCDQcRu88cXDEhOyA7+
LP1IRwmj3ArUEmhe7srGkvtPFvXhu+5sfkRFkcnLiHzcLCLFGWuPo4+vKMs/XO4GeXzI0wJpWJPg
lhLndX390b+O8ftSpA82+JQ3IC7548Q5iH68mhKJfW6y+mCDsGs4VlZFVo893cH8GmSft8s+4/W2
hK+KCMqBsKNM6dGmIUG/PD4NpSrt7ziRgRlNU4T/x6Ne8EcTTe2zlKMAlvQ4FEXWQpQcGjEqGnxq
dFJEnyDkKWFV2WdgrJYu0H3XZ0aoOdLXxu9C4vzR8XG0OasNzVJZrRzwl1y/caI9PJH3nBZbPnNN
oAlQAgXC7dVtSIY7axRNTx47Ab89+t+U6ky1jI8BYhVR07X+c8zqK4L72ChHGmgPQfxm7WPgnVYE
sUnC5WLTN2JOFeElIsLWvBUcNHntL4c7IX48/3iE05LcDRTB/DDKNZ/MKLnLlSIpXrO2KujtOVT6
YpP/VbEq2HNdZB07KbRgTLlUN8RG7XdngXj9sbtUDI7IvHtKXUIDJvNd4f63/YvBnbdnX0HDcHh2
EKTEf3sw100lM6PE/rCg6tVMF17+/oeF+Y/0NbEMwLTKNqsxkNO9OtWTFSZCr+6M7YI84PU0qLxH
YRrjWV6YlIimNLBYg3hGurBAbq5P4YdEXn3d8mMj6Q7wyq1r/eBnzz6Qkngqk+nqa3+c/qkSXKw4
S1R7ju96h5LXlHuMaxezeubLxrJSTKGMiWq2tuijQYLD8HODz9to5EcqNX+s1QGzNxnSAPH+ayFf
6H+zFpe6yLxDkqAXR0Evh8XNmLhRbgFVkCLNS1yBMwoL2px5hTD5gqLEirg065ymVpiCumBfp3hH
LUdUeKE/0GP5pMjbxhb3dK5AltL8j+AWzn31bpZIoxHdMPr0+StQOx6aVlFJ1UNBEI5ZqxcP2qTG
ncrp0RZchQr3Wg5YLjdeH1pocErk5vADMUz3vtbz3Ypj5MYAwScSIpDUYjai1moHuIW0MjYM8bfZ
abipQFYewKqISueAT5pzU0pgX9lZNanPg9lRdPMj/WOHVagfNoDrn5AWgldriWkJ1v3a1+fTGLfC
d/pwAjVeQuiLfbHmr8ZzNMqGgeWkuXYSO1O1ZIW05ezrFApoA1uJpMfgrk5CeCRKgkoxl+HvgaTf
tWKZc3lnIAg4XYZyAJHQB9wX/ayghulTH2QW3F/v/D/S/rLXbOuUSi1nYszY8U9me/mdA/USA4y0
BI27fMEFeW8ozQV7+7oU+nGcu2NnN6tabClzm+aMu52sDSuDwWFbL0+4jIM1vVGAPkzAZ95/J41U
RAWcYOPMGTuAgn5ksNbmNk+kZ9h9B3UNUMU54zSaAMi0/h9IWY/mA3oeyPq3TeqPadUkSobNQym7
eSY90VQiar+VTNG2rK0sv3noBd+crlgN+/oDpEjqpDVrehbAAZRuKpxghMQ9liy+YlZtpmHxvJBE
IBiQ1rueR0Y/2j//Q4RnfxGiQWKbVshybgS+MiElYhNyibs8nqkG+JL8zqnH4uPkswdqx0xi4fjH
uLj7HVhe/ypUpSpjcy31a3WdiyuR9csUOnhpznLkRhBmkyioI/5gFsm8L88W9pmROHG1d96sYEkm
6MUBuJyDUw1HbkQf4naIWeQ1euFF3JRBoyHfnb/vN1m25XS/6RlK4ePeXqefUNrq+p+T/IWx2AKS
tVYoYyPi/FUNqjlZm7BnpNF4eLms0XstoX1bsZlMytDuH2fO62idfLLw3qJnhRorIIoU+SLyAdt9
YSMpV6JqK19zLGdljyV8xkydSUXJrUHn92rUR/AuIsKnkM7+v5MwGYGjEiHmQ/w4IzjUx9TPqdRC
Hf08Cso9WfumPblq7JjKwH6OWy9luBrZZxi3seBFjs8le0IAHKQLO1pM+6jhASp0bQdcnxXJakrx
8qKm8V7GnKxCr57POOe4kzlHBmavoIAa7vCn6x57b5m9AZpR8yXJ0Hu0GbcZchCWvRgskYsmxTyx
5SyY4X+q2tcr3wrZZYmVBni5nOwF60qZPbsvl5qJHazk+qR5hFXyaVcffEOP0+ZgjZNASQvJ20Ue
6Zf9v4X77dFyu5AWh+6LxsjvQhRHwn/W7vzntJV8lV2qTmxr95GFdfITcbp1Scigk7fOqUa5uF9n
fRLcZwOe7p77OvlNevm1Yl/b/3KEUuc4GS1gS62KnsakM+iDMzMk5UHkEtPp2QuTO6aVlOJRG4pG
ZGVX0mYr55bVJwNGEgH+FkojfWdDn+J7pou49tftyWwRMIbFF1JLO49fr/HQQj/tkQfp+gmy/v8r
bsJtoVIEo3oxndnS4vq/WpGNUzIdQ2daf0my74K3iGFqvKHm/fZHkxLGbE3sA3wFUGE0thQaI6Rt
QxrdAZUj8RQ178Q11QmstW24Vywr0EVH6i620Il+p2GEaxdZhKkcKTWPg59mIM4UbOEpxk8LdGRn
jdF35kD6A4RY8Y/sQSqIWAPHl4/aA7ib29Pc6yKGf4MmjPiGSLKyj+UPiuTnH+9F+xpLe9rXDxVi
0gJUU5gVKZtXyw8Jlk7/Jki98VjlZzfkDWNjHMtydP31PIdqB7TUiLfCHa9Wn5al23ElVOqTQ6Mo
NLjkOofHgyEp215xajPCSlYH+FONkblKTmAxIGROyKklLF+GD/I3yF+zyh0LCcdACxjCPEM/xhI6
WEK5lheQoegcm0UDKb6EPqTwfgnB+hZ3cA+xyNojaAqAQZdvKu6HaCc7qINMqPr5oDqjcAMlFU20
xIb66Klmz9j3PxdOymcQIyNE0tyJ1iTfx4GoOxXw+MW6ipuj01IYBjJljmcwKyl/3FJQAYtoefgk
Q8BRpIdsZGcwabljlc6q444ACH/qRRmre54SGqg51mIriaFxA01v26N35pchfAfTeAKgA1Dq5sW9
d9FVMbDGRGoiwmiHTkCBiqfDkDnuKgrhfM6t0Sx/3YtvD+eYI50ejQ4QKquQz4CKrWMfZ+FTgrNx
3HB9eY8a3pIlJE/cqGcxHIgiaNyqD7XtWZQE66rajNSvR63XzfMNCp6A3sFoD0ltyixSWP46rJev
pupIwBiCOdP1qoJ0pOLkVVtYAz05Ikn+zKjpIOmb/tWMO7vxMUtIImPbuB2WS4PryN1TCySnych9
NRBkU2e7IHcypCMJ7MQwa1Eyq0oRj/kXASYctMIOHQd6dR+RDyG+rVOiXfiUlzGxIx4LayUu3EEv
WUGEz1N9LYiIV7s0QG6+7KA2W954ms1Qr7+DlLekY/s8ejfe2anYzgBM+sfidvENunyyC9JOZ1NM
Pv6WuALp3QT5lOE9pg+/2FQb2YhWrxhcvobM2CUFoogpHOTnQarQBjTYslP4Zc/YSQHlXw0U3Ouc
EBn+V1K0EcUj2dL7O+RdzQxlXzkxkTuNarzXZ5glUkQa2XHEMG7K/rDfOdH1k7UfVPvSmoAkt3Kv
3J3mR+nSIZgF1cYNtNVo2H5mmWZ3QQtBm0xbo463TdbbwamUG9nihNj+Qvbv2au1fLMrMu5P1nWr
84cFMd10bVZX7GcmLFm3EORlRYa8TLxw9VOUSzk6ndw/0PiRDoiKdVTOXmLaI8loAfPcdX2KznCt
gIjNWhD8u69TdPZpq1xB+NcnpcmRw1SJi72m72Cx9EFnm0QybMipYX3Om6osrYc3xWsquxvMyJp1
LghdxSoMXIHFal0088ccrkNLpaduOEwjq0JhDCiF02JFQDvii1a6EB/Yv944V8t3ZqjbBQ2wYqXp
vEx7PidFNb6414UITXhYIcdQrcz/8GSeME49xK69uYUv8OXkb+yOENazKCkGATiaVtWaKHSGRgPN
4vMRgB2lW4EP7mzjfGK5B1w8CohkXa3BjmzlcFASz2qls+pGY2oyeUdk3Z9ZTePRLW0EHNq/uXxo
zssPfjPpp9pfEE97wAyZZG3/xAx0khxCenNrhIJ767mBu0potDWFTRHnq7BImCSpTGry5hbOQtsc
rAwgofDRYl3mvAsBc5equs0rXzFZ0ca98KmzQqt8ePPjg9g7DJalAAodngsmCeCOAXu8AtgKpgjB
GSr1ylTFZ9AxLQ5rm5tINGMmq3db9RwV2rmi9PQyzA/Yi17dICfrpEvmahKZRyuommX67R7Csg+a
8BTjtOr3USonv5bIQfkAuIDzCmx2QGGyJHN0VS3HD65BouhLE2pNI6vdEZ+EcJY3hCRO1kZXti6k
lyJdZixr/JDVWmGu742OSQ7BuV8OteKC1mLFFVG0waZAh/MurpLLjMzN9HwA+5/OiuLx93qJpS7f
MRa3LPu5fnKsntmXhem7iacnn1Fuox2qUldzEfzPuSdOpDuQk/vbj9zLzbMsksP7mZXjvA/eT9Ws
eTZyHDdgIsSkyzgE6A7YIVx3fuIIALUjP9iXfzVgoE+Iwtkyjb4M7utWA43xV827aytapTXLOGHB
IzFbNElElx9MYPE/mPoNVNnUTqnWvRDxIxGig/7QqO+t4d6aQuG6FeXkEsXMxqcz4uxCE8zOXU8s
HfmK1BFJ3BfxUA4wA1csJbCdaqpYoryJXe7D5HeW7N0gg7B8Jq8t8QjepuvwACFVZ668W+pzZ16U
kRnHn36n2dLVrC3RhDrKGxU/39Q14uAGEGMZGxxPukPvzTgx/Tt05Qa+Mskj9wbZ4N9eEbwV3O8f
9KD5kIOK0PMPufFIuZGWADs+z2AoJtxMgrVizxMOBY2302bFZUuUN6sMcREX3MYAofYB1YhZY1dc
+xYNUS2kBy/nddnwcc2K5/6VtK8iEal1QCCXWfJPnVKYt6WlenomqspkRe1A8NI0Ji6Mwi/V6gox
Og0YDDCwIhnQA/iUjFRtzl+jhfEdr8IB3qmBuCE4BaRT6KBTjp22gFZauQstzxRTMM8uiFxv9SKq
SXVe3hVecCnIuwOfoRsQqhzYA3QmQcfT21O+PI6sLjkxNqTaTvLaDd6IrttEdi+5XboNmTMOsntB
dhvaBily/4pm5hg5Gm1oEYgn8Ab88OHwb1+NZuc9XT+GyA+znAmPgvlgwXWfC9uoEfXjNjZiFn7V
ysuKUQl0tcLIgJkZBRBLDFKiw7q0vw91CzwRm+aJB4Yy4BGz9vM2Mr9hXfFgQnnEjN7KBvQbpLWp
bYq6E656Q+8g0wyKnf/aErljiIlAkLMSOWqi2ZOeFyWoGXm3Ow1PY7QWABMS8MNA8oftDJe2TJOv
Nx2HiJvYyYrOCn89sPP9O/50sj+7hC4BA1nyogsuI9fMYkeu9pQ644zLWsqf0npYaLOgkYgWguib
zUc7D5z8NdebrxlHj3DIaOi9JZIMhVA+69ZoRrZU0tbmtqG9eLVg0+4rr15hhyV0ByoE4wCtkisS
cay813YTLPPLER3+Zcpal3AdI99C4sY2QiFuU8cpsZsFxsiUX68OZPSHN2FMt9TrgFJBQ/qjrRwk
JX6B9pbq8p0eyc74cq66Zej7DZojxaHbqXodkh39xFYrT0UEgVEocDQoRB1E0FGCPj5pz0Jy7QF+
kMNs5C2/Rdn+MB5a0HzDnsDpbiB/GyM/4Ji8CKy3Oc02ML885+asE+4kIAkp1mDJEKNBxlprc4fG
sXuxSnlZjVQ17fxLjDPof7/AXBmOm8Rw4/rbfkiujqXs1cv620ySSjgiyM5Xpt2OM2Ay65ptQ7WB
aiV8UpNg2lronPN9ki/CrFCaZKu8B/En0a26e6rXOfvW0XE79wv32FfvRPY0Gz5lU88QTWR8Pw1J
jgZGkcDjXTywL4p34raHCD0kSCcMqdZbXU/tt9VMocMNWGgrWNgvBy3SxsTMd8sv/E2K50EZW9fj
jgi/DB+mlQkmFh/gX1ktEyrRABcVSf3p0hhe8cvc08/N0+KvhFJ9Y+gi/ZgjKlBceZ88Z04jxkDY
2Odf48aF/Dkx4TWlqAU5Mu8nD8/cmPcgb5qdqYN2ND6Xnw3v3cjS8KnZrq/El6jJOeaLENMDVcjF
NUD0z9vAdrKfeZgXfwOMVcBVrT8TfSiDEkT/G3Os73FUgavIm5E8UbcCWubePVX3ZYngFxjdtq/L
CWMlwbICotgKXSnsbGWPgrTv45wMogGbEZ1jsUWWJ001xB1qqxDbce5Lg1faLgkPdxU3KVAZ/T7A
fSaXc6t3hl405MFVBx7YAAq8nmH7YQtWTYmU7rRqvmGIDWF+8VLmglhEC2GIQ3aFNVbWZfZZVWlU
nz9PlURzlRMiuW8u1KCY4J2bmN5m6wdiuGNuz2NF9O2i4VawABYsL6/ocMECs5Hn2X/b7IrR1yZD
Sr76/NMquDKfExx7wA9V9h22rSW4LlldffbRIxpOaCVnexrgvurwcMpavtmTL4/lmKsPZvrmSl8p
9GFIGMcUQFjkPQ+ouGmbiN7qanL2dW5t6RqSL5+1sRMEjrumULNbT/hBwK9qa8Gsg6oVVtWLQB2l
1jDEcMLWfOs9S7rv5caKbthwVo0odmM+3dkg7j8DOx28NtQidMZc4Va++TBbnRcB0f52YeBEMps3
MIUFSJA4hYBHB8XWW0H7/32t4kdwnaCpAtFLNX8VYDSK1MH9hu4ZyU9AzrRWZwagw3K99b+imiwa
qPcgGuXsnJK9wlKpwWqGxIKN6tFYiDzHVAOM16JgUMFiArI9i8fm2VKK/AK7bJVxk8gat5Ycg8cU
Uru+XHL56d/zz514+Yo4Ff4+12cCd8CK013WfJObMEcqd02MhYNzlwgm7u3clhdMHczYgkBJH/Eo
Z0HMNoSHRIFvhS83QVdyyyjz6+sagdbjej7x377l6tFdMBKa5NhCo+yh+FABNd0PPu+qnDU3eJKr
6+fKnws7vtnGCtTr/exee+CBzppouSwjBpVbnPg9aA1BHemEw/BQ8LW0sMdOBSReAEiABAJ8dKnM
IMK9wUlJi5K44/FQBqapPcEmnaRyS8MZgv13/Te4kXKHU2LO42uIUQaBiywJmkM/fnf4EO4SNWCS
/ZPHMSsFpXMZKHD1KuCG9BcETIA+CQvCmdmMrtiVYKpTy+D38t2j2AaoNVa9NqDyxVAvVIO9V2qi
LmJai1LC/2oNiDI2jdaj0Jhe9v//7NXxNxfOvyGVl3Gj4nsmzXeR3ZlSo8Q9UNYUZ8IUPeSNYe4L
WM7WHgJTQ13E0/XpUQH9/B3rvV1KFR+6JLpUDOKK4lWuFbDR5hNmrjLJe1sTE7AbHpxob8lRmCPI
K9LUexAuz3WwkYtHgqFxQ4yKqIGU3Y8jGgDDCuxuffByEk5uA5VZvnm6HzMXz8BeUjhE0/P81OdR
7gJGzECZ2xOUxcmP+seGvNTwQC7PqlPN4J60g2JekgYZoZhG4qciAdnrEa1ppf301E8CrKqu2WG4
/FbxExmyl+DDj9WJn4wuLuk0NJcl4l+OU4TvphJSNr2ddSIVdqt32h/ALw6t5hfgQZ9i2u9C7fWv
SQ8CECDr0Iu+oKXlbkIHLyYBLP0yiGcUhPG6+7rZj+W1clwimhqQ7NwAQmoeJYO+isOtvSvJm1J4
omYxVMv5+LjWVXfDap+juLPJTF6LDj8RPivlW9P1Vhkm9Y3m75n0Ka0C7JkICJ08MfK1LgE3FKEk
FOWy4cTF78D9eeQspqasxAU9oA35SXV+TCNo3k3TOcG8UzVDB9vxy+YTuOeET9Qqr8WDVtr6Of8R
WC4wmF5ks06rCDorLYlKBUoKgXM8uSbfUluXB1IeyukVhs2gRbuliOuBWVwsJ7gPbnUNnWjCRaoc
HS2q2fjg5eH0Dc9InOE/HPPJJI4Pera2e8Q7IYFntQoE7fXvpVGsEHKEUdasNkU6QTLgI1Nc37OS
ppBju32X3xv55HHl3ODEElkSFLkkyAJb03rLzTHx0/eqYpg6k0+nt1XPMqqsIQ9CFafBFjKYUMuW
YNo2a0Mu0Qk7++++IIxHpDVEbZLzm8nIiynPcvSRi6tTzucRQsPJbh2VkY/HSd5W55qwyBtpOQ83
fX/tJsRmie133r9a+TNCCB5Tc5gnjY4j1VtEE6AAfZnIP9nf2+Z0ZwAK/LzNnsF3Iz9+61lpo/6u
6Le7uCrtx+HVQ1nr+mxkm9Ezdbo/ZS0i2aKMz0gq1h0zZlQ+BvKEkh4ggarQkS07uHzt4C1IWAot
D578ucZypxgQBMsSnD7JhgWBZsIT+aSzFTdxD4lZ9RCFOdKhFXT8Q5t0+h5VdRQZvFHE+y/oiDKx
9BJitLuwkKgf/mBlw7DZmHMSpuUxz27j1815ae44WalPLLRIkQffginqdQEJIJVLSEv3a6qErrLY
GWgnDJaTYVkpR70KMeYV1GTG/Sd1ELjOUyEuDh5XKHJ03LC0tOmi/evs2zwBMd8WnfxI7gAP5rG1
7Eb9aV06+P5aFETGpbdiIFJYDZn9cbVaSCb3/ixfb/dg2Xdb9mOdkZEU3jKCXFjsH5Dyy88Fckco
yCwGeiE0jRLnB7IZT7X+9bp5IK9euZrBX1QYRfvjJrWr44jYiGB7WJqDqMof/6301fG2/wOy1iEm
8tAcp0fiNEvNJaqaIBveLqyzm1vqwnbSDCX1TLHLhIKy2NP8DLJr1T5ERwDrfk6rCrngaghFGNed
KSyv1JLHZaWbm1UZlahAtWhKXWqL+xGs66r5wO85rh2MMJp+i5+m9ccuFlYcbM8Dwuz+PzkJQTAz
/ynGc5U4/4g3G3dOTU8VYYrqosVh219K7gM60hTiTHbv7uwMIFHr9/AlIjokxPwatiEJYIbRsEyd
4gBcQb9UI6gcAhwC/Ai+Exk03OYWVmze059av4MQasvOx+8Dzv4JZDnb/mbGlyrquykyqpfEMyU3
Yz2Ddo1d4jbIEHpDNIuThTkVi/q7ydn1R+pyg5e0FsLIJsfZzufl8Iclx2AH94B/x3FxuMmvBmS2
xG7Rem8nQyK/u6wWfna3MH8J162D/EBhWlfksRR7XFJVbwjbTW/BV4rj1F2StU3w1khorPeYj8PH
Fukv5bJzovHOv49d/KxhKvThttHbCMEoKDW/AccMcvqOHg2WQ1tiDw+bstnxoYXInkK+hdrVhrsK
ywkGc+Pelg8Xhv59SVZUdLNaPCjR1z4lTzUVc9lrv/lJIGLutS0vH8i1uHIE07s8wdALlGTnrLG6
sFWnUMf4nUIMH1A0AXBzxgINspH/wKYsTxLSHpYRvrX2P1BIfV6Z7q7SN8Lu9Hsyz7AoNnQAGP77
FpAKaxRgtktOP5Gb8ANC9DQeFV9zaF1zgIxyCNqzFwasL3Nr3OT9RYiSZ18zgxFeJq/cShQIGXZN
dnbgVoO9toj+Pd2alGtwOwmZmuo4RUkGTkT0qkQ6dIFK9yrLRga6nUs78mHWaQK5jXNiWLoqQAPZ
7t/YFmhWOxbtEFRWLm7U6Si66evXLyQGaAo+OI34NLZu2/hBcBr7mhGTMmZyPGrRf5RKIsnmWm3h
B1PbTjepXIV/SmwTyf6/I0pVN5Xyp/YbvhojKnxAcE6BZtgRhAKyqvF19dqnHAl0LSmhMg6coYAM
+6nl36ActE6PvlSeEhHdODMVBoIuNtYI4xLPalwU7HeBwHRRQzGb61UhD25UTG49IY02NjS9lQVy
1UwTSly8T34vbX0v8glQdGOy1u3o6F6FOpH6BA/3L+E8pT+mXuXtI5FYnk5xXdqrJvJ2CJotxrMB
opqyHpPRL9kNtvVF/MvQ2cK3xfT8rbsaDj3Gjwph5D3T1J6XBTzvr+pDQJU003TYtEhvfhK80Apj
wgXDDH8kztJzw5MziCSwy0Slv8ZWX3rwrCx9wHxG7p2ODWtoybDTCNPnvcijC5jiwpnpAkWL7KGq
UdnpLycR5z/zZxz9YVYvWlTDrtr6xnkKBPIz79/J/wZERxJpLc23jNkqCmol9LngB9GdtNCEQ2X0
DCVEsHPYAT4IA2KCVtP+TlVxJAgvGt+Y7gMgXzqCj2pgYhrQvMBQUByiNnVcfC71X8BNJRKG4srC
k2WmridKIvJQCU8FTBfs9n0S+QLSOKrMf4d436BzbzLryOWJSjLr+8w7Z9//MUoVyBPXH3QVgI8r
+SYEY8wwM3HGafoU9ynrJtWAOm8nQoq3AmZnhbcVLAZcN/r0R7BdNWfeHR8DOMUfxfBxyHC5weK/
h6CnVkwCwicCZmMmsXvkbv7OBw9yJakd0bPD/1NjXaiNoAyt+AQ1HetrqGuEx+ocQrZ3gRjYFdYZ
kV+ISBuXHeDItTvTfn3yV5VkZxOAICljWLzC2knK6rGnOWG0mzKmZsFwsniiaNgPa9m/y1SwVMnE
/gP2A2dbsssjt/Ssjj1I72DKAi+wbF4K+X55GhOFh1uAuQpfI0chcmu1GWBeIckAm//mctrF3eVU
FIAgxTC254m5xrjhmqRRqcVMTVUbDQYi/OjA3qhyakndwPaOSH0+0bOnInTBQIl5DMYBV5rCEFaW
Qff4uu9j7Vj7ka0G4nopmEmfXKnAuzf38KH7sj1O9pfY9sRKhTj6tuEhs/g/wC8bE1Urk1utcEcH
xM9zHJzXggYFjyInHWSH29WqRMxO4hFSvP7psCtUuR1kTLMUzNQgBDONadNKSda5irawgejG0nPn
eGjB49sP+2MZrcMR1ni3JnGBz19reecUHFLrVQ7KsjjWONFSEM6thD9CY8COltNvdkrrBcDpjJsF
G376pp+RMZTMEWSPb4eXPhd53JHG5tsrzeXtMvbYPT5WAFGjMP5qMDXKz2+6r1qyNlPZ387QQRiJ
8CbNMFRPBLQKnE/0gokiKRpu1RXD6eza+y5MoOE0+LkqufdcikpA0c3OflGMJwZAd94kmyhql4kG
YLbf9g3ZTChwcmBap3OIijPlB9tf0opLCYrQMdUMs4TYDFKLs65kvRNAcxXfiBRXp28nEHyH7BaP
fhKW/2QsxTRkR4qqCYGN16igd3hw6FrnCul2/W3ZhwCxdv63780dVGblynb9noA+N5gywaaix4RA
t1zyX1vV4Hjf88y60HpVecRB0AKoLctx5AwvRXgjiS82aKC0u1Aroq7rSWVk1pHY86sMlSdi4+tz
TvJHKYJ25ruYO49KLzRINnG/yK7gwqnadQc4juB9pdmNYqdPqJSY95+mGKrWjxdJD7n+aR9+ud3i
jG2Y1G6X+zx4yJgWO+0OIJ1qqHIjHnTlaToVjA54iyaRMzm1hyIO4aYK7X3JlHOCyGiDyz5woGhr
JXlrVK94JHRIbG+W5vnpqpTC/Qh3D+2FGtj6xNsIeJGAtRqWThJBLv5XutJRVtKse6aN9uBNRpYA
NUMPT3QM+OuPTDv6Xh+TqJkc2E9D6uzFDzTw40Xh0EV5sQ/KHKuv9CJtagZCrdMOhtYdBsL5hc4H
ZoP+gMnOzSvULaawzziul2p9cKggXmrEXXekJWNNlIAoSx6nhL/sXVC6JRIj2JTCBvSLULduoscx
tKDgUhB0ORqHksHoHm90H7Nzdnjg2ru9lQKWaVHsOFr2tO3t6M1StvOPMhAYv2Q5r/UqwXsFGdOj
BOFtwZ/Lggj0JCYey25qDOdhTgCVxbtOlXTBc5GgPG7QZnYl0KDFJtRK5M+5xLyqpP5oI/1c+fvd
7TNZM3PJLXXoYNQdCrc1qB4lsu301mQIkwWwLbW0WIZHp7tFJnvsvn9rC8BbIE5fhPt/YFR1uPyj
BW6awvFv0MND0xf/z5sxvvatRzXjU6tupo6LY9v1423JEcYLmlEhdhO1eN+VSVk5esZd83n4Pxff
5dm/WN+Qe8jUdNLCUWtl1vJYEvsDG5pv2CcRRUBGVcEHMrx3XbjHf1TFPKMTpYR5Q113TLX0rp9X
9wJhb08MTBhhfCrvFl2AW1IjCowHRSICp6X+QNm8xjVBExtX1FrBpFW3UrBdh9xlDI/MygahMvTV
e08P9PdxSlWuRKYopmImUMZjf9vWI8jI5/aIbyK7F5BNeAEaEgd7GSKmeDjKcfOz7+kjpdU6Xqhd
Hx6VB0eDoD26SXj4GgoAHQ7dE5hTK9M1pJWrxZOvtty8zbyQdNfnZjY5yLF7EuPjm02nrLNMPaHy
E66eVT+4TrwNxnWp6fk1gF0Z2l+eOfXXDG0JbDtTmGppmwy48xXNeCs3L+lI2C8bhsvM6vnU1M/F
inejj2CArdy0KxBJeQ4Y9DcfWAgtcIYLK9uQfBcgvcEX27aStM8Fue5I7dwmThUhaFS1q205MJG9
jIV2rbrrgOoYn1PkfpBh8Dzy6c6jADJwr84sEn9+9XfDwgjBhDmPnyuq2CkF7Da3Pe/iBoZi14Ca
erBlMnACeZZWp+fgKB0v+4oRaISHaR1Pxob2DtafnUWIdX2ZjOMkxdnSMVTr+sBq8jfWBgTNz5Kk
egJYiolBKSHT1e501L1AueKydB7/USnCs34gU2IiXOP6Em0UoZLEb3fN/1zElh7PIqrNfWr+/oAH
/tUYU1t2PMASJ88JltJaxgE5T8LMc8OkoHdPpuvjLRNZhp7jWb9YEfKu6J7Bs+RUVD9gQpF4yBn7
LkeylPy6SUSDLjUWYav/UePOlBkAV+dNw4CqUGCKY8sPoGG3K8twmTtGjZzKzFzDhASPzFUsAqRt
3zdz1oVTKVa5uia23165lFXYHUwyf+MOCHwpKuX9JFoCSRraiBavjPdtXrolVK4iV+0fAacDqsPB
xURzmyiZqLkTvy36vJ+kwuvhAAarRYEZg+929VC29MSA+9d6lxhnvIdhMh5vRu6PK9+AXhZBQlNH
82rCgHQ0xM7jlzTgaUD5RBKymLNXxzEd/vUbo5TUbGPYFHPmR4U51eBNbT+CWGVgf4a4Jo3jMMKy
pHAqrSzkqeTt83aZhXss3AeQDHbP+NFQ667tyJxTRaJhmKpDnZNnxc5L0v0ch0NGOqfNTMMChbLY
HBxtWdOW1iG6iDiDUooabLqMK5LUrLHR0hF79CxQis8UDJz3BJ1ek0RPmlG4hwl3WMcMD1p07dec
y5jgWFAyiRxP4kin/qCPvkiBvIv/CKCQkPGz0UppVL1d8w+MXfx9yQHJLx1E/D9vflvgD8pea3ql
msmMjmbrxRiDKVaW03+vuvz1D/dt3JVxWZmGVr2E3+6apH3wWkVQLsdbqMYjqJDj7f3yiMqXpCGm
nRGrHOrcxs+OVnLAeeXho+bvzRky+6cpsfeF4eg/OuyLFD7ik6BKyZFQnO4TKaDArUM0yDtANmeF
doCWWsW9rtgaOhgHi/cF1W2P7/W2I3Esz6tiQBAfGq33mlZ9xka57jJgFYC261FW1RGr7z0Hxh5K
Rm3wurkL9qV6TSF51P48xhifPNso0S9MrwFldQEcL9cV8hM6xRol1sgogf981NPhgMRgD4bgABzS
t03P3xbCeTwVkZOOlinbRiQNatrzDIJQhpCQe75ZBL3zXjM/+0Onq9dv3GTMECL2EMro3Aw3l+q9
5Yx9pfQMxUPaB0ptgdem7ht15O32Xz0XJhLNxD3Iaxg3LjVtNezpc3TSejGx90+RynSb29Y4Smyk
yx9guc6JgIPfrh56sNJXQgMm2ZA+fbUcGxj6fiMoSmG1S4eLKNA3gNQSj2To6gX4L/XquuKtMzF0
cxwOlQmmYFOk8+inWTOCjdN2DG319TYG98+T81bdL8NrdBJiReCmHgAShKOtrTsUn82K4HlcFIHd
VgbC3FMHiInH3eIPDfWX1wmnHgd0WRhac4kjgNqadMmiGBgO4/zeZrNekJe+IgpcC/E4amE8Eutt
4vmFJjz+Fp3XJ9RE9IdLuAQQmnfCjuMjTd3Li+mgMYHrHUxPwew73U2Vdywj5sGzXqcPECR2LYCV
DIiVTsYYzsRw5VUPSvqFlJhV6anHGV7hu7O7TChFGGU1Vz1qETQSCyDsvi+uDF9WeHAHBedLQ3Uf
6Yy4SvQw3FpU54fW5FtyymD+dZVQM5n6hewVLe8nyVn02FNgH2Cb38ZnqPndhNDYQJZFYhJ4sTzY
5JXWxciTFjPdz6EcMTM4MQcQt8jzFlgVZz7NiHvDEz13BId02J1Xbmo2h9C2k88scLzdWYnYPfxO
a2Sg1Ghp5gtEGiECD0K+FuBC0rNMXWo05bA5Bah+7jfRNIsfhMdiT3QFUkclRv05REd+TicX3vOm
hmmocX4svGihKrk4nJcu5S+UUYST7HLpOhbQxc6uFEI290BDQ+AYbiTroViw3/lE4sGlOrC04Dgp
IAE6OOAfvBBLUfUM9BVGvZ8L7O7WcXkRaQAFaXBtTicBJCc/YBTXuTxPtr8zHI3s/0kBy9zMdxow
EN5e0kvzRmSVIZJ9MmU0iruaWweH6mkNkiC7FRKTEA8nF20bBLwHdoOX4WkclR24ldq8zbuhtkcd
mLeibTKJVzKaq2hsoLIu0mMf6rBWwjcl2qlr8QHWh7vJFE9Tk4a/skYCRp19TnnRbIVU9DH04WLl
dNUAAEHlVY1yF+HRjPMNzRPrBipJzlbN0keg6VCbAwsnn8COBwPrO0BRK+jwBFdMWHqC/kO16ZKw
GmJbYUlgS101EXkaPgILjeAF8C5a1t02qAt+aYK+FyBPlWcAizRwopiwMLbl4jP4WlRi288AnSI4
bSJFUvvE501nMk6VQc2a4MtCkA6rokkSb0M1dZshwg2wxQ0+iwgem4yqc3OPjOGdMBWTSO/5ecQX
Y+z69ea+kY20rZnB25PQtZfPG+jZRFGcRlYPKn5WlyiQgJbHTIh5PcnV9hjvPe3PGqbcrR0785lC
/IsOgiHvgMFQzKKONhX5SXHVuqkSp0RPF8NcAfkUeyaTKergal2O/najDJj5dGTMuygbszike2Sv
1kwJBoHMJEUMkICZh39yMoizAsFs3adI0Fn722Vrmg7RplL8xdE5yU6M8lzz2blmj2xCilt+IBNO
SsT2BO6l4ufjzugWRqjnWacYsbm6BcJ2i0COdDFt1YFRrJ+M6ZDuliNuI5u9OvAJYk94AD6jl7oc
IFoPKH2RlFUGz9xuhnBnFW3VUNAH5Q+QukUXcySVJ9R2pOnyhgFnXqvMYXkHMAt/hvPuxo4KvFVh
tUhb0p3DBJ2Vm8B+w1oo+YURG5Jy+2xS5Wuj05vJOnDjQZIihhFuM7plCVgIlOpb+ig9pKyCJgll
7pbZt3kENv4evMBr8VSXq6Cw7VqtSxy4f6pTcsqaGkoq15HDTVQTZL6YP7YoO5Pw393CyPr1vUbo
LAbYLWva16iiwkWdHaQNx7ILnW3RFnOqTvYcqZzxE29aeIT2gOng/SQZgj600GrrZ3yiUIzvWe2b
X8HWJS2LBRw4jRIJo2Dl8XVWz63kGqdevStSbjWEGY9bjDEMKoonaaC7jLFtsDu8piGdxAb+Snx1
aP34sljcd60RXoY82MUiAu/lYqm9Us1XsUU+t9oJ2D1le9r9KO6EBfLyjw+0A8lyEZFokvgQbhzT
fXWPcAe766YFPtLEQst++ulUiSOnmbGoTfdLCv8ju6vJuqO+on72ghpY7W4MNSewKxb3Q78EarOw
96m++gDpGHsZp4InaKrhIzzumDSGNT912ECThvEvdPZLBNuYh5ADOniW0pbfLfv9V0kW37lggcNT
a5D+1n8mYbnV7m0LvVGwPSkp5XcIzz7Ujz7MoqHARukZATcbWuAgEBCI67LGPnJzg8z3GedDgEfF
TxkdGKDr6QxTxXMpzrk59237R8Zo3fvtTSNmneUCEcpEWSIp0BAwWDjzTvM+cB66lWp06Z22lZfU
jvFrLc2n2CHyCvdGVkt99MjL7z6APNMkC89opX5bEt6WPF05sP250yeiyAgOraoUehp5UKJZ5kWo
fQwR+nEhI1ZX+rHBqQVcSB70UlKQSe5H8l0ZGYDFFk4sZT3y2ji84W86Xn5y7Y06ztLgk3T4AvQn
TjGpTZWwlTcnvm3Hii+qrWqDErXMi9Z8mhLZR+2xVaoZVJtqReXM1exQQocwLSgKL6AfYNJKG3Eo
IR3IYbbrL9pnCkAQN4oo+lv23QTd3BZAeaVBP7xBSSHlH/qOChy00VxCX96GEdpCm3GIOOLRXx4k
KYud1QYsMs1Zyu0zqUsO8YU10TFVYZ6/doXjUIjDayL29iSKU8qNr9IktBjnD7CRJ3mwYMesccbb
zi2vM+U9VlSp5lZV9Ub/QesjdzAUDyPZ4ohJyrrZei6Y11x7z7EbPsfMordzmmN6kVa+pvUom6UT
WuUpUr9PmMGxXq83sScIMH6Do/iPApjZOqzjcdLv0T1iU+0r7UJl4o0T4Xm3yBd9Ey/L3FgzTkjp
8N13cDPj+JcK2zrHUzDDfyzjHDruCOHZ9jJSV1xHxxzq2v4lTMJXhLp2pPwu5VEJ91kndtsUoBMO
KttTBmbuq/9q7BUSHpFdoMvqkniLJAfU5cUq8C00ywqIdbFI198g7zQ4BhN7FNqsQI1xqWwh4oq0
uKTBt1m5UZLJHK+foeE3o3qoj8+2ThGwOyfTP96Dv2vfuQoF8V9Pp5kIeBBj4MK5QNrxfCDyjQZq
KHWrLEoCNGtKT1Cefmgjh4QSTRpBtRG1rJMHe0/2AxAlSnNH5SXvVfzE7VT+h5KgjKMq8ueqftP8
klIXOgo7S8/aFp/MduMui4jPHEDkB3Vyp4rAhVgeMLVvoH3H3msCjBL2umRHNe38n5J7nj4WR/l3
q+5p52SoaZ9FGNGrmGN59/9W/kYhAaBiXQGxKbV7q4YgzEPLZkN1r+oXyb/yqCGjHRABWgAmGNv3
Sp4QWxcbMo8aI6VQEz31SEiQG9M6yph6DBzhKCF3RSchu5uQX0thusvowwKJ3QOGqWjxB2LgoKaz
yUV96hTq2Gbe0ZWB/svuU4KFpvQOYcS/j+j40vO7R6wmezGqwuxCkwJ8/JcPqXSQIMWASWjbCxKx
jYEeQ5qie65rTMtjCQ6Q+HUrCALuZG7SJ2uekIA8zxCsedUE33L+3hlg9S/I4BBcdURkbOheoxPk
47tA4RklrJaJSv37zeDy94alG3TnP5CVKChtgKzEYhyeB3WP3oyY6t84kKtZ8vF29SsVYB5l5q8b
8URTekOdEeSh1xAHOf17WH2RYa5CXwHIEqW6Jz6AKzvrjcqjt8c6ft+zU+tib/ymAOoEUMx1cJQE
HA0cPjflO5RDYheGVc5WaTyFSlNNh7XukQOJghNqvHd8C1DISN8mBcx3cX8oErCUSe58CpgyR5Nz
4NH1B/R+BRA0LzQCIjLEn0329fuLZAC+vp+B48Jby7ASEo92IA8eP3qi4/N9TMPXDgRx/kVKoYt+
bKk4r5nTRk48NpoXIqqUH7Bn+QjrZQHHWeMLaXdCqbS9sDglHtdDRqcqJ/Xv0vgtr9qd20Yg8kyW
o29OulRE2nP8VoySzYswrE/OudCh3zsyD0fHVAAoMWtl5l7oMip1g6pLeI9gbyBG+ypoaVJK5GUO
L3Sy2er7kOkoESsvTINhJYPrwt6oxCydbAj2FGa6+Inn3vBT4p3i1L8VdxDCPBOWfiTu4Z21l5CS
g18ksCHD136/5Ee5zTAot6fsVEvgdSkJMj5b00qtGSd4A9s/B9abYKk67aFDEDnzsY8NfPh4n695
VcTvLJp73ViUupJlNzZwKnWwt4miTCfCEZEmIgwS12naA7wlAMtUL5wPVdhxuxNChDMP+PIHVpk/
AU16aHoGLPCyqdure2lSn1b5G6tMlxIvd6fY81oB4WHvUGQf/+x3q47pFXND9455Gs3uDkChIWqt
JbHds0R8KfSN+j1Q+/ls6XkDSjS5B3ky6B4d8qUf9ebvD8EbHB3gPMeDuIUpozeEYJNdK2gmOg1a
PRVlWEOrBYNlVeIOYoz719DE4MkvI/4L8qOh8aUeMX7AYcAyvSyNu3wHUTKuUR5idYmYxbaxS8S0
/Urh6DiI0lrYCm7u03QzwIP5xLGjm5nBWsE9enjm/IDV3uJ5y6wZOxtVDNuwYELe0vHhiB52vP1u
35nSmLkRCiafDC5IEg0lfRcq4LY5gqB7j7VC12l3vtUr7b3WRV3PFGex9DQ1RY2xJ3NDOHEbvK4G
FfNOBwec8NwFO/80kOTgbtT6piYDf1NwTyaShlXyuxv7JPeooZgBKfN3r0t9AYe4seF1EeYwPwGC
HezeLXoIpmPDUPKmtqHlmZSFUFMJO7raFCPIFtXz5X27TFHaqmKNB29WkBh8wIH7edn1gWxxXW/B
jURo1bzBd1mHRqIJBuYJBiVA6hf5aGnCFXh9e02iKAegUv5759yUKifhBa2LIyGNWMxzpvtqVjfb
l4KQf4uB0qOqYE+4AOiohhzAOn8f6CWZ0PAg1+J1eOwOXbpwlxQnQIJYJQOwYlZ0E4OsNiUvaxFp
SNf5U+AC/DMvfHp2F7ec/mJ6BVdaBmu+cYLW/X9iCgjeefvgCyiWSrW9x1Ap3OFlJ3iwINjaRXLu
3H2o2Q3CYny1n77+jQXirL82U4te/G/myd2Isrfp6lhBr8biUsG3XHdDGyccUdI8k+Kq+ae0DOEq
kKBef7AfHXdRrH07hP0+h72fPAPQUYoJ6DcBNwRUDl55Nm7X5SObEXW3xJw6+a+9eHEBiZH7glft
UwgIMOqxpMr/bbt187k9qSTQEGEVrCajTxJqLSIQXGHxhY3y76zVi4wd9pdUb8JyJkW90CmqiQ3A
+HlVgRei08KRJlRjw/Q8K0nApMZWzX8elvkuT0P5BlJZHSacC5ljfdPZAbZvymrsZ/54YpA3hPvK
qaXRTLWx52jvZ06JF3q2n9PsceFN4TdGQlDwY/4IGlw/ArtbiBKrk3SOSzCPOVxxvVB0vCFEsO5s
q3OLlxi3BvfeUZ6OqSM/PyQxEYIjsuTmOuXP6A0XmWOEc5v/mIjZv25fH+vLaxwLpNvolqlsVgPX
vm95Qq0iuiZmsBppjeItj1/JaNmj3SpZAR+QQWx0thW2Oj8Jhn1+L4JeeHwQNqmgV9q+TOOkoSQ7
+Ys7C7H+GHsUECxe/YUFeCgGYHvbmU2D4P1ughMV3hhTof/NoBjqG55FhsLxL0y/xUalMFftsm0w
g3OTgpyditeJWw9KG3Eutosk9daJc/lG0ZcKnZsO2rp/Vu06lkSweHQjsILaI1vLZXpTJXx63adm
b54wsTyKyVsZc9R3CJ4S5xVQ1R4llj774PalHQsu0kcHu5ZoI801D0X2Zeo6C3u6EMv0EaJJuEHo
MDFNjEH6pWrsJDbslU4zp+X3do3WHfFYWGoiOc9k5OsKlXG045PXKPCQxX6t//sZMlyHTd2FXzto
ZFjvhdSBeeW8T1kaRX/XQwLlsUCicBA4nSjzGye3bn2XOqt5clyKRqIu+YJQ788sniY4tJ7R11i1
gg5Ly6dh024BwvjflgwPjH5kT0T4/KXESdkYF+hcFyQOSIIwnJEAfVCd6xPMOLsUPizgQAJaRGXA
jBmGAIq82RIOWle1RQgCa71tcerDIMbwB5aXgjTah3fVlhxPIE7kd1sG//SOZi2PEJyzO7CJsIjg
VJ5/Qr+VQ06z2LBN/LMjjUUbo8zVb0x5bDUlcGUzVI0hUx8HeL7RxgvZZFuetmCDKMVKBxIHZ/B/
OVWQ1YZLYiIl2fpcokxDeiNG235movj5uCKeEUVWa8EqDCyWw61kg7E3zJOVbMTTz4YbzoOwEAmZ
tHYdGzo8xMvWgnOBst2RttqWI8cGkQQbTohqo9Vt+ytLFhfJ8U5s5/4fU1UYq7/3Dqng9/MkIgyj
Cv/pnIp6S0lVh0Im7KgtHpREkTV5T+yfF1EGwDkEraY6x6fupAcNrRCOk4XJ/lXfi0UJlKVediMN
HyhH5WUdciewURKuAxhvl7k3LwumLn4EviW1IRqwHeFeyB9YVUD3CVAtOfpgQbs7NS1Zt+I1lVH2
XTfTDrIMQrktsk462d7WU1YciyCozVKnGqOLiaArmQF2JG+oFg2FlHKJbdhXeVSr9OYSx/6S5SBC
XWertg7QnFKrCQbNFJEepHdb67qtEeQ55n12UT9CkPLfq/osSMUq/jefLJytG7Z7BClbYQi0LpuP
Sp/eKLkZyN7gnrm+kVj+U5iCSP+gA6dYVLs66ToDi9o3jkwBIkFc0klqyocm78Zb9BoQntq3irai
DFWRh4itu4nIXK5mL+JNlY1240/FYxsUOg2UtDHXSp7lyTD8xC94GvvHaYPYHnTMSjHruOBHci0c
GvIrGh+eiTzXdMsn55PN0IlzpvMp6Hy28n4ofQxVGa7lrlMhUJ1HX85CuyVajDjBHCoszYWcSFov
RjbO0EPt6CmzME02oWh8oiF209Jb1n7/gfZuH5Tp1OrfYKPIUKAG6WaMVigMqxpq/O7R4wm7/9G8
jpBjOn3hKlsEY/f95kNpLl5C+wce3E3g4e3gsAa8ciAJZpkGlR/Cn5HatnVfszAPn84PvCf856EP
yBpmun0AqCkAf6LDoxP+9n+aXAi4m1m5Xhp1Dp8SGCiv+Gk566wCLWfQuZ82ELCyXaakzt8TN9Zs
TAzcAprdwIHVFi2+KU3HwpIxJAqcFD+lkCxcv+KxW6ZXuh9mqdcm1Qy6goIqCuJCiQIlaPCkW3Fl
n42rVjq1/hkuEMCREOOGjjMMeWTy2t0z7Le0v2u8kM0RyRBB54zQ4QNoXwafUKKx6zNT/F4fsJEz
Pn30I6FEIMWb3DCTHE/MDCqUck82aRgUoJ8gspLEHHJDoS5s2R/xzAqnquMCzdXsgBEFEhRRTo2n
WvH0PUui4IOG33Qi6eXKy5mMQLlEHDjWJtWLRrQToJzPD34ODEXvwrPlwKc+tfta8sOnvaGlzBpb
0se7CLNXDDkLbZ/CgRXLhJFG7GRd4g3fg/S3/qrkgHOPH+kOwtcrjzx7mkm9PHzwjWXffu6Xu2ja
/mGfSgCHS5Tt7vtvfpKMi0zjkKeNg/OVSEHgsAs3GhccCahKBpD/hn9moJXNj5k2gXT9Cktcwrig
TBkCUn1LTOWD9ZPo/bJdEvUMPyWyKSK9HLuwOjzEYNN3o38jo8dCOBm1i1rOYOcEQ6zTKRFA3bUt
ZvLI8HTMiyqbQW1ZCVJI7D4vhZCD9VLfyv/RF6DwjgSMNXkr/sf65bQDHpRt/QUX7lIzzQG8k6S+
j9WQkKo1gbqLmRUfxgBKW8Gkq+LwJoS4JBlxIkc0FjI6g3kIa+RGBR/c0AKbgXSb6c4T8d4nUVlm
DW7kssnKljsW+EzQc5PZ7bKluok0S7Dp7rjwPfdti6tV2dQTYriyh/tVC+Cx0L2J4jh5/t2FdUWh
AYtB12/wpYhPHD8mkuI93XbXzgpL5727/nyZsdqmyrSgMqaKa2WBSNPMIwYmPlykhBctKHrTWq0e
NI2YeHQKpeUGyQjSk2/tUPvJWBGySZl+sBrrSGLsgsuLbtdCZ4VcaizyTU5c2MRlxSyJvkoLECr+
LFNwOg84F1iZfofceeXKPOp5qiOdl+TsBQwexAul0tQ6lHghLCA/RU3nxTMhx0xgGmx4DRl45tNs
TjQh66BuZsu+BcpIyL41ys6MVrwg0GeABeAsLPuGN8GHIja9f03wCibVw5eSMlg0+pMFg8NyWNK4
KaeKlKYnUE+z96ALD5PgUkWYMblR7IM8qIsuVe1DqqNqF98BV0+XjfE2V/Up6U8lDsb4DLrzdJTO
P0fVsXeHe+2y8dhCC2IkM8W8wAM8O8vAiMponuvCo1N6mpJ4h2g9GhYu48dp/ErEfYvNrSR46f5L
wEOjk6/lSs/N9sMvWUJSj7lsWK5emafgZJbKyn+jmAIARWTL74wUxVp6yNJQBumn/hMNM/pwni6S
RaEmGv1Mc+DsFLKOgOvP+QfsHuyQOvGWbM+0hGFhW7otOjQqV+/Jst4uTTlPdekrKcFp4icg+Pef
pKnE1WEk8+ufCQsJd0HXIx+cslohtTvpKh9qD77BjDPpZTTR6GpOLdhamb1sr+ZBCSK98XF+mkEc
jOQNZZEyWgLvoL6NscQes7SeeeV5NlYRGq86WmfGyNb0BgStyx9ccUlQy2YVROqQq2XH06Z/9IWA
UmQ/QrhDLMLVxTRN51V2WLwMWVoENze9gcb7BRoJ3p55YogGsVPukRRHzixvkXXULTUvhMTFP1yR
cOok8/1JftcPG93PcqKJP6m5xKRJRWTORohRhv6cJla8uJXz7zZbWxRm3xXlU7++tkleL9olS2lz
oX1QmMxNlQztkpn1cICZF0abNFchz4iXtjOJZUgI9aQnroCWlWcGDNlAmRE54ahPp/vm4Kfbv52T
vXZZAdP89MUYxBWF2fTgb5ekBO88fzpzyDmpFbHpnqMMN0Pt3QTHzpA8AqOHIM53fBf79gr7VCEW
qaqfV4ZJmkQFcNIg/Mwbt0V3rxB88bU8NesHVv9ElUTk+zYe7hsV2gTXkIENoPGVJJy8pnPUjKOj
RT2g9tzIaQikeX3q3jMfsjH9V07h9fc15CSqk8JPkxgrE3264SE6MKr1Pbok7+7eqJzlnLbcYPX7
BicM+a+8Y6RUeZlYWINzFUXzfEE0iToOEoOkkDSWHB8RvWreDEa87bQCvTwHTqLowcyfv00YhshG
DJCkYKfv7R7REmQMktszX6QTsmQLj1dCIUB06xYnLlcSlrqp0wa266KRbMfuySXo2+Xv8ctzupwE
Mn5X+4Mqn3W2hvw+f2QNsyDGO0uXMjGnrgYgxqwtLexjcmw0N3PAlcVa59P2AtFEV2oqU6n6YwRk
0S81aouUqk/ejE8088QCbFnrR4P5wTY8wmF/Goq9wBpz6Wz95cm3ZNEvkJ5fg4s9COF7RvuxOpRQ
T24M0+SdBd/8OPUHFK0vr9YoDtEyTxm5o2KH6dWxj2FgeN2cACYPtSpATeTlg6N5T5hItBeJZkrg
aV0tJ2kcTsU0XfbgIsVskO4P/TIFN/odm5ZqeFLTyEQm398Fu5hiwmSR43QHVr3lS2gsEuEOp294
HyYfzOUuoperriZz7iREwp6jtNJyTIjOW2EgpZrBtTziLpe7WEQ805fCL2l4Cp3fJofSq8vvyhP+
Fm783HjAEpe2K0bu1fDRi+bIol1eUVu2dSUWQ6ne5DupREabGwM83jgvolecCXFasp8rzLzjI4FD
y4cZLOBB0ULge/wF1z5j8xX/SJXGKuloO7l09NrV0JDiXF6zp8BpN38h/pTERWQyK2dwJLB5BjNM
Up7YVEQuNqPivXT6skzfNS4GC6KNU4LuXH7r4i06UBywvzw/n2u50N9eezTK41h4fiLcziWDv/hn
YoNYCytwRATtoz3dgAXI4gg5W+Fh0dQLgqyVy5YRklRK5lWnUdfh2cmonQCLpOiZAZPiflSD5LEn
QQc+z/AyhTVJ6dAEc2FCYNGLaA0Aoks5i7Pi7K9GOLu5F/GBpoJvQKTeimuOPyI9FnYCbIvl+BpA
78XGsxcqKDwC7FMRQjfZ2Msek1ehfwx6DoJnhzsFmnBWbuusVjS4/CQ6DLN4ubsl+XL7bP9B8Yvs
b7Gs4OlL4uBAjxN/4n3h0pgKseUW5R3E2CUQ3vVjBH7NmdJ/4NTiOhOFbyKnCmZWNIOcQxzCn0y4
64pZyC4lNmMJ3kuwOaypQxh0/amJfFqxQYuE8vvTg/l7XfEyHATPBUUC8xfMGlPVh5O4jd7h7BHw
PQlbeEPIWQeMj4nRYTqT9VIo+WLQL5FjyuJzk2OzHgdkuKPhtof4rd6JeHCgpZmSQQtss8WCx11w
mTWH43pYOzHQHZhvFGSmqn+NybKS2kBG9qnPkZaZfkQJrWWhdWoGaRLQI7DX4tzCZCvQ9GozQBdX
jN5mb6djhvVoEVCiZ2MssFg7S1nU6YGnSRPM4qvaPQvLrYWcFY97HWAg/xZIGwOO4n2JIgsiKPof
mvXZzpV7JfUY64XBbhaMOSNQ9xlgWIpTECes0gLYyjBrbz0xgRtFJ1h91lQNzssjGJg8egDqixeY
LnL8J4zCiDjajKtpQNlsS5Gz+z8YYPHYaiGMAc6QRf5e4Mw+suqAYidB0mZ5uaUiV116h6Tu3doF
qsrdND6jZUW/Iu50/2H53we9Xxkk/o6o9HEQOHDa4AbPMXMEUFP2s3mqvzrFyMUPO+er56IUG9kg
A+OnvAgZ0QbVw30CvEhTHxOD+sVeKigqS2j7VPkmcPuUuhXBQLLmNCHbuMyQizpiuXpJ3qNdPhPG
XVzhdych32HgUj05hZ8cOAlXAUNpKLW9voWs0RmN5XUNCIXze58xKK4bOh8IxulqBQpxhIQoeTUw
xbkzeTs320wzKeAqZKZ3+EFGUfpxluNpa1lev7Vq7DAdp1b9DH0vw5xhMtTyP7JkIVDQwoSnHOWn
piDQZxZbYV9Edwk8PgBu3rFng4vho5dnEdkHAbm3j4xnV3gNCDbZSeOwRbYMfMvR1EOjRWCP4NQQ
1GWA/yyCe8Eq3KxehP3tdouZ+iSQtlnF/JOLTIKkc0R7QHUlvegcObu7EAAnNccAe2abriM9vHfL
OEax4wknjeZnpoVhnmY6MKubmPbVGgLmtuulDUOCrszUaHcUP//3vAJYatHccT7K4kG9adaqkbPT
P0oWUGYnHyFT9o9WDb2NrC0VhchbP2EmEsPEoKB2MW6aV2BX++GcyvSHdL59YxQQ9/unB8JGJ6sb
rqTMrl1tSKzgqBQz/HfBi/M3R12cFQHY9o8ryVtiQurP2k6uYjY3vIwL4NpkKNVxbnBaX1pMafmS
IB29QZ6YN2yxF8XqwbdRvF6TPcM2OUTkk/wZUJrJG+zl2pRW4togD3gmEROu2HL7iCIWUDjbvDPp
vhOQ/lPCHhdEr5hEFcblzJW+s8mJ18RFjTTtlr0uahAFXzHurpCtBQO1Gc3erev6xiI9q6Hc95io
wHtcvKEmJiRMCpsbkUUkRKF8IpQBKzxLcfqCzCiGmAqUXk7/a2xy4Cv3PASWNbAERKcFiIh5ggoe
OsLDtBn0lj28QJXZEa+pn7aTdRK4ey30epqxdihHpMXrXzb3TGiwtE1wXPKYesAFVqNYAX1y3mZq
P+JHNj4usWj6aoXDXGDHVsmXoWf+HzZBOvX5wBTuJU1+mmglFY6DofnXZWUNvdNgGV5CDSu45Dyp
0w4xRPRBhumoynfpqmXdIBM+Ae/XSh8r07tBiLCb81NNZ2xcQS90qUUWyRuN4B/vwDkfL/5SSx76
IDHNWmvnxObU+0szz6zl+Yl13vJK3/IcR52fCmFpk2TXou8jwP/3Np+sI/1chAWzuOatogWotMur
vevyNT0ztT27BQgSj/2XJZ+3SPDsxmBdQEoWigUa8f/if02K7+6p9wgRpnqGFdYNOfT125G9QlvI
nqarVAPmamtPZoaVymH+5VL1FaizJhY8/NBLBwlLfYgeqGEUuXNwlxP2qg6deQwsZQRPXceTJCpM
wWLN3EgA9Oz01BwObHsG2/Gu3Zy/CZ6tn9S65Ki0Qtj23mmr1/1zJncwtCEmmwtKHnqnoRUbb5wg
9khiJorUgcbVJj76Xs7vW0Ezgyiwsm8JBoZ8vt6NgrQL0Ki+8PCCneFAU8PG6cgqD4QmNgRfvjOj
FNgWckQGgD0yByPssEouh9qqSKeKHi1FPMQcSWdDcCOYja+onMoyWsYU6OTSUx5YkBA/0LQOSoyV
Umpde10/N8EA7dEwLo1RXpzatdRxMMMZ97y4FholREg848EjqygRCLbvxbzeI7J8IPyPtb2txoiW
eimFhR5ymkHIC5V46tvpVWjhfx9b7kbP78rB9WoT6FzA0iIiMSEDAH9u7hesz9CrMFGx7GNQlNyJ
m3ZPBajyvC1As+T0y7g0NbXroKbMKehzZ3KuMcXxFnFRMUfFLpEqRRSSBBTnIh4wty8ZiepNrvwU
d8uceXDoW0cJxQtuw2rpQK1vlZA+KjMgvMvGROnKAU2hJzQf1kyfj23snvKWNTNyRxqpTvdcV+kl
JhFT2K1Kb/y5OrlonrT0y9htg5HPh/knXGqnIjoknmX6h6XbKHh0yJAKTj6XOSNMacSgDMBlyX3D
I8HPYDLvfdhJZwTz2H42JJBTUNN+Zuo6GRPsJFhuyiwvbh3NKql8gwVX8iCSDSmRsbzmXl/SBNls
FkNQ76Ov9rLYHhFPu96+LcNYvjWkjSzlnudz9FW0U4Dr4ZoZkg/aA2N5Oo6KPSygNKZdj3JZRxzI
ccAv7hWdhWrE2V7o1SS94p1HR3McJVHBc03dvAUAkLdEZOyDshnX4O2+67LMMlu/qil/dHDpokXR
uI3D/+zVIXqm8grca6SIHlQWebu3+33XvKiOfZz1plaQhDPOM1a3xzxYlrY+EDXoOP4dEoC6FKO9
UvkIiOpo1UuI8O/QgdhiZYQkTO6yl9SigTVL3eg1QMdALPeWFGN+GghVX35A3BiHyxZFycDnc+XO
W0mu7eboUdKqa8bw4PSSmRW8JHc5htE6kVe4otGTD2sUfIHgXyCQdjLrRSIY/s3RjM/bJ4MfdloL
4OofTDlixcZEua6LiT2FCzL3PIXK3SRTXB73pWNw9gZit4tM+1lSsZMaHaPYNQIYhYQojKfNbPZN
NpVuF8S4JdMzBHAsxS/5STRXgGCezJ/XZzLiKoPoB2olTltkClTDhm40s/5c47tFZSlYd0BsNiUr
Uq3V4pDQ6+QERfv1xO7n7Rs85RofsKO+fvObLriYP4qXf5jrMGcd62sXgsXYMlGY76IUDOEcOZ8f
SRGWKYocrAJKZN62eF24uNOSwHmpiHyRbzdvurAtUSx4xcFd/yyp9hYuVfhdT8xma8D0Is+A5cTr
snecEulARpqI3h1/flii/oWk7hac/N5XpPb7ZKFotPcVZiFei/xxOLtYx2z+0jWkf4wQJnIwA2hi
mA4itSzSUkxKSs/ZhRCgesGAFM09erAdrDyjTCMHIq0sUjKHtuDAmOgMdiYk0JGgU9HVgcPkfcol
qS+GJwHd9YhZzc49ueBHq3E/J7d1c8g64J1j/VdnFEK3MNB0XkKjXUMj60K0kfk0t1H1TSssQek6
Sose3jqSnlgfKOrQxuw2VWZeXTSqFrvNtL2Cjq36dYuo4sbX9B0/lIh4tkw4siF0At1NBo327r5q
KgLcMO1EcgQGNqtWz32z1lsqIWvVgrfII6zi6KTjWBBaJ7priV9wWYzfTx11dSrIH3rRdGA9P+1D
maYwbHXqRK2WP8YbbN5+MGiDt+T+Sno4eF1wTSVi8yY5VZ/+3E2ggNLc/kyk5CV8TLmRkOUI+f5N
P0XscWP9uCyGZxSrYZzLcLAqt8dUUbh0hdv7CWBIZTde8MBklL8DPZnQUwfY7+uRq/Uu9ZA2Y0e6
N+K8cg7z90vgB9qu/GlBHpuaCS+mXtgCCsUPBoLlr7ILl9L3F0ZBeUKx4lwHm0VUNxRSff9mtnY0
0rpyYeWiDpgduGC9DqKQo4alVtliymEQ33OTULvkJ9MRk250qw+5IPH6xznHrZMf6RCEUZbQrdIw
xqWEqBBdf1WbZZv35jSYx/a6M+GDqAEiz+gPeExm/WBBbuR1WglHOqQOJEtpXfLji/8r5gxAXlcr
Expm0Frdx1sPtlhIfh0C0XQvRymedRJ5LxdCSfXBmpRNwDhl028ND+4xF52iY0k2joasE8BihB6v
uOx+zLvxvMU8Ossp686uSrHoPUbscEnnh0PabyhViI/bPljN4+tmH9NBTOH89SW1XY2WfL/hh6yh
lo9vTiDP7z1RVvZBan39drm45Gu3NF/+iMWSpMrUZTGNty6EMyFf3WX2UTzzxLImcV8E53jmGa/I
vj2ZyCiaxJvZHsoLwVteH/jqZg2x0iW36Wz/Vxwb0EdYHABFtR5A9dkv+1yXsW8nIPpk7ogItaEJ
SC9f6WWcSJtBv2/vX3pXmSiiH0AB1PWI55GZsGRdsIuWjzayDSz1tAvkPtmS6RtjtU6QpvXZD4vL
s7X5ScQhxGQDqni/XVvIribbTQbIO3gCPPwSbjjCM5q0gTS8j1RD2gQzjIIjWzxrcTJ0LxwfaPxg
eLiwxcENd8XFhSaul+lS1WG9/rv/Im8vQZflPoyPgw8sRa6HZR6pSzQIc07EBWG/zxSwWS/ycL/9
q6T4eMItQP+kq/6DdeJK4p5V9OM5PQs90iUhFa7jOwYi2YP6NMuT0xliQhM4WTx+8MwsBADsx4Aw
gNT/QXIOypvy6+PfZBrN8a9eVVTMigdpDr5mPYdJKk1PItkU005XN83OQQEEi9Nv49TeVW/xNrH6
LztZ87vPTBSKQTXaj6tmxvuoQ7DRWXA6fy4PPL+ok68gz+OgYhPJGjnRAR3Rq57NZas6pLCM0qyt
A+6LZhz1OWvFuuqCRfyfJwnENR/W7yp0FuNPQzhhGnt1B1cEWESXkGoq4AJFXqI60gNq4SCxamVE
5LeDEoBLNHN4ePcP19CwhzruWC0Vk92RygKafNQxYNg2mwJRkTrh/0eXGeI3Tef2XpAXR5jz9ip5
Wsggh47eTlPBe42XQdePzkhoXTxGxYdsnOd7wq6QZAn6wGe0pO0Xz4QvtfrSBzIdbqArVks1P6s3
xwSj/aPvdTLq5jPvZKq92+6j+L5kefr5S8IBHUuv6obq0DIgt27mTJ1q3wQWNtCHlWbwcFiCQzRB
rfbdc/Ae0oz9Ac/7vUgQF+9HjjqTcSvwRmEFB3Rxdhz2jEE7kjmTh1E8O9nK0Xlh8kd3ZsHuaSy2
kJ2MqolYQqSnaVEAico18fAuRTvabKlqcgDsCGranA0HZFbRVrj5AVmBxq2COh+Go5A4v/807yz8
nLIgYIipiWNx8iPVEq4wGUJu8a8B6L4nNdznNGeo0G8077VsoskKrm2n8+xVP5C33nL2LHUFyrck
KFkssYPQxu65AmEh2lYE5WbGwP0lue8zrxKLKInWJwVxFrCaBnM1AIG9FT52tpLw27dDrdQXrtBv
hBpNkCjIGpOEaXt1doFxqi969CYTUou0lHxxCbN/5GubrztJWIv95fVDEJ88sBGL5wyD1cvsC6QN
gJMDL3X+p2lLKh5V4aMOA5jv7dRap+Sq0m2byAC+JJ7Qq18lV5YckAYSlgIrD1yPGjZ1/FbmJuPt
1c6LoV9VE/Zs6bg/MLgml853mKeJY8UBrofX0o6POtwRck/az/UO9ndTSmquT2vSSFrifvRI67EP
QrjyKb0EKzveQOhI2V2KxiIt+MjLbYRvVbEhzIPzs1prbWg48RPkZfZS22cnJEOk1cljaHxZJCMO
QGhpDEtypXm4Khbmz4P0bR7wkvWzTI/fyuRNzcYSSGwD7b9tufUYAKFV777+CRfkHTJ014mxgKW+
4mqPcYPRgyUqY0Z5LXFHPmv00zvttoiUJP/AHf6DAlOhA/lm8wyWsEywNuFi6Tl1+5UetfcGYdpE
j3R1ZsOPWCjycFOgEiy6c93TX6DsssttuhxY67JijUPIQHOquWUy3CajGEWTP8Wu+Ou5WBg4BfvC
LP/3h8QqO/Nx+VZDhGHR70KQXriCT2fi05AgOyLFrTg6//iPC43sxf3wscrH+JRZR+K1Wo/dMK8F
6dAsDjXFFs2P38a0I4sEEEigTZxriGCNMUR7ERTJu8/je12VSYvafHnLo744nVLJeTSldWUU3LxY
LqxgPNJ/BwC2yIZgZM17M0YtVTdtsRPhl8F+yiw2pxEEg6sN0wpYaShNTP4hoUTX2Jv188dMgwbk
gnEQMm/UquqlboEn9MpHYQscASZbOT4i3I3qtsXJrIkJG74bcObq1hmWLTFxyUdBj3N2kyk8Tbsk
DwP+ZNY6NxR6WDwm+/yZiU5sSM3yddIt7jcNm9wBoQlVEuM4mDSoEYqL0wIYkAYaxji0NNxQgY0q
qvw+6XBGbNFOcU7i5kwgo4Kz0vB9chEXcl/+fYqWz55URN8MQWnoFXhN7c9hNut5Pz7yi4bfaCcp
yEaLI1tsOGwJmIchKFodcuUAE2/Uq0lw5WDbBBLqrg2gisDQd1wce7H2T00klXdSKwMI5dP0RUI0
9DEoFkRt6Isy8XmmDnNn1nZ7V9hhjUmlNcHE8VoQm7LiEOmS2U89oyUKTaiUAwJl2cdxZtJxrbJ9
kNvzObH0GOcr9rHgurzRU/f0wF5muu6D5rhPhYYAWnpsNel595bvdVTcf4ap1TbG9qNPgw4cHaYA
3Sm0ptwkMPsS2F8icZW0WTfrltLdWiw2uPSdvAW77tkcZYKSAMoMxEJrTQyGbmzByi+0WWEO40pO
SJRD+90hcFPRRMsrpxSn2hO7nH1uraM8b8IEjnIek/Su3ou8U2fIMySWXAgl92QNysRYEJDHjvh2
gtj7BeWvVUTiF5BfoVtOMWBvuVxtL9IiSRm5Q+LuSGxwWr+eFFhMF8RrZTcAHXLzeItB+g1PiYgH
3TVjM/lxm+VQWlxcvd99NAApYdyLt1UYZ2eg65dEUTNdskancLRn6Vx2lIaOzJwJTirzo3yFQXTt
ybhwliWLmqJ7+GylwHP5aMIhYtWArmLMpbg0xx7d28DA9CQ7Y8hu2te6mKuvWcW2mImMsBrbPdIO
hCldz8NHQenmiBVwmuRDbsJ3SSAPjH2sP7pg+GT2bUQJZJX7ePjyPMQEm/kEQ2hJMI4bPiQmYPQ/
EnMwBadBcpk++HWezVleeKPkZE+OgVCZlG2UZP9D+X2Sl2hNeai+kFz0QjTOVB4+IvECIj0NWE0T
JLL3m/phqUaO6ag9SqYO+5o4gAInIvoGkH/G8TitSdQ83FE7RZLFbbl7/Il8Oj49AY6LfKMu9AO0
4nQ3gmavImJCZ980j/z4nRWD6MT66yW3oQCfJakbVYLgvYO8GySclwOx9CeggEfW7nqGoZrEpKPh
VUqkPGJ8TWjk/oZsaEYoYcK+EPRgMYAK/Q7QOeQ8HoASYlahS8ZFbY8OrRJf209lf0zXkjx4Dy35
ZIbm18LSybhlYvY7VUxOpTyjjWGLLvOMofwnfuQTGRVekm4yjRBEWuWg8BTrSrYc5eyGFvpTJd/l
xJA85UDyRfOt2Xkc1Zj0vlelv1szXKzbO9GqUXH7t263famgIAwpEwjY+o7vBmeX9Pr8ASp6rTZN
/mJMTIr8SfjPnzKNO/yfDWPrbzjj5ZxktxKA3zGTnybW5WqpzXpSF58uEVZxeI+P5OxLY/hAVPgv
3XPeqrAuZmmWlpdEWiD+VIgH0rkcizyZcGuSVBIMnJFoyJ4Vy6p80WMKq1OZcmxT8do7F8HxnnZq
9BQcLqTzuI5+8wwBkXXyq3hUGsxKnRmWvBfeBa35VMM9tk0jKbQBeB4uMMVxjjY4IPZC0WqZqcFf
L7sUiUTjMgNfAG+ybb2pSzV8tWktBzlHwt6L0z3BoQfvPwiY2QRupSW9qOqjUjanuQ5wjktAXXJC
dFSPRBdzOZZF2ne/gfo7QbQu1PTP9PnlAnPnfpGfrqTJCih18D8c/9YPEJio2WiHgJk1AEOsQN6q
7f1sXrn0pYIG4Bh8IvanNUz92zWd90y9E57AZyuF6VyUxXJkk47uxWRKZvUYoyr3Kc+w7tBS6+Dx
9KR7RBMjufzgv52ANvVjHJDkT+FOKeVAJfZFBkNtz6al5+qIpz+jvpfK0FqOiZGJRcAdo60/wuqd
YyoFvr/WNKGzEGm6Mp5NdAYBN0YKJtDBapDRx58pp7QVT6UKpBT4U7/1p0gmq8Q8Blxc8/kpaLLk
H+N9f2PtaDcUFr4qIdEjIk4p6uknA4L95/vSQoqyLeQ+R9c22vA8uRK9+1u4NGF+BBKPQVMnpTJY
x1Mk+XIH2JU3KsBUeu1CMpeLsWpqN+iNjmrdeoZEF/6Pwu4pO4+DtAdEKPYQE/HyOig5JPu6FZ6d
9q2GOUbmuVrY8SxkBJVpRvVBjhjoo+MIQmSeGj8Lu6PmoDMNkQ7b12pViSKSzulZrkgFla9YeToF
L3feYWUhx6QclVbd/Bfx98egnRPNypy8oZnCyrYOVJZIFPbfvlDaDAhMpr4oThoG6HtZ1tXz83tA
Lpx+kh79wgYfK1BYWujc/INNB/t/sSSxvDpS56gnR88f4RUWVqtNJbGCvFwv4FQUgfmE/HxhzInD
9+CCAqYAP0ZJh6XPz0LrvwtZR1OIjyJXI1o85rL1uG819HCK8qOCBZDNN8XScy+vmK69cVsEY2FX
z5kWDxjaH0/6fLYYo8/YxXuMlsPkp/O/tiUg9MQ+dMP4CBWAIfVXTDFWzBbLsXEdYhzxQLI4OQq4
+2fhhQGWjyinJrTMVsKO8SSdvWYWdWz8X7645EHMfWdTpIS9Tgb/iD16lJ9Ei429dRu0mkSIVat2
4kRz8kcqH6H3az58OZFU1rsJPyqTDKvHcX12uJuOV1fiN+INSBOdXxlvSY4dYA3vqYa4J8VgayDU
MKt4jeTh+2ZkI1Lhh9CZAHjUuYvTQJwUF80LLZ+7yzNC+m94Jd15lsZQE+bmsMj43wIYsLWsIv00
K4FEav8XHIm8zQGIpOfDdjUr5Kd/01srFbomsMTNCM22au/MsQHSeR1jyFr3K0ElFowcRMgJm8lS
FlcrPuiu9xfJ59isgQFC/xrY76Gk17iD1Avxi2fGtENzhRol+k9mW9zrui4hEdnQ6uBPXTSj3BNZ
42fQa90QANiPZefXTJkxiQEDPEhiPH716FjSAJowRB46XPCAL90EK+wxmBiUKVdVXcZUe+qVQMw1
MoulLzKif8NYOlrEYJrLVV6sUtI+EhHNX0mw/SmYsyx042UgknfnNdjzPDK2pirU6GgnnwYkAMAQ
/uiEhp6ngnJJbRw/3WHF+/DfmlUal5Z9UmYof086d462SZ93//I7BtdnwgzM2U0w+IrQtbxN+kTC
35Tk4crVj5C1/1YlXtlkD6WBOUKXUjqBAGqLVQzJAN3DfGGJIxvYqVYac2D/qRfWMYybwuON10uU
gXbSfG4DC0qxAFNXVw2C8J95nehNqw4U6oPRrcTlAy6avPmdAI3gZjUJ63tfI95rJ4kD0ZfPEFxz
hD6yczWKFSO/JJMWAK17hdl6Ocu2wl9DKMqFb1Oyk1TJ0z4JAOcW/OogDJqOCaVavSPXFt1AsDPI
wvlfuKgUhBw/Q79N1+3JmTkcemHs9vtjYtYW9kJZRItUXWGJNucwiVJr9mwcll946imaAuSZ6QFa
E/FbZJO5k4ZwOwQgxSyigPvjNDyOXEl9JIMZozi+MoMx4suPLCBwfLyEJlsuQn3/tjYpmQWAKI+z
vFoIGxGoj07nLLV7XfPSSjSnwL28kjgONJn2ZPo+fQgjhepdVONv6aWokU8a77aHA+19EeApb078
l9XWxZEpnzkt2y8j7a/+dMGnADA8R3baYnwRJihnx8hZv+3sUBNTz09it+2kcZl4oNY2CNjnkgrR
ftxhTKKGCJmmIWi6MFJcfaj+cWombhzmm6H1hPQjoYjSD1SLOKnB+h2En8WlHn8qrZtE/Kzo4nA4
2VC4VFIlQ61ec5D2IvMi0HbNaKnUncw1Q6uab61uVHMmvdMINRvGHQxRrfKddscVmvLQns6sj99x
TU6/eqnae/6QUl3H7oZcYy1BQ5czUEehf8/apAuxvEz2bP91H2QSiNJ7boj0/IwLnTY68+0FfdVp
LVc7QQkdfvhF8fdyzPKPEWn9XqSR29YdxK16UU4sTtnoJnHAAUsuJfJ3zdot+R4Xh3Xhit87O1Eb
6gXzW0isgzeyx0epaaBF9Wh7mgD4+LHcmVuXxr8RHnoF/af1CsUqz581E7+MOVz98IhjZ2+nzdRc
oUxWtBwEBVAZkry/esYxptf+fB9DA6XEZ20B0Hp3Q6Ufl213K7mm5d9eKgapOtzLpMqrX5MvUwnF
YIy//EwRMXmVu5JIEqQSUP8XZUnCL6awt1JY7RiuOW/KQnlgz6ntlheur7njDQnrirEzIdU5fvGN
0ToBPu7oXuTHpboEmdGqOtlYxkqRuI/6YCEX9XocIC363f96byAu6YDRnSNcF1PjUNoZaEC1axDq
Z+ibL8nXwz3Oq3JkjYcbuslsMkuP6G79g2dLp7sbRmtyd4zQI/+XF/Nb+e1WYUXcAhL+P1Rl421x
0q7qwLDrJ809nl8x2cQG5cJSIUenU/hEjCbW2o5eAppl+XkP/vdipFn3C2oJackJViv/s+SiCgRB
Uhqi0amu3/8c58bJu9/+TuAHUglU48xAjgTwAp3KZVXhagPJQscOPuEqJC2IQJXeUN1jWMEg24sD
KkeHCMG0YQjcWM/vACj+XYHdo+O3F9x7RbCzAxdRXMkHN/mx1twQ2SGhaEnrXd2uX6D8oXF+FQOl
aLWURR4itNxQGAif30alR6NVZ9PO1Ai+YCHCGwgPMehBP1UKo742ZgOh1RcHH4nBmSFUgMft4ZgF
2JQdDpQViPsrwLalY7jNJ7uw+BXr3QECI8EAvLyjtOdbajUrbCf36gfx8e2sw0bUPnrSCzvmY0MB
4zW5dB1sRwXYKeyc6siMllgZSOKHF+iBxB9DfnojX1AVMbWEjRLjxbTp+RYvJ4bIGF+uXnmpRSTM
l/4Ncz13VS9k+97HCAFoLAIHpiHFakyduzWmKJ2poBr8MP4ZZr2mGDjBj3VdTHLOo5ToAfIK61K6
mpJBZRLfhHv7Ww0auEcDs35fU3NH52x74MTdl00ZHrijY4bxnqmUGXgSc8mKa/0CxnGU4J10McU8
qh8q8rxq4Gyjon0Ddg5dD7DsA2OYC3reWbfuLCWedsMlZwdFz6jQoyojL+wZDXdrb6MeX6zVizTl
lRIguP+2gn53CfXqUiyWarBasKXogCka4Yn/titgVSldJfZnXj/yDNeOdDqki5v8+s0mrcTLfTZD
x4rgCbtGwevlKMgcSkfEoO+AonK22FcCDp8juKfmwba69uZh9l84lpl0/MSPGAt1PrTOF1qts3h6
22yRLl9pb8f/9p7S89i2V76sA83Q4FD0l+52tm1Jp+aEp+cXs3vnQ+QgLX+7jpHD5KYAadBciNi+
pT5c6UO6rwzZcm6QqH/JGKlzlQ/qjcYdrTHwPr0hlHQgJkXxdZhj7zfbFBjVQGZcpAanqJHm91xQ
YXSlMSJlSvG1YYNUBYZNIvEPRtIsd7qPODncMnBulCkX0s5QlSNvxO6m5CIXRWlV3/VdqT13M0Lw
ms19OOfv2iH6mstKceIm6Uk/A5B3mdNTbQI/7qsR9DazcbfwlAAatxK60r2pgnQC42YIBaJQayFG
hdUT+vXf+w6FdKtmXETyRO+V1lueYpkKg2fz6htoWP5NWOmabrZTtHxhXj8dM2f3S05MeUVe0S0a
ReMV6kn3G7GfnWRYQId/jwat9+47lIFxBUa6EUjH4YPN00uBIaiCkRXYU99JlBaNszWK++B4+Ip3
MNKeiebfi+RWGFHe84QCSMnOBzE7ZGBaBJy4xO3Z7wsn2UeK/1Dd7wR67m4sbPcDlgUdFzOZiDf/
jp+7UtUrh3K37D3pruAM2l89by6C+hXC9b8vki4W15v5rNcpPlIM1ZobLT3LTPLKD/0ouyGEc6Db
kc9s3ApgvVn2uYp8as8piIn49rbCvTJPoyT7+STMc9DjdvO3uUKM8gWdqI0xtB+Lj4XU0BV4oqvl
Le2zKyKivOjiPPpsjtRAyK0sIdbhF+p7xvhlLK+mrKErGX29mTBc3fBrYNxxCk5IxgtHyFS06Fmc
Nxw0KQcQZWt8XsPonYI4v2Wqk/hesVYXEQbgacZm2YK0nMDJmhv9tsswYLHKJCeKrMd8bQXq1vy4
qDTzyW+oemwtcIZ41sSmZuyDoUKEE3ovWsaDMA7QPlTu6+gCJzQH6QtGTI75RjHFn07eEXyiIHxL
387ariam547LNOiu9PWt27ACk/QqYmhj7aQZAF0kxnXJ3mUE549Qt+tvKEmrTYZ9uoESM9UyrR2I
g30Q7JsrVJOiwZuJfgCtNBechD1/60vKj6qAT8inOwtqudYiTjsdHYgeyYzP2r+OCD8cE4Zbvfhp
cCIO4l0dRFhVAPa6XBcI2BJHd3SBS5qXprP5BrhKFrjXVMGaYzGzQ+5WOcAlm/UmVebF2eL+kSIB
oKLCVYu84NzHfsj6+bfJt59J+gBLUXuPieMHCi1Dx68x7nB0HIJ410jSYw412x59jJrk0xfWHR6a
jAG7A8KoOsw6SsruwzdKn4HJZtqIuTgOxCGKiWLrEGpVRvETG9VLZwXPvGFPUxtfNiXjsrtV7mYk
oLFBH5JnZ7TrTW+4Axjxyk04HJLEuIJNsa5j9ojTwYyLPuLusHnQctVto5uTetGiy52ITyCE5L/I
Bmx7OI/P/SO4hIEeMeBgPcq8h1gqpKiqDaA7BZKEL8KzrOpAumNWZUO/gMl10dIvsRUNSuBw3LOq
Y/CbAjkRYzWbJDaBAMM2zWQ7KM1Zs0BDCpZAzUsBlvUr/LqLdCdILcA4TayhdZ3Ab3+Uvvrop1jM
smHy7i/yeWlP3/CCxF8uKapkzSgCBfDTsEsBj+xe/yyxAM1I5hVLTJ3oMIL7ftMSYKOMjKAnV/AH
43DNgx37FgIwnusOnIQUkaQCP4TFSNOruwLnbN/D7rxme9wCwWVUb5S/rbxqigU8KtZcR7j4/Tjz
56axfI1m7opTN1OXwdL7pSXvx5UTehVf8ocowXul0WSKCPYCh0TABZpkKeLzz4GmTjDj73Vg1StU
4K8DrpwR6zZGsjp2zndqh+yMc+M2lgopORK8o0Ot+mq5rcEYvxbKzcvaJKB7+ORRn0qnUsQ0LCxs
KGlYOJ4LJawzyaurJ6VLEn/PFrN6MKgJPwPsJDWgsTKLDAuQVybCYoWUHbw5MJ1Lm3IdLc8OjC4U
pWRs8HtcL93taS26zjoiY9dLDBrG4mjOXLyEjSj2sB6TFkyN2y+dgsM9SFRgsTu19yA6kgbnWWRP
G4BaHOFOGjMNNGTwbgNDW9IAoeaN//QGyVSiZ2ZJCUCjwYGHBm0VSZx532QKzPRblw/F12ppwXi1
ugogivPfENfbFrWSoUUm8wFecxJKyELrXusO4VcgBtqDfwWqMCPgg8pLvj5Y5rpTwEYj/rKmy79q
aknAxHsXgCCGkgtYBCqfdY1yFoAhFvnUK6k5jTdIQAOCP6/mKVUxbpI7id0HdMWXeKU7wqduGwdd
CJfxEzcgC2bwl5Vh8lfj/uBzKB4TAqRw58R662p0lVjsksyIyZ0r0ubeaQSN6saayrPslOdVOaRD
AGPdt64md/0UaIjWgTwHJYanwFrq4vME0kZXRc4MYH3JTuAR5guZAZgsHChRbM4AjzxdVDHrVtx7
nVsUcqhl0tYc9RJjmcoTQGHYxtJ0d0fv9+fruk2MKRvwA7QcI+5pCy1YNPx3i4sOMBOaj4wVEtDV
kDRrcQUZRBiicOFhgT2Zwe1TNIlmKQadbxSLOMc3wsyvkonIMmQiDxbQSJyyhxgPtiY5mADM+vg8
UPN2qcywvq5h6jijl6MzVs561Nyqisb/+IN+pPp8wSJw+ds9hc8q/yqD5Cet7KxNfxUbAUnHkkeN
KRV9WKF5wBE7fQmQz8hC6bicJpk7NWtICCTeBRJaGVgaNk0UCYXOWIKQbNHh3N9yl17ve6MOwyn+
eOjMNLs0O+imDflWjCwRRnt3M4pOE2NUfXtSCimIWBHXu47fUxZ0i0PqlkfxRfttZbmO8OtZ9ZbU
GLnPkd+QU5Z4lQk0HR0lbwmwI79YrqI30D+QQYRxnQJWC6N60DgvjEIPgvmm5OpfplC2xcS2BZpz
XsyCZyiWCGC7Z/xCIKo+WCpKz97ghvqydc7cZc1QQKFza3VaqpUeFJTIMMymK7Pl0RMh3erh/EOg
Meb2A06/KEIoPLmMYWDnyteHzvQ/V/Ea68EvhzJGcXSOhVk80byYBAggfZB2O0ZNBJO4CbTkzQIb
JXCvce+eXtiU+VAIU4seaZg2x99A3cfY6mfuA08IU7vLudCCvnalmcXN2hVwACZjOyAKADCATJ/1
rEmlmYDyboiY6UUFOo+xqSiYeE0ICEx02TCKPTDCr/GndUG999UytsExsuXfLb8b7Wbk/yDsbG2e
1fmId1NbYbSsITHjpkRF1DIbgh0f+XiHke1TOsy9BZQ8KJGC8rcPcHdIIh2uQVGOkxSFgk6c1mwx
yyuZmMyxvsnW5VXqEz1CxikhTKuB09P3XgpmIAczpAlI6mKTphb/yKNrp07kV7IX6ZMh7a7ZQlHm
BdVlYnN6x/qh6BilrGbic8CaY/QR+5z2Dt6gE/ZSTc4PbjFyY5eVQ5qb2CzSKmfLtZzMiMatbN3Z
K/KYA5lYJqx7HpV5csuohQqdlvJ4iunnZmhzAR3GabCsobn14NMIgIFPmlon4RDeKE5Q2jzrgRgz
5oLOrbPETHnCjuPZ+jBH9VgEpexpdWIJ0P+KcrfI6nJK+IsifS+Nz+qG3NM2xOk/kk39Jdqt2uNc
/LhcFSg5IB1Ng/6FWGu24w+s/9IG/aSEOT8GWR4HAZgjt7Qam1JFtSprsSdaqRGP8l9VznCtPEoD
XCf4VT6oKDlUglPUsglPEOteS1lOYLe4ScYRcad2GqLfLd7UUvuY8VJHbvshDaBRF0b66jXeH/z7
prgXEztQvxIEkUEzRiufmVrx2V93gxQikjEtwF4x1Uq6KhjEaTdBCNpofoGJxQFkPTi8uF0BswdF
1bYD3qa8ZJqcOrme8/3yyrlUUPxmIrFQpA71P+HNIN/+oDuBHwdNQ8w/Yoy2ULjsx9dq8WsBsDCJ
B0Ht4ZDJEnP0IEBJhm1j61L+8cZeImHIbPzhJOOl/UoMc/qgU4+p3e9O1Tcp4Ak7RBgju6B/l23B
mq/e5Wu2CL/g3cHwAZJngHb1frU4b1+ES0Xc2bygAlK4z0jrT/2uD7aVoFT/osXPiMBMUhsmPRfk
/HNF6dodYrvwIlGNkvDU81YSPGiL9R4cQXUJA763aQozxvhEc97QUlJUK4gG6uCpsXckQvDBE4b1
JJkeg6HXDBrDoWp30Ap9osd+pptcUObKdN6m2RZ+A6+e/QKxviwvO1o+DpOwephNByqywlchxVde
aoJ8vS58rfJsypftu8TmtdNKMUrs98ffayEZxw2FXCwZC9WXNi0P34Utj8a896qqw3HMctilJud0
VmNyApEQURZ57CU0H3GFmhR+bjFuZJ7bQadim2Gx9b0cHyk/eWQXd5VIPLtVCIkLLQGLNuNqLgoX
eAGDYLd1UO/zj8jrp8QmS8g3BOyv/BnHHpZCmYExYGeirjgKbgxPamg1E3Tn/a9PK79Z4Ncro6K+
7IPOa6bM/IRBJB6Czr8aMC+eA37EyBiftpQhQfc9PpoZi8IZ8QHgOvEmlP7Iexfh6ND80mlk/4IY
tAUOxkTwhrs6czOLHdIBCa+jXdsklz4UQZEwxb1pyPvK5jzDmlyzRGGBPODrtTFU+WQ1rFoqnhkP
cAiTQeijRkjWYWGqisCiRU8x9RK5KwjapeqXotNrgbryttbA7J8IXD3Y05IIz9k24U+WJCNbaN5i
SHkl1xsFhMtPj3sWPe9AGH15xPupeVeb7lqWVugrdmKFo1DWWqhnPM9/vQT1So8VsGmOUnAeiEfA
t9NP915aEWl26cKOsWVw+r4qreq/QgZtoB6U5J9pJWZl7YTVE2rHMeZdXg3ngnTXDZEVTJu6Ak1y
TJa6pMC8fjsSWFjJtRgSyk3QcB37jQnHrQ9VQX3hC1AV+HXNlx6jmxsKvQvgVzOMwJs1M8cVYyYk
rVi0J7tMtH5I4rmMj5uRUwTQaYd2Z1Ioxxv4kts0ZUurOaKxAMkr/bdeowkn5feAebLD8FqTQTPM
4cQdAVji/IkR2zqyl7eP3BIb/3CQdkIwyiUS72lJsT/xJg4SGddyY58HHsQyk7xzx9Ny0VykWD6+
ClPsVwwN3sQxdma23joou3fRmmnxG49n0qTKKy8Mhs2x5rs8lN6pS064IJ+ol0GRV0Hlq+azBtH/
oDkttcO4VQrOs2SI+ogfmYzPmX/RIx14f/LdbkpvWcWtpA86mCQ0l0Gi4aW+ZT2Rsw2+WOOz7Wjs
w3ybC5a106bWVKIexUs+OtiJJ2jU7Yf/XKYx5zXTzWjP9L4GUwBHp7QEdXejuOISD0PeVqxvimo5
Kgbgx2/J4T9UPMgMGdIywvT7l9Yrm9mbzj7dq7NxJhwRpdqNfsS8Y9/z1pfXEhvZdj1LVBcXzap6
LQR4HQi00n/TL7ED17LAgefzIx8tAsUIJaPNWKUNQCqBatr2k18nkwvJWJ9c1Pkk1rVWuG1jSLyQ
Mus02PCzSIa9P+6Q1N1iaRPBr07BZtTJl0h5TklO0oGOiak6Od5GZ4d6JfCSe/tHdT+lL8Qrd97T
75w2v5YtZsbPBVIGuYht9iydP8Ps2EoLl5dT0633+Eyi5vou1Aojtx1s85Y2ICdcKW8v4iL44ats
fPxqO4mtf74EKBeJljUX1aR+LKMpvoz3EqdVczhblXERU96ZnAdYVrpOOEpbq+8ysB4Y76E0TPWq
XclQCYAeDCMu/diY3IWfr5OTV2ilXuam3ja7hWytjNi/DtGT/ub6PhBMob8AM47D0Leb27SaPpBh
ZurKmEteoH0RFx0sqk9N95KpZVnN4TBqav08osAlkjl6QXXppqwY5rsuTJtzONaD702x9tHl+pgV
k8UPH2p0CxDYipc6MBKC4EjBDmoWIhne54A8DLEA0JzYy8Ve8T4jpged1qcgg/dkAbeGSuM5Rf5Y
z7BwK0dBAn4qI4WROoOf86RW/BS+8upzcPbeUC3+QYiiWsUo9AXx+S6rHZFMfi81G2+paVDlwZ/P
nSVAgwh1W4Nbtugm8AnI1m1h8BnkPnglAjWYgnVM2X291czg8C4/w34o25VWfd582DiwJrt5nnXa
fcstOJaAtoxoIWgiTOu/hbhu8ApHjnqGQH/hrJQFWD6RKEJI6UfUDKdlSmLX8a/MoLPLW8A6nwY6
6G3t8ebJwl6s4/GzxEBdiPL6Q4CZpHdrYzSRlXZO/ga4CdGuuOxxw05etiSIJVadSfwMD7pzzZjr
9WjoNAbKa45l4JkAUSSNOkYOJpKU4+qcTsHcIOcGfNhOUBMYI9jHGEDexLtlJiA36dtUoK8gUj2G
q+SI/8ehUEckz7OSG+svQLlXTdkyYEV2svZGMMQ2K8eiU8R5zfi9lYYfMzDS/UzWJBrHemt4u8jF
xnCrW0PGkl0iPb2e9YJ+KAa5BiKCEK3SGsFy8iUyL30PwkhgdWvPk/pJq5bJNX8Mu4OKZwt1hfhX
2a4BZ16h5KqoMnQ+6krBrZqF0sSSo5/Ab264mOtMnGLgWblbTN4iXLbsVou6oWmIaO5WziXd2PWo
qPagVw2V9vLfTgThe1h02zA6W3Qd4KEuOubNSN+EzuaJJWCekf5HoGfFOcWV/1GwVwYJFGJ0ijQO
i7750AftF9Knfai1OBAnVUE7zbGsQh2ce+JauxiOBmLmHpw8wWucU7jrZoKH5GRT8SAM2mQP/x08
+nXZxGtLYvt4+LRSLrPhEeVAEvIUDEzhN70FC+oqJ0osis9PosWpHREMNHh8WJFQvX9lYVwTg9Jz
c09mlnAQsp7GXepW7tpcYMmEZJHQCG0JsyQtwNxvgD1RUk/Q6OVraCKhQvkXtEznUqyIp7/Iwly5
ECb28xkxZS2ooNoOEak6UFhaJjVnESg9CltKCVhaJC4cI7JZ0YkJtu94mBeVcuNLMB58AB77/AO8
YWz1qfjszi6jZanY1gLb6+cOFKtmt6oiwCn56gIojIrWQ8RsgbCoo92Jl8m5Ni/cil/PVN+rdvU6
Nua/2uZ7eGB4dTD/oNqB7GvnI3szAh4mlW2dYqUMOZ3k5iQg1MFgVm2qQu3l0szP3HJomCpTJrFk
wefEr3qvTYP7sdo69WNebsApFWdQUGqIJK+HegiKUQn+4K7TNgYXXvgPaf4R864dq3gig7p8/UPL
wVcRJb8RSEMx+rUmtjSQZailYACzLZ8/pO956+Eb9kIXSpx05k7HZqUg9F7JQBZhmmJdp7JHNduO
07npuuf1NryHaAsc7gaCR8h6FID5ONchH60Q/RAhsOrJSbrk7goR53eE7+5A8Df1SfWz65N3RCI9
ocSrUOY/u2VqRmHQMxgjxTOrJ29P3rENfVrNyOLY1+Ve3w+/EQVEAve7rcWz9HEXDsbp2jxe5d6Q
VkWcdCS8Dn+KnAtjDmMiAJXEwYGERjR2zp7NxXiWBKAr6xFiJjnvnmrCQEsec6r90C6AbJ4HDHPD
KdpUx3+PMVDSsdkHqpSg2Jtd3x7irNScGaGYgTLHd63gS/8vNbGVhUliI474vl6Cr876v8cUdWI4
YW1uAyvDjDTxgIyu/IDhoN+Twri7SGchMI6pbFOZFj1GMbsS5AsHAggXz9U70ivCiEDesLqpFy14
NQQHERXnNvldAKtMVMMQBxeSIftfil0N35HZmlwFhJ7jaWQQUA4SxwDyx20a4A44y+bKtoTzDJbI
Wm+e5FqUq0HyX2cSlfaZd/xFdZj7/pF1rKncd9lYKJ8TrMe37QQR/Lu3FYYS84Q4YYeweshTHICQ
7kurSy1SzjbJQIQGpHCCIrKWUdf3Up+TS8pS1B4wVQTGoceizrhbMU2BvqBl8CTfiP8Mej7kcUYL
0Gl2tZwj0Ze1AiBU+fVrINVA9o+I7hroLthtRJBbF6d/a2xN3yS4zv5qWM34i4730ysYeoWSBnyw
3w9U2sitYcszsC9/oTPN4TJYifOofDxINNJYe833hsYf3LvGMeDb2sXj+yqEcTwwFcGTcUNdmM3B
oLQdfAAoEOfM6SZ4bgHk0WEeJ09yBA5g3YW5yuYe1VsXmT/Gb+nNam0HcQfwKcHtniW3GpH+011i
JH7rcB0iYGDQl8ecoaUH6FtzUIgbN6Qw9o1tT1sYmAs1de1xxmFBbnUvxGOJztjyh69CVCaf5E53
qbxVnWsyUQkm3HJGiISfafibK/20MJeFCXkSkE0tGCOBLV/aBRSUi5+CwNC8DJIQv1dU1eCSs1bY
gLHA/Ub334YJEd9y+tgfC7XhFPaTtAlK/CF7fe4Ips7B00IP+8uI9e+bt6Xkpf4PdJKILyabRXPf
7LMp4FmQcxPmG4p5512eWVnGGesyRIGcs6YdVYghItJkLgCOaE+Mi5d3tjRLU1YRghfTIYQ/IIQd
7cwTpotsFxqg7hadbFHDLVoK0UzOAcUlCXIEmM5dXoSKDmZSFLrjouVuINAoDsW+He8wSAlW1YiJ
5oGd283eS348nJxS0P+PrOSIqiVhoTbwlhUfczYjUnGyDvInxKZ9QPf1ntHu2B4OkypGHrojvo/+
phppQNjtGBMXW5OLT7GGm5/D2RcV0Uc7PikNy6L/hDbgxm2lJ5fzp3xa9BRLG9Te9/GoKETeGeu/
Q2E1oOdXRc8Goylij6uF/ED878lN1qAzqdfKVxzLUT9pLJS1pndL1P9MwLs41/jSbkSqcHhfryZg
d2EeABYsDy2uBjRCKwF3tR1GP54Mc1Ztj+pPsYQ3AKlBtKJRmzR+inL9EaHd/SGotCr9lFSQiDIa
0E28CnIcJHdU+fLfKCGQrD2k2L9fmH2Q735EZ8frxamJM/iaCm+atLF7I8J3LN5pp6Dh3I3HuKYJ
l0gS4kZSIZG2VETcFl+W3QZzRZ0dX04IBwUjrY/jtxjG/3d3Y+uSvG3pe7yCrpKX0b36zrL9NMTp
RYlZjI/uX9JSbIh9C8a1aAw8lwhxMDG2iu3VcWHZD/RrCCr27pYoymHYO2P3HbPc3YEoAUrJn69U
hc/z3KrZw4qO8I6L1Ozj08gbZGiHn9/OCt2Laif26keAIb5oPvjhA8k2YVRTG8xYK5w8JC9Kklk8
v52GcG/Wjy4dtjOGz6WitMUPzxjN2twaG0oWP8aGQrNl6FERdpihkm+87u02yHZDCltIpUZe/T9m
NGGABfq00zw9PyZhGxlTGDa+UXYurT67oVPkqDgmuy43PaRe+xEiBbcF8I5oDgUEKtEUZ+JN0xfP
HbZlsb9cC1jxPsE/jrtIDFmuNv1RBfnCVwfCZRCrTmmAgwAqZbEV3A7fK5CiK0e1/tgcwvJUpdUB
ZTmIdq2xxxdgrEbzaSoXWObeNN8c6wT5l6NECqA6r1idn8nN845YQ1sWGy5a1PfSA03YmzJXltLu
Yueeo2wbYcwzpDmXxpno5DRY6/V2gv2IYRfJMzqbWzi++z2hyyKAbd5E3TO+hzooWlcRQcqs9Xyq
R9+scIqXdkjIN2Ue4YBrom0kWOUkbf1CTHV6SaDGQphVn0cKbFBjQuFo2lG41m2EEHOiq4Pwt7b4
9dKYbVgiiLE9+NUAJtEVvTq15QFKLfyT3YlZpdRBfuplL1qs7RGmciFRtQa7AMdXMVmHZhIYHvW2
I4cOQVTeIDz2WoBKgg9F7HvqoVyxp6GdL5axy5i94NYuh20Q6Okd1I9zRXKFRL6mPtER/1FwS9fk
hXlWO76LsfYmBReNfnjMoqC2fqdOecrMDbB8pUSYtfAvQ966BiidLR6apg+uKI3pLAX7ahoNFW1G
h3qV9pAMbEVz47F6YaeyTCcvAbktDSXx6JOUo6TrfW3sb9n1pF6CdqdtfzpvyUOU5mruntoZ+uu0
i3ZsXc6rXm/wSiNrMqVoq4BGwrNuF/3V4w+4SKm07sVw0aJcco+fOH4dzT7caszBy2UTMRQlxIyf
wOxxhpzJftI1Eys0p+uni83rmFEzbpIu+HNJYaZo9PC0A0AbHrzqcFHeyzxNN4IYA/C/u9JYLZG/
I5PO1yewZ4jissIqUnBDQGhfe2cUkQSzKi/feAsKkQiy+nYmDuFkOFe5SHHfxpo8DLKBppgTjqRk
kUgGcT8rpdAjXnjfXPmzPi6vZEKgpeMy/QfZUDoA4FOSI3L3YsfdPek/3DGbZdqJ5fAh7o59cGIh
TUpSv+1mVR/KMqNV9VbqsigdGLOe1bY98Uk+iAP0/L8uDnqycqNgOJJ4LWJTGZyVsAVCJhYs05WZ
ZtIT07EoqKiEV8GlCNBvQlVWwc0JuaNKJR4VjuL9FrOy4u6Y1tBbxJ5/iKT3tcIFXHEEatppc1GQ
XLtHGmoc5hVdJynSdZ2Fld2E+Kd5BCbA/HObnuNXCnhNjx6crGFuYfc2Xq8mLdfMK56G3qirh7Ih
GjNUU2m9p/LSTiZW69lOw+eVHjjWK9QDDj548k2ERbVBvztt5DWvd3UsmOQQ3a5XAb1xEyW9IdIK
PN8DLzYpVSqtPQVSNp3CqrGbKruc8AuyLI4W/stnFUwM9rv+GNZFK4jGlw0WzegbSSkkh9vfUEBt
HlNwh7YZfG1uaQIM40QduAOvP5O/US4p6alFwfBhF+0vpH65ktvqihw0LDVn6xcsaAqZYK/ppxhn
GZ12cmJMZA96p4nR03ggzprtXg5O1DqAzC7ozl7Tuh/JIsG/ixmqOea4I+ezv1nH+ddM60mcUGns
kee9aCiVjSIwj6O+2EAsroiUViuFos/I+YfrgAwzmHJLCmz+66ma6K7FPVAKIJEQfnkKNmeRuiuG
+tiR3wbY/V7dSXAkD1SYuPQxH6BM96FzYd7yWvLiKRgav16/0HM5t+PG8sZ9ZcYrNEwxCYConDnj
VB8GzupHgs8uY6yOOuiqRmqFBTAzvrae+OwIXbjQ2lUHHkn8MFwUv7KFd8fNEP9FC/IeQMqzyL7+
r7F05SEkJLj4XSE+fIbOxTGfBXc/iS1wgZZReTmRPUcy5yYvEnMRYwy5prgJAwtVZ+h0PxDHiZ+G
vlQiAQm7ji/zodwn4hC7KGqOz1KHrSqblD97b0QXpDkRf2c1f+vapBeVHWCy+4eAo2KPDRTK/iX4
ArjozykWH2pNUnxSiRnVrLktCio4Bm58lhFU9DIDFd+Q6dHQ/vTDaLtYLAmYJRF/a/Y5GT5Pit/j
bVhqhiBaU8gNS3QltOOsMhnRCEpVrX3TdXzm2SzY0SokqPVWSPHUXYsWEqJHJuE5ankE6xA9kljT
9TaCX/3q+I8KfWlW6pEsRg1QzjeB705HbA2zWDGjFfO5kcFSjlkz7yVSFxXA3mrmRAXwCGh9iT/a
/V4cacljatqYEZ2oLYSyO0wpIkJ9Wz0A2jJlF5Ns9i5jODvFFM2ZwMc2nZXmcyhtjP9cCZnciFAT
emcU0ecfKnr7mkaLRZlw96XpAhXinz67hyqOIlaVEo0Xi1/iDUbPgUt1DE6//mSuAG3A+6P5dXvF
YTUQ3nVuPakVu6ii3pSgcPsvIGOYY+dZWEJITSXAnJig3cHhpSd6aKjcvraX2WXPFUeKAT7BpH15
0UHzsql3tTvqrKdcGWjZx0mZI4aULjT9JK5hTf4tY+ghMv3ki+ak+Lscz4baepbPX/PcbymkLCdg
IAxglBTvuVbNN2IuJ8blA7zdx+dT1K+aLlLS0NaOwI+Hb6czykLkN56cwDP6SQCAbiv6sd4XYzsm
8oIkUsk8FshJjpN+YIdx/IpEF8xy5rksHfJWpRI8hL2u0scD9D8nURIlhofkwbVAJwsCkspuAvbj
KTrILeDs77z+YuIfS62XZCA81bgVjtsrj5vjaJ518TOaHacC8mngPGTa04yOdJBCP602QAYBTqJU
o1nAtrumw+qBII2JLJnWHcQZFZ2XgMCNYnsQ+LRdgW2xt6yPdNom/PAI6ZDu2fGrIdd3fKw2ab6+
HyXVozWMoo572KTPQYJ2jdMKBvnrLF83DKcrOtF3P96VG59rfB3zBq8vXlgttoKhfWhiWgjeJzA1
O/ff05jzmh2UmfQBtLaNDohcUbi6JTGm2G5vJJNVkKkMhfbqc5oSER8O/oSCd1aDgRYbC3HhYqO+
QDDnyMAKIhEZv52i0GvAllSl9OQsEvnGpyK9QOCySxdt8CEctjBjggYTI2eGcfHDomRWMPJDL4RB
nOkaknmv/6hqQRfe6Cvi159VX3tMMRqG20b3AZvhBH1B9w2vMbwe/x8HpsAASNp4fKJ+6Kmue6Ho
cpoBiBl8JebBfdXrbaHVm9mnq4CcNJE8el4+FyR3I0WUbXVlglaYq5tuelhyoUM/asR7Tbw5ffBH
SabI6TJEyWmR9zJ8HR5orOrGQEkErJljDNf7N7GN2esu1JR6y0Qursg4mOfvohFWNFFrWVz1CSXH
mH0eJyPrVjab01grLYx8C+7qcgZWSaeMupU6y5oj8nqo6f8RiYHAzxRPeZDYhcpx51fvH7Cl+Z21
dUNSVBeqjoPhavfcWALB45G0u1444yI5Z56uI30J/Ec+mJ9pLNRdStmhhqFM5DyhqTD4y7F6N3ke
+A3EzocIZxhWnh0c41CPlUkOmvcqrvHnly31CGR3BNX9NuPLVWfgG3h01FlFFpsURyIpPRPNaQaQ
sWwgmpzz66rOR/kVHrfYXINFgWh+TuqUruqSAzqQWEGeH7+ZsOxsE+Uf0DTW//jBhhz+t+My+z/k
8G1QnYXSCRUmFG+wtAlZSlMQT2Qq/H1QfxRsZPwANE04aWIw9B6Z819Wy1gNZ3ELT85fOre/II1O
QytHhazmRQ6Y9cp11uVYZ8nF0hPFbbnu9I69/h0bh78NjJrnCSUEABZbImoBROsRbKA8pE3XXSYs
3wImXjbykQLRWkaAACCRCoP/IM4HY+PeVlaWKYgpIreo6wIRtat8WNDw9zp/MA5pCywCfouOj08a
gDhPMPjVplqDiulI9yH8DLuWXzckfTEF2nprxrG68tMUF/yp8ar1xk0xE6EcpprB0ON1Xs2QtPOc
PuIlW2Tma2Suswk0EqrcGiu0e4azW3V99jdIVRWSsUznKOXuuBfukkQf4bYOYwX6EHTvLMUFMuSI
sHLUshF+q0G5dXI/E3X0SilLEj0vnLkHiXcgk76VQVgQFYnPCjIPGiqOULdf9OnadTBerwna4MOs
waQqyo3npdUw6EbzrxoNwY0m+61XIh4evll1PuQ/s1yre59GRaTrqd7tSm183TA89GJJCr4GsK7V
FgKW6zvJ/gjvHJStqwbwWhg8Iu++Uf3eG5abJQG0XfJaCzF2Qc7LWwS3IYeTdfTjaPqyeHWdxrBE
7xpN2iBL+AKoc3EwtV1C/H8rS/gP+Rm50dX8mfNBUwTAxu1db25rNeF0BX13Tixn+VW5aoqHQLDk
GY9y2KqsQbJuqXK42rXlPJq9wtuANeiGG4tnhAMv6ZDv7QQvo3gkzd1MExom2l8XF8FM3l55aLYB
uN65B0wvlOBm2GtXG2l5MaN7EOr+WzUVyKSXrP84VOt300ZcIr2KK1FCSIVgjYsNnUBB6Rnu7MKl
XSmX9I3vaLuJ1AQKh9voRzDyjV3i7OG5MKAx1tpHBNZ2enKQ68BnXrrghvbxXmNGB5NKK/cpCW+g
AnmO02a92s1BDzs0Ufvz8GrrdUf6E4nw9Gd5RuY8QECSrTKkppDncuwEICiHt0idVKJZwNTx5T+l
CyXM7TQGs9iq+eiVCxDguEsZJtJAATLIRkfE5Il4l70+P7eS1fmHZFW8M8s47Rm6gPzj5qGqNpjH
5LwNXwhZULeDJoj+ULJ3RmHQmAbOYJN/OsdmtM3eD4xRdAAiSAeSXX+1nMGIW2KnpEZiwmJgyg73
9IW0Z5MqS9UQHa+Yc5EzmVKH9XBXGQHxS1hsKvwcuZ/8QqALf35FMt3GHU3+ZecADRKIragP+oi/
UnpihkEXmsj76gq8iMPlF7b6jgmA1xCqGqAYllHnA6+T6ynXr6o8+J1smokRVh05E+FyHzPxFgOu
KHcZ1wm3lRwLvvdcECOTiFgDloEUhrc9VrynmKsEzuPWYHyBAdpkW5wd4i5+op/NGhgB8V+i5KPS
bi4G3GAUIKdONt3bphipn4ZAIp/DnwmcsmsR0ip/uHbxlKPlYwTopFzsfBgzHDQbX1AVSf+Q7y+2
N9CRjwgT3UqgxqpEnAdi2YOi7Q5M81IlCFRoQpUhc/vjQhP/cZXerkj1drjlo+oivE31uQBaPbJR
W2y2tzOanpuyMPlpRD7SrHTGZM3n4TZs7VQ/4vAfSxb63ucwHuFB1cwBcUsckDuX5IR2Rh7pA8aX
VSASpXjSi4yKr3fgG6oKGdGZAMu03k5nk+cmmEahhyGIonffOMOV43rInEmN3llm6fFptk25XvU5
2ftR2i02wkdk1zJ6T/EzlcxqerthtrOCYxE/O4Ytl9uuF/D+qi0QLNUrYaKJjXd0nZas8EmHkktt
Wi3GFCSE0zsaw/pNGayP2Yjpc+ZsjfsZVcsnUPED87PnAtTSW4Qmwbi92IWBtg3l1ow14jCQuuIY
k0aTLQzTP/BVwQK+m/5juiIxBQhIC8ZMRuUrnxM2EaxGF6uPRVCMo1ZKa+2Ru28agRjK/TFvbrPO
eyGuDLnW9zkq3Po7bFRhUmx0BPkstdin6blfb3F/XXkazokhZh++rPbuo+z/quxhcBgZgfi7O8xz
1pgT7tszIfo3SOfFWt0BUzH+bhCvihbI/6B5Yv3wxew1PIASB1HL0fCOOz4pEn9qAG1IkstngFrx
dhtnfVxxXvwPQ7VTFm6fmulHa+PidivtDWY/RVHgebaiPYRED2Hx6ssGDm3Z61l0q1f5pYeOR7DJ
ds1miQSgCVSja6KuGWQ6/B9wez0OweaRKy3WAc9Cr07bMZBOiZNXDDV2p3ceZvIYGRL7h1wb6fAf
h4pOpinwQsAUjtnnjU+vMPSuXL0HF4P3r6osGTY6m0+ILTln+aBUT0ci9KpL981O74JunL//vLH6
fG0ev8R+bSIfuMGGw0xt0JCBDP3/yscFk3wQoLHgJTkFvD2i7Mg34DmE00C4llFZHasciZjFPiKy
q65pPuL/f9Kh82yTP/JRHxLV3P8oJNYm7jjQkVgRnOS68EUb5z2Ic7gritbUonL1gA8IR4Xfvool
fSx/u/wH1NU9usqrrFwIrCSm4H1qdWCy4X7uAYWjHrk+wiYGRWF/K90Bvto5JDu9IW5jG52SF25a
60lCKOwpgcMVmSgdToGxTUzPV1Amf9vwzTNl508QVlEB3Tn7NqbCjAGiTGRvazSgnB/iqIaR5IgX
MNNRnWO8NgdP8JhcTaR3KPT4SbuB1192JgXn1QtiVwNWTlfGREjAAqMuGSgO5uIyNQS1ObpvaLLJ
WvdGB00DcqpZX+6AKL9RG99GVqhGobMmQDBf0LYuw5ILIC++NWAyaVgXb5MVft2Vvt7FpzLV5yTE
kEyhxK65t39Hd1iMu0YVPBaNGNB0Z+BepvL9OvQZqPAaF2PjmV38201SINa8v3dNNCQf4WkgNIa0
jA4GAhGgdoSSQtqccTQ7/8seExCfkr6HPTa70cUe5kuPbiP/8GXFt7xQXaHkW4bN0N+dv/Go5jKq
ougYTNKaiHIQATF8r27jDQUul0K+zgqYSfnJFQo2QU16r+5i9Nrk5R7r2dhrgf/blmjfXwSMBxR/
4jNa0ruBGHAUFhwKUnyoY+8g84P64qVUTENJUH1/BqbHDmuCZBN7q6et0KHBHn7UXIz93/PD1IOO
fLxPjdqrJdcDM2uivHfimMNlSPDqN0yRzNsWydxOJtqW2h8Z8Q4Bi2HDtOuhMUOBFEPCMgQ4VBNg
qeYsrw1FBk9FFnVIN00o8+vxu5FHMWGtE821oKw/RMFQ1SLbdZOxaYUOpvKY1L4MVcu6ytj0YRZe
Sp18O+6YlEZbjMOJevRDKkHgsNjK7fXbhfEqDY0Cx4kNZpUw8q44/45El+0QDyVDWoPlDpr1fZNp
omcjLX49knMnWeNvvvwiuJXow9Nl5pNzp4URG+/aYuZXfArQ8QKB//To0z+T1c614i5b82BSu25L
IB4Cwa1/zIeXnpE9bytcU6XG3dTSpvL31aanj0cFqJZgs34s0WfAkm3h9cQOsUNzU0QmKwrox/p7
a7hcejE/91/tZvfhRF63mJ/l3KkIQ2+OSdeojNyfBfDpROnyKKhSuQqTbQDxbll5Dk5WVIcQdMQq
rw6Dg3KtYtxWLPGXeJuHvE7+ObepyKZkFlJEtjl9njB3xv+7v/FMyGmdazd8uMvlCH8cikR4XmId
tAe2kp+JLrccpxi5Ja8LiU8B7jiCxXS7KRMbFqX3Ucj1eCaqwA/mqSFkn96NBXD54Cwukfko2VNQ
gW/ESfoFcbJ4fvfrmLoJJbeeb7SbW7Lz71vzYeJXbUvSF9dMipsc8BHtRAkiXhd8YZCrs+QwcVjX
YS86+dQLq7NP2F2lzBMg8gjoeUt0hf4Y15TuiK0WIgfCeAzU4LTMwN8HlL2sm9785WsPTjFQ8DJt
1GxvO6oP9wxOVCpr2KHFpxm7a3UUELkGCiBOurbRs5Zkp3ZynpAWxy3QZaD4O1oA24K3gIyIDkDk
1kh4cgmO0Rfgh1FYxgqYc5XcPs+k7jR8ZrTmf/TOaqJYElueBL/V/OaSFQT1Vvzj1HJJcgL5KWNu
ba9Lk8FikHfGviuyKZhqFxVTGluq3W6TcD8vn1liKRpbLVDEpAmOBHE2Oba5TTrnC/oUcz3hw+mQ
xQ/dD78FAslJq6WgEn9ftdmTeaBgjwcqX5s2RQ0rMa1aNatHLS2ip9NRtc8NFYpYjw6eFSN7ZZ79
/N5fYRZ+HRs2EX6WFSTsc8+zWD0qKCZrUNKV2LjRnPY8oReNIvnT+EBagRE/s0bFjpylZKgq6y3C
DTQjuHt+55XFsoyWkBW/D/6eW0FBZrQ4GeXl183YVxiUQq5BmFWkdosHC3E5km6kJ0HIyJT5U1Su
PlCHUfy6wEj+vND5FYDf75SqRuL4R6wpa9CBGX/HWZFw2zDYckuRSjy6OxWgFAmbdRmgbSfkjQz1
KlMGSrKICLjok+2m7UUcTDVhQIdHKUjWxw/tOMFNa79wqIKvYs0lkUMSDWboGyhKAWo2Fcx2PQfF
3ctL72xn3+eezTv8aPnmpupok16wEo1XoTuaXnsc6/GXB/EPh5N5vy27VImFknIi6SNym2X4FSJU
I3Da98aQZK9IlvDwtBcNiZBhxozAhG8fnYtjgDjwETgnTEzu7Cq5DwX+kGzYsRAxkMXe9nHRis3F
F42b/aaDUPCCtARidL+TgHnSI6Is/V335MZ7fX0o3xPkgPqoZ21i8Sjix+ycQ4/WQ8xuvYV2YMPk
JkUNg0MW9oq+/ICEQ6enCiBmeH4cGkajE8D/pmtCdjZt1KFFZWxOz8TKuyYQUsBhUqlwFYGsE7Ut
JexVdu4WBM0d7LHVh3XlF0x4PowySt3w6dd6dPi7s+DJf9s5D0WBLZIwe0zljzauTTICfvsqW7v6
0n8PXzulu64xeh4VcrerjXZoExWj3hAFo8zb9EJUZuIaqFEzUyN7dYcYHUS10VZlTgSjAmhiLJLE
5eWRrxqpRONIq4lxUDXwFcUeyBNE161XJmatozi1+CQY2Q5bKY6UZiCKwRenSJ9BnhS+Lk1k/CPf
ES33baEEoTNCjuX/udr4WrioinxuqdPQXGyo/t++/mLerh2C1BUU9xcPVwMn5VEcavmO5ayWzgMm
sEYwyZWiul67svmBXP6Fhh7KCvnggItFlTqLtnrov0KX5W8J8DS1eiHeGIWv4pmVEhWEbZnKVSxh
kKcxeDXANfnxjR/jt2hyq7XC78I5kAXQCUPML4GmRInBcumvtR8gpiRU9L+ptCnUfObLeHv5ZjrE
LodxWwZgMqKe2prDg9L502dMssgKwLvD4k/5z7TjaXr4V1f6sgZJzg4T8tRiqylGTlMngYwCfcbc
zMXZ6OeoNjztmeVBHHAdhmndqRETw9SLFolfcNkg6pgSU1qANyYArKIEbiAR2Jsoopn+EWSgN1Ab
v5/fQj6HFDNux37ov5tfzjBPThy6HogK/D1YPYPdVCTRI986d9cBM4WPGc1UL+1UhfhR5CcYG9sd
/Pyki78/342au+fJrSmI59dpWnfqLs7v3xf6whb4aSp66LA6AxsjiDaP9ZYdcYrnxk5wc6MNSgdn
tmfQAzYxTR08gae4q34Gvag6u3djWHCNfB7rAttAXO2rIl15AxOMsJd9uWPmqyu2iy7nfzwlcj8L
2mX0sLRzd7Sm0WnXLYHioZra2jJrr9ygvXD7MPjwrVKcKeqllFfLTfBCaeXiF4uIMgbz4d4VdiV2
Q1HEIv7Y7TPNfkzcybKQ2uZGFpvjufRZaLwDMo5ypQV272Hp+wTgonnbMvDYrWac5MGdA1vHVrZm
QZYCM9GSdA/m+wdwjd5MHwMwpMC8pq/egark725zCLipwJFCziNrwZzet4BcqtfH98L+eQ6xVulK
zEMwZAuIAb13eOLvmrpoUSgiqXFT0pzLyLnlCE9x79p/Sp1XyFYjDH38F7AHe0JqxGp6UvmWpVXD
UWUE0o2O7qq1DPnxsGle/ikdthj4iF5+wNS2NTd9mp2w6zLEZBzUUfFG/fvw807oaPQ316epwg4Y
uIQnfBJErn9l6hjKDXfgKkAy8kEM3rbglKmGy2x08mA94DYuNpdcHe558qnieQyTKlIJmbrrEOsD
FukPy9uPJ/yd0lyMk2PhB6PexVQmVLFkL+6cuf2yBdUgYIdddOp/hu9WFxwxezn66vgs/haaSz6Z
nljeoGgIxW+4mfM23t1+eXKEoNfAeFKuYXdKlqoxyHBbV8MsAjrRSx2mAk3QOE47QewJoksLnY+7
DxLl5J4xj5DTCueGGvM6qzSmaGHybyyxLcsm5LNqQPKaxFvG/+Ch3jql0JuavzkDwWHyVIg9BKVm
Ye+ZT60WcHNOUwZJ9Ack/M+7C+jgINTXfyQLH3MPxk++74UQKGzVbIUru3JaV7ztAZW+a8hGgHj5
TRmVd6a10OWd6JeMxuuJQYEeKcVsJSmmh5qM/Jo/zKS/cBVUNZcUJwXJGXRyL7+qWW/0ArxjFgfv
+j3kbgnFwszrgHgTC9Cu9xP17CQ78j6JT4Hrk4fjXFhkRZRVrnLO/x97Lkoz4iVC6jTsTwC6jiHx
mTY7wS2AfCVpb5i0W3DpiXaoqY6xBfbZT4CH0tNxPvCvkX8eO4ggbIhH6xojVOSMnFRQA7c1NfoK
yxTesvGbUZjlo2wwVNUPbAFmcpfIM+bJRsbqxJIOYOjMeoQxTIcNPB1hTtki2B2Oqa7kQdKaPKOV
wlrh463X4DDsGH0GGl2oWeprc/GhBX7da3rebtmjNHR0Zl43+p4RCGXU2bqeD2pSIM1Su7YeroWt
hbR+7HKgfW33avxeWt3OxegRfcjldf6wnVXIyKZyN68HvINdHlEhWp6pg3rXns6MT8NiLEbeZTtz
yqLeNrTDYu/Ha/lZMk3pAB97L3rBh749F3Kv3qJpy+8RSszvx6g2zThNet0lqW0TiKMpqu0ZNBPI
OZcp5BOpB4MF4VoMYnFuSFeZ7sebg7Q/gkXjY6U6aoYVJtKvsVX28BrqH337cocOVYKCgrssD/tL
fGi854fyJKG0ZsXl12uNnJnJ/Y8twQviOmKrbbsQFXbJyWPHOlObN+Ixm1VROh1HLi3OKGVsF4lF
i15YS3f2QZdDaRElbEQlJR5udiKTnVij4bUSsvTT30cFYljB38sNZaW6kfAfW2Ho3BCSvldS/ymi
wOtjs4vSIpWLptK0h4EZqav6wwuIuUmO3ZuPecLB61DNYdUpoZ66TVMn8uOXUN9BFvcBbPY7ATAB
PXbuNLNFfNadHYaV/HKKqF9wVnzCAeX2hPFTPY0adQz3mFkB2RDrQNKJVqjhoG/JQVmn6cxYGdgL
zyLHHUwA4cr9rkbM/xJMdogitV+cPqX2eSEsegKEzb1wi3byjJ0DihPyuBe366QdM86BZd24syXU
I2sCuxUZAFAUSu6hgvmeaRKcpgV2KuJ3e0jf3G7DryzCXGvyciEvTWJmg87hSg1n1hl8ko8IhpsG
YoZfoYPXhQIURIfPNUlG0I+ALJAGQ/e9nH1ygONUBTsrw0bQAJycsn0UL4wAp9Fp2zHdFbELjubM
BhAtBgfTqsCS4I6AJzPQQrun8qnoAy9eg39xFBjorpQje2YrNqpkFKpXjKu6xs4ynfBl3rOMiqGY
QZ+hd4QrizFxKKNZQ8m0QPsKfgavWY0tlsgJAuSeoSvoNifgG+T30dYDTyQn+aSW7O5AAa9Tn1S5
useo5+Jk01+ISmTGHla3X/6ZIX1hKvGnkWnAsjL6RQsnE0VHBfWoO1zRbhQGFJgw/TOw6DFa/oxH
A6EP67ZkcTW7qdumlblkQ/BvwSIXuAzwIIN4pGfStC5gPbE5Xr02GiYrB3XFlNO6K9XgxlUCnM/E
WajNrFDf00XEyacY0LlhC+EYadE0cEOQTn7CdQj3RA7J2pGyBCWM2E74VysBis2r8vNFxc6y7NMa
AUnwAhER1+X84NUVYG+yh0cOjZYfdSHo7K+H1MLJmCJZsZUEUjkiqdEoL/cvA0L0pDwmMkg/Gdz0
o4Fdy6vrHu1Vk321DqEqFUjsZ0qXhjrWjcF8iqAyfgyBTI7TAp+AtVU6c/TqeRKKeDUdbnot5vA1
aL1KEWL8CR/th+NvNTG+ZHy7nAYcxELPhCpXKVfcerDwp3IEztAZgcMqsX8d9Z2NpK4BOArX/7qC
hLF5ybbvEKMuiS2wH/MWILWlVaZnEYuBnVTGkOA6JYSQX/exKRLtW937urXU//Im3TXdQzTrOst5
qOzO9A74iG0Ui9LxWF3Q3fuNHET7dryj2o1bnsfkrUHOM+MEp3KbP/GPz7na4QGlfYX7tGy5BqTQ
v40WPOnE3dau/zX/aE3Za/zx/Ib4b4jr+jgdTc8lPUFvJeSvI6hZu9hpK1U1y2uiXxPBfJwTyFMP
8LGqxXPBknlvIVbEcHQiZ3zU5s5hgs8VTOGFesEIvmq6voiXjl7vpExgNvFJcG6361aqMuwiTDu0
Sr0CC/BWUbRxpFgEw3Jta9ebwtN6NAnm1leCtMNEtEy6ijLjx3OsODBLLAvX1HwZ6pa0pchBgDqj
bZEwUIg/V0yD0cY9fuBcAAiPKCdWqoFd1OH+0y7ZO07ylT9yptxA130MIHIDnooYRAYbDkzOW4l/
8YQkl+pvqxriJVdF9HkQmLFEGDbGFAyf5V4cgexDSkWopwqvvM3k5frNfkwNPzM9gzJx8O75eogR
iARyP1pdt+Qf6QtOY6gF51740WLSkfglDEon2F8uw1Y2l6tYGpRjtMZZ6p1BIq5v/TR/1BIDRpln
w1rJPxOH1K/GyJaznIa8eDYXWQxcY/VmSeKNz4DbxgAxsDKy3Xcj7qah3mqKwOX0n4nf7eyU8Nff
kDqEgcnjAExIavxBy2ospliqyaMV4EjI94eC4S0qN2TRpcSnuKCKtGWOXEycUkHNXQNtEDMupFB9
JmzWdZF5zukXsvPUTYNQUdR72X//UurzEsl2E/B1KSkGtp+0ht5LPYKMoBwLU6+QZ73A/rhXYY1N
3+HDtLa+YIjcWJemHvCPwZaaaGXgSxjTVi0WI6WEfSzA398UTLb4uRjCMbT7mdQMHyBjZ9nh4GVp
9M6KobarhtcPvdAPx7pNWyA55uLGDiqSuuCiz5i2vdhi/UuoBcbBqHQP4yJUqb2/GkdKRapq66qz
TcwhfENxRGOpnI92emPsv/iPLy7RJWRvD3QhHc2YBNqsjNn5X4nnN+AQkZESRZUVFLII3SOzGL8J
+qzbZLW0STLpr7kYHCelIKAyBethM4NJBhdMavZ7r5jNgFvwUoWSM9b8eQO8dvpakwmcrzJtSj6r
WseEW3ImohfHYROq6tuuaB5gNxc/doDcRsV2wCt7hFULZScq5v28RPNnS5i3NI00ADIJAE9YbwDm
TyUc9lniEuQ6I21Iv5iSWEe7fJzVjB70wMBtQjZf8qBzsiJ41RXLwpnyBc7kQRfHnSHt0m7u2Kdt
c0fH8jC6ReIjb3LlYF9TkuhxPva3yzQYzFMJbmnGxF4kO6PH5dtEJcc8FszrWbYxBeLIxMpjSGLG
U+KLbczxazzOISMFs4IY7qw1FzCzKjOQ/Pz8i3pOFdOTh2mIWYCZlZ1Dct2spNNbKnc7CT88bnEL
MtNGC/SA1uZzWFZpXtilq0Lo6nGJAvcV5XU5auUewN4DEG1aQeyuqc/WdymeeKUgofpbf3u5qomN
golqjMVAxSy/8xn3jhBxDbYpcwC8TVQGO7kXF2APag2SYPeRXNGQx3qxKDTHhRZH0oqqpZzz38u5
OB+p4uOETJxEO7ebnqwNprEZxK9jMUPPYQWMAml67NuiWTa6aSVyHZFGOIqhfbApG4psgDGWR8NZ
swT6V9Hjmj+8FkPKhjksK4V0fdSo4xGDC34w0BGF3KRSY7iwOM7v4SsoFox2iEUA0ikrsZBZuvHo
y8JuNfZ0cNEEjDThpmJKd7K0Xh0zMpx9gC/rM+H9F6WZdMfBKSRZrevzQgZ++sagvDfgGjnUaAoF
CgRiYxyMDx6mxY9X/phIASpR/IFP0dIxhpAdQJUxLq/VG8m7x6EEF89BaixaP496c90uNcbwM0rn
V739FHLIHq3tjfQSN9hH2APgt1w7QFx9cTBWyZfhd6ILc6GmnWci2qnF4kmJjA+rvxU9ukTw4NKm
DFwuB/RnSysi15MxRUiMR9NhQLSREsTQpTjsWBooZ2nD5DuGXi+o+L7ZReMPgoOx2mrqqZRHStYe
ZXIJKCby5f7G4WF4bRgVR1JO9jxvCpOjZ/iLaEXqU16oS5aNdYnBgSzX7nUkrdr742qlKrTshcj8
uPgECbkF0wenTkO85tol56iHZMWi/po8TO/d3hjIBHj7U+lqX/G/dx5IDSXSmmcbMsj88kSNTfOC
nTOu9NS83+juNHTCDwiGNn7NieA96G3p6Ms5OfjyEpCCBaRcGGo0IJEc0WFE6zFoZHTWyFhSRfbx
OZiNHERFG2mqaeEFgaohEsIHo3dRxPL4BVAQ4Sw7iZMiGbZ9nJavfwmGAdkr4qTyc01wemAurOPu
70tQiqsjRgsXAq9U+x288R0J46mxW+PaBnlxiueK/bKCpquot7xO7SZ+lCbwK58uH05MyvVWCget
UBqnSQzHdNPHLvsXFIk2DYw5FUulTi9MVV9PqYKNXddqceCAebXgoiG+7k7YzFirUn2laoUZF18d
GEPw8yh5oqF52fSFFa4n6fZ75z/6ZhAEvQF7n2r9EfFuonn8nfDvSDYNoC+ceOBM4F9ZxFWeknhi
419L5M6/1IbKEjpmT4AR0VrWJivGkTMIhNxbqCHGOVUJfDyaCLbNGhBJLYdeXLy5KWvvSHoL5SeG
YtcZHCRnUNi45C868Jhe2cIneAl9pdk2+73bFL3JFoykhCXMbXJa+O9wIOK5wMUB46V6UuUhw4yX
wE3gN9QOg4GsGxUKeQhOG039jt5LkyldGxXMDtku703Rg6l97Sm+8bfEt4DkZDZB4AWPKMX8/Out
x/y1ppBe9ma4QU3j18IvEMU2Ngp/GZ8OhXR1f/VkSLqjGki/V5dQGUJVobA97o21PoKHIpEjVd3b
PXkNwY5nnclJ96eizLFhYDYkf9loAT7lQdCVwoLrT+liabNXzNC8XIWrTO2RTQu8MdjJUXRB5cak
I3w9GMuOZtn4ZAhqc6HzX5E49O/mbPWJteNgPhQma301Pn9IKMWj3iT+SBaKV6rjE3K/dSyjKmPd
PjwJpShdy/07clMQ7W+XLA1jwd2lIeaHXbTNEKpHqIAQELa4Pb7ufoTrpxZ/BRZ6XkOXka1MAWfV
roBIEasynXxXsMNUpfv0+BO3ap6QMjOSzQ4RgmQu5FCVoY2R8FeUPElfxckC0js3ONVtZTmiq3od
xoEQfMyse7V4vGfWt13LffgVB/158JsZLtW2GrkOqUyHxa/tThYMGZnK+ZfveLuQRQ5zwwEydS6u
tct6bO/IQ6z/l0F5LGMeIfrqMa/pSH9dfM0u/NPGn12RW/tvw0Snd45iQDp3xBtCsf2nMFL0OySL
zR1Bivl7F4T+bsLCB1oq4ovtfuHFvz6xoYZsr9a7JDnSbw5fkoGs6CXKv10hIeuDzj7HNTw7zcoN
3VtehGs9uQ5Uvjio5ZSo9dM3Gbbim2tOGUVZ7iME8SmgEjY9+Zy2Arhb7+RivBIQ/Hgj5L3s/3eA
Iqhi0uPXZHwvKow1WZpUIM19Wgg8kYgQSKC1ryDXZ6MyZL6QH796ZY0BFDJFLzcX0UM8ajr5ocm6
AaKTUjOTefyiLLtLYcT7E5RcfGRtVtWobom3cglZFZnnGhC8X0kvREzCe0MntphZi0/Wh5cydHw6
BDj4RZ7leT3FlPXd4S+oNwCo+GjlXMqrjGRrX1Dv609CDPwwy/3Knk41pT1qby992XdJGnWaMDdH
hNWCjZLLGmtoxL13tMISGmuvoZ5q0O/rmZEsfvfN2olmAJfLfIxdU6jmf+12uPdtE939OEgk47+e
7toqoCMQFegDi7rQF9VC8w23uUTLEjuXU3/VfRLTsBfUlKZXT6pBLY1bayUz5evEHp+hofOdkTwj
pfE4wyyV7q76E98VH9kz42Kv8IVBgbjYlJeMAApOd/ctlEg48eB7/cxqLYXMIKLHBDc15h5kYWBP
1gfItcKCbXxzKg/OowYwBh5atVsAhclIRnnb1/OsdoZQdbox1mvbTG09ToD73c03hq89sFMBwXLF
/kANr51v/zqkJTnCRp3N3/4EqRD8LpRFl2AAGYTk+e5MvFUmm4bm/u3WyzgVs7rMZtRqCxaYWUG+
mgBtPy7MCYpotR6yLZLoUvV6/NNOhjY7KIXnGUkG+OTBdUr8Ju1b5tTB79ZftSnZKZvZDM7VL9Qa
Mi4t9kHSdrTqkCoJfmmwygRqmy8Imipvgxr6otJJYdi1fndQxcJKri5gfSti85HohWoor6BUpMMd
PtG379Hmya43vvg3Hvesh1bdOBoA5FZO1zwewH7QlnA5T0HQu35/ftyVEemv9UUDhKMzumsRqWuY
DFGS+ha3yiauhAlj1JN0IJ9f8Q8zOikbKc+w3B4tkCOfH7EdCMmJ15gThHqLHdRge4QVw38+Ea8q
SC2S+tGYJSv5z9Bc6ZcEHnNOBh/oCYEqsvZazCYcrzxiIbQUR3TSI6QYEKc/pU+Ui9tBOuoyuuTD
sW8UGdFPZ7zr2GBlBfNMnc2KgiwyqF2Cd5/cPH6NyblCJw6T+n8zffzzzl4Zr3zpQBShtw3ydO8G
dHLW+r0Dt1Shw3k80hib0SsyztxOUG3ePKgMDhobT/CFZsfQLkO8zRyaVFMv0WHv8njXgWK/wlrz
n6qjecgiGqilFHEQeHKbV42RDEqyEeoP0SbcHL2CB0G/HFzYxb7FuXB26Hoq8AKF8ElkWVnNi8DP
j0FNfmNgJfTSQkZ8lLXOl93JiYxPUa8T0lrnt6U/VndLUUecme+FzEhX37d9AY65tgVFIr8aMepC
hhyFY9xVDLaDawR+XWQMzNALIyznr2a1xkJR0S0us0ZyN1Xu4iMckby1zfkOyz+UYBSBBK4s72RP
gwlCysIIO3h3zmU+sMcTgg37/XUaCqLWuyMoaxZGZMsBlu2RIpbz9smnlo1ma3NUG+UtIvs1U4Gv
1FOHR7xyS0lGYfN0ChuNQ2LOhlCxoo2psjx4L3dPP96XwGd4dRO8HjFI4BEMB6mrNWLOKo9Fd1Df
S5inD5goH961rjaRaW3qtH9/m/d41vDoY+R1l0JBJRawd5i69M3ZwsSW6sbIB1kpw5LNJXvYwyF5
jS5BDF4TOyiWayIyBhwgVvqoPb1zj3szr3YTu6yRM+IX4nPc/MS+7EwjmENU1HHYShOrL83BhV6X
rZA57KBindVeWLt6LuodkYZqP/KU6rbnzFcvN3ybUXg6NnTX117yyzZOsoX4iDVCxYnM0mv3kgPc
sbzfVLRp+uVyCtavX7mzpGcEW0M70JPcH5fGhr0+/FlDiAuefWC/BB6N8U0tVIEo85RIzWV+X8dT
nIcLqwFbbthujkLgLHVEoCQvIn7oeoQG6geT1Ka3i8sXatHfrZWnj76915Mw3Uhl8E+/mjxue2mQ
QBMUNwUwFRzh9dP+/Fj4wKUdqS+iMpXoPeTmTNbm4mchYSMsSBYN8PZD6qRZcC6G9SP1kEfzR9kT
qT3y/5n2qm4SCVc0qNcCuZfK/K+5HkL7eMy+s1qVshCIYVTohYbbgBp5fKPytgS+hBiK576vU4VZ
Tq/G2A1xlttALUjLSFYNQpZ8S/4jXDDWMDWovlogRlvaAdL2ir+0Gpk5Tpq+E5/oqiUr0n+raV27
EyN8WPVEnmr/pGBSvGjdVpfq4MgGSHtap+qDjb0hx7rT1fv/UIW7X9rrH6ZEVwHd4Vpt652QcWkn
GkGHS9G54VgY5nznLiD2x5dEvgQ1CIMd3Yh0o2M+UGsgebOd2+HaQdoh5HyrlIpucl/gwOkazIvj
P5T+tkLibykaJxQujurGs0Iui9cH/np7EgyVD1f/Re1CEJXojHa7+huG+c6xKbGBUr1uE/yTdkuJ
JGJealIAK1jVEEOmIiPX10b0SesTz64l3TwwJbqXGlJevycMTcJfDSxGIpExWp4UaWcQvUGCp5XY
91HWlu2QEj1BmWyQfzKldOA4ubP/ygAEuDtDhVh9seGLAttuBBZgQVBFgq/hxCtHS3qe1/F5H9Wn
xp0CeaKOO8NZZ60K0RWfWkkLRg3jrQTWLUD+QDVBSWH1JjW0HCCW2B0S3efbiKIylAR8X5QbDJCH
A9IQKvr2xUZSIg0c+ITY8INzcp1hY6cHEaOp6mXFTUiSCmOJzGwSJpVthjjwh3Tlwew38NBklRYw
ItHJBtvxrYa6k9vRHlTG8tI1InpmAP82YbnfFkBeGslrp9pWIGOqRhZvROf/CX4MxSpkeGFgspnH
U+LlnRRbF6kx8RmFqa6tXo9/jfUqR8ERkl9rmxgHWRUjxKrNYJtHrGCO6iS8csX3eqtFEcgOqRKV
q/+jtN8ZmXbM7JzZ83Yls/y79/TeqiFI5ZY7QDhprNbxd2TcGwZF6RIq/cawRbmJ2Usjq8SwSI/S
Df8lN1Qy26+XICu5h1xBSGlDHIkm913+8nLGtP7LU26P8Ucg8qy/EIOJdwguJXspe/1V+SbrMD3W
L/QgoQ8mrfuVQAV/Gyl0HebHf0YdEujzdmCnTo+dCGIvbJ0yMAVGKnWLXcfzYSe/uZD+7HP+qBv5
X76KB/1tr0ZhmY+iJP6ygiAHxGLVEF4xX+8L05nF6yYW+FPPbEs6vPzQIiZlrNHLZzv+11jLXWOr
amLxbrVxUhXBdlfPU4riUxqUafK4UpcPpD1iVMBz4RpZOCHyPctwpvMCRdGnF6TR2OcMmiiXPRDV
0iHfKdfECSSF7ZTIqjL7WlZZNSdWRbAMSowxU8iqYtrOmJXv891nKo8QPHJcTLHQfiAnC42msWOS
FU1VyogwSQ+OCQGfsh4Dmpr4jigt0MvrpfXJY2M82ev3YrbgyTrYrt3ZF6rFlHRZKTRaRn6VtyDg
krQIq9luy2PQmzforFx8FnRVj0PI7LvOibTMCT0xFM2oO0fznaG3LTURVgDec1vYSGk5/f8+KYsF
JGgUBHEHz16QfklTSKSt97Edh/JGjZXYPuhCOoCtZ/JQp5WvU3MaID61Npxf0HHAt8uCt69uTFwl
R4JW7Pdlg1DB9UQQZXt7IB/J98F6t6LLjT67bRr9Vr4p7I09En5killrLkzflbbBOQQT1xLEbAfv
9H+UBBklyJ+3dF/c51caIbIZAE2PazAXuQe5gNjfvfH2otYib8DdORbpI77lE5qrXDmpr4G+NfIr
VFXqdBCwDQl9YPyi4i610Z3/CkCPZlwx0C7pLvYcOPCuqa51lGXxpnUMOUy3s/uro9QoA+41KQQ5
przuV4HsRDBLTr8m7IzYUhV0qoff83pNRkFg/G8OTjUO+Dq4myasHyDdbjq2ZlVQXZQc6x0sLTIH
pkxiPgGBXE9VBF/ggOD1OZTUUkw3oVLoUgXYEzHnUPlJMrIMPBLDUxh5g5LPt2ge848FLm3X7R61
dXSfrMvcCt+ZwO5UkBVFUeeNu6OL8RVwErAXDPNvJhwq3gbj+sXaijN9tSWt4Lu0h4d6G4tvOw/e
V4a0z+8+vECcVOekNS5/nRB2qvBa+R1pZ6EBoBWdF1Zj2Mj7adE/0y+JVQv8P62HlhcIOmRxISxi
putVjch1BGejEBk39D2hUwAaL90tBSIXl4uDAI26rrGVr87M0kJ3lPziyCy5jlOeF0/adEd51+f7
AiBiyFlKFeykyeiGzKkShmve+241z9my9jp7quTWg7ozsbYMwtzJgjAneO36PDs5hNQHmB6HVw1J
82Jf7n/45HbKVhH9aH5RoxGs5tj6VyPdLRhvI+YIIqlQjlPTuA2crLFHbUazRKSegODpOwmcZkSl
REWMfKJnMbKJsq5gL6DeUg1vBSyu7iY7TNOzFWUmBtH+Q2guzHmpOJFhQqXge8f8efbnO/AU4x97
CV8ns6QKT/GQO2eCk8+ExmznKFQ6M5nZ0vDxjFcX09gtSr3jbruCzXi8idmOpW8shlTVpWNuaaWw
JLB764nkxZBYyDGdUjpMiDVZY934p30sa6lpeQ/xFCDmSlHQG9Mz7dYaZmr2C7dnWN1ErdOsjEF5
+jwM2Qjzi9+oVlnjsY/sAOtmpBaZ7+nPk2fZTlQ4GeXiELFYG0LFshSzFDzDNzNDOc456ifu4QpN
y4fQlwJ2oZ9Dvxd/hqAMOU4uV09qAHfubaIH029sJF1Scl71Z5qpmhSStEYi4LeW3OkPDolJt4xf
3Mce9HEfPPeu/CvR9haLTKjtxcCdgHO1Fq9lvqzNTF3yOZdLVhRsj7nlN8KgUBAJPr/LxKGit3Wy
BSGU3ub3jJ/RRWW7cnWM+lrx+sVnfrwQNzAadbJdMQm9fCF3DT6cthkrA83ScxRQBks3fyREiw9x
PqAviEqPqP425ADmfNXmRdKJTa8crnY421Nzd+oKLYBTb65rnMJjCeC1ACQ7kF8nzqjI2VJi6qIQ
Rp51w0+jEFsM3EXj1f0sOij00+bbAToaaK8T+fy7GoxxZ/HJmi0LowY2r8RMMpdKRDoADHphvqrv
3MOwwbUhlsID9wlxX9z31A/2ka6kSRwpnCwZNm6AFs3mXC6xwFqYAfGWCyjmVAtW2mpe0mg9BS/r
XI4dm9vDV6CN4RiC1BjyI+6vPAXMPGkKXbKvocG+f1ziE3Voap4P59k0FxkptSsYh9yX1cK+5FVw
jdPA0FAYf9+rqu50kf79ePABv73E+C1PtpO8iLhUP5NnYxZcA7tjmtv16Nz8BYxtiz3+OJbR75yf
vsyx1CDITAaxMJ6ELe2QBzdEoo/7Z+8EiR5BgZ6jd8kUHluy5Uw1uzuN2Z5aEar7LJWTb2HAm3hT
qWnG2TJ/UMbwcFJCl+vPgluOgxwXSk+DU4N9y+BLNBI4EvWJ/5Egz6x9dFUeraT+YZZBLSrhyyNJ
F+szBeaCQbjvmhIlqsPHowroomZkwgLh33fWWgghLO7M9j+e7L2PsjrfGPzOAU3fh263svb1rfnO
xch1/CmU8on7ON2zUyBp74yoD4odIsZFreL0mFApUt8rJboA/xItJkdjSV4JX/cMc+Tped4rJ67a
xrpuw/a4xHb9T8jJR3VXTvCuocgGa81D7zvIZegWd58FUBVYj3EDZAvl6g2x2AihvglWwAF2alKU
lR6SGgEEMM7b3nue4xQgivRS6RLYohy1cE51JE8H+ScU8yci+dQExJztk5Msn+3XARu3LGieqL6t
Zk2Puj9OGKd3bsDazC1hy8V38cBNRa2/0GHXP+P+T8ZIh1VBe2KCbsBC4LKz67mKMmKQNdCdHxoL
FFh5qeeeDvrtfHUhJpNuUtEe5Mn0or242JrU3Uv1Z1XJJaqR4Ieigtcllq/i1T86SNY31Vs7dQK8
wNlNLzJzaRETmLvxtj8EIGd6mPHN8RmSrz17q2KB+QWe42vTpNo3su0Z3dwR57l3b5vbhfGSGbFz
htiijMXfMA2hjbbGBk2ptm2qjvdKK4TZ0ee9VCNs+D2AsZETo8tyArrUESbPHoq7/wWUv6XrbxtH
tja20/7FUwra7GlzYY9BE+qJrUzjP6JipP/7myISKA6jK2q6ImDBW9Qf5sqwRth0OZwdB4zYU5a7
h8PnH6oN4tDh+RF8aGYFq17+5yg6QNQ8VAQpbYzj6+WiEvsDi8MwcVmqtTZSdBxm7B5f3/PDd/PY
mqZgTuZbVl+b5Yk1If9wi5JzMvIcxDLPoxUn69O8y1WIzYkEhvnU7BNpGisJPS0y9miwaVFnAWa+
Swe25uJPBH7pNpdCbaXITgUhsj8zBILG/SskSMY13N9LDuuEYiHHbwHGtDrlxjl9umirQ9en+YSG
OKzeudRTQk2Q9EglR8/P8IM+2QfPxMCO6ALYFTuNr3Jb8NNHWP3Tm7Lw2iVAcnMARTgoWYy7sfyZ
vmZrb9cmMF0UNdDVTH2N2+ge3siBlAoPtRRkcn3j1ymMf6VkvutlAKyC5XLDwOd0a9Z2Azlg/0Wm
r44nCEZw0IBAibt9noXEvEwXzUxN3b5U4fgtyC8hncJuL7fYirbX8qrjS+JUCYwMwhlY2LV4zKqB
WxGZ0WbykUwSYS5rjV3aGh6Jjt0e5nBWnDdUDFnqYnN5rI49SXb0q7oMg4hkwSjluWQRWF27r+wV
uZ4SI+UIeGIC8YysPuN1ez3qJtSuUw+Nqk32cww10E2nMd/Pb/VXMUGZaugkvj4vm+LCyIqwQiaC
24bTUDG3s7E7B+czylnbMDX4OBlGJtE54zDOYlVkD4hjcXXTw2N9Q+MvYaX48cSymh+aO0/apz25
6Zn/UURDV/spQNcal+SotrRvgAMeo1zR+nNRoA3nnyDmryA2wrRtVpW7JoDefAN9b1bX+TWNCW0a
SOGwrcWYQYv47mmQmYiA25NBcryH7XnqbJ0sUoVn/fyesd5uu0BQnwVZNBKa2wwYdZRmb4j0HivV
3itAdGo+mcbT5Q/C000PDccuGIHJWacFbUI+oBifP8Eocd8AWVALm29KlI7EsZjv13FT80Shr+xp
XE4d1qCSy+sXUMC+jMegkPTYo2uy6S7niDhlCFsM3y3O7sjq+oYsIjN1tn1o0YgvvNNOh3plDC2Q
/JZlkvyWQ7VewKkVE4Uv14e+S6YUqN6g9mV2DLUcj6c3zk3QX/VE85z1q/Tr6D8rBHM1hO3iC2iS
9i2tXvb3k6LnTUObzr0lO2q5QYHKa4xd3U9cmg5652WXd0TIAny4+D+uMUbibrDlO9yQoL+ntgIW
zGTkqwWq1ojc842VbhhG6BwVI+ibJybuzmKqxO7AHEzN6EFdDq8gofAwnx+dELo0Aq7WLFK4Jn4p
Ue8ZfYIODl/cy3lwXgkVePKqU8x3W5IcqUdEawxSL07m4Rb6BuQwUXhrUyXcV5g+5RvhgIB9EFWL
nfPKuhQ6Kr/fAdFye3ZjP6ECmQSuFQhWyMw7E8oDLd35rDhqiV5P/FSjKLlLjPietnby008gV8QT
FQXQXaSQu0a7aXPoYj++o1EFhEU+p5f+BikJ3vNAmLN2rKWg1YimmNsZ+IoLB/9MkF2a4at21VEH
ICc88dSft+ZZ2Pwv9UAicssGQJ/9UarTpM7SAp2bIQmpEeFP1HBeQ/VFEsdOdtXk/6eH9O/U8Jx5
iXpV8W2ggvfQfY2o4cDRk4OhmuAtp3DGPfBsGbEpxdd42vWyUTriRu42ow8TRv/A2rJQJ2soC6Ld
nItqAsgmf3alo9crBjB8FWun9sL1BU+YKe7NVAOIZrlOQg1P6ZsJyox9KqNFCovgDp8MaPnGknZ3
wdbvr1gQYHNGvqagQurDdeAIKqsdgIF40sjvIFifWmuyHnqaCyi0SIeVLrGjDNjioB8k9XfVX8Rz
uQNt41U9AaKsOrRNA0CEHvpNu+fNtxOlFFdPUwzFVdbw4bIndkppecU1POxyrNHoHNOZCf0CiXj1
oaanzUYtKYEbM/2OPyuYX20orwWn/1SqZ5wj6rP0polYOKxLUAdrVzh7PZen43qsgmFe4irae5Xw
Lkgmr/tsakSBmYeD/YqVvn83xejYXxW6eSpWFtDGe4BDt3JaOPp6S9E2wikvb26liC2EC9M790NF
j0qu8e/1Ae8iOrytvccgsIKzs26MwCU/0z1fL7vEhhoImn3snZV1EW0avLOC3oM5A48AUCa315rq
TCi60i7pgLr5sB0PRYfpLLowt13ARyBh5L3lsNUXMBWDn3M0PaWdAKLqRMvP6J6Aia0n6ROUU+FD
k/QkQc0F5FJuLUXE8RxAhyZOFyXPQ01qQvgFA4XjhBkgpRTDdi33IqGBxr15lzafzbETsP89yuHs
iTDhXM1BOejTic6t1ZvanD8KJxbN/Y4KM/xu5J0/ma6ad17/F4y4D4vl49LcAkHGKxS50bPrPfQ4
8kyJbDsTPyvWuHgaRIR/HzBCciJW2VaWKYXLE6fSEXJhUsjVn1iQSrF7b3Y0tXw4VaKmklCX7LhB
L/8bJfZEe+Q+1fKqSli45rfV+fNTn4wc0wRZnM4KTNzmW5zfRepWAB2/W0Itrpp0/9DJx7CvKcZl
0npYccnjkSn6TyVB+S5SOmR5VknZ4TRMYUglmiCfce4s24cDCkZMyMkKYyRQWgOX2jGPn7dG16EE
gO9xRsrW55tq2YfmhCKtTDV4U+alg1B88nGu/KpJP4KfK3ojJT8UXuy9PE6HdPswCnm4Hm9Jb8C3
WgiwV5oXPF6TIJuHx4vwIzk5I0UodcADAiFZ3qnUcZEg84IG74HjmuhaWAor990qCheOk3hIuCYm
mkNSzZVkfjowtTyOM9pw6WtXD9qc3dLQExBm3THFq1XNYguR8YENFzR/RY0jm13cY1WPaW1AXb0q
w8NEtJ+G8I0VgjLxyQLW6SOwdHEqY+AHOvcywN8+C0ADuBxLsZu9TZOI5Iyci+GIm6huho+auhXW
4zleBbCJJWgXItC1KmNkfqPpkFMHfi4nktL5ilD62IEc4eHTebB/71ks5DpAFGAka+qjnB5YbGyf
9XGig8MeP1Hdsm1uQxjZY2TQr0dRi4N4C9/iAe8gSHj6uq0t8Aavk0I+fb+zjaRoeGy13ZiAHAiH
gW3E0pTKp5q69u8Vqm+riF3FbhiAX7GfjjiUNC2raGW45ybtgswT5fMAKRAVx/Cu3ISJQwGMcXUl
Pqt15dGkrNEtiKh6TnIQDGrW3UNZNLyhHuWmmvpwYI9fYNoJmrBdN6cKNh+k2AYtmeE9ou6Rf5Om
7Jju5CFVFPUm5ZPZkJOXnxULP+rVMoTMLqAWmUKRVnXqrhwkHc6vvUxisP3JN0nLXY9gJsI2PkBV
G330ZvWrlKh2oohysmrkZu+sd4MpUVFj1yVt8Br0+1PbKTyLMmRe/I6G0O8QHYBYb581BbgDep6C
xsx6wNRmLZ23024XodxB5spw0s541Fv4rO8zos5Qm1h+CqdzLjvJqCswyilCQ61atFGvnMm+hEgm
tMxVFbKruJYA0C3GWEXd5ZsqeB2CYb7BVwo4zgKjf50kqegX+FNYjgEi2NDwQK69OuSHLryan/DA
MJFhUP2rLsEp5ZB5CQQwZhY6lCrKq2YMJvTqoA1K/FqxGPcT03wDorKyoJNSOggN5qnXcZryHb1x
Gl1Nbb3W+rx6wBwnaoqpRU6xExELmQ5W7PNAzQNx0B2eiCPjmj4+pWoUvH4ua7qXDdbEdDf2eHEq
N2qO8qYpjoGAoR4qPGprqj9DzT08TXtlbEFRBaEJMIIocRw7bGt9egdTKiEdu9y3BR5bA13g9MKl
7sAzXnP8D1Lo1T/y5aM44SaHHC3DeUx3dJgtMsY//iv6qXkOjtCgziVwGX2+KRvByLGwFLjRnKhl
klxjxCgv9eY+d7yyl95INoqKNQvzGq1XBm10yq6OYFDXGje2HkO+d2jaxWZIVDbhU/13Yg8Qaxi0
yvnmuhrpEhuNnFUrbY24lMlCPDNAEjv7JQC2+JM1vpz+uaTqA+5XNx8CLwLL1OB2PmGcTBwvXkOD
99PngNLjkbhFLoEjU5ziooZX4+uSV1ytCbCHA3fGClAhe34bRk/c9WZGLi+Prj7DCFJRPxIhl9PH
U7qKzpIZ2YeKFZk6RncrIq3CEsOJx3cVVUvj43dk7z1WPDQV4cKJ2+7VrrQ/PwHAJj0UUeLVWVeo
0oNGKkVb4Qy0hh5L6qcWXuQ0stUMTAdyIfjN9B+04APQ3FssJ8VcVVLq64hWYJSetEaBIm8g0jpb
P0v84DxRvR4q+s+6IelwFLIp1awhZ/ez0IjxGRBzKqNfwEM+Rdzlv4bhHO97nRUaSjN3ZFlnl0c6
A10j59jtqdKqkZPOsvWCNZC5AlCC35vgBKQlyXiid+1Y3ThB531RHTY8mTzTenavzCzVlB2/uqno
TH/Byq4Cmrc9ptmp5WMHGg9B/h0jYstRg8BtMwJPLDtlB1KpCUzTpUsgsRLa2daRRNSVmhhdQRr/
YsoAfwiJuzY5HuPyz6B8kshwH99gdRWAA/xlLrxigyIpLJTb/ec00zm+wdn3e2iiaCzMNogY1olp
/RNVhT+OULqFZUf90c/R4zEHWk6Z2jXqhaL0ZMG8ToEhQv8NrFCoc1T3RyrmzaqdomH7co0/a8zd
utwB4rxZWaNWC2sVkPtZUqTROnqfAp7UL3NhhdITfn69fhZESDPSSmIHStf7bOyUUVVH28sCmhYY
PqPA1pZi8VcfMRTUtY6C/wApqxf7c5Td6icrKNRtVf7uQ5Zt2PcNWctZVnCcTstLY9hW3OHf4tt6
fEW+qYrrD4u+v/G880cVPtLah+5NoEByl7X3SiuFTtX0jgu6Bqu7cSmlbnoUuGPWcpgY4pq9Mmon
wo0g6MtLWG2GhUyayPV4VElDQxXgf3+XcQpw3q2Nk3O+hzaft+OQEo3ntNG5j9ruuALegWUge85i
gt4WwS7wBlcM4Jb5tftz6Saw3UbjGuvVbo0fS/WFO4i/v/LcyuF1gsPUU+Uge2jluUmpgf6JHP2Y
LUeBngy6I96rDsgHzdemAxLnak9WvpWWuUl4G347f2EG3xmPxGjgc0Ely6UmUnZ9SjOBSdb25d61
ZFFEkkysft5aoL6NXP0BXjlwhSnmQeztrCJZoQgKDkOyBlxl4hExW1p60LPMXrtpKYvIXUPz6CUx
PtPNjNC16cZNdPvb6ab2/VXMnKjkZvAPH5IDK5W718eDJoLio+1fHEXhu74kUKp8LJOUsNtnmfJz
6+XLbeYBRGbVvqZ+gdgKn+xK7ReHuwVg5pkIxfjzbFwNe4eChH8EOpbCEpBH3kF0Hn44nM79EX3I
GKQkuaFeFfAX4M84JVtdb7tOCkIHNXP4kfpKCTpnkOL64Xuf4BcQwe54bnStTKHrh1biPG+CQm8Q
OHW6thz+z+pe+x79WSYd3SlYlWloUhSqrEHF/JYVM7rgNmeWiHypNsx3U5y2taetzpd1uM4Na75r
Hi/G91IHgIX0ZlFm/mz78lwb4mBJ1zw9hjkH2523ZMGNZK4hbvYKSVmXOtQssRugezmUKBcbDijG
kqasVxItwP8zCRTuEWK7HIjLM+dBpdvM87LTrXdhO8lTmdrmJitErpoDUruF5nrPM9UEWVGLIhEq
J3ILrcHHG8mTfhriTfZJ41buiDt141qqS8EINLahWFuOQwHMbQsSs2ym7+z71cU8mOhvUlcxHZMW
j1+8IDgaRW0VLlvRSMjqc2Jm1v5etsXNUXQnfTzC6q7yHWDgJCzrlXapIr1n4T8Wr57MLgXsv89y
ZJB4hUEniUHFSCgaGonGsktqKzGdXp9PohvT8HHzXIFIYALUMdcqoZyaeW10FNaFXBuUCgg14y7V
GU89tbKNdtcNrLXQdLe+jfqcyLQv1UB8v/PX38oQfr3I022qqxOphCqMXy4btwwYspIzWmxiLeyN
midv9P5AMjwaKhFJ7SxL4uDek3qTyFhgLMeiXQZDAt6l24kuAA72MHTw90E0e2ikrEkKXg2iQq59
yZ8ghtpJQz8WCNsiPkYvR4tHHPi7K2gQi5fTIQcEkyP3o3CKNgUkssqjl9JbG8qpoueQxGN6CWXY
Fc7Bprz698Hd1l2CjftrnkEpTeep6CaEshZhrni1F4rl3/4snPGP0JrJ0frX59XZWX7JguSGAT4h
R35P5bQjeZ6kNzPOlECGxc2L0vi83lCfVQe7+Fb79g3malkgLIjokNNpyiZnq/R+zo9j4n9+EatV
EEiJfuqV99gIzlrglAihv5h8aHYqqM0R2G3Spkkm/M8LrAD3K6MbccKqum5v5n8/Ff1LwMhPYekH
6FjP4iURO1SJOlf9Z9gVD38HlKFs3F69m4VKySIJkDaoXltllLzZzKdlt8HzuGohcfRZFuP2oX1J
h3HQVDajJsFwPKqoetaFGwReE8AVUTzFBsbcOXRSDSWT5qzHCpgGxErqZ9FZVCJnwbrJwlmQMBZX
4yC34T4ORAlfQ8YMDV1N36UQc5ACJi32MdhJ0a1QUtLhMZV0MqQYQM4TQ2MHjeWyqkGpv8Q4dJbY
o35tAA2aTR1shZtG4R5FC/dvUy+OlYoHj6kDq/c9e/q2HLzNlebGJp+WS8VMzTvi+z6y7fSkQvcT
d/mwxbgA2DEui3GwHHFDwM6AmHSoYdaLlV8WIrWfuwaOvz87wT+nIIDWiB7ZEXCNuxMh2eOgVg4V
nKkk9Ghzql5GEGGI0cP90rZhgUfXcwSf00oerCvtRWUU1Eh49vzG3xpA3zL+2QP38DkP09z+8rEO
hG3Uo5rT6oyHqWVf1899IrVGG9pi0LRSpl0CbnwzNI7RplLutE8/7lWp9Nx7EJopBaJ0VeM/wERH
GuIsZrhrzZkNi16sRdTTfts3vIihVddMf3OpofuZBksFe8dh/DC+G60oSi54vFNG6BFhNDuAgWJ0
+MmSraWeVOTW12qXiFt0ZRJ6OfY41yNwY9U21rm1yGjitOJJvHR1mAafFOmWFSPj2KAehmhicKBb
QMgkQGnCrX6/7bmrJ/hReHS2fjIoiPhUKb5UIk/1W4spMBNkLZxGpvNS2AogbuDBM/DLUAaQ0doE
M5so0/xruH/4v1SXmWIaPrsjjlcXG1hWdYFeVD/RViAayje9zWeNZ3QMeefZr3B1GLaXwGntpUAy
2Wf7DSEYKdA6ytE2M63eay6R2R5RKnU0CkCgK8655t1pJTJjNagy5gL0gHDgZqNVS5ep/NI9kuzt
JFd6hrck7le5T1D9ifgU4RPcpeHaDgqIWKI9ZX96DS2HBAUeJUSt9pl9AOhUM/BsOyHjSy/sclT7
Qeu9bfnkq9XxErQ+B98aGRMsSq02rVeiAMBuPnNpGavU9W5SuGOAyDqku3b00o5xJQrutcrkvXqD
kmJujRo5BVOZvMyZt7UPXPQDvhDChWtwyg5xvyjAzNHW46cPmSb5McRVO2HAYAYqb8G9QrcjdzfR
Rsuzz8UayE94Gznj8OJWOo5wB7s3xvK2EzVQ9eKYfQ+ZdsR0JNx8l8BZWV4AUz8sl9ARAVHrD9S+
MB7uIMST5r7M2x39TzpvCsxS3zV//d+EBuBylg8QrgnDWJMbQ2l5kIzGb90RbEHSQJsRw3kJPIYt
e++/ympDwr8mk22GYYS4MEXoohdXMp23J3vKGbhvNQTDTsUHJcL+mzuHMe2oD65j3MD7pDOzdzn9
oEpYG6AZJ6GinnUy3j1YyMa3L1WDbGPHohTWVmeHI9hs4yQXCcHfR3eOszUxK7tabtBKT8NRh3dB
PqUum0ApGtaVj7VYvEPc9gHkjsnf756T0MAHIdz7rCN03jidIIRb9hu4K1wQF/jZEACK2vfp5wxI
bdBojwc+CParetIVcro0tMJx9bXwVp+c0eahC8mY1EfP3GakXvOA01m32Y5pxuqs5urmcjR8JuMb
0boiePYXXfyqUo5kYwEWib/xhOSq3ZZWfrxB7oTAdw+FpBmyEvZb432BCvvc0AE3jdY0YzAdVu7v
zel3PxCCorimFSQ3lCQ1MDj/K1Gp0sIUv60tHBqEUY2V4G3o2qGc81r8P9pv/5z/Xzhs2IIgpeWr
BWYpbc0hIJ7T1e3ru5wsMIlzNvKn3+eH6dvtAmM+dgCOJo+XpGQFfKYbHCSWtMwuaUFIr8gstlVN
Vb2sE0AasAllhFEgvX0HpYeO7cDkyeW+Q4rYJ86cnTl1je6L6VNds5o0WdfawhkfX4p3/p1OrBh6
WGY8q3QjgoFsZDRj1xHID4pbF1sK5l51LnAXdvwdI9GrlCQP8iaa/5aDYd/ZN19hJQVr+3CVkjFG
OpIt4SgD3x1o+V9ds5V7laf1Jk9qlJTDwjAl0YA1f03l7HGYIxQbslHtjUVCKzkQIHfalrydLRro
iT6/VZTFN1Q8gq03bkxhIHg/kXZHujqR51RVI0JoJ9h0HKxwlqbYs0y2z0oRpVLBAq05V+z3iO0Q
kfyEqfDcHqEwx6ASlo8SHZSbGyvxsSXxAWJIAhYKs6O3MxtXIx2morpnFiwQnghA0+G43JkHyn+q
v/e21jvHTDxHjyYaxEGphlTwHVdloSyhMlOxvVWrVM3tunrONTXDwNQv4jtkKjp1zwzS5EY40ylP
scimxnNsuWmqaAGhFXqvr5kH1G2fLuDqzDf8EVhopupmCB0ebrXjgXHZ5CkIKWycGZ9NiWifOUBb
x5vMKF7Bl2ZR/HYFl+m2H7AISbNQBuf7ZY+BLKVfvza82IAK5PZfqbezq7ivzZMNxM95ANmgxkjl
9L3mB6pNYHv4X4zwJ3wXSIQYwVJ8XxlGMQNQlYRyOpNH4PHft9qWx1SMETAPQjOsiTRtLTwfz2lG
v29cDuq+7yRE1NHDGcmX7AxK+aW441d0xn8zFlOgDrjXj1usOB2lTCXeMqrq/WbVGV/d5cJHV+Ej
r50G1KlOnBO9a6lT/sW7ggYfHlvMzpIK1lzraH3E6/d7pSJK05vzYOBcbC53Qrx/xaIN2OKdc9oR
cEiJPq0YUrxloNa9BrcgxYhRhOfCaa99413+GzQi5lLsg2g1Dtk8mBsvQGwoH4DV9qar3jo87piA
OgBscLzaGUJSwARwhFCkW+F8OuxOdm/oDo92ib/YYi9knYFRvZxS4cBuGcJcmYwOsJSahattcWO7
xyN1i+Exst0cCOlNmjQ36CJhslQUSv8G+gPmiVt4N4/15RDpeTBDUufw76GPPOzFcueUrFDalWKB
FHdJoHhgVwHT/YZLon7EFgJKzdex2GIoJnYYk15tDJ+HFIvuGqGbzkUJtItsC/m2ejAiYfW0rkd4
gd+1H9e4+5krbACPWdbl87rysBtdpFffNuF6RRFZQtH1EOx1/uSD/tJbPWPfjoIiFZz1Fbpf+q7u
xkId3ZGcx103ctsqv+/D/p5dBwBFUo771LDExhzVrlfcx0dtVUQR2bnTXcC3+BIapEZ0GIeiry/n
LwskX02aFWTiqNb93Rq5fk8dXvCDpzc9WqCZYv/p8z9GQhO9aaeBA/xWc895Eom3+s7EXAh5yhPy
opLp8Jv65H0ATUaGtyXA6j9hW6qOtF6THRZp7bdmuDaeOeZjLOT5qlyMnLESxC4dvQjqiHw2p3ML
YXclDFyIWJJbsbnyWcW4WqE2nCJQ2GEP86JimuZybShZ0J8vbTiE4jxDbzLbRFYknbTAfbXKPsBs
Vef2R0oev78RY/hRxV2HMj97gtB9UHcPpWiXRJe4ZuZwnEUzGZDJYojWg+x5eiu36BHLZgploEA2
Y2SvDrTGI0FN6KiJe/kJ4LZ6pRqW1pi+GazTD049HmIKTqRNFzHt2/5sbtqUbwJdSYrFL0RN8urU
8c9Lg2bPpnVY1n4OzXXUX6FQUzVfK0OapbgeJ7tkhs7sk8OrlmWrhVWxodQpEiQeoZXoPzPdKH7w
nvI09rrOLzQc0+C1alE9vBXq97ypZxZ87qS95JpGdOODPP7b1CAy15rT9zxKPo5/l17uqOYNQWM3
NycRRaFfi++yrWw/6+LuJqbKm6fp/TXnBK90XPsI7cZ9a4kIrLrE9JHd9ZKdOLhAD8O+vxbyrHAy
MlCQVXrm/MvGwzK0MxHzgpkHOFy0CaBC4dIM5b70PIHdYPrdao0dgwTZljax6rz8khldH7nuqecS
No1gqnln4D+Lkr4p6LpXGEOABHwS9dXELtRjZXSGFry1w9e9V2zRLCWDktsx+UtcHgyTIVdTr8jF
xDTBfxcbFwCKzeZwIwDZTi5p+4E9thJ9oufOwpbunOrr7vZxJT9w3GkEx/AyNA7bRqg7oJGjlW5J
eyDc1pjgXtlNR38EHKI1uRm/KpgqPzlYAnPdI4x4gN89u/O+nAQS3LMdRzM5Z3zsVKRkjSBKGfFz
wASfm5Js+VETg1dRFykpHZHRTtoHM4qKceaZ85BcphAYDwW0prMAjA+R/fU8DuH23S//toA9pW+/
38Qy3ihczeHrS635a0lsD0WvF0h5gajB/vqkfnNgKAnyCSm5kZnhVA8uwTImmRJCLV4HCfRzx201
40/9k9gQ0qDwZhxyjEqm+ZZRd8wzFu07Y02T5ed1tBllFY6EBskUtiuLOmPsL6xw8jI21Lg0rig7
9LgrOPGoloHd1f8pxi9tHZxziW8Z7zMxOFV8wBWrLvROybSMFNf3oGwapH2Fg0J49JNHVrX/dMxN
DwRuq2LRrfodH395B1XNxZR+8qYZnfNnpowOSm1sON/oJyuQl0afS8dMGzCq2h+czaVRXxyQR355
YDEQt5alA+r2A+MNBwU0mwZDer7PkK1u+sf/S2wMM8x/Mky2QVtg5PXpEk9atUsN+co/YvrK10Jx
wjgxwUHgz1hPY2YjVZ3Xm/PEaUwbtH2P03Qs+MD//EWeFx1mclwwMQHhBxGPiAAZYd49ClTkkbLX
NQiVON10Jw+8zvcjsHz+gYr4fK3fK+yAtNMErssXMG9Nbiqbzphu/4GjIJWIyvKKvfBzMtIxru1O
1dH4eITTY4W6Vq8iG6NM6vLnuFw1Os1l8miI00vszB2M3a+8ca/hiiSAlhZjyK8J/1OMvNO+e6nD
TL5TbNrZ06T3cl+waypFOpoNP8W5Tso5U0UdjW+Kpp7amNGH7uQy4Bm72BvknVW6FtAFnEgYMGQD
FxajZjSITybvFcb6AYcv7oGk1AG7HWrv+TVh/izhqePGmxparbF7hYnWP+X4I19ZlcU/GtA9m1iY
Ep3jqsXM6e7xuaAgfi1+LpDHXenLgiE1s438SJ8NcaT/NHyFmdAbICdrDpEUysWDDmBgF++0cfY5
hCUO/qyNuaLwCIZ1lOhDABZQguC9CiR606ciE1kv2r+HCfAwv5fIEUXwkbI0siqHVPsxAhw4p54a
qmmH58ipbdtZNK5IoO5+hxJKQjqIcZ/3Xlv3AEsscFBiGMIF4yMYxEpCySSceKndbm5rtpMT8QuA
frQaLVPqIQzEt9Tfww56I90q0mXBKKDvkzd8C7p3c3nqEmcK6czlGic6J0UBC0G28xJKn0ROghUz
PXl0SY7REeRG8PUmc/gzlfaY69FjbamIiEBPGor9sQ0xovLe1ljjxMJQ1WpSS9QPysvvtSEuQnkj
umKqynoivXhNNUtHyBDCFqABrKR6L/DAzu7+5ow2KavKa+M2ZxGBNkIHBvYfk63uM1mAnfCh6Ql+
YZ1myEmrMz9m4cgI4QJQGI8r+r0jzWXMHslPh/CrAvAYu9Fwc4OOXh3PeeaZxZRIKp/bGqfkFskV
neUmzM8A3oBXdEAXuo/2os9hrj+Q8NtwspDgjhh3xslCcRWRZQHr00C18pqBq6TOaXMm60VtBqtw
RRzDe5RIFPmaaCUwcjY72i862gdENj/KkTB+l3IxZSEtN3wcrRKFYbSazd+GfUAOIbjmIS5oVAzB
1O/uH5mVEAPB6xBbaj73SWg1UGih7YfhkMrPVDBS5KAQEJQRt7hgEq9rzIJhhQpiYEA3EC8fPduZ
tQ3Ct3onpsDyBY61hvSBw3n0lsJQdqrJogJ/iXRx0uzugWvDP9PfBkV6l7xm3E2PchkYclihNi4e
yMhxYAY27LKaJNZPPFcZAX5LPS9nilJxepRnoZmOwqnckR1cXpUhEMBp+hezExNd6hT9Rd5pI+st
pGFpv+6B3bCBuBfZOFx7J15A+aO3QufwPgPUSo8VCgjL8Stq4YZnGCOx9KHXT3BFx1BHqdZ37Qyw
JnEsPVlMX37HPRS4+5HlPejhClBBRr3jDU4Y+rDjVXWXwp8Ac9JIw5dtV19eB5JY+tiuNSpuJMII
93KZy+NWg4cSyXVL7tc7e47D+OCd27isBque74aiE34CoBjwuq8eVAA9cY15VRsVcRHEMvOMiGaS
YWFtkl76uhL5DjP8HNvn0/JbZfzze/N1+gZOVENX/7EY59tlaztKXxboP7zNQujRJVI2pb8OjEXX
3R5Lkn+QIhgMQBevKU3SN7DF8vCL+3/dk0XnoJ6P5JtJnTVnN9iMyYA1gEwvVgzssxyN5qmOhMTX
QkEVlh/NuGmnbOI6O9+AGeKQnn5PKpnEg9ZAXocy6DAjTFXXa0XUNffUKVpIuPePioKOPSnzgxBS
VMn5CrCUxhTxdW6V/mxzufBdldNiogomp+yMPClPqxnCH2Pp5VI7Udje//LFFJLdMF8YtXn4EASa
X5k8IoxbmYXPhgFBthDSBcm7R3patoetpan2cHK7IKtUpBzPYk+HB5Iq+mvRbcAXdzB73EwCoHUX
IdbzIgzsTz2bpou/Q1ZlPonQDgs+Oz3yAZHr3pOyWVivXjcBO23XDPz1cSBMSpTI7VEmKUvXCEpc
lSq9t7cDsOq+rOc+ZEXanITscGV4/v7Xy6mPzYH/Rg1XDC7dhS6jGyESyEGODGx/QlkbZUIo3dSd
7vF9TmyKOp/oCmCtT1hBs960kOY8N6WNrIj3VLNdk9ksNdb1HVNSrLkccGQ0tygP2h05rCJypT0z
3+rpcFvx8Hz060zKLBJ0XXV+SYRVNRFKz63RGSM2hX4HVJ29xkcTSBh/FKe+2HhofuWL8/32NM2F
5MyE/TrGHsq+dBAFybEVxNCtooZ0U/1TGK0xCinVFgFvSDgDCJW9f/v2zeIDWUeXQ7PMAZsXtoNw
180cdrN9aE6QSW1MWeqMYspcpE3eA+RXSEi1C80NZKogn7cxTmciO0AzSRJDa9wl4wTwfIugWH65
df9YWbY+Rrq+BgULpBtg/NtQuqRZy0cj8Bmx+csRr/DJBfFM1oe3Pi6GsLLFrTlAIsGU8kWFkgsj
Wjkibs2IgspR31FZiR6hJpP7UN9jhlN8DoD4Z6JP9Ttr/W7FQWUB6ZzPl/gwF6QDp+jwF+KHWDKA
0yqAgO3xbtxeRlbTfyIUgmvBeQBKXScLPvYumJQHwZTz6brqA5srOeI8jfSho5W+d/cXTgndVAnG
RvagOGLc1gpdhP/V75jlw45YHkdUWkllNxXtksWNuKJkBmOMrv+g/VgoLcwtmEELY/+8sq0RZ9KI
CxY19pcdGZgnNS0UM5+qQhdySrDFSYOCakDYijLxO54RgiJTdi8LJPV1sotVa+A+o19+SiCEZ2t/
RZESLX3MhzoouN20OnuPaq+ZThY9mXCv5FBNA9VUl7GzLBCy1Xp+gKpvY3Jik5hf07db/tDnJKsN
KjiA1YtJoBg7wRmNLlOgWSjg/EMCoJ/9aMUBtC4Z4VjNDKS9qYU1L4p0wrFDvk6NvcQleGUUW628
sDEN++zS/l+I0bTlX01BLfU4h/ebYUVMkGn+FudqDzDIdYNGPl9JNPH4MZ63IXt03aclnl0gpz1W
ohLTt3xvZcWpAAhNAy5NDs9HKkTz2qoSNyboSCvofTco/LMnx2e8abnMCF2wT5vpb8pvcDu91iwM
eWZqEgIC1VhX1wgPVbMXAv0w0RocOwNWTcG5EP+vLEu68OXYnR9J41ZCWvBep4VscVMWy7NMjKAv
SnM6A+KgcS3ID++4tU9P2aEX1PykTr71bQWT3QmeTt/oUycM2l3ftopiGWbG7tXdtmVyafHF9MDk
py2U+cYjVSX+aIBuiYvvirYNngj6Bc7p5a8hbV2HSW46z6U/zxoEgYtV5JafBtwe2GVwbg+NBm8/
UHefAlQ7mMa1DhDNkqNGq65gQ1kCUYdd3RBNxeDqZihFrVWCx2nz1gol54Ynz89shBPpkJlW0dTt
fSnaEqFEvUiWF8dwi7xH8XpvBGw3qE5MknlWoTx17z/q0uUtv68nhzyfW5OVLD6bC4P31QXUEy7T
QSr3pvTWd3VIc/ltmGMIziaUsKONJu4LfwVJxJYxtPaFYfF56mEzTtU0Bu5wK9cdlW8ugQ5r4Cj0
pmiKBGGf2gzqXH30l2COMWYeTVgLp4lM6dQU+nJe2OhlZgAXyPrjBIHCpGE/gbSPWrC1ebm7ySTB
JbbVx0QLPCdliD8hwkp3vbC0q3Pp85IDFrklPfNQS3HWBbDuQI7BxJuHdMngbcuDyS/tb/MIdOah
XjpIF+v+OC8KbKOSopbHyqjMzdJDqgOHd/e9HfC9p9b/2QmAFeXiHb1Q5HbZGh7aluZ12YiUZzq8
cy8SCIbHAnNq1qaGHWw/2ACZJE+7EG0ohUj/q/vMMiIuypuHVsnASyhA3JGVXL1urHalVRioASSQ
3EhRlyMZ+6rTbpShvXQWBzbS1zbQZydtrrUlqNzB9k53CKmyoU0Mbdufkj7241zyjksasPWsFfk9
AXOvmYPWFY++h2/2QsgWCj52F4/V08V97xT+pJPhZ/6UoEdasPZmK8jahTCjirVXZ7ht0A0qb53D
qCpxoI0wdTh9OV2oKoPJ1Lr8nt2NTkhI4v8+zsuElbVsNYw9HisRR00E6n4d/+VqOic3VtGmk02+
C2KZk5vucYCaDbWeD5Brb18wPFg59AOsaJscN9z0kz9dJBjj3r4U8U8one3SHeyvNq49MAoek/nF
dV5xmGCqNjJzlGrDXAV0GFvmXPgqAnuVylDISs4Iz2NMVJpntr7ZnCRA4WTU5ZaD716jXzw2nYAp
RYrW0lKuaUL6+jOQAyy21CAbrlqrlVwPbsvBbvRjENZk1Cjqolxv/uxQC0AS2Z/kW7oNIFBmbi7+
j4eSFqpkpAhKp3Iewii/6SZTDM70HPjlUSZcdamkG50jTTtOvgOU8U8PuT2TIrGf1OE2oGhog8Fl
4IPsxnYoXTrDSqgLd1bdXGhlvLSnwJIad1PUJOHyB3hf3Du8hlGGsQjVs5TtVvBrqVss8Nl2srJh
4RlVs6gqw0we7R46xyUxcllyuog7AVoPrz3RT5fCDlO2tRP+3EviMoJrpop4NUAUWRFMuNUoTHuN
z1ceGLBy27srdmTaaI46veN8AS0TN4W9Cb3L2p8e7QaflqSsgUVgJdQEWa2JKg0OyFxulCX8GKHA
tbkdzE7gYUjhQLvWn5kxUMcWf9MqImYlLja8VqNfuw9jXv2s4WEUNPohZdS4s4Giz9ArjDzhl6zO
oC6vkbl6bFCWnxAXsc8PgM5RaRVUyNKK1GuAVj4hoSa86YvNjBuFag53qibu4G9v3X10wTGWVcK+
LlXioYWMFiJpz2ON6KOyXlNMzHMjVM/+Y4w+Kt4tlDCofd9wvN+zCW0skjc+Qy99XNWxRbSh4AVz
jqF681dtimp35uLcrKjTuy9xs454ox5hPwtQmDrbIIO2xkoywrboEwn87zquxhmOAYTtSH1a+vY6
3lG5DMzL4qbUvuAVzupce+2+53nr0NXidzIvcu/YwK80uBI4x5F79462+nHBEC+S74CTEVuXY4Nj
S5bM113GFGbplp+wp9jRULxbmayMlwqfPUnphoWrwMBSWZLrInHAaSUADuB5BsTEj1K6A574+E9M
XJ6NbQHPRLMGbxbhXkIGSNAXzZmOYMVQYfYkMvaowmA5/WfybPrVZRuqzB+buN/MASkKFuaT+slK
M+hzaKqziXvZAvief5onouvw9N+D67UnpuSyMfiKb8cA9Ool7SUI8/z6aqPGW4aw3tX4+ZuaKQVT
/+S16H+n+rnXKt09IewT+pku+ead86RgThUMcEQoZ9SUjff5rdzcXH7/S3LRYyAT71ErjMpS6jL2
ER57mklOp6NO8WgmXorgoZkqupzcH4dWWRPGQojsVg6zhQUqnckxqUG6SFYTOYg4ZKW2gts4cawl
7PNHn0Nxkr4yOJmGDOZXd/3huLNegtEWf+jvBfyALrdhkIB6WuDI/r+v3B2x59X2/ZAaBi3dYy8F
iQGfZ0A6n6rm76g/fUVixwlbVvJhrJi99W2+HNDzuCJooU/0T0FYIdBIxwK9ypyBuM8OFTSJaNsH
FE5UrTjXo1j8FNLcxweqfMXFbXvOY+4rTDrYMwzjp2Y5PQWN1MwjTS+e9vwwbCB7b5yREK8FnNO1
B1C2fvYFyVdMQBIXwFE6VcNbUu+Bs+ehlwipBpqvQ3cjs3qT126wQYwWONXVhTR15maRX9pTe0uZ
Ft0SSjlAPIJb+KbxaPrOps9Kfioh2GUr81c+C5p39tpno3LLd5piWdRVv0lTIIwHXF2UR1KVWTJL
fxnjncqlbG83DCMrIcCqC9OFKAOX8G3cC6Hs42nZggRYhRFDGaB4vE30qm2ioOt2J9DYNn8gcG7S
5kRFuOcrZsZ6UqQlfvdxG3Ey9fz9PdTm5AMhzPVp6lnsmGmwJ7YM4u+dYhBZHdgW8jZg6dbgM1kw
y+WCsUAdgpX6ZL5qziaQ0nKIRxy8pI6FPtV6v5nP5EjP4xDAdiu33ZzQV7YaZF7eariYUgeItVc7
7aPLsRVUiENYaSYD8MWK3+uLUDeW9gdcqDKMdzSRHfbbYOSs9ToIMyVXZgKPWFGvMC0xXqLk05YT
hl8ycXBFFBNdv1C9z7csknHlIgh3IbtntERgp6juGoTBMjvOohM0koHFBNSTVi0h/qKMv3Xw0yss
DtBToQ8JF7ZB28p/67NZqZj5adz3qdhBoQQiTx7M6MNPyHfjbKTFFmtKLaXj1ne6d7qzLpLUChH2
39nSFdc6UkpRV1OJhq/mLOFr6FLMOapsk84LhfcDpeOvpr1rT5oj4FkI87O0ecUdf/X4Pat+/h91
ugJ9u6qE/pIvnZKg0JqfrcPDOxmO/5McGzyIqU6bmxi7PCNvXkNyhOmMK3MgfC23Kzec/qzMWJKV
+d1/B7tAxru3Ge1Mt2jhtb3JDMPlgOaiLs6BsuuozlybvRjlSJqCCh4lY5WlwbLfjPoTnAA3ogFf
jY/TAfwqmP/Jge6wk4ei3hoNfcOEYHpDABnaz+pXTTSmIJeKwElGWddpsUtfanm/qfQHwtfZNijp
kxkuoldIOKJNSwkRrMKsaStNN33zOCi7O0jLcxlhPN+PuarbPq4eSovAhxHiZCDbKqLiLNr2IC4e
iOB+BmG1FgDCKiOvRjhB37S7bmqUP7ZL+F1W40s0gR+UDxJpw/x3nZAEMPSs7qUXrdmuvk53PdQp
/n9ILZzkMx05aJnjAMu0GH7BkbfTC0Q6e/jOkY62BhG9V87+fi83L+eGxSiBLBWwPsAnN97mE14U
nl1GRUYFKhxErGq4wSEJBx3XKe02JH1ykrzGLt8plJ2W1cDHZ40514yQrwPLrU87PZUt5NIDbdDB
uSalpSHQmaQ6dOAnJSg3vSnVMBzTURS05+Y38UdTSieENn1yzHwRxTyvElwMJ/lk7O6rORMDSqnj
kDOps0s6ApUNiAHPIy5ByWWJa7ZG1s6zDK9ht1SeTtC8MFu25GzWw6IwyP733JKfzezXnxqaB9X6
KA6l4pSW8JzQS3+pGe7HWXn3Gz1aIF/t2dD/KIFqFgYZC7eRP+l9Jic/2w0B8KoclS5HVrDTJ05Q
nZiEpDY+NA/4eDmDt/lKsnNE2ptZtuCXguD6A5k2/HN1XH6xYia9rq6h8nB9hZ1xzdOcutL23UCC
I5jIPYbK0KSjJVVvSwbkb9Za10q6rUxMsr1tLL2pVcesCzF809mOPpQG4KUpEN7nIeGABlM6iVSo
EWWbAwVxf1thEPpGw5N8ZBt8/vVXptU0f5sGT6J1JMYO+xJQbalh87MHApzI/sY6iyPHSxRmNxOF
P48/M4M1QKGlQ2fsUYgaB8CCSOkWQ8XL66utwxm6bxBw4yjkUD5wAWQViX/+I3VcD/tZc2zfj0IV
l6V+PXR6WRdRIXcvrrSjhc7zACS3HYw85seKl6CucfvIPK2/8aTE/ylZ2niIJve4N3I8eeYS2UTh
QoxUM2jh4471PEnTBP299rUljOjWK6eyzmtJHI1LHUuUQiuBY7FcBb2oglKnAKq7KfgpUPLaLRWg
xXhiQX82Gt3Akkpa1Xud6KjIULHUeFB7FRp3BApBYeV2TZ1mCItl5ntjrklVxIo0mZ3W58cALr1t
A+rQjPTEaqKp9tGXKsVIDkkNKLFeNQ20+yzq5SLYDSk9EWa1fl6liih44otrGhbV0OtpoEpb0XOO
sZtX3+naEt3dx9GrSE66hvqwP23g0KHsY9H4har3bafecjqCUyrpufGKnanhGVPeepzZFjwSKHp8
8ok/Oql15PwGvCVHFJoHleWdFeZUd7CjEg/cyuZGlfxzn1CmE0BCG1Ih2fW7WfXQORLiA49Rb7e3
O5+TW/q2ORg1RyN9uXIN94Bwjg9j3SQNDW9Tcr67lhrrpPfJ5LzeiM1MXNrYalICfrOR2yyKg/mI
a8cR7RQnZcFCecHTWfZDTS4q6T7YGvNNoTxt5Nkhv8I9LSotTth7Z+c/NzSbaq7LCICrSFRu8Ctr
z1P+kUf/C6GGw5kMSZhEuWFEEdv0pgTYXNpZlJdIBQJjNBplbYVgOt1GjmYulRJUe3wUVUfYgnb4
ri4uA+QzZ+Hdth0axOKJrOlXNKbnZtIYFmEUtPC85Mj9ApgjrtFj0SGn2CPcl2rLoFULiL11LHht
Nvw8BTjL/4ravpuPCoeR0sfZP5aLPrJvdN1GYlVOboPmAj3gdauQvBZ5IY8POzi/35+z3FOgV0d2
vY3rUvTqWxwBclSkxBGf8UgY9raZ/PFOS7WPR+wpv2npAIml4YyXRq08/x4Irs2PvJE3WXKSeDF5
Ldftx57gY3N+FfArSljy5djt2t/lMiobrzwQAD5ZRIHc4IBaNizDJ3aHSMWdilo7wDy8qskYsquo
VnajYC5nzH9SsE2djdvlkvG0qReIQR8B1XIXuW5kyAGweD3hyr1VI2MhMA4U4cWFnsSahBa6jd2n
p+UItUbwfYQ8Y5MFFumGuDA+xPdOTfTyjRMbE0aB5Pb6y8xHj7g6J8zi+EgRHkpg11eEaTlAOtnL
bdXQa4gMUUfedLDnRsGYFnlgIhXLjugdH7PLKByXYOOBpEKiLPa0lSQVihcIP1XyHrEXOWUFoYbj
3f61IT2TzW3ThtjCL0ZCbShG+0eCdvU0RBmqnkR4aBOquGimMejIO5H4Qw7SMWRU6Ljh4goumV4e
kjYN+5OpNtcMZQM/6NydPA1a24OOt94/XWHiDFccyFPFKGqXIxzrl0knEk5+gye6ShVJlgo7ig0T
VMlYeR08RKeVX4bDg3cFsdNkNvla0A0t4WhNQZHcIqixnRbzb6KhHJlAxHe1eCr3fV7TDo887OIE
6SFJ1Uw+UQseBEsHs5c4srn9xzo7FgaXSuhn+x7hAIteT2yH92pQOY2HZHy+4Kca/GWUPs+ucJmM
3r1lx4rEf9F+rZKcnm6RO0QNWIHzriOZyub8UgbAYI+lxow3Da5QcVYl7QGwpFnTtA0eUSeMNlOu
JNbfwMtwei511i3Fc4LKRgix0V1hsLSIAEX1T/7meUAHM3fnjKfufSk31YiBK/QF8rH9NsK6wm2r
1IAyzBjORQqaYKT1LC/Q5agljZpPG8H7+hkN5jxouOWKzhkRacRVBRKNrh2xBS8h9mtfDXnodAPz
jkHZZHyrKru4YaAjmI+8vu5Z778G4fEVvz/8UkPc9ODZeOavihihDoXpyOUccbfMz/BIXMViLULm
/rYnuhqx5dmCKbvu9Un61R466PMbsb6hT+u6E6VDvWwGni2TFXki3yMQviHZVlu36ILgQmGjzzEK
vtTW9Rlef+4aAIDFd0hPUGg1ViVW6PKFs5THopbCLncBmuMMyZ98rbOH3xP2preJrSnR3SBCRKvj
dyqvtNHB3Dm4AQjEAzLTR4uUh7j8yyxZAQuXhOKSUg6ppQdHQCt6UAW+FB8sFBjDs5FPkrtZ6nc2
IWgbNdbivuHUR75T6xgXvPV3hvSHdM8jT0evh7dYR1d1kmWAPvpOen+OWbkRJYmqwMnVqj/fsr0H
sre+5hbqNKxzV3r3J0gKhItbPo9cNeFzBlZs4jkNl1ws/icYy+HzeF/qseeXyX25zuugqg4LutaS
MPZauUQgdgUCNly6Eq6tGjuJ4XHuSU1wB49mJm96BHWX1Il2V0T5pttSOfXYWP6jYRqLupYzCE9q
aZ7LoO0RUDSdZ/D6dRhvG4gh7XmRBV+FJNvmTpGNIueXUKAl7tRHiaSBCuHEZL7+YaMe4yY6ZqEO
5zv1Dh1OZVT8T3ozrJf3qzxAbvpHoQaY4kgsl5eKNXi0p6nz50VCJO2fV0IxyU2vYbaxyoLb40ds
LRHKx4GMIJymH1L2AFWT78CUz8FNdp4WXXKM+JHr8vFvPil11r/0hmoP2G4wcQJrABfHtcHMEt0d
5/xcN1/0jSWHlzYVvO+pWXEW6qAKGjCjiyAfm4o225t9BYRmV6XO5xdB97iPJgmFNK2tfn2yOwc9
BDcinILLBUPwkmV6O1iFoUnzF/fibzcjsf7+mfGDvvKf+zUqdgUcl4O+ZbNLhvcdiSoZQD5fr7C+
5okEX9+du4ejHKqK6hwbWNAW7uS4fPV8c3vKF0z/fFe/MeRZvkuaYayKgrytBA29vqdHQv0r0PAk
LGz1c/jdhXuzWAQntrRyoRes7CI/tM/zdqDYDiDhXQbWgr5Yjv04I+mfxwtQf06u/j1jtN/EV8se
6zxx8jgyBKp5bq3vDUZCdLIy19JY/wukvX5Eway7m7BwiDhbAFlnNm0P8fsct9LtebIwjE+KqCz3
YW8PZDOIu3y9es/ilOBcUUWlyhoGPXvRbhBH802DjixJTCO0xKpUnZUz+7qmpPa7+xFGUZ4x7XSM
LC3WmRyx1qhdG12kMPHGBhrNYxEOH0dE2UT8VjRMKfoQXLDDlGu6ey6j15AzunpIQ0nZd9v8zFyx
acPTvaLLeA5ZZxHKo79M2tRjjCbOUkUrGi7W8si+urrorjN2yy1dVNWD/G9K9hm2Z+zZuvJBocM7
b6BBcu7zDj1kMiAI1hb9ve/kijtljjpncdDuQJRUsLt7k57/SF29+CjDW3J/MZA/Z395JUyLZtSS
feFsx+Qmi+UCPl5gfsmDiFE1BN0YOtIILNYfF2e01OgKFshOQrTiG0quurb0Ce7Vu/9jWZv0hu6N
VqUnt1+bSXb9lUuAVm+Lu7+DZuCuGvlqHw8xossM23Ti46DhW7l8b59v7XfPpqpldYxbTWHw+mxU
+wTd2lC4Ma2h2BbSLiy6zRx02imkyaNWFSnrokbKh/B3TjHNpPyqlHyqPwIoVk3Drltm6+aAy1xH
xYrVTO1IVMcTw2j9V//fi3y4khSGea1OOu2TKu6Zul/PrP8WGOvy1qNWh/8z1Xt9As28yGl3wCOb
0RY4Ql0kFUl7+Wrt8d4RQX8J4SIE2gA8YGr3ZvC+pcP095kuCw6xLK9YUhvvqhzkYps21rtzb45i
FI6yMYDmyhpvLqfQ6AiISwrSTyqq0eA0ftUnpqqZpAnktWGTm9MthSYIoThZYjOgffy28/gEADeH
RWpDd1dCLaQakEb3irf/g/aGfAEWR4V1eyRu6SXDbqVlQ4arvjNSusJXkJX4sE1I+xA46ylfrQHv
GgJKXQe/REsi23Jq/OREdZwg0Xwa3/Y+7t/wmRt+OV1okbP/Ayf7EGrkTQg2xtPUMcBqnG9c6iIw
SyrtMNh/p+J47T8sXhSY9hnNC37CeQOwUriMq6/ajtHQf/eeBuxOS4Ubouit6kdLyixFPi1jkasz
i7L5n76iQnjLBsrLimmnxMcQH7tV6aEeLE9nSQo8EWVee6560f+TMdt48UMmuid6BrsBpHkCqCW4
Vk+JUQvei7IaXcanwzV1RDVYjK3wYdokzSa5t8L0/hX41GWW3hqjkJi66yluN7r0GiOO9B8ewstX
F5fAMxhk3+ayVfuiYxJz0G7nno8f01cUaxxGAPsgHBNDsGjzkUaf0Pu/+CP/haE0W9pslnpfUSJN
KuWIB44k5f8Vb8LA/ARfSMqtQOUdyxIOduzrVyglSz23jIjJP4TIk/sUG5fksi+vUBgJGao6KZeW
ChYUIVp+BVrkb5vGpUZ51j9B6loacJsQCvyBbKR1R9Hec1MGfBGsErqeuai+Y+PhCN48pmhhy3As
LTNarq3noN8Et2enwtDTnWGcKNf1b4HlX50c4Jef1fXPCGG31iZeb0stmO0AcbaZVpL3uVxmb7nn
66RuICtC3xGTIqMGcS86wvma3kcRHw9qxpMxF/9UFtRjc69JNZj9BFmVABZ86R7ptGOdYPHXbUsr
4OUO35t1EsyG9AQX8f5Y30KRfbzzMUUACzsNnD2EX8WugPNrq5rcmCxuJOsfbXvzP1kHPRXUIhND
mPGWWWTcBGJXJJedgMm2832FDsKeJoV0Uy9gtA+PXxK/K4/x8ia1WPN2VGIsFQ6Q6C/cfAI4Fv8R
NrH5qk16aQbjcYoqfidYpFJ1PZu0JZKnWz9dfX3UHViGf/lvl8cv5py5dHJ62mzl6XeqpcP7cp8l
VgcCGSyDZaBS8IDlosPdaVO9abisjwpK20D5Yrl5bFIhBT+t7UWA1dt0ly3dzJ6+v3qSlHEf+NHt
mo4VVY9RUWwyjc3j3XMTKak23Ou0q+htTzvuR6xNArSN6RVxJBVLgIIgkAt4D+VE5uDa8TYoOvNs
6VFof/dRs9TRgdDtft5rqVzFAkY8vfCgPKjAURU1EUWmvYElZgMpnr+WnWY6sDeEj0iylmErioOp
sw4TzJiotcrUqK0cWvmhtl9NV2LO6jJNaMU6GRiGHuldd0mxDeW6QqPMNNz5ZoU1bBEOSaxsDFaU
hggn/DC/L7Nois+7/pEVNGvHSisX5Ym2NgBbVAUZKzB1gqzRnaEyernGox6b2qu+eJaFPjqK2+wr
W6XK9oH+b50Uy8O7PiaxZn2mfOrer/7gMVhMuC0d4ekcGBRoRG7BYdwZsanYll0IUfdI5snWijCq
LYX+QeaDFHWrrJ0MTRbTPbEF6GMKYW3fsnntQDKYTlXGUeaVb4DbMGVv68341vXoyG1AKaUzsB0y
2/OxG2ItkxSyj5jenIRebQ/3QVzyG/1SvuvkTstnFse/3PjlOGhkrMreAeRbrjcgGTd/WUBO5dS7
nKwXJnGJn5iIuD0DFH5iCSWw4i68+4d2LgApqUmt7wjLuhpHU8Ld2hpzIGKuIab77zfRxxj9EIaF
16UCl6GyXg/zcY6GcR1tzWBtKoPd20/ytB0w7j0UzOq8H5NoLEqmaTE9Ab5gNL5c0dupLNDympG/
WNgMUiApvXsTZxm6252F9wOFhTmWBIC6pZQQX/FZwEYlPEJsbCxYwFng8Q7Uq95MiKUf3T1quI9d
yBqL6bqYt8egs/i+yy9yYiiEIq4qSbE9JyKloRQk+Sp4I+QV8AGE2BwWluYVdtKTJE9tw0Iio4JX
3niE+8gPu6wrgxwfWBdIx6sNqMEvdURTOYEuoXSUP73nxV5AetHOcvwI9jSkzAoA7oCPVVMGPLBD
w8tplTtL/QwesLL4GVMAHg9lpXjMWxThuSjDJ5F/9+xKhA8UcqbtTcfODoJWdAXxSCWMZeY1jYAC
A99NumYWyC2qIdbYKcZZWkCA/XlrMso+5tBXAgdbnGSmGW6Tf0Igg2tUhPbC4AfbvbBx/yF9309S
2uPjgPE/IhodNXhmTCx/kGgXsOsq/H2mCYj9ofDVWqAENSXz0LOoOtiwT2rm8XmZqYKOVjZuwrr2
hfx98sN78p5qeVmUBITQ2oGzT32fKmuOP2ffsBQjRYnpGcjV5R9VUkFnWn4qT0bLQUKIJTGD4OwS
B2LKQ8E74UdzgyS/Kv8/vRRPzs6dzvqI0N+9RQH9gnZKjcy/QN8gQNuAsQY15mIKq+//bGqBvDV6
p522VEx2f4tFwJpxVckxxvJC6ran7tfRweodd5T3PD9mfipejr5V3tQxZkJeMNgmS6/4/Nq7mUGY
6dostNW2EqfjtFZP+dIitkJmrtorqj3+wA5LWeAcz0xaTx2bwV5ZozJxNEgJm3tKp7kGAwQIanbY
IPwCrajlH1RrRcGj0GJ4gBZvR+wyc++pwBxyfJNA6Vr87VepO+fHuK/8uUwwAXixfuNsEblelZXp
0bNKOJDIttzOu+uhu48IWdbG2oKODMCir3SNywLSs2wU+WvqLvGO6es+pXF4p5cI+43d2/Cpxx2/
XeMs2DPnjqBwwk1K54Zd5GL7tWhl7xDK4OeEtrB+B2vfJLqr5gAK+hCgmB2zhkJ/fSnJ5ubBEogG
6WpcfKsIXjI49XL6iLFVUxxpp1P2G/y87Vr5MCfx4436TQKC0aAAToA8zXlZWqil5A21oBXa2Ix8
Woze61FMN53vamCtJDbGXmD3CfmDljp/D9AQ3mcP++JYZDA9gFlA3DmB07/1lT+E2bsDDuho4BGT
2tXSeaU7/YPNPGePRU0ejzMfvZFKTLvyKOTxwY02juQCg2Oddlng8QlUZhSTYcCQdIfoNwl1dE02
iMSaCwR2mY2nU77I4w+Gz7bSBPtXEFUk1xwJOAZSPfUQjyXDlTE3/tIG/yRKkfWyaUaauQipcapz
T5iR7bN0oGcWLq9Mc1DoV/ZKhrpgPgDTJSO96QmMkeiIChDIL7j1bDJzHaFgQ3y5pEZlBVBTqoJs
oKR1DFuQ2/e9c5EPbDB4foNARTfOuND44hi9wyCrnvqqafiLRJpaxHH9HFxkXBImkEKBlvVUSUqO
VElrVEs+9CCuYlJ9eVu7IAalH+uE6HonZW/10cUzYquwHmKaUOmR3wXam+CIyC8Z45o0dRdAW+3s
CMr09C+u7zUYsGw62ym/vCsZ+cd6ilw7sYvOKUpzD261GEFJ8Wco6Oh3UtS3VEB9HG7y43PMatn5
+eIY1cKki2JHCPfOBb0FYHUdLXjpS80GEs/3grQmSMu+npo8c6LL5aou0GyJov2VnFZwvdxJK/N1
4T96mKfLxO5UrlYkJ4NG+JqbzXJ6+f4Nm8o+orlSvVWUHkcvVLwfIyGOM5EsJaQ609HNqRG0ejyN
eZZNu7cQ88PP24jpxPYYV/K24zeBv6MT5dDgMiOWHVl7eyTjLSq+gbhMifd0XS1XYpgTvlDc/Ycy
QtRIHI6lhQ+s00T4i3pWlnOfcegIB7DxZnvXFdI70P1dVAiIndgGe4DZwwuAA2lYLy++GzaonEMm
PBS+kUre4bqWFOnGflAtk8lA/jIlNJXFh/pUpiUB9iG8HZ7P/6AHqw8bRl6k8e1IXbp8jecuPIio
jXl7vUn8VaCPKRpKXoKFI+PPzID1coPPSwfXftcDmkkcz7FerkHkazhteCsEp9eoXQZ7QnF6dsS5
4T5mEPX9HQR9ovyKjAV85exfDv+kD5VN83TB0ukiwKLd2/n/hLaC8ztZiUuR+LuYOvN16QWrEFn9
pW9gWuWw14eCi2nCFRgSxt3xsXyT5W4pDj5XGpHZyyET6quvf4TLs8rVJEdagBwb1DbC3NvYZDKv
022bgWi1CovNjYD9muoAZAcC6Vwk1mT9j5qbc4CV9aR0hAIL/BdWnDWdkP3nnoGX36RkgDiDfXcJ
URpwSS2dhQRZUxZMkooTl6fa8S8EmUT/nEhfTNDx02rgvfJK5hZuOpV1KOqgYSwvPsgh0WNFsYrw
pLevAmIIHXrUFtM0B0ElCjofqXRpPMjzr6QD3JQSJfbcPuftv/GQJR8Em5uOj83yrvbh6BVx9gA2
W/ey1Qq3rGYCP4KPHjm7POR+FgNeR5upEuScv9jijpJxqRdQr2GrJ4492AmI0+VPUoG/ejwjggx1
TigdnktwI270bkyrYeTbL1Eop2KPh5FEi9vLH/N4krIfCOJwXVi8JzeNJvRJm8bnjccPMqtsbmrZ
KAkkPKSV9IjsO01o5dlfCN91HduLFSxkVPawVZ4G8qFENT0xmkm/Luxl4E3NYeVO84Fq9BKUv/1S
yCnMRcrS+i3s9jzh30jTjK1NXbq+B+uR1AHChIl+dZz9ocq9QEyWLlPfTsDIHjn/gZ5ezbEelmsK
PZ+hObTSVaPs41qWs9BBRqSES8MJDcxqBt+TkNWJA0YfnOM9GGZU9g5wHp3ak/by1htLeeIvHNRD
47XkoNq2aa1c4qGsDLzMQh1qXeCsvLncU+zjS/RUD60HlpgHiQIsLRWBYxBQ2xNenKI2Y11ToIUO
N8ws/2LHZc7jwMFRtsrBddi2uuu+Av/4iKatndb7TEYZLLv7iY0EJ3rrJJ10QAeNHAOWOzOewama
sA0J3osPqESGt1cFwuYCx+s1dXd4YAW1so0MJieGGeZNhaDhyPsD6asYzXsVpbvg5CjxTqgpqkxY
6ANufdefqeFenGE0T5TyyKqOi6z2YRlPv0IYxoBxi9duOXWXGyONIb5r2YHpt05MhFj2whi+hf0R
QrYJGj+oaBk9/9SW/I90mfQ7cqim61v6om6rzxWzqEzq4PKpQaAX5xUEPU0iVjnbJdkdnu+tCKT6
GzcEKn07upuTEpcezw1roSt1GBdpVETDmuzPogrbGLoiNQTmLFPHAg1wcQGyYr4qqkfWDw0yS2Yb
TPX30IN1B33Pw4TBnwfLZ9eYHyEjK1hncrZeulRXLxfQZplU3KPE2egExD2ULOle5E0opJZoDhKw
g7W2MLGhx5TV/sIJUzTZY4Lahh0rBmi+3IVEV2WFFcQQHHIAfcYGtCxj6O+SOKfb0HEbHpjMMQo4
e+B3194t56DjPnXtH9MKnKmpnvXnPec9uA2wQFc2XH7UAm+lubOCAXs3WTQzw5z2I6Nq7mrpxPjq
0PO1YcJyBvLq/mFESBUrqQ8uoIsO5nWWCedM8Jf/bBo71XnSCdR0LweWOR265XqucBlN0Dia+pXT
5/7S0JQkw0JxOnJHpkuZYr1oFEYHgEA857WAgJRl5rTGsCNL5yufdpxJh7gRPGByXnbBG27eziso
ix/1BDz4IMYBHaZc7UoHtfxLLoMHOTfEnl9TCzT8f9zSzdI4WVypYJjQcP1Vne5BJ6PqjYMKLlXM
QAgrdwIbW+27QPBDBtMt7EQCAA6J4i4uYZJXW+2A1bt5S5CS7xRnPrMTIvoAFrDd/QHiGVl+F768
VpF1E2PK3nOXNh57fUJZ5QqpnDVYiNyIYZkuz0fGm8ynkvkdqL1wfwGyLIqIevDEEH9lgekUeCVA
SoVDYJjltwsAY5uU3dYGhJGUU+ClD03pfv2OXnLXo7EXQbFM6nuBsUatlOep27AKdkT3rys1A1n0
dbmdrab+1nekUQ8mDMXVM4/guu2P5/JH1siZqT3WkTlStrL3YfM8R8BA08Dj9mjviGKHfZHC/tYA
qcvTz0pU/buIObuB1t6/JYHvk/BocesH2UFnvAqjI2b1dzTTb5yOGNqzATSY6szi8qRl3ZcSm2dI
iWQiMPZ1n967mwpfl6Q8tQTzWfYNDkJZbROQC8iklPrdCaLYVn5CeHcu2OQjTggHRWLth42OY0Tq
Q8YKG4d3642IexXQUnxxjFcQiYdbKN5EZ3lpOqqobkxW3ees9mO8YNsh5y3hk0s9S+7cTRTTNo/0
NlpUg3xvFy1uH8uw0FTM+aK3ggqoQNjLp9CZevhiDodaocoXgA1oom19NMxcb08eoR+CvSVsJKRl
s0vP+vnmokbt6YE9Qb9YQcPwWASjP5AS67vhnpG1OCdqIRr/nf+Iso3SXYUdLsmpVy5RmKlFTlGq
HMyXGSOPIeAB9sByfnLGWWAXVvh0HTGE5uhtGLF1uk4u2xvhtdt8Ij+rmj6KKfX1bAA7yC/yAtWR
V+l3wT7FJfDv3YaxcBfy29LYulILJ4DlQVQulpp+pEogR30F5yZjtwfvfaqyZuw3SBivzCdR2enu
J97UD17Pv/PH312YYj5lqgR0mljddFTE+kKl3ev2WfnSoF4sEKNvVKhJZR7Es0bEWJjW6iXGtHgz
9l40T3qz/8iIocoywwvoClrk75ybiQry22nEgDcIlkSRQZqBuYiWI8A2Er/gwQDinzsAjNKeY+Cx
UbCehiQfeyVtUcZP+11hlO1dMee9VNpjfVHe8lVONzY21/AL+WlGJo9spheRLq3Sbh/VI4mGQMzL
6elN3hplQmpvV+JkMQSaeAFxG6FY15YN4IGBBvCDAqf8KGYFG0Ie/oOMb9lAEV9/MPEiHStnMpmy
bWArtyMC7ZH0g3vwtaIoa5DJDsMR0+TV+jsKuUqAbCML3yxRuRU1a7K9bOQylKq5JaJ2VvM0EMxu
8gnVoBl0Rw28e/ocBEuk1pJYKSYyy0GO/rcoWJEylIP7nR5wOm+II2qMfN0J14zD+N3VSTVpbKP+
HTgrMt0+NUfoS647uDhKULx+6BXNt2CrQ4ziMHzlJLwD4hXljtfC5pM0giVPLj7mR7Git+HzW3vi
LTJoHwzYt1hmbP0U/9eLAZkF2JQ6AwdGn/LUZlG+6duVduTEgfhsKW+waNDAIsBVizOtgwY8Vcr5
FbVjj2mKYCGGvMX2+6CzLtogrgBAjFQpzl//Tl0gG5kY70F74COjrq+pR9jm+dJp2D4p8fmOaxOg
hwQtluecabuQVs5PfggJ7ZBwKg4+thXKuD3sDZEAA0X2fmr2N9AR3jZvSS6Iawh1tnoY3Zo6dAgW
6GPajJEHXTP29NoLaQad+OR5p403BP7f7Fvc4T0ImM890/JmdHD9wAEuqH3EV0f6NRMf4dMGjSTM
dO9fXUgo2koVfpHA9mIF4dvW+e2zrCoMSMiNowzFFrQkY1tPYAofeXXr7YAZedEIgjzaZ6EI+0ze
W11Z/KSEj2UQJtL2+LkwBlUOcFStDPzBjFMz47gxpApns7nw/+VI0Bssugf8/J/jOR1OcIttqvib
EnIGoCmDXA/EUOQcg7ATS7OHS7t4ZQq423XQOK9HG+NRl9BjgFL6azBg925P6hmtgfRtjE6Ag+aI
P0d2UvuyMA5oaE4/Rre6nmDW7OSf5KEZQmxDmOhCY6MG8MdCEfUSy2EmExY1AQWe6Z4+lxd0sLaF
tqu/BUUI52e4Zo5c4fO/0OSA9MdGuQfFPziR5AXHzv5zVWT6zLlqogiFtXp+zkhuuRPjQc0WZF7+
X1PpzgDFcif4hSTOmYPUw1HaJyqZwAQkJgQd6z74NMf4dxldyw8vRSbvulU9+puS/BNycOZTONnj
/yYI6SDFUCKZuJbVXWbX1cVZDA+y4AUwHNxscgTlMXsUwwU7MB134Zzw34Jtf84CxW71sCcyfdE/
vATQN0j871EBZcuT99qVYx3x1LWC5KbCtrsAIc3mNmi7YK5IWI4gOQXEkVb9n0fNWXmj3sZX33Bf
GyKkEztulkmf9WPlf46N5FM/yk6qlx7BUGzcLPqqp1byYG1K7oQ6JPLtcoxcipFG2Ip9bytxZKev
NTZ2F5BibdajzPdEas8kVTTwhYdq/i3Wl8UNPPCFMiKsjvDzR1xaKGCohcrkWztkftjTqk8uh3DP
FPxdIJajE9a2+c92Gs07m9x7fbEkn73F8e9ONvgFr0dq5gRsj96KWjb+Ak4KlKb8CzLqHTrjKN3a
X66JIHgTXZQ0K8zvXKKutEi/VTpfG/hWiVL0ctFP1x+gLHFTNXKdJqMFN8hWTwiYwaYq5HzHXsQ2
4+SmiBYByvr89OiDE61tWIUW4T2mATacrXgJKdo5qx+Z3GQV1U91NrSHlw5RhjwoYFfutwQaEVsM
vje/sq5KTALWQ1rMKiV0D4ch4tpAQdpkH3oygw+WbpwHzq87+PWFpyv8wOYRhgHvYhowDCxVrYC5
vAm3LC/2stINPBGfHZBTpz7OHGrzylAFg1FYswe9zxfF0XM2qm8A8umsriqZpM4ar4ghtG9VibpC
hi1owAwCMj5bpigAPduuW472rwi4WubiPp/1lC276hQnhyqpCI8ctv91EL5C4f7VDzWQEIp9M0Rp
PQU1fzvJPv9ocQPph7e78qbaB3oEZ1KdSRtwVZLIUrJ7CzzKaJ2qybjziCmnuZlD9Ocyr/wdVxnu
qLmhmFVtxT25XYXRzYhc2uuZcxCpNwZsRnfg3x8kJX7vzSzJXLBtPBFnVstJpkwUfEzFf3uQ4r6/
6yd/xKKsA3WFxi4+aX8C0hLg2eCcu2uXz1awmJN4HkmjSCIYErNMZxVRnzyn4dThfYCIOd6BKQVx
IDpiK+b/frxRrUhvsJ1HhUouMukAbaJ1ltR5ettf/uTU5qV4GM1FtNkWOX0tBTbcIk9BKeQdgNit
5ghZr74Z68IPKfLTrHnkdAsPsfQDewwq2nFj7/nRtYBHjPqGRtxo821TlnCma87AxoxlXNlyzu8L
dYrZyaHqqU4da1l2hnYV+DmeOUoIcJbNnwpLE1d25AyNWS4wHiqgkTBpA+Aor/FMHTBvd3uDyUJ7
RbyIKnHJ6Cg46HfBXKCVNhGfSamxDEs1Vk4GYz9sle/pgmsgux9UsP91nE/iYKSjL6a3iCifk6hI
mFCtgv8Jfdb/3Wwng9WJ9usr6YWk9oHMPnnsZFJbyoFUZ4EF8mz19YTMLIXoGvBMAxfEVWxfYiWR
PYUundhDxMAkHEoUA1D9LrrekA+PBObbS/7Q0tkjpsugM68KZ72Rk5mkZ17/Q9ehPg2vHMe3XNwB
uN8O1he+XnuklNtkJnL+3Ln0C89afAbDdyK5gNt2sZ0KERO5YdPUTn9/Qoj7v6cBO3sxyP40tbqC
bzQoFocgWaOEoChOOAgwvNYfXICCAtns1WJMZJ8j8s4ueZKBxL/AkE9I4j3vym1bj0jg7ZbIXIkO
iiX8buYwbtWQxb3sUdZplB5baap9uOhk94PpXn66bRxPIW5utsBCb+9j7Z8q5fL8hbj6AKejyoeQ
pXwEO60suLetlgnN9KAUmdIOL+GF4XGEv8+ijciXxBKWPajc6Xe4Dd/ptPwk+LVqfYIqsyOrkqnQ
ay9ypUIxM5VOuUYM4KB28/5YMNYVZSlxXjBTbuAz/O3b1BzSFbR5XHtuDdKOlraxhrwgNT4SXsuB
CcMYD7KXLyjzBKubot2GZaDEZrZAhopIwhDCLT2W6GCUZu7CaeItfam5hmQ3iCycB0FhD39h1ckO
osFdsHjs3Y5cUcevPrtG8LPMAGDC5+UssOK65guOQnK6ue17e4ZOuuWfpel+jD9OBi6ajcqrBS0s
0JwjoyCMhWMX91cRwLc2CcE3zfv+HX4M+33j2KJ7bPWEueIxHVDExnCfSpVQIWEGu0nLXw2Md53S
Pfi2woUKs9rQyA0QSk7rjl7OmGu0T4NIAMUjXs4yiv2hInGWsG9mBpFhmj5t463sbawKlvsSUKCL
aySeS5O7GlgxGuMdaIzIprAeIK0X/+IFZtbLv9cy0kIrvf/hDGTJ2iANQVbb1nP+O9lbQec2y0dJ
Qk+h1pOV5GzxLA+6lpK2ne8RtpgqvBL5NIkHfZI4xe/naSrKz1DkANSS69g9eLaqq6lwtrV1e/Y2
4l0ObdZHasIUwOpFzNcLkl0BvJTZjgGuknCwPRVmSeeC0kps1pzHR9SPIDEywYBW8y/Czczh2Ixr
btbrOL8unCIKG9eR3D938PdlxsHulExCli6lzOjnzH9Xzd3XojiNEm5DNy/nfgwsHPRWyhRyTjyz
Aqt1XNLMOJKQatuCnfnfqJyyc/iTk7Z/mP+YMSDdbUTd4wLvpcBZKJRr2cBIrV+XeHNPZAWqSPTM
nHY0Dm53iJzShDwgMNKcHm4JHnjrHi3Fo//lc/9vbCgJ7tNN+f5pq1RAXfdHnpVecx9nHo4GqCco
AdSTGh1hQzt1E6Y8ad7FkljooY4jux5Z1l+h3if4PIQb8c25c+mpPXmoVp2ELzaKxaDSywSk+8QP
O02/ru62ZeTMp2r6xFbg1mA1qzkQhOR1+BUyvFwHQMvFDwGsYzCH1tjK0AIsBazd2mkApz037qJ5
tA+BH1Sw/4B/ozdlYxNlDdnpabfMTxQldBQ0/MBV455fbZ4Oww3q56DzYXHtI6nvZIvXMqHaVBWH
kkJ4AEMz4d1gvUhLu6alnqF4+LRbzi2ULOzOSSoRBsF1o+6vyLs2umBD7niKzvdY1BxrWwI1SDca
glnA0LyTh2RUijbJxuQ8mgDbjHMzKuITGLi/kWrW94UnczBlye/aCgBkYeErNZzZCQBfHCSQHjeN
ir7ZTm6kd1xR28xaM96da4s0EZ9k33COXod24Aj8cBfd3hEIL+ozw1gZQRGf1ogH1pmDZmrt4PRK
1jNVAqd4vfEfP5RQODgHfBcoihV81RTJerncSBeTy/aSqLr2uHoY5XjZTv8hO4mjzr2NvKYYdr/B
x9FcfdWCl9KhsDvniOC5qrLGXtDZcS4UG+BGW/2KJgi5s74iju5oI/C+yidxIfojChuqVwVUOqwk
3khuAkwqlcEKzNeCp6erCcEvXbd+fHJfc5CnfNmdmXMK4s51qzEw6m8+ULmkHWkqqT2einLXKrHN
eS7P4NSa/QiC2F5rUIZtcHFOYWp4DpMwKQJzjpLdqWETdBiMtJEL2hSiDCGD6TBJiiYaGRQ0BM9/
lOADx0/9aVKhG3tp/MYf1BEF8hLR+lZgpvZ+ECR1Xl9c+cw2JHNf3XXsQDL+UNk1ZZa1NzSmbVyA
9sJZagaLq5vD42lqHQ71y70UrRx0rBADMt6LZXnzqbjaVOMS6nOcTasLDneRO897hwoyVMK8HV1f
iioAm3NRWvIq2OBITR/lC0U3ChMV2B+MTyOIm4MBMhfhkQZZoxJ/SgwAe+g2PD8gkaNBFGa7DfLN
5wJkSQLGxU+vph4aH+G/txXmeEpqUwg+PhMlBOVd/frmeH6K+zckPymJcQIhhlDYLIeGX1edstOs
ZHPedRwNfklveZjRrwH9Kt/Om4MjIpbAvTVytoaowtckgMTEE7NZ2fjulCDpkLm7YRp1yu87cZZ4
ArwR3Pn2ShKVPSdlBJnSbDRev+PxPNqcAvXJmngxqWXP9/FHdYqThT+IRp90sS5F50OY5TZxxUdp
AHWhAFp3Ai+wAOH+HkfIfsIlMGdvWBtTcbvB0/5vnyPpmUJqvxZR+5h7R/RCqlbX2YX4EaiaD7T3
VjNd4YYnMseTd+hsSAbXmVRmd/LDyUklUvR1zOIbVYSJcsltFFUKiWErntbiHVnUESu0d45QKpb0
7TT0Z+AmapiN5v6p2T81AoQuGLPLsTjDUi9K3oLzLkwseqzHHQexNfTE70/1aYpfyl646tqCOGEv
XknKSq/LvwyoHuYNLEl/7IrX6Ncxwyd1BhHEYC1Pe04qq6MeUNC9RiIWUqvQYW8Olvh1j/kptqIU
dsN7HcSouvXCLABqgkq8VHeSFUW0Cb4Cf/I1ts4Xk7dW3wM6J0cySAkvbPGaNPtZlT+RVGBn2CMW
G5tBR+aBO2fDoNKMTeRtYhqopbZfze4KkgmbdF/yW/UjLpF5uOx78O/yl4x+KKBugdwdjWRmQ6q8
1eDroQShJ+6vX0hTsqwQ0DRT20+CwA+xHFUuV+OMwcMKWXcbhxdKmqKE0hRgolLUANrAM4TgeoyG
e70/SGdsPnWZm/EOjTXjpRvxQad51mWP5a8GMJSqR4o4FKyIDlVRBjyXugUSGckKhukuAJlMeiia
yMla6140p8Jm+DnI3fe+O2l0NFP42DxRqgzYDEmQq3bsKP+UQG+Z0C3IlFH07ZSlKs0MnmI8nVuT
OE9I4+qlmI6cRO4Ez4WzcIsO7bOA7V1DG8xWtT0e+gHbkr33L/Ii8WA8ll57q/QnVbhqIDeabrJ+
1e6Sp6OwDl7+MrpQEaF7DNGClSTLCCuI2UUmfrevkJvnUSGvoZr+XlAwgCdWUbtobWrDsEK2Fay3
srRB7iNJe+k4/uInwpIzirrponMIvnWVmXA4/6hszWK3lfdwsRYnuN4eycCfHhUi5eKixnn0LFdN
KbWYz6MjdBQjoX7VQfNfTG8KSN0vWmvvNQ8YqQpxpZdI4o542tAwzD29rwuXUmFfbq4LfdCmRAWZ
Fbt4pIaeKv2J3/sbjYXYxzvmIX3tlQjq5XN+OHuPDz9VjJgpmkDMR4fLn3pHGNbN7LU6Tlq8EZiv
F/k/GATT1kdKXBVBkIQ/RYiOnvAik3JPF0jlJu3vW9rohavRTGYkU4b7N3UCX3oONJGQGLs+5wPj
shZ3rXLKrEYPj3+iPSvqy8DCynSafr9NtB5KRbCO7Uwmfvp0rd4QgU8f/dJ280yn7LJxQ0ByDJJm
6Zv0f1eBAIZf0qGziAjvEToo7ngljSdU1toas9LOQgU6RIms5F+/9RNKlyj882E7FHfR9ADJGrRt
63pfHrJv+br6paqzpIulhqk6kgH7YZK5u99XFbSRwf46zDKTrnqgHRnOBtoDArgwJ708LbJOwMwa
Y/uPFSY+xogFxO4DzMJEbshvJ6CQvkJfQmfcD+TAZyYHYE5y0ESvpvTycnO/ZOLT3d/ZeKfjPXz6
N6EAeyTILu9ZckMNb0EdDZDt+Hh6GPgAZOzM/saGpfE4EmhXzLR9QK/d66VHd0n4kXBoElEQpXlr
wsDbwiBjFOb2aPaDe2s8hZniNeXEI0OuotS7JfH8dylW2ghJPjJJfuUNJ3ZIxIL3TsProgj9+7Ey
nuJL6CefPO9hYezOSnU50aSuF07qSYg9+iT+SvDOkD7gmAUxIJYvkG16XARpqmbN8x7EVUJSPloD
bgiN8qmFMeDZXkaZnyMNy/l0yz7urMVCPZi1ku8iV70nQe8UkAWK82MsiA3KWYoRG0TUe2gTGF2f
zmrRTeSfIFWKwx1TnKTwdwehVcKDxJxYyGfeqqGikoDeWmYwFKatQ4Xy32UldT+rsLSdS4yX75CJ
M7ihmWbbjQD1deaTW+3zQSCHqpVmoRDZlkB69LwnEwiMt2f28LkO2VFgbHmtJJg6spgOvzixl4Ib
TQd+PhASyIvXWhhVKSpBgVAIwL8SfnbiNOn9ub07mKDI0DKQoNlY3WKkF8pMoVtHJAf6/e5tjeF6
44fjt/TV04lScPqeMP0xe9LA1c59jUTHLI5/+tEz+l2cEM1mys/63atqPvrFdWyPbeRSeLVNt9uW
V4IkS4I1mmsnnJjASRvrV2mBWASaYkPez4D6tw1Z4Dz4zEYGV0eBW+q4aFNzwblOeBu7RryFB1sN
N6MijUfjMmNry68Sk2qK/lxsW2/0k4B7PZwe9LGFpsP0If/M5XIRrKJDWGiUOuLA9y/7d0RUe1qC
HJ0tKSuGnIpNCZ9DTKUWQkfwJNxaccgEygaZ+UTlfRRjq25ccX94KutB/46WApYKSH9nrqO0ct/a
QtKn/rEAIbunF/UNL8bd35gty0jd60JQ/rXzzB2xajhs6PXpNt0SsuLcBcsOmGBuUIUYHGAqc8Qr
iBvljYcOKF145uJA4+xwwzOv5OF43GipgLnColCphivUt27+JJClx6tbiKpBvl6YfOdgM+ePnuhA
repYH2PtZBiXp17OqAxNFpaYaV1qjnRxfUEaNtw2/4+vmMezsKQoQonisrQgyCq+sknI/Il9T4Pn
erNAGym5UMEX8B2uZeeZ42F4zkm07AMNigOZQMbxfvBOoxXcEE/SfHk9oyX/+U4F5ipk0mVUvEeZ
vdUC+ezAsMaDUHnHfztEWxVrcO9xipZdll4i8IlsLay3AO7avVNOtTdUCevbPP/vbjcDNQDRMZ9m
fKVV6zS8gLlF8JItgipobhpncVuTBdD0Z+BvlV9eBHZkM7uicowlAgALRpZ0S3LEwHQosk6fl06B
6VhYI9B4omXC7C783mkC1vQ00q0h0M6kK3ENeEptfPy3acUdId//PdRQi/+9kA3mKwWYbugU7nZY
fdyEb3DGdP7ONlpW5K8ZIju7IhaYTY2Vh7LxSmbpr5V1FcKzJMmx/ewQtjVYEJHJODoBiO3m7iZQ
AwYZlYvtBcDQ/LOVBKpOSBTxBs5xv1G6wT751Y48m9/WZuNGyOeN+qDEso3lpx1ZZSk66pKQJgm4
JiB2Mv981TMsIQi37dKa0nAvwPOpGTfhWMKmLp4/u3g/8nqsjSXE1WwuebFT1SfchRpUP0a5CZbu
n84rdoPEIW1OSLG54/H1rLz/cqsOxK/r9MRAQrQaI7cBxNabyptYVlCK8LlRmNrV/ymErW36+BdK
3PUKDlU2UzRwF1ZKHXS6SwVNbYFxJcftY3ZRXtFQgorq1T8UeM+SQgZXIfcwseea6j25cmFX4Hzm
VS0x7NvnRCFrbtX+gPYuFENE/uP3dIguxp4I+jUaYBxvfoIB7vYr0EbDPglw7Z8L8JQMgBaSqBEr
jEefN2h46mBr1SpTMXzMzIa+zBKs+rBLtqnux9024S07LeiwLn2bWFmF3Y4PLmSEjvQh6SM5QfQZ
ZujqSSMciGS4vJrOmHQ+c8LfH71Q1XcF3wUlsbyRzFkXDIVMgClwzPSSOMNVOu9H60YUT4Jx7p/E
1tvJG/jf4jtFCMVI2OLgSlOipkCLfOQNFj/bs3VdaRXH9vL7DFiS0udwT/e+O4+JQdo/5qdGmnu2
Tms8wGIOkqpaH2o2w2nVxsOuSVKB4Y2Bz1PBBmS9bJxO3yGNwm+zhd6nDS1NSfe6Y7qaWDRT3IBL
S+FxMZ6gOx5ilvT3ToeyT1RVieEyR3LmxipaHK29EwGw/Z/fEfeWb9y3mYLSFI61mr6tO/ZB+iqe
n4WuPYby9w5qNMqdM/55ib9I9BS/mU5jLFhg0KzKgLN2VGRSF+0CYJU40Fa/lxLYbXdvz7d/XWHg
3sVyrIRJnxc8RmJVJoNa6cM7lNMlCZ2nzJ0OjlMd8sl0mH8AQ3WIbdgz6M5xYqiaPn2hyhhxVXvf
dDcJRTgRHy2HTMBnPCn5wOHV0kHrkhStP9HlPVZr1B3cChvClA9BHEwQlxDOi7whjPkMlwB4YvdP
dHSJLcJ6D+CytsTPxhqnmCUeUwfCZWqIbCeNpagsJ1VU7N9/STAXeEUD8tXdmYI7Dp8iSIsqz8nk
BH3ukadCfbxxwBrtBZGSVcf+/lFsWpLC61jF0IQfiCPWd0WLLSNt2Uc1iOEuGfUNgaxCZor1UD0V
XpDOdSOVHQ385DF+kMCpVeYeXbsNgdelRXF/qTwgVE1IJBRIWA4Suj3iu4xqmx9x5w0+M1EV4Sdl
fHhpdKASPfyPRTibc+XsL11fGWcWQbZI3bTDVNnkomxj0YJyx4OrtjX5tm5R+fN6MeFubyOuFOFp
cjpuB5I9asIIY5lsKN/FKg4h26tt6XBgvnAveFmwDV9K0pffJRW5AoIk3RHb55QEKVnCgYc59uWS
aNKyo9HqDWjd2S+Bz0XWmzuSCZLbTqqCNFdWKB0WTBOXvUMYL0i1oovSmMa83+CcXixtZ/ORTIkr
TzjqvK621pRA84s6284JUyyfGgYr1VBYLSuiccOkHtahKnesQGbhXaHJY/Lm7H2Hx/l4b9OyPvyQ
91wgPLTa0v0MlDwT0id4CXjUJsY3KdNTJmNVx/9IdWJsBlZ+JdopE0DAWhx/J51eBviaYsyZWlhs
VaSoQ8MT0SaKy2Widc6tmcKMHSDRD5dA6oAd39M17Lgtzj5hoMm4tqiQ+ATBy7YCzW/Hr0/C/HGz
TX6KcaUpgFx/gsE0g3uRg533VEx7UaTQPQHmqo8pBG6MhCEeLsiyAV1CAfSNVtaya1VXWRLsO1Tc
YrdemAD2dSlwHQPS/m29MPbuFGw3wj0dvYDvxwISVVHvyoSZHCcEz6JxXm7kmf6IrnTnUA+2ssE5
RJxTKwGYH4aUC1pQILyQGG7ewx5WBnlfS3yKBo2bXcWB1CbNjMTEDw5cXypdqj6LX+rjCNlrno27
Zs7U5rmo5XW32vXzChVD1q5i9UcfgwS5nX4H0Q/Md66sOib+JLlYi+SpaExazWytID/SIqv2tmJY
oGxe9vxGrvHRmWn7VOLcDzF6pFZdLq5PjYPqVQxc1xJS8Hx8KifLBse1uDBmQL1H7ZS9FxwergC/
kj97IlFIlKsZSGd0teGEfA3HpKfjRMEtPMsPpmNUO8FQF9b1+OjewdYd2Ge6Stzxw6W0/zhrrQdu
g3cNAot2zWjk2tXeU2IdbiNftuKgwzGyV+96nYLdbuEQX+iY7Pcm4hfPs5LNc1lA/z9BTjJpr2bl
5xC1ISSCBNeYhhaC0/zQHo7feeDswNmtCyKK5XUuFY8rHW88yjkFsCewc5zDvnSmZFTzKOzgiR2i
+try8xE1cZwG45Ma/BlVJJeDdGICsckaMduz25pxonaHv95alAZeNInipn2tSeva3DLwLrulGSRx
bfufi4lV3fZzFVD5aVA3Gckkc/4jy4dPU7DUkj/LcsCnjfNflkZZbvqdEHm3E2w7ieHOyuYB4UMK
MdAuGVlFWPUMK1Js90ykbKLbS698NwRpxAUODaeJHH4xVG58VoOSjBQAhC6NqMDdXC9jyb+MEl/P
e5IbvFDyZRejrIAb3aXxB0HAhKx7P2X7G//S0ztO6Ot9UB3UzBGA92Cm5XhkGX1B5eiKIQz/oUk9
+G8srrWVkeKvpJfitbrdxK3Ba3cTm2mV7vS7vlkeGrdERp0wttqy45x5LS8/dJj+VyGZD9S9cXa8
0JVxU3yGHFo0dkHNM/OTdMa3OB1EqjQuO/JtRi793/0XnXijgPTkUJPrtYdxVHG6jVx5YXzqtkhg
wxeawDU4sQF+VxmhS6Iwc74Y89CYfRi6FSglYvMqSdfuQnPDHWt0eUqozDSUPy4c/6boSt7C+qun
vJ5wT9ADRqQoKcOn9aSRtk59ohTjOXSB76pcfM45vLEJBoaXBJCPGoDVNte9JiitxMV2RFLX1dK0
4vBP6XZGlXc8G4jWqj2WnJulyhKn8IeAh50erzYVIDopn8xQWdymu/Tp1O6OF6OnN5x78+Qk0xWF
2Ck0NAJUARnkW4XJiZw/72O+FMA1QFFHj6YtnZxqs99fsttaINP9upnTbexNnIKydAOsOlQiXRuS
76OJYsO7l3vn6ez9apXZ8VQCMhLZ/HcJgEra2fbcLPyI5WKOWl6UJPrC64EZ/KCuXvHU90rkjcoL
xG+XcoUK72ZjdUbwOCk82Jw7XSxfXoyUn0WYJq+IcB5YWZuRk9PeiMyoHxsFKjcH0N9ObNQxfPYO
NMfANymGtiwB+a+xhfUIJGrhmWNig8tOkSypCzSz8WXQSwMQWK2YWtxsg3NlAolKIAlX8ia0xOLX
dC2FrLjTnhL5bVcCNrZlEs+9tDOHHRl2wgxQ3cO1uuvpW7F6Q6GzHC8R45OG0S3fUxJucsufDTgX
nxd7qu/8J5fxmDnf0SXS32A9mo13L/9WxeyA4q2clDD7k0VrJuXQpcSzYgQbnXOc4ZscVZ5keoJd
WVil4Zhpt0Q3O4vTXXHC+ZIdto29mq5mP7MqppgNMqw8ZNwThjYNPLwUTfUmA2f02y9+0KQAPo8U
Va1uKmRZDXjBXUQ0EhQl+WEHQvTbPn0q+9Q4QXZ8t79OTdWoNTU44er3ayJqeS9YQZzvm9Fa0M/l
qcDVy4DgWE4GkziG2xUXDyBEYMlIEojWtw9CC243J8ahUcH/vZVu7arm8TeZHtod9wao5EyiJNYK
P4G4pRxpCjDEQzCsGKAVHPyt8tR1GYvELK2qf1NAisvptLlV/diIN1zTQwuYQnqqYgyV2o+giP/g
GOqKXphd5yvLSL0qjfbUStopomrSjKW/PDxtWRgLZ2QupHf+pThWNBSelU1XILIh/tCFF2BwaBUt
mYyXVovElISvpDsaDBD05woz1md1K87FkCKYTdQ8EfjdcrJu2izo8O9ZQ3x7t3qYkEkD0Ju6hy40
S4Vhzp37tKZKXE7gBNn0qwLlW2YhFqzoZyc6iRn95nI8kKIxuYsohdxMMiWsS7Rc0ybXDHi+t7S3
7WvaXohXm5nYByFRWKXrphTdBfKVWMuSFTFZdOtd5aPj9B52AgEb7oU9qKwPENaeLUN5eboC8vem
yTFyHjY95oPEkXHIPnEpmlGHfUKmUc9coQQ98zQ/IMJlv3DL3cnehQIK50VFxw6FbF3/zWgIqDsU
1ZfBRnUENccckXIY+5+3Hl0trnRQQvF/+WcLvavCU4yKN58be6SMACN5/IN6d31nIBfnk3/33kDU
xXAsV/lBD45dsY6VM+Ls9NarsfR9648PfDEEmaPDwCTC7PNbnI7KFUCNpfwHsrBVnjY1C0VR+jLI
vhF5vDFwaqd0F2oU0KITde3lbOkfGnN/M6znOyTkQvHnTQUwlpbhOAi5zU9Ln/g4Wt79RIQN5og/
BBVdAlLlSlr6I5ew5sJMVDtbO5sC4rc8/Qg4yw5wmCIlPTDPacX5oWLtaDMSz08Bl6AYUKYmJD2R
UMDd9jk66LVoVrXnGZuYEkFxH73wnW+y2GRn7VZA6jsIwzccY9GvnliMAz4APDckPEiTxip+Lffs
Fm2IS3O6Dl1lVi7o0VoRHNxs2//qSAS0Utpj94EsNH1m/ZHsLoRcExMk4o/pX4R/hMOphDD7kgzR
x/YMSEpcGDsRoWLODupFpPjuefe6BgdhcxotRwFym3jZ0Jc7rvUPq6EtlGK0+D708h05Cu8sfIF2
gIeNTK8YmEdZvHe+XbhOBOH0PbEpwCjkeCDOLLNTIjrsTdM7w+liJ+sIaJey+UU67e4wpikHQKuX
urWjaEQ7B4ao+NxFCbE4LIB8hxdB+/yyRast5hPVqs7avMiemeoDKLRQSe2cBW1TSMev+d6qQ5g5
c4ExZzUospn30RIlBVvXvmvDYNQjfBwaqmyZDAey+2xP6In8+MuwIz8AUPlR1rWMxxMXq3f4lsWd
TCjzPO7mpVknlKvoua5i/lJvVLg3FgfkK6x+VIOGIGM4+GjZAi/N2Ofwqeo3nzrzbZOVjG7lnTeC
ICbLCst6PPtsi/IOe76fwcGiCIlTHhWklhatwvGn3AoEk3zVR9xeGBhDGQmNouM16/ZGwon/ORnh
YgMHaGnf9q2HUgNnhObkvkjXUoTWoafbhLOujAwzqXk8WXwkXSjpMnE8KbWQUycaMw4bIaXjfi0t
QTPgJag0tKTEls3YHoFFYU8AwHU4wq7tVsG53oDXECP5j2OYoNYasKQ8iQZUqLgmVz/6BJr8zYDj
HoEeK0QQkZ9xZAFgmxiiKyP4j98OkHV1gl2RZMmCasnFuNkR4jrgsGw9nHEsAAcm3r7/CQ7n5WHx
TuKbvU7CuhG/IUEoNtKN5QAeeYhVfQ4oKna6dZ7pKddApVlbwqnReYN+p8o5jzHrzsJ6yelxtU91
wP6UPhYJBrHH/Styy7SXFt85+Tm3ee1QVnVRQygRj7QIjnQtyZjtbxjwWec81kGVzhyBENFdJKhM
8biz3Z8bbJA8JnwM2gWL3UoKVQ0C/o/YzbXz1H4OltEKNMCAc+ssWo9p9JYA7Tmk5UlFvG43Y1LX
5sSsAOtraszGqhhRppC3q66YmM3zY5/kDSo5GRyFWPQAqwTZv7okg6MTmbiQ7hPIdMyWdTOm4hxe
K0yzkVPq7Z/bj10K85ZfN29QzRKEz6/79IRLnbch/dpX1O8eRaOGFFUCGd87B1t9M4re+Bjgy0JD
TlFTYUk/tGUWoByDze9ZyTVvNVCW+yxWrt8AayflRkWUpZRlCHv98+YsyJ9uRHaCyEfzVpkU3kiJ
9z1d95luQkYaaBHC49WLkHTLafK4LfSKa1Mf7tpGYjNQcbYuifGxE/FXbxx7NypeCfDUyXbIQ0v5
WoGs0DZT4SlA9/adCFroop+bsaGt8AcXH57RpQBeqQzOQiBDjcrRmU96lxROhenTf4oCX3cYi/Ur
4QyulmyX1XnnXfjosF+yzKyz3jZVG0H7//qk05rPd9K9gCpDsmBZJVyO5Rpl6k+ZLjfB3EjDCFkN
nxx6kc2fE6APsIG8Mlw8sig3NHIW6peUULyIPee1DOzfZb/bLDjkwnDMqIirfsA0iL8nkckrELtS
CBpNLjh9Hg2d6HoY6g73G182G6TXxBi7HAQrAZfepZ5RnKtxkP6lFQ8z1yuwCrNGq1oUVmvQP4dT
E09uaLAo+0ASRED8UqBaBMg+0OxN/+WEHBsC//+O1q+IZgTiF112fRfqj7r9g/DB/BWZs7Tgq1MI
xFTMyUY7isFzAPD9xW7Ptau79uxz2iKgk2kFgTQMCPsWTi2rLCaMEKuBqCqc5DC8Bf+JcZVZDpuH
7S4LIepCQTPzQ7xSnic3mTnx7KXytqFfaDTEeEsuZZKhq9vvzyobO0iGCUulnJ6OGD7/xP7J+Aro
sPZFt/w5xU+p5k07CM/wBhr5DEWItQ7a+pAxAV2vOdznC2JDgxvRkerE07v4YtyPUz05eM/GA2R9
339uiuMXD3dduBd2CYlXn8IbP512oytxgyolHsnKjmecEgVO1EN3UMDGBamZ0k8AM5kKNo7M+YqW
UfrONf0WVCo6dE85t2shzLfZy5shloNlRB7T1ZxaSAiBAq/u6CQKFjk6wkyP8fwYaj1NzHuY9mlU
mkB9RxqeFOLKqsmo4QcXqJbqoDqOOCPCXSI5c8naxUYLLmscdALYGRVk71E3rv5gS3J3RMAt8UDJ
TiZoz8qRmhHS6XTVyulPJgaQ57faSbhVbfn19wIVUs27LxK7YkT1ypBAic2u4yMFDaQrG0v76eaG
74MCD6I7ruAvqJnVS5zXp7rcOZhq43n4a/IKMYmm7jTDG3jWNNO86S67tE4x/MsMcInokpJN7RmG
Vu85MKWF+8lmxBzVII6jO+zoDjVnFAjZQ0LlyeJts5HQ8Uj8KstkC7q7g54bzFZwwZAlGW9H/XpU
m78IdBJNL+4xlyaWmnf0V3K3fTsgWTSVsdvgkt4+ilcXAttEmKjgk4Ebec7GopScLOpXR3iCb0wz
yIwF6EhczEpbGhsDgp+l4AysWf8Bqn8P5QfkPpSlSpXleW7QlY4tMsqFZK1HT8tf6jiO4B6qz0gW
23l4RQv8ylND/nbVPZ6ZcLVdU7L5P6oyC0a/W4r53d4x2BDrzjbiCK6DLoMbfe/m8V9pKulvxioW
SP8ruBaTnJ4T2CTTjXhYzBqis8lzvstb1g2GvCeKBBSTkCDVH/+N7eT5vJFyIVseoPFoPau52i6r
+pLlgLk2QM1nmm33xD2NLordeZ+gVSHA/wflKVDzvBeq1td7ZRduKXOu/pzea8kAIlrUMtuCIDgA
Q+IjdZo1PtJRWtId+H4goZCbfcovI+GLV4O6/6lLKeYy5HTNKzTVTG21+G03l3NMmFKhf3qOsYNu
hksO4jV5AR8L8wRuf/Nfe32/MKnFW4WV6WrSLqf/+dusmQK4koPMUUIvkQMiDhliK1MRmz3Bo/+q
b4Gpi9ajZmh5Q2uQWwC86SFpU2Er+JXUbz9qh/Jdo/cMEkq4nX3XiaaggWaQbG1S7tJwZ8qKVqhk
0KTDJyhP/jtMBanEFcGvEFbhlnT8gQhgZhj2XTSNV0PgR3xuVZp7Odp5NtcAWulqXKh2dtgVAcGv
iKwXnOdEE3PmWRCEm290DHRZTGu7ABeumfy7fHyg+pWxkmXkCOMUCV5sLPP74JfaEZnsCBYgtKEk
AQ55sQT4j3ZIBXmyujE1Bt8nsNo1sYDd8rXNr+sWaYmJXcn8bLlM2O+hstmnwDx1JEg0CsyoHyFB
boUUioqG0cdCEcwadjLm4JIYdSQmrEGyQW8wo0IkbrWnLOfDV8Vr/sLuomf2OLqoQ2dTNu2sKElS
/CLo5hNQ/1EnyC85P6ZsQfnyQBLsTxbSC3jVxtZ76b3FuMJl437FeUtHIBSRDWkwL01YP8Bu9vQP
FuXC/eOnTViR+wgAx8xLIVQaVtxJ+mFnoApWf0t/rdMjhmGWFbbshOhArKWEXhSzMSEhcc2/rnH6
erz02IgH92rFw8jP1bmFmCyygYx8L+IWprLj+BefpIRV39hkfaCjtBDpIavHUuNIRn3co+0giPRX
9e9CSYipzO74WaNAy8SUkZ47w2DzovSS0kOKZMZJTaA13EbjIB8FfyrDOLDMKvU1zzsvpL1frtuJ
WEayWtZ7cYxEbwobK+x2rM8adn8jKhDQn4n+6ofIuoOrtLuVy6xXWO2JupYf/MChz1ffzA30dHJu
3yus1hlTyNDMIdgB4VNusU+37vni6NK8u0drqV15/ekE7G5RulKSkd35TnOk91/nOGsJSY+mdSyi
AKIYIxGIhBV+Lu4WROpdBUeftH9j2xsR2ycV0lzP0qz74N+WWa7doiMMfrmw3gOlj04ozx3fUa6S
hIEisJJdddR1Su98/yDIKriW8OlrpWG7KZB7ufqPx9oo+Q0xtwjBW7MuOlSePKeLlhQTKZP6PCnx
qB5kMjWPNI5Tzg6R3Bjdz9XHe2Cyu0FG8oBbY1rn28YefHV4CAKVl40iF6ZdmjKcSRDxlLbivo2z
HMBiPcWPXd01ZbTKdVdTykDEpDtwDNhYYfIzBXviHNTdIzbtxJN0bsqUAnhNL5eex5siWAkQKYwT
kvGso5aD5XOGmT0u5BmeIPwbyzZau6QOmWm9lr1/RQM+8K0BBmOtCN3BFn43rAn5WJBssI1evs4E
kWLLBWC4BginGcGTzZRPAL49PBY902NsR8o0IqFwuJdSjV6fZY709M0Pgl2htXxpnJox+E3Q75CN
5G1FBeKw4Q6sSeRQfwLvXSo7yl9ULdPQub3uHVSLcAaeKZcbb9F0Ywm26w2zbmOixANVDTUBg9Li
17cUn9VFtLhoZST4V0k33ZwPOiOsKtn0krl3t15smz6WIMlpWHV7TQcYFTVzIvwBuxOwRSFEiqID
LsQVlx8sM2sb3xQirRc2rdRBtjQAXSVrU8+de9te+ykqtCKC0P7uUqk9XlJ9Ax3aontG+iluVfPR
IqanrFPKo9S5lYzHqBfNukQsQTj42ikRTYJ6fvCIZBzJWKtVfFr7AMwPXXYDtSgSIIqLyn+ExN9A
teKRHexZ3gYunRFlQLhZsZlQsX1lteZf0ZO1HW34Cly3EtxlgBh4NNEBwRgz5jVHNLyeqYeDpJgC
sNgd0oNbTx8SelzPhONrEQa61lb+UiXDtplYRUeapkMl1N6C0KukPUqoU9ZiWgC4rzXNeRfo3zlW
h/7NwqUhbDOt7Igt2o68MRSrRXpFjwZ4pxC5MuhLqAlXVYe15nL6YenM5EjnWz4aApL/o6j/QnAB
fCMd5eKrUIeQ2YFBBkVKTHVkKVoRVPXlYwFv1RORGu4qgt3wiX9pM9CS1Jc89Msx1WoN8KlMzDK1
0jEorEDdCfAF+BDFnPglASPr0A6ynmXQ22oXTXZLOqxYVUSfBs7cmx/0rHeznUXvKRIBepERb0r+
PYRX8PhSGEPk2CJGE64EK4uUMzZfRNNb0uJqFyzm5vXQ8eGu/iCwHPZxvg6vleG6q0oquWFzu/Iq
+vqFKV5Q1JcbOkLDIIlhUDiafMKhQAF0ELQ0HClHF7o7y5JNRksEPhQokufnh8QlY3aKEqKWUO/d
SqV3cUN3+tvKgT1h/yy2h33aMSmjjhRBjzzK7TrOSYeeMTrT0eslNJgy0x+RHfX0YzM86WyokXOn
h0jcWa27YmiLttrdvj5SPO5pxZt2W9p+opOBtK8ain9tbuInBuQSMC3QlxLClif/eCew08wICmHA
axpLq2L9hckBf9ZQ4QoF+psOdoxDDmHDHWHbPmDvlcAOUmzkjmD6kiB92ZcHs9zgVPC8jn0R3cdA
IFqToYUK5TvchpZpKAqGtauJfcR7Y/L/nDhe+Vbz6NiVFrcsJGG2giplXLS0RWvbQVwO81TAYZP8
yuBUblhrjAujGBKN/t2oL+NSSNBvinB+HmbamMlQGBtuihpAHfW7CrobVFh6VjLxQKQMoW/v7+3y
jmwcG8Neg9zcWXkLK8zzuUW/5y0LKICtKftlyjbVFQqSF0YQf3VK5yJ7E7VHt7baN1YL8Q26m2g4
0nKBdDJktqZDdyo3c4HUbmgO8wsG/58BYhGyO3228bt6eY6Z+gTOr3pomCSHlDxlRnpweeAuG8+b
aurCU83lOHOcM8hmuALywE99f1i20ahjef6oi1+DELofCYO8Om+TQY0hOihE3mrVSwGBX9zBi5Cr
sZ0zRhDxoRAFy7bJmFGh2+LBTxx+kOeycXgs9lQME2kiWvcbknsFLEKE5G8WLn/u5Do/aZXfnQZJ
jWL5BqygDGtXt8UVT7o6AuUFE6YaGC88OIg7DEOkHtjDf+WYXGroJugVI5WEbgOPGVetMVkK5hxx
giMj7akkjirYa62SkT9nwSgyjkJO+Wdj8dEn36Ag4t8p5QmG6vSpjcs4ECl3p8ECu2ahvSIhNcL1
bvxEKTR08BDRdk1Fa9DKvQgBhA0iP8R4AV0nmzdMOloXNj1qRfm1Fe3u5Asiw7xrac7RANwG1yYe
nVY5hUl8TqK1qIry3U53tJl+ev96jAIv8TV8L59cq9USlzHoDgOqJ8dVnARp8sOfMmC2UTYsr96s
grjCTtT3cP+l2TC+BL+nmghzjZGHC6+SgDeYT+DJ0zY6iURGQkKcnBfaGgOVQvsNNUPP4/46TPcw
Ujf9nJ75nAuuKYm6mA9+QD8zwPNEm52B12g+kwWyBxolfeu3kY/XNiQhZcJvyy88ZBQQvSf0q4W2
BndrFTasj4S7OEZX7Im3qwDxlRmWYS8q3W3RUdI0aLE2Snt7M5dPz/m2A6XQgR4RVNVINqagN5w2
iOOKUaaw4quUGZD+m1Y3nkyDCKLjarwrvb4JE5HNQmmKQRfWktMG/xlNP8ZinyyoQaapgFtt+/Bm
4ahqmF6p+CknLHmkgwNn9pG5qML022PCjUJeZHWObqxnU25WKfm7sF0q7NtECJWmoPc+d1hiZP9t
7/c/IDgfknjAfJMsn7MwxiQ4/Me2+nWFhSQQrDBdsCOzjI3BC3KBC5B+5jC/IQunbpen3YqD++TI
ABzl8G99xjMMb+KdqMiRYakBCCXu2sK3VQxPYl5ttf2tx8r08r+2WFi6Zn+oWxCS69VLbbuMjqZj
Mh044SV1qEOMMCGpqEsD/g3Gs3cFWm84oqAzlXY0zf6uhB3P4MruJC9FDm6l0CjmWFCbqq6AHy5K
AyimWCrsmoOr0eUKO5y432z4kCSjptsfAaODpjVn0yBQgYyO+ww4sAybWDIb5DJJkYhWW9k06G4i
DrqFM+gqR7SYxHMaWZ55DAfJpIQ9T04XSmOBee7nIHPcyO1jE722pXihDAvs8xjikczR6WCmL+G5
sIvDvcsYO22XHgBZEnzub9VbrPY0wkfaFDyTHeUkl0Gk9bCghQrRcXjcsl7gmK/qHIi1hryGOYem
JLbYArJRPVMrT+P7AcpvnM339bVmPrO6+R6AuzsgwjsfYcORPxuvR5NKCkPnHHWhtpmRUfkJkxUQ
dNTUxRM0kcvaZFyti5cmSavYSZ6Bv/O/immmjXA8j6/FF56b+XBrkYVdRUih3QpqQEDM42AsO9em
QVoRs5Ev8IY/uMlvlGb4l2tUNhmAE14YSewRRnb9b0p5aKg2sfQ2H6W4cm36kHOnMVm1g0myqoZs
5ISjLNwjPNHb6C5Ej7VF9BZGE5IfCupcrUl/ku7vjNmXxpuSrzNuGKWRl1nfnz8DUV6/8U0WmLP2
8aKh85J/Gs9w0Dov44xCDK5fCX27y/dnuCSuyB7PvbvLz0scB4lcb137depGheLTs7mFiW8ZA/7U
9AwvcuhvHCeHqWpw12jotq6cNr4Lhf+CSdwbhZoRy2GL6PPoxfa+NmRebhemJsr+WWbCQDeKPv+w
q1C4JGGc4NpOZj3OrXa+Af1AL89n6UeMG3heDn42ohweD/TzFWmF8Ud/NhPJcbskO3HvPbj+p949
yS5id6P9L5phB8S9FZmls1+I+UM/mWT4uWHBQUwWIf/JvLsnIrI9b6LVCigJuE4xiWL7rx3QPOYd
uYrDILuJKfrHA0vCCSI0uvRxS26/Vgs6jNR9Omoewk8lA4VagXUHtz2SBmaAJoDcfW5I29KvIKsi
3kb4FVJEP4TKAC4X5uDSBi9CXhz6hR/s1n0TduQmHbXYfvWahErvehhyjdCGk608uiw/APaHSXno
+TRFRu96M1jCGOOfHuB3Uo+BFFyM+XzMZskwmVJ1fqbzVsryhViH5jnXur/2SMZASE7ePiBDPmJm
pq8reU078Ws5EsK8sjBHp+c4Qfb/a1OWnUEM9B7UlQHBn/yu6iitUCcYs4M7Yd6HbSrFV+HvvUEK
vw/+PhznY/+sHtUo6wuKnmes2I/9NR/sdWCAeALfa6qZfjIJebEC8bunn80H/cCgdVh8R6rS02MZ
Li5RS5vxfV4JSENHThatZCWI2B6Uoo3XYfYTzTtxJnvvgpaeE5/r4jtgRu1RyPI8AqyAkYtaNUcb
vpR3GF2oCrZMPSxMjzQwsyTkIl/sJwgYR3tlvd23VKyr4YOvZEyBzUR32I/ANDajhkgaiuIkvGCe
WR6Y9qmZqVaoEHs4AwMHSXlmeiYYJY4Q3cCugoefAaB9HkxzEekNe93daAur5xu0HV6fc4vglUY5
IIoxmU1BKWcYg7bL/meN1eevGGu+TceAr61EbNlxshNRG9VbhIbMj/lN7Ismh9udnnZHsnzgBFxK
kFqbvbqWNz/qqUJNh3cxlLi7niWouNEx+SBHXH7xFf4EZr9o6TcykZwOZd3U9Mx27JN4WnfJNmLO
iH+m8C9c2SG9UNt0cSxhlcV8qimJMm09Rdn7lreieUfFt/z3bZznFeACZfK6xn8B2oDf/680zkAy
1VgrAMgG8jU4bdIk9MTn83rVX4x57/fR/aZL3g1wQYVanCauIKtYHoYk6i8/Z2/r25fpKVP+3/8h
A0icQuhYiz+yiaWEePtzTGNqvGSMGldWG2xIICpOgzgb+DhmCIZWlsq5FVSG80ttrHF0F5ZhBoNs
88uXZPL/koVcVevmnmalP/w30PtnvDfcHsloc3E4OULZ3j8GXUJeupYmXoVqtMzeza9oMfc6ZKNW
1++3y4r8ke8st31iQmPivd9B9svwJNlblo1DQCNNePT5TQRDaUc7Nhyryug0msC/gH5GfP7L13Sk
Qfn8Tbn6ECR8WkGucqFtSAXI26hg09QpcbMbYgbcRIAgvDzo9xf5UPgJq4dwDk/yoQtxhogJgcti
NcHa8Yx3t4xZ6BZDCJ18xNydtc9C70aLUYw2VxQgxnj6ih1hnheDe+lIhpZ+aViUmfJlccyU/nLx
Na8leQ4/0yOcVV6EcB+dQmCL7xvGxKP5Rli+bZCUR5k4a5sVLwaBM2SeJAF2VuddPiCFmdxyv2wU
FFu2DuUpsCAQclTZfBuxrcOA3ijGA4cIzO987iFMeXg4fUyRNQe9Qz0iZZDj+EICfIqvUaaFk/pq
m4YIvQDdWk8iq4SJc6Lk/oM+JSyy9CB9V+ZCld+j5qjG6dqbIGiARR8c8rn9h6FnxITJ8UgmyNOc
of2fahB/Wf2CDL1OlRiuczOhdG3P19KDyZdxK46xZctOa+s/ogvJj77CiihHb6Hf/60MTDM/WzLJ
bqhR4AIfrU+gshtgEDs0sNFOK4Zu0Pc+iRDoeeK2rf59ETlJ/BHLUT2kB2jspcnqxRWqAbRlmOQD
9JRKUbxmn51EMfO3wSZkIZJx5KMq7abbWQXMQ79Kyno8I/fM5TJMRU+hPw06Fqt2Vmdwc6gLLFZn
2WitIzh51cqDg2zGW1jpa+88Ig985Dhh1vN6VshLY6TzSCDho2MHEBdtS0WIHreou/Gixl88zJC3
91PbyRdA7JyNOJpCrw78bOD5OUSJLy5RWHTJSXZofGjVUdD1oQYVRnCo23+n5tCOpimORKk5bBsN
ydQbahfsHSZdR1iboUKqI8BY+ZRleIt5AcVKYSewr4TVOOFCYLQ2oZ1TRw4vlrBK1ODkWbs2mbSO
wEUhqN9w+9kuGU6dhQ6/AjZYQTfFHlxbSEsLyYSF74T+YcI1c0yZyEj65i+SUKU9RehP6fmgtq2W
0A7aBKHtjhHDX5lBaHL14o83pyYN2WWPpPBbxw4AGVb/jk1+Z7zbzz3itBTis789/KygYSTfQmvx
w/N1YH55C3kLu4frbGFfbEg6PMTt3FRwO45pod5caUVab+4ZM4vlAKOtrw50EhZVMIsnBKsjteN+
W6vmeF6NRJNgpvxWF9+DVK/Uu2Ef+rIcfzO0q8cPC6N6iR3sjZ5/EAIWb9+Mr0X7c028iThk7O1T
vmfimUJ93vC8ichdiR2z1mjRQEpW096iSX7avSKJ6F06GEylSScJrFlNsHo2wrHqCPrGVcs524cz
lAJk+DXcmppSrv3Dw2RQ75S2HJ/ZAgqEk6Nw52IZOAa0Q+/i+KZHaIEPVhSPjixRTMxJ5HUbUzMg
MiwOC/5Exz+ulOqE4MJp6bHCOF6NnV7Y1gMzMLCESm+FKB6kFL2dFRuztg1JxxMm4cfKMmydsTDr
yBkcrsScE7Gnp0WLVoiDmTICHDB0l81vAvd7OILjXnHNiTXUc6+v6gilikPG5yxxd2nwRhcrUSxK
GWU2i6pmj8VlXLiwww6Rd8rmg3YfZuv0KSkornYdZY3dWazaLdNUCKA0NEWxF/FD0DEcN4GDmrkB
kVyurmyszFd7VZJ1V2fqfRmkOuvX1kq9dhURkp28sB3rmdY41UYJZJutTxUlN0ysTnFEqeO6H8Aq
CauKgpkBV1tM9qctmjpezEOx8JoSNxKIGOzek1UxoyRbQ0gK6ttjZr1GsKFuxhNMHHM+MLBADr28
JsOAgBwZDj7aTFrz0MgHwXvSBNyzIBG9+VfKUNIAut9OYQBqD+UeYWA2jsO1YQQ1L5yxNcQ5Dqi6
KFE6Np489Uyl8s58ThQX8KCeR5EyOmtJw+IkBsjRzbFoQaS6QRTNCTSvIiT7rk25t1DbFKSVkZoX
lyhieuilzvnQUn5FZPctVSfC3qD6K5+QX5w576K8HAjH6ERIZOrR9Zh+nW6ulYoiw9Y7yQxRWxYm
FtACHPxP0aR3WUFl//CNmMFewBemnSDV6AzEqsFGFRGMibHAo3FuOFnnrermJSd1HZlQ1NBG2Hp2
tEkwnM0D8fN9xxeWWFThJuqwQfHs+Cb/Z9KkFasxM3pgBfRGDDuTk6oWmUYop44eYsHFxhddFz5a
zYwZ0dKhdSgjd9PS1CGnZmdL6Eh/TYjVFBF+5E8EL9AQdl/I72MWotFTmxfaKio8qOWFwJbF9YZL
fI+LP1rqzGx7HsN4YMAmHcmS/npp6MyTPXVz3sHvvlIo9pDFBaIJSVaCzMagvXBcnY4NDe8682Ag
Zez43BqOR3JbdS5NM4NamO+5MtMlY9DSt9PW3uhbv5oj8u2njMzYs4ydI6o6iS2wKJms6oa52YUW
IRNoVfVZioQgjCXUqnoLhohQFgB23gr5va4m/EbU5ns4mt+ZY1Z0U/rDs1CyZtxnISf+B64OoR3l
3OX+ojk2EfE0arSVZdXkYIYmeWaA3JgYijk50RZCbZiTWwy2yfnUG5Y0oe+4Ks0+stqu9+cB8Ubk
5v8s7GWptVA2TEyi6ua84TQBDoJr39V5fVjYZCx1v7Q4w2ji/25NkBB6SCFQ/D4K+xuu2MckuOa+
/ZuV40WX9iBT30RSH9AOMgOH8OrKw1JjlW6fEKM23cn4Tc2xd0/MLEyzEBSOMqJ7a4V1odCZvWQ+
t1IcXpizi26pGKc9jr/fSX1jQEOa0Qi6h/4AnvkzwVAWbawd97c6PKIrvqo3Kh80oe8YMobUZ7Ko
hnk03YCXBYYngEBnkxNHBeegAGz1mxHk8+yeDbdg073awy9cQdReyw2aMlrhGigz1iNd132FuYV7
Ix6QBMQv9hkYSqXks6FCtoLjrZ6Y5X/LQaDH5zEWh6cs7vivKuS7fzzBLayXZFnyL7ks6zC3YAZ8
VU2GJ2tca/P32H/x2Lu6aa3PJ/emmkyKjOlpKsynpnA6OIK6L4jwGqsSFsV7jdcQRPyt4KGCWDDn
k5hSX23OOSE3Rz6v51+Xc9U/8Gvz9KDr3/a6nQ4U+ntCbJRKp4Y0/GjQvOKfwNUU1NIFyB/tnDzU
+MZQd9tMEzul9e/TaRDf4oh1Ps6BMPp9iMIYzcn1WLBssJzR/O866CqyPZDimL2yXs1XD+tBFIyU
8NsLJljHx2LX8VHIjm+ZczgpPfUqrrXSZ9h4HiY/QSNVer1D4o9TFD0H3NrpYmtQTkPP8FfuDVPM
nrw30DVZ22R1YA5e1V2qqTW5grPF9wODWVPDTszAkrS+jRx4k9ii/Sd0OZW1PXTl/BK2w6LxU6XQ
aP+QGopUspUVL49MPqyrnVjaEMn5Rf9m+K2AQbx8QDK2vZh5sAx3JLOHzL1C6lvm00jGm38Ab2MW
CXrTtbh5Mi/aZlyNAmleaq+QegjIZpT2OBLNswperda0ebAw8Z5scfkcAeqdy1mgUfkKjU2dO/9m
JRLBkbIRRQI7cVIJtybydgbdrrB5dHR7lTl73MWhNT6iXbzphfYBG0E1NzaVHRLckB6FXaCBgOl8
YtrDie55s/lEqY15wrDAuyncOePh20uQ6+FzDnZf0vJtbMSsXFpLxZsOl8x+rIG1jk62cjP4PujL
9VHqBKiWN7OYSDbIS32Hwx8KYMSG5rlmckvfZQtjMKafZ48lYhIYZHNBCx1N5xKc+GAQU2ruqV2o
DV8qi7xUbEtCs56TuREcAnYm0kpTSk8YPVjr0OiA0fRKDISgdv4cpcJLGavIlI7T2ha44pp/K8bD
+KHNM26tdLvkL9kYB5RWGM9W8H1NpgRzkvJhVFNjoZ+LWQZQIBEzu92gMkDkG4L9zNIsYGphwWgd
xacMDRo/26CEJAFy8wQhBBNmGSPjxvAcIr1vF7fPfegmp6xQPaDmEqA2Uw0Jc1x/90+IrIzMgXOx
YoDHWtDHG/HVUnZ2vNwa1UwS1xlp76fWAP5PruD0pv45xEUIlWr3syBxpauA6ssio+KajSXzp3Pr
u4Mauhv9FMQcmtc1OxpZQbJHagAy9ZGqmN/eUBPVB/0O0pE1XQzeqWkBxJ0YABaNdhRGVL6iTJNk
R4XLyVdqiVfUkhqHZlCZIvR3Od6QUL03Ulbv5MrUBA5s2a/zw5r0A4Y3Qrk4m/DLxrcrJqSTAJcm
KIp+9D0lJASibVfmKfX7TMDWVkF3pQ1O/piwmxjUJswl2X/69UDl0tLxxR0rplX9aK6lHMWi2qCx
Sxgxxp4XcmBmOUxi7iclsSweac6F8AvmDCW2B9uCzGUsf/CdAGOLlahDO6EFMZ+RxREKaLc0kmOh
IrkvHwDfIxF6xdjeAhh1nFF6Xr7LyCGw2N4OpfWfP5S7BfXOf29obTj3ykEQmFRa/gxPHX0jPVps
h1RjNqlZJVTGLVainPVEzhF4WlbrDdFbRhP35k3zKqo4tJW8/t1tBppyZhpQY62cxyaotPIxwOnf
jEEkcBsFrd+UZQKZXaF7OH61APDF1dqBh0vndbDyNy7hqVV5DSiiq8faeGqLz35dd1L/cz4yPLMz
aktZGR4RN9b6A+SMbLyiH+5BzfaeEVEobuAgAB7WFe8PBncXGCoiPs/HYjYpqg2Vvi0MPHbSZ6VA
N1ApXY3JkIbpigoAzqBPPwYXQSM+LBOuMvDnfoIikwsv7j5NNwGWIqQT9E0Ae9A7PDPQaTOTAmuC
9mkD5g56F9jsJ825FGVO3MLhH6p1eYkjrTQwuIvacoQPdtgrXOmuwn9OLgFd7GWPVFK1ZR6v8ztt
EdbrHzogS15zt0gjvthKxD0OLxD5B5odFy4YCxUWnPl4QuG3SIXKN2Hm9dUSEyo8/33f81JVLcBR
2YHr6VsqoPD3JEADrD4dY51hr/tQexyaGHb8xbiad5+rlsSaXLQ4IKJAhDx5OVTUD7lOoGycmrHt
DYD9wnc6ejUtjAVDH/YuUSCAkUMPTwTjkpIpBBlbmETDfrDlHRA+62i6UbswiRuvxJSdvKagkUIz
lMmykEuYeqkvSIwQNpap57JJczdLGpt9OhVRWI9NIUzSV8MUXXk3R6j9jpk7Z1W10O+7yFdYFFxh
A3efUmptSsXuE+wgC++Emj1o7hHotOcKRvfuuznN3+F6NV5EpvRK64UgzH1OvLVAih2z+c/hSz2R
qEaJ87veD+Q1DedoTCN9RXDBTxbmXAZM1csDXVxacIXBjCuoRDb2N8xDfS6394oG07ugNO2hUOPR
OCaX/x7GvZ84TYaZx8ZDLjuBnnzo4umKRaVNoYUqpUvwz1wm09d8eRIQt1I0jkC96hkpGDEFW2mz
DH8kkONfyIGuHcowo071BdxB3vpzTTVhBms+eXH2W9J1tpdwUQ0CPuTnhmxJIgRPcS5XfKKfSRkY
a3LS74Kouu9h2oNnPohINXucQqu/1oe9e2yYyct9ReACHbKnaynOABtrud6U3LuNEcmtpRbx7GN3
uHv4PRlZ7rx6uIawVrHTgZopUiJ1Fl6ibflBr3LYsedzL2iDPFF36R4L0mAVyRUW1kkMSlFRTj8Q
mVbHdAJvPTK4OYYPqbDzQe9sVpgrzTG/sjaoPX8HX3Dsx5pIOivGSBoxdrRH3WSYD/kVxk4gvk35
AIzQjTjbo79Qs/IZcl1SD0DiT+G2jholzUbdCrxzhWNzeWQFOPUD1c4ZX3ZB9ozj+bPpeD8U6a2N
rSdi8j03LeHl+YzKfXB2BUID9VcZQSvbIlDMDatHDhS6vqUWyWpHZztF2yjFl7b977FTqO20vJM7
+ZXajbpSKac4pPDCWPgso/A6TL7UqAn24e4OBLpRz+WSLeU45gJggPNXwkTh8nKcDrochsGZyh/5
yoje1bj7ADyjyN2wsemy/fdBuObOIIScmwOgLAnuoSfXGyaglUKvU7PD5SNQp68SgZmUK6ekH46B
7qXYj3kB8zwLGxPo0mZmhjN3xlCS41CC5WGGqCdIN5g8PXjiE2dYElPL8DUFsat9KrPesVyz9rB5
H3LTUGLXbr5Vgv4/3/0qd7BIdRRw4kCWoV9QRc8puzmlCsnULFqrIINS6MOoXZqWlVfXFSheuAkM
x/Ao5KSrnby80hMapp1iWYgw2UXz1IwPP6eSqGhvXTGhbgrNeYQ22hmxYPTTLcTzYSHU80pwyzlV
8SXxWOJD3FBSe6bYq+pHE/dUbaiDEmAkhUpW7Op16+QSqKYR9m5HXj1BCcdAXS11G6K4blzNtrTe
XjYG3G8X7aKhnt5e6VMebliIw3Qx4V5dHtO8JQpx3o91JKjqjl/IL8ShyLOYm6jWTl3atwLdSFN1
e60CdmUtSlsQPMq5lFuITQ8zdV48z+j7nFumfKtoNgiWdTNFxLdX1tydWrMkZXO7xZBL7INNkq+3
SsofneO6MuhTzoppJvkrTjx5SDMbUj/xy6OAdDQ0R8FLieIEXRzcErndZDsdP2qjGNkMjhP2jnGU
T2lesnzJzihBTnjjt9s20ALUBNKzc8HDI+KVl+AVRrLBFtBz1CZlXn38yStdAzy8T4L/QLGETiMU
kmrK5ziEb4arAMU9WCPoXHj6qBg14fm3xWXkqQXT7Z2UHSPTcYwtrEALa1WV3ZZv1WGRu85viUoT
bkTqUXzMdX79ZGxhokPgZb4AzYDcUIkv2642OtSAoQiFzwaSlnR+5P0a/dnNf+hhaJSJRbFHyOBQ
Tyd/mdfmY75aaVSMOMHMm2/JzMzOHygZcyd9ML2W+ClMWURmhw1Oj3ZYe8w5hs5YyIWdVM2tvKfP
vmsYWYtYEb6eUkDcLZ9m8EzEK+MZGPsiSEtF37SbbqfWUVeJo0cxTczEgFLUQmF3cGEM6oIc5GFL
KXRowYImryJtyqx7D/nRokTg0PDbNu/NjUQFEQXbyqKItgGy3HJOmPVqBuZfI0ji44kd+9859ipY
nUj8LZN9bOsVNEP3sG64BpNGIVtPuOyqJgMJlsxS5KFrNx6ovje5+0MwB1vEMtBvWWM1oHEiI4wD
5wl6lHeDWez3dNYFt4RMySKyANnczZX9K+HCrhBx6h4JvNuh3M3dtuUCjWPq4/HQFpVl3LYw9Hsa
aHXAiAQwxMkuXnXsRkQ3eANYTkUde6+MgL8YT3aTPct3ulMKQ8vHAer93csTpOGzz7RdultWP80I
isYwKJTwf0h02epTpWPGMLkNQ7q+MjfyYnAvXySP+R05jBHaQoTLh4z2CGWkyTSYoQ2LosNIAyKV
FyZ1e/UfpLqIFLsnJceu7GADZcb7N6pP85DJUzq5xFCOa4O/jzRYz0L/GOniLrL8DU2rTIkIEB8t
ex47J8XSlHakvXvngP/bmpYHc1YrTuprbSp4Xs23gz/kF55RrEsf1+ufZH8+6UWuGpT37/vSJ7ap
9zX0EbMlymSLgWGWyx8DUz0NNjPoMZMeZ5uaJnKHtE1e1mHeFbV9ZMEP5n+UItPGbnb0TwciIzUb
iLYeUPzCg/dk4oB9/qNslWHwU4AtR0etxxaLJP9ckvKCgKnewQ0YuYWFre0iYGgGcH1ZxRL52lHW
1KeTCIztnvhhi3z9pq5eke5RP7ld71yXF785oR/ow/uy/xVZXA2Kd9MOO0Fq8/CQf6rUzqKAPQ+4
GZVfg+XWYQQAtvU/pQMiGkKemnJ+MsWz/6bDFneC2ZaHFSoy8C9cc0khjJ/qfNpoaoQCrAK+A7qZ
PFVRYmHQCmgUbnBpwb8tOoW/qu0r1Ikd88eNr618MWx1mt9cCx6QnQxbMYKTevq79NU77FRJ3M8x
m9Uz7JxjdRGMLNfHP9++8Bd7i8Iie7exRSdiqvawyDESWey71RzBHJc93BL32o/8Kx2z3VUAkbpQ
fJ4bLAd7531dpLzsUnhRsU1MR5b/n6ibu1Jn0+DQi7u0ItEnuR0d5mck0T3k46EBVPABpILcYLkP
Zxax0MidVbtdxtVsBHclA+YZOVX1QaNBwCOU3DvycwGJzfqctXO+vIS2H0EhmKVPB9rzfIJOPKhE
AWoN04oktWk2G/UH6+psQOTd/qiZTaX1TRkTfDVnEHxCAsJpLDuDk8C8MQZYadQqy0cA+1SpjbKX
SExBGRDvEbXMIFa1C2V8bOJsIAA6hag46iqTUc4HNA4uw5vOxvfl7YbTeK8zznh2bRdkDsAUzXUU
HlHwLAzRFrBmZNecXeEwiJAKXW2uKKfpyqkub8ZAaqvM8I1jItG9SMK/dr10VObkArppYkxRkKuX
s7hIUDVlv7vsg3fV17RaiiIAN2KpzsJbxpQw0YzVqF9cDRc/vR61RKP/aB9ReN8Tld3O5VorpZw9
eevk+eVbB4fRZVe/Ot43sgpx7e+K0GUc+XLFmgU5r4Rl8mn0gkD5t4FG8PIEWrWNsvX36PRpLiz0
5TE0f6/CCTUok+f/588Q1A4gOAYgv9HdErtGoYzAG5jiyDSJ12T9uxHy+fiTmnoQ/S3pWe3S3Az/
gTLP1ghntbdCJYNTVggFtZCzMpMH6QwWE2euDExMNJDRJWZOs3fFZXT1CqzgowHdtTlEQDyogd+j
YaB7zYUUfk1Br83lxpV5yhqUqOOWBuicQ9nR0h/e+LeycTmE7XzlZ3CQgOrHBFcF7aOFl5GH0eVL
3mey4/rZiIk/b4Oa3pID2oQUQkx+ShjdR+Dxb/zELiQE7CKjh167g/OyiZ8VfOK92i1BhopSjalY
soTeSOEDmr9NmNMukFGTNEpFYz+Von5067pCnQdrA+Fl4+aSc43eWTN0kBtm5n0iXyP5C8oJx34b
cldY/VhJ8mRtIOg+/bS+Ceu4zo+inTEC90QckhdyvJ8PJ8wTeQdeIM++ekMbeIR3sRlgRbKmgmwn
9C4ORJ5GbnSxTybez/xuSEmD3Z7XOoDnQv5xhaDzSl1Xm3BqPRoTBQRf2rdY6+IS6sbJyiM+ybpj
tcr45OzokZNWLDIX1261fQsE9op5ySd206qBMI2H/zzAO3DImZeqad7eTfcKYqbcbujssgdhMTKe
wzivvyflIZRUImiU4vC4NU0kTpMHgTTJkBcFMUShMxzcIczj9/SizcTSlj2r/Mb4FYuBP27Gh8vi
S5IthhaNIbUkKvUoHdjmw84Lo/7rvW2qqTs5Gv6hzZC93HFL2Fmurmn3CzFkgJ57TfJvV/WCVj3Y
yTEn4scozgtQeL3ulm0WRZPaRe34Vu4iuvp+RqVpZriaK/YM0Shl93paolmYENNd3h34iYDFeYk4
FB7CIh9nyswNbJI1XC58sEa559tIHU2BSqsT5sc+GjogPWReRlYBVncs/cl/uZZ0AhxNWJMFQkf8
lM70SVrMscQ8TFQtNWQO8u0ltl5KLnK9E7QcxqkaZbT0gkBAFfNh6Wlho1MimUBqM3Uix6Crvhnx
T3B/sCiSCpyWJOxOu+n/ffFvsRQW83NwBepQLBgvaKd2vQ7nqWzxHDLW3kowwDdMLUbNe4/iMPll
CNs3agrWlGqSaIPL91+5XyXbCe87b+RevPA504kZywcqjrOy4YTh8TBeYyHdeC2srM5IW06+YftX
ZOtVaLgMuNsQfB0+lJS8+JH/cM+MXKEDcYoJ0wcjUSRnZ1DGyd+2B71e3KgeknWb6Ii8JMbpJ5j7
URcf37uLYAJhLpcZLtkN3BfwP/b6gNHxNAMHls1hux2/SrKSFscwxGrlr3OSzOObO/nF3cLbm3MY
WPd5X16y5VaIEcGXx+4jl58MFeszcFmMoHkUX9K8V0V9iWLYkA+zn+SbmMiDrPuud0QQJNXjCKSH
lU6E2eNEIbXERU6txqLseyhYeAuHfOdWNt90tcdu1Cye807eSKD/7pN6ZmNwKKvT4ruSWmCL2LW7
wXNlopGgJ5uq/ES2hmSAtExQlx7GaM/wWBxHp1aA17gtNIHfSxzRK5jXwpKB2dBMPAgRctvcPu+C
vMoZ0BMxsvrlh7TsHNHkvvZ/B5MEoiMBKx4mOrKA50JfCI1BCmejoCUGRLo0pjFaQTHfEYWSeVS3
3KZgrZUIVrfd9Ahjy3624TqNcelrTJujpcpyyJtYtiVIqb2GH5fkjgunmR8c80oBFL3QuSv4p6Ui
6r9NT1yWGKy8s7qhHCJJO4KwfACUKrcHtZwu8daS/mMJ16tYUbLfz2l4WNIGrpYFawFHCRpSETqp
Kw0LfC2YSriDOSh+HLn7k8dC9P4FRJATxNJa+JDk53g8WfAl9JtauFLTeGTZ4iONU7HWxyqJnrXp
gpCm6IB8i22rLqc5sWXtgrsKTTeCOaqCJ0h2kfQgaN/XF427Kd6jERWmgQiHKusWup00TXvIoUM3
KbP35FB0Th0GKYo7ySnGSMwRUhyH95wKpD+1eAbDc++ypFZeSN84OeaAyXovIwnQg9VRa4X9BkPj
s+9768/22BkuBRDE75ccDsPSP/CgOytFnbQxTYVyTwF+4glDBG20lp/aMaIQY7VA0hBYvUpDHSS5
6/O7jseqTyCewKYq9GxoWcRaKyn6cBIPyQi56AUvoRka9vxNZgJsx6Ij7bqj6XQHMJ1ifNKv9q+i
vFsWaWkk60Xyqyx5totpSF7+VgrvFPo1x//qY9uF05Y5WJLTWw7CMv8ftKLB/EK2kTe76KLJ/CBo
bNIdpGZydI8M5RzeYcTE22lESv3/N4LYcJ1faijkrnH32pTAKWnAPAorwVj55DK5gRqafiO9e6OV
0Qo6pzbE9CaadaDUxwK/BtHqIMwBSX+zBpguDhEi/Jor49U193OgOMDV1LxN5m07gPVaUA2qOwrH
YYnnafW9WGew3SeBP+ygFLwK21r61jWilD0LfBGwakAMv51fsvzxaLU5+ffIGw8Ls1IQIJMRU9xF
lwgkq6YmPlhdRinnRWKG28uVPC1YsJEPV8mU1tsEYoOGKoxx6RQl76ZlqwmVmVklb553cnD1n+Vu
izEfyFa3RxcP+kydJJl06ssQiiij0b3GB2riByMLuFHfLx2Mtnqw8UdujrymNyYwmMfgSglxObTo
nTUK0GWqpYEmptMUTm6FdjOyK7DqtkrtUT1pDlXeeiW//+v0kwUSLlomSaY2ShVsj9+7SjpLbGg4
OcDNgrz9Q2kW7lWFQ+YPqfbJSgceF7QGTLoxpdPqs6h3NgfFPdhUs6pVTxylLLt/n7p+A/0SnNWn
L6pDbKaYWZFRRFGAclZHYmSjk9RJWVITGXHJmP5whjignWEeV36ukhSrM/IcBpkRlsa2wuNNRntT
McndE8at7Kkcd5NwSBwbfhxYjr8KyD45b6nlZm6H1cJlR1OhL970SsX247YkvCDQthPR4XubDriO
U1Q52zdWQtOMGmivJ8fIVOGjk9pZV6aWIZptNPeUWuG1NBeLOKLmhyPiQ+kWo7XVVYfdcqq89+0C
eSjBYWFpMF6tZ4RMAH1MjmKJXIadHbTF6babw17Y28+tdzvOWT1fbLQqc6FLwNgZmlVYkqa/OWLR
3AzBhqa2pqBKMm0G4dXnyayg8yAkhaMnzSsamsRyK6Q3N3et7Y9RW0+fdRfyWo5gZhRBlHGg0ngq
yv8vqlYtVhAonz3xFYDrBnUiN4TpbwkkH26TeHP7VKWaoxQZzCbED+qLZ8YCSMgXBPVgfMYFltgx
ehoz3cxy1PyTn5eqjW2O5NjJqZ4m98QIeFhoMKny71UJ+osxi1i2js9zZmTy1R1TLxNbdljZRQbi
HZBP0BcrDMSc2xPzfgxHoOj00JrQeH1CBgul5Hq4FZCoVNo3HOKp6P+Z+FRB/gO660Jp52Y9XV67
Sqw3hRT2GuOgbET251yJEwiE62TVmg0gqH/5Jtd8Edb19pHCNkRFbgfpV1oRFPkSv1Ery9GOp2EQ
w7TI1gYkfc8zaSOVQY/j2jZjnDr8AxFM+NwOQN1R7Bnieu6vtKKSz+ngtb/1FpP3Q9B3VdhcvbRt
MAn2UN3ihpRs3P5wHQbgt5V9g1itktFWKdvyQisHX3bcJFCYIlCzDTCFsFlnqa+7VVBnRKm9INxW
2qumcDEZovVZOvCmNUos9EFGs7/QFqOpqFy1i/dXmStUIspMJM6Cc5QB+OBS6r6Y/kyuj3dDA3lB
iM6UcB+bTt6y60rNWc6FJpe7QCly58uCzU/lWDb7Yu9QmfNTOv4HQNUHRFpuKfBSlN7bErXDtdb+
ikVn/Mpey8CaMuV5KjG9hL5Cckp+NMsVpR2IuV/R6mYMYdS4n8KTYvzSvzT4miX8BYp0wckfMIDM
OrYSCNB7wfV4Uc85h7Of3rvWPNRLEoKQx4JR1N+phZig+1JMq/PiSmBPiHoSVbYsmmDpBiRqtLqL
TpoA1dgyTtescdNmGItZ+aZ5CMbcriIYb4j7HAs1VS3sMAHPfWBmROilkLlX51JI8+EZ7AukzPxV
MQkJ3E43FcXnqW4uYZlt7Vibbor/igTxS60WxRpQe9An5ddoNyGFMpBiG4LR/6fGsBNzpvnhFBKp
QXpTT45fX3b9NTC6LUpATsmem54tqYrbR7TqFr49NDCiiTqDXtm8pqZ1fABdevwv4LsNmY0rrzG1
QZUr/fuZJSv5jACVarDx+7klFTpU81tOj4ADRGz3+XJTdJnPsF/5jTYV3tZs5lbm3WMuN4w8Qnr7
hrV+aasQ2uv+wpGi1t+LdKDP0XAEFK/+bIhmfUngxw7QllwuF1UHK9TOT2jIdFz6CD7AqZWS3rzU
fcrpWz4U2iDhQTu/MFSyDRjhUV5en9oe1p32J0RQHIF3clqjfbErW87CfiA50T0uig8UwMDfB+E/
m64ZZr4X++nj1TNqKVJz4Dp7O82wLvlwqDMklSwnSZRsBraG3oHc5Jmvjcy3q+ZB+pVGX4Fb0dsF
YIA6C/mjSJTC9DW2daIf2Pez6iGoz4/O/DqUBnvNkRwiMU4tuGanfSCSKOvh3HwPr8XiOUnuA8Zn
UDyKRkQpE+kJkOI8OiTXsQhn4awor3iIoF3nQcN5zn0PYe9iriLSefMIblyYUDwQ8EkD+C2d//1J
ZDzY/rG56IWBj5PzLm1MOJ2XxBz7L+JZmoj1BdQqtOpbBdNNHP/8pu2JXEfPuOoAxDe9bNKqtEVF
NF7R3rXgaz/YZtma7uetB2ENmGj6WfFug3tRj864C/hlRT7G5IsC8dGM8EX0IXtvjpFBh6DRw+QO
6jcHYO8s1HYJ2JkoAlGnX5MzHJAhKXVNJB8axyNe5K+JEr3Ge3bO+nJuCIMNaoyrOAWGSYbISXTe
srvXuiugrtmyh9+BhGxnIo593TVUIsYn4hO8HGJ/0KrMK/Dbb+lFrasljIhAG1Qh5udO63+xFtf7
Oa0Ntuskbdmw7GiVerkyMrrIY5GQ5dUWu1Pttr/5TYGL67TrkDb3NS4F7Qxku16hoYJJcpcy2XPQ
5Q+JUBSDpD8eAIvuKB8xOuW9DJaDscHj75Lk9el+yM38FniJHcdWwygFQBvEjokM0w2Jr5Q6xTWF
sxhASUrTCdDedrF/8CtUMq4rCiT4M4DK+R4jFV/t/iyhaz2nqF4FR44Ustn326OPrIHJydCKby0I
t2k8Q+lIbiCUfglZJslNMvUj9/gS5u3KJyEJpns2KJrmInbmulZUu6tHyjzQjoBE+l4L8qooOrgf
vpWlz1FOO7mRJC8bVbnDGIUYvhaRlBHTEsBKdpXGCm8evkBgVQHM3KmkjSkHKTuvu8sSkBee2bdU
mEa8sqv2LB6i5ayxaDDEqCDjgOZ1w6QwUwDs28fXjwR+DBTEjr3A7lS1NUz/0btaABpU1JwsMs48
GlpaPqpNYkkIAwnhHzMtnT+GlACeQ77O2/KCgPp+ei01Ewa/BZj75GzQnxKPwNdp8yFXk4yIndzr
iB4VvcVppy4hSm/oC2KviGXhTx+ljRKpvb5mnGq35zeYcXSOig9WHC/BK9IN+WZM1Wq0lcxO/vSZ
EdMcUOAPA2cN/4xKoJ9nqgSruGjH3WOsNkUNzNiXHNl6NwSXTqdAvKXondhupZLjxc+l35OogxJc
CDQLmzw4f6bC5WG6oTC5bCX5P2iH7hCeORFObi6gS8DpjNiIKFgGJMi4pC6WNCGxv8/+9TN7IXrK
AbiqAxpwyA9s13/Xb9YcQMcDf7jMOpSjQuqEHOgX+QvymzJA5r0Y9av0PhoIH2p8sh7bBVd4dP5Y
jzfrccNuj16aVJ7d7E3R/FPymWko8fZ5L1IoycVmIynLXuM8dLNt6P/1IcXaLGAgly+HbAIIxm9c
dJIDVjAekJiO78LBMRNrq9DzrNH1sGr99y8wQzL4obU3/iAyJJNOORRto0jyZlwKMCbFj/bFKb2Q
mDGEiyRWRL0jBNcTW7VXgsB1sd2mdSRP+tgBC24kjCsKb8m4tpWBZuv746IkEtIexOyyeodIrWgo
KIq0qJ9r5UgJAyM4CVersdt0lCJAskIg178yGC9s2RLIrlfaEliWfNrXEsnFrhViyNIPzxmcz8w0
ZoIrImMbdv371TGszLi0h6Vt8IxyV4aG8KotwtqQ8+oe+6n3NuC9naGhI0CrlwK3j/6IuEKNnI0/
h622EHC1oxVZkot26uYRIVq/R8a7kvPExJudfhotQSDt+kRryhni8sKXcKd3fFudafSnCUPMmzlp
XNyXSCwN0HgOjlEULNNQ7FrlVinIRKvsX3GXr14PT9/twm2KCCB7P8/+wP2Y2akn+DzZu5luYoug
kDXPws/o94ZmCeijYbMH+1w3svLPD1iA0Fs9s5yRLzq12xXEQufGzP3YFqGAr/cUWG/R6VqkAq4/
oVm+PPS6ulW96hEKQ3Yd+c94t/IQuyu9RM7t1IrWKnoSCURXnOKd9FCZWjWNfN9oqIVO5kfJb4yz
e8s2Ey5JvXgEF5h7dSNooYvN2Yjzds55mUkBbDoSz0glxq+i3fkCle40wobJwh8FkuSe8xJanBbi
LJXXqgnuDGBlg7Bbqpsi+jvRlUeqt2LJdxsuorySTJcCIqLEj59qUslvf4iFs6dx1e8CvKEIam14
BtCyGxr6ZWV9Y74sjIzSIAUELra1TEGcIAMU8AxEhAPcW+QqdqBFJTBRkssxmaB1/yScJINXoCkw
kcVwd3R9JuZHe21vZZxrHxlrjmRADqn4//AGu8Xw+iI8PKv5O97HXpbDLrXDS40GrJUb8fmIYRIf
KOXgGbPa27RkYYKBYZnuLRahewk/ERElDKX6SN95e3DQetCIwOlsyRBijnLBHGsYomZ4raS9q6Br
2L+4LVqjkYSko2gLa+Nbj9uSdnN+qYons6RRsSZ8x0ADu8Csh2k47bxN5n5znlDAb+MYc0bEX8Gu
TUaPlTPPoL1Txr2qJxW4Gl4IYc5W5sHh6xEBUNdT5sfQPnRPGRmrKLEYqdm5eHEtrrLEn5Z6STq2
+ucN4xaPSVfrCoMJNCkUIomA62GdL1yBjzE+5bNhBkvh6WuALms0O9bS6KfElGGH3fDVYcNJwoM8
G7O7UoVBF/LJ18wIEDDuFb1UzDqd7kuG2Se4mXrPayyQjLOekMMP7gQ+RuezTMKAXw6wVbTq8dEl
86kqjZP+jmLclrSCjsLLN0VTL8mdfxa6NB175Ikr7CCiivCDSZz/g5vA1lEseLrc5OnLImzTprAC
odjnD1oevWLprYe+FJ3aCJpaB2XzO11rnMAv9ZrXAG6UwLrPxBDmYE7hQDFyVJmHivJaDdokCX7U
S4Rmt27aY1WkU/LwUs5mO03/5FuIJijiXOw3CeXBzQnpQoaXvM9CeG0RHeEookr2s/8he4E2he1h
M5hb6NM9boTMTPt+MLlqe8fUG2gO50q4zP+sxNVfuxhSMaNuGsIfxsw+2DI0/NHOw6CAx1VtURCX
fuTyp7ico+VS8ypFS57RaWvaMVthmVp1dflR/xxrcbzo7KQFG2ZBKtnraPvB8a9qs422nIetK3wq
yOv/PogPIi0eGjzoxGesH+bVU14hG2Jgb2KbaanRHJtNDW243KCgRfmphoOjt0lChiLMJI+0kEcN
gkNKCpB81ISSu00k9d3ZiSZ5WOZMmeS8/26+1ERTPrxxj38eUfC5qFgyJuBwUhuyeFBm7iV+PQrQ
3JMGskF4erXi9ekmClGFeLinE2rbV7GxHpANCoSMy/3+tWciF/ujzvc5xUKNTzErHIuA+VI1EV21
EGnmbbmw3gYPMQAXLEOkcAc6eQwfUUVMOOtaFYlMuCQKAyL07Tlh2cj1dbUaNjrS+gLhrwjrxyuS
y9LiXq0EzKr9OdaIVRpTg6tH8Fjf1pcn+llFtAHDnuSOPgTWBecAXwBpOrggKdVAq63MIUwPwIyE
ZHujOfiZGpdomfa5xCjknrmnxpzjAexBdJonr7iNM1VnxzGN3pELUv/38pqafLD1/OPwIaGXRflf
Xrnj1sV/2W1DMs13W9kzMrSuOsj+9zM8lp/oRQjlP8+wmrPqElyHxpNyaUk8GZ1CFte91TGsCNzM
9wxWPq3PIq5ZYE+OS7KfijeteMveepW4OPiqDAdc26Z2RC01maj0RzR3HfYkiaz2zrnY0M4sBTCc
u6mpDMagzGO8iwKm+3ENW/R5RdsS+/otX8R8c4l+WrYr3+S06W2dkIOnbGCym6apx3ULX13o1z4Q
2bH0VheBN3MztV+FnrWjvd934bsnu0BB2S1LmvBGb+MhrTw3LXndCK/tCawpMvqa4DsnDnmftk9j
fq7gTACFhAf+vZriXVwc62dqw1w2j2ONxtE2hJRxGuSVtyE+n4jJJY3HOIfo5dCkDglVLX30pKGK
b+WR65arQJceEuQY0e7/Dxp3mMpvdABmPSKGpTQ4isbU4iIuGWY/OFJESblFSXp/tXDLpkpndtRE
BdMZV21eUsahin6CnzmJWz0RfPMF5Gg4Eb+sDgDRsm90ysl7oyja9hrIF7P7Xy4EbC6/BxmwlqOz
gsXEATMSpRtjoqg5cdwqWoi6e1PxxY3ZF4KZKMi988dVtpHQLljdbNo1Nut2eqV7BaMSY1vkWPfa
5qkMw/zkxZF2sNz36D0BT4U235fI2hTUiluJtOHQq961dPm+SVmQpr3SOvF8fIxr4EUDsKcVvT24
XM35Z2Krz8qtdw6dX/4PDMS+31mR1bpt6dV3NrcF95599oPqIQthxCJ33J2PWbmZmnYZLnuMqPKQ
D6N8qOFD9lPAj9UTAKHc6nlCvRS8yW4IuCHzbxXf8HRGoHo03VdrZ7RBj5C4qT6asqhWW4EVFzXr
+YcI1Gz9Xt7u0OXn53+tEtuIz4nMVnypZPidLJHqrT281sdWr8FqM9P5zDskPaTW5zsVPTozdnqu
+7+TX+hGwmMkVa798xs4KIKC+QAbaQEtQwVwV+XIUCAQDcAFBhIqUBQlnqCg4ZDgtHhfcJDuMa/h
fOhpdZK4wE59/Gmfmo++4HFzU3LizNuhdauUVlD8HdMykfV2f+D1JSU80PNfTtzJiADPn+Zp+PbH
Hel8sLdP1DpMhv++mhPYrxl1uPXHUCNCw8c+H/JrTfHsEX1cdKGcOdAssh4DaCDAMtFUGvVSdmfF
0/N9i/eiFQkofFhjR9xrF35Uz3I6zyTSGgelJkBD1Eix2HHHgqrEYXSH8JsVuvlw1OYG/NsLlQbK
YT6wUOmBk7VD3qQcDSLLCD302acLrj6toAx4H04YCEipQ9VyLGMIV8EiLOY4ljfXO5MjaKb6wdUs
Con/6BX5AVNlW7N+j0Ozq2dnDgTtEQMh2Ef51K1O5MCmuiENsv8HjGPMLt3cnQSvE/8m/VggQDSF
ttjp2BUOeFNetCx+YgMPWpSvvWZEDngXZE3aEtl/MG9Ye7g4TvuQ5q9vjd18pj8WsTdc9lMCEHUj
BmI73keRd9ZfmYyYRthNm7XzrwZuGxcxyUCJzhB0cxIHlXMyP6xr2+Thzzh2WRwWeS81Dwws0Xmh
FWpj2uLF57YZcitT4HQ8FV4Q/r3JI5db+Qlqez08Gzgr9EGHD9+91LThu9kRVfnX7XsIoyMRQ2YU
/pSUPB5/eTbJQs1z8/tKnWyN6NrPR+euG22AdaCr2M3wb4DjvZvACpbUF5VXMZ1SFStnTitS53vz
HcxH8IUmhBp9epdtB7NvPke/LaQEBHY64bMMsH99qgs79/APgM7tnepGYjoWg+MIEKF0ZrfC0Js0
foRFloWJSh3Y4329o7A3eh9GgV3+5158ZH/v4K03/YrjE5TMTSx6UcILBLlOaMQNBa8M0vKDunQj
anHyuraETfKQYsv175n6UvdXlEFOQ0jLuBimY5AWykj+vGxm0n80/3yOjuFlBfBQdgNryobX9qgk
25GU6N0bNXzGmFEhVZsiyqPwexArwqmUVyzr+VIqOprVIy/oIc7XguJ8Z+XV7PbUuiE+B+LdgDVd
vWS3FixUh2Aaud4hZcMZ9RGB8/DRbXgqhN5BQU4po7EpP7WJrpE1ElUXOxdCsuTjZbe4bSpZd6B3
tBQNLSIOvlHc3tW20yUQV6QZC4/JOpC8pcrssqetO59G35MltqfLBmkhTZPR4e1c92IuRMUAykDM
dyRMG1khkCpjqTr0geBSdA8diVo4n9aNOPyIzRqCWFjC+zBxKGJxgVebS+OGv/66e625K+8RjXqz
heTYRrEc8AZSc8RMaDm0i4lNucT47BxvcaHh7vKA41FqxJRnebDNiu488qz2W9SwEdjbTdemEUS0
Z134rfg15NqU51QDNd2HJqcbAVwK6Zhei/2/lUQSCz8t/sErAolhp5I6wHf+yQN4+yF3cQq8lOBK
TP6igDxyyXhK0+BkNSPKnMpJKV9yjmmszbQ8o84ceAT8OcR4j3h9oVwNqCSEtxc1c0k04Dhh6z2D
BYC7qiKWl6Xr1SwODBtQRmZUXm89yrvMm6Rtm2tGfVHcfrwGYX8duI8Suu2ClsIxZxd0mxbnvoz0
YSoT+X7LGpxiVB4hjPz1j1t2OHgPillM/MAI6YEucmevaeOU3UGHrX+jtVdFP3s4hMu16bItsbgo
5WyohN72WpVrcV/5b6zmjrv/heAb+A/xY+pCr3CYonwSDAh1c2BTE7x21XJlga5bxzm/648EIZaK
hdFSww8kPgCHdN1kqje3tcgv3Qg86ZQJPO5a7lfg4uQLZmhST/7d8H9VfXQmhN7rzJvGGG0wSatH
1R7ZmR2lc/rh8cTi/g/dCEBMpJaD59SKTuz+9niMONL0zAXF1oTazwrBeFEn7Pk5IBto8T6GHzf8
qcTaHJ+u3erkT1yS9YCPcK6w8tHHpVViJxJwxmFl46Gd/NIToDLwMUwiQYS9dImET66xobY/3gSR
E1VAHJaUy9yyPuk7QSm1vTsnfsf4xR6xAZmEaBIbfN6UnWy0z3GlUAIv1OKbtZrw4M6u0E7piXgS
BWOrScotnTXBGBYcqA8h/vwUyAgzv1oGucWIxztaRyf8smSszVxE4nV4QX8vt1j0oCxNBOeF6QNk
QA91GAs7IPQrYB26DNgo8aguTDZxaM80qRuSw/yeov0RhUGuhgxHIScT+KGb2+tfSkAA+MEowIhS
BGPYqUcvXXS9FlyEfBHSUvvlcjXYpa/ZCCPKqvH9bR5bXlunG4p21PEmQTjv+WSgK2nHd8Y9ysOR
YKbNv8Wsm9w3NqHRgjGxP22p+3EmrJpRKawrN7uQvyh4v+t7Cxog8i+d9b63q/Z9BJP9IE4JogkM
wtoTmoqlvl7cJInqmfy1GvASXaMtsELAmsIA8W8lzjVZAbWZONAVwtTrSkxPypaaVmo7HRTtg4dd
GYzMdO25v2fUC3W7FjAD5pydPGdISHquRCeejwlkqVdeJ28pjvvudbjAYFnlZWbaZjqX2Ft9x+8p
rtn7eZ4py6hg//KPayR1N0oFpKAO73wsOItM505YPY/lkGtxcbvKYcDLvC42SobMGNeNrUSbybpL
JFApFkItpUCH8EJZeWuaMJMe/YHv18Kx2PHmpIuPhtZBPWWgNe9wFg7az8XxFTX2I0xLzgpSIXMt
GfC1JzBzioaQxlz07m9xPHc6mvPdecEE44qvYRIcuNhMGkPkPWY5+GKOvsKfxmkZWAQ+FhQHRiJJ
ypZO4GQwPSureA7XQKAxkhhCLFkLHdgQjvSTDWNh2IJKCW98gnVavx8wZcw6iuMidwB0/UE8/D0G
Eqy0IUwjSRkRG+dKnb0OGdqSwwMgo6jVz+TMlC6PhDbH+3JGLNN8H1CGHP+sRMJ+AFFS6NuSBOYr
c81dVdk1Z4zJZwRTVB7j3lpZzfOeRsF2yfiu5229ajEH7xJym6yVKvJG9LKMbmw8APkRbRaqOZC/
boj9fE4BdJ4sArHmR1p4VY7XLjH5oB/RdQSGd5kYf3o8XaVozklFmURz3hg/182DUElYFJrWyAwi
TJSN8i52QDPX1pVvst6yivGTZEH8oGoPT27Ug6eDz04dRVmcLNweINeQHS7rA39UeOgMujJLjtVJ
3utTcjvKYdJ2T5RUeaWap4x2Su3lJjrmiFEcqTJ6pWEPYdpvOHer8gkZlrBtuG8WkF/QPqFXXsdH
5S7lOMpJopQU/wFUCkkFxfX2SNbhQDfR7+1wigatbTKAHnPea6k+LQgLHk7Z8k1lvAvt3MEJ5MWn
9fQDFCb8Fe+Fk61hnLyjZ+DRzBwh3cAHHVpvk89+sNJxO5GJtwQCTJcDZv5Yi5zpPecsPVcTixxP
vCzlr8/qcOCIkHN3Bs3PvzD0evrbyFZuDD8Evk2NJ892XnpuAqe4aQ5+Hg8xyArQ6Ccc8RPe5Cwc
oHbKzqvo6zkZ4uGThrSVrtBrcKIqe6aiFYULyB4WZKDHAR08aPUAQDJtzBZ60t89SH3dAB49OKso
i7RZW6CeklGKLk2Y4rCM7KnXR7fNuUdtbQYJZ7r2fbO4ASflByHDWtS1AiHSs0ZpqaqNgNev/7s/
nncG3AH6ChZrLCp2u/F5/8Eh1LNnsBooeYwYMJGK9S4IkTNOIVox4ucqnM1XBg7U8znvxtLnfy8v
S+uCMWoR+PC9xOyFdD3k7mpFQyAIl9fjf9HORGFZqlM8V+/tlnccuajoB9FHRgbvVJTGsUHJRWXJ
aAhhApLL3JNg5xBL0F7EughJEGO7eI48/8JH7YPlzHNYNYQDeY34CVo+enE4v2saPNlyxexOVS1J
hfiubyBZXrfATm+6Wz8OGvn+6ZO7oiBqMtlX42GivwBjhrc+Jw1QcOKUjgyiYkjv8OkAvla1rXgZ
pZrS48p81dLJhA6/k2NLvaUeZLspPBZg8t7uuCPDq2ONFzgM+1iZZlVMQPQqHx3bGWZLvGn5vwLt
s/KyJb3VSyBXCYqQbWyIA9lpNKjW/LIGhj7pk1mpjIgrjxLQT2kgZH2X2fW2N4HX8r41zLQ2sYOS
urGX7zSndD7nYjwD03prMnC80M6IiVG/yvLodBKvSgyVOzX7FG+7JTsBmVI4bpzHViUnYcOkzbq8
sHpopsVdPqmHITazlilwrflkau+OI1odM1heyDa2Cn+o31jHpUcTlNiMJEahHLDOmhqRa08lyJyV
QH5lRRkbx+jAIcS/Ic/+XQGm+zuTX4i05RnEWrtn7rH1wBpeKwTCc0DTpihcvHPEuxl4cDyhvbJB
bpMDCA9Q5wl2Bh8Yiv2jTUA2d3PUhUHbDqk6gqatObUL0XreTMN7vsVTgHn2jDhTVxTdLxzcwA3Y
Lb67QOvGRssUX7hz26VazP5pHU9HRs/MxbKigfeD6GYEmcSGAVFR3RQYT0vjoM/O9ojyWqK78aOW
lh8P1//Bg8KteefYHUrbRMoFB3ZzrXCRvrNEdQECkQyXldivji+sVrmbTIeW4zSeL9+qrXXALPLS
IXlF0QFtB/Iakxlbse1fIEfUzBdR6Ow0kpDimg4ZKTHMNq+jo0+hWy+FYxRT7AHw08Nc63+ubw3B
+vfK/Nfpqq48oAxL5VR4o1WNGiPkCWA5FWSrIanhPFC1KrpPyQx9lT46Tya/YRVdN8q+WpayYzZa
S9uBjpXLmnMT2h6uOjBaX15K1vlEowsq330e9lzcSXYslDuQW9LTB+CGcIbQfkjJ6awMyGTj8rNc
G7YiQd3jly0mAmBqMVe+xr4Yny6Vcpmduh18gUMboykPLZlSevKkRhGwaZguYthvYeITFOAdBd8b
bM2WfOFGXo5l7Kd2hKk0QLPW9AtjjhavBisBweoZXw1aZUtu3uZvl7ssFVaKiiPfuIwdsWU628oO
/OkOX4CW2TCozW5GSWQq9BHBIjsfvGU8ITfWkUytW4LFUZ8JbKy9kRGs0RMfTiXgrL6wsb0Fblaf
yAA4MlhWV1E1B+VtVrk/zhQhDeUAW++znKLAapbCq8H+JH7t0KAuHb29IRQt2mNpw1h4ANw08f02
/e36Hyko71RwAkjKvrF9fYIZIkXr50lzwzmEVgbvKPFGJGU90ybjnGqrx2q9WpCerFUyeIKyB/JN
jRdXPrgxszxtX9DvNhCwjETMQ56p6z6GA8q8WV3GEzwzKqD2vJYuH3imZLRh2UYF7r8RoG5REZLD
FO3xZvvuv1euehsfhaMRX+xcjaBQmVi3cF11MXHZpgtyRYiXea63MxTpA9Z9bUmrHe2BZAA5K1tb
kDBINVKV1ZdxL1Y6pqjLZAdFkagQd6o/FDGWat2GZ9kr5BuSg3yLpakum11wkXUXh8d67eQM3sOs
56Xl0aK14AYKG/oaUaUiQRwHYN5+Ihn8YgnGyumA7yeH+fcu5uelqICy3866xNvwQkWsMJeEXKLE
cvWKoW9TqHUCiHtgSVy1MTGU5OtlAzimozBJEGXE8k0whSKnpq2Ak18Gq88VXinYuDj25mqRJNJp
zm7SC6p3jWn7XUqxfZhbUFqMtgkbnpti4dg4SmkSM+KhOhWK48EoGZ1clVUP5ckuspYEltaSFTMp
amxS211eAu+reOr1ZMcaanURln9wT3KvP2rgDgm1pOrKTRbJ8m1cRrtvRLUtVDq1LWP0dmbWWnDv
04xy8WG337qSvO3IED0Xb/dokuRkAn9EfnXwSHjHTsGWogssm7yjnapmVWfDLkwOEUa8nzjUyglD
ZjtcAKKc0VHyyeVAY9pL66OmAMgBRUIDqkq5jbHZU1zYeY6jzzuGjd51Sj55ArkQuKJy8y1ORO0i
cuZ+GmLqjK9iW8geSATpehFGxPBGYorj1p0+58NBNKtoGkZLh7kfpTVEjXZymqKhUk3+NL/8S4oA
za1+L4gmJebNaBWirl0Wx5g7rgIwTKGtupJMtjakG+TXiS6lRaM7ShsKs3Efj9c4I9G26wU32AhS
YRWEqH0P9uj92LSIys9LQ2Vi/3oJdSBMGS85bFFZ14zgj4eGfo7N++/9oUAhi6BpLmrncYj2Ple0
tY3ogjVRXpvIZTHtYsPaP4yAoXGNq/fq4j7eoVCotXYPdyoz4Ml2LeWJyQU0PaQt0S4knd78WsML
CIhvqij5BgkLy9zwP/flv5mMr85hl2mudcLYFwDOD2fua3I61K7Pmd7POO+7a9gcV7hWwIiPJIBr
3F7aeW69ypfiX5bCNLYijhGaOUIgnThiGsPv3PjpUqTcWHqHnMYGuq1dgUbigEhj1oUQrSy9Udlw
YJxdP/s4iY8CowrQJJrI1YJCFUaACHX8d3M8DET7ZK0jPQJx2h2mwzxWYh9N+d5P8flyWeh8cP0e
gXvWyhEBItYehZdMVg1XBpfV3e++zy8/36VoFpnqV6Fx1FxCRIrhcRKk//PFBn4KPc73fFAfTgqZ
ZluaT5Lp02PPvLCo99xtaVoXW509/+Q1rRTubTDmLrW0mXidiAuGCDGOiah70bNS//ReWhIFk7fq
dlCgFZr0JT1Xd91Lu4wrTzG4CS92SoxBZf1fOgH3JJZZ0vP2kXjd8plCSrPNz8/Z+cEA/YH2jc7t
+7k0N8wVQkd2E2Q2o+dCjTucnjJQ+OWYRQuIDVe/Md5LDXEjEkX+Fan3QTyMrWpL28DfmtMOsOgE
7fX0RarwKMtLoYwM+vmq+K7ZvchPsv+c35J+uOKMHRKIaxI5SyS3lR/KAMpoXp45yOqbL8k2GzPx
J/le+Ndvpr+gUae7FOOc53LW2NxfFYAVrYd6Eh9ddA4+TRzxPyJe1BcOJjPq7JqVprg3IvHzHWs3
0MWSeehYiNoMxgsewzyushJ7BEUQLNbDQs1DKG9UUEUbXPcsgS3sfz44Ox8yQoaRYu4ZxmZEwBNz
mOjCSiV41MmP6ycNhiNU7BFHGhScjGaCOWf5PhX52M+7BQRR0UhgHyoJelLzXbDohnvLMv5roHEt
SVjIUTdSqL77ckZe6DQ/vvDfwUpPw3XsZCMh2jP4xtlZ9BeFD6jaXNRRYjk/Q3qJ53v5hlQY9DJA
EsN/R/n6HzAFEggWc/CGWVjcMvbd/pkuSiJZ1IKFMPwIliwr999w5ILJVUVh0fMxlisVkLsJ+DgI
cpzcwd9w68XjlVtRpuyQtW2RZTtM3xxFoS9O3oPmK0vZ0jdMsotQlHuTY5FkSgLmyogmfH8PU+8x
QZ9m+Y4ilAWaMXbR9yRiuM7dY8crObtt+QcZc6Fd+rWZjLteRzD74khs/5fjQ34wCumzxp30Tk9g
FiFwat8tGuXe+JCbZOa/AO9K/iblRHX6tg1b3R3R+N80712K2cXQ5GRIcnG+8z99D3PLfrrIzW9F
PxFXIGbvGyau9yHCCjoTPJsJ0Edy3HPkJweeLRwRfT4bjTbO2knHgBaSlC0AYLLuGl5qb1blRGMh
fLqIWPrprROi37itH5bejRnBUBxU3v+lWlJIDqcH5pWKvPOrpKPLVxil7UGoH5yUg3hcqZOKsNj1
KrHDoIx28FOxKEITzgFNnxX1YCRsg03sUCNL4H1vK69WAtat/7DJUGPZaSeSCF9i94Vtv7x+3Sga
aucxYGp26f70Fqpq8jJMx9fRGKHAiCrtwdTSgnsEr3vDYGRlK8JzlxR5PCSdwoA4FM6tayyeyoiP
B6bj+ne6duny0jVhEm8l3Mp1thYt4XDObLnRE/oY7G7k5aw1g4o3kZTOSSyTwulNOtYHg6BLzkbi
LqktI8vS+LvlLgz6inctrP45pMpdxTF25vsM5XKVE0y182BGtkQiva6yIiuaXWIWUY8zwXGf9tWY
BaWuOPxHfNSRkOyJINwaci0bG9Z4S9K6wb/lgYtToICI1JeK5aoFiJXmtriguV/qvETstXGkM2kA
dFcp5Pak30AFNVStACwE4bWsM28CWOOQOwAnXJ9Y2RckSgwT0jOQOeP1ILeuMa+LKJLW+Y90gLV4
RDikeCWV2LYi91egPaVwFKZeYabXIBYauQDebPRDTelsAsVjmi/CNBo582D5ZxUZWS/GbcGOyk8l
9xPJqmjpsC9+7mPaLv778Y7Uz2c16rJ2qUfIT0Fi96WwXcUG6T7CAtz8BlyafGrZMvl5wH6FxkHZ
pnh+xF8vJKQ5bcw/rXCWxSzootrIVOj76WSAkQe1/hUDfub2M/ywXQBwBQTdg5XWCcQtST7HzdDO
rW5gzBTwtsWkCr33Y2Lud9eETzs4z2l9qRQMZzWmD4El1r++ZV5Dqg0Harzx3vTWFLFU2b/RKh/S
cWqI0ET74AiNKiBvjDHqYcjBz9bEKAQG6W3c76YDTYy6zFMWfO04Cw2Xm/Z9nccRAbtGZQXgY1Di
hTyjzC837e14Mv8S+OC8pI/UkLe7xL8fhNTD6O32SDh4jGUz6CzBdwa6HA7q0E15d55SUN1vtDhz
I5pH4sxAbbAoGASSQWF+7ceXiegXY0OUlxBFW+rCbEp/AG+zZOHlpb4MNXSk7MkloM932Bz1CKF0
PiIoa0eUP58RlKjPxNuL59BRoSXhTgd1Ouxg4F8AirV6D1v4suWaiWEoE/RSUTfL3skRJWHd99GQ
cgfjDjSKXqpnMzeMx9ZSGDkbZ9/a7nyYNKUQAyU1jz00YAa5j9v9UzEnbnHenjkljx0Eop7YgUcc
a3L5wKpP46/QNJoiN1LLzyn4C92V1DNOTw8KX33K9PN9cECSiGhEr/gfNc0heol0JI601M4lOgsy
z9Pl3Fqo4ZluMGerpOnArxHQa6CgVu9kWum37eJ0rXsDf4z6HQp/3HLuaY1XYgY1nblC1WiSEmWg
lblz0g6uEqiMWvVxikCdTGca5az13ByTewyTaIgQUZ7iJHnO+Y/w582r6H82YRKxKLGfAx0xhlAV
/2CpgPTMZgIcfKUmML7ouR6wTIF5IA5iivn9SlkIxXwW5i2Istw0QuLMHjQDupgs5IwQNrlRrY7i
0jkPhTd78TxbJI6zxUItUhsG4PjO2Hzpn3EWeOG+wmHZapvmfPKtetmjgqqpXgprK294O0QpCSBi
gNNlRrhCsmVnhS5e2bE6u2SGwHLvIo1YGJNV4/5GbOHSsBfkjiBSR5aM0/Q3frpmPyLXhxl+CZzi
3WjaNDIY+VlA+6UNdpEezVlYY8exWPqVthSzrmXaQ2mXCcCwZ+4SicxhRqJVLJ7SbJKfQaJrFzPC
c3n3ICJSKPvbnh9MNVGHX6JLLP2MmsX/yvPhFsPoUZZK9xYGWv8f6me61CSO0stAA1FxojfvWAIF
1HAFFLwNRoYm06fRmmGr6NfEppSc5iFSvViWYzk9/QzdxFtQ92oR6CN5xRI8ew+sy36fFhBHcYh1
1sYnXaYAhhqDbS+t1J6qQlvydn0s5hh8jBVYWjLhQIij1hjgaUHJxzr//6NcRTKbErgjlh+lf7R9
Vo29Q6gIeqo9kNFiSW21776oSE5g93KOn0WLQhs34s8NxKBONmdGlBc0uxA73Xy49w3C+BrIjTg1
2dsSkfUa8BG+7bprViPXHUsaIUx0I4KdNOVdRNvwpjXeAuP/oBFMnFNIAf07qyCHQ6QjrpOmzXMb
josmK1fQSlNZkYmPCKuo4wTxh3dyNh6wxPdV7YoUkXSNCZUPDDF4p2aCL5Jnu9gb7mTUDcI+ltYm
ejGQBnYX1W7VHwmd/5M7GcisrQ8/oY6nCz6M8HKx7Pp+/8uXLN5hgxWfWptdMaNYRkO45K5Rf9dz
E/9NLVF5AxM41YkPwqJNzVMKPkFKs5AOFa8yM/NkVmXy8ZHvJDJeLXR6fcqMxPZAh55ILK96GydI
L20QWjd/EGgadNUtj4hsv07NjJwSYJx4wJrS/FrV2seg/G3kYREa2mU/LBtplik1mOusPVj96UHI
Pv6qQUIg6E4aoIAQ15erZQ+Z0Ayk8HZD6hFpt5cH0lbs8qiNZjmrhIe6zQh7i6aSl945p/6P9UGB
WBki0GKKBOwyPBUfj2rr0YdvqhFDmULKb/jxV1iDQFkqhklTRhvNKfoZ0yyuGjvdIT02XN3cUDZZ
gIg6NO3J33iqTgIg+a/uGy+GKQBim2VPHE7PwM3wC8DcgY6K+wqNvy8PedG/kyECHLw65lsFbRvh
w/MLBTX6n+rQUUKtHz74ACWePOy0FxSBBclelxx/4oK8dFsbqTYvJxK5KqSmpYIwGvKqKfy3C7ur
XjD2ZnLWMuKmGq10CHBjg6wqb1zLKpT4NPmC2CpL+BlY6y2/9+ZaKWyY6Ntnne5reCFhc586J+Of
cHQsERPxy4J4MKxuAEZ7ysGp3LKePT+Ur/AmXqvMH9QFr0G+p3BVjmaXQ9NIdija0tLlaVO7yK64
KkPhVffoqRad6iiHGJFsNAWOzAISR3/L4NitZqyVrw4FnfKCT9E2aVSsW5QJOiuOB/GRRBXaORl6
x4U1bSfhOoMNuHPK/OCyRtmQfqNGEunycxs9oe0hUA+KP7X7SNin5AQxhwAk0KdwHqkFI0cjuVAd
+l/eCBuTEDV6nFv7kUNVSxYzMLI5rb9XOoSiDSqyb3yIn86MIMZ6U3tC3kH9lWXVLbof8TxjpPWd
Sm+cBURq0y3+YWcX87cNWxwtO29bXTdnER76lWk5VDQ1+a7HhGHYBVqJYdQbzde9Wjn7JQ0kH3T3
J4/MBoISVUwibVNNAhZ2X7Q57v9i7ZsVX5hVCMrgjwJE7bTWJVyilFvYqSow9b2djflVZoG9+8Pj
bfUjhNNjmT9Yt5zcyEYX28bIaaHxFcZuuGbPustH8syZp3oA/qqTAB/VitfrfhRk9F9woBTZbeh4
kvxNTg0wWbEUxXu7gSOFm8buE0SCqf8ihGPS4o9acz6HrNs69sbsZWk7Ynu22bqKneaTDOmnM+jP
6vLuAao8fE9LnOHMyjEhH9pbLI5jZ1U0cEu/lJUCvrtk+zMebxvWNpL73I3St8snl5XTq7wZQWyL
IZYmVwgfazfaHjChbrg2u6BqGV4gYhSm0siaQsTCMXUspOvo37qQ3dlOgUuuUW/Nz9hsZgIGgBRi
ZpbBYF3JIZk0NSKxnFwBOxdV6dfD/NH/A46maN0Eyh8nIpBq5c6MtaJ4CegEGNOLQJmJeP1bqyLt
y3d++Uc5ZaYtQfHoTThrZJL4dZv15ZpqVCL+vMTuUCN01Ze6VzzjDW/YJm7WHfIhayrIDEMWw2jw
ThLdsGikMLhqbktKNtL+ir1Z393XFd9Ulhc9/sD0nVHU61fHADSWp0Df/rsXmIzhv0QfamVYgAvk
6xKhEi9iTBtgxjRaNFyXDBpiI1/pK/Q5ZXQ0mmmFYN794QVUUAYhfqraS6Rk45PFlHcLDTCmyJqR
vXPSXwtBK1vVOuTwByeQuWozpdMDMbJ7/enjQ9GVjFOp5MHGKhgAHcJ1nar9/GsvPVV5Yv9Y5hCA
SaSJrGKVq09nTW2dUfNPIDc607IcExy+ANoBErETKk/KBp8Naa4pIBIv/8LjGVWcPpSksEMd/iAg
/sPMB6hIV9Afa05C0ZT7rUIRewfdkUJP2qRbYBOgBnDyLf7FIZoetcp7QVczBUJDemZwDyhMGnNc
dlPx8bMxbvqgp25HRTLbDsk9WeLx2nc6lbBnK0SeMtPx8M2PhRdsDWYB9aaXGGx4QKGbSec+mWyD
Ej5+j+jCNTVBfjaE2r89CO3kdWeIfpX4Ce4+ZIvg7n9iI2Rs6iqmm7JtKb6G1cE2L9h89qAs1TPD
4vQDciMLgkjYce6Xien3S39J13vMtER2ovvZEzlu+1+KeCQSXf162EenwkustNwO3q/FkOX1m0nB
YNVhvJRW+JNG1IKMly4JQmd3LdSD+o9Wg82ezRGjBHD8JFT0T8F9j7IXgpX+6mBOER9ek9Ueuxbq
UjpcaGXT+y8DjUPyL5TL8IvYlp8vAhMjErGDIWQFC2YCGAzTmEQDabs1sDHSdmMQ5SankjLvMi1w
Z2ytWKkYXKe+B90kcwD7Nx3QEutikJx+XJ+iVbmfDcGR1x69DcsbkI24YOCsJaqfGnfurCkow6Hz
5CGXF6Zw1ir8wsJWcBvOTOoLuFvu3l5QqV6dxRwOKbTZh5FcjXNDiIh1st5rk1C2vcpiGQfGXMYD
gdYNvAVw6cxbczuqt9CHrOog8EyynEkLnDhsvZwk79ug79VQvpKpqVNMsaCbcweqDprMhsVG6Zgz
M/dGMLbgSsj6rF7dDBcBacGHGKqSmqFj4lERLwI2khTSVqn1YXRJ2VKP9GJMqnWiE2FHB+IK45qd
owN8rPrWyP0zeYdN54S5TQVg4Jg2bE2qKuRz8DEcmwZMgdtRODeIq/Jnz3Z3J/3Ws4/L+Hy1hDmf
fF0AOe1MSOqzowKBEvr7gbRU6tZJ08X5uO5EJ5SMUlf8mYcatBoBvV43tWpnpEwSusPP4a96mmwT
rjKagpRjQ136KSYkxd2jcmFlx8Sjsp78tygy53Ep8ngxpxX0+JgDloWHwjudQmIWWoPjWDkUABsH
XnLARehAAL6zxkukMTSTGxjVnFhqq6OnGw6jHqc8ZC8YY0wHs29TTvmqWaAkJ0H7o2JeHLuX0MTp
Q+YbnKYHQOPkN6MD/FfZvzOF9Dez27ZkSxG3NIKzf2GnsXL2o12COkvILitlYMoSd2iPEt0qRsWC
BAJC1uWpFpq37CFW2bx6QvFl0ftcMA+2peYO2gb3Ecr2eXRUPYI7+3mU+McXmmmtj7iBfN/grXcA
ITkuGCFRL04VafTWPSQyRouO6CnOw7+mvSuAEwxzTrv0YoDuhUto/u6lP7QpmVhUz7GRx5wNv89D
JnrUK7SoSChm16pdCDnsU2EL8DvO4KCQLqShlA88znXw5sBs9jXX0YX/nOtHbX1Nn7OoG9QWzFIt
+ecWd+XDyAR7mvi2qC/aXADOHh4d5GXi+awZZmhyMfdUtiGgq0bxSUxXDkd8nWZDVx/qDuAQbxv/
lnHJd+qzLYY7nKYRsCcll5BbIbEYanGyasknUIOhtXc22JC/yEjt1NslQnyZ8+wnbPH/cuqECqlX
NmM57wIeYVZEFiT3u6i3E7AeqLYCVtf9JzlsncnENahGUXRZvgtZ75BWzsKoTA9szz2J5KMUVfCA
XP2Dcse7YIRWkjczVMxXOb2dxDflrRx2882yYGed72tVhvHtPM6qHS2oqdPJZzK8+xVTHKRnGUd0
4PBMZDvjs8HpbHwvAiIKsmQUp1IUyeh+YCpDTuaKHGBQ2CzRbexR960+nP7dOmDboCdNQ6LIe3Ic
q/BMpGUq4aWCNSHym+vbChWG4ZORYE5ZOlbHvgKjtGj8zxLSI+1P5QIDjd15NbZLJPZCKCwpKR47
uahmaHvBLJdgb21rp5KA+Gk+9PGsznwsWglTAKT+0cTtZ9FC5VaCj7aeP1uwxWwoJIBeJJ6gHT8B
Zux99N9BXOV8U2G2z4oyRuRXotxRy8Y7/nhII/Xyq9bQHnRyeVO9PK0XprvYHFAHhKG1K+Z3SJJ+
EPcGaybJkH+KkLr08prLZp75qOlNLQgZ2SM92gxV/6zkqUciczbujDS4dq10TfDcoZ5mtrWCehHr
8q3iBS+ZrRAJZxa+Qn5bKbvngnxAZMYv0eBwMNoxpx8lWAz5Rv7LS6p03D8mxO6ixlr09L15thfh
H52dAcjooN8V8g30LXiCFJXaALEY8DukfPSz6/DpB1FTNH0l7EoD6z0xDA8JMEAVwhn9tzMxDfpS
UAG7dykny74AUL6cAaD2Z9WauNNhmDA5w6SyltB7tdTodRvHmJKCkB8A4KSeO3YTNiiN+BA57+Wj
Dd8JA7+EDLdwV+3v8WvCu/wnRmLLy99WbWLPYOCgILkNA46Dr9AmY7B1p8TNLcOrHtBM4RTpiu2E
a3FTCMolWK5I8IjcR0i+m/6QpkVPry1EWn4QoHBe6hkD71pWB475Iv+EQz8ZMDQBiHoAGOfZXW3x
TbdxIRjWXLiqwjwqx869uYggVZusteSy3R7UK+IcPbrTlUNkueasxtDZoywzMV63NUP+IEOEj7nM
V5jCxJprL5zR7yzQranebZFOXvElgUyTZ4n8RMQXAKo3ODWTreUsgTinft+MvgSStji4glGDBRMy
H106AQ0gGFbAPelf85vvtXYINCrADWr7DOKMe0K6nXH+Qzit35c2t51LM6d/oZj6lfWdGsEwNj4R
ne9iSQ8CgiJiXAp7mw0bJktcMpLxVdEBzHCxsUblS9x+465fjTg+CFaK8Up0+6xD7t6AvRvoKU0M
rfQmBLa9Abf53O6UR1cUpxj1qorbO5OE3/qlQU4yCRRCYk/4okZtCzDVvq46V3h4JSpyktE3/hBU
EYFCxR9NXXiwMEffX22R79h5n1mIqiwP+9TmOpfNfRCl30xz18wQnDZmdObQrlGTLo+pP8nhlL9B
PUqqOJhhneyd4ASUOuXpEYzXrhFoD299KxT4TwS/rG6MOGbnXYE3gLxJVmAi2nvhJVyoXVqny7A6
jP9gNBSH5CQJ2zFV8CEnijXB5potsRr0ULqSAbhCNxye1vsKYXUBqrSVNCIG8K5Gwd8mYJlwRsSZ
E6SDpur4iUgJ3Prx66hPNMTOidmX9PUsHWIT2cCm6FovVIlfj+NVmksoOvATj4Iu4TgwDk5sMEh/
Q4sYFiopyj4WHHTK6mlq+O7AYrvwvjiJXyl2DeMCblk8iMt+o1CbVlTVEW7KuNe6VY+DcXHkxuP2
oF3obXkLWDA9M0t2HD85Y23ra1fKheX/bYdmWy2ZsIZWtfnpGE5A0RJYvDppLBhUqZdYz9280Znq
wxkw5YM5sCjA1mROGsMzo1Zq897KS7b+PLBaHJKQWGMBmudjWUYX2IVeuEh6HCSOa9+hQwjlFE5+
B7nPqkpui8WcAUe2+njpQ7JmpJpmUhAYDmd3M+I8Sd4LNrdU7k1tvaqwoMgGl7FnS6sZzYO08HFz
NZ4Kkye+Z54UMMnbTzhaZ+infOBDeXDpGUFagxP1JiNXeXL5csvx7Rscoec50xYNc3NKOlav8g1z
/RNcY0qkJ78iSt/OqqAqSz/oUpo5ZmdYM0JHmDT15ZozgSS5CgHpqrK5N3plwfctdzwWiZ4rzvL2
Ab5iOiU1bcB+TlVdtRpm54i6vW47hEKAWAQgUPYPT5OBYMZ0IbwR0qYjc1w4+FSOU+y4i7gJ7Vhk
6NGNQkur0noc7wY1SbnAbzS2tmxKeXW4elIBg6YPD3tquhpec6VOnyWylrUeUJL73wjofWXvQg6l
CsvkSi2ODC5k1WYLkNmadb5um19e7FgP4wqAYs9glXX7h4iQaES5Wi8MEfTxocUQFf9ltU1P0mKX
4YmAEtgiBylY93yh8nQROQ+V1eojtM9549MzTUFJPglneJMU0qyWzNs1TnZeH2f0Nlz2PHBC6Wmp
MMzUu7zGWdUOJHoHnVjgqFbYZfpALrr59HkwJEnUTAbZFZ7GkdfrWl0lzKlU9VDRlFKIEnQzK6l6
7IflEb3vQ1d3/bnT2mKdFRjv9nzuHPGCvk8Rl11de8aFZ30vzpsYWkYH5Z9ckc9H3AKEdI+XzjIF
xKWKctMloNxUhuBsteNvQhVcYxyxVlAJHMQqLerz6Dow0020dw13qCP3FNz7I9+oCtFmVBHUFXd0
888yTXNUL4w32iWw/6gZ4bzoylKsZ3q5AAf2yrLwy22qbNHJKpdbonA4OIQy7wFaLeQv0keZqw8H
Ny8mYtZ3/AMryIAZDXCIBRPrdcbI/JbXeWELiibrA0UKk7whpwrNGGfoG6+ld7SBUXmw9gh6mCEz
6yVlQAHrl3Ra0O1AKVclEG2nHAefpZx7/yCaQzeq69pABOCPQixQHps36IvF+VKB40xTNPKoee3k
I5AkkCJpXE6R2n/SL9NvvU8SeZyeU/zQhIuuxpmJnL3tyXAsOMzd9ZvKoY3bMj+mYIhGDLBs7xWK
/5Xm0J5H2ABZL5Xg+gQDp4Ilyb8FutXAJ22JEInAEb0tSrSgiRKdtYvQ88FaAIiuHYBeF/KoNou9
HaMxvJx7O2U/sCzcolgtTvBmZwMBByqSZO6RnkhTksQTUKznn+VKlTuDIfyYaEVT0RVEC/iSVt57
k0jkYNbQw7KWVCF2NY8BkF0rLeYljKD6YJQnLq6YO7xudhYRilCggs5TsUPJeeQiaTbcHLvsp1T2
Ao1Uv0JZF8UvWdImuWzq25/TkvkWtE8TOAUCCrG/FNFrsSwnFxWOCYq963jxAGsGtjE3ePUHE6Ph
l0CwDgtly/w+BpdEVP5x/KUUFdwXZqmV0GVij8anIQ/j87cqDq9fnMu0N9pmpW7X56YjkGz+Zi1N
qcZBm/r+NP2EmYbFAlP4m3ZyUj+SClIHW3/LJfPQUbqpzMUKSuVwebshtP094LaHEqqmtNQVAMdB
pGAkqw3k0ZeMIFtoZ45YAxWGpykomv5HGNQxC6hIWBLLWsz1qYrZBRaWkTbw1/zuAnuKf92J9dTC
ptWlWSGgdrjEfuyEIZcQGBDg5HL/DJFyPxhPqMFck1/uztNxBajHP8qqB///R72IdTIhBYZ2cUMT
27oQjhDLUsaHiFq24SxYgyGoUT6uCHpkupBTitR9fHCdcsTItBIGyOVKRfVw1Y+v9SEMmhZCOGBb
rvUpVC0JS3JjRZRaucXBCIVGJ8BENBAUVvkWP4JZ1ZhugeocXm+SporbsG3r5ksWX1M++9iwQhFd
QuAaIi91mjDxCGYcmMR4SfeyluC5cU5aOk4KRO9FsmIDEUBs+3BWOdyqLGdmQC+NGJzxUpQAawWL
+xkLdYy2jXtElxBSrVtlYk3LdTQ2P9eQvIJFaBNOK79Sg4Zt3uBl9F6s4QOvPsSDneVrTs3eP+l8
1o4r+y7KdYSjUtrHbhy1VEFsmPljz5LTGV1qqWCFZjDSMMBnErobfsTegOqgbyJJ+FzqDMQc+aSl
1LCpvqBvboUDR4XjjuJs/n/MYET3eMhyj1jHVLiMHyOL5c8kWT3rHyJlyZSWGNO8RiivcHVSdgso
2Lw6VKWHZWapT7BlFBRluPLdTFJeXqBHhoHQRp1lSgj/Alm4CSFLRn3ovn8wCG496dgFrxvi5mYA
vfk7D2OjLO+4i07nLWGM1mLywA5Kn0PLznaJcEUzRvdJIT/LdeDgoxaJEEUeVlj5QKEdtLNJj9dA
e0DkYjwutPs3wqD7875z2bUyeuuQBYhkkYZSOmPbKRZHXxlaKZHf+tGlAcMBb9xFstrXENhgtnPQ
0SOw3B9xlImJemWsXIUls7SzZUlthSFegUUOxy1tt34YOxSQLUy6iL8aa/MTK6LYbeQHc4MH4KHo
/86YvdjbjRlZrhKyJ8E8Av4hUY8S/TPG7bjU1JJmv9vFa+Dr5RD3KwQdMO2RKHytla1W8NERvZDO
YcVjEkD9j9il3yJwmweGLQXboopdSiqpmVpdp7+JwfqvpDo6ziVnBshuZ6XigyXTMmsIdyhmJMGj
mHDOriTY5RpSS+9lMS8+4RZcbMj4brtdbfpyDGt2AxzkHWiIr8p/YqcxzIyeGI5NJcQCOcWmZNBh
f3u+isjKSaOtcK0XbSTBS9KZgfgD2htcuD0iaUYr2XlG3ol2w/QON+qj9y3NVZmj8gmKyoz106mG
LiwoAp1jlfozcAXr40LzPsS5ojrUA4OtnoJbyFn4OaYWuAueby1lvUYVoy8dwLprrEdqB1wa3jZF
/UoNUWyNZyvaTi7XVoRahq6w2gH1VthIrc2lvdbbrCCk55JeQdzdxv1vGj1YscyR7dwnxyPYgwnF
sIrdAKUrCwkBnIn3aXvRTdg6JSEqSDUQ1Y6/fy8ioyabShXtrByZOj8N4G4nFzLFDQ5bR5t1rPmR
3W1DT+AD5QJyYJXgmV/0u/E5t7ac61Gnn6N5NdRapJ83N0KonTZfIr+RLfdWnzy27c4SVKrviYtc
4OGz8HRVgfsBCY2AYfbAT1Xp/UXdCM1621usauxK4219J9UXQCuGOAqZW7RATAii5KK6iOTYDiKU
c2iwNI5ko+p8pf1WD0c1q5sKrI5BQv15EJ53ZZEjxBdShz1HTjTa1PO9Nk7suxb/HqjH+6Ux6KdV
mIFp7kHKuBPvBoSVLSTx/uxuskzWhD0SfguF+UCqtlnuBxLOZxL4RbBhYLZTvcQAQSML8e1J+Yz2
iKvYAEIKBtUcjqVXnGPIIKd9uHWtSr8VNfbyef/bPQp+Q3vnp3J8GTLM9oiM9EmMCFHtOal7Jpw3
2Icic6Fhq5QdI/+bFryT0wkKvY8va9vX0p+1y1HSQb/I9c5KjQyeFPgF2iAH7b9zfAlBaOtIfZp3
UZuUJQXyZ7Qkle5fOLU7dne0nQXsZ6Z9+9gQPglXVZOzy3bniqi1A6HwG5xu0XyBvTKd5ovI2we5
ODENEWwcw5KEZ8p7teG4aQ5tbMx+3pjcIpuUhfjPeBmZflhsjB3UzMs/Hy5MO4SCu9KYfF32ipmd
33ULsC++9Cx2dR+fbfQQ65+ToqkYLlyKGxyaK9lAWCIbT2lXeNKSGTEx2rEhLO6224Flaqd86muk
UXGeSlPxCincBD6saSqiy2bsbeIm+Rkwqx+eOlIUpJ2rcyI7ImvtYmJQfYSawsX+bzJwyycE6Dmv
sa906pAFDJu1uFnlSafBbDxdl4g2STWQJ+262vPk+xQ2XQt2wBl4JjzZHvLmWa1Ans5QkPICBwpd
7VQAbxGGd/75azVVWFKF/JTkUHKEmHfI66tT4tHsTbYYfRqFOqKkFy8xK9aj1vyTvsTIodKPA7OG
0Zk9F+sShqf05XR5nshBMrIz65IQsJxOGcRjC0p5IxBFCCFFaYN+G3TauTw4Q5sy1hS+iA8Kk+3U
ehKFTKDymiRot5GQIIOV27nPoAAfRtKtXgz+RO5q4XsNPkNq3HcI5rXq19gWFO0t7IZltGauT74a
XnWUuEftOPAazjb9j95lUjm9ZLpXxdFGPz3V9vFcHh31L+VPQjEFqOAnUFvDzROqB12QU4NeKkzq
Wc7/2oFsKG5HW6txA4BOCELDkoS3cUzOUIIyuGt64EOxjfRo3lSs7KvW6Ew3+ftLV+SxYUyi+My+
csqQX4MvrcWlvTT8wrQL20/RpM6oq3eCVNfupDTEHyTjSpIoCWd/KbtV1QaUXzNRDLTOLpM51sQu
KQQUmFTmyRAf3vCrkpyLD9OnTFr2Rsb30lcnD+rXUasomj7OMTmzrn7xit+Dryi9HScmBStBDlvn
m+O3t0b0rtneFHdonTJS6LtBGUUMut7QI9z9Lww+4rV3FAp+Ybn7LjmNhW6GPxnzfBGzbyVGb3bx
am+avdYfiR98tc5E6H+HEXyGGEAyaiwb+YOj2bQ7S/M3pmiLqwBSmqp8w4JCXn2kZEAYD0gCVzDl
92WTUpilY8xOzHNaU9bLThfTwaeeWsdXB17MJTjlcPhut2kqARLNWD2lc277NPuse2xwwtzDi1zc
hLG9F+GllLr/IK9OQFIFWreFy1k9InILJCFkvYvCrlSf6xEsxswQT9mxpD3hqu07hLVpodyMBkV2
VQkveXbEvKLoY93LfJUnnD5NCUhBTFZUnZvT+jxEyYWWVtemulVCHD50Q6FRTgkWUgi0cJaUyegi
cyCjq1TPMbHTSCU2M+6WitLVDsPTi3uBl6JrKAQMSkDWI7WrMwKm5BD6jrCGdQSt0MLrFYDR+8vl
ss9WoO3QKh+0xNg7Ba7a9qFTxhjwoPCQLWBWrKfvqe8VbOxtAavx7TK/x12X4EbfakJVv0LoVHVt
KYU7B08RSlHAciXtAaSKYhnmopyG7Wj9nzprU8YnMeBhxGOzvF2RGXG7QL0MkrRPd0/1aSWkyr62
8XTWMTi1rRif1WMnBoL74gg+TfacgxQ++jiYX+vyCk05D1m8jnEHFR0JrYUM2zJo3tBP3Egp/2Ye
Jkxx3i5suVVXCQT04aOadoxKTrEj9mWK9gDX6YknCEwxLJ0jYCqs1Rp6MAqufXr2JwI8DMoH2qBA
dxwg9w9XNzaS2NGXzxKLYe9m3YZigc3IgUisG7ZKxHw6hlLEQUHbhguQF3DVxJBCVET6uko9osnY
j36ed4zqDKy7Yxry8f7nDn8xFmCwME6DT536Uc+oiA3PjjgEHIB01aae30da0gigkpGRe/o1bIfl
ZUTbFA69ekJMSTvDeuutZ5pZPspE7EXHwh1yLu9jVR5zH2D1zkM970MWTyP2BuGFILAzh/Jg0Tsu
zond1a80O6DCSGLPaXVpvLaV28xcR0Qr01UnpF7JBpsmhCdaVvTGmiT25eTm25YVeWc73guDCaY7
hD6myJax8C/d8HfuGgQypBXn+G3iQYQNp7LnsW20QIlIH1NvRoiOTUu930P6lsmKtwNbWF5GS2OB
sFCZBXwlcdAUq7sF/DwaFx3VODKGIysJfW+ypdEpkqmMMJeSB7fq8hNjATgeNozjqC09hFkGQTho
umtECUMS0d23wF+rGqXPygE9fspfXUgQ5dS4z+ZZKskQUvd5Oeu3sAaVvCd5n6VJK5A7lyRmHZhc
30T//l0rsQqhUO5IZG9PWOtdhfBH9EKH+DYxiNCiWqRSB7Hb0KITNvcw4bQe2UU8CSb0Qs7z9yHy
8obpcD1ZzJ2Qt1tx6zsfJGyodqNwA78Musl8fnTUYioP5sTTU3S395gtXK5J0WjLljD0nvIqKs+X
ASs9K00gkpynL2X06HuDrUw2QGC8P6n0mq2ji1bz5ECKyEK2RlF40sRcigM146lCC+BqlGEZRze+
1nZlHUDF+LGwGrbat486ghBMTg9PTbC+MSYPOUA9DzXkFn+Sbo9oMMrYkpgGE9I6f4vFnZBZsU6T
OaQ6BstHx5op/+JzP/PrDKRVFRYMKFH/kSIbEMZvaSwam3Q40fsItn/k4buD32nZSjLHRtWsdb66
tCuO1EQragujI+3BUGLTlN9iZWBFTTmQIPH49CTjcZ57596AjIyBiYTlZfEw/f/mRJbRBRJ/2ALt
BDmbJ9S9qePS3wPBPqn+aslF5FvPPlX+jgk0fiBZFqurZJGKV1nTUi4uErJ5ilGxY292Fbz+OUvj
VO3wLIaRmSXSG7iSqMcMskc0A/kFLzWwvKvinIZC2k9d2Vwj08M+Cv13i/q4BpAgSmZvw1lOyEBk
T9OPBjV7iE+g6NequsVq9I233ba2XYJbPR0gIedJFrDhV46bpunbyaycsBzMHwJg/wu+3G7NAVwH
v1VS49C05FP9r6FSBo6guAj2U/iLQJX6VpJafMSqBQ4/sLFB1rBMo6dnjQVQCcIqGlJqzeaxlQa1
UN3p6J+YeXKRh7aKXUUF74luYkwxE96c5ZbFSOrBuyOqpXI7X7Zd0SjzM7FZsi5dbBQkFr8l2w5i
NndINx4Bx+4hDzNYXyaHMzRkoBLgduRn/f2tpKMxJbuRtPJLilfeK+NXzHCy141VM30oLJMM7sLW
4Q+bHrGGbijyId4Q7iz7i6XckjIfv1xaomS4rhblHJc4bNN3ceRSuNy2ZM5poJuua7mqeg9nHUI0
5Q7o1WYr6N01u9oeylxySS6dJsDcNBu7no6xKrO2UoVobiSekiC0/Kzs7tZQfPRYrqa/9/G4JeWW
D2uVgjCuLpEVqdUh95neVDhA/mUyA/krpLAKlNEd9PeO7nuC6a1bnbcHjOevXO01P80BMQVj9zz8
vXIGQ4BT9JJFL1XN9nYML47I9Sz89jMSnu3nXGf4DcWTBWyvEMSbfWV1vpeNiIlt6VG0qY84/tBA
bpCcbI9FniQPAAywirByXSe0EMydwZB1UiNLLyac5bh6ERRAfnACUxxNWGFmPje4hPZsRO1U92Rq
Ac9+PKeRJLERUyhpT3fgYbzcatQ6g0qW+DFPxbCPN4xs9BBvJtlM87FohkRkK8rDC74VWUMw/pkF
bB+907tLgIjep0mr6o6TEVtIespmkKoEhTUu+ydQToOaiCNRC4z0Anfl7vGfnduiMZj/gCcYVvcW
80yJbVbuEJANW3pZzmvLHg69O0wR9VrWBfFDzjiIbf8uTQ9MEaY6j4NHCGqslC9iXGiDM/W5g6Ss
bImhSrLRbi+xCnAiKPnxCTXNzecLy58Smab5skk5WBg+Rxn1fNfuZICfzVKqJV2SYQTdps5rTMP8
CGh8CmAwUwfyw2+E8lwg3DfTi8CRnxgICBa+fP/POIdRrAc4SXg9i41PGLnXHPqMHMgfAol4ezp7
dXCqou2qK4vUmJbgcx6ijnJoy9ek/WP7ErgEv7AzGR/T3ecw6Rj5GQ+yX8KteGKqKwBVuoYWXOLG
AcHW7rmENnGL9Krjw5L91z9PHBYIXnNtlyURF0zkknnrCDLEK3iuBP21BEd73kecmP5CED2Wc/7j
v4mDtuX898VZZlyWBqQKmuIOAQGPA1Af/wIYmzCjrICkHAoB/cj00FDub+wKFXwvocoiWd3a9DW5
B+ZKQnCqGsgvV0seVt8k0PfeW/XjP9Xmga//R35cavoF9Vf7VOx7muQlOB6vg5am+9bJAfTqqwCC
irWGtWWoWw2K9u9qr2SzSpiObrqGums25q/dvj25VrK68bKULqtQYkul7rFhWvCVJtb4QL9AmwuY
MB6PEy121N/WTn3PE3jNKvrSkMtuOJtDsPeuQ6rc5twuB8fmx5Fne8K6jJ0mOx1BZuL38gRxYwD+
3fSF0ep223LzKwV6ZBiAKCbP0f7SZchOIvAuaBmryQUJp2dqLESkfGyglwii641CPiG/FFovCxsJ
tdEmKpV0Om5yoiFxA7ttX7zdQk8CPHyCwBY1laOtRqxtb7HYYHdKfbkMl7eeW5UjB3PVfq1+8qg0
fcXBBX4T2JH3WXNZuK0BjMWSOuEhA1a2aRz/rU/67pVfxQWW2WOo6/COMsmMAShgk8O4SKmbIkqw
O/K1X8IzqnbOeMLVlPADwk2lYZjNAfjjvSOn4ORtgAKh2hYBocqRzcsuTo+l2hNwS5f2OWbG+D1/
XxhCPnbCHPFGTFtKrPGssy3a24uPNSJD+6i8Qjwygu7jLThGj0NdLjaslE25KbBdZDczJ+9YQkRG
2NcDz0OwU0iOEroNx5htbb5/UXxd35j23ii3Bp/caP0X0saivWVIxQkyML+5PeAV6/JCk7fcSf4v
566O66sbavke6NEYL69Y9YkYNifwbYcKvoT3g9zxMwGLz8Yjsmj2knRy9kvj+uhLuGN8wcboBgNZ
EnfEye1QVvzkgHj2bKsdTHVxp+vNm0I3huPeREK8Hl44ZbYPWfWjTvwCbfuhEG3fabzTMFLokvR5
N9HqZvx3V8jyR7/WhMZ8n7MrcCTUTWz31U2r0yynBYJ8n5KOrm9m3MwxAktMM4BJS6MGoi9N38dM
8Wmjyc+o3oiMl1CWXLL9aTLH40I8GUjVkTjE1TaadZpxBBkksE6VHVIfwRW07g56cYhT+Zq6SXoZ
TtBkFL4epk5bbQ6wlcSP4/wD6V087uHYdf96XjZCcm8LOJX04UmObQ4xSP03JHPaa7cKpKK5GAp5
p6PciB+/K415IW+sKNmSQDFWeURO0IZg5IK//UIjteyqu8oDJL1U2rKQChUJ6G83Jz+p/LePE+y7
itwtjXyN7p8cMCi1itfsmRpro5n6j0Rtor9VGy+U/C+JcZhWP609owcMfiVZZaXCyzi/G35gGRte
erjmmFM05e7bkfZ/J1jj3/PZSKK8zxvtgkf3p4KbCwC4fKG27lmHSaOQk+1DLDX0786EUCNmLi59
ckIabAbuGr7xLy9OCNWiDFvXrSTooxT/nyjEUnaNCeoWWN+dfD1ORrKnAgSYaPe/ud/wbQLoIZi0
cEktMDWhIDdynToxvPFUap5O8ON27qGhNgmfWlhR2iujKIGCLVujNjKC3WZpqLviKSVMwe6ag65e
2q4BJGokTWbeg0mSPNG7OdUoTGl8JGJHwiyrNbS4+RcacRA6riXt1tRa9K81zk3DsOvSWGkQYY4M
bqEmHmrO0cxtWZSydC7/8dU90N+Gw6wJG4/efFPRvfuWFvR3inUbYtijX3/e1HwCDLqPdbCBgq3q
x7oYHOZOFmCOi4RqV1DNzd35MRdQTk3GuVBbUfnee33N53He2oxtZXFw/BQ3tGczAw65DlzxsWQ3
1OSDYR3+9P58f+nFWe4xbwgtaXZh447wKNK5Eqr2+RFoOCqzTle2IyguPYCe5MNQ/I3vFON0BIFC
dizvdU784Afo9rqyy7EKMc3K6VdxbM+CLrpAsaYUtigQlWutew5GU4wH93luknVDHBPKOqtPBd4l
q2KeilELwtrHNOcUhS7YwUp+E55luQvuzCLQgDuox9bWR65FAXWUPqi26fjLTcxEIU7dG7cl9sRs
+jiuvz1B9BSHkEbdL3dvmP4k9MyrdMbmeFWpMudGSi7554a8BCYAUPjJNC0yfP/QgD9K9Pptu1S4
RD3M8YhX5bfio1M27cnBVXUaM1ukNtUqhnDWRnLS8EmBe4i1OWZ8QS9lXMDDeDIqzy22FKw8t1I8
vi1bcySn+WS0x8eICMXe8lDT08+ZM67+I0IlBLrYOiMZjpqwLszIQTjxksh8aRUKlkPEUmtReBSM
h7I79PNqz/JKBCB1+Uv2ZuV6RG1ILiyptEL2CBtLnuSediIo3CJ4fOvtr/20PKgwey+fyPz5APxr
OHsb2E//kthu+HYD/vc1kLentZPMzT63O4ZOmN8dd533+UMzcE8UHziqAy+vYOUosh/GTWLFY3NF
hyaHIJzGBOT3JMeUJR1Bi+FnR96hY61dh1jcw//VKVa8jfPtXWOTKs8RtNammqYSrpgXb9EtcavE
FTwLFdDj2g1UBRawF0/1C8V18m3JJZ0RsCO1Go84mvS1jDWh09Ej9JtnDLVii7ETFQe5FEFLYT+m
JdBvJGF3nWdE+tRgHrlD3V4y5YB5mQcPNET1aRnzd3HNBgrCV1O2YqWLb13dlYeH1Jr7GJkf4m+8
VvjSJU7Zry2eyE0Zd2CMDo9PsTZiR0a5RdZ84VEm883Fryl+V55fZHx3ZEtdhM8c3BBovUSEo26f
R4jGxojrjjOdzOIyHBBKGOM2yvqzsknehhKnI+CbPFgoCHDPsRYn3uOBitQY4LIBvnG1Jo4qq9Tn
mYkZ3moHatG0tObzr+iF7pBLcus82IfwpzsFZXyesuhX5SAV7WT6D56Ohcoi/a0i3jAUZtTV617F
yb1FL0lQ9QNCszKNB8M4ZgCe3+l18+zgKUtUzR/+/ByTGOmxFB60oSD0ko2K5RZlRmKydadOxxFb
wgYl1HoppmOlZFSs6yMj/NxTIYndnutwW0wP9/K56b6lNW1SFsJ0pYTJ6mDG2jkFx+gGKxQYFw8O
XweTu0KEzPjmCEd/HAgjYx32mCOE5oTj49DMCNHT4NVKog30Od6yxpIKteLVLG5JdAjASR7GOOPa
tpgmGzlZv2eGLkKZ3XvGDcYU0obJsFw7ps8jGE4wxT8MoBmVKVOwB25w0d5xumwv9arCyhe1yTGm
tEMbK5zz4XE2sEKIzmxO9V5jhOI5sgnToEM75V7G415bUOpIL144uzOe9sP8SRzQmBTmlbMD+xpX
vFmrHbSPB6zQQPokJ12syqknZRUpwfTBqcTrreA1F5rp7jmOSa54P3ogKl1C+tX6BQa/6q+wx3S2
umwV2rmCM2RWeyvnsYj0mza9uRxWLU+KiKuIiFcdlMsdyY/s1IemBj98/t9/ieQdGn5dB/94l3L0
sC7ej3I7sa/mKjiwZUq3PB4BNN2aBQS4ocgOSGq+AHS6HhXHIzstAw3wRrHb0HqtMx9Tjzb+4ejw
/b2OTD2BIS/9MxtcDsfX7akpLGo0pygk/QAvxQ9O8q5W8h4ktuFj3tO8vP+0tZ9mdn/gikRVLrBE
5fR/xWnEYdVL7k9CfbxvV9Rhj3fOZ2d/14qk72kJTX0ka134C6Fm4LeTKDhkavstCeHpkg2sqFUI
dqfHAr2ildExTEN36cIK+RaBRe0GKzBveZfH0sv7sLnpdpAwUn459Mfh37B1gh1nTXcPeUTkDiiG
Y7HCfHxSunwmy+Fw6ZfRxTYs7UGDNtYRb+maphdKVg+709RVBdLwfdYh/53a7lsblzLVEawN/JWP
76EYkh5GT+mys52Aho7UxMwfj2UhfPEmS66Uvly0lJcHUSDCZiqkd9Ge7HEu3tVxGDE/UbqzT1Tp
CpvqJS5zD/U6kDu7yjg4THp0XK85BhRcCgsuHjteEAux2wRWVTCGXGXIrPPF0UFJz5LEMuwFOcOE
uktr2ul8tMDql+Gau9HLqoCiVkkyolcN6HSrPUv2vquLafluAs0epiXUAyWWeHj2Fnk/POkNnakM
nFXJ/aBNzTBb4QBLBgXMv4s8pikQuyk57PhhT9gy+2EAG77JPL2Ffw1WAPKDaxe89ELCWkoxCnuk
h0+AJcpswYJgTu3T63gXlkJHVJcb9/SwvwKNgfs4hg7Sf/a4tlVp9Wr+6WV9POS5BC57z0RA9Jgv
Yi+aeHnx6DXm5piJtPiXh3VbSUOKpPSiaR54OhwPEEguC2AP5bT8GYWr+WY0eqTbyU+ohEN82/UB
bne4kZ79GwjIcnRvyF8EVrBh5CeJOIF+Yfs2McT8vTfzrPWAeToi0CvA7Pb8A9PF4YHinXMxhsCU
+h/KkWwlebFXKGHl7lVtJGYyvVPryvrKhE5RRl9BuIxFZFkDSGSL0szGIarR8eze0q3IpiBxme0r
b5PX7+Uiiv3r6ZF06yUkR5l+KFPrV60rInLuG65VotAeNh6UmEPVIB0zLQPQCRFidyqKrEjlZa0X
plRURLAl9cVyxlISz0tKIXoRetxzjIujoqwiArtO8sphjnXNTavHIVebEGVh7bGW6r4pHomUCXGk
qd21xDtRwTT0BKCC3Dm3RLJ+gsTGiTGA9+C9jDsf9epEYlUFl44Bmm5JtjEZiUhEAB27P+wk0KkA
v+yEyqAOK+XmQg4O4VdFQE1KILv0Hcd6MGjFQhwPEeoNkUwjIn6mLjVRFweuedjlrK1wCqK7iZrZ
3Yv/1qUiAoQhYqgFdSwaFqSdl4Ms9rW4QvIl36XmtF1EYqSHyIZF9JJr7pGG5t38CrwcUpSRoWWN
eN+o/IkRBvWTIbMhHXNkgrknwlH4AZLLS6fB0dNrRiuCuHuhD2cXSS1uZabnuewvxdw9AkFLHcZX
31ApmE2JGAokg3KUVx29Mmlj0B00NoHfpgwD38UU29d1fAzwO400OA4FAF/IuhkNQCweNZUc3uVD
b8cgkRbdx2QZyRSN71PvxcMMvFkjIrlBRtihevWNmoORu/qMqfKg5xSCmyA3dX+FcijN/Tb3PIpZ
Wu6KgIQqe+OeReRsRQ3wATqGIQaAxxkJypkfdb5d4Vt9wG8eZxBcSxdIN4fgua3Fr6c06NCd35dc
qCF/CbQ3U87xlSZ9oRkw4aj/1fwysr45x8xXdfbPIeuhwXMHCBLgDOnYioGJqLTvnVkkZISsmDTo
IMmVZPBbA4JjfRZclmpJ20FlAKFUJkHsw92I6/SMrbHkQc1ILQwow3SLxQwLOlMSTRpT9PrfR5oQ
KwCwkEtPKkjAjV7PFzFq2Xphi5hoitlers//SjprNXG2oXhRRqK/WNJDsCHE6+9/g3qlcKjpY2Q/
2r3Hji8t763Yt0zUjOd3P5mn4YMn5j89lSgy6yoBZP9K4gnExDnchuoneEqplCbObPzmKlKupBL+
WPChAJR/uv3R8D5PGhsd8SWGspp75Rims9OUKao+LQeW4obkCUGda35X1m+lTAuZjBcJJ/UBq+dG
cN6sy0rpHuUZ1vPZ5yHkLntG4Dg51I+dsjePbeqtwiizD2IyWqiGWH2v1x24GqfGiqQV+mWv2AzL
NLww8ns+jhhI2X661MzMc8ecbyG5YiK4VDhSC1n82mJEyxfUZnJuYDsDqV2sGGPj8PoKUVRhmaDz
4cuxqQin2MU2FkSJfK54Xu8zVMJ4MMQNQ1Lg5+AljLsLgo8WcZ//zgTn2SSHadlYTqHo8mKezzJQ
fFb1bPBtbHB1Tn+LOF7zstu/KubEMWrmAKwpFY5K3z6/MySUCGTDMfgv1pvlETd7EK0tPedp3G0k
lTO/Cs2OrZMnJxBDxtJPZVRundWzW9FavKY9yrJbx6OixFbPQ4izIvBk0Tbky04B5NTltgO2belN
s8v+fsM1/AwkZcrYtCNcvBAUzafMXZzLFUpwVVBb+wSpfGDiULxi3t9aR/6TyRI9Bd+1KNc0Qqe5
8H7LaCCkfhtjyj/Oc/KJfJKgJLmF2n1PIvLUqBV5Dfr6QAgaCSZrs9B5Jm9HUtYQUFj73Dr5PRji
sgKfY9nLMXuPULxoDmOqD3ZNLuB/iYau7PXe4W9L5H3PtZPQsHW1LVgsKdVy5RXgj9SQoDca++Et
x0v1fgMrPu/Q96hn4MjCvVWNs955Doc9rw9j+g/gL7OU6LYl1wELxKi+ib8j+ORHh7K+kWWWfKoO
d/vSG+iJiDpVFG78jZaE+6GndUoXwOAKhTZ6uGFqIxV8idCVXe1sA6hERHTAW5rwukm0IjdVVC4V
5sHbNu/urOS9A2AwNWT8XHQo5MCzjIDB2RuYoexn7n/lmvxqiG9Z200xb8LY1Ttdb4Tmekc9IHUj
EP+T3Oa/PsiAqYjNQISmPXHbURlxqZGmOEGTVwipk4KC4fo5yvXqxIWCV+7BdNK58fUMVMt+z6zX
RskaooGuH4jjMsD4axBrS6be6tio+Y6Ct7uPjKaF4ir6tHmnpUGApWG6prvp653SgQEg5RMPOy60
u363zSaREB3gkFUwBKfBeThSYp0gZyTDAV9GjS5LYf/OhllM/FjeLZDXZrr22gybSDqspaw6Fy7G
jF5leA42foSOcIRcG9OroEUP3gYF7eI5vkoMS+cu004wF6E9hfxHzZi4b5km4iHSVnNCcUsmaQnH
3Um20cu5PuSKMb/8vrB4YTqIVS/iVNfr7giFs4TQyZtoMrSgvidSOmlx6rJMxwi2v7nN3mB1olwO
hkx+h6i4OpNtZx64JvfTzFp3whLTtsyWn4Lf+YXed42NkFEDueS8w9149vK/b2mKg5eRdXYANdcA
jpKbSXJqQfuXyNms9xjlDT4uh6D1GP9AB6S/afmmAfXsAj2nZiMz0FMXqhRI0W8W/tkpesw5a5VG
Po3ConRU5ymPhElp7DEnxhu/GK7HZ1LZtNPoqnaRNylCu7Tw2R79lHnFXk5JMJcLl9NCBjYLDvpl
OEgs16RZ9nwJC2Dq+1aRJupVrihfGYHF98KgkLrHgTqRCJxqSwRcEftWAjzWXOHwU0gbr+uhMB6/
9qqshz23UKr5qAEnTrIh26Mi98Di6v9VtqM07JlgjWt1JdhpTbxi5LuSZ1SMcf+1D+9V09RHC92z
Q04AbPlYMlI34XPPS1z1ZirjptguiW5rEjVueOJ/mETKOqWACt9h1qo+PXh6nWX9NjjxFdwtq29R
UDkU5lLeoMtfPuj9e76QAALGZq3XPpd7kfdGNrDyt8z4Mv7jsPk4f54+s4IKsnYVfZVCC5Bfd2Mr
QzxbTsds/w2XxUTaZUEpsy5wSoOEzuYxixemC3tOAAdzos026yLGeeRPEtzzfORoMK443X51nuc0
/CMCho62yfUaGJn2PRRvIjWM1GZvIh+GbHurtYDWZ8dtFIe/wFRBqgadqwAQxPKVqiNTMBG+JDQB
zjUwoxwBu2TALtrfgqgvygyvhGglHLUyAaF/fgVg+EvsvnzGZHYsCYeuwRQX1JIdwJoSBxyXasXH
FdkFAM84dluw0ARxgn5/0WEHgcfS+XnQQT9CMmyQ3T6TPjdiPtoOilH9SmtF4QhdzKROgUqtLw2H
J0NFzR6Akzs5hZg3h/FGwmb8umQ7y74Q1TBOgPdssZflhVopFSbYQeIQ3Mn9aCoD7GuTiqIEzkY/
jLmBRZhfVVy5rcTqkQs0E7VE1WDl7vtP0X2WFDQNcPXdzhggm4fLRvzSUVnJ/37MnwuH+iCNQ2ux
jiZYh/mL6Y98ZaYEvO/9MetvFzH3pz4LePaQCih+fx3h4e2VrpAkuQY4klzZfZxd5z0C9tFm+OxM
bV+8+j60Bxe3+2CEk3ftSIOij1Tam8YQkQoj3btxWQUuAVfxBqlouUSKKuhofci6FmdHElbXIOQq
08fcke7Am8PP5k9wAkUHuLTSJyMCOjd2pcgzV6n92eXZX3j9jM9vb443PJDPL5q4dPfCTfjtw7MC
y3SB9zJofIIwLhD9to8cZM4Ibk5XuYRi3RpKD8nqLqJvcgp3MoMMSrWJzz+1v8U9NIx6XhPL0lzp
vPLusUayPJTemdALmSUy01ipDxfGQx8pAYx2bKcRfltOxLKQArf9eoakf3hBxbsf2V1DCqub+Ak1
yFJcfI+WYwkwQGWCV9qV6Zn0El9jzqCFyyZhWgVhMo5d3dz1EIWwUkRijwSugv8GAGBnix4/3Dk2
nxFx4KJLbsST9X+l5yQGx87EwO9AMInjNxIo8Ay52DwRub5HjJkXnGC2NWulbq5VM8b8PM9eVqpT
CkX5NyoLocQyA7rPJv8EQE2kksBaV0loZmheBa+Hf5axIydj+4YUdHkReAXodXy3D8fwJNgBCaZo
DEHxNktuEGmGWvWnSD1XCVciG/CPwuXR3TaiC9j7tjm2iaPxxfRky8lgzzXBrcCISiNSiVsw+FyR
AhrXDrId4QKszYuVKQz5k+1hOxGo/lDHNnlW5vI63KAovGXzqdsgg8G9nt2+5nm8Q2WsgX2q5P3F
Hh9I741DqP0jaqpONrxVTYsKHDsIoIz9CSKKPrGtqwUaatdiWpBj6/fqPGsqbe6uhrBHDWRXihm1
KAdo2XykyKP+mfN3Er+vLvjGjZ5fAf8LEl+9eQtYgTHSty/+pa/n7MPsCITmdqrJCdrFPlg11JjM
vrU4duI2y7mC1bTRExVaFNNNxN4oGtLCAFhmPG/DQl51gTTLOFeFVtU6yIglIBAFrdzKuBQnPeWV
qTnv6PRDN8PhYz3/3+33gqE4ng9fHjbyZmGobcu6y59Vyd/MW0IiDDy68hcNOA0O/gmNLSZ50xzv
ScKNaXpCD9QyzPo9covUQMSwZ7YX7v4nctMfsm9JooU0Tmqm59CYc2blXstOi+LrurD2mu9fSqH8
RheUhRxIEFJCWWWBcsDHScRGXkG7PMFSazb36YCfijSt+WHCyUuBGTc4dIgc71Vwg5m7t5pSNBdU
M6e2lhxbV33evWj5+uSO4+3ONETuF+I26wvmOntoiVES1/Ss0/3DPkD/QIAPp2Z+kjz+jlXRB/fD
vU1MdH1qSDxmLZ0OLIupsEZAUJziEOozcb7h0DiatgKbaFOQS2Ca74cC32Sq6Cq1MFTJ/o/+GLux
3w5Sot7P1ZV8LBEpyvxRnbpvIFoPrX3bAuIadIbjZ+0e/Mv9ppZjEyPhH3EtkpqU63fTvORTgA/N
ZKBnqkS5EYfqPkd2xxuUavy3IEgl5pIU9mLGYmQq0Bln5+uUuZOAVY3gaZql2N3eIkS3GobJlki0
R1KydKzdbv62zLc+BkahIqbQhufntaSk0y58n9Y4csee9pW1HVzQuDqIZkq7RGFKfbFzEpYk2v7x
WB9/XBTucPnS8glug4dZjD3wdgN242wJYVbS0XfC5Vw0/sZwQgxRetnEjcODJjq7nDlMeWK3p9jM
3chkayn6o7Qzf+BhiNowIBt+Mn49NxM38Dwk0UXYtbAVvF8SJDg1kwCTtjyMQ+aZxb9C5eT8gpvM
gWsc/yRLHLuYegMFQ250oMCVjUcrApkzwp9KhtXtvOY/b3G0XBOagX3ppLKL0uNd/5zz0cnAVTu9
nm43vMDOBONmPI3U4H3YovclWysYPK0T6xAEmpbyWf2TweOR14en7npJYkjJ9gIipuj/LRe7aL/2
gGy7dje77VS0ZRDERDjgbLsfdymXWJristcqnTDdqIrJ891QAs3FrG0cRdRfgnT3EcD2HqQEFYRT
Cf21VVuYgbiyXlcfCAsvQQDj3kifEPqlenDmTzc91JesOqz+/waDJW9s45Jd+XAa5r74YuorZw+t
kZulDxPD0Md9lnQGYD/NBZX7oCrtFsHQ5NTdAcIwtxNxMKbcak165A6cYJOFdVbh6hupz4OQ/oJy
MGbMRDhWD5Sobuq2YzOgoXymi0ZsaEgFLBR1VEVsdMAbyDhhpIR+V7bi3NNWMd23gwp/ZWyjRGVi
a3ti3zEPeaaODGLrf/kCe4XefC5kaPKUHckoDqZto7yJQopq4IpJtvzOhXuMlTACpq7SnC6r8bG5
3DRFO1JulU9si78omxZubFl1zUklyhMipgu3HLmVbeYg5E4YPHQKr+N0K2zfp9r32x7y+PhqaFwd
KDfEOQfKg8Z+muLjdHWUfUhMvHFg8C8O5O5QgerLKUziM126mkiPtlJjZdeU+PO6EeVppQLvjRx9
dM6kNA1D/5zux8E8vf7W8YZy3RqK8JNndsHWROzL3gkUP2hShBPgUTMKd5cb3AbFMI3FBWPX45Vb
NILlQjLxnizWzY/wygN1tNnqtRlTL0tlMda0w3jQx3XOprGsB7B6g109cmLThSfdQ2VcYnUn+5pZ
wJEPZedxXvv228vVakQG6SnsszphJUbkgdTSMdOnlI2h020zNUn/zRYCb6WPC7CGrpocSBu8gT7A
8iQ7x5Q2m7XyXkleQZUrSkPfPxUZ6ii02JOpUwF+P+f8L5hNqQH1rlcXMJ9awotsapK70WJVsFwO
Kh3RmAOiDMoG+HfF7GMW291Y/1pdIRRT6l9F9zS3owgu/hkLJDp6MWgqjhew6eHDCmHdLR7fcv6T
iknGFE68mUzBMt+uvsMqkz0peT9N9vZIyxxUOZkvHu82eIqsU5byI4EFYAxzlVqMVvrh0d6yV0w6
MblocBJf5KDii5JPe1J5PVlLNHGvnDIjHzLd4CcJjbPwsTlwrHGbYiSk3SOtUrdblZ8xLMg78loe
YG9Qzf3Nh/bBdM6GQeCN/MbctJkYmqblSeJEcKITu+h3s2Cdcr19I+s/lo6DyyJg+cYmtdIdC//b
aw8ZlQL7O+yYFI+1kiVcseA7sBW+W9+yFzCPwYRlYdZjMRWMVKFT5kRx4d57No9fP6cWr21xClBD
fWO/aKRFEXJ6Y+6c4l6yBaOGc97LPrSUDEjPdZVB9rLh1hiWCqjQDAk2VtNcJhSBUDt3jboFQtgH
R3VW6SfkGo3WWEKwJTkVo09kffhQbAenHQhA1QSaGfXkZdnxczICjO/rIktGnUhyzrBeLOS5RBJP
WJ4/FBfpEdAmAx6HOkqCKHz3gXV2DTR3YUCVlkRotqaWwt1vaL/D3+mEiA2L7gXcYeeKyrgaM8Tg
1VNvOC1kg1+vOwWKQGjZqqvkqyF1EUe591k+xTXu5SPhLCG+eDyL0D6gVcQ0sT/myTmjYpa4AyGa
FnPiMf5s4QjXT8ssuPGoxrr9tO8HUVfAqYNmhrBrY2wV5nz6vEZMXiuA2iCNyBEKrcjN7sJJq8pr
ltn0S+n2okiNNWSJrp+olIapWM+T/QNo3VH0mshpjCV/AkmjyFCiRog99nhgXzCs6C7Yy758K8VI
qr0WEBmV6pOyPSA7eDBTI8k4Hu8pOqDB0gcD/dDJ9nsDwCmb4TK3DgGqFM2pjBu56CvCWgn5dktx
fSsFMnPD59n7/tNaCkEVcflpb+P7d9lyLoJSiiaa2j3484AnmyJNhVErFRE4weTx+3Am/TeJuPk3
0AJcgU4Uvxu8xfJfR+JoltdumSvikifuEtsoK+FyaiV7Xx2KS8GNtzWWOU2XqtCBU4B5WUaehVMe
3NmdbW2Xr+EL5XJQD/0kASGDXXfKpbavqy764rmkrBNPLFFdih8IrOpY/ouSmstJLe/b9L4XujRo
HqxSn2c/VaUBLwlqqvajLeNYjmMlKXU/E/dUzXXVWxBg72P9Arl44/1+C1ROoyUFneC5XVLbiSYs
eyovZcvneUJluTakf2hdFG0WF+on4QinZulPvgTLC50T7VD4phmxDVyVO+w4/QO/SsMpgr67zcDS
7RmGJLN5rKKiFItoIzu8DCPr3C4FNLih43ItiKDEfIYL5aKjP0TL3AKSAZPlrFR1fXTthKd7KWKo
4AwHPPJVg7ft0odmKCBj/JF6INX9wsxKLYAu1wZfVqMZo+jI2MPHzChbWVIzOLPrI/FYG6zzcwa7
JbFcHPrQTYXt4KToaNOeuS9qHj5DygwADJZoH3CrEnbaammxCrjnwDwm/KoqNzJ48JZNF+hFwSNF
C4k7iVrHRRE8kdJKC5ErR/5bccnIgv1MQZn5mgC+NQFl1D+UJEirVS3fjVd/RbHiy7+zftitd22a
MFAIGeUaIsRWNTPNF9PsHmSEX6Qq9s+qt5CTixnun+hZoWQQkmWqCStwMH2c0DZZzt1huTQAMgfA
43u92BnI2VN8cnJDWmI1rGX/80a3woEdvSQ7qfAbXrzv0xdddI0Pkt0PqQzGhd507zh7pCNcMGCn
/vpFpi7j5gRDVidYUNjSqR1I0z1NdkS9wQAyCK7xyrRSW3XtkYGVmZFiGMEZbU12bCHXGmVXsp7g
yHNn38lwrgyu1GQaQLCCGVtT5EEYmz32L/qW78QZ4MF4A1772/DLSPbJNSBMUl7tbAbQd77K6I3w
5uwcWyHS/fQ1c/HGGNK4jKFqEkUb3BBwD7vGeOPZJdHXaS8hjjxjA89U5ywpKd2BQuWXPBT48eJl
U37YTJnTzME7fFGS3s7wLZ6sbBkUrY8iLRGYit3twc13ERaIHP5tkRu/gL8dyP1j87u6GZ/CqyWb
fBOVLhaSFGqkH2rdQIqQk6xfpIJznrWTmZatZngfvlAsQrkxnCJNklELNzw9pBOT37zoRCopYO0U
I5nHLiEI/jBFa9Vsa4K3dmQZ/fTTE2/ElCK78YhxclaJmj5VSQAeeTHXXg9w8oaSHT054pSCJU4y
EnZoCj4Uf1RxesBDVBdcFwKo3RuvAw3glidFfM08A0dJprkPapaiNhlb/N54eu3Z347H6cBjpDzl
gbKk4t+rbwnScmIKFVBLiUxL5z7Xfc2q7tttwUbmLk5oodDmNERAY3FXfwFUaetLlnCeU1I01rO/
erxCU6bZdYUvbgBtTkIHGE/wq1GsKjrZvDOONdq9NkRWcbud+s0IpHd+23sysPK6/2DzVWR8G6YQ
HfawC1Vgsd3q4F2zS8nmGhlIseptNyn5/IDvCTckmp1+F7J1a4IQV6xSlqCaOpydV5o7pG3ynjKh
EgTCdokmTDwbMqgTFepjqmIuII5DPVCUGajDVTFeRGaWzeHpxccGsz3bj9Oi4PU1VTnIRG/EfaEr
ulTXsVlcPX9gmpBHrVAweNuBrdzsxncGQvfDv2iwc1WpJIVrRE/sTLxG32HgngBWfaOTHMImtvaw
3gh2ENFg77OBFqZFQV/lZI0GPX2zJp2W+BXYT51BwATYB36SKXrX4x5z5SyQknLKnSXkFF4mbKnL
lwJ1WE94AcWlrkUQNAY5lDJS45XZswXU7aZZUP+gVnlQT8twURuPSyiRYdfFjC3W+1pakyWKOFrC
b3kOfCztfm/iX9m3Vje+4HmAUof6j88XMEZSvRnsGhcd406Hc8RxEbQRJe7a3y18NjqN2NBm4Fjk
CuP7GwEBMZXb+urXmqVg5gJaU1eYMBa50SeqyKiE9BKPaEEf2put9WLa0WAStyu71q95YP6/qR93
lcMI/F14Dj5M+6yOl310v7dF99ijOtsCt+3gwzi5cEfoZhGTecSEnx/DIWCiyqAKtC9ZxnitdNn2
HP0E9rdUAdq2vPl6+uFVH32l8o9VD0IFAj5L3kwr0FozKqiqO2UjMuM0DwjgRtl4clFD7FwVjUxZ
r5ZaLWCI435YjPMSBuRXmhDqfAzXpNDhLvjHQNZYyweWMiKEU7r9lCV5WWfjfEPez/cscg8FthPr
AUlzxECXgKDI9aaR6X00F4NtuAwFFFdM3G4d7IeyC6+y4ednMRqIC+80BOA8I+QOVHhTbaAjKaZ3
BDNSrANAxZ+ABjxvSjKBhkTuGlAM9/8AY7phwoq5+MG8HlbEJSpmLNQ5KyFObd24YPig8qYbp7sg
Wkiq2lTXqMDHg//nSSgO2qr6BbAMBs3pv2PUmqE8/fsmBNjmCZTv1SYegCLTmtYpmyfWD6xzP/J8
iPI7AXf1t2clkEi5s1Bk0Y0rzsMrIK6w3f76A7EUU9dJsmb9kMsXj4x3UBWzAxZ/bplHKLC/Z8Wv
wuJtrmGOG6L3lZkxde8HCoEVJBV6EbDZBgiMBSw9Bk41PHvdSK1AeVS9ogDD7s1dotpKVm9G90Ws
bQbRBKYoU3oj98y0Wl/h+XR4TxkZ+iUGeqrfJ2+SjGmExX2navTDULNPQWJHXhVBE+bkGxh9/B8s
pnWYQZ6kGdDEkH9/iahgrF9pK5Hv0V6yt1YoemTCtQ+5GxRNYOAXuOOk0vC+eQUr1vBSsEw3QOLG
ZJIvw/0XZlVXbkSivEmR9mQfuoyHJC+C/v/4iltV0i47Xlf7awyRDrHwd5SnWCf7afHZvE/r8DDY
vL/87yarKjT52Xas7yEC528kr/FsBvgtNaabwTnnVjxmXOBskrtFJzuQe8ABKEUpPqOu7N5ltNB5
F5xOVUJ6bqNzEGSXJb3f7L4wVIbKasXqGv789GEQuSkJG9yPCq6zYiPqTnhVnXw6nj8fftbYv6Qq
vmtNOKeNIX0nBgjsB2NOBapCLMkl+fY6hkFZPB+IjTV6WsxjldeWFk2A2qga026/0Mb08JEYZH50
AItLgST03WEwVu8gZMj36lm65vhP8ikn3MS9w/DJsrlhyPRt+oeqfonc2B0dBztzgxnisQD8Tlaz
lEiAo6gOD9CIKffiCjT8fxt/XkIjd+ld+F/jpRzRNHpwdkrCAnslu1xviRcvvWdFQMq40/4dl0q1
MZ8E3n2XhrqF7ranfraZMDVkj65nRQy7MMEZHQz28aylBbTxeYBgdyt95/Z4NT7csnhroAsPIVO1
QY80wowElFTTsAE8RVrQbTyKdFOb2hDdDVbsz4Cji8ilVvPYod2jfc5HQ23lQFNv5YqkWoAlLftG
wVUzy1ZkNMXVwR90TmddVqMgRjkqBzgm+ctCsotp0+Bd7cn8mOPt+EaMzrcT6mfurboiHrpKLvx7
qthwauhsZW2oE+j3yyVctw26iTcM0VmaEvTHm6qLZv4rPrjRcEEb2NtaMKGN/sOw2hySNnxRQ437
ksC7njrzzRsGmxC0UbLl0cc0p3dBWmsQ4zj1kJjkxYGnzXDGrTePWf6Pq+pyhOaujxGhOKISxWhb
Bcb1comSo5dynJ7S+k36vnFPBcMFU3ts/d+2OJ3/3tfWU9nOg5Mk5NJgN3glB7tSvP+65NXORiOI
amCstPjFvM4HTZO9zIjTtMGIGen/hgiP9PXVBk7GGx5/u5wt4wqBDuSiRAnGDYNSs06rBIM6cHRG
cCyt1yOliNWaeSrQTiuM71qWo+8W6FOePBsUzTIQgq7SYU8dKxu2UJafw4G7A4kiz7SCRpd6V6HW
0OjH+0YICSa7DTBSt8B7+moXmhPsdHaqmdDWSMAXoFm8X9FMD9neA6IRc7gWFvbW3vmdqBxjKDY6
Lzem10VNB2+Qm4jcXA8fpk5su8Bbc7zT4nOp4CeRlqpuCqoTE0WWOjTVOQ9kG9YWg+8z2B47xvWq
AYpeZK9pvBmtwCZm1L13ZHb2M8k3vBTNdiLJeK0Yv4fP/4IGP5wZNniYQfn5DL71Fpr0T0Uy7OVF
utIECns9TMkETl9zgybI+u9aEsAVvsJ9cb+HAn5yThT4xw1Oejpf0xUCM2e8o04xOXg/c9exTKOw
9jOhn2RbgsqcARUVbBLHvznbxxV/G7tcGvLFcsj/vU6hvBJv5d3y4fQD0EMApal1mRwac7djV8zu
TEpm+Ox64PbknOvu6o0L0WWH+1fxN5beP73iG59OMg1eqXIFKpxpVLdHqOmwuvnnSyZ3ht6qSWlk
XxUuG3WgNsM46Nbs0PYQKrOHryYa6BsOXpYJnlLSJs2mHh+eXo1y7Otdmbd/jRXohcc9rGhJiy2i
N/XjT7vABShvnTnBXtmqUAob8adAiStD0GAL4MlPRxLRalRMweVj8Lk3YVznv+aFUP62ASE5yvtE
22IFTND3JBORTSKniXFWaEInNwthF7DIsj5jn4R4TrzDRdiC3MkvkzzF2DVobTazEGz8phXD3MAV
hh7dJR+tPlI2xFZVF/MSh7aO9vCb7il53YHuXXSs9fOQZJaXGY4wA2aqclrjS+HlPjq4gF/ZIO54
o6OgM2splVdcW6HvD1A08Gpiq1awZUqznPzhe0iJozeGeEqkZNj7qkhWFX1z6dFhsnhYFA/LDfZy
juExjJP1NUa7FM8sRHFAFShWh9ptuqCGD+UERJH2IPDPp/PHf94oSaEb01mPe+8AKMh9ETe0lIrf
LLpwDcqE6ProlCd7v9x0JQjEw451CW22pLo5sLyWCU4y2IISjlx/LhTYytb4rqiLGoEOlGc++STQ
gDZP/U08Xf2Ja0Xc5PIZxvBb/QClcBV44ViGR5ikXLq3Gxm1Bh8ajIpySL/Gp0HKK268/+R6oQLh
Jin7LXr0HaxjCZXw42Lbdsu2hYYUFY8kI1Tz4QX8FO2X6bA4rFhuJ999dcjdS9TffvjuoyorcX+H
9BNHl9gABYjz258gIePES0BBLju1gpNPatVoADv1C9hWY2+ydDvOAMQNqGPEZdu3CoQziufZe0L7
sv6lFColHjZV5DU/GtZwBefgFld/lvqI+faO56+6Tc12h7SLSPQCg3kR9/PZTeHAJaFLUajktwrT
QOoiEP2MjoFMXMv7O6Dw8VoiE32m8/LvUioiqcYw0qkOZwpIdfv99zzPTfEGVIKBs+OoyHWnY71z
+7ATbUwlDw4freVLZzgD6+2v9HKvCUU8MduT7CbS4CIMgZ90jRo4MpRnUdKuSMa7+mVDO0TKz0H/
a9VI6ZYYrvHuwqDIrCnDSPtkMReApe6tazLnQEXfwdIbS4wFUCget5VYGl/1LWQpVf+6riX4WnN+
YoElxApZG3MYLmAS+n5H3PPqxSa91ZEgIrRNejl2qzLSGfdA66ZcwzcA88PAGkmkJJ58gYrVlqD6
Pw4qwbS9qbsXwpcf6br9MwjF9wl/FlWyGeTg2zmR6I4uR4MwbyTVwGRl3M+UFoV/9grgPAudeYVF
ToR1sHtT1uD/Orf8CXOfw0uHSme2bd1NGffHxd7j90OsDxmvBIwxkDPl7NtDiu/WkE/gWc8XKogB
99Fxh5Zt5mE1R4piv8U5e8ysZITotHyMUfPGoONgjKhJLcjg5RdO99IMJFEQF97R6VpGgGaDyjf6
XOUvKX1G/hooTpQ1Fe6H62yrXt8AnkoXgW9S/sbtI1SH4bhYf6tOr76AwfOcZB+YQRI+cbAS2U/H
xgix0Li9hyFhM4/KFD9CyPr/Hko1DB52VmyVYPPmdJYVZ8umr9tV7Fafz6xARtDDG7de6iNBf0dl
ibQ0g4aC4BYh5d6eCH40KdlHRHo4n1lGjS4lharg4UFaIgYL6i9ZF8XXc/Ice2/Xf3ew5A5rlbWT
xEnXaxnuUPKn6QGy1qPpf5CCOnR7L300DAUCbQIIpDQ9rNF5uIhuwcl8cHduC7XE3uXOJuhHt+rN
KY9OmNMo+aF+Suj2xFYCS4TSOmfphxirhJMofatdfwkvChkN3aHLHbjLt2g5SDXQj7vff8nZZ709
GeG/lCtA/wCeKGdPu4EDVNlIoPoRWv+JhHG4ZaJWYLwNxYJ3+vFtwhIuy0wV7QGxY4Ttq9QNqBc0
7LeE9C/5gr7Xqz1sQH6IgV1Qvyje/jfxQAvn7omgX3EF2ntUkNg1EYDfT8DC0ZDbsiOiLzj6U6u1
q+SCRMQMmi4/7EZtSl3+RMUVWC0MEqBPobXE9+A2n1kCsHDE+tk8Vjfv0PFzpw9TUImfwW1bnbRC
ijJBjozYEddAGhuffZxTWIvxIjGf3tYSaOxuIMmxLkjjXhW5u4wjwEdodFH87VpZh9dFia9cm4ux
Et3zbVPYKch9WBHasEAZ/vqAvr7tMvMv7dHlkZSFBHq6RHLgBNO+EHCz0YNnbXUAfIhd9aNjrFK/
6hhxOQ3EqSURZHHm+8+wKfgOCqqTdPijXd1tvYQ68pd6CHvvtuMzbTWbrq6Cc8m4+HqzXwqX3n9o
bAREddHB9mkkYUSAIFichFBu/rtvfc18io1bLesHePydyL73FM6+Vpu7tiiATOCaOf3QxwxllOSW
7Ekd/G7IgPSRx2/c4JBo23RGODPdQ2BHv+8TGBvmk5Ai8MHYl1I/As+7vpCVK7MkngUQU2zF8v8O
dHxVbaC7RT0BV8/frVcnnPsu6FTHLFqgFEJvlP9JcC3cUmC/AzZkMiO88nYSX6R4UthGD2/MlU8i
cpbSR4qXksyyHIEYMrmXd+jsvwAgwVs9HfCa6E5NuZBfly9ejrYkm1LvJvUAAQKFoYPl5ARy5hIe
Gau3T1sgXsGMAV4P+C05BFyjq6u/wVHLhif65KnIpv0mMKb7sj5h5z69u0A3F7M+G4kbUsQfLSAI
zFILY9wVmvueDVTJAvl7BFHlhlpUGQ7h6O41AWuj8qMcsS4jDsDCKq0qYVDqSUO7iH7deCcJnzxh
5e6wz0aNqVwv0YuXuckJs2ygY7Udg60zEpjd4kRh3Y6boeOI0Op9h7w3c4Hka1avqAam4lZwXCMV
XT0fngeLcCqwQctk1FfZhoLNXhnwGBwzrTkcY9KdR9PlDydP1mm7YtgxhG5BMccGmxq2xemd+pP7
ouq9PJLs2X6O1DXrECKehO0OWpGZjb2uSwBIO87PzqCl9imwHcWof3hoMAlIyV92bTsAfOt2MbOL
MD/uryx9dIMIFRJZKRMBBJec28542tCcIDjW2aqNc/IdGpD2Qf1k6jCg/YsRAl7a4OOGWQaX5Pcw
stgzCViRrYiYwVzMXi++3BwfzKpRinpk8AwQh2C5utOWY+qNff9oB+NU7jKtVtVBnbQ8kzG8hPbJ
f12MxOU3pKyoYh++w4u8hceYoQUipQ/jYTrxQ9i5ac6jihP8i6ZoTuEE7VTSEvrYVBbw4hRTT500
kc4IdduAEIvGILOlzQwC7YYQd6eprqwX0L5vcKwsgaf/GZpNTWvZiWShm6ptFt4aRhVLSw4J4plw
tWg2c677rjizDA8GzU7Hbx6VukFGTSSSB91fpcgClEXiAkjaDtGhahVGytNJbVj5hibnWkKTl/lB
EwPfqoXJL5yIEij6jgre/lQK+MLxNlsBQfQCZ/Y3WayblpHIUvQ3l17FKYR3azuKkZEUYkCmEaAY
O8VPIhXsBEiMxmERq5axERf/2x7PHImTsvoWYSD4t636Ck23usR0/kZcpEK9FZY79wAr53b6eyzq
E6lgXNljftfoj+yOfCw3y7tSA14uNE/V+llkOf4ciLySUI7Tlwgv9FmqijZMbjrEFJ34GBKaNaBq
lkXCRoe0kGU/81c1D3+YudgHVXqNrwZhP4j8iNfcIqttpYxn2CCCuDiKdjR7RGut/IgUzaubD27W
Zvg3jeF6LlcNZ2/1wYStWgAuBTEjCUiW7VBAFcbB53tpJF6DFMplgX3YUzxyrgzisq8S2NRNvqE2
S1wjv9bBuyetQIjTYQNwqf11y0e6JY3PiJFuoQaybVCxrNd9VcoM+zDu9eX3WoilYa4HqAuR5o25
X6SfE3EtOE+eCi/1OVzR4G/cXRYRY/6AX3q/BObM4I1RJTMgbzED+cJYGF2UvpFVOpsRDaiROQ6Y
F+jIgQJWUWn5gRsD2igM9zgthrD4JJtQE/4JykPThofKcDUG7srtRYj+FxbrHwoqJsd9QrODlVhk
ijgUBDieF1ndxEEz/iDzKHzdDY1/T2EFMy0TAXfRqGAKJ9tOzRoR98iN7gMqfpLLl5om8tEG0iu+
u/Cd2bnCtNx4NtSrEdmOJ40jYi0G/3OdqMEX52ALPtGpdlj3ryJin0dsOsV4pWRKK0qma6mLrPsj
x+324RC2GCpsIBE7os5vFXPHeH/sj10cfoReINTFWn8+G5ynfSx3csZ8m9+OM0Tm4s3TkPsnm7Xo
NmCByE7UNF39CkZKaMHxieS7qy1aikwSMi8T/N80j9xgiY/REOF5hez2bqsfiYkiXbXqyVUzXAIl
Pqbgdon+OOSRVpfvVFSvxLWXxCZlpJs8NBPyRwGDiYzZE8AYAOaoDXt2CIbUvAjN2vXgyGzpyfH1
tZWgBQB9YbDDyY4ra+c642sMl7lrrz5inMfOJWbItmZYA/radSHXp5vmn2s/B7RfIOW7P38Xk9T+
VUN7MG4HKU2XqcDM5JEDLQUTf9LFr+US0YREE2WLwbbRF4z+a3pTdxr0kaiJbq/sn4Rh/LtLL7tY
BOxaFqD/gB/rAY2ENQ07TemfbFpx2vRyNJqGbBYwwXXNItNf5DfwNyxrex6pMgymcVgMWlxuZ7fk
kusNlsCJr0K8Lt2YQQizTWO8CCgJtfxlZaYLo1QvJ8AEJyYEtezbE5l1kmLiBYu1ipH42Bwsymf+
0DTsW4fHI5ujhF2ZPNfqUT4Dt6ke/J5pwOvwyB7d06dKxPo/TqmcA5wWre7m1gfN84EXNFjHLpVE
dniVT/WSRLm5qIWKFpisvdmhGGywbJe/H8DUeh7DFoVQ3RNasYLcFYKFxneZvI1zRo6tWiI3kW7+
yzroMN0uja9B5noc04aqvb/u5EgtW4ShUssfWVPdCYl7Q7STLDhXjcpg+/ZZ4JCjbZQruGHO2tcu
oeQ/E19LqMEnZ5DNlMYs+aoyh5luJ8ilTfOTEjEe4WVj3HTTIMrHfg4+8hLZXwV1LjvfYnE8HTDc
buiteN3hcNMTZ7frEYRLb5qbH70jb0PHnYGABLUy9fCsLAYcZXrhCneQlLSSETSWd5uZKKe0nm/N
R7e30QVtHepMVNe1mgSyzVo2xJkpDHCJ6y3zO6HkIB5jHJVDFhcUC4x3UzToAEDuWpssr+RzAWcx
m33mINo3xUvkI0Ryi0yxcjj0T3q3UW/aDXPftoOfqzDYWK/44KMb5SV0cP7wq6JOSFv/7GrM1+3V
MzH8HWiRG6XN/nJgfpoXwbbUsCjdbTO5aOiUi4jwR9tu3XduvLqrgaS67vRTzRzFehSyAREaBumf
MbbJ7K5i9Ude15+H/FrqcjxBKe0GUusN3U+nm8eyNXC64q3el34/aDLVvOe9eDqP6V91unQRmvdw
NmBqytn+Kp+YnCm57AiLhg7V11YLo2JxqdEYyzu7qFyXjt0RJtIMoVYZdCO3yWHCRjira4p7iG2G
aiJCFoqZcQScTDQIbG3QUvFFqNpKUVcZCEtNysgkzv+f3s7NDKGXNmXWhJnQRvPEqFGBizqTTS/V
LIflCxrIQ7GLDuvCK78zC9RLB0EiMDLiqiVZ7CdhtHsOZTMXKOCJqM7VI5q8D5QuXQeP8Mk05wjV
+TG9YMU4UAxgoCTX9LMEex4yN6ow3ZFD3q5LcbiNnDWDuR8RbZtvHYiuH+/ABZ+53pmVALH18+sg
NISrxon4sb4X0hx6AMO5brag2yfFb6bHvo/+n7UaCQ2kbmNrI9UvULf0hMRL3p38btSpVrOxwwtk
bm9VUhsJdQplwnKTUYc+cDLK3B8PDzO80MJeTUXWrbgWIhzIZxT8oRKgyv1gNLrVzgpOUabxOxTS
eYRo5TYMdCI27JnVT71HwqkZilmsLhs12vY9dC/ehQgaShjPTKhSB2e0WG36pR2wWdNGLyFfcj+f
BxWD26tSSt4xcq9hGgTLOCnUAseQfUnwQHd9em7TB5FF6ajm1d98P/iQPMvi7R2JGqXC1oGPJ95W
HGnz73Vh/haNKfTaQDzoy01Uqyw704cSs9p86cWyOCfZUSEkGBWgUAlDoTPCwX4vhXHytNarIxYO
Qm2cJM1G97FQ6lX4WfmifmgfhHPqN8q0KU7HvvWEGSQkuHW/GGgtW9CGg28jGBALw6nhGfIgJVlJ
QgVfR/FlaO9M3saT+0b/Po8+g8NlDPlFXiRg8b7uNoqM92XhzehD83Q1zoRkQcGStw/Ze5OBb55o
LbNnrNmFLhX5rUJiio4h+d+HYfQRvTBE+APySX8U0TVzK8eu9AspiDpnjR9jlDla4TI8Q4YnQc/I
W42UOWyiHycMzdSZA+f/KLoYKlDXeCuD5a8W84058MS3s5b7ED7XC90HMzZP5pa8Kq/PoDGMpHiE
+tc3lUDhjR3xZkWG5yLb/QFoX9esUr4XGOp2YyvJQOf0nQ6v4ySDw8IVFbwAbwnx+/mu8Dey3SZ4
tu0EegK4Tgn3yuCJVduK8cAL/wCG4t3bPIgoej3OsdusdbXNzbfMeNrpoRuAiYH2zQRcZltitwqd
2sZg8izKiPM3xidhn5LUYyVLPyU4rvvKIhijrnNVW1AShhJ+/0Tyvz3lKANCnCr1kF5krVyx9pZN
qAwuPHbYcOFF6KvBixh1N77wNZ6fdtNbzWxbNLL/eUQg57YNMBzYVJXqVjKS5LspJYBENSD881q7
iIQRcviQWHEtgQowkGxdIjGiJPQ4mW4IkdSNKeIjHhdqsvMxAMzAfYA1gsocj4Lz+vM+xESed8Vq
1wxrqreQB6kfZboy3EMd0R+SpPSNzVlZHc9LexdVBqVQBwyEqdfpvzNNHFqvnov4mpsA/zAydzhy
ZvoJJ3TpRMm5e+L1Nc3zqQiX+NOPIygBay23MAs8lR0eo20sKK9cElcN5fcHwqPCfjYNU5y0He6Y
1lzMo/Q+uBWEI/et9pACwc93RP675Ardve4T2C1QqKHShk/wexy4ugw23VEVwSobl7RwTbvZbCp6
moSVu271jSt2A3tmd9eCZPrIWN1nNyHgxBhU+EcG+2OCzS85GvwQ8qCl72s+Dxx13K1zXKhO60xb
nVagl16E6JPLClAJ/XclYq5njlEEgg9b7fgkkiKFIwrEuNRwD0W2fyDoZg/J9kprXvyLbTiPIQQX
Tq+MsOp2cETdCVnb9EQRvUArEP/7ZVGtByqpE4aMrju8RTVLmeOBRDGHblLptzCSUeon4DkU+H7/
hyOgH5DZQndQtiXUNssM9g4J/ONYGQKJAqhusrnx7TsW+wykKzBaF83nu/DdK5kcLC2s2E2GKZXL
UnbKpqCAgejGJZBFqmGW7bYLtr8tNrVBHRcGVlwBE2pUNAwV29OQXnTbczAJNsZF0OZlBZ7O6hcZ
SuT9zsHGVv3t3Wo/FDUUq8hugRH+lNHfEhxURkrJd8LSDaFSsZ4S5XYojP3K6vcbF9WRIzqKXigj
Wen0TJxp1R019XoYfqOYep2iczEPtUU1pKaXskgt7ZqzsQjhCFolLHjZZDhNdJAnRZ4Cr4q3It0g
FvKKtgD5Pq5ImE2QqcFHlIsSrLqlAIF1tWt1iTpju/wIXO3JDPvqu+yqtFbvS+z2BacmUosil0pO
QwqFC6WOtHdVBPYGGAwPZpE5RGkH6P1JG9zXOXuiDKugY5Io3S2UhzrDXduls+s/Olcdga4kels2
NjtG9Hj/bRf8TJI93E31tlhw1bmfvPLaNRABTYHTtIvt1ib7JYFYE0AYLgIfz1x5bvBWX0ijsOLJ
BEl09nAwngOnhlvT5IR07ccLXIdbUMkFNCRN2g7BGPClDBEn1iJGcUDowe1tQ14XdyYzFeUaUMq4
3h49wRm+ViIbiygzUH+e4oqWsmo40BlDzetm1S2/uE9gjBxKyC9l4Bba5voKURkH5i4s6fJUQKoD
Fu4QOFtm/dSkfStfwul3wTvo722+M6q/FMquGYEkg3vZUXjYS89DDMxMSDBcY3xp+7bcjZ6/xd5F
yDure/Rs/l6dneUbnW/iuHgtATVvgPRuinNGxqhCFhymdxE09zHmrmRHBUkW7wqWNcDQf3a3Wxd+
3Ca0tuHb+02NcRAK25SvYCyX7a5KDS7GNuril6F+AjVoiCQMNS0BmF/r/xbisJD2Evj5Ret9t23Z
0QM0IIcVCGFun7lcDIHAaZoDj/3v8CmHAu9QS+4Gmm+k8wWFwbiJepwzU58nW125J/8xJuWELcm0
cYwJD1JVCPgQ+ipawyb1XVkKQpJI3T1LRbgWqpZBbYUr5yM+pnEHdyLxbooQifuTNlFdLdyBUMVa
i7D3siz1y6Gjc9/Hl0VcPzRyaen2UL3csCMNZT0RMs7TSKhaWij/985k9kET+xpdq4AY2epX432/
sqLBOyteR9eFOaMebMbpwvmFZ7kbYtxM3vQv28R6+l5QkwkQacsjZDTywTXIiPb2fzY/pGaGqS1n
IXdm5qu3/QqnKDG2NLUpEd5JswqukhAfHA3gzPj4PXgDdQ3SCrFNVOQ63pMr5J7vVP/4eh8K3f+Z
09bYpduHgALX/QduyPJTsOrvIu3EcK4dxlrgwrJM3KgpaTC3aFrlXVnbjGZmJQMXhlKJgx9lVY2c
bHOoD5AKGTwmuodIclnTeysiQrj4Y4fE3qOnOVm+md2C62Gmb++BmLZn+jT8zTFWBViyUxsASNU1
jHyxgmgDbYp9iLwYYgW4QoPGR/31XEFLf7z7pt12PUIKREuLr4/AbLy4lybeLs9Lqf4G5ff8n1tf
m9RQKmugoSrV7xbFhZG87MFIT4xRwCrVa8nVEDdGPQKObA06ljyArXb+Ppwtd1bmtSGU3DaC6zvP
mG7SLnZ2wseNM443jpZVwH3IJHnfNc+EcK54Y3dpXp1N58kcjNmmr00z5WjdsSaNAbvELGf6Yt4W
Kypgz9qqOdE8PY3+IUDIo2sAuGOc7ctqsUJEOvlIlU61aM5oTwhSt9YPyPXWIC2ct/KrSj70C9KS
/+Zxzu0gb/2G7jVW/xrlgTBFGS8IqC8z2ZjAzuHBmTYTuNiHlytWNs4PWyJRc5U83bi6EnHTD/TW
eyL6ZDVK0L8HXJQAQrnLKmK2AX8g2P7eeMsOlC9WWvunUdLKAiFarTB030qnr9raJ5CyZFNv1cTC
vYMM5lkXlV6IyZYzQBvL84rWQ/0Kq6MOqcD3SByYYfzXfhdz7lJRWCiNzmgxgViGHWxPDqiznIxW
lHjbq/1jIKdNJPasp5McuMkUWKNbg7+qnhKsQTCPnLLyqHnV827QXq58z3M6/jFeR7I+iccv1s0F
8qUbwJChCYffo0mpU4SXxYcY4RU7gKEZL9CksI9ooRYbKc30/JCU2MWoylsvc/bnVDvRg0alixtW
2rgSolDDb4ClW0GDe4lrKB7A02bdrQd8hha2nz5fp+uU73Bb6Qzt3gztbzxVimD4W0UGuaL2hthU
WbLAXB3+ius2VHsVPLl+s9ZoN9hDr0uR1pPd8UjynCBXzcKyfJHSD/M72fMfvUtV1jvDO+gXxhUQ
z0hyQHFiqZNzX1lluEET+/ASvIyod3JjlpGnyqIOWOukOFSVu390GdEWMctQEMNi6mIc7c6B1e8e
kJCe+YDDtqYgc1xmbdh/nDpeNLtgSUZwmKXxCupl0fuvWJbej72J1gNcTkDFIxUsW9qhs1CLIYIK
S59yLJIKUshf0tG8zd9EdHY1mHtsbBfFi3mD7EZ0MuNzZcCFFcprNOYtUcLkp02dbMGCz1mhIJMm
PrA8zXzVZ9Bp4rTC8sioBeTM+hd8bqBxOTzCW/w4ARGXIvUT3dYedsfCUAPXPmd37sVg7U6FvvP6
Y1yTUCqpaTe0/+FKS9U29SzYNzm3IDBHJ2Fyp6EjAmDZYwa4JU1nw5UWGw1ZV9Wa5tVOnNmKgU7E
i4gJAcHpADGm7EFo3DzE+UNaDAw5jt9iBdLzBCUkKltXQsxmd+72Mjtf0Lh6V9FkBBKAq+I4N727
YgRx9j0oyeVduDyatL4X67w8bze5xOkTfGtukt8LhO9nGi/FeYXvCWYjs+5AaekJUbpwATkUlUIY
mrJPclbwE6Pz/nicRewx9i/Bq2xAzhwLisrgd3RCLoeLIutEuVafULgwCzM+mM8/7AlCtAPbeKQx
6dnIOeq5LpkEAoIgLmJPUwRpvrIL5CH2X6nN/09CMAubmBVXxUv0nQP4/w8f6eniq8AdvIYOkB8d
HHWylVnmF8IrmVUdNJGSY3+ewOOr7+FWjHcmUsRMn2wlCByrW32HQla+hj1K8wEKybUnWV80vBCF
aAlIKUvTKVzvrzG3TiPjIUO80eQ15gAR0TNSxWJLe7oupY/Us7FOjYatL9tMAHpDC4jqAYQDjVlo
geZa57FfqWiD/GSHpRhqDfV/YLJ7wxQ70VHEiJtbHgv3MT69LfxLPV481rYLahkXpdpCbHqrHnjl
GJtXfAhngBXz6tok6g4P47Y0hrgZXO6afNEEp8R4J1UG0zLNbh5gzWzLvJrHTEdk9mdM4H/KN1x9
aSi+6jlOK/5W6TOIa/0RAbPetIEW1S7CoODSS2mll4VRYAi/I1o8t14y5mkCxnoF6gluOys3htEj
MQTHSRZSS30bvhjLliwG6MJ344IMrcWdLGBDViCnkzLY/hlophBygbVO3P/qjVixSblLYV/GNZtn
0Aul0Hw6ZvAXpdzaAKC3JFsdHE/O7hSnSnaybGUaph0wnbRpMQh6TmoYdg0aG3/rerXtF0QeWpoo
h46LPlUEcmBVQXQ4er4V46ENTtAdYYUy00dASf292Wisdvj/iFQwoWR04aQ2/e2fn7ntNZt6pJ35
OaHuY0qopVzNkzozczkUCdLrk7b6o4qmuFkj2zkdQeRGli8/e1Pvoq+1G0qIM5PXLKqvDyUeSzcA
cznEY3dG17Wv3hd+b8Ns5Y3N3q0YZFyWVt4dZXDxfYwLXv+/Gp3G1I1MDkzqhWZN8cbd7jp92qX9
VKRKNofyUzi1Ijfn1zjLkxg7aE8C2FyIe4YyUw+M/Eq6feeSAgf0rihMcago6H0D5V3jSRt4w5g6
i2bkQapcoWjZLMzRBHkzsaFyahpKS7CzDSEWZmVBPsMSRLdikNe3unlbG9EKhfMGnvdJ3TyJssYt
B+QFQAG3ztFaYzj9OYFN7APfCX5hPa+NuBgNAwfGuTRpf0uZttwrwxVDDFi0VeFnl6MPjtXp8sqY
uBpo/wFBwUFqexGLrbJJFUMqsCSbcCDnys6RERKs9FO3CL487eplEgGbxTyWYxGNmN023qYv6AtT
JSlrdL2WwWVbdvVefC2ma7MDiy7fdC+NLtyct8GZ6mlFUgrHdPmuVu11oTZ35DuKq6yWW2yNKpeD
eiwqMVE4nl2H3ohlVFo6Djyu0HjQnMXS6HWcMuq0O6yNWOXZm/bCk5uQgBITmPhgEytbeT6dC+pm
zE02aVduyle03umpXanjrAGvI55tyLBBwa4oz0BXmAkVMfLUJCKH0ZIXbsBU6uoVSwtolZKND589
JtaIqH2SQ91Q/Go1yIDCkzQAjiH5ioPCinMQIyqr8B5losLf4/xmJlBZHgIkrobXV5PGxdXVHvKA
Gq7+fFQGrUDXHtS4nJLKVpubqFKDXhLcD8ngmvX+YW/W1PK/HepezY5svivN9TyQdciGCJQ1pc8C
9DsduuzKqoQBHta4sVnndItQgmWyb8DvDms15Hxm6V3XZWMC5Z5WClNuwYPS+HIZ5VZkSoPNtJSD
Ux9RA9XBiJme0IDASxb7AtfU75Z9PsgU1yUUfRtFKD//kxHE4AaJRCMmId6PCdIux1bXE+8953j/
Ly/bXzFnIMbrVYDGitgSGNa4HEmCXMX0u7O0TGKwELQPTnJUsXdsK2/oZjVOSQIsSNuVKu4+gWeN
sFBDoFZcNJ0fmTqliNACbv7hRBmXMfkxMva1EOfdvt72CfMRSZtOanJ3oJjiHq/VfESjFFcx7qYT
eKjuiYq7PmqOOtgoFlKTKpPvojFkv3XN24EKfkDKUC13N1xUbBFMiXMf7dm7/vc5buvzSj6fBZwh
AUi47v3fZQEeoVqVYZ3I7UAUikwPUUbrEhsDdTYAC/lPtAA/R9KYw4biprrI5hs+r4BQbN37p587
76i3xgY1BVgCeCj2MpCtgz599xDvXGMO+tHXYEfwNIRr35fewKfKCUMR4795btHGgLapAjBOKvzs
Cm/VuYJnQDuOAJujvSdoF+ggEWvgwFuehO8x1hDn64mlUL4FyAEaH4ONnHiC+zTHef84vVwPmhDC
0HuqnT2a2/isbHbFj1lPwcZFyN2j+4F8cXN8LA0XGe3WfUKQNlL/skp496Hthmb1WrnmODZL368Z
mUG5racniiUWPU4g5nW25IRJJBrjC45QHKlnFTLz1NyaRol38DEI5MohxEMFIkrJ0MPcVdAjlMeC
6NKIsi1dzWEa9UyuAbVDrfFP8vULOmsfsMyEqRdahRXfpPREqaBvfM/ikmYGEFv1OOdsthY2DxvO
HkAVIcZcTsmUYe5ZC3LKo+uYGGELIBbqv7nyF2VUPECwnJ9Ifgd2FZQx3MJU9piG/F4LwkDY8SP5
kx0/dZ4vMYRrEpkfX+Qxc8kCZ/MP6hto0yUlvuREY5gSW3fpPNj3JLhGcq7iaw9Gk54l+VrZSJCN
uBlWxEU1AaLLv05X/wv3ZHFk9ubNQ+zaig8xWdgrQYXputzJoD3gRJLWB2ad4aulnuvRJ2mQqFYM
+qpp3KRBDtiA/wMcgIZXlo93VUSlF1lYM6AAqGu7zt7edSBPD5N0SFlRf3JKLYKukdgJbHAcyS1K
izDMv2GquhbXWMka7ML3jCg2siAknSOc2c1lWsvXv5uW/L9sMnYY7mWAGhn0gL1eO4LoXJb7oO9+
5watTJTgowiHQ9nCvZevfB1GF+xSx/ZNyDL8qOE66RPVIMu+KTO/w6aVOdd3fHxwYHnJnJMi9sZ2
LmMAGdpkDAfoEvLNeJIFxhjief2palZyfdqeQjaF6w1KL5IfmVmlgsDITJoheLvN3JI0yPYAQsCz
hK3TmJVuKjbVr6RznNJBTQ4Sqg22N35d9Dq0R8UTBpGlg6QdYRSxAFK78JELifgZLRE7VsfcbUfw
+NArs17lZvBijRyvqTVHTs80400dGi5vcFqFlrhSlDo3veWJXlw+wwPDuimfjwpsbEmoMnBzzh3t
/EIEK97tLBdmQIFA4MqRHdr/bv5eDacC65I5a21ByFmoaPhUXBkL1qeDopcEtUUKPD79WbMxuyKk
t79SScdQlZ1P9oI8wCYgbCU3mN8tWcwjj+Pw6Vy2a5i0SfzBghfYsNCccA73GwQh2xdJVHYD2LX+
M9ETQJJpvOvtWRAo4GX/cD9AgExV9z6NS/+TM9nO9ZtOPfNMbfnHKmtZnauHH5XEvSvGyM+TnPTo
7RRIvax1zs3ebi1SunnSGv+Er7QKxkvBvxRTzFO/Jc5hWpN3W6DW4ckwsPVlYDG6l6ijpJErm+SD
vT/mlF8ihINIhmWXm//8SivMiEYEhC/Q5mz0tGgIMX2AFCLSOt9V0QUApdoRqKxr3/VVmTCCM93d
eGYaY7Bm0VAlPVY9aoc6QerfYC7IGTcYE6d19bRuFiTVq4rX2DljK+IJF6UKVO0WxUo23WNcX+JX
Y2SdiMbRQtHvyWtd8l0tqnaxAQY3A4r/0ho44c83osQb66faurbI6Qp9p/Y5o6HUdc5rnMvRO3qI
6r3AxOrbT+XNWk8P0beiuE73+DHPIR6PkpYDifKc0ObecEBLGrn0rlWRoXZnXMy9aB270eGKm1Cf
1RrFcbsA1BbfVZTm+tL0dyrrMbacPliiJ+HXEiaiCSxPXCN9kK/nnPfcVmGE7e5DYn7OYGsTW5RG
reRbLSJ3edgl0RBHCxZcc/e/fdn6vZslaBjWomMECGqEfdr101ORzlQw38T5R0KLWh6VZ+ogtlZ8
ONroZaGowoyzv/cHeL9j22xyXhL2ej80CBHE1PKqmAhUYq5cMOSEQdO6bHkJHzHjpIq5Bl7EvwD6
RNRIk9n75DBKEyZiYk5Opop6MpYVd7t4oz3TcExoHYDYmqUz9mDxxRH6RUpu0JRjlF0LkXZaE0/L
A6kH6jbzkLmdaKTeKGtiXAnaaciLEA6k1O7xgJlWHBG1dz4556B9LAfrRAhYzlGdDbdQDcFwUf97
jjn1mLF7FY4SFI8vrKZCpFsPiMNIPMSJTpKVXy9GnyPoDiMMg3snsRMQRzOWKoN9YQD9ZiMinaFu
5kzUutGcWIcSkrGYYcfqdaiUWYjvS3WjsjhOAAlygI7y0AbfPXMqtxk0IuYdxbfDK4cYtjznDwRO
c2vkSIqNwvEL9u3xc4VkCVwV7V3F9AxORaBE7COZfJjB/2YIL2aTbI6yPKw/Yk2ohwjU9FRWjht0
1xOoig0zTBfIMmo/g3+e4+yjApV7DoshFN1+1mr5yb/IHfgUgkz9YHk5zPZu2+Lcd0B8Mp7QLs5Z
Y8HhXs/4w5z1IwpuHqc/G9TlMmNAwVqsFMCy+dRr/fY6Wn052txqZN9w1qyjStEYPeTwrbmcMYF2
gdLIMKMzQu5oYBRggaelGahAvWXM0FStZgvmohrJQ6POrXDY8OI8LBAXVyT6gomoMx8jE2ohAGeM
gZGaxE5K9Qe1Q8mhVd+R7m+cC/ASv6Bu39max9REve06d2VCI2WEOTYro+8JK52mwAgCUtuECnxF
IZf/55audd2CBMzMSP8Xmu1xu+eU0anSPpp3QtosomfSOei+AT6pNdDuE41fO7umc2RR0Hgl6eMh
ku+JAphQtDODkJdFvx7zLPJ1cihibjWPNzpERfR3/J3uRDiIuhQdgR70MlFHLVThTzGRACfwaelE
6smDHynXh5WYSoDLC1UYjrLHTLOvt41BD1dj5xX+zTFO/CgZgBhF2T/vjROMvIhtRznltxn3BJhY
16TeYif19NoBNJPxh7bTPis8roS2GXlJgo0Qk9Giw2MuklRsd7M7E8Uv7BRs/NPH8NmLwhM2CyGx
oL1PAxn8bOU/cX46LO4k5/bisCUokRKUgjRnRroSrnVejtkVJWpWUxu9MVq1/nMq8Lh7OM/4VU8B
rIF+OKdpuP+KClITMsCsAkl5CQlxWZ5hftsjGO5+1M06iMzo9JKnHry82phhtPIMmV6ljgJrOSen
A5MTa7ky93eDFI8CXEKbEQERWRbWpgxfJf8bnO8VGA/DIdsfE9z+yzBw4KOrWzRyybkglUlbkqCp
VfGbKuXvJtr4yVx+FVg1Rt1OagQuIn5uEsIs9yQRUfK8jvycmwP3fXwhCA/nPeXcZst8efr0sCG3
dMEQHfxITKZx2xgqzpo9hyd3p410Tk390dmcR1HcCCQdLZtNN+597ludr9g6tkcULSLDHMJN8ZUV
5rWPbbTeq6TJBEZcnmp1iTkrSqi5JyUuY4PIZE2V7gIcG6r01AnII4USMFw1g0vTPq+7Ph7hjVS3
sQ6lKqmJKxz0jxMCFa2/xdpaDjVsHseaPEjR7SC+PS9VrZXpqdSzueUaCpk5HN7lQ4exM8Oom7Tq
/QrY8xy5k7jof+qe+TJNEZH3qMnrDxg0fXVx/ZlXmgee6gEnCunLLj34hg7JEnJMkajloS9dDD8Q
cIH1tHHlXy0f9e796LOviSquTv2u/fIzM1dQ1ojToOE5RyanWad584knjHVNi7PxaHOYv7QY9FvR
gP6DjssqVnZPoD2dvY+ZYEBxVkYfUKgRF32Kedeh0DFgDt6Lo+7UYszwRwcES3MHRCpTXx+x92Q+
eMA4wLyl32R4YMpdVR8+zpSDvmLZx0dGD/h6Auy0JyJIL1HOsPa7haw9lKJn7DGAiQIKkmEM6wtJ
O9KwgVMbXQGGJtPtreNbzBdzPKQPAdW3j89zQhFf2ybSCJ+w1IQiIt852zqH6SQgb/IkJNzg2t0O
IWdq/081QaEJcT5MdMNQSmHgMpejMChm4xrZob30NKA9nBHL6WO0ZAcMUtY8jTJMDbMxEf6rqX0D
SdUK56RpqO/q9VVrdH52zDohncwowWMMiv9WJF9qAOsACQ/XzWF17Clvm/1tc1CzZ69YU23k8bdv
HEYZmEZTrvMwl7Dosulwe8WhoyGm0Ot4aAM6/4/wC4JZ5Vqwg3sR4y9OYw5srN5UHWlYoIPUiqqo
6oIyUi7/++HzQPV+u4b5pEan1da5UgNbnnvZIBslVdxseFDixCnDPG4okR4do20X3z7TwVHr7Uh+
wceANT/RPWpE+1b4E8nSuL425qhlUu7MMjVQvsGOctoX0oSVa1UV9+hqfE3JAYD8VBa+3Vb0p86e
p6g4/iOrapkEzIOCcsvXumiJ5wtNULwj5lE/cQsAZbso4m8hrTOOGQfopnSUjCdZI77SNPZ4KYhW
t5eih0PBu60qYcU5vAZUUUsva/Ij6Q/gqjNz+MEt+vE/xDTWjE+x7DrKhj9zW2cwSvRzsmMAsziO
JbarBrFogiYtT113pLWwaP2GuHltMnYh2XS8s0Ho0XRl7lNCFtQTWpfEmwqE6AK9ChOLkC+qZmW3
J0BfEW+bgA9GAUh/JlwL/geCW1JbpaQi6gRwsV6ibN2kjszR50cfcmOf4WJaAMG1n0AjTo8Z9arF
CdnxDn3CtPwp4NU/cSLavbxzFrp3scQRrc145pCtvN6LD5rf8+HcUPZNDJwe7nZ/4P5aSJdy7KEw
cGDXgH0cSherjhmKkxxSqs4FF+15mJP9teKgWQo2hGcILYAP+IaCYmkh/LJ0AvREEBmbew9W3cLF
UdAkIDwYqHsh0FxBb33wzikaWdroo1rUlZHiniCc8oJ/AN5RHxcR7zebowZYzJq9o6gsSXgyrR53
2fhG0HO4eyB5sxthjL7rgB39VhS89t91uCdEB/8cQ40K63eTbwRqHDx81vvU1PQmILFRcbyMr+/I
tuXB3gMfbs11bgH8TtiFsQuisBMPJSujyfIjGEKkQ6ZXw0RV6Xs2CdKINGhv/xtpzEFrAvIFhaMH
aVBZzO3cUAEnhK6fBQtOkGZWNWuNEFZ449dW/C1UY6/U39/G/pavp4Th4FEKhVVRant9SbBtMbBy
GFyP/aYPkV8g/gV9pr4RnwdYaj4XOvRrwHFrlGI5QMiDWfxvIhdecgFhBTEdO1BH0XEKTi1WCnuC
Yr6bV94c0vba94NoUlxwk9HpwtJsWTI/7VNWwHSKm5RlTP/TyQXBcR+/ObOWY3PPBQMBdMbbVGOR
+dAohGBSUYKWTgeGGrWEzk8PH84MqS/2Y2MvJvIje7HcSdVSmQRJOQl0SB8TLJJEHiOcYu6Z7iGA
NHYGIkuG7ar6Dhjex9ZyGvoCCwbQxCScoWUOQ0/lzbQ6GnXoBGKNj7LjlXsEVa/50gxdH32xzGRI
b7b+Hae8yHWd6U16cvEVqeuhpy3t8DFGKe6LK6z/zcX0LZkFvnTb0aMq7DAMgqESxcPMm21Xdjiy
21EoczhFUBDR8Ap0Uaf/CZpv0Kj4zeBFhPVpqpc1pj1gBXQLNMzM4CkJ5RcJHCdupExVO/UD55yP
SLSrLTpI8MBAq7IHxHaZVt4zr2bYRtPYQGkTENGZo3KBgquW2mi7lshcJvi+f2SZcvN4yeN12Ymd
wmrEHhhNKFuO1lU7mo08ovlLIYcygQXPOG4+tvzM4zG8M3sNzGdGfoC4tqr4UiYVHsIBkdYwH/ws
He4kTjvm8dWgq2MvhNx7KuGY5pp8iyK11tXKasReLCr3klttd53VtbL05/dWlvR/uAvAyrw6hYRJ
LPkqOIz1D8TCQsSPfOsYsj+/XvKC9+tZS4kKXhkfZWKCe7fxkeaZEqUuBaGT6Wr06jHMEXiKUraW
n9w3PGXT0RBzOxUeH3UzLXDNsKpVed1eD4lXSG/IeUTNxEKsxqdJJ6R9wFj9RQluGxrC2swwifbo
cRCMSsqq6R1RGQkBb/9F6W92UMs0WhvO963qs5AtDjOxcVHyOYd/AK9zW91pHIHbjXQ+WTdbL/AE
tpTLdCGiJbr6G7AbhELo9GftqDL8/UrerU2ube4kh87/HN65VqNt6z61w1xkU0Zv6jGo4QeMHsp3
X1S8yNLGuPDgW75tVGjPz4JYLBQ+qEZALCF69RD3gGlqg/Dw55C+hsA8DfiKb7aAP5WtywI8TBKI
b4gq3DMfH5NjcAbN3zq/dMgyght9nFz1UFKlTr2piZ+ZfjyW6HpQEa4B5UDXOkkufD4/3tSeGTph
88XCX7L0rBWliAkkgIXnWnsEBAmKNtxOe/eFGuxL2pW4zGFNogP9su1TpMAbQDaQ7bufIOatjlSo
W4z1snOTet2hIu69XfMihCvBWfgUp2hyEAdZ8al9YtklYA5VZmbjQ729RWP859SXCWbYzITYdyY/
hsTRj1jwA2a9a/rkvzBtNJdXL54W+4y0Z2VrgSkKc1VgLDanoV8VNujVjtDF8qBLOEQgCQlLwBfy
veuliUSHaP9O95b/nLGTKd5jPzqAsaigAV00A5NOHuyl9pIEoHcaoI72549y/dPqrPuudVR7NTrl
dgOiXZjntrRdYdFWG7ezZlNiRDTHB0jWo37QePaZV3yx+6dflQN8gVTuERaRHXsvjSLHDOlnhM4/
1fzryJM0eJepKxlEr+A2t2QsD5BdREwV0twqeaGv85xS8nOXq9iJdIHhsiQ/ml955tFwRclWEcHa
U1IffojblA75Pz446o00W++IkVyPFM+k/5uFoKfd8zWtm3WO4Fij64RoNABrkejzqVvfVYWizUDh
QmKPljBSf2NkPZ2opbrkjTcmGyZS/Rlec80oGR3Zu2Sss1IjWIPWSlkCccbokou8szRDGOnMOIY7
ajVl2o7sLiLQ9FSSGL8/6wMZEaqAorx6gLV1dgUcLN7pKpRkLbHHNptCpgcxYRZI8C1xLBTttjL4
qMqG2JP4a/Al6i9dA/6TR+0l0dS+wL6cH5EBS1BPiMHj07UfIioU5ctgmFtFwsZrf3d/c0QKITat
BISq8WWHuFVoS9w7VdD+BLxjm0efsZpFY88coSK92i+Yv+kIMwpTLrEh9cQC48dsvtXR9w1jmH35
C2/7K3uihrNODl37wYFw+Z4q66l19vpW64+BEIekL1MQzYeassW+CdO/4Oa6GMbeNYngKYllK55y
Z1hwPZ/nsQXqQ8PZ3WTH/DRcB/qtbNdn7fOu+q9ztOsuxFD/54EQk9tUSEC3bTddJMB4V2SvMFYp
M+aBBPyC2W0Zaz/OgXCMjtYoi13lyKaJs6dHWGD32e1JI4V8+wldp0idLLFLSOpFCJS8CaeuR/Wz
TQGl6Nu8SBNds6MT36YygzUCb846pWjcgqJXoJN5Ayqe+72xt9fhCw9Vm+ZbNRnFGVY6FOJd8J61
URhYMLqD2BHkjoZ6QiHlR/xht4vsEvVm0NLm62vErNRLWCPxFVKRc+GFeuFd849vzBnyvMjESh2N
+gFOhm88TphBa3cfK0dhxuYGacOsUaExCqDdqSgVrqQUG8PfreufF4q43TE2TZEDkpLuV5pwL73M
PePFFQpqAPMyyR8PBjW6XjJH27Efzj2VqTICicFIWrGEfC61dZVpHPy6olBcqnZ4Mt5mDDRfPErJ
BIM1hHdmMWaWorkhNd4r8BaEbQ+ssVnaJI9oWh/AVygI+2URkKREE4GZwk5kOAnmmnlFxypyC6ZS
svAnXhQMG0F4euFAe0C18Mn7MYohEAJnlO4XIUKcp8bj/W9apJ/hIQV7ffUesjild6dZz71UolWl
iqDJXkALEM3Il9RSl+kX/RWS3NIrRVonrkNdVSDeQrCg+7vpDyLl809AKFDVBBPHBBVlZBjHkukS
9MXozc0mIYVp8rj2eYp4ybSuCo69NdX6tK+XMSTpI5/iikgeZzzcBSlx7ritS1TH0Rh4BGF/mQgz
P4+2J8LYvGV8utlTKIlhmzNLstjNmiI32DUkxaY2KuxY7cJC0EzkGIPdbSgxcOZFrpSJv3faVLOO
YYVoxWmjGuVTQA/dCHT6DSzUhppk0qj1E6PpLzwcss/rst+H0eF9LIWE8LW2Cw8AigLLD6D/R9ia
i3R7hKwSV42z8rDtBWwddOtz2sC0E5PWYzTzVdPnOrufQpsngg4a0yyrZsKQMijK+sF2YNPfms83
fIm3NlY6gtV/0IrNfJ+nand4tpF6eri8KMdOroLRCJviXM3Q0shL0cOMTaYujovpHnpAAkyRrfom
+k5I5GP2P6+MsRtP2+EodGIkLnt0AABG5G/XCmnGtgxysHivOV/Sl0bWFFqcz8hldHxr4+p9AhmZ
zAyMhF2rAdnpyzCxxDnvKG8xs7HB3hp28TLVjstlp8ynbqiN2Rh/T3PlJ41uxjPfT0Ko8z6y+PQ7
w9xI188PiAbeD8C8xbh+Z33oC/LFIUTpHysGGFHoUxz7ITOnKuqiD1KEEWYxoBcKUu6CCeSNy+bf
LiU/Y1EuVKKLX5trr7T8SFtfqBmRQTyTwA2C2oBUfSur8hlEnp5RN4Pd4nT5/5Ba1sFdV7v53qor
7XlXCJIlX2i4yNmVXiWgyyPZ4iKQ3jguolvGEHNIl2YpECJkwfrCGIi+Xmt2etrbIHvpjSnF/fIT
ZI+/emqbjCSxu/C7Lc8jy2NaSo5hqR/cFgLpo6jd5dFy/9tD32PO6X7ccOaI8CNdFRuNKj2/ZgAp
IQhGi++oJQqnovGd5xH2W6qe7+8epOuhx4/eE5L5hc53rJCBZz/74zOAkU3B+aCXTbTib4i0r60f
a31oOc2KdtwfJ1IqfB01c4x2vsB+ivMpEM0BBd5SgRMphxZWpr4Ff8sd2GBytBlvMFv97wGw6+kV
hm0hQ8YFVYj6tgXXeVkutxnlZs6NjCtFc+INpl8OwDSGdcNqTUL2aAHzUkRv3rz39B4S5yxLpPbe
txSQem/TRhFGs3RE0HP0whnSuePHR/yaKsbTNGAjCKV6wGWEiqKlagmlu09hGDKP75t33Rmdy6eT
uJuMg4xFy6BBcxDLRAdDGino2LtA24lTA04KFX/AP7LhqFip8Q0rhfHAnOHcQpCdGONbAkOHnssj
plg4f+7P2Af5w0jBgK8c53gaMuHyOkzMEAsgbwujuFprttaMSDE928Dhbv6YeAyqYq9kKzFj6dX+
hQKuhHy3Cy3RB18i8QxIJvs8560yXO68npJds9P0nKaNoJGMyYagz8q8+h1pg6Ecd9Sf1Ng3fdR2
O6/YAeZlVn4JyBW4GZEGv0o64iDKSnnZbCZUgmkegROck+o/t2ouS4fV6HfZKYC/bcOEQulAikn2
UBvcnLR3I1v8IzXbct2xTXLvrWZXWfveKNMHXdikU54MVeVCGWA5Rmwto4wSIrIikouvwklPyPbi
AhfBmTO+2j3hZUYZQ4PVz+QCCUdpOwkaC3n0cQ8CQslZWQ0x09IRaiHBEvaJeNRD3JOMcYsuqtNn
MEcRwSB5R5HwjHR9WWnkS5N4NaQhO1D5DhBX+y81tz3NTUD9Gx3VwPm7hJDZeKhJvbtDtlj+OWU2
wjmlyinQLddEF1Xg54D4LV7j3kIHW1G0n8BxOQyiGiZYVQ1QqT8dBCp+38mYs+mVUY576gbfY63E
F9+YLw0Qlu9wWVihKO839tObYe6ax3+RHxv4gqLu9nKI8i72ecivFO/qaPknYrlrhvd9JXFunExP
q6ZRzkJKcankyqYT1ybZP/MUmO1VWOg4G0+ESasTMM6aXPS95UIprt2mocFtAueQelDgL8llnSlm
q9n6BmrZuxk8rHoLt3GFXfOHltAdCVhNZFmGfHv/nCOYjWGNJVvMz5HN3ZzIy9xhKrzQpJAyBMwI
RhPltmfTuIdbFhouzt+XK1YH0Q+af7n9eyHnkGIZi9JG5P3TXDIJbkZv3fa+3ssK2ZgQ7pgRz48r
lvD61nOqxyieMpQCd8EH/DHrjy5ZQxKOAlhw8GVCuyMF0HpPyDDLSS/pLN0udNVSD6rqL2QuOqEJ
bZfH48lpyV6A6ECYQVoAQX3ARmsQvFOGVIM/Th5MxWFf81N4oJsoITRt0aObm47MNYyHKmdjsdUX
0Su060lkLuQe8AVpIGJYajHluuzMWL9MO5urnNZPUlxquHEiDK0NYynKO4tfYim03ddA1yTX95WT
qdcfxB4iQ3Xd571g6Cgvx6z4ClPXm5+ubjma4CF+r1+a51dhHw16E+xwKzCksXX75G4/b+sTl/sx
x16dOQ9tTwwgo1gPUktggARiyJaLOcbvURUKEsl/UvYNQYYIIXPVU5/MWENWQoAqGEhbLz9/WcEI
IsFJNYIw4BUOIqbju9sbV0vsaV2tgv7vrJaD8Mo8llz/JkwQqyeY+mviR3otmrtLJB1fL0Gk2rh5
Pn4u4sM3Vnyr0XFQ65DoyP3FkN3w3yKHRr5BvQhCQ1aCIADWaydODVOpsU+qIiWpLLyqJ74W9ae/
oZ95og3PpYNCE/XyGAQuLb7tt3FwonS6A6hs+sz4vl9V2IcRxarHFQWFC9j1TVjwtreeInw0H0Vb
e9HEn+7RcPcfjhNx6Pt4Fhp62FUdt0Xg1LxJbrg8LGqEaSriBUdBeeFwCPi2BHPlcs8SLc3Hwk1Z
dlD3D8XJtFlfRQogrkGQy3r8ej9EyliJwAQdTOPnfNn8/K9xgU3rX2NuL2uIIgWkI8l1UN93gG+g
dMYDyDqrjPX+xApfIyLxliNyqgxUge+zFrTfZQj/ITlsfplTbE2YKsgMlMr/LbAiIN+jzRcNRPim
YWAsmkZJvcK5KLpihIDbEKEciBT8458t/XQviJcsw/K0SXd+Ggm89V2KQAjpSgUsVguJQYLiy8+U
lS7mMrcqQS5DG7RwGdNSZlCNCH1mx7Xn0/IeVnBDF0sIv8sPBip0F0Wh89ouwOomriXOzu+jc8/0
UmJbg7aZR32rNQgVuwIdr1d0VH0GHlP6/TQIJu2qwkez4YreM7WP5MfBSfnAccOf5wfBlMWSIVxN
m6XxpHhkg/UstSaiIIlkvTrI+Eua07iDhh61yT+UZ6BRZRikvNiWIc8MkOGQ4BzGRRLdM4vUCJjU
V5APk4m7FJ+MqV9mZVmd5r2Z7UYP/VjZqogjNiVGpOWvxuLcQdyQJmuyB6XScYCvejtXMJ4FPcVm
vo0df0Z+5T9I95dXjlUzeC3oPnl1Kd7e9yvlDYvGH/KM+b2Tjfnxq5lMynAIASJ1deONRcy4AOzh
OLIxEvLwdXffJKK5AdbJkg04CHCHvM869/lE/w+U+DxECYeKSUQY3oU8rNxXk24g/MH8VMua5qD7
q8/4h1nQbWjo/5rF59f8TFkX7TcEJqNmD28w4S9eccjHcqLhoWu/KoP0D/IbKokNWIjOuNZVPJQs
5W4VoZRFV+070JTTooGgrfZSHRSrwmx5KUUgeAhP7y1GpY2FmZuYZWLlJdUxRmDGZ1P6R22LS9vy
Zzw8VSz4YrxFQVWgBVkEwhmUVoD6LpGO4vnVFrxyQDNUNySeOT0uzyWJP3lMqjGTIxH6L96E8jQ8
TYgoVMRdHj2Ax7s8vWnKa2qkrNGkGtGzVWF6SK7TgnZkhI8M0MjT3TW3n4ETg/Wlgc1HnsyS5dFn
tVfojr/trVoWa2SxjGSQMUDjTcYTxCwsn+kG05aSNPgDas4GwTggQNah6nwYQp51CIrzyuUiN1Kz
3ryw0GI6ovp+QLyn4JUdWpxY46JS0jJUqUaRETyNnXGXbuolpUjg9ndu/wXc7Khihp8O8K963eam
PuGhkef1GJ2BPIJOR9900tiR0he6ilHKtG0GgzNK1T1Nn7GkgpvCO/9Del2GgF5HwBTQpJL5x1xb
AdteJ5s8GCwnwCzG9uOUQH4VAJUr/0oHa99uAIjjBBa7Ea7jrL/SPhYHN5vifw/kO1Hm0CLBwq5X
goFtEaR9vem8Y24cUxEzUtRpe0YU7ZAhmyotm2cCms/I3SnBANnJPBErbZ0FXOW2yqu3+mGFxQLg
xcAVIW95++onDBkSPnAS1VZa4JQkR0ThVSGaWu8pC4/qqltuwnrUswjBB4xmExB8Pe0QgDnb/R+P
0TWQPzPqlEJ0VDrDONCqEZ4704VHhoFFV2mGDSxGUJ0BbDrpWHBUVNEdv/0aydfxtCXfG92CFyNr
f7Q4Y6+U2ofBfw3tMaMoyqBulsqYVlqD6Pm2RURT8o59q6IlnHJIbY9uNXZABAPVhtAy3bHMd0Wo
F0eiDThy4EV5IkxIIMcxti9xhebit75Tbtd1/dFdJTtmIkl8umTUWLBkg07yYccyvzy9F8U6LmkV
eoKumpn4SSae7s5YF0jLnFrdhh4TsAz7M+wPCvUv45hKI3Y2wAB9ztGlJc1BmVi7mfF42ZGAfdc6
R877OsAAf5ZFeMunIpJIFOk+YdfRfRh9Hbbfl8QO532mMxsf/yQcsSuQjNylgX7obDN+SWMxG79G
SxeLd/aTJ2RjVhgb27P43HjsQmZhF2dYrc3ccapR5m2UVFidmE/PH98V7wQ0Uy/ebePl0PlgtMTC
S72y00hbxPsnDXCl3AhtVZO6SSyoTo7jjXztJCHKL8+mer2gBBaEP5bJZ6AiVCDblpkfVBUfUeWG
R6Gi92pGGc9M6pI63Knzdgm+QtYksnJv0dxEHjwJj3bw9zKEJ+7ETDHTmZ6vaEbQw+XXpavJP6PZ
8iCTI6suURH2MaEnpysx2Mg2htmHDHTblyRhjAXKHv9cOm5CAoRKX+RN5Vz/Z1RCrVnnhRJhtMyK
cf7XnVaTjVxQzzH5TBm3l5TB27BFmKyTYtMEGQDzRPnj1e4hb/8BEk4ueTe3UhkLl6Yp4b5j775K
AGPwclrf8WUzvrM24UsHVh2mk4taTQnshXalts/ZFQs343vOgbFkXUJ2YrNv7Mj5pwimzYamks+Y
vnj6LddeC7EkAqVwewezolooTOL4lYFG+kedKnSSV4uBuhBAgzDqZsBpfgbqg4B2/G/Pc0DPbJvz
5COrYqRFNWxik4bcAjfKp6/J5aF06GFiNU/PyIyEFKXN/POoOekPoY9BuBbHwoad+slj1ebYsHr9
eSjhm5jcscjijzJVhLgwS5WM8Jx1CrCMAIaP52eYf9i8Fg1uinMeJWQ0eTbCU2wqLBt6sIw85okl
1UmO3ZwZer+6A9G2U6IDUM5d26spKTyRJTmppAwwBPZSWhdVMaPpHvlkK/LR8m/aPUHHJB7TLX0t
sHZPRJHsCwTkYX9IIPhh5UQiQYch/Cmt7wbTwZNDSBxOmrlz+zlUrUCxImw7Bna3dK8NqUE9CXyi
GcaVzNJYvYxbclmAaqtYMjtNpjZ7fFqKTt3Hv9j0ig5yygh6hJbSojWNGYlZpUjNlMEgPRgklJyH
A18opZet04WkWioZZYuE10M5gTos2wWHO+ERCtgHVlnP892cLlxMPaTulk+LgDjMgbB4o93aqZwl
ikukyNW6fLw5s/3jdikfy8s09VPtawvm+b2JScB0LAbFPpCt1IV8XLAH2sNWZ0txKWkQSR0DSrxC
AMTIXDm0YtjcMKFx7vp35HjQfs/eDI+zlOpkSJ9+iXdFgsfPjtlQE1d7WyCvbKVeiDzGGT2pgcqh
YpLrFYp0wiyiMRk+6aW1+L+I9TjnO8FWg4mPTqJuW7cD1jdAMXLhmzAlHB0RF+dpfOsOJqdBBIJ+
vypuhU5D/XunyfGw7jxbPAWzBCUB3w6Sc9AtrBi5UpcWL1Q8cdhYO2EOwvrkzpiWcidmt4O5yfdB
a933PScSRogO3cgHjwRjGdmGZmAttGkzVy0l4Ky7hUvag99/n4k+ZCU3ALtEDuTe2yCF7T2yijw/
iFTEdBvosMa5HUVPGba5QfqKQBsGWIq/x4voQC5YEgHy82A2vnPpI0JX4VQcIBRiD5lKVtfJgvt6
l71056vuHKQu/VziZuErxnx0m5LS+PiniFB94QsMmV18R5rn3anUJqaJknwEXmdR8e89nvAo+fpn
ZD8y06CtmX8pHdd8N5DJhaw7Ib87nsaFBj1JSL7hd5M8PE8qdMOqOufOfENOZShbz7mlu7XCxN4/
cn7TFeqRmjQUF1e+1gCFrjbR8goIYIJ1mlh4NUVg6iBrYSElX3w+F2OsPAoXMXWnIvNLI7BIR4dP
zYVlMyhXpf0vhjVTe1mz58858qoL6p4N0T4Aqtw5u573Vaya+SSkreHzXaDxBp0ZbeMfOIUJPXVb
08g7Hb7G5IBAiVcqW5td/GblnG52sBDrDjJsHpJaoKraQoG5hz9oG+Ir79lSv4ymGibnX4J82jZN
N+Q77VTy8MBY+NEOSjplGEizO6Cm1Szhe2Pab/VgP2yWbJsC7WKQqKmu0ugtckbj/U80RnIzCbZU
dlBUszyQVCj9I6Tey7wFq/q8ySyKrHwtpA82qtilnuUgGPCbTYEcsJ2+F6CQNrEJFlpLFzT0wGWC
vDtuVHQkJEnohkWDtd1hzqXm8+g80fIqHrct4aAdlpp4Gs9HMLeSCRBMsfnko3oCtFNfdo8np0Zo
Z55XMxDrnr+HyjxWM3PJtAjSXnJi+wTmbMOFN+DaTKyOc+49mFovWWtXcTwtestQVNIkklgi/5AA
YtsebofNuXc207fH/Rmj6Ps1DEJDtBubPoSu3Bu8/A/CFrauNosRSmxJX+XyDiJCDF9ODRDXAasD
YGbcMfdv+Gj5JaXOGh3GGJhyJlaGq6vRo559jxoXBFch1CzezCEf5R8m4ygDUwSaBj4DjuK/m3yc
XuLvfutDhW1dCeIS4ysaw0oeOopiGgBiTR6D2BOi+i78gksJKK9r/Kro4cIZSArfbtbRS8hzgaC4
qHU7z1iryIqOqDxbYYlfddXa7liX9PRWSf/LVIdYAZe8kI1j4Tw39OW0Bdfne/F7a8jp+UxYlI10
gu7GABvYe/QwS/u9lpDQV5706YbRpe8NfyLbbRsXlrT1/ZouQwlUhYkWb9eZwXj2dCUkPHxHJtgf
rhoQv+ChVDXfkGyhD1JLR9Lv9WOlXeHFhZEeg2ZeA1BPaWRQDw1mHRpUSSfN3KMNFQMqJyT4mW3U
v1KLApC094+VXzBHF2GSNt82gLqR7wJMWycTqUYg09CDSZ2RAjd4rSa3csy5A8vswAwm99pDq3Gt
bU6lnGPQF5G79NJe+ninIdg6VCNG8jNAuxbH6/wJ8uArpMKcCEBBeAqcq+bJeNhlwRDl0O3cBK+2
vNx59qQYa48xa/8fhh6QE0DFrszRv+4tnOwqMAANoE8vj6MnmydGOIByfm5zoiSks6XDEzMZu/C+
dczFvqp2WM/UJ349ceRY/OqzbYYuFdLOqxsY7aOfidt3SViJ7U7VaxnS2d734tz0tA5+iLZG310a
ATcTTdu5p4lA7uAbCMi2reSywy4xUEgmGjnYvdnYO8/dE86q/fV/qh+Y/pV0uAmC8aQ6syCdmPEj
Q7ryjJKFQNrbt0osIGvoMp+nxIkJmyqtO0VxK+dPTsayKgwFY5m0zYUJIIZndYPeHgJfR6OmzEko
im5oVbE+N/UpCFZyiGmDN9+bCoAZw/dpSjaNO3SejLecHgJJqlVCVwX66CWuqf/HjjXDRGo72Iu3
qsPZ1lBloXiYV2sSK6YSvTRLzfaXoX89UHzhzN8tGLGBwz7k5BDKCqNtUPqrOe76Ud3APnew8b2t
dwWYGpo4U8Q+n+c8rYnBUqM6komobB97sonTOMxZukXhhZFb2AbK9soDjigEQJNYVce7LaAG+xhI
yz7QHcyep8Z4euhQ13xiM5gg0rxLg9edbWY7VCSz02E8MR5qLl9GIj+3rVQctr6UXOFrTbp2t5q2
wXb2ZqA5tviE1rdzR1MpKKY8rc80ID8jA5W+tnHQAZVDxnVwoh4tLpoLO1CxNVKq+Ymx73XddJwv
xT6zg8k8agO16gdHhCbB3Tf/OoiGonhfjQiH6Q88AswWJCEGwxAmZODTVVFNAaJcpbZY8NstKgQu
tnhUtRZ5GtmWPEVyvtunPoXeKUKMDbVXw/yKvrrTxC9Y94GJvFTjC+spVVJPoUXIpg6ksyEogxIF
UZL9amXWPD/Nx9WfWV6oes01LrwvyUsB/hgqXZL42iJIBOOhX74LXD0H6Fgfeuwbs+o1DEmrsPiE
CcgvTTSyv99zO8groaggiQAUVxgrHx27wtxO84dV1+dT2sWSQCfifTr6tMLsFafdkmrSPeiAdeSc
K0CeYqrIWMHiBWs/077pDEXCmTZT8uHwaFf4mcHmlnQv+TgzfUkNVbzfs4OTxCxruoU2R/t3FW6N
6onUOPZxveGJgZKSlysfFAs8aIaOo/K1spLigozVFpHkIsJ4CMGf1ZdKhmanj7sHbzUuacD2T4+f
6HBPJFDTPi6BGX5QE4gD4dq3fM3/E7SYEmxHub7DTQPyOzXG62E/q72lyg0jWdqXUQwnPYkqIxBB
MuoCaZDhlzk47O5SYxxt3zdU3VXx1++ovEeM/gXb8Q1prjNKGgnDUMjgeBp/348NvStQ8tqXKsFm
GU0Tbg21XXGdyzQtQtf05rV2Eu1NCyT/3WErQzmPg6zAOUKippxO6RCBqol3v0VwYoGG8VtZYAQ0
LClb1ejO2Vj9k1sm9HleiOnkCAX7KCQ1DiSiwggihm77nx2vuKxUKmaO60MryXus6KwCIm6m01ts
gnyYS0ZTTLGWZhNR1Wlvy7OfkAxaHXy0JYaFiLVLkoHB85RyNvOY6yeAPSiZX83Xu1Rd1pipa2Hr
ciBOna29yY5FC3CWu/S3WQkcfvdLIbuvDvWiFxvnpNOCDhXtNP+QoMlt6olaukuKFIGBlhsChL8u
x8qV0LQb5QXFpF6uWT1PdZoLuNVTyW2uklKT3yBIDguAL3nxvl9xJkGYUF/CD8Rh1NpXPFHUMFF/
Pi4rCPpBQn2Xneds45s/Fw6VtKOxADYb6G1GlpV5lDsazHhOAxAly2SxgFd72LALQ5ykgx3QHIhk
Omko3lyNHeNMs1Rh80b3u6lqBxPBjGs5DLkIhFGHrk8CA0JhvcinEuwNkN2sKm700AaE9ghY3Pb8
4S71pZa0e92yhm1lQe6FAX0acIrBUwHXN/IkSuH3nRIzKYwI6qE+myDq8+Oaa+TFDRYL81IZwuMR
vuUkUQYOuWdusOcseFEFCn3q8udMVvIq1yvqw+blnjgq15h0ixXce45Fq8g39lklqu+AH8gkmpLS
JUlx6fiUEcjCxPqyGUhcFMC3Wp6p484oR8b5XTsPRJi5JFGpNvbfsLoqyX9e3/kUGldntlkCx55s
itjhLCWfOvxduQVw8y1vQGV66RHS9WPamaTFc8hI60SslWPKyDz0fvj9T2OC1nHy0xM+IRdQu5O/
5NcReez9wyy6HVuAB1kmaqz6SP2BgINE8q2tMsen4U5+E8XZwcCAZpfuTsGmekMXBEp8qHm19cF2
ZDPWIn0p9pBwksWz0ePnHqKX3yCayKyXccr6iH5MAuJ9/Ngm+4NsMcO6NIsy//g5Ruvo45AGvQUF
ZACmxWraLgMrLBhbolsFFdnGtILJGoEa9iEjwi68oQPoZaTbtB75CP+PQaRc+Gwjd6LodhAI9He9
ZFTZjLUG4139e4wBT8/NjqQrzdJ0ROWdYmQQanPr7pp1i4p7bhXk94AEo9oJBgj8gjO66xKIhvOu
a69taVa8duI9ZtRy3IF7t7lDgMwD30lABgpgNl/IAUHzhUmtKVbuB+yztjrr4BdKJOwo/J9sWYJ6
2Cuqr6jJy/MjBG5Y2JR2pNW3y+JWEHrC9d2qEzUx+K3DFXE6pn6g96eUbgkaNSVSs+KFdZ3v98oi
cUy9WK9OMNhR3PfaHtfZZAekPLMQAHLyqPhis563Rwrmzuw5x43X4Co6J3ZxfRiG8ADF1RCH60qY
fhuuhxGqiLf11QkBDdSiD2LBIY47GpNbvqheZAxx7l5PY6Q802RAMKRKZTkO88TOYUwUdwkLuxOO
5sKafGdV4ntfbNCDzlzqT06Tm0cDaNUXtsbXEGtHjQXRZ22To+opZi1QKq97uSysxD1xHIm7VT/k
IvU1yGgz5vHlDeb5Ll57L+kXt+nignZymWFAlArMV17U1mDiTSm+51OOFWNMqWIGTcP2SdctsTyl
O5iQ91EaRyIw+PHvzsGRIlKz+AZbnMkyMwFEAjMZG1n6Zlq3I4SH72lXgW6mHLqaBW6e6Mdp/Hvr
nr01c/6pziweoo2vQ0BLsnjEPH/zguYf8uuoNBnD9rVS3MA9w5hxHBCwCLxQdVupDm/DuBnC25sz
uhu3ZJNZosc/m/6pmYzB+ZBhHx6eOJFtT7/NKeB4iKqz25GotE5/o1elcd4H16+fXNbk3Z6cjbFf
Tk02QOEoqbD0o67GZVM8NyCLytvX1Ox7k4byO879vft75W8nr6mFaVNn+R7oXdBOuWVbnObGc28A
70ob/WgU2BC32Vmlhk1W403OgznHG2PUpkJrg2O8d9OH6xkz2rUSRiwSXd6xO41Xjud8rC+ZqvBO
vuQEK+QLy6l4jsKF6yaIi6PCak4VY0zSSeelLU70Q534TyN7s75ZIjkq3PNoA6LRPXTtcNLk8X6p
0/QCOP6GzaJTkkYesAhQGymQZmccrSauSYItLwYSFq+ti2rf1zRp1KMtAGtgHGw+jD3pFRSIVwR8
taALgGesUeeM/RaVarDh1lk49XnO8sOy3jmSjy9qwYPZLBeMmr27MxKYaptKNGtjuJGXiYztJP3P
ush05stfIe168AaUMzOSgY/FOO5cLLk+za0bY3Iptbft+B2Oe8PSZ+InidMm3sclcyb6AivoLfy8
y3ZvhZencfi4hzNZXcDnFY0uD9CexaTX+fmY5MT7hB2HESjV4BH3IGXrtz29oxstW4sXQa0odf/Y
cOOoANtR1yg6Eb11/Ohrd8eSjR3CNDniouoU4wTsjEP/Fct7Ywcba8LydDkOCfK8DwwbBKvt9m+K
f2yLNlmi6+zmxhWXHO5MyTMlVH+uxfv1epHzJPh6dMah+Sm79J6k4WClq0rKOfCUx3mXp1He5ROa
eDOBdM4BKFqxVG8HEW9ErKg5g033PKm9Ja0pllKiTa0zRTfrNDMMVwNeOrK2fp9e+9DVcBtuwtFG
qSDI0jGiiWcKZKYnPiUxFG70z5qaWH9pnB7/mkbmj0RezvexKI4KuHTup5hGmQteRPMTg8IUWKcF
sgOfsvBU70Kpn91hVO9YnmRB3Lh5TnHdW5KdG6U885VkVtMqpVMfxHBpgpDHJjVO6M29zqmfFp+L
jlV/if/xVc82uHsqRUgliPEbWiUKp/DlABxyJipKAniy9ytFDPbyRJZDOfR0hE7i6msIsgpaSIvX
fYUkJ3GzreUgUNMUSEC0pl6R87hG2XnavlGSAuFp6ibPg6LzTqmKBGgSqHv9VaWvZ814S/fb1j45
qnw6JEjbM3ExMg5HDGVBuDXEEen2JHsFjSAJZx87C801JqAWyqPszTHdUfgOD5b756VpONG2+dvW
RuT42hTx7kmtNssaus54VaLCFDvThye2PEICrLdQ3HoPjz+iMKUOs9E0EvnlnfkmWQqs5lVLuHjg
A0NVP20c4VrxUE1J/LeiWJPJkhvnt5i1bObfxzTQ6xvyFNWQMQFvn1nizgKcL1aHy8Zux3mQufSa
kb5ai+TrbT14r3wdouIkc+KTf99S2tVbpXg1dDlxI22rgGSoE8/ug5DxLp4cDoDVBbKnq59xt+Md
4Kg0rtLmYhnI9gQtK6kTdMRF+e7Yckh9LWdkpKr/TMDfIsnraeJATVqhl15o9mAX4dzl6q57yXt3
Av7ARxLg8egMKXWAQop5AfXPfuoRJs2O+hf3VBQdxcd10WF1JlkfFc5k42cpxMLAcI1zVnqp8i/M
hAl1iNaTwrqCk7W98rYNLgVFFOZgjDF+s0Embkh2+t3r+PtIh5IBGHc1hr8MDCaxX/Fx2ThU5VX9
IvghF8gbSIjuXjfGmabIaQ4fCJ5Wx+rDUhok5OL3Pj9Uu9MWNUlcGrgRhpq9PsubSzSCPx5HvZvh
UqY3nCxRaLjBoQk/QJkOc1Nfr/VVoaxPJ/31EWGgxSFBYr4Schdhp2ryTGHOAwkK1graiRBdnBNp
65qyKr9ke/ZoZZNTBBvdHHN4eH2i8gwU1E5J0IfvuRclugHm2X9yPJ6zptZt1qIrHeKKH3scwOan
AY9KpQ48s61vsuU+J9GuHZLECBoR5H4ilr0Vkd7nY4Gwb34kypTNSc40h3f2GCcjO5DK0OyFKWDw
16c3GweuYLfsz7uOaVkNncs9cufQoYg6GYdCjyAV8mts063t3Tap1nfJlob5jcyGW/V0FxHt1dNF
paBo5+uA+NAHBD+QltBO1Mxur5ycgxEmsyfxsCS74zUt/l1mkiEmdND7osdvtippu3ldn1cPn1Di
FvaWGeQXR+vL+yXtyOq7pBJY6JB+ni9uiitaMmZD33Ic3GGro5jY7WVuPNwh1Ckj5mg11HD1+1pU
rfQNMSWotYDswDUoxdvDb0ZDYtIFa+QLZv3QkHIwZQx/AQf49Hl+RXHWe8efCsdnIUAf48kgsOEj
rB2Zv1uJv1iUOCEtVT5daTokqtbG03slsXH8E2WHUVrt28OIJj99f0oimTpJtZdcDYBwTalB9He2
sjmFr5DlbhE7AW2QWhudvdOpfi9GUDWCDVXD58PkACPjvscG0gQPpN9x3pGIC5bHxdMAsvDsJftw
egr4E+s5yBIr/PHjrPz3GgfIo5JChxlokg7mPOohCbWxY1KcBTe7igEj3JbIKxUBxOSkhp5bz3/o
w57LU1f+/tM1jJhboz/DP1xXoF8f7zhcjIZ5kAdgti12ZcJIg6mMa5Vl8EnfP9kR0BcCuVX2D8hS
uWYhIHI9vdmuZkSkyxVY31LJVfZC8E3/iXcvPrJSM9AA5N8TRUN6mUnkxogJC4SFyzK7IHbJnJJG
RQFQxPmwL14GwIVCGNkkgk12HJRZ5sUlWd04Xdyixo4urPnwYPso5grLmPckzrBKxBieZIi9iaJz
H6IHRlllH1aBhrM3ERwQ3lo8KvtLz/N2oEe+0JQHg8iLhWH97o3Lb3Yrdob8M4ISieTrmc+eYkaE
OmWlxqMRbCQsTC+KTZ+ig8fz6cVdMGaKlOErP/huVQNx+yZXLHolEwaNaoV6NOZPnOw//7ER0SzQ
Gdke6iSSOnZGS9fGpYEyAU0a9bEpRdbmKfzALhcleeCpF9YE6YaDlbnIHjNNQmqAV4FRPC1PR1i9
DoV4xaNhNzPnzXIZOoe4ial48/Yr2I6adJlo+jjhkYDEvP6A8f02TYjrLeoWWdmmR1vEKR5C+CbK
aNVo84J0343hhiR2vtylM3Pzh9CP+ddEWt4ZyCh2Yat6sweLxRR9QjvlkIx1MKHxrpl2MffeeBhY
KbemDupvorVgTwzItHl5AyWGyx3mBYK/40XBQ5GS2Q+UHUxWS661nKPcso6A1Xbnq+toSqFSoF2W
Y+0dEyTtFVXnjs6ja4jVs0KjSz/c3xoYJrE99XpVEyvGNcWypb5uGRP4mpakdbggxFOv0YVTLOje
W4FSkS5zvOYtlJaxCi+HFIHkzTiiv7Qvd6RkF7uByuSNGCK5OYriV/thrPOFk/zv+xwovLZJrSBT
jeLmIKdFywr49wpqT8z+90c+azI+6nGOpOYGDOnncH2bgoaQovNXLo96XQ6wncGihJReKFrncRNz
cf3AlZLHw+jIXeTwQ280IBl9shyqLkflSZnlnIGh+BhBe1kZQwDlpCbTnluS7+C/rNdubjeuIllv
Xf8VNP7ttLjio9VUPEQ4HCmBzx5ngHqbP7/HE9LmHQxEuZBt6phQSeH5KpjIhACf+n0GLUS9zJ5S
qWjdtRBvy031K/o6vRHXxF13p78n0yL0YoxYUcScO9fypDbo52bDT66NJPzCBmlkaISTkQzo2J4S
IIPAyXPkDiLah0beok5Kcy9zMMpgtHXku/NPDg/nGpFisvOqZOVNB31O3J5s2IDN+fBnIHbHqktR
TvnfZNoTab1xTzsZBxqWMG+ejNEiqV/mHXMHgKti4rFVK5wdYVM91DAVbR0ViDsuoqFLBW9gbfAf
VJh9LutykcPQMq5u009AKF55KqBMNKR0zy6s+51CUJdOYoAoEOye3TYFwhVklu1JAnzmVacWP9fl
6YFc8IgPZDPUNpylUZIRZ/ngKqqOmaZzQeoVxCz8BFgRtw9lZ4ElDKXwi6vRERpxdKJHgcJ9EJHH
shZvZKCTsDSxkgG8OnvQibTwo9o8LCdPuFCznGu5pzl0PLvVeWvmj80Tw5Y+Wms27RfVZs4naXdw
GCDyfMe+5Zn2ota+4DrxZEkKrdIc/OKRCeKgtb6m/WJ307uQLVNXWXSSAG/Y9gr8utgEwn76/cGD
hM9CAre4FrFvOMTA2vG1uWk3OTz7E+iqDgsXdPPS2hfbU48Qvunblc5N2XYWHhUaoxM8dxqt0O6P
82gtesq2RSKwjzqqACXbfSsktQr3VBpCaKwJjS/g+4BzyMARn7MPjITO+mm6XuVQMrMrn3FybU6l
fQXaeBOfNkQNgwcituAkRj5c4VqAG9XbVNj+OSHcDVEfk7Bb2WuoSXxk4jX2TpFld3GNHtvPI0LE
DTvEjkDe4VCEMTEM8DkZl+RlAjbKUmscVbKGdrpofMmIVeGyMM291A4xRR2npe7qAgrKLS9+vz7W
pqUi9Q/MV2j5kTLoVIHRnw0hvCiXn+HFMFIU7ewBr3EI8mbnqCJ9MPqj4eRYLCHssGmEFxcd01lK
pSlfnjkz+zjMzy6wSEZ4xAb2QgrUc3pG3akU9X/Bp0yFQE4WTNDhbt7qyzYTQDZ9VHMT3/9MAvTy
kpRvG4c5gz9S2CJZ6hSwEUm8f/osHzfhpBQXorVmB2JaWbnA+R55N+31tpOIAY0XjN3wkni2AVWE
4gaOY3FOu7c2VmH3QFu3lCD+GqGF+2HDAMeiqghEvn+LIGs/ABEEpKeeXGDq306NVSefU+7RzAsu
R+p32fCVxEocGOCfLCLLaRxxnh/qvKqkg1JEI6t2EQcVBLEFC+a9UOJfRwsEsxPdG6Eq3tDXlNdI
+KDZHdQf7dPifDE7DBLKpQzUsOKeczkPVirShULLdwbE+uslT6FW1SutFsLCA+9c9mnq5xCt57/6
EWXkANHBnXzfHkGrV+JkyF49o0aXTpcp+JC65GdUOc1EAU/wWYOZP1BXh0q6mrjiGe2lnPhQbBUN
hhyF1gWsW9CiuxXXeCd22WmG5rlliWuRSlsC9TTcVVb5RtYTR8ZvzSF4j2LhR4zq+N7uKDS0df7p
8q2fLCx9BpaPkqwptJRvsviLIl5ZkOkNJkI4CTNZit4NlrNZL+Hxet30proyY1fTMb/KKTg+QpUo
AQ5ol+1UY+xm4L8p6Feq/yhYB6vHk/+wlugpTJM3VwnEUPG49fIgQ8LK4dp309VHoPbQk2HXsg9n
j/XsvrFKO4W0pOlWmSVHcmjcFfqpJfxUxQGI3WZxmeLkRxflkFUguJU4vhrCQCj92ZnCDRiYZUCQ
ps46QrT+mz2aYIK/yb4+nzwaXD4QC4wmrOMw8Bi8MpPw+8j9Vmj88zYgZ6Beq3okOtZV4YCy0bJ4
nJEB+m2gSdT8TdCyHQrjPKZbZZRrv8bUjtwPYFgYZRdxosPUeJ8a9Z47fp08wKODxj5rOwuZPi69
jSsUIUPVq80dy8ukHO5B00z29ikbaF4kLzF/zZrME13bQxO2x7BKGmSbGpR/HGDDexBeeTwVWrkq
40AMQlzj1HhVMFON8jF5fS9Ghx0CJFpof2ftwWY9Q224emJVe2j7ohZp4pjN442P/7uDQ8i3nLMa
l7jFbCfmjyyT/WE1sjzbIXKhSdckwkNrmJBVRO1c7W71GP9b4CXQHNna8WYdReP8ViG0X2a1e1Vc
047v1UggqfctPNwo3N5xPsKI4EJxzZFqcOBhwjcGjByQRsKs6uwDDC5N7GZj3sdEf8wdlc1pjyMJ
P5B52yXJGYXsINY94XDfDm8A9ET5fOf41bh4uuSJAlCcn5gnbPLfYajSIKAaLt7yM/TX5wxUH7nm
R2RmzwYZbM1YdLhSAtXEDccmXzB06Bdn1qMUwKDT++A8F8YHOhQPDV3yVPOxWGcwzVJOwTNNucxR
W7pFZn5Elp4DcRM6/bPGE18dShq3QMqzDM5hpXGHsygioYcn+BTadQ9ILGZNaj3kIMsDRMhVwOFz
Oax4sJrAtIFZs14UWcWt1DcqdskkuC+un66qQg1yby0RBOCwGry+YU09ZgT1sn87rypTeYWefhNK
BJpzVzTAjjvm3bu7UdMd2y0K2kj7SsmTSwPbHRCJOxON91qIwGutbLwWd6Ch5ksyM7DVJK8oSFtg
JnX2BVaSagdX8yj7YF/Pzs2l1/MUnXUzT2Ak6z6cGOFu3Ql1E41xq+6wvPqu/rkahA7bIQUrO4ks
NfxxGgxcsynECC+KC2JHM2pl4jY7OSEsF/THsY4LMudelmzRpBHG/cTPQafMA9xZtsxgS0EtEiIR
flvEbXOxwr+mSmhF4omSgyLJpUaYCaYS9XjUdeR7gUqkU6mgDfkji15BjxcxGqrpf9fWCD/HRv9w
bGsRcRsrLZTnpKZt7oQjqPgTNHkOzA2VoSUO0jHXtsOt7BUSPKMRYQNaaD6p6YpJQEm/n3+kBuqs
CwDyFvtK2eZ07Zz4mrex3HJVM635DxlqnxFAEifyk1BGktHHtKE2/APPwyuCENXCKw6W0oMXeMYp
LnbBThGF9HX6hAeimbVcWCv48PnnU+UO4djm0QSivUI1OtOCNolUKF6Sj5QPoXY37ZXeZt1UMfFa
bKqo8hQY4/8axn8NvrZ7nc5QOkgOAIccgd+2aSEphhViG42jToiCpjE4bWqm72EveeUtJ7E1qUnf
n6E5ZjpbJJ8KI2/X8dkNGKEv4ZHj6NAE2axH8HRWynGk1XkYb/S0vt1QDH934qsHhFg5skx+ETZt
bCxWEIAXmvAU2stSqTFgcfk2G7/OIjWSEI6G8xOAMgGoHM9ZArDck4ggfDw0eVQ1EwMPZB0KLXPZ
6sDseFNDxSFmMjavFrDhSnrmOJ5XN+0wdCtni34+hbNd4hMBwQEIclS91Wju8CSCd1IHuLM1jtda
hx6UrvoWfhi/JmEmbCTH+SWEM4Vof+5mzOFO9EwYjrtuu0uEWzrfjRDUx31mboFo0nAgdCOqWHXk
hJfren4MqMjq4Bp/5kfjPigDu83br6WPX7ztWd5NqVw+sCw8Rbb5p0Y0U6ociCBmb1wj54aD9zSi
m738OmUSb3zlS1Sy8f8ZISMPzxeRKux/PoxJv3cNrdTaI93cPqnikydz9JpT7jt718aoPhvoMN32
GsBhEGZ5yZAdYwE2I6z2g7OOkJLVHUIY9yKXEFucRX152026rJ3+STuyNFW733k2NKKkFOPpcfWA
pf/lJNeV8njwOheVn5x2jJvIN5oNhUrI3nUEdUwq1sZjolKC1Dt311Gui/eFFGckZIvVXGQSsmWb
EnxyKxOV+xXJqWDVrgm5Nm22AAsK3OJVehIQFRIqne995rc0AWj9ikHW5rG0ZBxAkMjM6nDEV0oS
FX0GjrcXFDJfCItEogko+jENb1xShfr4rjYjBFhrG9BwK/lzTLwDMFabp/BuAcOKGJa9Uff5HMTP
+kap4ECzgi0oLD+8rwRfu1wwqZJPBzRFhTe01RO1pNaaPKIhMbT0JFt8NZQHZl02Vr/rihxNHt5T
U4d0VLyLAdGia5hbCxwRa2JBjKTkle4weLKx60mrrHnb8oap+dBgSixM5Z8TS27TzxtgjiC/jw0C
eS3Im/rLMsnJ0RuLIO7N616DIRzCsWT5oe/GY1THbopxeiO7Hh2sr1vpO++oGvlIvoZHftIRrNxn
JtH6aFz3/sFl2lcmtVOmKgX6epseqm3jGm1dMOGZhJKazbRI6QsK65AmZoZxtokMIRAHGeXtxasW
2TqmuRowXOvG7rEabW9UPKfJw1zBk9L2E1ZAKv1fl1OOX4VH6vTxXZQaYhsixcrwlNWgpJKHcgep
Uno++wjQaHXlXsAfkXJAqq0Ljc5JBYa6MHCjpeIxI/YlSws2fasSr0f9PA0bqGlgwpuiDgtdjqAi
foy7jjlmbcsx9E+4e9LjozEWCKgVwvfy/cUS9S6+3a0udHWF2UMPb/ChlOPM2ekm4lmwEYT2MhAw
PoHSKsGfEcrHmDRCw/P3MzYQtq+mSROWw+zzoPqvZ7qhFzZOic/oUu4XCU/ivzFyvsgYYu+zpXzV
1Z7xG6v8kMtB+Ujb0wuP2pUOC2sQvVtPKfrz2+xZuz0Vue1a18hO4udCNtHCZt7/WnKh47gYX/wR
4NnNMUpKSbQzOy9c4ePckWXsl4tf+vtacYC+p/YO2sKgYAwPuEVATR4URVVp8ujudhMiOnbxGnKK
pRsvo5l8QgJOUVYxPQfC++UdG3cGSHoRXPTenFwZ9tEQwtVLSi5+nSBQVyaPnkdKAtZDnvGeDBSt
1oZwl//FQeDDTQKBjhmkKcDPPOHiXJR8VCArcf0SRICrbkTQ4CjkUaR44PYjwxZphwSGsBb0QkBn
cm0beEGAP41XDV80qKf8GHnHtmd5X+3f0wIvhy7hpXumAaa+F6RVnd7ESbBdTD3/Qiwe6MOlFBq7
/YDJ2d/sHDcZwDz+dp7v0Fn3r7hMvAUo5iF7D3fdRgicHwK1jgU+VHxSUd2+05cQtaHAfWGyyzwF
NdUla4ZoOcyXAf1IV+OqrKcJTAzSfn9CdnrRe2ne4750sywZxLJXthubUejr8M43EbL8guRPt/oZ
P6omswhOPOgIRPl8SrBndOY2gPQSkRIIrnD4J/y5xbqp/Dz/L6nXP58JrAM0Y/dsuGwnu0q2NyGW
9jPhTj80MIHzO4cWVTsLy1p8S1Kyo1D1jGh9mD46EHk1aLFZI23RajnS2MahzLa4Adq1FuGI99Ge
Gcz/JeMj1V/4G/VlOb1W848NC7/k0/k788/QksdZsWIkTekvgHQsDBUdhOoMbKP8SDhhNSavl2CW
E0f9uxJVBoCLpcjA63zmy+L2mPDizCHregw4sbijgjdexVzRNzXLL9+xIxOwb2P/upez3qc/B7Jn
s4k2XVr/IP8aACOsYyorJFhHC8W7VJZIwaQcCSx9zqRDAFgCGsNLK/fOjwSk8dojcn+COHjlnzNO
raPhP42iHenlOLDvFKsFg3x4nP4+va3+w3Hahn9y25VQHiv8/6f+7suTRR5KJCcqzzokd8iSMvgi
q3U/OP8zZzs/49h0y+NHt8GZ6ixIzt94EZOLWSwos6K2W+0neKnmJtHsovJY7Txf3DscKgqSc7tZ
0ESIuxKq0/EUU2o6km52hjAvg7V7752Ap5XBdEgI4Fpk6LL84kp53ocJnsWM2P/pv27CW2Le8m1z
dkHJsDoxCzzZ5bYDjYZIXdFYaOwxiYdbAvA6XwNJgoOvZlsMM6DrXo8Xpa8Nue5ITBLB7URqj0Q4
AUnrTVLPSHfPYG60nvXD3ZT8k3YPpIIxq2Ds2XVUKoimQpSK/MBJC7bcbxqOK3YNXZETv8jtf+w/
csYyTjUGDjunGup64Zy9ltNzgtCQ6g/2QyBw6tM1GxI7czX3ELkHtP9wYcy6wEx7W+CYd+7pVvlE
ouk1uzYkRaxY1x0q2ej+fXPawEHyvRwhRaDfD6j+xonK/3HufHu2DH3p99jrba/ULqPZkHPfeNZg
6dQPUdNSA69I1WE8hLSzx6stkUOC63ItH77pkX4Jnr4+a3gdJ2f6706+SKNkIGDTQH3KlpSY4fv7
JW5SY6kZRqLucO68z3qIfnmd/C53f3AZqVBOxuGir/qkB10SRb8FD2dmsmLsRchlGzr4MecD/e0f
w2r6UkMQzVOsG16uzY4zw+p+0NEZLaCZL5rLbDbeWfZlQGCmXFniUqacJyngBPI6o3KICO5L/fdO
nvXmR7M/MniLYz9jUfAh5Fa5ipEu1uMlLpY+emLMTfnjCGWRr4CqEhUWwQoYYmHCtvdR1oVlJUiF
AelmRbZYhtY89B2YllpvScrSFqR0A6EYdYtbA9FwJAF5SnoKBG3g7H2CsAncqc2BWc095l6BNHv0
VJT4LDBeAa7PEkgb89ufbbqW1PxxzTIeScIZqP2UwghY0K6AtzcXsLFj5mthcXO1O5X4Pheuk3J+
r2PbyAonHUXHowkWbFf2FyV68Vw5eLbxGkE9NttAZkSK1AY8h6rqY9saUVciDpoNUgs/bPRLRN/g
2DgPd549irWJKa9L0RyW35oGPnf9PYDllORigBJs9+/RuJ/1hfLp2DJSoIaREjtcVrliG2eUvs0X
ok5JFirQmOki0XdW1si1tycAQsdstPfuEoLioIcAUxtvhaKa+RvnhN/VHzdue2kNWnhrsCyn+FWC
DAWHAmlvn7kM2WW1HZgR7qjn0lCC5inTKeNgFFOaLFcoP5Ghjycscj5hy0EqgxcrozqP7pYowg2u
xEyf+sdk8xN8see2hGqdednyEiuw5gJ+j+r8q0kVFIFMKsctb8CdI8A6lVDME4R8ewX7rJF7mRlt
8kzmRx71M5ZADZTZDm1E2EWyIJ4FtIgOBaAvMjVy0/YRJBo6NBZOWB6CO2lxxbLfUruzzdE25Jcj
H7CTZFZncn41tCZROnBoCLl6lQaLhpJalYT4mf0bH0rLWXz5cVZHcLlKNr2iEU+oCu3kQYMu/iVA
k0tPu8C0miT5RAmOyBPMx2Xxmgj4yyQZoaz0NywaLmAnSrqMzTIpjh9KnTvtUIA9d3YkRFoQCILL
7nFoAFrgLDmMCzi5q3shJ3W0cmUiPlAeQqH08DYfSqtKQQtJdG+AjeO4axa/aOYSvv+mSTbytquZ
eFgX1ISbDj/EYLC4cTclE/1Pup+QZcpqrnJam4ZCVxeQUGP5vskuR802mI9uWRaori/T4/qHxPOZ
9BvfROGVqcjoJWhzMdtiCK5awxRcihmVPXq+4mygGph4YUGVO5v2O4dazb4FC5Vf3eFS2MWdIWnD
hU5/ITS23WLNu4wCZ2yolz+Ak7MeGIZF60MW2nEKHkf1klRMBcaxsLgUOE+4DAoXkioc8J5eZKOR
FE9ub4z+Wq/4lTPFOgOZj0W42/PEVc2UvFw/a34YD8w42PWM78yDQp5W/xHc9SbWua8h/aokrATl
EXmANctWYDuh+ZkhrhRUnqojhKjNnjQWmx8zctUT4vBk2mNDmgyhriWlLzYU74kFRpjQxwGPZ8+E
63YkHeQ9u5hnew7oUzHKSRvHWaXhmClvS8ibrWATBkuE9uoOddrhsfo8NDozyjj8+McPF+3DyX2C
rn5+3TvlfcEJURR7SNiGvmmv3vzY32f9hcMGcdHZ2vZZavWRI4iKiZNl+fK6Xl7r42JwQ7sGGXBA
ch7MZVn0Kns92N/58oy7l38HWSxrBLdPncPNOfcAP+tVZmPXk02iKdUaDcaGJRoRK+IQQmLRmIOf
dOO0+yZCk7ccEpacKQobl4m3swjeeyVw2zWjoiXwD7gvbhuMae1ZPsNOe/yi5xOZq3QfwIzEGw4+
aX24iPXNIvf16jOCg5y6kZe6+zqLIFNjYtciJy+G0hxAUHAMCRQUjYLeJODGl/9nbHVEKVbgx+Fu
yoTHE6i17uxFUQm9uFn5jkHSljpn5YuqIMhgs846kCCApVQ8BeUV9mnICAxjqySuEyLgRxgJqaw6
2dAuLAWMVNBz1aHNlWbhxJorNbD5EYfa/eizDosjIW3rYivgI1tQ5klL+IRao2LhYZK7OJ8nSTbr
8SF2elg6MQ6FA/9R6jNf3MEHgMeaqYn4kqj0pQZPDHeIQ1mcU9JqIqDop5Ee2tZaz7Jmu5dZDUAj
jHZOtnn/ymWdDsrDQW6FHM7ARy+cyYLOek1UjE2i6wjSrIe/1rvWeu0HMez4VIqzLeTf4psahPCg
3wYE7POVXkeD7A20xBGk9UEmanK/GoFtbVFQlu13NLVIjVfGFycrDMQN+czrf2NbQ7qZWE1Fi5jg
voHG2EDvIt1pn7akiuEOEep97FG48s40tmM8hkWqf3QbrW7YH8D/z4c2i5JeArI+xm9lnq86L3HL
Ep/yPRg0VbJRyYcZOyRy9AlS1w3nYdi6z664D7DrEKzGe/PI8Srk0E3PApsr3EAUx9UtKvAhD9eY
WftXgc1vGLEDAWXdvdbZVIb397Jg6Qf3rPyF/egWkPN4Chp38TE9fgTHu2/q7jJEHZAv8zbkgP6d
/oaXlmPv3Dnpa669S2BoNTOyaiScn1SpK9rY1x9hvqFmaQTjEZ/Ks+RxVxz/KwWv/StCspyp/Z/4
rziE9m6CxqDUaVqtS1dl7WqkDprxb6oGswWxqeJq2qCPBQzbouBOMzyk5N5thTJJVNFg3vsE2h8F
vRTmLkXxDqwB5dk3Agoa3V2kvnQ3JQhg9XAY5cg9pZbVAm03jRhKSw6OtJKs8P0cFykQDOBHQOWy
53uq21dMbWD3EkSHBuEuebcN3B5JyB75HF61Ug5gJwjcoAFCsHRv7m9uciQU+gW21CkfYUEjTMxr
p7AoCS5LHMoaA5pWVrp7aLffz9wo8xxeLdrmxZ9RLx0QBfctTbFvw2ZAl3GSJnDHgc0rxT+fDdzh
lm5vZZRuI9Za2bwmIPHh3TynK7zX18KRnZSxcsbtz9krJ7lZWsRVqy+VSw0VxNdywe8AU9jcmg4b
3ceI2d1v0sdVmGnEvjWzjdizCd0IMvc2FbUsImO6yZt2qUhLzFoPGpP2bXc3btXFb+VhWXbEFgZN
8cdSgYqVzlaqrOz00IeDN8dqv6ckltl77Hbs6ulgd61mPiMAapmcTp4gEn63zAx5yXxlG6i7wtgy
ptI4TL+iBpoDK3LAS589SwLrhRi1y72vbPgTWvAdGJIKPsnXfLJfYEVZely0jETTok26VJhbahUq
gRP2TY/tuwwCLt+h2F17FOfqmXw5ux1erdiI0G8HDyolcwAtbev0Mlqbtrlzy+Y6QiM9m5WrFigA
wWa7qdhsfzcie4Pmpbnt1Xc1FRWxd6kvHfdd1TX8/NTP6K6o8NG1EQ3Z+0BEkXX3VG4TWB+6qfCk
Nhv8zWeGCE5C/D17xbV6rDoZTRgK7OmmLODFEWYWr8QXFBym/E/TQS3QkhDwb9Me39AxGtf5lnrC
c2g5zCIStVTqaw7+UHZVsg7+h0BmLsw4ki5Bo/ziu08IILz7XUoUeJAkXA9/92iuup74vwghzoau
K52giS+mo6lXvknKE9YKJyQehCYPPb6hyl4/KrECwF5m/lGy7myzL7SYpXUzhv9t5VT8RCokWaVu
8kANcazvG54DuEqyyn7T+CrcLnMjZmr1n7Eg2GoIbvVT40sBGJPGp39AEWXFeJEZR32RI4R0FpbB
W0yWGFDKpiDfLZBxvEeAwu0wRdE9ppXJv6csyK7gCdliqlIgSVP46SmyDyZoiixgbm8AUfa2axKO
V9hhJvsbX5XbPWnf+MdrUJOazOIeDYwJUIXA5ws+wnADbIS3sB84KhPRSsFENYVKysDquXZi+YD3
OKKr1ttnZelDNh1PA2Z9U2TcfTMZUbGhYnFXxEPo9ZuN3ha+vXFI5pe/qKOp/eGWcUforyn/lFhi
SVmBKGannplqSdTb25cHYKWRV4vrXJNAGJgITGurY83i7ya5NC6YqvNn1wgyN8ISAFCM4IA2l7cU
G8biFHSq2VzJ1doqhLmZu3v9r2Jf4uukxby0griokdwBfa9t9n4vKz2+XafNRA6k0naj9UQoBVvK
2qkJiBbpCEF3GNP3uJORhg7qZRdBEKGRrolkBXyoaKZfCmBzvAxOku1WKBPB8AuoXjN4pbA1ns7w
1VTfsu7V2YMQOekMbwz4rhSlmo25kaHB28N/Df8/2jB5jxCDoR8/dy1aCeMoL/VngUxk3OSCzeb0
Sqi0zTmezCoZDPPFk2kaWI0B2Ts+jPUpHufhqV+8giRGiRarts6Xu6mm3qPP/7NZ0G3Pf0FwdyYV
OM+xNCjJNuNrSUKJe6WeloT0BsBNIKOOl6EzoHLjYCnAjO/A307BHtekdeR4DK0HikeBqIoIKSwk
UGN30a8Z2MptoPltpOB3v5fn41UzTycbGOeC5USKud/8dlJHqxJNG14dG7jkgCNLunkE3Z8km1/a
7oDoF4DSZDyl31CLYIGU5ecdojRpz2bLs4nRITJYmlY0haMuXqzF99SHto2/gDHNbhn6xh+dIjM8
dykg0ConCy60f6f/VWbzG5Bkv0l/EmWK7cC2ZCh/un+FgBxAH6x7ePHFXlAtxLbWNJ86JoTGwBVF
SD73ONCfKTsKITQX7b/7IvW5+DKoGExjP5UPEiuE22MODBz0i+gtWXKve9v0TmgwljBCY/x9oghA
DN6BjjU28krXF+lI/cE8z0aMk+GzKRAMzHu0KCQh44XMgHUOQOkAa3RrAWMSsLozS6r8IfxqlPOI
+ddHmDFlz6l7yzvpEzdrwHP8F9nk1vo87Vgbcxgm+GfPgAEhJWMg59AnQqfBkWdynRu1K8YWHHub
kh3Azkh7nOvndzUNKc4JD5O3OgsJAxgWeMQ0dPJbGlyJmY6kgtQTzGWOedTyAbldagA5xLQT/pkq
o59r3PomUxCaIoO1XuQdZd88Yzoxf6cp3EMZgmQH+eyrrUuT0QzAn/LavrhzeQ+78ZI7r/dIFFXE
tnB/oeGKRhiaYWO5TZ2wUU/77rD5CKvJDjaMvYHHo5/7dA9c+8gIV0YLk2KM6mzs0wKMOJAG+A7d
uYt74NyGNlOT0/V5URtMKfokHbTPpb3nVM91yw6fSXFqZE/wI7p/RUeDwrhg/bzcYi55rAQHpZcr
c6IUTHOHJp8B9ez6lAVJ3cqAmIW1yJ34apjoHI/BFpID5Vx22nJhHN0kOCpZHrcMjqf8+fn1JFoP
374NuqPq7U3wGGIqORpTqsnH4FXGqqpKIqWMDxvNwWXsqqTvFByvuOWhzU7+9sI284G9oN0dTp1O
HhW2qBXCoOh2vmvyeXItglB4p2xcn/21Fx0QVhqs8QeI0+K3Hq+9oIdoOmMnwenNntxLJallaUuC
VqOcCyhWKbretf6V9InPrxSgy2E8dcRQ1oP88BHR0DEZF20m92ko1AXten08fUwySFB9i4DAQr+Q
03FmHcfEOOoSrUzdNa3QQgkWyU5g0a5OjUs5qEAaB04HjoV1EVSYZCO6QnN/FpujVU3CjvOLtthZ
UHPEQ4tx32hjeitlycv5d/ACnWGQ0WSAu/3QO8csu58TiZ0Y3IJW9maVxlsnq8AE3KRxXT+aDtEu
xU1G/zAqV41GAGI7ElBg5gcPV3PmoTBhS+rxROdogdCkGju2i7iV3LitjAF3L5ly3YeBD9kNHwBr
HNeup3aO3wPYarNRYL539VPPF4MjurlaNrmxE+no0CYAO6ILRYn70uxfrBDH/kBP0T3eNRgcCtrh
sCq4ku6MmzaGRIbtJb/6uRc0D2DOJ/1h0PRpgI0Ch+L45Ve3tqG7+cepS3KmUqIwxzqrM1iBHHw6
8/KFHEQDvputmKt90aW/O73WXGCDkJ9WbqBWXA6od61HntINYVd0HDzIkqd/2N53b3yUolvAsJGF
KFhfE4w0Q5TBNwAMtcG17Xhh5nDgdpTdJgTVu3ErA7uoW392coXzkfkUYzeDSLDfg7E6eWokL7LP
c+PnjsR6Bxx7MP2C3des+iXApNEj8HieOO1C+lwYYL1C/f+a+4J6oLLnCHAwUHQxAERRgLJdkUrf
R5jXZyuE3eWFKNJ8/XZaB7t14rewW8P3GBRhyVsJjgfb7ZdCKrkxxxN96SdARu7S1+JIuOVe7Zjk
gOtfMiD+Czs5SUonjGpvnl4x0llLWEHR173Ln1KHK8KDi3+kzvXevQ0UXQldG5wPAf7fJaf3siNZ
1nh61sDkG/yZTIDXdLBrEi2QQ+KND5U2PKtkUaOphzpBhlaCwjuNIUtf9VnH3Ua0pveQlFZUkJhA
JlPe+FjLoUPfycpRE8oPyt/IB8ey+gnxY6psoWiIWY6w78QaxqoK1F3n4nLuDFhYManGIp3tMh0e
ZZp6iKVDbRgVDguItRI/hhOaqQP5ZU4fpquR0R/sOtrUwsMkciz9rkKcgYWzylI1j9WSKMKPAh/Y
UB7e6FoYojM1XnHC85Nm9ng+z/sHXSjFiffrtvbszaKf28v9KBkis2TbWm8Q0ko3BxyEvO+Cv2Tn
zs6FMDsbe5n6Osy6WICfduVhRAZbft8ewT1zHC3tF4+qWpUQaDsTve5nH12JPry9I993w3kxqs2u
TmIz+EndKdOQNUMbvBnnGxwm8nJSIpXzotLbyab1CViCKyr9cKxsxZ6PxpT6eLh+QOTgUowzFsiB
/iZdvTq5hcxOdKwpnhA0kJc+6AsyRkbHpwNcUxUDKQnDknkiTKK4ewRGmaJW+SWIh1ocwHcPf5e4
pZcBQxv1gEVD4gfvvaN+GgcCEjiOnuPYqlpIb63XKTfWNToriuP0p4m9ZzxtUDgPmyYrfgr6d3hh
o1mCk65LPq3YuDMCSRKjjkr6BYfIA0G0I3Le5tSKBU4gcOxT7Bh/UMir94Xcqh7ypImWvV+FtZVP
h5nKQLlH6zT6z0rkQRMqhNka28hHxaQIiy1TVlYFd30HYB0XCHpeHVevkxBvkUAXwimxk+1018Pi
koDJdpyhLVWIXD/YgAQBwS4UY0wQn+jBLKtViTUJUOx37UR9hZntKacz45j/eVgOhOnCCr2/I3uh
1educKikiZPusTR+B64dKieqLHNNG5kSGW2JXzzJWvFpLz9jMKtHybaRHD/dbX+hEjBTNV0CqKKb
zXT834b3wasm9yBUz5RBFtq5oXeS720LHpVx/VB21g7585m0zEbyMtx7B1rgjemajGPbpg3Wt9ZT
Dz36Bi9CbL/e9uKa9xriX/GBpcVjACOLvgo3WpFz1niW/3AK0t+oM/3dGN1CdZtxy3QB+qTqC6Xe
qKYWK+YDynpOgY3HupwfXardlTDDOOdzyPB+zEoNdxcSPvLSkWSVBHCHe72rsWvwQDjVezUS1dt8
x9TY2PrVRKQzUa+nhhIp5PK9tnZbfFQKyq7bKJtaQTjf6GBfBTLxqjqTyl3iF2/n4A8v7kXTUJni
fTiXpd29p7aRmJPj4BG55Gl+92LL621syo8ht3TaPncneS7p+knF7BYN0YFzCh7nAoeEYNZ+iUm5
wzD+S7tMa+q/35RMd3VJOS1VJj+LmrCViqSqjntU4bszv1V3uT6LVxkSqudBLEejOIGgmhGnRVTQ
jzauUuPDssM86Idy1eVQU+Tbqb7TzTyNzbnyzRCEbH0Nm+VQKI+FiUGnH03gjXiajWQOZvzl9ef0
zBI943oTHlsQrJiCA28yJ/SNH2YF6QPHmsUt1FYKnBbeGi4DAtRJAzPt5ZDL9gnP/KRcpzI13Dx8
gh5YB+ZeMBdEpi0YAJs6QLpcqgJ39Yu6Totj4bad4irEE6yL4w0uq86rQGoSLj+jmJYCJhbYwQPy
203M3AHekJLZ2EQ31jw0Ha6dxLWF4wczPWGXhDyQYjnxF4bS/FfTr7p2DbMW1D/13oO1VzKb9Dqw
Tc5lxEve4IIapkMRGBoYiFb4Y/mrFGU1+/vp4YTwRpuxQ6Bdh/kvg/0Qc5eXzPn17IilF48XXqmH
SdA/6DmqMUhnw5kcFbWZCPZ0xkbkjPqH2ucgpACN9aY9MkG04UC1w3jiHHIdVTIDOBtLOZz/uwS2
E8r+yqWl+IuZEhCJj4hayiLbUCPMzTBhqYdbvYugh3qxupknXLwB5QN0AMhp3dAfdi/TfF1C8WVR
T+fDeJLVeyp82MQPDnyZ5xoNfTpcH/nby6Ix5uUCrDBmqX3U/FPe80sg5Qmw2l5/t3IL0Z3Lv9kI
1y9jWHjItTz6NQHIneK3c0rqUxU1123q4zl3bVLdW3XhFxMhaKgwpZelXIZARZ06SZ3koDxSNIYe
ZnhjuRXJFqexO9tHJo8+j6Q4XPmLftGH9KFvBthibEql+xAKWQXVQCJpCbsj58aebEjufJJC8Yes
BMgMtR37kq0Vtqx4+s7FogwYrbODJ2PFqHQU8ET1yQgJuwXh4UJb4Qp0WXnc8ZpMeB2Z47FeLqFu
R2Ri25jYZieh2md/uFeyjPGBXnZIvz3D7RUAanjBES10cUsdcILr2eeqbsvgwMx6ooP7QBAG8LtL
S9ntJTxvT+5DH6ZotVryw9z61bWMJZLLNofONrIZF91TELrVANEA+cyzxvSqDcArpAZOhvZdbxkG
09+ujn76dbcxMgrcPgzWrs2ck4pqkm+Y67dJYlVkROd5nRS0+B6JzlpNEJob6bNhyGLMwQ0SigKC
vz8zX3ud26A+FoZpk+D4dzykGhYuaxkjj2mCFeWRG6DM2Ism9kackGcqJyHQQKcenG7Yjg0QPSYk
y6YrYpU8Hi9x3I6H5zgHJCtYJe2EoAXc++/YN8SGgz4CDoDgVxsncImVKxuyQCoyv4EK3mEwztrc
dD6b/FGu9o5SyCQl/uff6B4i4PzIz27IpqL03N8E47xtNApwA8Xc6gE7FuE7PckyJR3rKLH/HtsG
lD+67z6UtK8B5/XVfbv1quOF4XwL0sCWJD59ZJXcd6SsBtw0TjewdibX+UQIPnKWzROtczffPH3B
fyTYQiZm7uJIfMSAhsSt6tMx+Y0Wg3FDoMO4gUaPbRTmNCvP+TBkgMN6xVhB8GxrQnzPbjtaQnfv
7iapbFrAVY0fjDQLN0oEsCR9Mrk5InG+AaZ6ZzKiXSNSynHoaEckTO1dWflab42yV5eU4mfl4Agl
HD7Y1ZlFZ+gWvohs5ZPhQqHyrP1BDysJ1tZBn79KQOZRSxDEclend1YUtcS7NYC4pG+tCbJzXjNr
fmP7t0OSJTSWe1lPezJbZmiEEy2Jt6R6qpw439EdJ+KuNStocvLyJ07zkchXtGlsaj+DDKQcOU4J
2gs5gQL7sMrWY7mEPBFJvmbLhCPPEJp25WLBJX5iifluc4a/GD26pltZkOyNZQzdxhTc5HHGQrIc
BwcDac878ut+SNTOtOuLdzKvvXJg6WuBv+v99UL6SxwGEEBxgR/uiH81jFgAwEFAMerfkQkODcB7
SAcAhjKg1xgkUIWJJ/Cr0MjwiKqZwnzQEyU35hTyizkQpZMipEshFN2uS0dgsMKZ7R+9IOQjZaDv
TXUxcVttGWzvCZcGTrBp6xNEAh7I7j7rW8OfXzCx7gY/HXcarlaVRHJ/ZHalhqRue7ljQmVuYFbe
xNMCtWfR4Jhdzk2oE8Q7nboVUOCH34lWYXFX1IZhd39SduSf8vhB/HwciL7leOizRbLSYE370Kjs
WTzWi4cMWY7y9vTHjkpYndVANy7ET4MOyAf/5OzhuNRuxx8nqcHhCgSl11jzLRj+8vco/Z6R5lrh
RaxOEBW6uuatLv/2ezHEtPoZonIKkaDXh9K5zYGqtqtqat05yZGA6g3sapiP90WPGVJMXu3xalmV
HEjiV9Ca3AK0u+6idPGl0EuuUDgP3KhU2GLZo81r4w5chnaKS4myof/KG3uHJlfmQQ90XwEBwfkA
SpMbyE6m59C1ypyPAOMy9hUKEJMLllT6vNIpiZ/R0lI4yW9C/fo9ZZHYpaUHRceakApYYkr+xMDK
yvvt15T7sE9NxMxXoCLlkt0h9LQ65mWjdBUNHpBD0xsFuLCRqQCZ1OjVzpnkLMCI9uNNT97iqO2i
kXMBnuO+Y/2i/eD4IeVHd2EYe5ybWwHGfw4aWjaldhiWhWDqMMHyp0VTXuQTN9+fo1Wp09062Chh
+kR3llsC6tiooKno7OMmNE76uLDftJp9zmRCMmUop0JEdezvtnbCyJ5WrIQTxqP5VTCK/+r0IiTf
SkytAYrA+ehh6Snn5oyTuZuN41hGS1Z2WfIXivQY+um7Ozw3KnxXJirqtUqtLQySE1UuOgPq+ZVN
eFykg2PDFBuPUQF9UOy69dP0QBYBpyjCrhEd4brDiSuJyUB0rbxCcQNG/pSVm9Q/95ZGAsLiMsKA
5VoMZgpExyunD9sSq0mM4UapQTrz3ptLB22kam5Q5hdcBDbn4yTrN94if/JoDWFqs3dxstLmYP7V
nYHa/iy+CE94eJcS+UnV7DtruKhqlw4SSW2K1dauJ8mYsDEpjxj6Z2qNpwVwPElxUHC1uECAShZb
fUpEAbqeaoG+AN/LwGPfiBmbwFiEaa/Q/V7tUyx+f+AU1A4WdBsYOYBCtqIcmyRa2L7es1k49ZxC
sZw7jhNTZj+7oFdaoZgxaBHE2QbWQZQuzY0/dVc2I0bXzzc3L3nh12K3vfc1qhkV8+CGneorRtZK
sQKJkpu+iF5Y6Fbm/19rUwcbgQVeaYIWOHP/XXn6OaIPL+dPrvZhWNxk9MKpLyS4k5NKTaWHozHQ
kQxZU9d2/PoGWVdaZiplUqtnc7+kxx9WcNzwqhTyvDh0PLplpLL9IfXx7Ap0gM35wRRgaL24kJTr
Xx93iehzAtacYxlMVlphcqaQXuJlEAQuF/rVe0+CwUeq57dbDEZjLK2r8qlYtxtltJQbUQWqzZip
d+XBvB/j+pRome1bmU3bC0P0JstfFpMVY4/TU3LTi3yVWEntDz0ADKi+QBOPpVexfrzjtf7hS2Cc
LZ6bG4WYcrHKeeWuPEkXiWmfb2imVBKRA3/ORNOvUAQBiBjXtALMIX1mcZx+abRcThgqSTtSH8gm
3xkic3AhLGlfWDis9GYgnWMDHd14VbS32ZuhLCS0Lh30lJkEtgX5fJEr2Q8WoL83vcGLqfJ2lbgd
UAIyTf18txEnC6fQJp+DNKciUZ/dD+qgvb8SmIfxwt7AYxgtI5pNW3WiUJzyINzk/5DoRhw48K6v
NcT6VooZnaEF7wEBkAdtxp1hlMj541uhvMhuLUtAp2lgxzUNlGrYMGYeB2L9A08SjHfE9wiW/wU2
daWXUVfS178T+JvVHmHVRr5oWUqTDjbY88oJW4Y7j/Z9xuKT7M01Z5KRl5bMs64WCOjMqyFPdqHY
IPlB5JDVxWBMmH6VdMvJqN8xM8W21paOfB7dPFiOYzD/V3UarJoPcMedpayVxMidnHq9m6La4rpx
GUJK+RhbTZxg2H1cr3rayruOMH3goYoqEVbki2jsaXnZ0erFE8tsIu3RN8ins6wBw5FqyXPHxp07
CbOX/NDmLyPEWqWG/oZcOVVynbpPIGrGfa1zGc7M+97EYg602ZZWAp4fEdZEaUvQ7cXVhc1zFjZW
vxlTFisQRXzcytPBfPMFOAHM1QET+FWavj7bPafnmMef5LEavlx7Oz4+///1GuDAhI8KIvdADvc8
hX1ho5dJSjuelc8r//d645Mjz+cUp9NKu2b1qIsniHon0MIzjmCuNyLXhABrb+yo71WA3BY1/m22
LPI4oQuziR5Rj7WUFwFpFmhe6kHUKhP1vCbgQiA0wapDqRbDWDNJTH22DELlvR+t4xvR2XPClDCA
VV57/MYisnhNNhutaWpj3esqoiZXP/m+NkRXy6YgBOnka6u6cZ8qmgYjweFKV+L1Gs2dL9PaXMfQ
7qnC3gNR6VfOGywHeGJ22rYk9QFpbE7gkwFXaShXtR1io0efmpL0PZ3+SmC6qHPHnclfAkwh/l/2
Vq1Gm2PyhPs1mfYc8CmlCkJ5tdbYZZEAnSyIbtWmtxz+NgHyC5zTzRMWlfTXPHBk/+OwHfVgonrK
DZilAnLBdvDWqJ/wiiF0sgpXC77jvuqao1QThwzWyQNg1ZAozWIYsClMK4uZkpRo9CtF9PTCo29y
8NkvDP7YRhDy+DVgkZa4EO7UsUhUJes2vQ1aCpc6LOQJ0O92lfZLGlDZwL0vmD6cxggoyLda+B0Y
5m6UtvltIJgUGbcBuBExEpu61RH9AnACv5WoqsAnaIDHUqFHXBboAMPyM4I7lU6MYhcUKJEKw9RO
nKXv60nLqlWkorcWtnvg7ssPSDUvUsHfDjJ06KFICZNKmHXOBOKvKRKJ5AX3u/Vh0pC9Ou3sZk29
ap4NsreowFbEZZbeKkqFug9rbnYfZ2qmxgBw/1/NaTu2UiHwRV17oeL+L6XOnLFeXQoG6LeYmHKj
BzoYDAup1KP5a0UFAebeGSeN/RwKvDncTS5M17lIONQbuiid2nx6QqL6aLmmITeImp+0uSo5p0SO
G5m2g3TcpIazMElb55mgU03/BmycNbvAsOo9Xmt0EMSAh24P5Rv/HFQIlFcPFi5XhOTu1yZ7tASl
dvqeooM2zbIWqAgjAUbLEvaQx5tVJuHSDu8uOaHTBjgzl9dgpv8BoYq1w+nliYRhtk2JFDyHWudT
lnAbFcFrwwlnWs+2tIjmvkkcbvE1z4FcfDgk3RUvgRgmOcrFpFGdJTmOTJJBxAcOSMpnXKRya0qw
41lJAGt5oLJyc/eMMYcZLFXwegY1M+ioX+9G20xOkd+hEj4+TPwk+3nHwzI+/Cp1G11hijY6pVQa
gFFTKjxD89CF4S2AdjO4AInRbR7kExa4Rn0TE8gwCO8fxbOxnjeY8k393NR9RGpCHnxXWs/LtBNh
B0HN8Z3+W9JcookBtELZlvmeIqLGCsMz5CK5Em0jqJp8gNNoq4KywwillmwoBI1fOutmvbIx5Sle
bJPiLXeI6BMo0a0lu1NZdbvCZVAguDaqfoh6HqxKz81dNbbpt3E8VA6YKjgFjqixZfaMs4zsUmr4
7xFORpSUWd9Zl6UIOpevl+/lbTkc5NJqYs1U5clXDqJA0rZ5Qq5GaWgI5q8nGR2Nv69QJVP64pwM
kIhSPbZtpQL1o+kXAZkKos15VApZyujjTgOAxp+TqUgx5Etyp8226BgqHjCO6GUCyXscL3XN/0Es
qQjOKbrNsrtR+J2VbFQb9LTNB9944tJ+aJugoMb9OVf12w2ihgyhyGLlrF1hNnjDn41meygEuvCn
UvRSBAmOHyHjmnvhxDnXetcHBCZSkznyv4dUGXVHzcemkQeiAUWUNarbgTg5AbA2WsFQ5Wmv7u3t
OCZhg5euST5xKFC6Vi+kg+GpZdX0a3y1uXxDMsbbH4gY45RAxTYZJDlnqgN0nLi5npiSnSyKlaev
OagQ//nhbHcLpfluV2KrDIcwSmTPHULydr7wyW4mOq2yuoDZWbJb42zYT9s6I1HrS1jyIhoX15BK
3/0Tf5n1IGx4CRi8GOwTVg8MCA6glI4cOyAor6b2NfjJ9QAsIzaJjbm5LlzMARu1qKmi1RZvXjX2
4ioS7dynlLkYoZWBu8XSExwe505Hb83K8/YcHLOg6UzR1TMcwFoQ5apYrhoJz5aBiz9RAmUth8R9
nhZSbL/zXsu03/F6gtRfInOdeuFTEFegRQXCGyln03G3fBUcBY2Hv6THNyOQspSO8rTwYpHDLBmA
ObUhS+OAhCVaMlM5EgJwsa0/fUVmRGOYr/vGEyXGOOpkPKTy0TNiRHYAgNPVEq9lbpT42Uc6kH+t
oMVG8dfAQhYter/DVb56qwIQn3ffCPQ6fUqmNGj5L/gD/cjedlASbHivjnmGh6RUKgc9Pq0eLmBU
QplUt2rjepTDHJZdPUYwJGSZfN9vyMjRrky6nCfbfKC0Ke7O/l3wwhFhED7qhhi2OrLE0xYsKwgy
PZXzXJkgvSbyJ002T6WjUeOXIC0FS/JOfsjJ+1LpoNhJVCTbkGb8dRAMnuxRMUc4WOfw4xSv6Ltw
b7xItQGvU10ji+7LAL+RcMcamohIyaIKZbpeqSjy9y3RwUUm9ckGNXzHKxXJMSiLCF24CYsiujqF
hDvydI6Z35PN73fjY/SLnzU3LTd97J7cwMlCQ5bOu9n6kQGclSCoKanGj+eoCAAMCTRGy1IbjQCA
PGbK1VTw00kMD6CYM3l2pOv6PXUd7cv+Xk/Cti5KeP2SMV373GGuWhOUWJ/+Bww3Jf05txPQX3RO
NDIDRjG1knswzxiw6c61zRSlG+P1n8zU/3xNxeDK2MetsCQ7QVBHALPcvzu2THRzfzUGmzGKTJ48
gVlk1F1j2BSgGFi2Xfjz2t3wM4D8pShbUWNx36bq2SzJy1SAgqbmU5ld7VSvYBxeI/H1Fdb59A5L
3BzpqNH6PcM9gZPq+DHHMRrCIaQCWvln4uB4qwM8ZFlJUXygXEVXgPWT7H84jtH4zroPPVZ7Vurw
++LDSrd3JwYrQmitpSwQkWZsEPPYKtW6wsmZtpo5ihuKjyHOAGEHmR4SCVBXojGd0uhqoMao9W5M
n36tumXKSHOusveFlpZND7XHPOoMbrqb9xqQ21FXGIT9FW11qErfh7JgywHJpsdvGRwt1RVjiEhy
IlCtdTNCStye/pMsxtZcORJbhYtSdcp2KDu6N1Kt2+8jToMTdFOQns6F7ie/L/fPnDDB1Kr8XaAD
5vsUuXdZKBytAcpnG7CUdWyowJMN7Pt1ZSc4xsU1kLLBb3jpqhrwDU8y1rrCYIzDhRI1H/gkfyEz
BWv4G033FKIsUSF/Ryk3XM+5ofoelTzlCjmat74aA9U15+1MKQl0HMTe66JH1kHtSue1U9w9TX5N
8Pq1z1vK964U+Q+Qw3ApB1iaVvIEIcp2NokR3ZIVo9oH1rzbCfVjA1o4TNR0W9rkJB9LLpH2YDdC
mActI8sUdg3uHkY178jjB6Ujzf9gQ17ni57J/ilA3c1Rq6YAf2T/MrZbP5rvXbmmaFeAd5Q0f5vb
gWyszEs7Ub6qlYwy5xWA529QYUcRV0uj0BIISqW3u3rdCfBmDrOlZ/uFiC3W5fRsCs/YYPPoCkL9
dm4oONj9DYu+39lhbCZD1gx/w6I/X6zAdI+f4Hji3szGTz9p2BM6v9qkBBKlWNdLRa3srWG4F9w4
hmJ826X+7RoPh2r9BJTbwThzoKfLEQ3unWmnlbu87Jt4jgaTGRvlenaLS4NhSqV2qOhuR5U5m0cf
5Y47Uez2a8mwZvdL5oET18fAkjpIilAS10EvFAVoGFQ5NowNrq2wF+dTaSIViGN+YNbA6eKGuaMM
HYS43SF5YL1zQmIDzNhquUtlVc8IyCOH80/Vk5SRT0D7w4LlZ89/lj8/Kum5sFStfOhR9vNx1I2T
bt8hdrNOQVw3Fot0Iyrm3Vp7KbuaUM5xJCaKb+/Z1UsLtKELFPSr2VCaNMsWyjm6sLj2OMvlZHjx
JpqzS7qYxSs5jeoTjtw9Vkd+8GWHcdP/HjB/mtYeV5qNRIKbGdDD9teHHENirCiFy12ryrMk7aZ6
bEEPpgqS0Z7tF3TMHCvMWPeXRqsJHVuhj5Uus1ZORXrbDRpMDYdoBGoZwzInI4EOSVKJ9RGQDDY8
BYzE6Ipd0U2fsyu/xksTUTLRvgD5QDyYUgfoKvbe1W4qNozrgRF2flxbp/F/PeEFs3Q+tUiJ3TxI
6Zj2GQSeG7K1+82zFrHqdsK11/yZUgfMwjiYPm5NY42SjiSxiOQfLz9xE2KeFWDLK6YRgZO3yP9V
l9eOonF1/CKi95NdRAVHXxV9UKmq37odDebKpFFEI7m7c0Cf6JWyQlZ+qX3v9OL3OKrUI98ahv4s
Uv3j8D+2Vv42VmY67uMu0pWsGhObsisCc1PKAurdCs8+ZFDvMfjHJEQZWU4j7l/YCQkT2nuI0Bx9
YTB9owzF9+pQ8CmywCmZjYCXb8dIbKjVbi1SLG3RkjvM941HdbgbrTLcCuz9o+bcTuZt0CvzmQAi
nNUP33QDjLPXp6WJKKkRQTdm6DrNPkhazbjnr7PKgBatns1a48XrVoDytmSnrU3Fd/6g9bFwGKhM
c+Bdx3Rq3YXD1rj6oB3R1IXZ9+QyqdY4hi/Rb2c0Hnnc3weYJAbS9CXx7oEA9CRSMs4iN66KiCRe
IH8O95clOamrhZS+si833oRlE1NQRkyvPJP7dZHBIuTxBeLwgnsHr5MVD2shxqNZ7tk8Q0wqh+x6
oCyt6/LP7Wndz5bre77Ip8bS2dmTmEWkWdhMm3jWVMc+su1pqLoRRcDDiaOgC4MQhiHB63JS17aT
m668A2CFy2cU/nLfNpnHCdxHwg/0wRKoi/fxXpSdDUPaABRgFyASzGRqmuUYopQ+F1TAN2Bvrm+3
cTFx6acpi37Rv63EEaEQ29oUeRS3PqtDBcecFLCtOyAyQghtUpU49hQUdWIosGrcNj+OhnS0+od3
cC9/WY5/a3tK1PikL+iHUQpHcMN7kl7RxXYf6MdGttohbcpNu2PUJfxhypL4SEpv2XjKpSMTv08q
sfQTPwX/IzXdql+QPLn+Z1morpKUs27e/qYpEwZQoj5VQnNTX6tFog6FgXstTzpDpD8l7bme6AqM
lOhXgMUrcfw5Ac7ZECpHTuPXoqypA/omPBaz8uUoqep8LAil4Q4odUTCwZCiauqqVdjDFw0qs9e8
k3KLGXB2Djd74tuw+qEW1Mc2w6zWoHf6erE7FtE6xNI1/vWDJGDtp+UXu+9ez21P6KSKOy+kz45m
Ksz8so/rlgQAFtarLmRUaDkpFBd5Olhtj8ql+HkQqoQUQbPTUIWis7BMbhFW5eaVIWqdIKd9DG8w
X5YNcH4C/TCXqJ4WkPiAfkOqfg5AKu1p8oi0vvH2Ep7jueMx1XMGXSk7SCObeXH1jOpWaDM/wxAv
LZ9/vKqUzv0Pc8ihORwSHLRhg8zdPxDVyLBY0MvOG4HgD2vWQe86eRNpNScviMuT3+u+11kyDY1q
VjsYh9S2NUmRkUQ6XDOi/wwdKgCq/KXYI5cavgeDSUA2hnorxqLj4JsFS+OkuxVDsqTFYDd+msP4
IpnRws+goMglALRHEN7XpD6CW9Pn2u0/tZtUzZirb8jlG1xSWjNnOmGwHPb++vPccTjMT6tURp9l
nY9gmqsIBqx5AHliRXUNzDpC7TItBBRuMj1jLEv4r2eWVAdvsUHgp197LW/IZNxusHTDswpppJ0D
5LuSAPvQRnIwy45V4FKJd/A82KlOKtn0YOPMe9b+mgSruDnwW23Mbv4DXE+D3Bhrh4OBaQthPwJz
bkyuS/jvykUM3Idz0vbKHjuL0+rH02PCtdhr0vT7R5JkUH3YR5hyghplYBLViFpO3LKe5/Hs/0sB
8rvogAh/WdKeHkfGHrs41k91G5ZSAKYBnuMB+9Ibl6Q9As4/tMcrCVzVu9GqShlaaFotWuEPtuQQ
tejmRAPdaEXz+a+3Jgw5hhih6INM0AqdSkBPORjfVwGXfQj0bk1B3Ajgh2gkOXVG4L5Qg+WnC3Iu
KCPH0UHItpFw8mDagF5/6eYQXnaecO5TR8m51az4Zk9QJvXftJlDF+FrV2NgOjSMaz8aL4lDdRi0
JQe1ji/AweQsGgtaqCSfckNNYUoo07Y6OSg4RvGFTbjmf0tr7OcyqmoYsJr+Rno82LHnWP7eM3+F
fdN9zu7Msj0NQhI0Kow1c22BMTVjCPMiBwEcItbFJC4zsh6/8m+HhiBDURAvbOnjyldalJ6lgKLC
VspTRVCvM64n0eR5Ep+rKH8kY5UNpSfwGdr7sSqmmapA1jef4r+vz32CvMFaaxslJU6ej0r8nkU6
wQjQJtYoL3DkwM6q2SxQgasK8zZ50nIzPCulzAsSlngDcbiQUqA6ZSmWyj5nNDbSFhzUBylR9PC+
sLJAP/liptaRzkugIkJ9nfeRDT8XZUniiPdFU1P5HMhNo0eUnNetBYrexwftIxgSKksyGGsdQ+Ph
sm3wk7lmZieF9g99NmSHURYuGIzPScJv/JKpSBdEy/ZNVteR8mvqGcYz169Q69d9n2P569jFr7yq
a1XozwsgYmhcxrQKiigIjTkLZxi3vGMZY6Up5+roXGtnPKFduV9nF6bWZrHezZ7PkHAqW0B5tmOs
MrcIrPxeCnuibroGLE2c+B+XQPsu7VUVq6Q//UvcpBDcy90g/GOty7FL/Lmvi14+S7CCy8gnbX09
K3N3LA7N0GyQ8sOl2HL1hV6E/ZFhin7WJ2ZCSigWUfArfA8xFO/2Ovkdy5BaI4wqMGdVAyxpUH0g
1taDDAfRAu9vlgIEReCPw02mXFRVjcOTG9al24HC9bEzri5SbEjB6DZonsOh/77TCp6TsvNIvlR5
obZGyU+6ePpjyAgtosBR09m5t3VSmSexU7Ta2E5qHhT1jgeh7bq4CRVrT3GBpY8aE7rEX3qsFz2M
FYqIYYgwZETbmuj/g+7a8SgPR/9C3Vfxt859p9bb989BOsjxX2mdeljiEaTeDO3O3ZXAZbejS/Up
0KBl3ZiApwK8AFnkC44KhoDgm2rM6aXl/VhpKB6DIzbMBR1dLRNVzudOqqSlhGAEeuogYT/G/OPJ
k+uzbarbjYh6NJ8nIxzoQL7Ww68qM7ZyoEsck+dpLRJcjCpa5U0we8ghREEAcoqXdrW4rJkaKXWo
rKFpXam7iyiXhn9fbCXLOY+dIEvg4iYtOocwtw6Lx4rIfn+YzaLFVGDswD1jNeAxyd21KM8loWt5
tJeOCI3LmYG88V/w7elkA2JV7lJCiTJ23ergpaJf+8J4RehpAqiIzkcaqv4oZoq2Zotx7Ik2Mx/0
ioUTbK1KfrFw5uBI5UbNCC+x3ZUplQ6tV658/qGWOd+v5WQxFo1RU2rPgPu9WmJrYiy1rxl7TFAl
V57MlN9s7AY0eF6lpPCYgkBO1krjZLBulaqHVGY7uCIRTwItYdND5/1t2Epusn1TOhR8SizR1XzJ
xMwZedzwy3iZN8RQaWf1KZsFNbY8wZ3KbBomKxGcOFdWhUoxJ3GABrm9YCVvlpDXmoNE4hTBGFd0
VWt+qHVbLsJYVfN8i7+/mQ5Scc4u/1Ljt1tIdw1i6ru+duwR7Wmq1akpR48Qo+6+byzPNR0UYAOu
8yL7skhOml3qV+e42t1wNcidZ2Ot+h/1HNiHFE/8eF7QBnBnKZ2Y/3IpJq2e8NuK6rIw6UNaqdL7
4FCGi5covkA/zInB48zPF48QyxSShrXGb1zaLzF0Ngkw6GmyYluDibQ/im2ARvH9s4Vymd871dFp
mZwS+eLNM6Tr4Ffnb+A2LGKFFtQT2Ua5w6NqdL1pV6wLeTlT2q4lXZtii7L3Lgud/zbisxEj/fPe
40AZx/I/V9f7PT4VB+7IJWy+hsxaXYHkDkc5adZTM3q6Nvhgln+cF36qV3o1/lakNulruUKiJrc7
TJnWGhyxyudNGp/auyBZ+UuNPTO66gpZFFP1PIvDjlmPArC6YdEqQxzPydTUZvAOk/b21g0Ra3Db
XG3IDIgHJX/5jwE7//qM75L1s5tDzX6bGH79uFYyQHPhpPc05Y0iyAX7Rf8a71cbTt6NJvjSmbgq
61bxEuJ7X6h7M1RM/WnxMZ8qoI9ZQ54bRZNgISl8tAs6XGmGEe8KY7kymmUYOwLrYUcJDRSwsOdi
Lg5JsP9g8JNQgSWMxpHuhuwCeWLvDAfJS3eWWrPMtFGBQi6721hIoMdfL+nEf7boO3PkKZ7zYrXV
1JLcXecb89fNtm11l2yzBYSbSQh52/KGx1k8B/tkrjxFCjj3yhv/mKnErdPgRFXOcnH3hf7eGIue
0mmliKC1NhP/C0Hj+8ZhwuGRAsetIeAoEWHI1NNLaIjUMcJHaMFc5fKafkAKoeDQoBCZovBVRt8F
C0qGbjQMX4nFlEGD+gCdwwg8tBKnw1a3g/tMhds7pgStHxeCtBPUJQo95VOMMJL2pwHPB1pBHfi1
lLtn5fX+jDvOEpY2kqEaukEpOC8E4wk+7cS0NkODNpDF6o3Jy5pahMWFui46FLuKe6bJfNQyQKi5
4KDFFRIugyu5VhYQZQObXxi0sEdq/BC+yaj/2x2dCB3XgKamxjCtqbbWqOFsijoCyX6oG3vY2JE6
idjfQYWG7YfEahPaPas9jqvDlwaIHdcTu/COATuV0i97GwQbn47KW0j/okwhuur3e1Wv/Um4NjL2
V+41HQdwarqarAOcq7vjuAlg+YwF9LfsRhAKrUdPMzBltd5xfmMcBwNBl8uLnIxIIIjEwbbW3L6O
bTkv5auKsb+B1BSHKqYJbkIzbk2f1xZkg9cMNvugVarPNj+3Tc3yQo+4aWFX0B2OCp77BRK7FuEK
CqJf0oefw+RZFGg2QcUx1ouES2DtFaEYqRg1nbOc9fdOTvzroGlt2h2g8FK+xiI03vcfA2mvCQeP
cNQYHMb22CYcl0cKzFB/9gK5IyGE3i/x2CoKyLG/xnWPX+wVtrANpHnndZHSMZHMlQ+ZkksdfmCi
ViqyzejplDxYEaje67RYqg7OkYwzhlqUYTIqCcPeL/v4v+bFEvn0TQtcVyEDDoO9LdJUv2pE/AuK
2l2sGsLvgCGrjPmdjBt5LOyJ3zggTrL14C9ObFdtSv1C7rlMJ1yddM36fs43hU6dkIp1RGMbPYwX
ReOTVn19iOA08+OFOpQx1+kloZBo9XyeMSoZWSFO9Yl9lw9zQYa+WnqtvXJ0aFUAKRHBnkOyguoh
ftq0Ig0OQb2UJtqE7yZOUc2Uv8gt8FfPXet/WBhtZUEjN0C33t+z+aUYWE4HE9KzcFe/OqsTjfyA
VVCTB2yI4lxLWLYLe4BeJKOXZrtWgZZN6gC3ZcJCzQdvR1s6/wk0RLey6BUW03FZHIHK5BHd8S3Z
KGQg27N2uffxqIEogMcVe5ewIDzB8d0nYcjbT0JB53ZYsLtcCa1k0yh4EGFGA+hTeav7Gu6m3Fig
ZDJ2+dkRydOXn18u6WZvXEbbaYdV5m7FJ8ExLoWAHgagm1MZyTk+4Gxmk/uP7uPC55zcaOR8MqLw
NUSEmpDRSgo3wCGleMApli+hZg4lmwbQ+C6yrfp41eVeWSJqA1VNRs6l76bv+ymCrlWa8k2q5mm0
gxGyqlTLwIpEm64+fQG8MNnS3SP3EdnJybnFhRQO20o/vM/thPNeqOXheQMFGtWNg4qJ4pEU9Uf6
Jnd4hEcZMMOlxRAWMWfUQ1IJpOBHV5OVPlvaql9IHIW070N/H28elY1DnwC8vogp8Nog4/6iAH7a
uT1U+kKuwQQ/LSqfuD73TReN8c3ITzn5qQHSNy4Eej0hV+/sPPPIERUxj2HjM9iM70hP6UmEv1tU
AJA7TgAi6HsiidMDVkuxeAUIbe1PKmfQNf1JxtFbQsxFTVxXTE4N/Gvu/z1Z2Iv0bZ5Z2nWcS1q3
KtltwCzbkUaMYnqj0g4KnMxOxm3KkgERWjAAWA7uZuGkKOLIuLJAoOyAcP1dmQ2ZSVI8IyFZQ4Zy
uPDBrWi4YeFiaxcJRV5UR4rbpV9+yqsRLq1suAEKcmJtqTP/m/lF5YC//xXEZxnr5Dh7HqX4ScB0
WUW9IrloI3LCbEY/rxHR9sjIHZ0ugvLiVxyFWzbKdb/RzDILmiwIdPjpDOpSr9DJC7Rw8qhjN4OL
T8OauSmvmqdUeM1zrZnelEm7nmTtQ0iqpI/ZYnamHNWm5+2v7xFGnZ/qEX0DprTL3ga0ugCOTKvq
jLVWjeLe5G1aHg5VuHnK5LnbgYgfCVXXqPy63Jb/0jAL7v533Wd04q3qK2Scy8N3IfNGj26CpIr/
0fMGUPpVIZFpJdUts76MBPOVLQKR9HhI2nDqpEtFhuM7zk/imA4/xTzinjF03OGfyliWklaESMSt
elr10M6nqfDfZBCPi0dfQBv6dAX2AOY2g+iLmk84SEVEqckmr1Bk9nANG/sbz83Xi4ud0jlx+l2a
uX8JbqJFrFQtRlKxtXZJRYRhruKREDSDVhW33nRsZRaUjHVKkCq0CmtM2bA5ZlOhC3Klv0zZ9A9e
+B8pJtEe//bhBNzo/0VcGSXhCZqdTX3ZQACYW/tAM8Ln2JeZCKiXp0tNRs/4+xFz63U4b2vhNkvX
8n8Avh+1yqKminf8LVI5NZbdaUoOEuL49wpaiBkuetvXAC9AwlhwhlmzaNpNAe5A4A7+OmU+leK0
+02jfY2is6HNPmRXCzwDUvZnwHYnowMNKpOBIDqmNHJAv42Z2/NFeI1WnpNl6eqiHTHb96Gft6VQ
mBgQ3alRmgA5NBEOLsNdAIX77X1XSF4Z58dMtL+2XaMJmHKQn7zITPU4htwZHqhbPHpaZ8TpSBje
wlVp3GB0O0L04QHEjUClq6cXb4u89/5jqSJ659apCyFq91VlBco3G/RGODB4plbr7ELW65GoR0Tw
bWSVtYPP9ANiUJUYY/I8QvCral2Xv0L0xIetpeCnKVoW5w8GeSiB8NsPnObdbzhLdQiZ3TXBSBKC
sXIf9brboXkzGwZAD0ZmGSMfjjaVxndCSSwk/exN92mM0QgUFFAmpE63PyCxJwPdcK2AwetxP/GN
DIK4jkMI/fnZG7WKBBLlLPnFhVwnJIZUSn0+7oLebCXYdCLu4AdrqPK3Sy1Xkq4HqqOdJG1wPUfu
2TnltoJyotbBFr2eeyOPN4eI8Ep0iLpLrTeFq+Hznaiz9PNrUOxQkVanYiMM9zw3NO7Y5nLdRmS1
0GrlbwVc5Mmho2YQvXq22IRxgunSdqJyeCIegeeaXMXuQcVOjM1RWJikKz8f78Lw/rwRJYv4fCYl
au/jgYIl7uIlrqwQhp6fq94GNLF9sq3IouLhhVTRZ3HnhMfHNXFGifL8pervkP0N8FH34hIyLBww
ppt6MDpEpTVTJ0ZjC0Rjq9uKjutqlzzA5fd1qxvUMSR3PNYHZJnXbjmgrCry0iBnNhJz0evbcImQ
+bWpQ99+fRJb1yFCMWt3dqR0TzeBRXgVlvf9NVqvpTCQgVqU4Nz/kn7b3kfUI07EKAPIkFDlnQrW
+1poHn04TtBQdbG/K03jzE0i+wudEv5RJOE3YGDSUckUBINb3g+tZW7rQTlE2fHOyMnVBGgoV13q
DCVgLXIOGpyE1WDZJjYf1gjxNBMd8l5Xt1KndkUO3TtHe/W1PqwDwZzvRn7kQD+iLz3wOPCC/qdK
AFGgV4Yf2u+A2pdwkIEoEcHwauEL7Ebf0udA4w+N8Z9v7hB5IOizgwVdZ7mQCakCkVwmxdRO/vHV
80R9MJjsDHvaO6FS5D5Tc/OQWnUcVkzNPy6u7L1/9yLKxGqhAGILaR5wsfqmSWWpPv8uXbdG6A5v
YqhbtOKIfUk53Rbxr1IAPqN5YnQn7xuXU5caiYJ+AOX6H0t4Q6cFT2MuooPSz4qtU/KPK1mNz2Sm
7G/pQqxRlE+yvZv5a08LP/gFWXaGB6+gfnJ9IY5nBwQhKx1kvjmuftb4S5gXq+H7ykzIAWT2us/0
2x+goGxqQSwKXmhfdS6uCW5kH0Dsevbmp3wLRbxcA215m0OXLnNWklWWUbdvgLCdI78drae4yA1Y
gnxfOhLKAF48ki3UwIuabAvXE3K8y2pY+xtXyina2zLlCyCZirAQ4g870jRU5CryUheEgXXmRevP
J1Kgbck/42fDXqc38hZMeCrMmJjVMb6NygYxB+lqbfowTPbfDxRDwn6yNSq38R5AnCMO7g6qnmLj
zeab5GXU1oGJYZytwzf6VoK37ZurnAehon5NWrGy2BiP+X8GR47KuT+3aHBWVSKEe9m30IsaIJ9x
6FTbrd3Y7/zYGZetgc+NskG1iEnCQ9KYEzd5S1NV/lWfJLq7chwnjwfgUCVVvsCq2kqx3N0ezWxz
QCPSCPsX6nxT1pJUuaa4BTqJUoI+QYsZHRGe3Sfl0bLXKWwKyzz32eD6Ht8O6AEhaRnZVk91Jp0D
S4S5HRcoxbXELkyoE2s1Vp47A77yjG4eBJsUl+gv04lUanWS+S+kPgIxWRebxwIng/izAuUmXgck
lu4N8gWvYyxBt05LPh/orruRLOMLl4DLEPzlp0fl6/01bRHh+XjRUpOafSmK58nbGFHxLmbqvho5
laLDDVDUIwbkK6U8gBrJRYvXy/JZqq7O/J7Va0XuThs7sKGnFd+pGYPj7ZWZ8R3c3PlAJsj5K0ij
LB7H0kt2BuekD/WN7bl694IyqUPN7BpKFWUJ6n2ubGSt45/cQlLcTRsQ/lsEFsXzENSFOKLatobn
1xrUq0sC1iEoJeAX79fOp08aReI++izTOQc8WWmOCFzgYJUSM2luTXciGWSrm82rCakVsKlzUGQa
WSyMAFJKzfcs2NFv2zBqAiNbA7O0s2M3BeFmnTyh84b0/PfwL2dhTAysudxkRWcwGMNtTNO0Ora4
JOP0ewbvAOybbSXF2eWIzrtKGiaFOU5G0tR4tgUoIdrziKp2algbqkUNShxb/N7WolIMLiaL7r7f
1WDZJeGQNs3xUtz9Ee3Q7/GLaj7f6JeCCJTn4Uvs9nFI6kBstZq0rCpnB/smTpTgB9ym7D6300Q4
WiDX3iTHVq5n6JcGIbCnUgXpnQr31KNCXHdzEfS0AuWVpzijN4y3vbIk1TF/UEdDzNV24nj1sOls
nHgXsDBS2OAdzTf+VuSPqPfPwWScDgLz4Rp0ZIyquvrSWnr8PV0DiLmghR77so8Ml7RZ9q5skoSt
ybIhrfOupjzjfFlPnG3D419b6dk6DZsCeSVlhlvZWhwD3HMXp8LugBoIpHdCN7au+1QWB6Vn/+Lv
fxweZEngB8J0XenclC/mRB7SCOjDvM3eGLe4lf4UMKNK3O+5rZSQRvFB1OCubzEtMkrLbkYu/h/L
o17ZJ6Bj+Hr7+g7kslukhUzuOMQG+vr4e/B+Nt2tk9TKkk1o5k4S5kY1ausJt3Wfs6PTPeiFJ264
YbxKl9qET1qYTUbahjyP/m51JPRZV+VftEvRaOZMw/chWqrF8uUwrBB1IcMSxdsq7HUD1P6SSM4n
O33TXUYNNrpTU+mhK2QGvpyzzVB5f2NaJkCfinONOpOMBMIqJmMTqc7zRVsD9WCIaL5lNgf5lJtO
2x9B/JdRMxx37i8FeQUVBkiDRzTwprmufWjiv4oh1Fn+6gc0YfeEQxNnQmKc2S2xwWpeV0GEMKJI
YLW15dJqsivjHn0+2O9VBd/VscgrifqmGoZbW1eTep3OddSYiP7P5tKGgu6FXmORc8JrjKE8+PSH
fH0qm+wK5++LuRPtA1LqBldOPWGIYAHeoFUxGsdbHgK4Ceg9ibE4oUe6G2eooNKpWObcOssi4xg3
np3UekWwcjXteozi1Fm8DqKG7ilNOqZzL+9w/IJpP6JEw9e57VwH7l3ltnZnH/G/3H53R+vMkT5E
PeqxwrSznxw1FveKPGZuZiNQvqLh3Mnd6Es9BJ6Wdb6PWH42QyWvjKbzUMs+pmUWMVquHcmG1LQT
Iw/1HnCJ2cPT8jJ8BAEv4AlP0x/eufJ95jT/IQK/HutZYT3vSogGOAMIdUvs+cw6ID8j6yet4fSE
kBL7XYQjqAuk9uD5q2a0uu2CJcJGkwxe14HQq0NPC9+1LRLbuIRaCELOdChxBCPKj/Sfo87mAnqa
jw0Gm69rDa0uyRf8cb2wygGCrzUsWV5vmucM1zniVV0/lsVxkgdn4K3tV2oA7wTy92Pcx3Y09oIL
tbwD0ayN52VBBAKrN50aWrCFeVex4JecaE15K3tcur5Hqk+XaafmBcwhIOUxP3GhrwvGq0k+mTre
GGAUjxKd9uUJZ2MoiATRtX6Ge0F7bc91W+KzpvTzA6YAMP85FI9iAU+MMlYO2cN3LPVBywtYdN23
qZuNAzHAt3j9YJnrJiGFlE7kFJ2xGAMGzvdjSUSXlB9C5FVCgYnnnpsbaSLAMacpZPpFKzJbYTuA
J+PJ3qEobQIdcs9xcpMJrCILsbCp/3SZl/nRKv/cHFMxqP4BZCcp5iu9qB4fIGBMfxEasAYiwUi8
nK6nF/rxFJM9zHI4vD11XXxnfeNiEJ9YxY68HabQKbnQsGutBko++m6YdaAluqTXGdMqiJnGzBc8
+CxSKDX/M83EoPS2HvshQI3QGndpCgsUWDJ5ZXa5PFFT9Vltg90lpmVVwOuJV6zjWU5lothcaD0X
hOVKtOZevl19aW9aOZckQUuEbxdx+hrBerpxJSLUNJs8MD3BK8HNFBvy7+yp8jPYJRS5CH6Umrz/
SnqjBGqjglqV2hwn+PIT937c7iGgCpTtiWJ5bvrFOqxZE7cx0jEWlCHW8VC/UqakmIPpVEJyiNnR
i+EyhfNdRXWpWpIi9GOsgArLCoKC8nqrts/JJDPH/EUwzzuNsyxoocmf9YREsYgDF7waNOenoFis
83/SYPC9iv9Rg96hbh2nqBvsXOlYn+4BRFcM9cx0JkvyIEhaHoL75WyZ5Q1EpiuX+yGvg6rW2QoV
tmJF+sncKDJk3gPTiDXLQLLBgZT5brHzNloPZTbUM/UzTMckqLBwJFniI/K9Zy1F57JJ7jHZqdZB
Nk9CbUoqsSgt+gcNSHM7ixK4iRH9z4StDgunuhm3dW1sXB0qADLQq47kfdlZEwO//ut5iIsp+OJ0
48ANbCGvydtgGMs2q2WIi2l4Cd9vKZ3cfeJH+BSE40Y/YfUYW0XXgjuxlYfGzRiyUZ+2Uz9EF15d
k3CwkXGFB2tfeleOFIrDpWeLvKNGGwKcy3oVoLcGA7pmb0xZp/cYmFJ6A6ljmsaJrHU+7D2YcomU
8rjLADvqsQYxoMjnfpZVvm3oiIH2C2JVG6ydTwz1K4Y2oGMQYOB5+oU+EkzLYOZmibWAOTJqSpI0
00iG0uVDnsD4xmRQ1C/wsJNn//uLLnvH6Ybb52y64D/6pdWtpm19a5NrSwVhU11Z0XMeZHn2AlS0
96caouPnem5TPfItS4+yuZEq/DgHJGxPs96Pl5ipnZga3AwqwgTLXbp8CqnMfKuvGqx0ypq3S9kG
Mvvpczm/gbyfzLmPgMz3PCXLcApDOA9V6DfrqTcqlZbBgCPEBqy9a68n7isTdd5N3rNkmvUBwwvn
P/pWrNOvML6cdKH7VUCoE6W4DeMYGmzCmjVd6NUEK9sfRD+E3Xexuk9nFbKMRAnr5d5HLCDNBaQa
Wyr7/PHzO9brsJyXaMukqp68krktXODrAIa+0Ez4XhrsSw3acE3Dipdly+0NN2ZY3esmmp0p1D66
znTGaeEe1biMPnO8YWIs1NhvDC22vJP0DwsT7Nv91KlQAhfPDjUHD9xwlR1ZkAA/fwVZ2JRAjAq4
2b37hig1GWdnLbunLBKY/V6AUB0UWFJhDaeeGjeLYY7/K8C5Q/WMmM35tHBUfIO3KDJ+kt8eMg6L
Q7VEXRFucGXNmr8lAgy46pGVuVUuSZIaQscvVkHdi7bDhfPZR4SE1zEEUCGSLLVAzTHM/RZu288I
DwY64l0ND3R6pXbLpPM7Vha0K2r4LLeMdyY577dHAeWLBQGsJWX4QVIIbO3YMXUdcRyhdlDVUrm0
3QYl0RS2c7nuMMq75dEZ1EHEbJyqqF+vPePj4zSVGrcwFcQ83zMffM5E9YeHXhA3QvH0T7H6Yxtz
ZsGcL/y5o7MSp/eUKLJIi/Lxp2VHKxf+ZzC1R6LM5mOfJ4t1+RKe6J4sOFm8QmN4WyUMPldT4mmi
XR5QITpFuBcaq9HeO/RDnBA/yCAX++kbg6v2C4bXbk8Upmz3VhoGOQnRp5l7xe8kEUGWwHR363/A
gj6h01EgYYsT+FIEX7v2MXCgD9TJ0+AzxUR6+ElQwC4utb/AwhASUKZXprbZARCE+8vjzBY8crBr
OjwrWOtND91/7iNI3masEfEWQqYvijHY1xsLlYKyYJ2xiq06CJVuUkdwF0rP8bKoesN7brOpVfxI
Ce7x1BirWuLWkL2mBXpRZ4qPTJy4B3Z1s4OPiGs+GJbZ8fgihAcSy3/lgJhWJ9wCUQvqrkyFl2gf
jQeE5iDlAftmW4gx8cDxM67YSpnwJTfYqTomXMRfua36LyXiEa+Zm1O5ZqK1AJb3u0e11khz1rnD
PDUYvwIdCqLT4TWD70AK2akHpTZzSWYk5h8OPZAB5BAOrlo5x3Yd9IMrCYlelYA4PvPEsR084lI1
La+cOLmbkdFhomZTmDFQgMbBZiUJEVFhSjvS1kqXOjFntSsonzGf+u7UrYBpMNJZGhWwRqrEwDLE
U7GsJZ2nMhYdJdneMpQntD2Srq0oqq2geJwriHOb+0AVn0cjS79QYQvnnKbWwsMS8dPlAe48trN2
lUj8jWYCvg29L8d9Nstr7SoZIXFOvTZfy5ji6CDqAJs1ZofgQ78DYASHH9mcRLa7X7BlEzjTkn93
Y+qwEZ7grz90ZoGiDqgANfFjzT5afsYkXILxQtmNfPcXsrz5pyhdHSnKvUUWp7od2XBk5uCrkMRK
9+JiTA2isSJ6hQfClBWgf+8/useXASXTH6DTMerrxhpcr3ofrYzfwAEamNmAQKQsDZSgAdpdyoa1
EgHdugwvMLLw4sPsTSm44UzNigG9t9BkntbhC1FmwoXMkA+/SY4I+ChNsBK8bBuOHvOSrrEzbGhq
X+qvi5D8LY+49kOXRrrZp9B8/65D0gNG3dED1CnJ0yU+QuWY/sJCC+NPOXevOZFi5I78gOEYynaY
w3dWUiYmGCa0wUUNrM8EHvq1e5uuxZXiXu0DXdQS8vdjtbtj1Wn99pP5F0CfI2SKckt76bUZS3Y8
iliUjb4Fw0kz8BfpVPlf9HQ4sSbKdOdRrV37eSumHtrVhlYgUCthZD0vKz9lmfP2sUy/eYltgMMc
ZISGjsmnIAubEC6V9HltDlqBMBz64Q3lwhcYmV5+jrh8Do1vDqdN420yiA3/aW6W1wZj/T2ISgZ6
1w7LYGh/fK7sLJG8ZB03ba38pkHTzC0lLoontJ51Fkd5oWorlKak4IJzcgkpAAlvc+1OxqLX6efZ
ldrkGdtetn0pEaP9z4Loe/TTyB/LKyXbQV4iJsXv6QeWeyntbTK8TvvxgMWcS4aeg7HLEiRwzAmL
KObN8anw5vks54l2QY+CroAgK8yTWoAqqqIzflsKX7DvP670SG1ULzwncEfxYPXNcwYDLyN0Rkuq
x6tjcSQLME6V4jp7/+LPLwDMOY/8E6pkb7rs4kMyi7qemHxUD/qHDfrB0wuGYzw0YH9nML8mAZkU
7jb78MG9Qh2TcAbMiy3KzagtvoHYDz9IKtK9osKyBsAOjvmrvHuw8cbEQKa3c/0it0bJIlSgOXsj
YAclX6MTTr6ONK5m++AEkEifDqv3PbXrkbMbjVgTM6BGUePqF0smm9hLgFFb7gz8PXNr8V1mscRl
u3Wx7e7WUXj61g0Y4i0FNT7IJHA7hLO7iLxwOMPARK9IhFjHlFQyM/WanWGa9g6Vpebq3OsBYOiK
Yk4dXkg2ep9K0AjOMz8uf4FLtyfw0TRuuGMxNFyj/qL2ZHvzqiKzSS2nQOzbtANqZ9K1mb4rHBnG
WodEtmE1mnPW0kFzov1lltjhYyPCAOoUzhFTA7e2by0LMDi8JTfn8+LV8AP+Mr2ZdLvvx5T3k9PD
977/yLCmS9yyphv53mOzEN/4xrTkK8yHoCgY5B+ah/F5OHDqcF0YzZRX4dR3FGhKMLYjQYCFnx1i
ccufaH+HqTxbqcSF+aLGIHWjHU725ETNxZt0XTvYqMFyHnrRLuV4SJCvzTBxQbErVypor3B3notM
2mOuUVUXZ2CjyB0bB8EvqnFHB9O2fl9byn8Qj+YQytDF7nu2nV3S0Dei0T5/gd1vmjCvhvX2qCa9
ezpcmcFXBa8GI/H+Lp+k3JQ9XMIG7HjFUmiX1+AY4faTNEXXSFDjWmMBSKJsLzRHKDcEfMrgKqJ1
BjECx/CJL7adek2b4jZ24V1lTCzTLaJDuWozUFJHgRUAPyBDVIZkiY22g4A3r2hLItWVGJ5y9Psf
yxmHrjvgtSO5TLP6j1I5iSqgrgou133Uw7HSpo5ugdjCH6eMJOpN2OCyqBt+DxYf2BKWxObfrkRj
eLTq9n57TFKI+ZpVLZtakceEAWpkxd/5b38fNZVFGGMwYdAY5NqREOaYur3yQFOFaRjYRe806jwS
2D7e5Nm+FOnNpdt9hPRWLYHhzsUaIIjvPi9s8mLIhdBh8g+E3aWfaRYzFhVlK+VCXStg8wVNKtEp
nCu+XoXhfkp210+/e/0w9ze8c5VPicpqOpNMGo2Q0fdw/+fHMd864yj+h3QAm3ib5FJhX352J9yM
9vvu6dWmo/LPMn5kBKGGWWMxETP6dlDDHpsPjFdwrhi8pAg7p5Qslj/OG4RjqeyJIZCXWiqwyzt5
zeLExwE4HaejKcgs90EumQihWfLBDdI3IpQtrG6fP5DjoeET7nPJYGz+1R1UH5z+h0oGhy1kKjoO
+AXWfnO3Bvvk+5ZTxK5dJfBvQpqCeEDEqT7/2UjEQiZmxdjzKRvlHSMvpqMYQE/qKAedVrepywOu
RgW5rYmece7L5j9bYQQSxjYm9/z0oOgjGop0BIbZpPLfoCsbS1cL8aPKclq9i4jJn0KytccjY9fk
UcF8nYYqSdYS+kRnj79wfcv673Ma6tiv6rQpcyev12I1N4sW9Zn8+rNt9NmJDjAYMKuUSA0FQXIt
UY1rqPhc5cTb0Rmymy98pi0Qo5zHDRSRjZNJZPVhuelTU4+8vt1N/Z8uS7/8VTsw4Hgx9f0FNDaC
z6mri0lyJXtqsc+lxc7UHUR7CKIueUTLHJ9k9BNOyGgnxdhwLaYpsVA1CPMxvK8ouj/u99BPj6gM
kscs7e67nR0CI9sInGUTlvPIKun6mj1Z3IiDfQPqaB2oyDmcBvHF4d8EUyD1aTwoye9hoyKCIERX
ViW67CHVfughjs9VLynbECLhrMLdIOsP0pALLeQmeeuh3SGYjSmGL0GkGhIwZEbtZ4wvB0he375c
NOi62aqky/JQfDe/SnPziDWVQMI5cGIafBxm/46K0pwlMEOJ5pqBmnnPnV/hWws5Xyq3S2NEvPJO
mZ3ktE7RIEaRabIT5repmU9aSz4t8erFmj62fS7Uh82xM/WWLQCWw2OkiAmqzHRYw9yQx0NTGyZS
FUQrJeD5tyqNu7+ds4YpS4hj7/Pj+XfQTImohp9uN0MlPk8XsE54Qo7aEZZyUfpKdpFvgM8nz31Q
fOnkqXqCKR2G7Poii7o0C/ivvKSqPL4gd31d+bbqb8JBXWu9XSzOkHzhtJvAf/PmI1StOOZXJSVR
ft9HGIyQEMGfs6Z6qJbvEHJF2KalbRiBDnY/oNXXrHFvsC1LqYbyUF0Bh4LXHekjyT3ckJKdvGFD
jVg0/iv6DqA9WU11tTByf/khcR0gHaIEebfzMvHkCSoPeW6oDFwlH2w1AZclYDk81DZue6uUtlpc
C9/ahYLKQAI0ZjMjmIrVDhvGaJtVF6lmcKDrjc9P/Cb7+5yWOX8BTeKiw4/wkngDgnIZXsDiyG8i
wVg4IcRws1lMN9h6OrG4DWs8uXC9EA5LeObEIzlTdejpRug6V3JEem56WL6+8O1ft2FNzQwsI+XC
PvolBHewQoJ/DyIkZQao0LzINhyXol9TJWN0pmT0rmsoK4LalRSJYLHkfUZJmfe/w4Rk8zv/RjjZ
Q1JFH0IgEHW/k1cgsYwIgOAJS3w9PYpNOTghkzSSBAFsaUd18ptwVL8iz10hDlAG/D7lUQL2/w3i
/pJG8pkO8BgQSSj0lMN9HG5OJKRpNOkUlNtConQHvK0RcQQTP2r1DSrMUL9s0eVi7y59gRcLFZXA
tB/OPn1BHi06NBn6c1yn2KQlBdAZ4+GwF/kIasH3A8DWgqy+GAtRs7BIc1L/OFOGdCkG6QpUpnOT
ISO9qKPkn+T/PMfY90PffaxudP54HT8AYJW10XCuU27F4p/Th5BEIvF7aq26dRWmC7f5M56AeA5a
xAe/oFqXuOZ4ZnCYV74FLS6CDmBpEqmjfjNADTzOv5xCBg24i7iZtgNj6/nNIKT9oGZo6KeqLI0m
8X9wrw2NsoEIBHoKkSSlxuo0pBm8PdCiz8Uvin6Gjk1KB3cdvVAJl2KqWNbb+2of2LQSJZQyynW8
SrQRWqaOG88cI1bDg0RhQKjRlOUbt43eobLpgIiqahIZtoqT3yt9/8mWNeVrQ/8hZbtyjyQrZNRW
Pjn+2wAPCmTqKq1N6jwiSwpO8wcCd46GsBxg10O2LEjRoFKpLIyXRBQlfGeQ2dnH4FDCKZ5Ktduw
5c765nv8OhbWkSa346mEtQFjEMcc1O9uCJ9OnL633M5hH/DD5+TOulx1o4q5RwZtccP69NRAZfr+
EYNvuusF3adO02xMU6EkZ+z1cxT6Oq9+UTBITUr32Lw8uygo71Z72vuHXuo+xD5A17HNs7btX3Y7
8hHuGu2jjrkdRgFKtntKalyGHz4eIXdLvlO+b4ENr7xdNPMr9Vz9LCxe6WeY1MB6M3TLsFOhKYTF
HVKZwLvalaioAD+C3npIWLp/KcwILZv1wh6txD8C5wOCvT8MIUtWdZLKdoKvr2SPZdCkeWiX21tv
rkkS9v7zzj+af7Cxh/wVqLjkrT97Gok2g40IHVmM9gK9oVh2UfbwBRQQnTo430gCheBGqBDZn6KK
IONNPU8A43u5KD5JBYOyPJo/oPMH7pS5XlMe4fwDc5RkPQOMkz/TLo5/LgIrYVEkgrSIQG2P4LON
r9lHHuhONzWLFwxuulOBqfSr9tU5BrGUkLxY4cBupRe+x58YC08envrcZDIo4vCglUhw9waV7lep
MndjYOn1E0qhyDr8WQlRUjI7YhdLS7ZWI6iyxoBZAa9WIfFn0WMTvTMZat8m6e1AqoqUlDZwoebu
6QrutzePFp8BoPMi8waU+DvQsSJcFUgb1X6bPjvYku5h8qwKbHC7zcEF63qSwSfI192sBEpxw/u3
DDcQwpFWVCWHi7Y/m0s/NnWv2i/qS61rbPQPTsQ6YFXaiRymlMTg787sWVX2/+5Bx850ZcAYi+ZM
Ct+aS4zzAEC1lLUInk3r61r9yXm/BzZ9OhcuHfFzYtNduBo/z192tVdCBwCf/qGOfQ62rRDSmnIC
qayt1uzT1rVg/uf+raOKlcJgQ+DTrd3eGbzN+cQLQS2pKnlb1yPAzDnqzl4emMjXB6TmZf5tlWDh
lV9GW136Cmjzu8Z56V9gjRwMAxZERrlneB0lxVSRVKyRwHWa6q680/IudWF3zeefmC9nyWua02ha
MNKdpiOrA6wg+fZlX6iDPhO/4g8K2DiKtsarXLR3JGO2RXPhya2M0n05Q5Hey9mSFN8S+jRzsQSn
db8ZTVJ/el7ZN0DXfOJR1zvlwzRplGXV0pdCaeq1Cx8DPdFPMt7JsFWc+ktrO6mDk8ChoQjNnlJG
mXfuoKdbZu2iJ2sy28kVVs+O9/QOS5p0yerj8UzEwxhaI5k1JmmJJXHls2Y/2pSD/cc6SrqQffXX
Aluqf/BzxVTRkZ8e6oqNr/VW07wNAX5SSaOatkC8zoeaQaXeJVzVXaFY/0yBx3zFzgJOeJENVmCB
TbUdMjsLfaDiSyWhG0oneUO5NORyBjRrb4RlrFow00IhFPV9fR7U6Z29lG/bBy3ojzFMEjXcOcZv
AjEg6oLEgo1Gh7cET4vDTs9bnPbcNDC69YFVKVpcLF9zxPTB2nARXlgUy1p4YL3yDv453tLK1hD0
KLKSV3GpAjXy9Fl6whZZMa9UZPmNxABLUuqwdfDBLP1I9xPAohotj31UcyyKkjbrtqhQHnxgYFTM
Y3pW9EPwACxBqD8AJ5Yq68WfgdeHqmlo6Mt5L4A7zVVTcYq0+qZBmqQvaCA94+vBcmLdgT7SMsYI
Mf+VOUH7v/H/5rXOxdD+vnQBnCZD0tEl2y0+s1IOKSxTe1HPJY9oK2AvhjneB9G0RQa229kqr6nf
WK9cDcc0r0OvfoIjWi7NS/JYTUIWwPBwP/tA/s/9ODpFEd35pnQFlc5mEh65N8zo6QRV7DIepWhA
qu+2rdJmMfSyTExD4sWu8rnPubt134JyvCCU7+sZeWwKZBQTF/65KHTefGxGE5c07m+sYV62e9KP
5j/Jd4PV4AWXHXXzzVUIGderZOyOy5uNOvQltF7bwOy4MrFxrjO+8JxxoBkMP+4ImtW+c/WTHlNN
cO0ulDilZZ/DN5obt7M5IU5fUX2Jfe/2AA7dXwpO2Vyv6nyn1vDeuYgWsnYIwcLvMa5oAr2n6o1e
Y1o3X2NuoYDLD7g2rKAtHkCECEikyHWZgZFolQTyG+IHXUAk19SmI8UYKZshxF8kTzcMS/bdKAOd
bWmB0CPMH5k+12FTJyy2oFQmvYGs/tY2H2dWlMLgLMylSXKVM2zRlr/E9Y1rNnn5SA5wdoq+aarI
VMbOq8tLTobQFpgeJ73YV1ESXeqIJzkDXlbBQ1emdRz5m3UCEzFCoiamEgPg0dyRiNqpgOlx22ON
j1QvvG77t5jTZfW2DBu2Re9OwPQE+DRTMWmUN1as3UDRGHygdWJtdnA+6gv5ZAkzJFB49i2VsLx2
Mr1qS8op2FriMCKjKyp4+yrv55tGSz7e6uJ9LzcoDC9zsmH2BFJs5e3QDqS+5MxSiWn3vwagVm0Z
Vq/tW//BYwTfkRM+FovB9aSGvBAY5Byf341/koHt7MRmZ2SXJ2uXF3YmHCDQ8MhiBlDtxRHa/VJ/
2Tyw8b55zM4966+iCOgw5akztJ8cVx4SGxVfn67KR2MvGRJFWNcm7dHaE2WMNtts4KaZqMH6C4BB
4k0vzKK/pyYy+xsTCVtEEkRupVhtRnUqXHdLcGKET4PIVn6UDYUMn9BYO+o3A9GjBeHx+txz70em
e+R61EsOHGESXz5suRqBmj9EKosn4oKqb+d3QJ1OY52YTZP5lqexkEb1XBnGrDEatEBy6XXpigUf
wSmcClR9bjkgiWXdy5XRvw7cvT4fM/etAQVWKM8gOfhrwJGH4j3/fxl/Qzk8UUTOYA4/LXUqHIzc
dohp2CK+vv3EeDxa6jIljkv4HvbutNv+Q6uqVJyOsO0LIEyQki6nKE4Nu9LnDGsHxFAnUYZQVd+g
8fUpsMXEjM7t4knJ7fkDSYVRYZGmfxlUzjMq/6VZ1whoASSDDCk1F3Omsw80BxUiOOZ4lRNXgNlV
OsCo9ADqSmIu0TKWj7JrFsvvSVUr2GQP5ap1OD1npqHfAEC11Cd+3SzMU+UNd/tPoZYiCfogxD0D
W2xp3VInfJhWONGWb/5v+AugSca8P5AiPAn90IFojOEAKqThet6aH8U4D+LvLIyrEvZkzGIVWr39
XBT1cPUR04F148llfs1oalCYa79M8x8W+tL24ljKvsuDANGPMER9WsRmCM7Con9SZm8yKEaXlaCG
S5L2f5HFQy2NhsgtFbhbLIpuv9Y8T1dHO3zy4Lt2Pg97TYKchRbCI7/Wc553fXxwywYigMYjxiAH
aiyuyEvINgfqTYsnCvq/F5JIkvXF4/kJWG8QpimbctC15nNXzCpLqsA5Ng7EhV9p/zxS2ztKJ8tk
aDuy6CCS28UU9mQSB9HkHJSSUVyPFUdOjvZ4D+z268xn2EKs3dHVIk6oTveOcJzcFAbpSg3Kzma+
Ystdxm9/lzna+vW2Dfx/C2LOxFTgADYqWzPT0VEicXNCMty44G4VFPm4xDSXSukaBG6/TLBPLBw3
lmRlkJXliMmtOvuRrrwYUVvIculLsRyoFtx6+NIrUZigsBwE6MhnDwCKd/qgRYVodp6GSf25WKT2
oLX1+4lfn6c+W/nK9Kp255ciH4tIXySmroVIcLKhfWiTC3NEXu3mNAQ1BuZZbyIcOmiUVLdxUgXC
LYbwm12u8BwWRWP4vHf561qvQ631LdEIzPD6hROvwOKf+aLOXZJf5AQJQDim0dzow1EuktMfg+UM
+nUWEvtK1BdpwTsORpI9pz+baeI2p5TICnXpw7ve16YsIunOXjeSUEX834VUUM52ivu58W/cW+tG
0gmKL0YJ0C68DEVbh6FIU+FOVJJqsJGDL6m5XNeQ87wqWaRiPkDlyDx5mDo5M0zhpBryEK4LXf10
loMF9U7szWIu/tSYpCNfjXOJoAmlEfvJnuJ0sU/TSGlnls32YITZ0TKQsXt3HCZdW8/jsIoROEor
nwQlVFrKQkhN2XT9pILCLdyzWRXXq1tuylJkXmjieAJpMZ2g20Yi0tVQHX4MA6uuxNnB/yUsHPYO
Kicuz2m9OxlVQHuVxpX1O80W4bIXweN2+H0WjKlxymgOYyHhYhRCVBBtLk5kZqcTjQpHVCh7AUCw
E3fhRWrb36VOGd+7lbA5X5+IDBptrNsJGXUlv5lWKO3GG9cq6QXa0xzk47qrxU5HPJsaCDehQ0qj
CpCUK56vcZkhT3SXsCn810+r3NudYo2hTqVye9XdYnbgTkfJ03q/be/JDELfJ54TYvN9MLandnF0
1od+QWa0HYkKKGDCZdky0AGld16m81WFEBVh39kCXnGWLoQWZsXCwIRS8O8XtyU/HvPZWDCaE/tn
/nvo/GbyMBg514QRBQ5/vP3YPEjdpPTp0N52qsrTAIm8pKibyMGuOfSKF1h3QBhMLneVE3kuGtFb
xRTu+qkUQxOB9FyfcC0RSHBpiT07L3+lJPnGF0uwtwaKCfeXHu5Nr5tGqBZGYzSmKIkF37xIPe5y
JzWSYCuljB1dv/lFipS66jFKKuUIqGZ0cYeaNz/4bQ2X9qbBrcUObRy7XqGZDlLPoBdopL/ncnDT
5VMgbba5mLLo6LM5d7mTNteqpwjuDIaEl+OC2gDawJOwqFxRbIbG6iuABQ5/AORk3MW8y2oE+6mb
TNm/wkBmmIvHkm9tBUmFVEowTUiOqsMyfUxoELSE/Ch9YexDc3qnBltNZ2MAqSM8wZjttqIZqAjX
+2rs0wmHewTkcoxJup79+K2rJISmNVENUQX5VljmUd0XVNWDzqa+pujU9pR9zvPWeg1Kpr/AhDPy
QQ5EH9vqPKQqapNCIlMsygXQS9IYNwlZlnCTQvwDA9BFyTtdTCdLvMkWSrgBMBz26/s29EU8+dHj
BsR3UFpZHOa1+xBQwaeVRhtM8Plspv2qGnZlPZcElHs6TgSp1lnb4lrjf2xCZmBmGEEgnVXEVd0S
aJL+msmkQ2jLRz4lRWFRWApgVOC+T0p/BukRYuxKLips3g8sJGWbWo+NwT/fs6jN+5nKxmPwKuLH
Al9U8hZ/QAE5UZA7qkEAbWQdRE3h9aUtxarN2k+l0V40iDtPAllyZF8zowiQ0DUUlEaSdL/uHQl1
G1aBT5DgLgD6R97pXU4juwc2ME+MySn+RJAkpWqsie1JpRKU2Xscn6NkKSQkUClNViXac5uNNcPV
N8uXD+LiMcsLUmiSJxUxcUKnq/D7uvGp+tCUJnZboOr8+ibSzkuoGyWdOUjMvf4ANJRhPUcd6rNO
k14PzIHXiWOCl8WAzstRW2c+SwMvtskYpWbmsFBeczTAB4upQ52j6VKEF6pPlA0IWxP3Vt6CWnxx
wTx6NxtDojDpUUfRd7qFiN+WJTFKfZOFXRRf35/cWijL1U9sKKyPEVY1F+sB2AbiFRDUsPcr53PA
dn6cHoNCLxZxhTjoz1vlSwhlnR8QhPDyKqQpR/e94fKIJ7FJNqgoEQvpLYgRf6VEwtR3C3dq+yrA
n4Fsh24Z63BQIui4IYJWGJo6vJ3UAM5xiFXPbJboI+qPTdAwI4IVojz1/rmjq43Wxo52jj9JPmcM
kib/vGYSMwYPZgfdFk0Uy8kMqCk167ZyDvwA6gNsaX+8zHQRv3yv2/+8vjVs2yd6x5gfISrX30aC
QAxtboI2ShJo9zQCiOeiX1xqwDzCCJL6wdPPk4YGpsgBqZx+FbvDlA2gvkU0LzKlYCXkiJakShrd
fRGz4Kef0dmXN3t2kbkm0FGXawwZyM6Gd9eb37Zem9xOAuA+x2QrKR2xGTCpEFUSz0Y2tDWsGudC
m+p20FsG7rQqn7v+aDXoIiMA9KcssvOgdg/JYerCkfLz7oudFHGW94iSYWTLHcemi+IWkCYg/Fxy
N73Q2Y3QJcPVabmbTyKxb0V7R0tfQ1qZdhqw/YleRlqywFLbwBnEGG35azQ4hS+OiYX7xpwTAke2
gRCBxpsBd/RFWaOeiOGhsR7mvC6V03MnDtfySfNygY721nNPqmVN8RVtl5Mcc9gBuNsbCj6px8F0
r18Y3zOSRgiKpPM9HVaogiwgTWqnV7OPP4OKoQKRKtgP6/hmIuuASvwMni2YrOC+3AOyk8U42O9L
lA9AXi9/aP8mOO+5p++kSyR5OhKFZKWREGK5v6aPPnFxlYrqrhhh068InrOXZNSwh7irQ+/UU+jZ
nY/rLWFniqM7tW6tdU5ae/MZ0nmCfTe5fQHFw95oPpneIAQNcF33E4ydIFOoCa+L2QUzk5buciJ3
zlwdhyThfe7oeu3ZfQxm75gPDC0segiUGIvNsZf7qApLNAbrCo19vpbSIpHSvvet2sMfUii0BiK1
2bzOlY7peqn2tGkHSpf2vf29oTrB3zc08PIe0sC0H6LSEk5NWNDMSUR5CVSwq6kKpEqqcs2K7E1e
V9RuFPdwPMs0mkXxdSmF6prhqQd/ppcuye2MXJcTnAYVmAbjpQP1EUWNFSF/IHsvpRuNG6gpvVHy
STNfM7i74HX4ZCtfJHKnYUQGDbFZwqcrjM0XFI5S2UlSNB8d+3gV8+oxnqWExZPGZTXSiDSeSWRW
4JtJ8owxLzqa7gkILCxZSWe9eaCBg0pwvoxUpZ1qzexo6tXu0n8T70tyJQebUp8fg4WA3HY3ra12
/v7k4FHOUvi6T1ozuTgSpblOLF7kqlZh/41XPKsX6X4eow+8bcEH2LbvgQXY13WGXNSjlCXFqcaq
0HR96YLCTE+WSoxOFJyzmtbfmlvBZ2ljrNZfXYB23xvc4PXxN3r3Zmo8eGPybVA2QUg2R0P6SDmM
Gz6VnwgN/ur54VXCTluuqQyH/t0RyEthb6Y9VmN4/N6kBXIDEAkhFT8z2Qfz/g4ARdXofNzM+aqL
a6Hfil7L+n/oROJ9HP4rs1HPnlASoS2U12atjIyh+AhfHRzJbs5eH7JbvP9M+Gwt5aDgAxEjnT9g
HzoIqm8u00/3H6AHoQrgLH0tSrO2HhwU2DSXtNG55zFWdu1rKTptdO3TN7NeH08LvXhmJplWaHLJ
afpI/27le3SJm1/uAop/D18tBpSKB1O5Q0yPDdLZawue3QQzdNuuzPRaYneGOJpTV9Wglwiw27pp
dg9q/fXe4k+jfdlZQRghJZbfcM1D+CdQv28aDVK7Kjd2Q5Ty05f9EcgtYYUzdBLSIGmU+GrZiZAn
ZuB+SA5bKbaJ3cj3llle7jO+xLL6wAwulTij8YnZj99z73MS1d7T/QO5LhSn4/kN29KAZwFCRgAE
cCmsOdhJVp2qu7TxT480OvOtx7Gme/WNJNinp45ttbqUiKXDiR8DxXPiSMVERnqLbmbLxC+QrmsH
2nK/LrpCRaPFef/AGQGIBnURdaLWDOikE4DF0gHt90di0f8w3Ym6sCjp5gtTCy5a80Uy0LdSgOgZ
6u2EFNTs72KhsP3u52BrLeUtmmO2YWdBsDxlpopN6CM8iwKw2p/sq5TQs8Fy2/7x4SMDT/9eTQCN
ZsD3HTRQLCv6FHBMGl5IiQbjYxjr7PEa5zzmysD+g7NwjI+CR+q5g0AVoadUl8K8VhIOxTBhp7Zf
YcZBXKlXAFr8xI7GwOaS6CkMH7K437iJnJo2QeuHQY1aPWduVXET7bC2yCAEHKUE/rAbijTkFrRt
Eggwwd9E4FVi8SSnbaiFLvwXt8uk6lohaodr9CUMKXJ1lns3gaCOZmEwnHbo58OJn+FyqxxK+2BS
woGUZXNQQKF4TrasPhSHgNNF9TQZyaiKTFYs3yikX2u21arvR/YrPLxG+VFLTx5fAgN1cCadf4qb
s1BpgDrnrTQe0XSCL7V2PsP431n7jxoG9KUciiQ5w2MC55EUPBgHHG6irmq2vOKDt/93a+GKb8Mo
Az2HWNywfWSMkVl+bpVsu2yio5lnE8NCts+rgdzqlXEnlEX1keKvxfCDTAqbkmV6lwDQGeCuo9K4
IJaPM0JFbgwy/dKDk4z8Oe8uClLwt8daUHwIVRXIGxse2VZp8Gx0qayxOjlG38EGW/YxdNyXI479
z1aD95LLWRXI8r0EK3VT/zRalKa5mBMx1Ggu2GvoehS9MFzSjr3VRwQOtWN+ahVjbjQeK4xHfjnH
KV0v6G4w3iPqFMGfkYkx/5zPmRxikIWn0HHEvfAatiGVBOkHojoxPZIRUkG5lrPp0IfYHFo7znHt
9TpAbhSnHRAxF0X7EQQA83X+kUd6hUFp9auD9HRtY+aFMrfwHoQuwSjQX+/JHc4yZN5656eDPdGW
91kZQX3JENy21J3Sbzj7YxQLwTiwD/QWHBcUwTylA00XPtWMh4JF0DQQhnMfqJsDOnhicQAC4tHp
FO9jg9EqHYf2uR1AI+sObdQtdNS8HMigwc4gLdo66bkzpjgCETPAGhooOMHer2qyd2F13H/1nDzj
ZPixTM12YjduITNe/UGivO0BqjIeIt6NdeFTBv0FVwlrDm1KLPHD7CRuSd9mKrbyPiqdYLmYY8Gt
cnM7PQOUpQXDttHlLXW8NLDRIkShvB2rCzdXCRJpRu6MySaVdJ2Ndmii63z6VCnAZipj/+edyIuR
HXJNK4I2SWp4su40neIFk7oiti5jcg+3psUkHRR6lrULevR6c8DLSPMFcHv13f8ESvomiJclKYId
GUomX0O73Xpjw4LdPUSH30qiE82g9FLytljZoCvAQHAeTchm2XyATqkEwr751EG63zvjRc5rRdrk
6vzrFvSWRkYkhmQ4WRHe6wJ7n5EXNeq9WtouJrjddsWcOj26v134i2UP/ipTvLkOMj3W+pcqiHN4
6ab8inO2b62tiiNzo5S+f7uquia3wHe0l37jmOVyhPsUXHcS+D2EXH/HsjQpJteJrEfOAvJu4GGS
OJ7j3oQz9lrZAAx9dfdnggMckBePBSmR6+fWiPE60GYM8qTui5WJknhZAa37FPA1b9Cz/+tmNNOl
+DrEyLc04Q0BQEklvsvd66JZ8QF6fSSggn6gGIlDYi6FgixXQeqnaqtEL/baJoYWuqEECgaqxw3u
Z5riD+JftKb8EG/6y4JoOxryTKqCF4QN7/0yrjz5zOyoqe8KQKkqPR1FYucJ1FXCpBBDE1rsUqGT
4ahZD0fzjrlTaiBAXEhroA3KLfa1tmS+vCDjniyxtgabf3PZd6gg5XJhmd+L1kVA2eSmgAcUJVpq
Kq3GJfZEDHpa6d3F7NoE9HxrL3ceb1F+rtklVCa4ZlJBF13QjTRbQnVSlxE0mhTUhGMwZ0N57DrY
eM6fTRz4wIokXITuZwqdikuFib9TVvqWDEHnY00BwuJbDP9JL1ol6+vcznt9uV66UkkffJ93us0r
2xIuxVeXXGL71NwectKrvG9KS4eZnQot79DLmHKcTTGbW2EerZz8Nv9JVcmqy+Im8WcnF5Em5gKd
riBwmSB8f4PcsZ/Xm6j2dVhhGNjzSOJhbXopVxPh1KHRMttdPKmPWDYaZPg5Rbv7A61YoTzIW1qh
W+xhU6uTvQ4s7Izragv8QVWqhTplRHYf4sd+9DBtDCyi9UeCR2ktB4imdplHDzg34RC0iq7iAnD+
OdFCYrVnf2u7BVBLoaOvxpN/zkK+3MkbajDlFzQxW7zXfQk1F9NqrTeuv5BwzpHNVz+U1XLxpxBJ
59PthRF2dGu4IJyF8WZvFIEgpedIU/du2YWCsQMyu32XOpBaDTaAXHkY13rpOQc4wyk6GtNznXg4
kTItlmlKTMHRWwCSkj0vbs3zbc20YXKfMDAmeB4pkECF20I0+7ilDm4ysz9x3MY3EgiHGNs5PmOY
p2VyiCkIfxX3Ra9XDvZSzKHAzfMaGy6QSh7KRBmcbaUQfthjhz0uNs92j8AegrGcJ1pNWOfW3fm3
rmKJN5c86PQ6eWH6Qh4NHz+RzGRGXWqc3UeOr+dLJwyB9BRuFShe+Wg+Kgg58klTN7Fu/fvYahVg
Yl/byQgVl7aEzGd5/ilmxuIlTdQbD4ZsIBhrPZDVz+Jww5im6bbRajcxw00zdb3gr9BX7GBcix2D
4hINA4cLu3Xs3U4E0Mb7J/fcrgSgzsvLJXR6TYZe17CGdXJY1qRqFgaXmWpA5f0hUTyXhU8Pe/J3
WADI+Xq7TzuKDJikku580sxk9UjkOxrxxnamThbUYioXJYxPImh84PsJrzPFsJYMe51kkHEkRhsr
cJXGKlKZD1RsJITs2uCAFqmKIBGRxYYw9vehDt4EbnqoUNksZEJsgaWG4re3OwbG2298Zwnnn3jI
zNVhDH+97UNwvxIbJmq4uU31yFMwrXOSCA63Ks1X4d50W1Qqx1qwx1DlXFmdurpLBJ7oXMVQ/qh5
CHhw6Oj5lD2AeLuYrbjuXMbjSEp/ru5K/uRP6q8GhpjP72eT0Fm4l1DeoHKyLwY7FwnHrHOCxX/S
4w9rnia9c0rxzuu0vHk13NOC8c02N2NLYRBihAM0nuk6uF0bmVo9ieRCeLvniSzi00/IVC9LWBva
auAXXd4BV7T/UGp7GxiX4chJuwqn00h8rPEbDeR2bTpBQkeFCEDS3fFGhW8tlCKs57OQ4zBQE9FB
Z0/kQCqrwdmr2PWS3rgaP6Dmw54Fv/oHJftVXESxuD2IREPPUhKsbUojxMfMscurJN9hIFajw8Hq
eXUnLuUEtvoVIxceC+6Q236XwG/+xn5qZCFaan1uC/aTh2Q/8skq5PBRcRjw3DMpa2RnfMzLIPcc
TgQSWn5mC8nFWjIR4QtKHTx6i9GlvoXx1QR9M2L0T0KlpsX96Tuo5i5hn5vEXEk7mdsqJob7BM/a
EsdJ/w0TiQgWzZUMIuVcY4iWxdCpR5pZ+9vzaTwFM4kKfchiYVopFzzX+9c9GmoHUkeL3y+jUo/c
4K6YnUDtJQh1GXEaKgsUMEUOhTFvt0wciJssQL1X1LQhhVG09q46sqXrkYa2houtS+lUQ574yOVq
uOuWcAk8/s7bIqOqXZ1dc3jRTzqXX4COemcWKjY3GzIEWb96q/sIGmiRDKV41akxE+S3hBybuUmi
EJky5mDzCLK7AKOlZugTDG1Ep8MuNrCTFShps/4Qe1TeOFm4xHhhH+M8I4YI1mZkpavgSAFJfhHF
2kdG4UvDc9tmNNgsxbrBDtTziI9CvSGr8WrNLNZ1wyodKDw85Sk9/hsWvvU6l8wbXJmq6n6RQDN8
ttT7TpoEmMxD+E8IUX4PyuDzGR++0jlez+2PfXA7x3HB5LCs68aQmMgtszYUKxRfrqlHVRhzeMyI
yotrwIcb33cTdZT3Skg8/S6xd7YxBsUPMBHJRDXy6RYPLLwQ3cO17FeIej9IIFOxxaXti8DjGBI5
Uh+bmzLku6b7rR6wB3nt1zIFlLldbCY9O3PWNb0FRhJIxr2BpeGrjBzUTrkcPMh1urp4MsiFYEZ6
XXp8ZnI56fWEpRtcR0cUHZM6Lvm5UzBRDHP0QivtvQSDj3BlQyK/x1OTu0EwAMbpvjTgk8S9/Pzu
/UZKE2H+gsuJtpqbEUq97OpjD6fbM8fHmI0QHK7zS4UGIXixaTvaXMntGZNrSf7uH4WBnWjR1bn/
J4Yl8q7juHY0ETbZFEfTO8aGUs42AvIhmtbC5wVVVEjeSXW58OIRORPyrHiI1flqjL013C11Q6oQ
Wk9TUlwPbMUPdQVHW388fHybyxizM5qJyNYkncr2GOti54+Cwh9+PlKXzssVsfHXDivs1BsNeTJI
PdfkXl8jgBtrvMjTbibnDneW33tC9rJQqVgByxDpP1uvyTW4dljv/3Xas6J4vDhf74Rb4Q32BTKn
+04csxWwi1/qEj6JTJuivO5jL8Tu6Uv24lrQNzrimDfJr6BSngpa56np5HhRd2Vq9yTbUuZY8Rfl
NOsAGnJwH3A3fRUL4cvWPgVhf9NEmh1iLHt+0CdOO0PzaiFo+w3HeLuZJNwiW2diQRBwj2TR8t+k
gId6Un/RIlGLpfbdF2OVnZHxp/wx6iMNSirUlStA6QjOoV6kwn4v8KiqBoWK6NdQWxSReFLSY/O6
Yo+9XushZci5aPuUAIUOP7rpjHSuQGuWHk2YHxkVjt1SLwj/tMCTNjNEc8Q8o7ETJQaYsZ0yqgo3
ECfdw47igY8jK1lb00DdhcjmSZ0b6/iqmwhBOxq/X+SPcF3qxhVZbRobOkl/Hlw77WmtNh8zE+Qg
P+YdizYttgUoLDQrv+M/cQ0aVAxiLl6jXAuRgzGoklHPN8fe8RaQagq7k7jGD4zsCpbOOerysDIq
756TMdOCfQQltHY7c7g/pCOj6h1VEfOliAOLsJC8kWW4flUDITGB34aRupHq9HS6vjIGmM2O5hO3
0HhQOdOzpAkdlhe0LFcR4NJavpdIYUSbBjPGWcdFSvj3trUpSiNZMjYRyNF6VuK0MdIGZoMnV57V
f+wQcSQKzsczOPbJbtCCZTfC0ADkAwDqHoiTgsXniWcZUe82OSMd+/PrsoKcW6RHVD6s+f7mtlEB
7JW5PoCuRv8tYr+cH8ul6witYyr49d5U2phWr79JAoYFEsHDxHOMgTkbEDHoaukLGEwwd4NfwERa
hjcPvSsYNTSl0JqwQ36tbnerwa05AgnlO0cVTmOLIuvS14Mzm3n6iigR3f+9ofVqa9f5E6ZZti8a
3szWoxs+qk0lnA3lemYKBGbJlHeMVYobKP6GsuBlpXAOzkSisxmBeZxV3dw6hl4NAYMaH82YLgVC
vRcQipheXfWbxszAKM7X/ibXqX2vyl6UqLFLSx305U3INvRpJMV4Rv0aKncFcSwO4gRAMMrIXMBq
dd3MuK8oWqg+iO6usxrq+3Sr7ARABVE7iWLujV0e43juiixbBHmGqNyjCPyBhELLqn9jHF74AE2F
Z2Z8ndZw5eNX4Ix9r56+qBqTlITWbXSjVShnqKCpBiXlpvP8H4/xedh8Fjg2buNsUuM1CoERxSqm
So0kumBcmDtSlnj30ouwfcXRCNSHFBgk7tQz0DeO2KZJg0DsZ003vTohjkfL9Ay0uWLTlcBf1/Wp
oJ+97Tg7U1irTSMeGJurSSh933bTLTp5+Htgb2DvHSJOK0ceeSsjxUVopkYHkBzE/KXRDMokPI+B
tF93rxfQu6D1OfaelGRth3ZiqkAmV/rJxYbt19ncnJnPp2Rvr97GQ34IY2gwvG4bFghkjfrHZfNn
AuoNkQuvGpNW5XBJlvb4fRkPKFofaW7Aevt5qB25BA7ozHdQ7P67xz6AcVbHQXMtrABRrlIT9FWX
o1wMPUY6tnxVT4+OqbDSL03wJ9tJ4OCYglJV36IMGqSwW3Bae4k34MGWPd0Atf8/B9aD/J1XKmfA
e3nHIJ76786O9dhqo3Sfcr6P5R8Ya27r9lTIv5xS88V8T73e6x740bA7HuPJFwfxh0YbXAbTIdcO
Nwkhhlntg2N6W2ES6kchOBhS9GSX8/CpIPHFt9YU9wLRPx+InGTq1wI0HHIkG2bGH0qNrcpTjgv9
Vs1Gpm0ZPM6AL2mAo4MJTzDJ8hyQlzus5xzbew852NrDUO46t7/naqEZkucWUhHBe+E5xhWD2vqr
R56TYncidzh6UkF5b1qFDkXUZ77Cg0oHeA/6jJ43hXsu5kDQQTuOQT0GYubhM75GBlf/EXvuw2r8
iIVPrEwaYRdNWW79sQqpDcJ2HTo+sxheRZmUL7PHswB//afCo0jF6x3P7K/+I7xxJ9BRPaaPHGKP
Vr8cupUkVcpSJXkJUwhzZhSb+h0nEv7phVAfPWiM3n8vkJeYkDKQVcMovDfYm5KgWV7znky6U/Fn
Orh89y+FIxW9OxYJ9/6ekjaKPxl2KDhkYa9P2S+YMMbfqX6lLUWW6KwY7BJXiXjQfbY4WyhsVBJT
5iyCspwR8Gq8tok+yfXDTLFJXOUDXNM4GUrqW1MQkYLmYosBqiDv7V43vJ6Kad8He1O5X5x7gtvJ
K9Etbb+htgruXJABzm0x+VQJLfQ0rnjcv6dnL+KuFQXU9hzuHNZHtX+cvQQhoM648rdYvaEKYatU
XOTiK6JOXM/SMUJn5wWdOMWWCM+UfQpeZNvSc91yaD5GGmIu0D58p3PN7/Xb+EYSxTYBLqkkdBEx
5Iedq9raZjX413s5ErZArk9MdxPMtSx/7Mxknc7xLh2KUFyQM4VxNW3wejtlYLT9EOhq+Lwt9nK/
tNcAPAq/OXHxg9iXAprM3MOgBLvhU0+cbIKR4jLq4W4UcDsqc9AJeLLWxmgl4DaMufRRY3bflkhE
+7DPY2svywcy4fqA90n+F2dmGHiwMroYlR63pwNauxxUZLCzPAnH4J2OrEmybKVa5//XHyVyG+UM
TvC6v4Zq1roS2StGG+hq0wVOvnZjm7mqNrl1D12eBG6jyvfatZi2YxbaQQMC+5Xke9aC/rtMUDIw
Fl+Q5nv7KVrI4h1c5y105Rmrnp1Hc2l0KsgdIiHrWhNZ9lSrILEIr0dmt/2P7v2xLOF7HeOPfdRi
cAWKz/cpq821P30gCYH3RqqhAPO/2Nk/BMXNVLjI/KhLIeMCOd0twiX2Ux4TbVhZt+Ilu8FEJA+B
rykvqIgPj0TUWtzFBGimMypDGwN9LEGRjMohIxRMLSyRDRfYLqawiPjp9FCUDBLvY07t7SaNNhFY
F2XJWOARp/ihdl/+q/TyKE2+A9F7D/GwJvgelabnQ9PU/ogdODKP2+icf02azOFOMnBh2SNb4nok
H3teMsNzDVfDm4lwZ5r/bqDLtPFWZxa1aTSah88QHTe+QAz5WC8oeMHvSaZx7DHQ5JYDHoF0sYJK
ryjL6aXbtGBNmW2cilXY1IUc1StxFaA+1bcqKkiJ+UZa7UC85mmmMx65iQQp+GK8G+e+ORnnogPm
BWK9ctLQ7hdBm6I+3lDHAZOaLrvflbSUewC3exEVmoYa3Ba/LW/1spXZwa1dH5mpdK1wsNtq3Be/
WoEXfIcZyuimdKK3zBwgZXKXaI/FFJbKCkB07WaOPpUKBB9YLvBdFxsogASyOS6dpVpFY0pEqYhM
9PuzYJn3KatsUyHof+PSbGrSwC/xHy5PsNyweTuBp6bYpuimN0s9ih518xz1u0YVKwHfB1cAjLZX
vjFoZUqAUcWix13M7sFaIcpaNyfKHXFY3Qn0sAmNL0lvdxo0dSVj/G+fCXDaVC4mv6LlvK4TlPHT
lS8ocdQp592TMs9VKnbUv0tCcd8vq5xm2p3LkUb4xzeP8TvKl5FSrksw/CWhQfXn4Lsr0aXg1Ltc
lTG1VUQTKCaKP3NEoTgnj+Io4ZyAbvBLcUrd8plYXPHCeMMtYRd0vIoI9rlq2SX2ZZRAC9VLa8Zw
10A1hmc/GMZndy4FqC/PPWNtUax8Y3vDths7EHURbEpYTrf35H7F8T47WII+AOsxYSk/qB2y+3PK
DKgdv0kYY1IR1aKVlp/hibimxAkUyVWMp+AWXuiJ/nkjMYJjjS52pX1NCiDwPTFuGExiGWw2k2x8
rym1Naw9NH+4szhfL279+tH5VKARsYoB3utOqbnDbV11KmVmIDVoT3V2suBpjOyr8JgRAYMNXbkO
q/CRPj2kNwleq46K5xW5gZH4z5f5bCqiJpIUNWwALKNz69oy9CFfvxav1bf65lqf8iiNQLiMqFbq
WAZ21aHmPWZ1FWcDL+hFAmmJVa2Nh25LgKNeK7tHyZ2cRHpz7xE0APLgKRY3qvcyVx0GDgb5FFjy
bTLlyNYAkS++iFU7zhG7CJhazW1qtKUgcaTRDpRAcptDEnJ6TXJJE3Slog55mAV11ceth+p1GB5+
DDHc0PlA+iIqfIoOD0IghaFJLakas66e4U2NryEEyFHH3gqvaKwX3UEd1ekBNAMcfD5+wjZBEBFS
TDo7nlIq5fZZzU1/eyvAWVOZk/QQJnUnuUXm2xBy3pesbFncSdi2QO11qjFjdT170SM5AAepq6lj
leGloRlPfAn/LUVjrKtXzPmb94NQU8/hvvRJeNK7aIX3n6vTDcHj14eoFEy63k+CQNFFWdT0kWHq
OJYvibYdDOFrzVOxIQzDarwrqtk4xovp/jXbPlIp1VIvoTWkyGQDZ+9M43XeUSlsMs5RrvDO2nVQ
9vgJeyMVSHRb/kzQovfuG2Im+2e6n4nh55UBf0Kp8hEB8AmlxP22UOlOJNUYVh3rYiRzlH1jCMMJ
TCBQbD9Ly7UcgEVy0CU1aFAPtjX6uJg0kcUQzR3wBCtfjSWuKX9faFTcPU6R5nG+nZTRQy6t9RPz
7UCf9mILR7llgNV+3E4BLIXtEORoMRyyUdbQWpWIG/LMTp/5eLOQ3wHY8ydOqkKMV5hdAs1S3OEj
NYTVvzjo81Wiffa0IDfLSLZ+YS/NdobGtD3e77WUMky4cZ0p1OfFAF6lGtNVV7yJhaxko+on1IX4
tdbg902bKNQKkdm4RTsE9SsuiJ5mvHNHUnCepyUZ/NjiQbD7Idwvs98rWoebNammmbTllweVsWUI
yShF6pRHDxtjjlutDgX/YtDRzVTIjXSJ1Ot2ywJZqk8qfhxaqfWl0xmR+itKU/wdp9IWnzrmrh7W
fj2LMSKpG2twP7DRRU2ej651Fxagg55xzWA0Y8l+LRdqruxv95fXS15uNpsGvAgkbqtQE1A6jPZN
Ep/fs7SJZAfD8KjWFtL5gv8yg6H6tCWVElH35wMjANvjB6XYC2W/Z/v9Te/gF55xUCDuQcBeuNfa
DSnnWvopBcYkQs2nR6yXE+XtKrXXy9BGa2y8AkOaxY9+asD81wYddemGie5X2B5ynXl3nkGTHiTo
Ex7Dx5EWsUM+RLbiYyb6a+yvThhYYVK3S6GhB9gy4L27h1uElXsTBwYtVD7d+bG8MjzGGBgw0hnj
gklnv6mO/DsSifkeru5LWDpTC2Vq5p0kwME6XvjNJfbM3Oc2JCpVMvAZOMDo++9GQFlOFDsS37O9
1cKI8p0E6lZwldqrf7DZ8xIbef4NTKmd3R27iDjQGpnKG/c8P3tAOxCa3bT0rdtg+w5vDmkWSWpQ
7p3F1mEFTvbMq19EENRvB59Q9If/SB7LncQI59/PNYGno9VohvrPqgA1SGpwoJH3u5lH7yRYDeoJ
ADMe/3Cu9i964q+2t6h28iPXQyDdE7BSm+fnJKD9o8Q1c3QHN7rgwYZfenxA7iGxQJPh7C8NBrTB
Tts7cDE5gVqt8q+gFgk6+sy/Btf8X9MWFdGFPHi8/ACkF9bI3iUV8HYlAZkZYjt2JKI6KsJmZt29
FAwSU2/LUYx9kujpENLXygGtZRXELqJ6WIjs7eOvt28EyXl8b100WvifrsBNQLsGhnTqStdqvM/c
/KoACFSy1Xm2TwBqBl1UlFK5tbaFdAD19IVVWM0byuyAgmGu6K63YROBe2QxzBA0a0WHA9oRJgBv
2Mix8jtiUG3DiWI0ODWVyMYAtF3jt7tytwlfS/vpTyZZUARzTl4iSUbZZ0E9Y6yDvcyk2a4HH2I/
/mpOjsSAhvYO87WdNsMxNWhysyYHJKxw14EDhF2XnOi4MHM9Rl5EqtZEn5I2DsfgwWqilAZuEBK7
AxV8yNKFLPbHxqminLUyC/5P+czzvAVQKOIIU+FDc8znfr6Ye3EL+t85QvzNk+i0JNS5KZqt1F9K
/DGJMU829zsdJwiNJ8sktqrvQwC96eAff5ovwuG3EaAAQnKWBmzsX/SJWZbNW/hEGEwiVdz4gzB7
uMkg12FsglLGOWCEXSNuyFc7X4YRcx0kCdyYuX4DhNvUCZK1Nj6fuJJVCkYHpIKXPhFQWSa68q3B
itkGkSPWrdN6wSh6SqRgaTmiqeKnPLdgPSYUDKEgnjljdPRjb7QJmJ5RL7RlnUGG3PDO5Oe9mL8X
VwbfroDJmAUV71ECwvjPJkrHRyIE9YBMOzaM7uMDVHqLHW8i9TAIlRO8n1xZiatpUl2HpiNuU9V5
ivJNMPl2XCc7S/6b+00MUYVwEpVh6jNx9Pn+TZzI3C8mqwP1UCeGIxk6XEOkrAU9lQwVzd6iJRXb
AIpYDDq/n+H72UTPS/XTS97eB2XyAR+IRvxRILhFNSRTFs4B8WYBWtKh97On4m+JZp1cv287gvCD
NEZ1Rh1GRhXgmaZ4RET7TNATcIFv8CWrKJJbKJr2uC61m4gIyHd6GQMqM/g+qM7ytt+mgHU4GxcZ
sZjrSR5vlGX3cGQ0CXQaR0zrVaNzt19R5cjOZbwHJTz8dD92T9sEkXOw3xIXITZknfL61hDOqKSm
82prpFRVlDSNICuVTd96Vb9Ov8O78FeaVz7rj4pHdQPiCCLYbUPNuaWBwwKp7h138FhlZg5t/ho7
qsdTaG99h64+q5uEoLFY0qg9cEEaJCLLI6CPT4OJjWScVp5+kHmtHAbNozB0vTPEwtMvp6A5hEtV
fqQL7YDCpOXatUKbVnELp/CGHvQNdlzJ880gaOemj4CcjSp9t8M/8pt4yRXi4mMMB/By13tzrHNm
RTnwNZx5FM6Ye0RD+rpJKDQx+gXBldRRWOQ0LYqmlTwABWPousAiPt4D7lpbKMc/oBvlmS5NWWa1
r9WIJsrvE3oM2iJkAJ9eu8KdkNHOsDHTxAEXL/2LASlKQ/NLQuEVZjPn59F4lQ9t0eZrVBaMfBBr
f9iZzgk4byZUoC4BMk2NsBLzH2ok3PqNOmFWClmv8QewbG0KbWrnQoT8zgE3aqMhSM/IIY6XkHZb
St1jRRTVJEt4IvEUNLMWkFo0Spay8/f2ANkKJ6eAVH4ifejEmMTTGy0SPqmRWhGFqTzFKqjXl/3O
ZCeJRRApA/j1Z7HGno0O1nmiIXVJ9avaXM+hLr5B8sYLeJOFqGQe5aNzT/p29mYZOY1jjQiSc4GG
p67eMNckzwUo+rASuz82MQQyyKsoCLxA/yNXiKoeN3EFB5RNyMCPYJSD4IUI4tIUIQqn/euQfpYr
s2zJzWP5V9ghCsEo+CGykpKGlFGeq/2WKvwpYMlEv9zDzLIPEa/wJaJN73ua1J9c7RjNUeYTNlYq
keuZSgJKBCDclKGkXF5wH+lgQ1NrkvJJgz4Cv4+qt64X7fbQKJhPz72ouL0c72ppiuSRgYmPE1Tc
nIJ8FrFYjjMlArEvJwS+zSFYj60JVopLUSbAumi2JClK0jTx0pCHBixw24rZSOkL+W6HL36/nnNz
/4XIcottvSCRXu2cPIc8Ww06OCovAgthaAo4l2NK9KwULxct5WL6mQtb6JXmQ4NIs14tTGqbD1OQ
C0vCEqEBn8gUYmPbNKy9pEAGZ7O/ENxpbdtiP8H6glRrrS1Id2uB/ikrF6UjncAtjKtAUBMX5vXu
RpTyeLzT3+tdN8EszGXBOXIiW+qhWL+8W4fa6EsuCkAJ8ZI/7a8dVxKtFKVIrj0UUrMJqaqCpRDG
VXYul6hbUK8Thh4c9X7elGP5rsZGwYeRjicdoyow1ECwwKXQPz24WIbVDT7kAhQT2Qf6N8xekjlG
1PoKe15yaq8XSCLuzCchY3KW5FcE0qmJ2gDh/f7aESKT4jStzLKUchhiaw7FrNsvU2QHYLN6VBNe
329pyghejQVD6kFcb0fDS5Z7TA6yjvv+VELGEb1O2qz2R9Jm+SSEQTKldxNJl+UGOwCbsGA/d+8d
H+9WKoFICiA9/7AEpzzuPlxW4KkgEXJnGqs0ISPszMi3uJV3m8DGLpf77/jtKh63AKRSysxV4t0/
Qf1chc5gaWk5ygWSF0f6Ron0HfgRwQwZADR6rjoD3CLS6KzhRE9Yt9BYc3R9HBsHqoU2G0gSe9DF
avSdXWBop29sVtSalS95bta9yvUcT2lSKXxQyZu3wcvkbCPc20V2Fyn4pvQQoXIAUUh151WrL4p5
0qXFHD91cL58trgYN1MIa9RKMiLuyCanir7YRkBrKv4qSN/9WGLrStT8KZfJxemB+I2D8XTA+2Sa
QkJUn7bZpgPraBQpgJnoP5FenG0hljCvH3GdElm36cb8T7F890/2jxHYv5ow4pIj26zZh0HEZrtV
mWdBWxHGRO/PUboKtKW1V37D8Rw6/642Kn0TWe9bCMyt4JVDYlcKCvb6fVvNieLb2B6nrCGzknp5
QhhRorK9/4I7QnxcYGaSvoqAntARA8INsHO4F4KtLTSTuCIJDL4TSb9h07FVQtXONZ3VPV/Z1k21
kw7alWFsumT4xjjuy//VWqY/1mkjriTs57KyNGYipDvDHUsD21KV8Ulv+UmIi1DHWZJxnleRv4g+
z1NXUaQ13RU/1ly0hnfvjDtKkE7dIzeQbXN9nWer8C6Wqh0WrHQU9yuZ0PQe1lcPR8zuB7wp0JJM
yHyaylMrrwK5dW7Kih3KOEgQ+SrC8KMxSh50oIjdYxriarLVcNSjtsTfNa8QVQwPFj2xMW+1JSco
Ku2VCOmhSQ2IaeNpHgtRYYy4yUWQVieoznKdPk1LfduzTAPw15DyQniutJYftiazamjU7vtCniBx
1WIOFGLyxZF3NtORZMWM901AgP/KXK/DyB8bCck7e1hiozJ95WFKr8AFnh+G+XRNhankUmSU/0DX
H1ctvaf9r2feHGEl2gQD4Xfs2ICQC3gFLd54hbctIHOynQGR6EWHbOpjbV7pkQ2RVvzkqL3cjxLM
gbdmgrIEupiA3KMCAVZElKdWdWnljhtUrkzQVBBwga6Dahl+SOsNoJUXKkbPxdwNqiiJ1q/3NhKo
2Uc+zaCg0rFvmm4ET4e7XgvAoWCxJ9y4Zy/n2gg7ag/v+5XFCxImdqJxZAtAhHjgo+wyO/F8IjEw
9fCcPebKlKZd35BFzuoX4Tlhmnwr28leyw36xKAu9nEBpFjFrH7DuSbZEC0khdrJVB2PEHQHp4zV
9HWK0EZN8R+uLp5WXxNSt8tNFwQYbCaOqZzqzrtLPSxFGXnINF9YhNZ9szWi7A9yHqq1P3uC8UKO
wYTxmSpebQ/gXSg8WIDU6jzWEmOPHCP4ybCV+gBmCxqUJywAqbOC6URTBCVBgKMo1gyUMWyHUrAJ
90Etsi3nxCERihM2j1BFi52oLX/vBouVM60lPkM5awZlfJKpR8ICAmpxbRRF+Kwgy74uZ5MdjPSm
nBJv5EnHciScXSX0EZ+39+8ZviaCiE0a1edZmANdG4+hEk1n8ABT/H7BIX0QYWRquq4fzwRW9nPK
inEU+5BeUaWhZiiznPGF7NDF+RQQBtyFvm+2Iq+fcTRMjIFxmPYtiaoejh+RjEs/EDfllBzFzLci
jVpFuPfUQKmLXwLlPtXTEeS1bLQhwwS2t8SZ2o3bacST84Sl/ZN+cwtMLZeb+XllgzxCb0fnCVi+
XHGaI9ssaaQJz3p1gukBaXIVKrBpMBG7o+JJcnSnLNzGqVnZYxmCAOF6egTwqYwDArVeUYqCabui
wi6g16qMCBm2UVAISVchaVO4Z1DWh+P1VATLBmVNTITwi/UwhlT02qVOD9S1kBjK27sfU+ftrSBO
bRm11/Z9QOL0RTfYNXqhFAz44nVIeE4IqJviljoq21PNxWMMJQw1cyzYOBCcrR3S4aKH64QFK8bo
J09iv3eDxCSJzf+tektoo+FI8mH+vwmdQyZDmpIJjMe3zrLQMmxD/5ZEZeu9SAFF9pl7cL4eX7+T
dCgggkFfKaJux+ITNpJVf5cosMi1BB8Gg8qGT55VyllMwdutxjDfHr29zt7GVATyoKvudZR3Wuyh
LyY7OXawdGnT6LRrAHFqJjuq4/Pj7n7vX9OnsD+WfMyrs2O/4wmmRHgHRopMPwaeswGbb3Rk7RoP
X4nQ8qBx02qXZKUXppJmb4mRyzy2yuR4UgAdWowveMkYFItmtVp9X0P1sNqQmZ1F3KzK27U0gN2I
CCGgcgp01AFQxu4kUDZEzo+7BLWg1NUllhN9unRPP+TE8TSTkI6tyEkWjhg8k4zKiHTYRPlDIi6w
anC0Rf9+UCECrC0puPyaz6lxkkkO+GeIfcHq3r2ZFifSKuhTT3DosrCQTS9p0X3EG2H3RTFljNhG
DhYHFmdi43TZsmh2R3NHqP2mZs6Fxv6QOYKpDGJ8Rc6C3aPfzQcFmjssNJcGLuvWMRCC33eqi2XR
Y2QdbMHTsTxAgUvUAV1frzp7vxAlUQf8N7C9bNwrizL/7WTsavSuNDfbaoLgS2uAMe4it3VaEbJA
O0EpMGR6RfV+ex8rwGcKUw50oQwPOEBFLU7UAOTgc9Qaa8VkMmNF+stsUBJEeMHw/1nGwdYZEqjH
MB54e61sNYZBU5hOBAKgUt08dx3JJxzUkWfWzRD02mwCdw67oVlLV882FBF4Pch6CrqTHU05EnLN
Mt8JbwcQJgYAx3PgRz8XwMNEq2vPv6hKOfumNqTi4iBipsx3YJ0krN8+WsJ8QSmiEfiLxvxqsCTq
7OzhLhdoHCqFCHw5cXUqP1jyRe+XU3Va3X/P4wcmnQE0zam3LjSC1kpdbvDmoUaQYHewZ7XvsNs4
7yx26BQ6b3xaq6Z20lJyRMuOpUQzTNF9BnpkUxNJDvVvd4q8/nYyaI++7mppuBN59iFauXQWIgcC
4vreBUFbivwwgo6qFq5L3aOVlsQKiHR75MV7r+pASAtqL6daFJXTir/IqAux/XDAr0sh1Ihd/kxH
G1wak5WS+jAJv2HW5vyKZ9nW7QQ4zB4vTI40uMNl4ITWPiHlIcFeFGcTPknuoLGzgJemxno5263b
VT+isvi1ZV73zFyHqnownz1OldRjBwJPlJ72TR39ZtWuqXZS5NtNfow8NWY4jQlnmA6hWXEn4nvy
s9zg+bvBZ0Ls+E5VKCPWlN772RA/GULDLlgviIdu87Wd/ba6tULbj9ZRh5/nkNVXQmsqGfegmnE4
dZKzdJQ2I9Atg+cIHSOW6cmsFVoGX0Qv41fMVwA/0pnWYilHLFpbtSv/f3zddO1/5x7LXjEJvTMG
giR+ZsA4LUhQY4+aafgtElEsee3gGwzYyoKcjgXmkCYPaz2d0oos+R/TlJRQzVWj96FQWprGru08
P4zdeA4jAiTF6olUQjLxIQ+UBcRUyVQTDFftROAA6Lr47k68bUp0iJ5fDEz2WJlcPsl4kxqKnxCg
tUiFEbH95v3PZc70VQFbkL6RPhpJSNmUDMWbh9RK9gLikHzFG/EcNeS3fZDwnrLJ5FSKXcWyFnD6
FJjtnRqBqMPI+b4gefVwcLD/MoEPbZzOnSHHkxSUTCgGk1CbFRjqcsiLUYn4FkJZAda8vOu8vPs9
/0bdYfb1Kd3RoWs2Zx+pP5i0ZKpE2Hl2Ktz79Kh9KkMzKFCs29ib/bQIFjKy2CGvoyk2ZVnNq+jx
ipU0ISAvaTZrsvSXsVTHE0GPsUlgilBeoyH/gQdrMZKtLxRjUMkqpQfj499K3Aroz/DAP6P1GFxL
fFXPSZjMVwQG9vRB1igo7+K2TG0stJie3uzYIeGSSsTd6KduB+linFMpYM5hXguTbti8bJobqvxR
5icYuGx0hw+yTE7hWx8mCn61t8WdZl31Pz1ZC9ubHTSJ/QNgqAHXgAhkfKQutqRdTJ4Bmv+GNhk8
k4eQjLbN+LiQwlgWPgDTIBzkltdhnLUZ8XgFy8E2lpUPZrnb9hy4IN7gWQXcPMEKjj3aCJzKg6C/
d/hI2P2m9EBeMSRopuZo0PfKRwcq+2WO0Yk0sVm3Z6fLGQxnCrwjBH56ncvVs1Nh82Vsi5gKvr8u
h3do1fBMCkg2DqD4Om9o0G7f2bZzpnBSS6PQBwOdMk7bUSGtXElrLb3wV3H3h5e61uJ1uYSVJN+V
As7DfOzn5ig8nshW0rLJWlLEPoU2jtLTYLfj9zdCb7CS4DnnBK6GUnCreXY291xJGZmWBMI31wYh
6AlBfXv49frUOxK2tgKTFgGBRicNbtaC9dm5sEV29Jl54IHvdPQdXwRAC1cYfIN9SxHejS0Iyk/x
LGSaFc0+NE+I/kKhEW356h582anvM1umhXp10W/6zRB+P9+Sa7tJOYl2zQVVGStv8eJn8zIpDTn3
+ZuyVWyJK/sduRnU31q29E8L3ohANvXXFQPUoLhlWP3IyeJqMhwNQfgEBTdYaCWbHNemRpof3LDU
/zCSYqe3irOnbWsbwcMiciutvj+Gt3jxB8iqHpvums1G7YIHGsAl1wgu4GsqiL19ysFk/VjYFE7t
Pmx3MN3TemkOfaBWBaU0/CC7RkjzUlqLll3yiR+OM97OO056M3yuD8YehJAJB6Enn6g5i3r/zjxy
yDZUj9pGC98DLk2ERZroGLrOfG8Sr3FdDY/IymZtvTf9n/9SVRNXiZ8kufWdT0byIPmzI+t5h8YT
w5arf2odN9+yjgaqe5c3bypIG5U/mFmcpcOkX6ff8IIDGjnSVwuzvKrHYieKXSDn1BInVropIBDl
S/ksAH282vtC9ooTvn56sqEBwXNYUFOI+I9tBi8twgT39y4ehHHcvQBDldu4GS4VrrszhVKni+Bo
4gsaHv6BXr7qaKBqLkr0fN0oDdgeMuNn3gJyRBajSHrMM5sJyrfxGHviVUbqEDoxwOxrIt8FJpa8
fdCoW7yS0xAYKjFxkMvDFbsLns7oiWN97h8/wENvQhSX2Y+hlaAKwFl+E+D2BH9FIIsOsvegPJXh
bA5HieRpVlG6xxy8Ow+923xb200oggPEwnU9UU+WujIO4guxDi1U6bCutjfPBnvFqVt+Oe/R5IXk
9OfS4szcMZYoKyAuGD40lin2SERrryvsNr62WFZCPi4hhpcdGiOycZxzHn/eKXfME20neCKxP33v
/VmkI1rx5/dMTP6c3LBHQoopOA4Ul+GrcbCMxPazs2pVLqqDKRE1ohltuGTBNNjLg76zDbw6IYzF
LBZa1eMXZGkIUC+siA+KqwymYep9rDvQOmBhpMtjNzzw6fj0zDXFvc1AduWzKNAIcKBA440e6mzb
0VhtZK+PmNrGOYR3cGpFKhg1OovdTMIahoGRsynvDt9yzUWW58iNyBwamKbSrT7vyJNOmGIZ5Hk4
Kuj9WssgsnoJbV+CmmOC4TS80WqKxvfbASTOl3TwjMWxBA531+5jrl7B2WEOov3ct896yahYTsq6
xvXcArhrZypQuESu3H+dm8FQi33133Cws2EoPrn3SfpO/ZAPkz7wfy2B1rR7M29jzRYXfHxrkPoL
pd984gGZjXA3dgY7JuF/8KX8vv6vtI1H8nV2or3YjVICIRzmyMv+39Y7L28dBsnL6MXdfPTtpTCT
iuqsm9BrAtlcSTBjMcQ2m8yCUOH8DrzfdYXTA7fM7Ii2QEUsFKsDaSJgXvfOAgAH+x5bgXfzdNut
IO/h2uc9MIFPmIpw9EwcAiEr/vfF4NzEvaMk4/AE+dskahZksezLtGshEEL6CPZVbrqPIuO2lTg/
NoboSwlQ6DkZTbN3mI+Wl5kpqNwyxtV8Et09dR5SlnX2ZU26O0hLTkT2G2uQFc4fhagPt8Lhw740
AVzTV3x0T1mw2MGqbNrH5B5vvo5W/1ncNUXSRT94Polsl5bPWt1Eur3QtpNklFUISkSN7ZViJPTt
RChGE04DCIvKRCqONccohhcCabeRD0HJLbisBahkM3TzAupeJMkkg82D2RC/OQf61hgo6AMWCp3N
h8wWQ4GdBEEFayg2Br2k6zstRTNAQbPIc0nsKWBy+mSNMX1RkynhtZmyMuPvTKRGnWRCfs4VUAXa
E0CwLrLYCCxjpld57fNzJBhH6u99XzZogNL1Vmr4HubBmTGrquRF12gGaOmUproVAl0mWfLIB4DK
mVkqpbdD43pEz8F4Hn0FBBmF02Ky2UrkBBAuAf0leeh+/U7BUAMH63Aem0nX774RcG3vy8jRNCzN
LMrc/zkq7T+h84sDH9Ua4ZjIJi2U5FG0cXrTaQWPKMF73g1zsptZkqhRTzAfKEbkrUFmDtDNVCGl
VI6wtIJ3rJhlJKn+aayVw9gLmJTaOBwAguBlLwrrBcp+p62ju2tFfehi3kMWMSFvmud2zgTeewWg
s9Hc5nPZDDTn/vBQXXtOCyXeEUKrdmflCaoMaMbqhMF04vN/P7zWm5dBN2+yRLpmGxmBDPnTbg4B
jMuEcpnp3j2aCF0fnTlyhGiB1URUTVt+GtlBTBbtAtZG+sxWZSCchHpDeuN+ux5xbZkyXcJCi5c8
np48n7SySDz4ea1f+tsT2WF8GmmmmoTTkkfWuAPaSs1HIHWaQ+TmdQ0cyl8qfImfbz8N3YzdhMPF
H+pg4fIHRVsrAENQ+lUZXsR46aT667Va9MElItBWz1MFY4XJ4mEUC1YDELjUYJnAv0BpFNpcb4Ka
Sj98E+3M9Z94LK6Ohy6gtsQ4tUhX3GvSELQQfjUjs5e3EcbPKpzcclQzy/H/TkDOLaSbJ40qxU3D
lw936G5/Dzgl4KC9HBN2H3pEC7OxkPZHpS/AWyIP9z8lFtdP6zJYkzQdspEqPtXQO37yNn91imc3
1PERRYOfCqdf30URfxE0SiFpnLvKp6/dangtRtCALksIryN2JNzS2jFIuQ7lYaRIhQv8LBlOL3n+
VYuIalxs6hx/nuE+bnnr66SaxwyEgz/NAOxM30bLfEnGYgWKKJoCXzgQoayD07M9LS++nCK5wdj5
g2ZNGPummsrlDIR2Id+vFETj0jU9aCfJ6gV5lEhYf77/4IeamXwbp4Q4KarQsdUZ5Wq/4DsF5TEk
bXt/qqOTl645wMVW0HLGIFCACzkBkpY++gBMtUn3scS2QD9OYbIJfkVspI/bf1fJEk323C31nhmd
8O9mH80VXBIGdEeiZb4ZJatmTZfHBtEZ3WiPteK/d1qaaS93oYUMbDdaSBPzB2gORWPIFZ2cxIG6
8X59WvUdIVUaWUDOgVytCJoKegrfaa4xhu0CQLguzDnyFSxgfpkug7TeKgHwq2PxiOjf5xomivSr
MqA0tKqol6X5FD3Ce0xCjZy7ueLNITLPnIC4gKvxDmWfLzaeKTHAccoY6aZ1RvTVBjx2qWl5WtA5
A764XoeMFHbeGLyjzNAuNvvjnmll3gfq11grzXEzw0p43a5XWyWE0vkSRSccyjKIaVdwZweeZR8u
TCikpkWz/XimqD1gfJBC8H+JvrwchuVS0h/0iIq6JlAk1Jut0IAFbe9hkJkvPecMiNkPv+melQaG
cKgebHQAMtfpBsgJuQmZNXCLrQYaCYoE8NCE1g8XvG8O3V7kU0PeHXoddqbj2XChPaTvc65LihFS
cWTlppRGZPvpggbLmPTRwydSsv1vRR1sS8tmZq+XJaTkjpwVDb2WJ65bm4OTNrSc2WrzeUIdzfVh
MKLGBxdmnVz0FAYO1nzMJzAaiDn+H84YmHRPFJC/yj1TEtBhS0CTkzXZPxN5/FGIOyUMr2r4LjY4
9sqYlNC7uaEr7DhLYYHLzCl0QzaZqXD8EE3KXXgH0ZXxQgT4ulY5BHc0C3kP4AcRF0j49jrAfiVX
1C5TMEBSAdi4YFpCLETSaCRMRtG8n/OJXHNWYT3I1Iozq8QqqSnZayb8t4aDpBB8wTsvqcWDgTlf
63ZJZOqeacBmNefpoCkNJJC7dmT/P6bvm0TDjY9k2w5F0KyBVz8mG6+GcjYRG6TkbQpouo+LutPS
XW/ZrZW0PfjB6XZRk/0kssDG5GO32N+leLtS8qwJiQtKYOQxgIIIHxVgpnfN8wP13bRb1p1dnRCS
Ji9wWnvLsvWe1UPBTZeVa+Tz+nRO7Rk+d/NRol127jqKCF347GCo7QAZmeC+MfWOSCK0SlyZTVUs
XaPej9CvQttxOkwQCVEVC2IbK4+D2CoFmGYrRXdxQNZ0IgDwmMgJBZRUvvhCLPKJW3FaNoMBe/df
ii9qB5JZnPontNHyyVhP7N77DzdUZrN0dIqtNp5Q4KCiplz/fQnPfDvmRt1VS0wDjTJnuE1AFVdI
q7EFzOsX80MFcVpma8KU5ykq6wiDBgKop6GRF2iVOWd4DvF7P7gIC84GI7MiddfPBuyLM4ulhOMm
MBYVk+83NqgY7bkNeUHOvqHgIHe+TtrJpmjfhzS23svqK5r79ei42te8laFahiQ/0kCmt6+w2rWX
jheXMmoGUD34WLwC+YmQFTPimvNnf8dm0dMAMTa4Ea60x4Hu7CC0ymvE1DPH/4ianVAqDIqDw4AN
YAkRte4RLGtsbGWhXng1T5aLRI3zhf25pSgA2GPimCQ1cb2o/aX0KyGtRpsRiTWDQegP0vgBGLLO
11PTvJZn1PV2394id64e39pEbEmoUgYq68Ft42XmElCW6iDqyN6ATUJ4WKVyzjwxlBY9yLC0F7hF
G95X3cPkCawfUMAIcUwVI9eSrVV2muTnBgnOWxvZgcGuY199mDR2+M9Gzl6VPVXDvSWfZfkUZBES
rjWcrmcoPlJR0uujJRaECjwjmUaGQm/lu6SpV9PIVy4+VyQgHEg0RlR5pPXpDeBKazJujwQ+gDMv
1LKPSUpRjFquupSF71jYOF5KviBew60rkP8nzzVb1jGHiLRegI0O3TKSqVuGRlwho+VIThKjldRr
QCG9NtdgjwcC/US9U/N8tT6Ljy7QfMM1KcKIbgSs5ka2RhJNZvOihu8Uc0CVNKrxotxHu6YqZV9Z
nRTCDITlhGh9wbVUG9nrBdXjhcxTZeru9Tm+dU4lz26S9IWRE7FEDn3lV1+gHZ7f00/C/iyDxXlg
Nh/GfHFXD6YuHS9JvH8a62+pLQvlW9yIPAegNBPBZ4+iTwaTz0loEkMlvNU082AQQ6pZC13I054w
D7gU3BEIkK6IYpb3ENcNo1Kf7TcyLfpedqH6Yzis2AEqsPIfjzAoo668KV62BSYKEEQV/DAFOOb0
t7mUFiGa+yCEwvyvIT3LEbPIsIC720n/TIirpoElD2jqPHQMApmh13+3MVSbOM4RtDPsxaO97p7l
YOEDhObcMMU6nremMbghdTGxiTj1R2KvAGP8LCulPR2Dmd+jEPdHdRbS49w2GVZiyhj/86p/Co2E
5zMjet8VoOOqe4a9ZUn2KefQ9SBKDwRIKpDQ8WAzuqI3LZ08lpCAsET6wLbirJ1PP5kY4oNi2pfX
JT4dlnFssYTT/zGuIcqcc/H3XOcuGyBYf+rIRavPdAiwa1hFqLscXbUFIJZVRDlMsXZJ5/dhAQRE
lZJIx33E82XYEB3RpI4StpAG0mAWDB6pmUBFQyOIfUtLShx/x92LeGDCqGRg46VSYRlSYydonThM
SczWV9xzJU6jU+lMwZ86gO1Ef/fSZmiY6i9LuBCj6lCdrs0Zon0HNyehrE+VtKeaJkxmxOItOek5
CLQsE0XVf5frwdROkKq3/uu1QCRwrOX3ac/AZu2/cVQCVi2QF4zOzCXPBIy2AIlilUwNqomNdHwN
CVgyfqM8Va//+gDWDY7P8iuDjnW3r64Oe2oN4l0lPIpTS6ATDli6d5bAdPjFLmEYdsof6+8W0DTo
2QT4uDbLiH354zdQijqVoJNwCIuD2SRuFbRp9Vo8xAoZ2TGccmVEPPWy5KyYNqqw+LeTaOQcljxX
wjY58nY9eNY8VZWLwexJUBWQD5yh+I7/HiYV8O/Ep/Tn++JA7r64CQp05I5iWTEbMQvzFOxMc4io
sWo+HexXRQVWtZ171rMTfMe/Mey77CLsa2a3d4i9m2+w8TIsTT25NHPLfCejCA9CfE+UC+rtrP0C
KG56qL5d9/s+4mbpF+z+TTgPQu8N4FBIOKRNQQPgLJlsa6hBK/IZiyC2SaaJFbWPvuN2Ia+AF3oW
Ncm22hfv1EKZv4XmTUVxKev9d/qrrh/+6B+Vgs7tbX0ghOfXiMGd63/Lqb7uhzSCUJKhvmJRoD7V
bsGSTJ/gp6cFXmkvNOMGa58E6SrZOWfGFt23X/Yj3HIpz25kUUJvm2WX5TYtLEXj/PNk5FuLOBW/
4j0T9aM/3W24E5lmYGj+a7vBrqlwx+hU9w6Q0Q7DVHTmJ+48BxGqQV9Rieos/dwNOQrZCG38k+rM
r1txdn/r+iCf88q/loU/GOCaLTNDPQ9Jvzcs53YqgTO1/By2whfnfi38lNlXsTuw639KiI6YFg7J
iACXif8+0ukBaGixew/XaES538Fc5LMSw4eckZQHCXBJK2sXPv+li1RJFvsCl3/sggqAxudsfe0U
HZTwpOAkq30E4Ud+gHv3aBlyGg421nadp3sPd69R6Qj84vTQPmjUnkjeiG3LSZDiLKbRe+iFd1bo
kbqNw1MvdhRVuvtnpLztWZEzmqhHe/1msSEILU03ywLX/IwS6UaJSuXVtfS5D4u1nxjozb+v2nJE
lIJimqMTujXyEZrVQxDMLVIgvBD92QcVc5nAuVEVqOPJln2uDDuKIzYn/yOMQSLKkXXrr7ctRoiJ
QLIlzKVW+1b7Wxgg99iP9bLIUmjp0RjcwAO7Uq7Tt2sR3R5ku//gRd5+GkLvl0GG7gS4fJ5ozw42
7SVNsTfAj5oG4HQ5H/AtrBDO4Tr2MtTJYSHwOHvRtSl/gMLEg7cSn/fypmR2mLv7t6OEKXaDZ6hY
hegqn8h/vaQIUGQ4fjMo07yQWCUmX16Q/PEwnW2bVInUmTkgzTyVvwlwpnL9FHnk3vqBOyVvlDiK
dJcidGQj/aYSVkwAy2Wi9/x0EyTWm01KBbrJrzwZaR2G+74VXA+bp1c/LvSrWx9Ekh0LQLtRWtQv
jvgGotnpAMOXaFskrEi9HRhrUjULpgUEgm7mSIc7Ei3fn6gA64zIcAf1qk3re7+Xi4HQbR4lu5Wf
5sEqCMc3KBNb7R5zy+YeJkd22y+OhjKNrds7G27YiHOp8PR4jR4f4FXek35ks2eNcttjGvVrW/uH
BDbm4xW2TNHSoTeV8vKO1fN5k24SZmj4JkIma3u6Mpzb8uwXM5UvpL7UXQ89z2JwR9ThV84jf0l/
cMsh4oycwImy49hOJSMPjQIRb6ZCE/0u2XieSFrCHItAHtnQDoS+WqB9YvveErKFuT+sysW5ZagX
0ckGBiEottvADbEam1T/oXa2/sgNhhE7TEbxU2IAxxzbfm5XfxXBrL7KsYuWBAKtfKBUuF8bgfky
t7l/CuCp+Zhhm3vJ3WrHFNxJU22PLyqH07QsIu+fixvgAxsIx8lH7pa6kGAkTgdnI24cZep7PORE
Th4uPyZ+E4ct2StZPbHzdxsXrMXDNTLZDWhUddG2nuWhWtKeq6w9an8XIj5AinnQ9k+dvYmYI87N
AW4I8zUqb4AJjNGBtD7zpcr+FDD/t/egpzXxHmhMo6d5qoCeu4OJrPI0OLfQnGbE6NuTrAQTPTrw
yrvZXez9H4TwRy/4U6SDBnKXbipOqermG8nn9VifBlg8z3CJs7CwpSFHWh54vCDGLEdq/hP2UAMm
ZOmIdwskLNU3keB5KKTRbRlaK8Hp7visKvndV57fnJVJTimEhQKHb4+Utfs5BDwzpOVFBEuyNw58
O6OixXdI7EKcZ9J+FYfQHzJnAGPIoYMpUd4dsFf2kJGijXC7vh9Oz3F/PqjUTFl1+3X8bW8c0xuk
MO3jPtbNcSoel0qSqa5NB0EOArnkt3mnAP36JlqGqjbci5zkycGFF1qJqgWVgkl4FdpGeAP2/sIQ
79joRwvbWgAHq0zxap0/e4QDEX8QtHMUY48xf1N1nLo5Uy/A3MXto1U9ALr5SqenJqpPAcLS5MXw
+5NmQTXQBCkAmEaCKfWGcG1brZqrrFw/THR6OKFeT5mNwqcptuHC74Drsh8fdnVavILokmC8ru93
pYEI+KJbqaIiFPrfEtQdmY9QLltw/roc43Hh6Upy6z7LCt9C1OfPUf+ZQSt7AvOm3bO0We8JG5wB
Nor9G6CPnE4hdKDA55/Tj1q9gcDEu/k1/YUXcDOxCxCP+uGqZm4RUexg7YZZX3HtjBzl4CVCHJbh
Ug7fS4R45+421bpQnBLpZmfz6lHqodfNINsoXuaW3YxzV70g6E7rDn0R6zmp5GYBNs0W7hC8v8Wp
a1Aas1Z2jhn9snnlCzV4k+CLnx7D9hYA4YLmNHjebDfKdF1HYwluc7mvLo8Yi9ZqV63nnbMBRkeF
cGQusbRpe3cyRiLnjXXqwO3SAiz1zW3cg6+++Ma3Jhm8tm/vDHoTRU2rQDRddczMI2/OqHwy3qWA
9HlxoCdg3buaVNnhmMHmSeeIljsytE1Mwlu/+sbz8pUC3oX0WKhfE0TnIefKzRqNM0j4bZGMPmkp
KUCekkyOCjdrMwt/fUJLbk8Zst+ZAdnnkKDfUNclari84QnQ43I+IJfeGpzVyb2KYj0/6DissSNp
4h+naC3EZGMKpph83lk3lODu+wm2nSuXA/4LLd6K1ICazIklmbUCtBtWYpDqKIUNNDojzY3Y4EuZ
CPpL5ScQa7rq5kU78E4kKAJd+x73MmTQGupWcMYGVFga6NjRzJWgfa3Vfg//lMggKHRzI60cUumu
PAtLHM/7R2FD+haVdWE84hHULxt311l45arShJf7QaYYptkG11Uz0OGVOPgrVNP++XVBU+meQjOE
6wjZnENAqkefSviyQN64bW+J3pHa6/HyglIVTChgW7C/Iqbvo9nW09/tNn3bTWjHINhV2OGG62wb
vIG9YLSS6DgbyYTeaNsRELRp8XzqDTFlV+oimNVLEXJxlv1zsWP1OJYeg12BxIRc7Ezc6KV7lxla
/rC9sPzQtkTFVhCBM0Ewk1FXMREc8S/89hQ5yJ7iB8njIUxYLY3xYWA80/AjzOTiI2aN0befdk2L
H+Q4KTc6rPYbmcOCHx1eixj/GULvZGhVNMUlTCLMccrQ3Sb6hxOOJBm8Y+GSmkPqNJStPyzLh+rd
RissiEp/HCG/h9Z3lGKTM5BAs5ci3WbIfBh5h1nX4wXOfKrFGG1C0i1y2UMM59j3YpuAun4Taodo
xW3dm1nGyjBSdv+CIXCbGM2exeooATc4QoMjRaLfbAE1ECr5KvPzJXbpBrBrRJ9C5+Dx2X7PGYek
iRRfOSWL38H2XuTRow4BvHksf/GrzRtIkreIx636jjFXUQv7jA77m7tEOExt2M3gFC2P1xARkDrC
VshoNivhTBSvu4a001HGD0PZk6ikvpaQSKwp9LI6mBqaD+arIZmXLbpy3VlJeFg/Bl2PfB128+Kq
2VToeIv0dwVsvPfH5INANTBrOIJ6C0179RC/W4Jc5APLlA/AV6vw2dFKuvm/fqj+9oDAv8kd5HJg
A+Hz76nkHOpHlldreBeWrECJHpp7MpkKjscGaNNzGnSo1uxngO24j1B7FFfAR4fnrnad8xjYyTt5
8JwWjlYGcyoRohIOjysoGJ5IFnh/3TgWPOdUXwGtbvkVgITSm0eWpOKuvP8UM7MEVX2qcRpRMf7m
4sSZkgXvvvt6uVJIzrj41ruG9FrVsVEw/dIkoWT+Mts1E4cQnN74ajtQOgn4PtJ2+ndomrwNyyy0
9pVJ3VMuKcpA5P45203L+B+TC3sV5RO2QwFJGsJ4+PmXX0gxUn/Ne+oQ/sq+8gwpdkC6SUh6IX5M
OP0AW2aCCgvee13qhu9a5zpMBFR9Sc5lBcvQbOt0NrUZXrPXCqg3P/AWxf5ZPvatnlNBIWvlCjNy
eWABClXU/MWBawQ9m/j4hOFTCvuEt2xHubLlD9fzNlep63Xcqj72ddASjcyLMDHI5zGZuh9WkV3F
YROYFsaVSkq7MuRGlWHl4CCH5OC0THdV8GkpJ6dDRW6ImZj5d59N99sWc4cCgizPoPj3DbJXoDgT
kXruoI/EamdKE6CT8y8QgERkaD4sySQguE21ee8ljIMU7LbhniKlgYoIPwCzj3/rvmv8Ohqzj7/W
oUijWW41jJnLpmKxThYVtpSnfnqfQh3VSAOBSbZXtXeMJPsItfHeroTx/yxV/nj+7uvlinENLXKn
H0DMwvAZSn9q5Oz6ENGgjedM4xdsx+afmE2saANat+25yci8GicVNW+tS3r2qf95IdCiaz5EwQMZ
bqRBvt4uTRk5riMrRH6/vToO/XDpbD9DgoFCPs0lQqJi8DUXs/LzFtO3DDHx2qRYcX53x/ugJ9ju
NvkZiaUZUCAJ7KOKJYQFQ2IvSrbW70GKK1fiu8tfe/YaO3Qs63aeW4OS3OuPsuNBpY9cV8/jpx/H
D7IyoYV8th7rmeCgnbt9dCHMpxmoATZEHosbx9deo8BIcZ0TUXc3mtnFVyhQAn4Y76c3ddKpaZBS
6umP5oQP3FKEWYhRIQeTBcWCVNfwL4S0KrJtKiwK9RUx1Z45X8XkN2hSqXGq8YVUumIDFT+q+I62
WqJMzQANUVpDkuNYRiNQIEH07j+Kmd5/M5+2VdLLMJOrfAtzj9jtIeLQZzF2D5DNA22qHrrbpggB
RBAswfQHIJbkPtzYgdDOBtbWFypZ3tNKyc9Nd7cGjlSw72jVOm8Xt6iYE+hdXBEpT8CpzBUceqUO
l/dm3sUP8WFF6/FMVQv31GINj5zsPcSxaELUpiu01j8BaxgifuNk0//ODDhs/eP3F8W1gjyFL3Zj
xcTBwwwPWtCenGMp4wJNIx6hXMawuZG7PRBdiZrwmmf3cMSE05u7tiyazdB/s/s5IERHOwaKnVa+
n8HBHLiHcXJ2kQmx/CpLCX7bCxaKuyouHae+HvkGLXd8QBmX4+uqDFAGt69Y/uMYibXDcg2jzBST
/ZgZF4mjDJnziNA3zofnG9uEuJWPoBXsjf53Ei/54bM/+qqvQZHJm25Xc4Gj6FnUQQd6wOnF8OcE
T9DfI9fr43qe7AKuszKUkgeCzrDb/sUmHdNRRKaZfp4Wm2AUmDng47rnSYT1ur+qFrSlnfC5VA1F
jJemFBJAOjchVL71R3sYbwUXoVHhmg9fAryfMusmtHHajThe1pECE8BgkQnHaXjOKgAf5Vr7FaKd
FOm3FKug1p4BAvwnI2vXrpa+/6lCC/8VVfMn1iCUFKH5RcINogE68ceizpOlmIqE29C7KDPAE71K
iGVxLRjF6fZUDRfghJCJpmgKiG5VlEYgSnR7GIBTUwZRFTKP1NFAnhMo9YE6y9JS2K4+/DIzf2uS
Qica/9HmS5Q5eCHULHuda7VRGa51lbZPTgb0jQZSA4XCf3EnZPxea1/xMMV7rvuIwnRBhJUgab6n
jNrELApApVdqynBUGn5AR/0uNXyomZfowREhEukGacy2XnhDiJT94Y3wlbJ3V4ruRqh7BZEPAle5
x56MA8nT1QUgILzcFC8zBHg5GpkDldW69TczpAiylQYQ8AdJ+hHPVWiBgRIOGfmiKQvc1UsIlDDT
yZVOONGTqsQalw13hK7KTxOS9IXIRU2PLzbly5uykvwdpIl2paDyR64cs7zuL7WwkC7yLNKMM8gC
6JAvGwEqfNyEzeshtU6gvTlGILKdTFAEHrNBSb484iNqWdpaEOgkWxc+wAT3FuhJyen/TjPyaEvv
W3LV2l8QvgyEkf3BhL4WRHVWefGw3CCGeg6l127BchKo0HLty6nmAVLEk+NkzTUGwMfJIswkvSz9
jKRXYbQY7HYctW3V9kN+tm+ExfEqrJNZkBB8haZozCwC5Yqle5zHJ9c1DQq5+bE3pyLxt6l/3L/r
tKNMmHe7UebeDXkTZw32EJW0uZBEK3km7nRaJw8DPgfjETYezbl76ih22L0j3PHamzaal9jjIyEO
D2mSqx6gFDr88lv9LS84R6wqDaTuVE++DMBfUrrgT/Pg8d0RQeBTBd5GK8BHdgWANhvvGhbWT261
khmyPWJ2KOP5otTQwdTy6sAavioyCyhqfH7LwBP6BvUoW6LmBGWGGIHTsVOzr0eN4dAGVsqBg/5G
yphmfJFVgh4AdzK3XSdYI+6pkth2qv/SNR0Fb5WW51R4F9AjhDpiyYaiyFy4mOa/7787MLkg6Yzm
/J38ORmQHq7BSb4UujHgUAwol5YfWMX+vhqxBYXYs2Od0ouf7+W6x6iVJCDiitXzhhpUCthgPaWd
u6mEtZMkQwAGwJERL9YjavSNw774OEZPrq//u1gcj8Q/Y1g+1f2QP36pVTLUHDxhnA+lskwRiYfp
TjNvZRFhZ8J+Ob5wCbbLQBy/jz5uAFgSZRP7Z1wWLHxCpaVJ4RSGricXq+bEgZD5AZUNgue7PGb8
AGwGLH6zBFZbVpQ6yPqiIABHZHH3wLr+rjGiHs0P+WeSOmUxl0DxcbD3WL7C5cPBDg46a8C2z34W
sMpvGl/GNYFmrc13GMFPei4LWA6teT8AvdHcSvpiyBEwIa7ivFIIjj2MpgGlJnFXasc5Hk2figXn
dkYEPRsMZDvyH4VqnFxKUNLxZzRP6k+OrRQedCqHKUVi7qhM3QCIBU1vTFTTNMVVob7n88kD7KLr
TI1uXUyMTkH4u3NXpFAcQFCkShrJ+E84tHTTeSFCxCx2IbfNxuNtQ2WDQd+qheSSSetBLiPnnV9Y
UgOeIJHMpRRYnvB6FVEP4lXcSvYbetg2DtCDdVCRPRWyCmR1Sqg4YS96t6YZCx9KG/Uavg4WLkkL
U1HUhisL9zjRdUWPPJDmEe2xFkBjgl8Jp/o2+zJmJP3nxP/Efm45RoGmdRPiFEhuSR/C2gKd/8bR
0LJOQLikcN0723tYNDvnahtOiOV0UmwApEM7+ksx/6Dc8psM9cTWJiHilxJm9mADLJTzmBseRs9A
d0knqasviaeC+u/TKvFnqWrvckXvm6irWHjRxVO7O3Mi47khI5uyZ0dXp8jjDDVgqBwZMywleR1c
RQmdQ2PvwOrz/6oExZkMMWdtijNVioKGgOHMnwkkdKuMZonoIko5vHO1VEyJx4QJnrZb9HIOPdih
NHsKebYOLNmtZQR6HSbTjjSkYT3MOL9MwARdjA1+UvQoqKbfbaZSjrH4z0OjGcKjH6oSs7qtV6mL
WmwUib8cjzJZTg0v5Xu3smFDLeG36KwRjW9D4gP+e1hjlys7/6r1aT/WZRj7A/oqypv4JjIMnFVP
r62BlELu1u87SBAtY4NWUFtEfxMpEuI8SIMbZvwHTbwdn3axNh8fUD9prSolPzXMTEBmWoWf7fKf
2fvIHSx+Yp5lPawMGZRErJi1+ReXOSk0cMVnAAR8SIF8PzfwFkbkuhWLK3LGZ2GpAS9vNdjRA9MD
YibZZdm2JZ13VwccJf9rrE+xTrq+80d+Wmr6+Anq8cn4BRuI6CXvqqkH5cM9PSz3Jyg87rzc8yG3
6wjXpbfNv9rrBG6gTCV5sU7rVzgkQEmbuqWL33bABXZrU5hklxtWA0zL6QPZIFV5+VqAkVbHc0kI
7enjbVR2a71ghOf545Vw3xep2Xnzk7A/wNtY+k33faDU2Aj+WpBIpZ2Ye8OkRt6nwbA2aHa5Z/vd
wrjNowCwOpiZqSoFeIvvxTn7BZifRbCgEd3EurFK7WV0ZiYgGfN+EEppsozqxnvMA7zjUbkSVSoZ
t+oc2vwj2F0ScCgdiVKR6sFr1e5aoZtALn5CiNMPVqux2WWrkMmALoRQG3LsmE3xAOVVJVgd9jAF
YE4PiABzf0aocsrPfAqP3+CcxZKikhm9kaGJiZmGzTDsKkxUzYzu19r5ZE3AA8UIzwQOLTAE6L6z
WGkAwdLeC+VTqAofY4cEAT3kQrTX/oS8L7SjlkPIc3VdItstR3+9MQYxGt0sKNq0oRa5kjItkkO3
LExZyqcksHsi2S1HIW/F3Dh99mCi9dloNgZ0drjId3kJcs4uLMHVKVYfGXsMTHrbMLRDYQJotBgR
ISOZFZu1ev/ccOEWW78ooRXs8t7wEWVZ+isA6LnV2WOzfUBqlM1HiTSk4GpnGuNYpMvUAj1AEerY
ZXnnBGD9TjGPQcvkiYjnVegvM3jHVSR40/Ex0xkyca/Mzju8bdbJLa6rr6MsphwKoh09hy+2Jdqy
rMVS9JlR2xQXbZmyUTbAcfeD1+4R9YOnhc46r0KC+Js/+buXrH20TqjFdKjHgt+WRerZp3bDAPv2
yqESplEFCMafXXU/gQ9sLSAkIQ80jvGK6RkKsoyJMhvau19adLuyqZsbmjbKAJlsBz7MlfOv7ris
igFOJcN2uTwgrK8I5XEmHC4afq+vNBzXAqfsczEcYWl/TWKFJtzg5nyqRPK2ftTyVwvCQjLPAifA
CvgnJxz473U0S3NEebsJSj776ctCyNlqGeRqrE/4EGVJvmXUtgStShXmL58nY/Xs46Mh7Ug0ISE4
fiRKNIASS4Z6ka+dIUzDaqgTDvMhH9/GzK+JDeGHU43qcJ0o7e8DQfkdeMPxkuOFSrxEMhZ4FYZD
uM1EdST/NuyCe1UPrwZqujhh6wjPyjRBapawUUhz5Z5M0wJxligqFafIj7CbxE9gBjx9HhTWXl3e
HdPVoLycQfVrrR9oso+A9T+UrUdKpGsVGCIZxscXSdwbiW2kCtFx2ztRF7xqjYRyrRKCscCMLW+h
DAEzWe3TmZer2MgXaj0UTA3GpHPJ316N4ck7bGhkk4LJemEcIFd9B4c4QcJHmPwrMoME5nSBidcV
jqjA8rrkknhlSS+UKV3XY5kd3Ow0Que3xPud+NEwWBAahVHAQSRqkJA/sxNL6MKFPNGR40g4CE1R
FqrT4Dl7XYlilgfHBI/AhxsOzJ6qH+dY5prZcoG/++DVrjoNt7xLYlIPI842yJn+asspSsDfNYLy
htd2A27BweOLVBXi7+TFQWovjlvFqyudVsmbr6Id0qdMlGL+Lx6prJEiFbaFSIDW5cK4czMXy6rV
Zy2tsc1K9tXk9RLnhhddxVVC3nTuqZ34AsIzLDGNZwEheQbUbs5RmrINwRQFu7AKIDJv9XQhoqfE
aXZ3CU6QGrjdcWdDCHMURz6sPwBBC4PLacePUvFLiAdE4MKze9+CrFT9XxKXYtnrOeWDgNtNneCX
Qnob56Mi34ssebHGQcwIpzlidjz5Apkp7+6Ad9YniWbEDH+6OGx55KJu9xd6TqnnwA9BHcNhpaT5
IPSLaUFc770A2AlBcph0elhIVd3xY23up7Xu5T94guk4oJu4gQxzTM/DdZgUifc78NvLjtcxhPsT
jjX0z6JRtCVEsQE66PgaHHv3DtsnfgN1NWLsZOICdn7rlPo7dOvl6Zq9jsIhGwUKDlR74A0MG0un
6iDVEvQnr+KttFbQE2OOSOhNayAL+v86M3ddXdcoxh4wwzJStLDUQr3DLw1q2pxBG5DKapzR9ghN
EHB2NaLvNpGWtYLLO+TvsYvuBL8KR3ot63hy1Kn+lKMr/RnO3iKH7Bj7hyrKkH4RtDGXaeNkV+l/
XslsLfGzEOHitkc3tsVGJIYYqymYprr23QItWGDJ68B37Yc9YZq+O4sP6RIFLrpwJ4B4DfdAgrl1
AL6uTYKWBJcj/nxw++OXAMukLdyIncDKmCrFB1kDmRmDGejlYlLK6T5QFPfVQ5UO094dZvzFew4F
ff0JpEZXQTRKUMC0RdUEA/RmV80gI9569UaaFSCfDBFgc0uC9dBLjY9f31px7zIsq7yN6l8R8ggr
aiQ5lGt6grm82mM1gjGVUN0F4YlgYuqYAY4UIiJXfIH5ZNlPyODScSTTmUHG068NeigTSyH0+Fgh
2Mcvw+xhmKnV/dM9HxF03IJ7SsLOgp0qauAYvmQT20d1Q29DOV3yju/zoaL+2Bkw7Y19Mpxk0y9I
ye2JWQvuNFKSuRARUxmd5G6DOeDh+xkzxj96YAP5gHKW3NvpPPI+2tWPW6ZBm4TckkD3wO0Rzt5E
gRASN08qjURk5nZcmxDQibhaNbHIC05ZhBTp/RZ0L6heENhSSGz+B93bgPwZ++0+GVcS7as0ciIm
mfptRtmtx6WxSA/FNpm44GPk2CWFtt7D+m1gQwcsSM8d6Hh4I7O/gb9+t2x1aYMizH1Ab+04Aae+
EPG1SFaXK5IRn1r5ENWAWdVqHhKAi7iWWDv+t8m3r97ijzh0CbDqv9GkmgVylQI7IJbOewbw2Bl5
Syvn6qcC8eBKJx297OSDil6dBo/ZSiLr/MUg/9atVmth2G6XBFqK4tEXZ+NaPvY8Snex0GizM6gh
AYkYQKBYGEHJgxJTafbRNNPBDrMiz+fQTz+b/g1XDo9jmDjiQPZaPrdCi9+z/6fSk3COxOJH6rhM
bZWe3t7ULZ9s7HOtXq24zwus38eVQS6nqCQGbSh9mrMVWhwL+SXUDxV52MRo9enLgewxpb39k9WD
ZO2IwgLTvH6xyLjmfPqvDVIT8LmZztUwYYGrpunCT7NspQBEeLnk++hcRex3fCt7dq23Z6310fax
9XAQTE2EFZOPMPHQLue1gxO/XCN3d/K3D9UDDpNMX1z4Q4pPj01D6/4EDCuv5Y98CO8YHc0qYWMm
BPrQ3So5/CpEBgvO/7ISyApPNBQ6wKoAItw+h/htOw1sj+MszMHAwskjpG9d/lS0j3nLQZoVsWMX
zQfStdLwNAWT10Io/QB2x9aDuxNxRqHdEZCHw0FOndNpHWD+fqcGzS2lSCZPyO6TFSYfoFxJRW9S
/ky0PwjbKT0XWc/qPA0DWptI4wlC0SKF3v15BhBN6Vr3nJxwWagRN47gNwvBjnyK/HyxmSqd8vXO
U4FCeXQjOkOhjQnkkL6TQ6msXcK+gZDnqxyLTk7qsMzlC8YCKw3d02qDQkb2jU0uv9iLAkW5fWpW
Cvdty6EF7uSGu9VWa9HhCdfk9zWMwFNYK39W5pntkaSx9JAn/hamO+4gVGAgKqFGR+v7NBhtb82/
Zxkfng2zi6X7laGlkXcUX6yQi2ffrKydHD04VkO9DK6E1p0tgva0wwGc1KpSpNE2XilxFcVHmJ6+
GHrsGfrDaWjEO1VI8gc48m2veSL/YUnWdVLAz6T21BnVKxlIGR+xXwzU5IgRQZ5RwHKzAm5ARDOF
GXFWRE0su5xFcA3fhgdsB0yhaDgQg+uNfjc/wbU54pQczdwzGWB72aWFFI+/sp0x6sFNBjaH7fyf
SIv+u6YQa6cOJLASs/Y/QfGe97Mfv2CQhaump0nHKAICiwUfpES7tm7p8SoTB3ku5L+BmX5dZE2g
bYes3E0fO+m6l7lxmHui3E6IX1B5g09DdD5zC9zy1HdP8hDS26Un6GTw8qzSdF0MTnQOV9MRyK42
FbBJsVkEFHRu/UTRe/2Dn8L1sngjmlPDHv89s+VuWL9sFDBDhYNzFM+0aMUt3JtKaQgy1VI2BrIR
vo6myfiVsr1MaZt+bgY39ixFFum7Z+2S3HPXJmGOE3rX7iGbIyoEdwGnnrqeOJ+MK4Od5BM9s3B4
A5qinrYcMXhZywAp4zrFQ6pylN4iC8wnmubdiJrePVeV8cMuzjZlCYu07ZMu9OHEl03CW+510Wqz
QJPrN0F0fpz7S3tmyjwONCS1cZ+li9+1lsUv5wU3oYbF1sZmqEJxezOI6X/SCvvW8WB28RiCGH4M
TDltDphMW0QYMOvWEhfauOVrggFlteA2k5oxp2S1sV3rvaQHe5/ZO/dr6IPcyh+DZb4QgcKVnx8M
QWoP4C2NvPtBRnGjgH6W4DPOj2nL/Xa/O2fbAkMhs+QP5FUiLdWINIWiRB7ZTUd7gd1Co+i9zRe2
UxOZkOCVad0w0u03GGGAhfBmyNksyUNqczXEkMtHfUWLSFGx3FumYlEe8wIoANGkIp8pyJzB0BVI
YtDbvoJzlCSRHJy+fNVnJ6lnFdjIUxp+jHJtyJKJhv9nZ/FZaHfmejaFbt9RLWVNnl3HgHNI8xmm
gDQ/6NLcp925+t+qmIOT2DlXNRcGpok15yRlPfts+Nx6NHb71YUYH0TLa1WUv+jLv+zlUgmPn2/B
CJqIDQeXVwwdQqGFje5qfTd/fXXgYErSAHs0Ou2vhXbfzMRo1ulX2awQnFs2lq+LmacvXxvhD8WA
av7w8Bka1waNA6mdBPcz89oIj0vD4NRPIfmlB/T80UkJ8n38hFHQSauPGgu2+NwwIYqWMPB/m7ep
6L//kliN1WeDeJTb1F4mHOPWqRWzG1HV/Bv7hA19TTtNIbdW59TB/EHW4uq6r0YobXU+u9k4VCnT
7DNfmYg/amVTiz5kHuZXt+I7pWKbG60fh5OB3OtGoI3Kvh5HplpeFoEtBo/ZGvNt5pAmJ+dPRG/U
CsDx25RPe9bhnpu7uR7MF8ltphy3ZUPQqE3f1T5634RcMutdj5szslTYyPXz3isu7U0n616xZ7Ge
s3X0mbIGnsTeUzYmaSZLf1ZbyvnxPa90EHWff65m4CZPJ+GZzJR+qsgdf6cWtX+SZo82KIViUQJK
Jjon+helg5gASX6fTle4Ctu9wctZsYhmz2Md1M0y75TgT2vO6WTxG2j4B9t13vqXCUZJrFWB8o3h
X58hV4mFsuixoDcS3gdAf51WURut0/hBN7JB4lcQZANSlpWYTKcTja53OouoIDmeK6rvK9PlnBxK
JWc0342YUTcz1W1qkYnonfq5RZ42pmCGIiDFfcWncydH926vM3byn0vCavy2uIBq3nHIO3j5YtPD
S59ncQY1KKyK1W8nS3UDiHZcDEs4FF1fNgEtrPP1HDLbEbJvq+5aIGiieW0bpiVotAB0EhyCADIX
pDIjFLjaYx6dhmCbOoQjNhovwQ59AtfoCA/IThTdNNe2zU1HEnCVa22GdHUSxjFE+HlkAN+vfj+E
YOB60KsX5X7ARh0Tl2yNejxKn3DxBAXZKVq1FUS+IR6US0qq6YC39r7WXdMJ1gXq7TSYOmxTSMpr
zOJmoQqAet8D4gnpNYVWRUmL9wxX07h2ZctT2Jj15b6JTLS9WJZJdC5lFeZ2qJjwbyH2p+Qszsvc
FXqz0IR4oQ5535iv6i04RX/eSMdm/+D+Onsd5j34Ptgw6580Ws1XSTxSOMRdtnd2RLMOiqpwcn19
z22w0rbObv45Cgu0lHtPcmbii/DzEfjoYu7+p1lZV4K5x3EqyrCyOziRxkIKN+5LTugjOyMMKUVX
PYCMvk51DJpvaJEZ3YywK2Fnl+0rdsU4K06sSKwY0vRwdXbGB1r/znTOSs9Vp1mIiY6M4CINBHAH
vAR1vDY4QN3Uszx0/YHl8erm+ZPe4pGICdpFwcTrksgJjm4vYs0woKjt6ujP+DbVbVttMm1GZVEg
CDypiWWQtzD+NRq+iGEvUu3fjF/KcBo6OgMfJXhoQGcnYHAOYW/wl4GkceNXeoGLeQRX9mSV7zL2
LbNnL3u8E8iqEgarKfV50fRAubfToJrLF/3ErT0nXirGRxPqD1MaMqNORDwA5A7HJF1GaHu17xgo
o31x4+vxs/1T0vT4qrwhLEfQuonBei/CIohN4fpcz996069pVs7BssbtEEU0wE5xzhFiHq52pT4B
KxAbjfjTTIbX4p5LqJkZoJJG6E2Bpjx06rR2vI6+MK2RKVzLafP6a3OPJ1d3w/QkaMnOgh3oEf2e
CXefRghYytkhXgQxa5KZDUv/kGi7EOvd9HWkJgVMUBTJG8CBm4FsYRmX/uCDH0ZAlFYerbrQ0h6v
T51A96jx6DbNWoSZuR7OznSUqsEcJQRVok8sPY28y3DKEmQEngVRlyJPwphTBCVrPuBMtkzUhF7L
ffEFB7yx+C3coBIm2lTH6hJKTWxMB1bIb9v8xtiay1Xr/pV02rfm7gn5RQzDeZxxyu1UeSnBna2W
NCdsF13E9WPzXouId3lar5YWZjGBcfZOAeAdWdlYyEcxkgePpBrgULj5eVPULNED/l9eiVzYJMA4
TOmKnorFttw7tYYvDMbTKKMq1tFqrOb1FLYihN5vkZc6E2+LEczA3WLoKgEcVc7UO1Dpm/wpMCBU
XIP4O6T90QmqomZN7mFbgYaYfOWJIZEn6e0PXKAcBrgT1BE6AP20fXOBOSazz1mzeBWz0KGKJt3K
GgaRQhn0PUj0eSsRxaxjmHN1kkSJ2jmyHRgtr3Cfn9WrfotTDLdqvPHy5NBSontcyNluZgkbwB1l
aEp7K14PYqXQ9EMrazT5kCryE60k1jnp+BpTrPHSkHvCw9OkQZYmwYYbBrxcjftY2TfoRJLQPlTF
Etej0tUQERUI8jJ/k2JysN9p+O/MrRhfTBA7f+tZ6J+C2DoUKWBf88nU4CBj3He7hrbA/6pIYRXx
rsj6frwKmVLWOkhaPpAx7QrA8WzjBS5i6chipZnwm0NVZnF4aWFdLbH9kqlnSgnLtfKe9CtMzJp9
UuPUDIMnmNUVTkdjR0lqtTLuBQF3ZtEpoReA7HOvoyeyQoGmU3HURPmbbzQ8F2rUee9FiEU/Utjw
Jm+kXk2S/TbWgbSbUp1VNOfqyhs0auMl+QPKaUY7LSVzMBchm+K3aRgki4LnH/8Zg26ryDNxEkab
nTvRUWN6MbkQC+EEkabcaKRnexIcNasd636Zoj7DUkzzvb6H08XxABtuNaOBe86jhFf/znjbIc63
JTWm2nIZcPI373OlcZrG4r9o1Uzof1+gSXGDPXt2Z/VNLUsRTYa8L0NxlfHewPnpIBr7UYiceNxB
1iWlkYDqH0L+seXm9QrmgWtyvk3GOihBh+BXsosslw2xCK0dDv12FGZOKQWCs9nbuLrHb5Pf9F8m
iCLfqN9DDyic3tXie7D40i9FKuj39jliF07wqBQyzEuzreBuGa/PUE7/rdYqeydJUHCKoSNAMxvH
0UH+0WDmAob/+ubXAJtXEaNxX4BRer5x27TjUT7RyclZ/50MwdBjDz9IgvsglDqd61K+xrMgiyil
yILO/WID2T6QSewDgsI0kVtBaV3FxeAEDPUUi6/TvtEKDD3qvB1B9wIr4pLlGEuHQ9qMOmQfWeCt
7lqt/tIlIilCrYe8LJYFQ9gP/GSVNU5EvqTnsHN7LEjqBNQTmRHQPhpCCWpkq2OFscYQ3WypCYaT
lD6BjldyVPeQ1B9goMua+rzCgC3nwx9kX4A3d63fEZgZO8uUHL96Rx8DupLF1xgK+qkF4F58PKxN
vz1LoXeKMpz12r1usgiXgjADJvQAbqyyN4Yxj4KZmQktOl0RormLu6uJTzaB/+8bY9Uk5Va9tRqy
4UGx7b4LyQAWlqKwM2Q6YCG/ADQMoOB+s4V5C2yisX0rYTGmdv6OAL5U2R4wytMsKmDPN2Fl19yI
HAf05Y1n0aAuke6i5wwqFB9GhYBwW82ADaYBGnh2+qLjqQlKeGgGWq5NPNupVzD3JKHrCtJwIxAx
KD0TADAo7elWOQL9SMl10k3MZO6GJ/3uH+kGPDSyj9KQ1hrfqJbqw+CYDkfdM+m4PyliF6z6fU02
Dmd7lvXzBCeJPB26e4j5BjuXPJbAKoVdvBdqr9R45ju/Zs4O7gKc8BB924fakEgrT4XlHlLY7QBY
CaHdlI6+C3rrv9+ijAcaBAA0oKisCj+4tXH6q69BkmT0x7Mnzbfm8kq6VEi7fmUEvJP5CuePxCI4
6AQuo25ZdLH3avptXNOKOG5d4QQ3ED1W9F/irGeo8rFpJMWSO6dUmaC7GhYObvPKYIvp4Ud4KlsE
mS3X/ggl7JgeN5Ts+T5bxLCDV3PZKc61TbbKs7+uuPxGy4hZxzGvvtb2FCQmCgCVSoWWa3qTKFOf
0/aQ+TlfI1LuTQE/6byCabQs+R5pPM4rOFAYq2yktJjO48yTwoXuJmFrAkkrf3OK6r0LvWmN+Sez
/QfazWYhnQWkClOYAh9DYin6rzcQZ+v45Eg3c6HFym74Q/Fx5vtB+EEFxYtJEKsBEaRDeFj55+Q2
woQcT7w860MtHLKcuKX8TsZLtDMUayhwJwJOigYEe6RfEZ74W8+QqWYQBA1IekoT75mCgbPlOZx2
xPhxLbrdp7LHLAWKwhmCyBXuIntuAwL8bjZkH7+bqHzJxlysLycGCZx/E1rdpP0DK1F+sf099AcA
FrmhwJFboUPMAAqB0vl3KmEm0ddWY+XGca1xr0J6tjD2/ioXioM4THxveNErrimTPnw76eXjs1Of
6hFGCOctqw4eK0xsL51YMFo3ykIkgdBBNhNuUszlw1bdjhu+VPeAflPDKpIu6xtrW4SRsyXn5Q2G
Owdq796Hrq6E1gANv7jCvOW8VEypVotjJp4nPK3ADG+Qwu9QEDDtPQ8r0/cV0t5nu92W47gAw1Pt
Sdnk2JTaMwS91m6mN1t7FTv5eTLTzUOoevLnX3hAYAtsA2k/B3gKGb69mp2aBfuSdjToMzSamyKz
x6neLbUwj/GTIDydOVewvOp3EjAI9I2okm1erD120zGGZgnUijrvZMDTvJrWjTZVaPowq+zwW+DA
WFCjWmgjVTGjEyRtbnMLRYsxHudnhlMsjHyujykKxw8qXPMyjQevpjzzx6ilpFTU49mEuEisU+gM
+WMXcXpRmfjqjKdb56MD11PN0gq7k7KhTrje7otIINC0Gw8CVrkMoynRDjXSaAQ01PfKDDFsPE4n
O2w1Ov04Z0Zv0/GHO2+bb2sB7M5LAnoWCVhSm8lwUiNGqUndUyh16rWdexoCS5pxYyJaMCT0aKvV
Z6xnlWcFvuLuw+55SRM90yenkJC09h05zYGuxRMqrmrnCRt+78WNpj8TvhF+TrTp2I9EK0mIelWN
vB0GHJzDjzRrRZAt+tmE0khYUGo6DH/zC4eH+u7ViLT9L+eiD5rGeKxbY9hl9vDpEdbRW8Bh+R9l
pHHRue9n/g9b+YaHDhrEy4tSO9aySwwoQoojYhMMJuP1RcxqVHIJi5E9LFmDsKvNK9rB9nnqZ56r
waBBqzw0bP7BOV8HeNJRuXgdeYNLc08gznVYMiiymYn7VpExIZO+TgHs8pKvHXvwqPIf+3kAGFi9
KRdJX3YdyNQmXLNKuYRFEjAebogu6KflT3BXgcGx0gkHqFt4f9ZLMvrTsJfSUlCHB0rZfvDoDO+X
IHmRN+TdTs1pzaEUUB+dZGAvGRXMLLXuJ0tJtCEpU2w8ujQ2zz4o5nEUXzB5XPIN2XuGNxCg/3xk
4HOPm/HZ4eETa4C1L8AqCcXZCjU5ZYBhWhdnnytnrUu4Dp15j9g2L/qrgt5d5GeQ97/J5JXxNUZl
Ywu1479dyR9OAcR+RgYFC2exvxKkcxDXVWKlrvdgRtbR73b89YSE2/ukwy5ojgekDIZCJ/wfzgTv
iZpeM5PYMZQHopkUiTe2MpzFRfCsak9KBp8Ql86Rc+IncmCf5pJi5U1quL0QOn7d6RgJB4FoSp3I
u8DoLU/EZL68oi3Wbj/WvSKECAtk1ot2e/bfYV7inf5AI5PTXyGnAXF+lRLeSMdKQYGY0ZOmoyOC
hsoNy+0QWmnoXqs8GSo/GWZe6x1WbcVVObZUKM+HSV+TXOFC78bVN6eVW/qmlGo4lFmWu+LqKi64
kHiOgI7LsnwbK/hM2O/u7fk1MjcUHX4HyPa7OP95mtcF+UrY8tVBg9p5jbgfu3gOvDjgg6u1ow5A
rOZMMXgrT6y0OQOySVNKkmHKNve9U1RBrEHT6CjalK72BziwoH4ODPInlEzdxjLeY+UIlIRxNzMn
K1YmOtCpqLddO4b+hqQcxO2BEsuzTgDWHb5vcA3hS5NyUOZEwySjvlzPPn4QfcWtesVJ6qDLDKx2
YwJWZWRuuWi2BCiXtBGiPeKm9tN5taksxmLg7Gwf35I31udMg7z1TGJIrD5SI/wR60jdPnoJwGpX
k1BQaIrveoSWdhVDwH5cVuRHKAxf5AtCMve48g9c9F/78zezct7oz55RZE+FOx9QB2BA1kvJgrBO
KeAPt7g09OaBkrEb7X7MSvO1au2mc4t5Q5R+clXEzAwsC4xrxXplxZIHReXKAXnERmNybs/sE5LS
t3VL07Z7xHWjl2QuKCaCgPC8gl5wbiXInR3sVRMO82iV8oegPX17E3HymA4RxNUHiWWyLYPoPCbG
WBEwgy91pzyFZzJfhktPMhCjPys8EOzB0kJEJQnXI+vHKXmL2Kiu2Ywtjf51//gdU0xvldwFXqP6
4NhM5EgQlV8dH7ut0Qq+EejFxSLa6nzWydufsRC+Fyfy8myHoNrc3i/5WaNrv4vkWQqBOknB9cVP
+XvpfJhDyAQSCMkBlv08ZiyRgnImGW1waG7142yabq3fsqSuNLnqXaIiDH3kq8Z4L2TYsD4h5P7g
3jtLKK164LuhPKEovWNokneN8yLMn4zSNvhmLhJUj/jlBIc+Lw53MVzOJoU3ol/vOIq9yNG3fOVS
ATiQVWFq6Dky29W/dXRkMKJL6xIW8W++6l6Svrmu8QFXM3NJgrYreo16yqKZlM8JDufe7m9rAqch
Q/rZHlbupZBjSwM+RYN4mPO4Qs+FyWbekFLuGTUvz0khEj3q9r4gj3MJ0tWZzb+mQ/KnGC0aF6uI
FEitpIyKVb6kqdo1cTtxc7MzrjYLimlrIHJtOn8ZEXv7EpYSEuoKQqxa1vEdQAchT1wxo3bV2zNq
gAuxTkbOWJk/9EFCOPMkdWbTMQdmvPFNDDYVu2+mGTu4yJ0lADMFc0oXy9nEWgmsEEZTCeBBthAX
U5UkRV9LAwUe5L+thca5qENVXTwh60Z8kwfE+n9RCMmbVJQhCnV/Fwl/XM98pJTGiP/1BVORZBhP
3SGllhB/Tbv1RHAXhdGj/16l7ZtkdOuN0TBbPNR72KU/5xIqBqxT0zQdgDlWhmokAsZiTFOAsBr5
bjZT88uc8EsKZF+kq5GR9FZA2/r5s8MSLVJxVpeahNHN8wGVEy12acB/ujb0ODjswXZVqDOZ4h+R
OdAP3NnbGTt+r18nWnuKCZMpigF8yhuanrRCdHLK+p/cybjux7JAiGvVZ1Tz2E6FyuMco2N+ajG+
0xgph+w5Qxq85DAVUkV8cHdUFrxhMIpj20Wu+NaD88y8EWYM1EFlHodORD12E3tnj5MyPL9he0mj
y/qnsmYkC66lhaSqLT+VsOb+S32QOyqk4yqgV5isHyRCO0aEqOmR3YaBhMEqd9lGtPNxK6ehCwai
Nb+3cfvB8Pr6mVLEJ6ikevKYHg6oAqrnz9FhfrT1H/mejAm9z7tKDzWANqKA5ekvp91svktKItgh
WBjLIZ4Kis0I09RNPXL/vOGft65pI58nqR1VZOD4XEKzIcIOeE7cxtCgVuceHdax+tl0UVdf55LH
9wjYTJn1m8zoDR4Vjj5wZDq7eVtyIJKejfFVtUVkfYVhGsr1USuwAVEFZz5NJ1iUZMir6cvkXDtL
w7dAt8ZsSZDJzYhktfNv1qiFqoxJZwNiV0w26DUT3flvULL4IuHek/HGA5Nxixite98ufCVjNIq3
AQN5SrhJPxHtE7ka9UwA4dMaTbhJa5nSJaWW0XHCAF+Z/QqrcTA9fPdm5upodT7iWhGywgn2qE8i
piXeIKrS6/8nsWqDBNG3MEP4TqreGA1jsfp7XMPqNLY/IojHJ/OC4MENnV3EioL9KeAAxH4gS9j7
4XMq0rvptZ+f5/kEWhxkR4JZi1cX7W3g6Q4Z+8k1i68wmrfXp1/beUz6OOMAfMGiDuDF5a6+ZNsz
tHLRlLjj1jIbM/77V2MvF+hxqs1bS+T3iA/3MG5Pifyqr26nx1Eh2cMZEJ8mg/rO5lsZZxzjpr8c
RheAy5tE3PHEPG2LcAC/xi1b+0J/AessPLWqRG90jd+BYyLh/mUpKAFmgCJCjwPtU8ktIcD05yZY
Mu7tu1QS7krJvU+Pn1rDDP5fCXlWa9aiOF3zqr+LB/DjcmHkAQYMtJb4KcMQ9FYpFgKv+3IbaDeD
BtXw/jTJYia1vVzKnEPfPQsgpHwiw1WI1aKtb211mWCZ9aYtsYTTYzZrjaaVpLIuhVFJbqYBXURg
X7rjcMR2clcUmuHnuBEmU+MUQBhLCg0cgrYGzkv9bg7T8Ar9gBdufJjjTpVA1uYzvAEY+pb9XYP1
hdp1EK7RHOhPh3FGe+TP1IJ49TDMZskRS5a+BFjv/P3S2uN1pC/I4QoDUywdW7a/Aj7xwK9Ptd6R
UPXBx+6vtRi3jHKuIcJ7PbI6cJKjwsjpU3Fb3kdYEFwJbI/T+mXQRwGhImLtkos+Isk9Nftw/iUN
ogS2gHNFnLtDGuZo6dhon585DoAqKUgV3yORF+4gH8BbPsZdTmnCrSqSIYMsBfFsLvrTj2TUhFZ4
4tad51ewnyej07UDK3lRJtrNP+8/1Y2lRM6dXepmbV13u6IUuNTntkAKKYScb8ezM5NBzdubxyjx
ZxRLvMzaiItr2GqRKic8Fg79Rydh7vSxUjU6M9ec6ZTsJ8716Pc/IUFno7OQPCc5m2iGisSrXBgQ
X+D8w1wq2dq++rYE74fysZcLuSiPYqESo+I9G57FxMh8brSePVY2YZaJHXnQMij9Idd5pW2PLDbj
VWgZDsG7oVWpWwbiW9OaM27vZIDpCr7aKUJv4KxTjVmNosfQomKLRt+oo2894YfOvJsC0gEr3aGq
reLUiFgWJYzQ822qiwwxggTmfEjRq+CTXppxCkL1W8DqVzJ+le6Q1j83+kt3IImv7BwklI3Aa7JZ
8xWtJi/1Dvf7MDRur9h8D5CBtRR7ymO5wD3TiPuNKaxgm3BI7Jt6F6T+OvCTjVeIt62hIZO1GDT7
smD0JtIAKgbmsxb0u5Z8r/ONDAfrlzxc7aMK0Acr0CuKoOopyQIFW7vBxxZ40zLDsvkMHUGh4u7R
+4hAy4qBJKrPK/Y6AEsSHYTRGOuMvoUgRQssMhkQIH8ufpUFh33Ll/xfGNkFrq3RvIcbUUsiwb/i
TXYRC/Z7yrbtgcG/freUJb+dWEwjgtTrdPTpIyJD7H680ETheNg1Ib1pWNij6NcqzgozkBMR8S2K
/yqHIcmdQ22d4dCtoct6gV7eE8m3o1NTL/ZdHqMyoI5e/jG9OOSQW/ZYjaRvs8i2zu/ELQhhOC23
TNj0axwgGcFxRQjfH8iVMO2g8E6THjI3+TasJt/3FHX9umNTEi4nXhJidfXza09jWBVrLCNAYC1H
CaJEQE/yrhkpMp8m33nEKlgXLUDN00nWWJ/s81lQKl1/XgT9xQLZBPiY/Y+KbGqVpo8SFQKM+42L
LWyPNJdAzUw7cv7qeWhHVuG7G5sDi6B8xZCx6R4700BTMEnDKKl8OrGGtc7M2Wso8KyYMPz6vcBb
2B9673hlOGN+39jKOinv5yOPg5qRlMkKwdzCDg0uxeNbM/mR99Xo80vnR4iM8zrpof5FxK2SGWJm
/PXiClQmHf/PsHqo5VHCe2yeh6k1Sm7nW/i5v2ouUjdRGaN3EbA+zXr29mQIvmV1QwgdCdHwbHHT
JueLIMnMbJyoPhzlXC8TEUaTTs4AswJRiWJtZW34CZAMTJvLKw4/tQ0shdVEqNzW9JfEhDLFlTOB
dJgwvCwxSTZYYFfgPZ/0a+0G4r19FsxJYzyXm3gUWSTyAhAaF1UQqpfVxDUpqkHlvZhStYG5DUav
NgNs9UbSZj1kfWAT3gMdbme2ZwtJ8ndb7z7YlcBYqaH+7UYDh5ekDfHc+43Wn/AdeqUxPzWmLkO2
lBqa9ygCBPwFd3CA+i5lshGRPo8zMteHNdu+AI0nr0UmV1oBNyDtChmIpPzNYmKAaGRy9MZ99pny
ThRZZabAS1VGVFBZf9CLiIH9UhflA218RtGAApxDdE5011BKhD1Vk/QRBMUqINtYsKQHwTCF9EgM
HefABNmMCbDlwnBetQzHHFiFXZ2x7/2Fp3g+CcJs+eJtR774X2pM4ahgwzgxFh5wlXWG8UfC/XuG
DQZlUHN89JyWBmrrf8Yrm2078+IsnxZAlgDH9ME5B19A0N/r3c30ypJQCcKxZbLYu4SpKKxAWDf9
/otYBjutEc477rIAOe327K5qmsAybhef36DgNm5fdFP1u78WLzQQoJkzOtKfDZjHdyZ+GQRIfF8v
YDXPSA1hey+eJQbitHB1OJ4UPI3Ao4R/gI3uzKeeAUKYaEorVaVV4XLqcBYOo3FlF4D0r6rcsQv6
nVnaZ96iMx/SrB8uBki7PXOW8vX2sl+I+lRTSMi0rOirhKRLR2/eymijkHxScICPYumhVTeZRhYG
M/+H8h5StRaskLS1d/xfF5xBP3Lg/JHwYDirEmJE6Nc6R9+f3dPn0gfB9c9RLATVcX3YzDninHF+
I5QACmGiOpxb5Fm2Fk/KXJq8cU8VaxOQ1JsvBGoI8I+YVMhof3WjeJGAa7xMODZlxu0NnHDKqN5T
nXBDurSiuF+NwlSOMc2BqifxuC1M5gl7+v7fVoqz7+zNRj0c1MMxooaxGLLlpquITywxXo1S37es
LFYO68xLN3Wtycst6EBdcMUImjZsh0+OgJIL9FR2wR44hYnZ1Xrl8KiKK4QQZRPlwndEiZ/a0I0+
lpVIaXzTCX8P2CEO+s/RoJwE8ZlBmest7a69b8i61+aZB2a95AS2U7pPTcu/8pissm9O9Dx/tmMk
3Vpx+f4ecBmtbXZsbyYLy6qgTqKkJMvux4BPvILhbtN1Ugz5DzuHvPANmIvaNnZCnaWbLYUeSOwA
oSKl28vA5D2SDorgNJLW2x6JeHMWYmNTG7yalrjsg8lHHoKG12EJFSZwGxCy1hWxPxSiy+hwDqeQ
5OOhKebUXd7P5d7Z43gHXfpZUBwd2ZOFHvE34JaQWqneZoLSht+Ms1xDrYqnwQN9vQ7pPF0WheZ4
0Uwiz1uz8WVYILTfGIuRw16GNkiTiiHu314G5+L6cF9u/3ce9GFql+XWA3RTkffqa9IwNyat6Hok
baAdgzwfyoEHQe5c/iCW+o5WVlt0vcJvFN2LPLDXIemQdDEEIizt2q5Wz0jSR+R66JnDUtH8/u8g
/aJi8TFbZ5jUHVu4h9kcosja3BxzSfS1JGmOkV/BukPsWP3AdOPjFLDtL/fHseU5qMtwr3SQXN0d
NRWnITReNLBPUbdMinKGW8qnfsm433ZyDT41afc3djHgjQV87UAFuI9WpxSoPvu+74myjuBlt3U2
ks5uIo2+N9b2xhq0ZozpiQ6yXf2J2pgpQEPnkk+huRe0emvuF2qcVDMMHB0d9MWbDxgAqOaJiS+p
Ah2NDMfbFqDips0gNBR4mrGlVAaiAhSXgpZ7uE+syz9ZzfM5suaRxgOoi75A5xy7+KbDmo8Ib+gP
wiR1kgt+Wx1YmEdre0KheUmAMhQbaMQltTipaCMhsydJ9MN/1LUoYhZ+pccsAzZ6VnZJCdOpuYfJ
l8hN8Q6uvdIkpNl/u+0tI69JaAHdEn83DBL/gYQtYkKewYZB46v35Y8HMlrCfnE7pdEy9OFPJsY4
Ud3E8WF9+5Fbgg7e1S1G/g6pvPsAWUJCP2MxSgi0FYb+H1Gb4NNYV/M71Mo3LrTvIY7Ogd0KqEh4
d9Hoq9XyaQ2BqACj+DQLNYsN58gAbR0CJ3WURnyHwD8r2d3V8TMWmvmaIL7EMPkKcBYLqPIForVl
q7tRD6PqqLfEHRG1AJLtekdJcH+yDFZ4XejrSN41vP7cxaJOTn5nl/6L4lbabMsrVxV0Xx+uJ+/X
W0BCtCXfFde0LecRisKVGTQ8g/6bZIaKbFuQhxOWqbp/xnGnQKoO/EEQ7LBa4WEmlYFDLEZlG+WT
0VI7ijIUvjxn3Sv6t4f61vGHiJhIa8QhRer27c0pGWGXtMTJjc9Uuu3nHDYcozKnyv0YnZ0PXbyA
6RZKPahOlGVXJV5cmJ/9Egr1TgG1p1+L09gxDQKfdlyLMOYHxHUFYCo8BaLZ9OCyvPA0RF6GBP0b
MGBTLLmr7SQOnTgcbLFdRbUCllr0yn5PgQyPpw2En6kpKKbQZPRbhn4RKKhaKx8LmR2A6Vfi8QAL
Fo0fNECWlILdLn0zUbB/KioIvazXwPNygwkoZk6twbt0+atjSyq3rk6RqHbgPAQr7c9LHoUpTFmy
rMMJ/LgMoM+akfnwVxe8rnGynrDZTc/KeugrCrpecF8iMGrAR6Q9X3bLvhUWqOg5O0jfV6qLf0lV
NJH1rw1DA1wrRKpmsnlWe8NibTAoyKQHi3GD/9yExJH7mf76tkO4wS37MsA5pgRYuUn3xbI6qnPY
Yg5r26zFbBuGnOWZnsXBiXVocPPp6AmwW23H6a4iKH8D+OsFXS1JGR9MS9yG35NELo1EbttqHOMm
9OmgD8K+Di1XPFA8RoS1B8hCeRW1/PNGdDNGk6/PWWKH7xCh9tMPcrqGMFEBu9krmWPIDWZVIfcg
ZLkitB/5MpbLHLAs7SNiwzysq3KBFT8CP43e115g+cYtoeit78izFxDKI3uLQNXBbTpNCarFT70W
INmsKHTGShODb75h13onhNQ1pj+oeBWzgl4mBQyly3czsbyt46aLPmdSLhmyOREuVvUGfng97Th7
8d50U8e8aK1nu7BdfSjKY2NcSKhPO1h/E+9xExuY+WXyEK3OhOeEPK7Ed6ltPeBodZ1S3BlMbOVF
MpdatnNicTk6a+k+Ntr419c0pFqS1RGYj9hcq83eWvfPtMGiG9/F9VQKXdWp1I3B7bNVycT+eVhl
lX33xgJ+3M+GO4P+a3VSUVfp79nO/4od5YuF3yuoQAEJyOKoWWwteiRjPGtiXiGB/kLwiz6xsjJ6
5ZszNmV4BNceRtzJfRuw8Xq/EdNSwPOqJS3BCMTmgdGmm2bTC0HgASPS2ImRO+p+v7JGZU4U7/QN
nUGZd4gHV2/rg/cfdUQfCCmp/JsFH+L3J+wxauuEIT6DHIToD0RC4jep3JrVoMc6eez5+trW9lWQ
7WnCQWXPetEkKb6FL2KGw0ULaQpdYc43pX9IvA33QtqOVFIhNQ6DlDVibl+6KgeC12gXlSFlmGNp
9C8QxfGFbawJDPP3xLW+Nsyl0MQQ4F+5OS3IJjapGs7GFzBO2+pc8Z/BhSvL4bXTtQAlLSpn0/EE
HO71hjwrBEkQZ1nDTjJEzkMhzPoA9hxxNQwLXxP9Ffj50ZgDcR6KaUILB/hioLrZZrAwkvfFwV9e
YdB5Pb6l6SQLffHTCHVDMOY9qs2c5X9Q2GBsQn8TQ04QFyO5k98FqkyGyXVh/mJUjdyuqKiJweCY
nX6C/7vG6UVH5PbVwiVW5WEDEUEIYNIist4HHdfvZtuYyU32I1yKESbiiiRV1/A70Wy8N1QUbZp+
34mQIkRusN8tx8qqMykWWYoK+49imOlRBFvFlCyaYqyAaMVWyBGxD70jZzQ5aDxH7sDhEj6ehc+l
aa0qx/daVzr4NH2DDq5pizq/uj06RavyAu+9LvNDAcPdC/3Di7KNu34amG9aHNv6+l0MPaf7OBMf
RCupublrzm76uPOwlTxqLUmPqPmIGSEvPHU0xOP47La67FTwCgz+7/rk6BuUY1nOIwunlTtLvO2X
m432rMturZGfv64jZO5kqopDwMfn5mv9vMmSUx2vbh0jU6/SLMPyRgiCLZjkjRFdtbZMT3UfnBj8
h8hV8bzIYGbrdRHYt+E95LhQectTvFYg63qvJLrRejFT30VJ8jvT6biybIiUJfdsSCghJ7x5XX/G
QNnCjHYC1J3TkX+lZSpd4brb5ty9EKD6wU2QTSRw59bzXuBgeh43m5YAMBDyfjwnwQHjdm04HxaH
VjUGHPGJVSo5GZwhbm1rs52QudqWJt1ktYt2almSqBG77024j9nloZzVQFk442HXFz+/xR/qBY+u
TdCXA2cNatlpZ4+5yii5kCZlE2U5TVq9Bd7rICx3aF7+yLO5+2RZtX4jtm/V8SpmyWVQcgTzug0e
cuSkppOkh5UHNAnwhJHMvjFAQIscqZ7STSx1zsuZbNAIHagM7Uq+GB2eTzK93UdRmGd+wFlYK+/m
GHzi5tqqJX+AJ9UkpUy/XjwS0v5i/UcH+l1FMXpTtaFNEppML35odrGIRfZuOdWC8kykAROctlrv
PCmlRANW1zToOGWLNtMDTLdK1lAM8UnrBx5uldyzTVZYGoPusIc7voF/MyxYMsXYT94t2MRkEyoV
YDoPHY3VPhNll53d3OKjTUZR7JU0HWLKacp5K8uhTbB1p/xSrmNWvCvnhPrnjNsEIK53cr9bHOHT
ukUBrGd5tSmhr3MjW8ylcZ8ul8mxGJxJHt5B4EqbyXgplBuqEnRp1Z809iDrKeDuqKs/KtAZ9h08
UK488ht6V/1jTa+pxHC8Bb7GUoeccZ8Grum80s+nRIarQz7Y2uqsh9Yv7fBBOhyd9mI4y7/Ros3P
AwtmDilzeYFOIhmkfG8i+2N7K6BOiETfYZInNn0PgH/emZIW0R7U/qyJa7UkwY0UJIU6uA6xZDwP
UQhmmmxuP3EO+/KR3kZhhZkfGyHoQxyd2mVvfcNw5tfM6gPJSC/+L9pdBaiBO13+6h/6gq88HV6X
NXGq58p17o+JRc2Ye1EZOBLU48Exy55lwJ2y7EDyjrql9dmPemFVJsZ7e0ipNm5xhmsbVUK3U3qB
Aj6c0SGnjt3v49KXWaQfhTDdlARm6yG/4UWTs501Zf3AQcT+gsjJ+Ci7zkYBls9WcbxRqkr8bym5
ZFkODS4nK7mqHDCOpLlWiZi4Wy8yTi6iYuVCLr/A88uAISqN39agMxUs8E5k6i8OxXuXUOnJEGuh
0WiIe4+aXIIjGeU8KpXjZbzF58aGs4OFDeAHltTVH3HxdvjEvEGVmiU+9bT7/yu7VQuK5fkobitV
PszCyyXibBTh0LcVWdbZy6I72Iq/FGf+71JXnOWyi9YInpEY1GQ2FFZY6n/xvtViDwIlsL11w+rl
FQ3rxOjdh3Z6KING7HTHyq6XRW1Yf1n8cHavjl/RaDJycXzYHzeUnDIIehYEX2+3ncBrgrQ550XS
jI9VVigUemzesVtx7tVLrcd/dE0c6x9XwM/MOjtmOgJBfKATEKKjSger0QH6qAvcMO2ta2d1X34I
fzbWZxqzLohT5doS2Ph1uy31y7Mukza0z36Vh/KiOk154Y4BN2EsULC0T7nVbT1Y2cCJPYVZ4zDB
WZsa6xQfR5hfSseQAALjScaM1bmD69omzcDORWUSJ7rDt4gAiDQOBFSyLjbrOxRRRoZ42F2GYMtS
ONgeY9k8IjfdUh0w2uPcz6NY18q7VjT7d9SmuMZL5xkD59pDcDKvq+DnZdOSWRErCZVnTsXwjpbd
T5b9uOGjJecmVlWJyrMhcJdqEOLHwUKtRy+t8PGkSVNxl2/RHiUP29VPpTMmECdF6hhrvMzkYa3g
AyPYxUbxhNW6BCU/ImpVS2Brhs8vfBwvP7NXcM3Heo9Qtm+DTdcy9e7mnT2A/pSBhy0M3sszTKqs
GUvqx2ilT1wIG/9aSIrvwv1Elff7HrbLIF41E6+8rTcH5hsJOkyekL3ftxh16GCgcwa2JRs2gZta
6bCpu+J9Qn8aGveZcXs3NrTPcaeHDUnZGpQugGxgDx3jvXCd35zN7ao9wB9R0+mqAsDCKjFbdV6C
Ek7h26FZWGNNsqBd/f5Ht/8+sVRO9D+zqdFxbr2FFLmL/MhYc4F7H9rKZS+XgbbAzjRsU81uvPXp
Drvxn/EhXzqIQHv6+4saJ1Mey6sMOAsl20VZRx7Zesb5XpAKq1/zuHcSs0D3ClKL4suH/3DouXoL
acgHHP9gNDxFQ0E35541i9cVDuV9WBetNKJeW1eHDbaTsjTfh155COnyzeeMxMAuVE6h7k8NSH8X
AecG7VSsxWifj/0FmRDaN6CzIXhaYZEH7C5QKGIXVpyi1NBGvvHktsItNnaeSzrpF8Rr7CWNRyms
xg+rsE599OJjKRwbNk9KFOQNLHqEhVlGeCEjS4fIryhIkTGUsPKSD2cIYJ/uKzIA9YibAJjV7xLf
W/lIovtyaHzK6g5e94vXSFwv9SQxFA+WKGfD9cYHOSP1PzaYni98mK3PcKIRWmx2RwLPeY0BkTbk
YmSB/QVkFPpTn14hxmW1E+CR7i7thrQMgrA8IW+T1MaFYdTh2QBNsqc21BHmq16KJp26WZJ2fHOs
P0H2tD/rsMNDrykqRtlRuJb6yNEj/82XlfcxPPm+1S4ltZec1UtIyQi6c8U9KBFr4ly93wTQm6yK
LiacVsrcX1ntxnKuZ9idhJ/wncvJATZnZ/YR1JP7a6VtzfAPUqBq6tZjOYXCbZfRiNvB7KgDfDUm
ns/xj+Ey9fe7YOavP/n8Jom5/twUFx0yG0y2aeCoYdJbFKVnLGZdRrinYDcIc69gc68FLOUCL5R0
UCjspKsY0n7Lgefb15JI4HhCqilfwErbPwSJvSlYYpvxpU1w1/VM9eMYghxP6HDQKpVgqfoMJuF+
K+LfnOxckoQ3O0nTSDgUaD467009oJTztZp47P3iIPySeyECmGkZTZtr6i5qro8ykhW9c805Cclu
2TmbTPjJPV+3b5voCgYdcNkv7SbWd4AJDAc9qkZu/9V/dn8GyUhHWgWrQ0yKmoixiSVI7E0s7/U4
jVCCumfkYO9Bz0CzfeWtQXLK9kDaPIoh3Ot389e0arq+5GiDAl4Ggs0SmZwNur3WiPhZt+v0/xOt
rkD0h2zgtNSoJ4iNrFUGI2FsgvNWR2GDhzzL41wVvEsNFaSnW3Thsn0No8eTG3M37kG8DHTmcx++
ji7bHUgB5xCUiI2u7AE7qq4fuDrH8kIQ7h6/jDVqjmH9lOMRcpOeMhX8lIb7Ian6qO2sYrk+g2D+
cZudmJSNql6RdkNdDUbtMoWQFSLJGsTfjyiT2+G0dflgMzqbRlcgwq5ZK1CCVlMSIdJW8IY6gmuU
3uBeTkDVcsJkWHdb7ym12awciM1qs5LFa7JGdnZAkNdMKZYEBw3x1xHppGLqwdDMF8ec2Q33NhRp
Pp7J0NOek7JG/H8TYBPKs9CneFbjvBzpXnRoOJW87q0zozZaLX4Spro39yvgEKt8yWKg350Osqbv
Kg8UVeAfROC5NmPQBLE/Uanq6PQD8jneEV7+8wZ6bYE3YBWe2PuZexwVXFQBW3zJJUDEWNCi7isV
SjsKhnZMhzgSZiBO5deXC7OZSBbsx0yd0iwAfSUTgitBY5syhF+tcuTm5qNImEV/jHkqIbuFSE1B
EGDoJoZaNEvTFLkpmbvTkE02tUjxW1/BdNMU4kZPdNKj8wxlFzwf9SCugqnYRzRQSkLjgdYYBJ2x
dhEH2QX2KJLrgAxANkJ++a2/PlJPJttPr0xCilzVyCJzJV0NWKewIFIBmz5HGLVjP3CC6E94oAlA
SIpFb5+Hrw6fmrjFE+UhxKn1C9zCs9VXq+T5zqoSg7xJRCl9SaRAzjJzySal9dwhcwPfvBT1Gxfy
mi9WBWL4QrrX2JNzKNTFz9jHvFwgT8jJORQsrCes1rGlHHMRqZ1OgzszTBnp4EC8BPxLcNa985kW
WNZB+0lGY6P2hqGYrNLLnh3tvmAkLa5wXySysOQNSf9LPnxuwqgcboQBCfxuJzKkV0f/3of127Tg
tHA8c3DovfFaGkUAFQplVLGKY0lLk92TjulF714J5Q695LyFYA+4At7+UiAHX77xWnocaSPfGDZn
ZuFuM99TXnGihuzyM9N1Fpl1WEHyRhi57YizBumBYcXavGA7ze0HDYaAz3Vbbbfv2oDKqGOlrYRK
AXVqn+4Zva7SYFv5aJqzNAHfQ0B6zAKhnzm3NP5znW7WhxlJ1ZEddp+sBxfvhBkGo2KhScgAyZOt
pZgANiCKPOkPApM3sjoggi3Lc3LETWYFw0qrj8Hiid4WXFIdkztK7eAY5YdDalZioCX7DYQ9ytaZ
umxgwsNjLX1i/LMUwAB4OB51LYLl2dEGdjcYzv9zYDKBpU6LNRXTNnQAlSL7C20FN3G3LInJEGlR
5uOhXPQLyeTommPhqM2t/KfbSXL3fu3UnJ+Qh0rWITZyOcCn/7rqYUuHGiUbvwngbfSnDn90KCN3
6zrHoWAdBBwt2IHWjFyzTbZvHU9jiBp4T7hrBiOfaWAFHl0QYAldqopXZ3YyNPLd5j/VHx8dTbz7
Y2fFefwZjaQPR4KIdCF0mY3DQIiKmcsDQUrpabzCvBguemaBIEhhWtCzjbdkhwgBoyvogqJjo76i
4lBmGAXUrmfWW2It+CXE1PbE3XMuCdf27fbhWGhsq2635eEY7KlvYzQF+Nama9pJqm/Rk4CHs5J5
mbs3CP7Q246JRiD2UNyZArMoLvN8ljL9Mf8tzUdm4wpWbfF/k7JmG2yCb6xFW213nttoA51QLBGS
p9iHshDNB4GOMzjdnFqfozkRo5xsN/aRUfuPN6mqCrBNr9678RC3ZT3SIA3NwQLK33HPj6z9XEI5
NgiX/TsVkGEn8oLj1Ooo07oaB3Qq6xEqSH6dd6JBF+AtYamPqI6AZYXQPaWQ4V97ITYRLdAh8T2h
SVb+NCefMmc1iYd6WxZn3GfGfWhme6etdUL8lQdSEf2C+Svfwcn1JBOLl4JF0WxH/9IzLz3xbq3q
j/A3AnnBfqhTYx5iE8UjVFM+SjQm0vqeV/OIM4Cef0+rjrx1NxRrEfkhsTlpQWovNI5zRgsJaHkl
cnz/lePByt7KfJYjglRThNosgPfLYJEChfV4b4VGos9tpvJ/3onFug7KUyxIGK+hG391iLvy48d6
nBrQLVnrf7IjDAd4vf4PyaJdc+Xi7wvKtLYULgu2nH7j2METiuEL8esyqIzUpeexlz+XNPRC8J6B
lbY923ol0uV4zvnXp1Magwu6dGkebz+OAAlXbowkoOncKty1QPBh4azH+q+YBlfLyXIyaccq7hr0
eAP97EvyOKVVPmSJ7v0Br5MXVXas0kX6kURB1kDXgROlqimlUby0WudItzsim237Vr7h71gpEXYR
wya5z5St0XnVdg75f6SwH81QR3qw7NDOsGQmYEJkF8g89gdeybXgMbWCv2OUQBjiFJO8hy1vUiwl
1yGVfvo1I3afRHVjHWCNAorQ3/NXX2KFuS4C5iUwlwM/12A7mrRtpkuS4eec7HrR1rCfvxuv1/vo
CZprQwW81uxom7wJ/Req1VHGPv9xCO/CMW9KTubUvCW7Sq1OzNsRPEM9tcuQ4MW5imsROt05IXk5
PZkS8g80/MRSnY6rh92oMuzbM+AlROvnO+g8nwAV8L4EXidg4vSZA2fj7IG0UuSBMO36bMHM7k4N
10nmOvKcu2xIc2BcNqJs+lfcsgCSxgVyTw22SPAmxr0sIVGKz7j+et/VJs9XHY4XfSIXVJoctk0Q
pAV6pCyJBLY1KOp2fHqNDts1Z8ERvsPLyKOf1Y6+Fe0ITU4KMrpDAOItz8FhKlDGv8iG+WPTEOon
0qWADDgnFHsLULxG1fU209Bvg5H1GHfwIoBmDycLV4oKG0ECu+meIV1+o0fJ+CPfIenkgbOn5pX3
iqsrAaXI3V/zSp4aCJoIBvo9DoJxmEJL//V3MKhcUqjHiWUiTdA6RnBxa9UouikIW4ratKxx8LwY
Q4Ryz00NINQMc/oeWpJsbU/OrdLt4dtVR4FRi5eLeiBepeYseSEIiRbp5vq0aYMWg9DfjxGnv5Qu
nUdA3NqcMN9JfKBzmtgy7tmCWyZ1tlLRpV0vneuMdN5pGrE490cQIM3myIkpn8cmkcCnxtV/KLcX
JBK2G+rIAa7jbXvHCj7UWHJMSSJv4TR+kE1esPtS4x3CXXg693Zg087z0Vd4JbeDa6RmNYh8vMX8
DmMLeaOSEoUxFPRI4NpFH0saJx4omEKxJI+qc+LuL4YLOfQr/Itn50zfVY7goqHvfRBPC8fdZmsq
a26y6I8WjCpZdxfEDZcBZ2sVrwqm2xJtGn3y9vKm526V/QUBxxp5M8QaXkTVGauzzmPEn4NMQQP0
bDlvcdnJ3ozxB52ljij8w60g6ACqV3+cyvmMKvhBkuu4hI7Zw1BTV5bKxBNDZzY+5Bt1EpeVr3Cf
pFpjks/FtKF7P3nnNU6CBIUA26TTaidjYoEVXC6fc2jcyAuflYKE+mm5VK09ZUqjCh21h4UECm4q
2oMci4+Hvvhw9PJydb8nLVPGwXLB7jsM4FqUfy3VOsmDiDk1W8jM0YT1NMWAnHKGxN1itb7w/FCL
tsyn7HTr9au4+V3946NqyvEZil4WLur4Z2gFJu5gf4N2UOfFULaa3jc8T3rMW3Vxk0QfOHsblb7O
xbzDG4W/Z4IOJRu/5TejbASJJdMNJVchnLjUTmSDL/6ajW6koCCpFJOjvSG4/1poSK5AVJg3hIbh
/PZCjriMWd6xgWbVW0lur2uSTtZJuV6DzzcU/bRZNsI53bc4lYNjTP1f/65T4O4+uuKCr3fKV+fn
p9hVMykRorI/lQ7nEdKrwkPf5OHc5MLqR8VFJpFRrmRowB8oeb6sI1jjyFGNtVS7R5cikl3HnAdO
qCqY8fOwT0PAxytBT1FaOEW9TmA1D/00FbOfHP7itopxMc4usuP4lGBycCCJeJMLzFZ0V0RRJSsw
5z4UCHddSlYiriGLnO0ogu1BwjY4fA4eRsUHR6+immq4T2Q4qSsnWIFCWYa+sru3MUQConK3di9+
pAB55RjNB3MUV38PrdCCLI7h/F/hB4nvo2DoXfc/6sldw8aH6ia+frMDEmg+Cec2ZVwJ271TqHDo
dsVp7YuY3j1Jl8bpKNwFdP+k363NATJePytpo3tA1YUO95tWVCwhaYceBg1EU/1u+YK+vZCl5djY
OgVBhBQ+qx1UQbVAH2Et1Pa868bnmM0Gmntr7Vzs7NtsWpY0zekf87tZ/grO0XJTHGqeSmH6MMDJ
DMKgqT8Hgf0vUWGME9vWygOYIOdkypYOMwOxQ6MGnXlaze0TwI0J2tsvxKmlkh9QtqK65Gs8YofM
kCj5dADE45BZ4/B3EeLkTcG3WDue9J65qHwujme5QoywvZIQlHCE7gArNuwKaRxGvVwUwdg9DV4i
+Rgcehy3HPacTHjUYktCCm2ku6o1EMR2NpEmfATUdp2e79N36dAbV2kDhh7OVwmTmZD3QsO6bBa9
SkXkx+/oS6PuLapQU9bQeaianZzfPdxGqKGQAHrS880kJjizd2Pdxpq1n3xxzrSI62bUmjUUxxu+
MdrTt1/e0ZVdli7vx0CqiGNWbrAah5TwgL37oEEIVNtXSxkv1M59c9DzaUuxQplLKufNzGt2uD9I
Yd/VlSytCixAqcHyvlvHBqbpDOBXX3hnk2jZ+R7l9T+Oe9j7j22btbGmKAj1BBtOwMGY194gFPOY
vF2bKsmXqS8txXGXy1dGSOAcwBrED2IoqFFywYf0CVWBkTuwCzUHcVvOd48caM1DXiKpphRxJIyy
Aim/3ItjTUlM3fluud9AOheaBGhJ+4ndAoPcW0oeAKPsSkN6kZX8aUWocJxeObib3J//qh8/5rAQ
7nHRvV5XM0qK0rdVHuhHd5fwINY9iqj53BZz9xeI9Fap4bmCNL3rpfH7MMEfrG5b3gy+PmvjVgqb
YxexrxPNCB9QQgKtmI4GJIe1KkheA3Xpmp5cYQUCaG0g3mYu9LZqG/hur5bYW6kqZ/mP7NGiKbpU
sk+pBASJTU6/GpOXdlGhqwYiIZi6vxhxaKv+8BkdF2zt9gqpj2OcAAsUDJIkFuDJOviQZHMJl1hL
Ij7ZwzVsu4N06h22mrbtcLWjztN+4ergAa+mDmC25rRhFOEKGoQPwmLIJ4n5kblioaOBleUDwN7F
4lrYZYNbHDVhzzG2YO4NICtPcXGbP/Wrdn+DjVUq+5oWMjYOZngXBoWug4TYtqlvkIbc2MxvoPDM
Sed+4cnnYSLoIAMpiaYsAcj5zSa38FnnD1yxmq1pxKkXdYt0O0PagsPCf84wY7CSipsjTL5rWi8J
J1CLWp+vI3a6EupDZumjK9uvSqBVuf7kWWUi2clf1b1dbgVLEFP6Twx0YZwOco8M0SBxH24nWCvR
VqdAcPtYcRwUtcKPDaUwBpUCBLIgqNL6TlspJvP2ZsUuri+dSOQEcqoMcnI5hExIVxvo4IDO+PSD
tZl7S5YuAV7xzDuH/v18VXn0Q2KD8N/49pjWu76EJTeFnjJU3LcaaFrq7cfPQCk/jaXtj6zm6QW4
tpVwwPXYf8UwQ5qpjFNWivheLPPU+dOvA2bAJY1913QsPqT0KDOIFstCbyfXR28ClSX4GVY0d+0T
1t6xtUcwO/XjtfNELYbw9p+iWkhAp0DdYC1K0vyl1bowWHvC5NMiIeZEWMY4EK7FC43bTCHHNzdL
V/W9y5+vy/h5k0uQlu3nii/VljMN9zcA3i0jscgDLs4YKgaYwsbfY7ejJXJS4XNagjb/W2wKmGSQ
DL4Ahxbp8rQTqkSkNFYOqo1XUchNQHjItafllq88iP6oMPowO/YHlfXZyic8t9emzqLw4W0wy2RE
gjesPYyAOUAlSspXAf8s/PZ7z3hnz6DZeeVvP0QWDdvMkNSkaE8241gxHwza6zNW+unmzA4zMETK
E3fk2g7XweHoitUnc5h1oPj50QUXtYDFwRWXPAPFR5SH1lGSvwx4WBy5BZuU6NGS4Rjmt15L8+I+
ZZuyYiuCn4sJP0gAYhYKH3dbR2Obh9RHQWZsGQk1JcxbBtzWuJjD+ktg2KEVr4JOKvIaoWAHXSmd
lQi0hRSVDgf7x1oRDNMG8zEDi7Y/Tl6hKAxTfDWAG40CLOSyR5cLeq33G5xSsG82GBKJ0VnVvdht
ULG2BAsNsIi1vaupTjUamvUlgc4phICPlk1y40MjTKXJsa8TVmZONysRbx2oiXGn5hQ9CkVkR19J
yAoNd/BSLxBFvpNWusUukr5qRQQiPkEVBakteM5RBTYYaRkGL5u58tSJkUv5TNgpB7b7ka3siWHV
23vS4tCpxbDywPEvyw1uSG2VRcZwjkiuVyQ27ubdGUAJI0szuEvwcy+e5JgZ4bAXehfVegKLHEDC
PfGbqCZ36pbKEYvBy0s99UoxExg6K2HOLdQyOZrDEtoX6uxDOlJssfnbzOrPa4GgD+4UnM7KS7cp
W7tSql55NwZkJnylb0ZaUL0G/n3BXJUV3IOafpVWgjw3W9KbUoNUnz5BIf+64DTv0Bb5bwHQO0DY
7e6Zj5zAevuP/Oix3JpaSj3DAUguFFjLKwT40ptdcss+ZMsnUcLTWa2GSZg3OZCR94Lx702VMyqN
pV7/bEKBauQJ2sGv5fivJNiTFQumqe9v25YvhYkZSD+J6MA+Q3OifAY9GjeFJ8hz0rqgdCCwjVmf
5etmfEhoH4h2U6jhnhvFhhxPiWug82xanukccocrUlOTxGTSffdBAqZ37pWqA4tgesSUvq92Wcou
qEpAUrfoeyhV3ErTOCRP9H4K47ISDu2AN6KKF6sc/xtW1jiYCofWzRJJiOoFWOHdXHghdQsyf9bg
sT++n54c4U6atvv+rhTgbvJsYxr03YpYaaQpiWHPFxOAEuQYgLEBZRG05FhapoDeImBvHD07ba2+
T5BsSJmhflHAkCcqCtlsJLy9QmUQEl1cOBRhVGWhrlsQMaPhS7Na4/z/ADwDAj6T44EjfopK+2tJ
gR2wn/mfKvj88p3SwzPboM6peNk23jJ7tilJlT5ZRV58s0SB2Nu4l7V/OAzqf/WgCcog/9W8N8Ls
uhaccnShW9dRImhjkQumVFwInTBbUdz4achzzDKFmDpXPkQt85mcfj5BCxjthZUamjvkiy9ZuORF
Oi35BOo7ERXL9CPQ0QOFFNc0QT3aW8q7ZyFIXXwemLVT+4IHME0s/ZNdYvCmevICFIV7AABwB8bV
2BN5xpoxQ2XCtfjte/M6UIXMgQnJUZYeeWaH+9iuPubjklsdd+wiZDrF4c3+V0uBFMuWy2rzgpjv
nSRwWM6YNC0sakICuBKnHgCQrxK4FwrAF8xagmrb2BTKvK/eY64bM1Amvux6dEE3o/oZ6nRw9o5V
laMAueREkTKled8q5KRGoTfpdwy1+Iz6NT9hTsM6Nxtz786dxF1zBQMfKMzawZRur8VHBDmvq8AB
hZVjhYiYHSdrafYOXIAI/QPKY1+HC0XFTbIVONeAi+RK/0ZRby1RYrwZfeJx5Nc7oFwkU4RD4atd
T/l2iDbYMwDjkOMXT8ON59LmG7B1C1BK8yDKvtT8KMi9dIl9q7X6r0njdrH6ToTyjJXInUMrtC70
kC8+ZkqfIZ6xzE7M0TVcL2VEKkLzVXRtKt7Wv1Z81Zm2tztWiNgMPJJiMLMjbcvoKPTFAw0Fhb1h
IFjDoO0FqTst5LhPPGO42t5fH9H90Mh2bmWUpTwuu0wha9ZSJy6PSs7oNRFzapQDyJQ9tQYOGZ3i
0almBGahodqfLjQxCsC6DxR6QOkpnPLrlybrjVWeombR/vrTPzKwsQv0DFSpreFVHH+npgEjabY5
ukx7vfMgVhnsn9svSw8/OpvZhFPsFRNg66xsw5wWp0jIbGOdVMx7mI2q7Y9rv1k2XR45Wzz25qJJ
WLYBA2KFtDsMGIjRri8ahY5ZPuSr1utr6VHxyZuhHyB/n4glkKoCjNWLPGRY3sG/7XfcMrx4FDtm
lnV56VxDaqwmE60KTmsl+ZmuEGbh7VaAUXUnxB03BuBN/uEzyyT+2SWfCZMw1h96IGb8o9wAfbYh
TbH5re0IWWUk9gbrPXKZmF6yAE0xAcq0lxlZHw/6o85uRSxnhfRwbZJpHwrvQbDrKmCZ7J+uGVEL
U4FB7+UVGXqQoGAsBvLNehYMuTXMfPvk+ZRtCwrXVOcSkDKQrBdc6c0OJRCm8XDdAKOt3Gjb/R/7
wxxS47ycP5fxN/Vk+0bk9ygTmB/mDeAiEYPaPScYpbfgarFnJ4zzUv+7BMAcXwmnykTQDe8i+BeL
XjVZ6BRwNmUACRxQvU4lMAqVjIPyZ+i19YtkGtZVor11j/ENCsZUH8RTL4vwILsWLKUdcVuvqIme
cppWdILR8rucJU52vi479wvZVCjlWIUEqTpwVFCH+NJifzcgyEUCD+RNEyONrI0xHOrPt+C96zPJ
DITOvA5ogrCiOEW6Lazx9jMk0xNvOpxfgavgBR3+lKMNz9zDyMkU79TWApEKnVqKyfD5dVqv1y8k
NsFOGdbtRLreNVJWwX69DJdO5NUgvHLNmqR8dxLl9b7mLMMADZ19sKcy6xroWqdMZ/5AL3O6SDnY
w/lNJSTZR8BK6POeBqIIdznuKZADA6vR/Qgik1nWB/3EHCtFK1Q4Fy3K1nUYfXeWw5Hf9OSku4Aa
NXYNkI64enUf9LEm4uLdAU3Jw4knXPcF9e9rduiFAuzR+aTOBX4iv0NAbDDzXto7RMc7zuXOQJZo
nuZGa3kXMXX6oSQWFm4Shfw1AjBmSB1rodZefRluz0FE2oVHyDBWBJ427XHaUBdq28bA6QT9M4YY
CtigOcNwMGDsLPWZb84m22h4SxfYptzYa+unxUUaRwf0+ec2fMJQMpJtdgVl92rOTZu7/60ukmEa
NK2dllvV046lRrcTWaT1ZGA7GnR+NFuyvXk+13FbUgPRTenn3Nnk/8UQNdneuJBs7gZZes8rrR5v
sowHL8WnjenZ5ozfNd6WkPv3ONEid9n8eZ3XtrdqBsdwiT4UBV78vudn5yjd8mAbiRxsQOI6n9U/
daWsJy0I9rJVlqsG/tn8Q0FQ6FWdAsvwZHp0LREtIh6rbVf0v9yoLyvNwxle7G6rZHR377Kn3sLp
EbDwru67mlga3HKzzbzAZHRz/riUyDebA2w1Ld/M2UGn0Vlt8q6T5WVraIEGoE7qqYtZyHp4otoq
OcDIFa/uKJcBRk/d2ZJ2bWr6VWboEDGXKvAJ5qg2AD75Wy+IeZFcAUupZlkCUWKHAi99QWd7HhvK
eohkfqYY+2yP+004SNQpqGJivubpWBWQYNV+CfEha4i0tWczAcVTi8NYkM30cGPs4tjGrGzuUnL+
oD5Inf/2rz3BCsnpuGcdafKsjFutGiels7h+itCR3PMvmzij5UES4C+iwv4NEDZBOVeaaFOfYUXj
kKmlS5Wqa0L8urFnDLiqc0OCycKhVQzmA2/sZXvKEFic0f26kE6PL2neXJHaZImEk65rt1+cxIyC
/0lraAJ6KINO0Oo6zdzVbqQcbsJrX43GSG9Ljb2IbRfljTFghbfmvQPjKpGVAm4f6dAKPi2Qvd5l
Q6oOFVXg3CgcyMSP7qQ3uN9vjWsn+hXh0vWsXek445DHBnBn//BRaIa6YCWdxsI0EDNCOvfW15am
GYYNTuvCJj51vqM39xQzbl6Y+CW5Fx8uxxOQWi8VLkObpUoomJD+AgsDc3UccdZ6md5jfGPBzeqI
n+vxH+8rvsBwKvTh6eZYvlMl6aZBKhAJj84ZovD2R/dkK5XANxa4txwH5aIBHIA0hOCBi+opN+T+
TXbu8By6xXIr3fjx3bFv/0yzXfP6kqvxzpDOiqtXS9AZvvCHH2H/NyxbAXXVv5JnpAKgmpX3a4Gl
GOm7hTPt4LlcmuShi/wKV7k3xfKZ73ACiHnMtkXRZT4L5zc926+pG4jmZs7fvW+ja+KDa2ouUX91
NVpqzPR2EmxissaKRmQx4jbxVSaTPfOGndnLw6NwjIAo87x6mYMC3475Ruo4I+oDD/1c//PL5ign
GNoaTmn1bl5/WmYrEwlhzDD68j19t7d3kA/ILseEbtA55X0dkHNEKACEfC9Yz/lzAhzyY01g5uJ6
+7leeTtvFnwWSgpzDbDyfZOGn/J1nt21hFl+XnfkKgksgwSypyC25KFwC9HGJLpZKJPSvbZN3fWM
jz/Q8ic2bppy+FxoqeB0e1SyimUA469qRxuV+Rmfab4pZBb3JWM9owW1MzOQYO9KsRwBjuvlauDn
eQj3ZGGRuf+h1Foip+HGwT+Hmx1Zv0Pgb5kErKfpRg3DqGQLbPYHjStWaOMDFKLkyYGxamcrlKzn
uOPPRN2NPPsZeQRtxdBNBwdzlVvfTWXxMO/8L/QKMxBNPCjfgSJAKWPG6mEnDFLK75Xw7Oc/K/VF
IJnqw5pKWZo3KcBr7Q31I2jO7bfx1RfjWt0lozdqB6sBlY/BeK7RvjYxKsxGP3tKi500HpaYFae+
2Zy/D6axIK3cBe+wyu52SrkhjDjBYVSGgZyN7HUznvxVmK8xVdsQNQPjwgke5UVr9HkR/Zv6lMS6
127SBvG9Panj2LOvIV6Dfn2kcJH7JkWskKNSfNMd5e3KgZYch9/Tuv5fB/Xq8zRzVIRIRL8n6dby
b/Q+AfCGlHFJRgr+OAE5tVeU1BTNbiaezfMCZHQNJjKIHSBrzjORj9Xe3yVbc04uH4cg8t5hGfdP
t9cCFvfQ796AjxRzDBFGlnc25lFa7mEl7K2QnMmxk7jVjmensEel2CrkYsrtT5TeyNNB/pFkxtN6
o+1CaHWhIfQ1l3/FCbqYxRkWJ+A1oaPJXT1RxmkwtIdssZdsIexz51xSTEZnMdpneZnn0Jrovx77
sJVzVTJMeHGc5GIv1gqXfR55ov4gUTmV03c47b01YbsLzgajxSHUsFXZcEcaeysRJD8o4IARl/6g
FbUl2xzu6xd4GN+MWJnRmP/LW5aSCp3+8yX2iaH9MTdPHQnuEkazPVDJQxGq+EfncIcdOxka6pgy
Vwmiwi9Z8LfnlvzfzUHHhQ5vq7VuIAjRLN9bQFDbTnGcTOvewe+lNzxAYyhd7ZvnZEvr7uojAfjj
pj2hh0w9zZb/D6R6iHSJEAG2I83uMNHiy/V6MoijWNuUHA7edUZZamHq+cGnAxuYYhdzcCrhSr2X
S/a21N+IPJNrHt+24VhzaVl0my935AFqESDorKGlxfLwOOHgMR3nYojrwhxZ5uU5f1wvR+WMpsZF
N6xHI/puqfFlHAV6eePAI/RlGIsowCfDhbz4j3X37kWemuw0ZoCmpdxm4bY67JvW5m/Hba21OJoo
JgZ4GrCvETd5DYm4AGgt91VkoJ6p1+r4YLczrHRU4r3d1Lx5V6oi1r+kwRLK/7KzUAZfxVKneuC1
fzr2JepWsQparOd1RhdWLUPtWDX1HTWsip4dGCirEKzxx9dwuQnjeUOHIeU+vRIiNz0GlzUU8wph
bjS9UOxFKbkVvO8wEQpK3ukxhBjL+1XYD4NvKJ9vuBvwLVxS+rLW4TIBVsS33ksu70JXn4kyX4AK
7ZGK3ARHyE0bwk7AwVr30Ri1LvzdLOi6piTn3aO2fU2/1Np2Pdo4tgX55jsIuIZ6oCzQTA93mjcK
yFNJaD4qE52mK1MrydouBhp/8fEH8US4dB3vZHaDXmF//Na60n++lxtPWx7/If9aJ/toDUUwp9IH
LDI5RyG01XBBw0kM7/K3mwDldt3e0kVL8qlwHnOMebzc29XlzGXunUTJNlaXc4RulxMKUdv/gNqp
mQiyM/FgIHWoUTCr6blwTNrsUfXzwjLbA9NqgeUCNlm2VS5Tw1Cxd6uCWPs4TVswIVzFCmyawaJi
ETw7fiL8McGYFD3uv9YNE9q06Zy65E+qqdgySQi2QBbNjoBxa5hcNittRazBvG5F1VHYE37OHrDm
t95TLtxOcKlDp6+5hqFORM+Am3+ICu1/QKCW658SdI/q8qvzo0VgQVTIplxpSncHmRvucd29ySEJ
mh8QxHD7Q7q0s3mxmyEiqimcUe2cdicBDUQJxu/OIZHQqgP4d9OE2CmvQYbZh+FC9Kwd7+aHtNvq
KJvlNKsxPxp+/oLGysAifcRX74Cw7xqCD+C4G2a0VwjHuip+le0TpUE+6FqqWbY6ZhCKKQrfq5ok
S7JzAcQdSy5eQtVEgyLk3ZeTWelw3HMj8IPSxQ6vHYhBPjFu63N8qe5dfGtLTKGKOPZtG75jItWj
10KZc6DrU+ihhay05GgoXB2FglxQO54o/hRvIobDqoWGKw+maoGpmHJW6vw+uv3/prK87hASJH5x
y83AceLg1u/q5QqTVVHFBMELm/qG+Rdcei7Yeqtsrc+P0E0AziCjBZA0gBhohIJKQIzAWMSAhrSM
0gss0daO4MlCFsrLbmaqL/XIAXwEScbXHld85wre+zbhE7fCFEU3lnd2t7pfjHGZgtQ4gDAn1Wgh
gJ95R9CY1oEGYIYW2zppaA9YQj3mmHikmmO0z+Mpkvs8LbJDgPXqUp8Op/GAVGR9g7UzabJZGDaw
Rzyr6h0zKH4rZNn8LQdgEwsUPelLb7lmuiuFNcwvOvDRvLIIQhb3R4jyFZSlGtpnh53hnM6ML89t
QIb5U26HsTgpIp5wmmYCzyfGwP4iaA5Nmlv9y3lo4OFhoIcHKZd0Qc4z2tw7WU407EihqARBUB4W
A5UNR/gJF/I9s+u6G/GNlotJhMlAYRn9rWxL7nZOzDTgY+em4FhetXIl+vZ+aabOeO9OdxDTHWgz
dALqE1SZmSxqq+jQBLj21HvORbN8CuB08GLw52eN6tPEZx9GV54jG3IhpjdFbrChMRhCjV9etBsE
XKG6CliA1O+kw/jI1l8JJh0e4eLvp02JS2HoGFBxdgh100GxNM9SGx2V8vKemIFY+E412A7dNbPr
VvQWOEavUBOx4PxI+bx27QfDAVLDzIOOH+B+FqdBwbYqfjbOlpigG5S6iEZiGD+pWdJ5fagqSnU8
KcCJ9UQNXc9yBNps5FR0Ru1qBY+d2gcRZJ/03XE5GEmKE2k/QCvFZcgeUI1rKpF0ifXV22COXCW9
OuYPmdkO04h8j1gRVJrbgPi5XzFPzfnj9SbT/lQnrmU9ctHCwujr88yNOhRlvr6BgH+ZL3WnR7Tw
CQ9XvmEpIwy2kCBe9A6Ghpf6BToB8UJ5aTvxkHlqPJXm6OnDMBxwWDbvTbleuj8H+OSaOZFBxx6w
0nMX837qy6oS1YyseDrifvZvI5zgPstXxCWfQr71Ti8vkSjfBldJZIQbm9ueYl6hlhBOqlY0ZQRS
OCUn1K5qvsGxAC3ci+9SufqG6lfnZPs0aUKYzBHK1O4DgJwcGMOJlHGi6LKSkCfwGuM1uHVS2YwY
CuKSs9iXyulThQGUqzgBIvNe+nJV4J3B5YWH3MNEKTL6oUoyGdZC1zlLqBTIb3aYF/+OsUEDHGzG
9hyHc0sSh95jSY7zADLcVKOHvWtiyOR3EVMDXh0sqzO7BSWtkyE+rvyTlOrrV/7Uu3FUZYWKnHDk
EOmlYGpNhxzw8lJzlAwd0PgcmiAafdcl0x/fXcyZeEAtMt33WlJ0WyzhSvbvaubT7RZFSzCrZ69K
5QXpb8bjQ1gH0BFbBqJeUuZe/IXR5l/uXtxBPtivmiGoERYSoncTzwlOMFbnDCY9lNOH6KwbiNYp
qcRzi1lpLCvCU51DuH8B8/x4ec0oHQklTd2O2c/3u7LgkcKIuORwe56qv/cX+ps45O9AwdCQWs/s
ip9/vsm2sOS5cgPJHey402H4VVp3S2j6wqkcZoITUOSXRnMuHbpRVtoWC5kalfpitvT1mGWLSaBN
nW/qFhaH8m3vzRiLw1tMXXIQhHXSfDxQQ0tJ942mgt/SUfXbVbDt5kqdlLxKqMXC0p96V1ZYfjrw
+NhQ3gbu9shzhbUTPdQ/7oszHNH/5dHR3CV3+Uk840rEIgTM3ZdplBcNz+8P4S4HJBCzv5PYw/i4
AxXPXLUitx2Rg2/q0+UNJmfm/mEXBsgM5AE+rbFj6LEN3R+uyutko6f10a9SPKjlfgwx/Nz+7Xvl
R6yrUsWYmtQ6kbeSc/zoOCUWQQ2vSem6NK+VTvrVEz4OI0RI39UzdK8tgYs4FWfrZOcvXBSZtRRd
0lKKE3eyhdUDcOegzmEx6tbu7jVW4tIGPN0ZHtyVsQksQpBF5xPK9toYfkxQC6xBPi7lp+gmki2J
L7dA25DWaNuhFbh7Vw2mXw3WuXmtzmCma7ENPqRiVrqtiPTxhIMxtnjE540BV17vxodSQSQZJLK4
YUQ9x+BG/4mi/0f7gUByV3t5cItSwqe4ndIdQrdThcXdVPaEyjxPPe75FPgpdzaZ9MeoOqbJGEV9
WxGlkZWVlkfCfAtTkK7JqaEIOCZ7v8Rnom+UzSS9luIvevOzkUpuZUm2SDPEtIREi2rZ6/rSI727
9vGdc1/E61jQbrg7VJZN8cZx5qhG9Ug3CKHmWAvF+HF2HgbWOj7pBOENM59J1O2RDVlqY3W5cf0X
iFFxq/DQRU+by78BHwWsqAs/TZ+hMZoO+I9LNtfanKFfpr4fmf6N9nBcD4ct41KN9HayARt0VtzG
4K5Qslbj0thQVXDz9KboZ9Ox0wxyhT77bxaML3lAmVbBXSnicgWBE/ZxcpkGBRyQo2ZhnBM4tbjt
9/KzYCjjng+qwBZkGk2IsECvve8c5pYFPfUvWmoVvbM52ocpaVk8QKQvq/UoN8zhwIZujqi7y209
i5CZ8SN2NbVWvRRomhkB3VpUVMI7BYlzSwfteZm7APaU9eAMGx6r47qCXDEj7q1/7ZviI0+pvfAM
A6UtrrKpms2bfkb1cYWTOaAQ4oJJB9ns1u8zM/rOJpw+sIuOKNpAixeMAvowg/YSPu9pV4XQIpOG
vdomgdJlyij3bZWLAArpW7c8XtH+aQiDBy0onTlxNc86fsO1g75+HfoeiizAOWNwcJQNBsn8wJQS
BKUZFiOHoChj11TBuGIow5bwsHOsNa9v1Ds4VGMUxMnr6Z1Eo754DyEutT5qkdseHwcG0f9DTgQu
Zsua3/LjobhapFkhysxi3gpeQkp/8+AeAvLSVZNPC435m7AIgvykc6Q1c+luvaRDMJ/343NHpDr1
FQTja1rlbKUMFDmrNg58Uf0ulVdS9YfivkFkfgY0sNJ+zdBh1ao+xa3sufGdXw6K5vlWVuAXUcL0
SZ3TB0bf+RPjW05hbRMDd7CJksq+l0lcUK9n/VI3ZA2pfTFMHu8y6mpGslSWNvSRjE7GJla0IQ+c
xOAe2W3bA8PYoAyWbCu3xLeT397g3decct9mnX4FHCqdRzJcq6nOH7sA7/MJv72vffYOP0NSvyvp
qi6/Z/ubqhfZO0pkdER6/XRibpqFIrNFEghdtD9Evk7NFJjsmmRDwXvglgdGvSfoKmE1fsUhtA3t
YJeQ2TJUiEnVEg7eKG/3rFGa373S2frAMVV49eA+uDO1tuZwVuqfO43Wf/6QDZEUGRSvMz6ZHTaI
2HCbFUP45L5wghPlrQ0Mv7XY6i9oh118KhrIO/rbzP18ni8D3swwCx8mTicgBvvHfGfDxZ9SwYr/
l6ePs79pbbFjORT/xBDOoRKBZx/ufGNK0YLj+s+ni8G1esVtk6+IxhOSb8zmXhHHjvnwfCptgvv1
h4pk7DmiVxzAtvzZsP02v7p15SIFnZoMno7C6NxhWj9tiqEmK+GGmdDW+1kD6P9pAY8k69LiY9G8
js47VGUXjrSyblZrQQq7MsKYHeh9fb+WExw4RDEovzIqye6kVA3SO8t55rrFfrVORZU8oXUwqRjy
+hRzBnamYthEeJ9oxCom/mHKfhTumiLCy0/89W0HWr8oVobM68im+wxj3HOyZxEnlIYIKZAwRJjk
4DX723dRKUCkDqK1OXQ84sqavYeMP0LfOQ5vI+zaewZllp0YzRLSZnA8tEbjO/sl0cKaKRtjFoz5
sccsIlCXo5ljoXWRSCaJ3xPd36aI6wymV/uU9Tm66Za6gdIlLCTcu9FcSvQSYXTqPp3Dpzx2Kj1v
UvDDACT/4mAyXIHok6qUvkVzcfq1YWPMsrsp7n8Vj0BDwbbayPH8ZzUjGjUmAaZyzceX7xrRGPNA
n0uNTR3J6muNEkwAA6RAyxnJRojPOjdhvaYX+MyvFrNcHAUIEKC4/51O74Vw7jZXalAIdE86f5+C
V36GZc6cs6MU0u3WxeBo2YdGH87DO4vQa5FyhWP+RUk+pwOXR0uqzHXxt25iciHZxNaAg2/SvLlp
ADtWeZrqNg1cK2cTB3DOysoTgFgVLsNlZ9yrQmYtRacN10C6lOb7/WB6MqJM4ScgVtrmiDa+oijF
sE6XtnhfISNbUH4KcfC9/SjHAn12zKj+tY8MfgynxjIrH3T1N4oO8wcIN5uyffCjr3zrz6qLflak
F6NlS/HlR/+7OX1hYw8JySiqNXsY36UAVvz87ayjKfM1GlTbqDb6Hcf3SuSpBK6VXIYppPYF7t80
9ptz/8MZEZDtqIOu2RBjkR9Cu+/oF/NI1uICO9CVKw0GIINRL9fp0MrfNYyPhvh+nL9eJ47+9Z3t
AageuhyyjXUDmUQ+8lh7dQQThU0vnjxE0lEMNWEUSVyfCmRSUfdOp5QH0tTOTSYLmMDnGwlWY/Ec
Q0kQmPeUtazYilBN1vcMLGoeVozugcaHbrIzoDHAMT0//5fum9F4wNy8y7F1SWRWTHvvlflh5st4
mRW3z5HL8teVrVgH9i1+k4JQGqMSOkePckCoj/5TGNF/1kmHvuJ6eqjF7fSdhLW7hS+FmdD/ZDGF
fjDJN8XfmMG5T87zZ806f9EEto1Zb4i3ILB8SMnpliDWvyCEEIH4iyuQXWQl9S8wZiJRxh1+46nt
boRXKv5MXR6+AowFZIJKUcD47kNPX8wgLclFF2+ZTLWOIWLgDMl5FdnuH4QsduVNhxtR4SXhY95l
aZoHDrVfZqIQowd9dEI/m6zNi8X5TCCl1iNp6nBEa+oaPBLN+PGi4vJAuPy/BeOYirLuy43JpqAI
LcyS98NZ6ecL854hBqForeBAjF7fKJkCn28+5APXvp0tPyAwPHlEpqS2U0qNzQcCKmb1tHqXDzFf
5dsHZoM0Jr+QhvmJG2deAh9/deJBFJSQZbcrxf5LsNu+rrl1yXGB2m7Hs2QxT7J3phNFDPpmoHp2
M77sq2PPJb3ljkB76c0Uq6kGVUMTAccL7r/VBogM9/Y6YeNt3/cLg3fH57D5+pLmFk3l7t9/3UHS
yEqHVBAXP3JUMDBNd8aHa4b0RFWvNHdtIED4wPCLQdEQ3AmY+6/3v9qBiCoAf8bxuGi0EutLmXe2
E07vmCXc12zVFAFkWwna2OXB3bGgytD1tMz2phcWWYYJJtNuUJ7gWAVSURaHXm0FYTYkj8/P0qMJ
Xo9WJW1zEAOULK8zRfae/r+M7oSlYM611RScGo3Yusq3yIAGetgQz0YYw76ssjvuo/w9uBSBZ/ea
RYRoFo9yT0x3nbvGF7EaVteppwOnrQ2vJrhRDsYxyBvM49yDX155v6nhTBgEIM+kdCI9u7itgklU
SYJIFuoGp3UzFEia+biBceWbI4bWghh/E43/KxALj1Ynw/k1raQDcn8MRWy1b3gu8HI1QredaQXV
MFMCJFhYWqBBkmcpZM/qAlhD6AWPRWP5brVRfR3/0SzuFDl1LEifii5CZGm4sIxKa9siVKSdJrQd
a2gjpAOl2Z2kDFZhDgx0kkLRhLHCaeHJ7N5i3Pqt1EwC75lEx6BL53gjsYJMBOMZHCO+E3WFrZVl
37A650YLlbUfZPai3RK4pkAV+30XqG2zQQfdhTy6tJAEZnTGJwfPtdargX5kfNWeD2YxNn2/Tk6v
kYTOI9g50wqEU7hh+0tlO0QIdjbrkSFZvO9NHyFys+OnLgZRLM64ZFq46KoQRHFeO1k1Zvi1Wge4
CMznn1B0sdRaHubxotMAUWOSBZ5zqLgan76pn+Qavugrq7dFXn5QMf01AFlyeGs92iGRLQEBF1Te
qSbJddZzF/l0BZsfZHkUEC3pA/wW1/cN6d/bKhjgngNyymzzDuuLCERpVwYiLo0ZXlc7tau3601t
qKdGpAfR7N8BrJZVQnF4kSeX2rtTC11ECj+ODoQIxGIw/6Qwwk49BLiXynvLFIsFu6d9bmRmIJoe
AqScMcq/6ZuDRzRAb1GJSuwX9xlap55+kcg0DLqQagHKi5bapEDXwyQUZMWweTEjQJhVNU7DO1MW
LdbB1h58QPSX0kPiAeH9XIjU5nnN6yC3piIFfc18c8TyFin14A1A2SscO8pN17cqKAsxneT5/zPc
2Bfwv+80kEniHyrN2d0uBO624RjTf+woaP3SqmR5857a4Nf6HrjgXazLF+atbTcIjAyqUIJAvtjm
DpMzRTZdhpuDGrldHKnRXMLqJ6c5wgwf61bPnoE1PcJDjafm4uXM+XJVUeipw4RAcjzu07GgYLKg
ONTRp7Z7FLiT3n+yqA7Xus/+RHAgeo+IuLU8/kAPgmUeerAOiWaXcj9sM8ac6lBCI+0dPcEw0aKN
BBNQgS/sl6q/efSqZ+OgNZlE08wST0m3sMw9SVHHO0fjb2vYFaHeGbN+pPfpppUUWnmVRqzBiwTP
b+V/MuP6wwTTQvJl6zyVR5zAVvScCxtgYRsZczoRMsxBeqhGsCAKAT0W/0RQM7shDBtsO26uaTxy
40W79FXuJOaESCgG68ffX9dQVllvKZo+VPL4eC4EHUuf4NL9W7lQm6OANftZcZVQIITRKf4Vaok6
j0jceRu21GweOVU1cdn3HPXZyHlJ+pvWw4CopWo6i/rJRonSsed+DccjdPmq9aQp9vR1ux1VFMTu
Ll0q8zd5NS6qbRcYvpM8bhAw/IC+BzCWpy7y5yTRd0EklsXAnaFoTOYIcAZGfjLM11gK6t7F9Cy/
mYLvmFFYG6wocibinnczjvJpjzGQf3lsib+yeXlly3GIAJaFF/txHKBWSTMSP5VNyFnRmwvXXGql
ulV2e3Nlaf36J8FX3Wg74usHvw1DXWyp9jma8tjXvb/ro7R9CnIKi+/otIVst57rT5Mi2cSeqc9G
T0Wo9k9hPlaLEtA2IYRKL8RSz+YxTGdwHhwIxfDx8D7c7u6bz4gi82MQvzJc5wpK0USAPXqOT4Ye
5kVloIxPuA08aT/JlyuqVS/QdUtsr5Dh3jOvIQ3TJCfAwmEqL0GKWga3w23KpXclEj5hqw7sRvG5
YTASaqXOAQYpyqEHWCfkh4r4b64Za09QbfIUCfrMqDnBNFLqjmkDGfoLQYvAAfaDlQIBP8DCSM7D
nSw1Qbo12fcuxoIjwwm+BjWR00RC9WXlwg8pzrwb+Wsnocsk7frv3lCJD2LTXajGlTN+V2wEoxuY
TUVzkIOgrRDlv8LHa6FuMfxr70BaVF3vb5oHG5XRPNLQhQ5aDeuN3enH6pJX3C7XrqHwrmsj4J3y
HmDaVBa9e+Tmgk5h0sHo/9ghaBZI5jyIg6bMciB3hKDe/wxr7poBKAys1d2A6NPC3qFW8ECbTqdl
FwNAVuuL1D9wS2OUM4CRV/Xnag76lhJd87iTuGFyOzh8z6fHbyOWpXxKQPkvWR3H29rfE0lJX3C+
FF4rIVtINOc/w9JBcvf1rkf4Y1zXiWvoaeRWfuIht0ZBqvzqKoRvQ8Y1g/LF13goFG1dVaPzwwXj
FlFSdICGyA+FkKVIsNUw+9bCLo5+gxsKp8xg1MQnySAs+dHmBN/eIl2tI2JprKYAUbDzd2UaudT4
NmYiWOw+MZF1TOc6mQXcBkBoYrS08+dqIT7D7qqSxkxWNAHpcEAHifw/syk6Lb8+PEbvX26qJQtD
+31+hhfuZiQApgXYatZKjkyzYJczY5wAWbIsQjeWj3DxRgfCDxKTprJdD4QwEvF+v71swK58M4/Z
J7ao7CXTXTuoEOh15C2oUwftKs5WEXKqkW0xneA9TR2B/kGBTPAi9PQUxPZpSIXRcoKvC9cufitq
ic4DQ7pZFumjkZorJ3MMaTo62wfaJoXRNHi1IhgRaJg1zEPwt7G7OkMW/AXxDfkBWwovdFBaS0/z
UKl+o4i0Glj++jf+990SKAWgkM810Bp/RoQ/y7sMiEi23CvVNhawz3+WXbbHHR0/2Rxmdzg9C2nw
KI2gQlyE0FumZkBaPPnJl054znRuolZElnCR9p+IwDDKeKl3JK218rFG4yVptN/EedyGV79JogEd
B/HiysVNY8JN1EWjdBw0HNrY6zdeZS8X7viitqLwzIQrhIgh1cbg57XHDqoz5ypk7TdYT9mK7Jwz
xAh6E7Jk37cIX7ZE/R2k3z+loYX8+XxLbGr53+jOQJODYjbCo3bW3ul3QQ2Ps9GuFg/SF5qFsWLs
W7hg/yGk02n6KlqnQNZRnUilEjD0KP26CRxIKqSYUu6T9l/ALsNoQLsPkow6mOGBRJxq+WH/007B
/El3ie9KfR5+KSWTNpTgcTgnkQpuT2pzySj1WZyxomOkf9O47qHPJydcVz2IbsdqqspFWhsd34dE
9jlZu0GhmYdeRiDyctlctl4SFuWRZf+0zHbIvwsJ2AA7uLrvUwPA5W/dZ/sYl9z7FSyjaBqXrRyq
51ls+wWZoCl6dJheIPbKc7OCv4x+whj2RvxvkWk6rbK4rg5hjV6dCDjka13/tWOYKdftvRJCQO8M
qQj2hahxVvDCUW3Ezdgb6ie+ceWinGSsl1/tsR5paoP94qNKgim2YO9/FNNq+5fpDRywj7eL/NRw
H1Ltpt8PtcTHmTsntzYC8kblth28VUYGtIwFurxzD3f4BLfslHnosU2faKoUy26p9CZVXTJHvkd/
9tQEGh3OQ1DDwTV2NZchn2vuWbOMw22TKM3lsQE1mzg7LjjyyJhJBSRpmTwjSAcaGM5P92/t1jqf
AsJEEtBIQjY/PtqoFcsISOXjdIaYVikU+jPbftWKtuLLKhfUHliVNizTq0DrJuC0/8vbx0TM1Rox
3heZkFr7epjjYTU8dCWMPjKxwzsS5qJfgMSOeerA2oP+4I7YQNnY2OJJI8Sgkde/XAjmdX5m+FDZ
JJ+9PX8zq57hEqxEmAL6+bZ9yunIlumB2bNy9AJFKDMHyt6owhTdQKJiyFsD8OXDFr/JYICYxrX8
xa6qRaxNxykyuAkVfgKdqqVwXW2k/hdnyjZg2gBYGU+tc4pTx0xuZRYDUSc/c53Lt1H95vTLnzix
EczJmbbw4l9L41wguGeL6F9a9kUg34lldwCrdiE87Zjug/+3xLVdG5wQ8C7heP0gIrDRS38AWKno
HvooD2puRg9kGux6XbXrtHIiwfkXxkeU6kJQGPtVcxfJ/t/MrvF2ex63lw4N0zbZG/YZ2s83inFW
DlxUK8fZ7NS8IS7GS8LDis8GfwYzTJqhVCkxiV/Q3egQF+SBcy4XVuHYxXE/Wu15/vmL+roJCzbO
ikfIq1EK6ona1wgc1+Lp3GTdqDJJ7kjGuKRhfmlzMScXPgyB1tEt1BSiT1uLwwsH/+b8nDQ3+M6D
WJ+QG4cZu2S64IQUa3Do4VQMr/teuoFyifHDpgsjjPEcrOq2VIXDjjSV3wVnAt88BH/iEQkEDhO8
wJe9qLR8sFUAXrj1uo7PfyTVQgo9eXzazFaqTbqD7Nkp20+HX7krPH1s90PbvrvmQdnRJRemp3F/
V4SdQ/ZPegt2a1+sp6eUBdCkLSC5u/31P5kgL7OXiH8fGKUhMbQoiZxJYmb14CdXQmgmAaaR/iSb
7CfepoOAYQ3FNDLi5YquUaPBn5oe0yfP5byYYu17mXCMVZpTP49uQKBtRwcdaD2KwlhjIs5R5qpg
e5yuhOJKb+2ZxT3xyPdMhgVs7/pZIzK0rHBD/X1yPVXd8/604/JPFiu10WreNJIpye/VUrUVtqmm
5TXhDbuldgMTBIZyY+06Le3WA3X9Mpw8ImnHx+XJHt6l2mI/zA3uVlnCtmEKizHXzAQiJfzc/X47
dSbnf0c60sFGjCYcCGdPfRO8wLARBAXiMTpM0NvBer+Kj4Jgrs7Mn2fnjXyDk/EM54SB/Z9HDFFt
90xMfBUIGLxJfdVB1L95N3f5IKW19ovwbH7ftb6p9btKuMHZVdKyZ0QhT1B7PSTFoQY+/tz7viPX
APuluyWlwtvuPEPFwDC3nhj8/k2hpu9hRz6sH/A7uZov9EBmNJWVmmFLaXSV4VKmGOdSE8+P/CJq
yayqhobjE7FGfN7ZXb9u1io8eYgnbHUtmXJWQUKTkzjWbeTY+g/BoAT+Mc8OpyCoAPb922gHDgnt
4ynepsiB+CVDFGSd9SFMrCJEfLxnasDXyyosa6oWUotziHnx0t/2RAsSq7WXC2KVcutFwqcp2cZh
EX1yEKR1QLnmjvTDkHRtbYt9cIMyY0O9yV32R5qltMmkoTulaZOKapEo50qgNJmaLJaT0+XMvecO
cOP1BKc19MxN9aKBmAuUnobpvRCfJv/4YZXWR1d1LxvT8prDo+ca3voXnV+JCJtxTRQcq4Pfw9T5
h/p0u7gCJ7IZDzKV6U42J8Fo1Ul8uoLmcGqBKl7pvAEQOFe+1u8hxMZMtJj6d4ACTTkD1imKXuCw
HWLz3X8QhmonFGCvOYhfx3VDv7MSzg9T5x+E3gVEUI7aQOtIRp7XaKrf/28BdaiDu4nJlwoOCdLt
QeaxobSuOJ4pmIiz9TRN/oIzoowjiymJAGV/UF1Lk0E70LURBjBKkaeNp+PWq2gpw2PTeVXKHpvp
Ms8ciKHsLVFcjmitF567UYbJRFoOD4jTBYKWX6II9sz70bRFKYT+SXl7JG8fR255/ZRn1Bx6UGqx
yUzSYKhhwTV07FLOlHxfI+Gj1q/X2xo8EY/Hurhjk8HPGwfvD0jdzzlnWvwP3z2crplj6nA7N8d/
RDLQyvSgtySYq2nTzh30Q4jv+LE2iSelZzpcNx3F3acm0I9EoKwSpih3ewjs2fqlK8tEC2d95xgh
w5cMby1QpDFZ723IUlLpLnk0UERddSBB+NweioNBe7lCtOWh9lHFPYG+FoaDQ9QfkAvt28frVksY
oNGLKG8zl+KF+Anm9GyBGrNIrNIXngOVBp1HfNV9vLgxvxTLuW0hOxbXhkPuJHCfMNH9G6rcECXG
a3vIlsP+Hw3r0XLt8CKgX9ooP8IoXyjtnnCcaoPGdtDuWrcC3EFmPkel77UdVCfiZHcFiKXBocOy
Rw5oRdcfKwZ6l0RkXpqDT+i3qDHmZBC7VbDBCIpaq9NkBfhq85BRtorhm+P4tAmrDPGBPqsg2JGP
lHU82u7akHiecV/Tl19vCPOX58lzHOE8e8fVh9EyJPXfvyPEiESxQ8dK3Ylsxg6Bnw+0GUCoNdGV
Nll0YThEsUikZalTHHbcJkyLum5e5gm28zmG6XsShCnsUu7wQ+oF54K/rzkfUJBVbnTQs7iTY87/
LroTdw30X59RMHb0Pdz9rTKu8ghqh4TefS9mGcrBbr8Ed3rHQnXvMjxRnJSCPLt2uRhHcrLETT8K
PQuYG0Z6+WHJDsdjtzSxfrNWvLUZRxH6ph6/kdpG2NZPgB1b4WtoqCNU4UeI4zGaGu/S5v08K/n4
yfNYwXw0eQIPdtJMPtXk6JeF3PZD9A7uOFDk/4vi1ST0Ti/FJjSjCkqCunbW0tu8HG0kpmn9YtMc
yTHu1sURTFEykkGKoVJR9GEt3DT4ckYu42odN/7fKdzCIqh57UX435y1SBCcNdj59jPWDa8swRFl
nP6i9/5RL/1P8/MZ71HqZnExOv3wfQlmfROWR1BSQhsY95/OjSnsaZnI41c8PCBfoY/lANI/pzFY
/zzZznivBKPRjQpucJvU5ynzXfDVnx69hTNHatM9m+6IVPJXziVZzZ4sZaRnCszAPTHVCAutQcuk
5bG1Mr7alStKEipR7ATHlTX73KaGpAqDT1EJzIXo6WmA7LkUjDQ/57YyJpgoAASR1XO49yJa6J//
ZJv7AuAoiupHO41GAJkIs0DAjr/fZVzOQN6x5hsJCNyEk+UxspCuD285mGALCnWUEkaPUslIp74b
XTIq32FnnEJSHdBHCZ9PyVSGfUWPdVi1O6zQCsOL0aXTX4tkj5g0P9m/srpobo5J7Pqhh+jXDuAV
9XKCSgAqRIHed3XTttl4KCnmOOlaS5YsYxHm4tIXH44RMzSTMDM3u2Ga0t+cxTsOUvtYPIcKuh6l
Rd8wa7RLE2z+iGUfu1ZdsOp33zx2F/wrLeq+cVq8Qxgry7FFRFQg7S6q7AhWBAn5vPuk6h6+ztV5
JdJZZyxj03iQQKj3KksSO7yVmLjlKVSkyJLJAZpJhTzRrLZtDYmK9pSRZx0mhB6FxqLmDqPPDQwL
z8aXoLZpFdUOOckP9Kn6KmiUYuJZt1/mOXR428L3rhVDRHCh1q15WVOOQrbCKanRxlg4+LnEQhuq
YgNFhXUyF91ZPxZTpS1vlW6kRvpLClJiuYTqjK+Yxp0bJRZn3+Nf91iRtiE54dmROaAsfUvIac5k
Zt96tGe1g+Sa5nCOkfNj1xBPTtkZRf6xURlDWWEI3Sq9zfVmoRvAhcDYCikrRW4S9oMFOj6pyXxb
kfueZZ1q/BksCQ6IcjoX/fSgznbhGcYVzxIAXoG33PsuanHljJAcWUqtfWv2bvoYdhcn0HIFixjq
RjbqFDT50Mrsf+sW7RgnEbKAHwW1gPnn7AzJdDIybgL++Daz4aFIsbfDmMZ9fxqTA9xY7jIzuhfx
ls9gIdrNpe8X/dIUtytpsRtl50tgf7+Nfht9hM+owPbPd7ZI/2J0v7dvE7aqK0OMMVC8hYma1P83
hmEZfgPMoC8hat7dLpEhXQOKFGWOOBXTsFmIb/M/S3UgYohto2cPLlhoH33DOFmavMZMB9IOfliU
MygbUHlcT4SmTB2GQ7bW1hKUR7ElhgS0JxKBuxVuCPgDX3Ikgrx00fpFTGa+ZH0H22T2LNhQLdGa
6JRjZFd1LlVWiti2j/5X7t276spU5SEpeM7Gwv1y2Mh/0Q9PqHoYhMgOGMkJADcrYZAjkCmFEJIZ
81LGAXwo9SFzPBDTtW29J0MgKAysRUbSMrnp5hd5JR/rqVwn56Q0VN6o1aCHn9GIy8b28jUBv5a6
SKopXxBKbI6ad1RHG6vZKACmzcAZKyaX0YGqkD4pitKTGDqXtm7rcje5cVEow7N47mFuQwlBKkXs
Z3cFydpQkBZyXHcRpKUQLGFltP2AYm1vS6vfQbsiGARs0wXLE19pdlP7fBnftrP/nAXZXb5SY27S
rfshIElsxlv5UD/wOt7fIwB8zC/q1z6x0IdGWO76d4ZBNPqjAjFrQ5jd/xIyXqrs/Q/7sGNpPo1/
ckMA6XLiIZBsUnF7Kfxn7jRTapOz9VP/bxA4HLqzl+B1hX9qs8VWmbIlIg/bZ/OAvBTykUPB0QKY
6LCdn+CYZKPULzj+nA4DZ34jgYZIaaYSA1j+4DmjzNN6Kn1Q3WJsQiTPFkq20KjqLArkHAaHb06K
TJTAVCxgHFHqXXQ7MC4CNTel502ntM86MVNNRKMUnp2RUeCmS7tzg87FXIy30RIHb/2Y1ir2CVKl
S+2Cf7c/IAnrRY9fIQSe0NzNRbLGfE46y3MEP/a/nQ2Z9eS1pzxiAtMx2mIRtPyOEWyVpyplgZB/
3pwO9CqBR2w3QnpeZdOE5/G5wjoUNFIjj9XcPgMtIm0lkhBZ1dVSqORXDagxWi89k0Rlzj6EqJqq
eBFr+qTAyjsBKuty9iVAeXjCzhMsJdGsyg6inE7rhL4oeiSdLkLT2SncGdcJpVpk3xGH+pbOJHt2
z7U+6lDu7NETMdJlVM609r3FwusAVe/SNUb7KDZaeCZ3q85hOOj+ED9tsUqPIRUY91PcZGw3EPlj
kLezB0nUJswNYs9i2trM4LqtxWPjzG4fa0U+4I4XRZyDAB/P4z98CgTInAfEDZnyGQfCOMcbmL8l
beFbt74NQpAGsq5ZtITv2n/9q5/1F9qCNRIktVdqWTzvj+aBvl7VetQyx2c+jMt4H7iWp2iZFoCj
MbT3tSE+yKoOYvuDI8YL3UoYMGzLTMAD9amCiKD4qb9bATaCSykykcWu3yntY9JukcEeube2/KC4
I8ezS1CwnQw9oZGf0REC4Ypcy/vg8z6/oNT7YhLgaYjeGjKu52j0pE/n6ai0jBzLwFXrSXdYKOJx
48+36l8oJfSkeiOql4/lxVYWMmVfUqDLudjzlE1x5HquHYNnmNve8uI14RcPN8yFxFwY92ChFIq4
9FXfR5R79qSHxS4x4l+UBpH06isJfmYrJQT2BsiTfSYKpaQs3iI6IjVQv2djWSktKsBUZ2HuUT09
e2+1OUpJ+RjSwrh1OSYoCUXyTDkVuqJS61ipxT/wH1C9+0vI67HKTa5t+xkG+ofTRAeDs7YRM0MV
Hl6WWHTZ3XLTTO6BFCrVoXQg/cl1se5IGptGgQZM+dwINTjfO6drQUB8POi2GjuPhEWYL9nxJIC8
bvtm6ZEMthLroFNyyEWShfUnLN5RINnygb4Yjn5zDPNh/Bv6buoXSTQVT3n4qQXQ80Tjl0pPOu1O
K1XfEsFmEi2ivnXvU0oEDsxwpEcLZcma1U7e1AZcoILm4KZfpudTrlGdsuPqgC9Ux/Truv1AvoUU
BsLHSrJO/P6ZKkCtMKxxhISQoi1okasBuHFPxDUt3xcmS1pAiud/Ip2IIxsVg2O69ovno1+X0czu
BSxCzVk/r87U6R+ntLlbMuZHMgMVDLBj8MGs73x6uCb+Zncve9TRSISGzl0Hmou7mbB8IgDtYv6v
mZpd1ZSYwU1eNF+xL6WgS6PyXRAAHUzcMgUscxcP9tja2Yp6UJuPz/l5EjTQDW95LaY8OMSeKXOa
xurTlB+R1r08mndWzYYazIHMmR+xhuszvBJP6mATAPwxaD/APrNHP0e+wknvN4XOB8HQzAuM255/
JyqVMYvevqxR97Yb2qfFd3Tx6vNim3rnt541Ue7mOJce1qPmY0EsJwojnivUpA0NQATMiEV4uqwp
mv4HeuCfXe/y0ipaXFwEUWvDtaJSLkJUijA3T6Zr2EbIOrBVVegca/Vh2AvqkDjbr7K3ki+hnjrW
Msxa5j/8ZyHlLyc6YD2aKf/Wpc7ciwDSiE5hBKv/DNczRmj+ADrPS9Omzs3/yJHSVeA9NbRULlMP
UcyLst2iFS7/Uledc8GIRPSbaHS8aHfyMqKi6ilFB7pMgY/8JZx38XPk6ZcLqkCbCORkzIEGnBeN
ziHnCFLMVmifHH2hX4IBFOyYR4osZuzPEWIffubmZy6VVAMB9MoH8dFnKRfH7OEwd29EJYsxXfsb
PD5DjGbyQLTbwZf3c1fAHe/U5ADVbx+dWc1vWUBs164DzxOzCZ9PAUj3tLtNLHD3mBLH5ycUwcXg
qJybMJ9uUQIhoSJtdX8wUWpqpNoOkIvEmPYKPw8LJ3g+emucIRQqouynqXdC7iKIpu80FAb/juek
h+uWUxTTg0kgzLs/Y/mvhq4X9I/NGiVq8Gd/R8jYE1XtJtLVm1w4AFPiDGC74e9ws6utzr9xg25J
O26gC6cJZGQ0Vgi82+f25yZX352R41zyLSneej4EQu39h+L5FKBj02KU5gdgFt2At01YK/yRoGRp
5bJF9SnC9DngAVqLbFovk8egwMQPopMaV6TYuFw5ftQbvEmFJKthNmAuBOqAKyOOYABwvsfbzCOS
eCyr4B19keelgxgX4+zVB3qb6D30eQmWCFAnSc48AF05dVLz6oaqRrfEFsr+jLf4W/BZUW1pzili
bMC4uPsfzMXyVtbGlKD9iQFT2HI0CaVCv16McXs1tAMG8oFMJ1YpAnwRF+LqxN0jvrlssLmPi7Sw
QkJyWIZ0/kzG2sJSnCpwD6kdoknA63oCwpYi4AKoZczXeRpRGDB6m23sRW0WJ1cOIuUsdSri6quH
9HPzGpYRo6b5MEEoTsrN6KtB3wRs71Xjx9CNR80Qd4gCU4XN2muLnW6V0puHYUb1oJSBDTBXm5Y3
VoW5EmTo6eS8dacN72HML58gHh3L2fqigiV79aCvJjObTb5mnWluiWHHombPEIM6ga6X8GUl8zFD
I9uwXJLqtlHMP39tIN13I/EBgE0Nn5veTNKGVlRAbnAM4ySYtIJqJZzfPxxZLtNcOGzf+eBqABq7
fQ4+jyU/DwiPqHkUX6brSbWiVXEtmr6XFBGO5bl27spegnR5HALnYsUtFwxzm7k5DMJXqn4asM80
CGcRyJWGttExngxZZ/fKwUfdkzvOVSmxLoO4YtjHkdWUrTH3gdEXYGqVKK1De+D3DF480D9HBEBo
QaWHyG5Rir3+fYtTkSUCbYLu5tnYgA2OgF7WdtaBAiYSAnWSKAAgS3VEwgP6fwC3q+WosxSMSJLM
SmJNYHfEAiQW/AOxDErVBdzZNAnNLVmF3jf1dqQDRf9nzBccxltDUyopGaJ4mFLYUJgO8U/s3a3v
W2faKbb1yXGrLx/g5Qp8e1Obra1gaMgLhntOvlU9Lze6PdGidShdi7a7wzNRd0FPCnLpxKiN7cTy
PeONUqjkdggvTJgfcreisRdBzh52WI8BF8uvnHUvMpqPNxhE9trf2lLSVSSDpq7OqeikiYTKHGd2
Qr0NtyO9wA+PBmukqk49M9sqJZG60WRfFzw5u3yzieey1ulYjYlrTL3hKYnRQlFUo0xwx+jG8+ak
f2izLDoFJ++fnvflvdhMTd1jT5cC8Q1ikmTMEoHYlo4OF9iANWBIX822if7NQvzxz32ooIP/+eBz
dcbZX7qGicybqSoEFywpFGOAfeHbBgZwMvK9G1QYyosziq/Vc9kgAanl4v8HtoFJP5avaw9x1kaw
u3Vq2m/JjgaEwBFvUzRCmuCTn9y0zxRRz5els553psc0UQmcbo4s2uWD0RG4M/X8srpQVWpNORmB
Tu6HBvy0KHK/Gdn6NI+jGuPxvI+z1zeojuZFqPchVL5yQp6VTIXGUWXtHwnV6FiPLJElszvZwV++
uOxQfZ800rOmASbDOjdXN1Gptj91PYg0CJ39YaIsxaG3s0Qexyt/ehJiqWOEQDJcFaZu29vApXFk
dR69cws71l28Z1hv9DFmISyKjxKq/D90NPF5Ba3pSQSYtyQHOqKBJKi3rZW5b1NVzzOp66hEMW1J
T0UP08xKA6t7ZXa0q4eOyUxiXY5tYtwkGwA+H8sfE36eeDeCbUtAl4uRGurF8UiBWhRR0cC/r8kW
KVHAjIZBp+Xjvl+cgM/yZJB4ulEaKZ5gaQsJ6vA8T92HPx08qgY10yOTAiW4lXizZTpHc6ywXnvu
3vVmFvIdeJ8pJHwtCZwyL2093ebSHTugsZVpRUwiRgoWcKxABkOyAjA5GMRCLr9kYGmABRQHYMT5
zJME046ztP+Pij1eJrlsueykq0r6gnxkBr59cIUYKpPw9CCalaR6mbpPkyMyWKB05yh7iiHpanup
3czVkiYy7kCa9QxtVPwaEcwaeAK9d6/Q/4LUnabybdefEHA5Z2XAEhkPhvdtF3Wim6vKhddH85yY
CUzP6TRXBo4a0RjdCe5PwVBf6EDiST9rDLmJRPWjKEDunA9wEpLXGYotRF9tv+d+MhMunFO1Ajb0
mEnMQ+baMEQV2Q6KJXXFMYAptovpLlqmUZxdpTvZEv8xFs3rh/kvv62aRjw1tOKHbMgEYPPacwSO
f/XtIm55luo5Z0wtcmm32eiyGNnp9S+kCthC5UUB698s8iUEs8JzSpejZnFgCHA7K5OtoMhwmxwv
5mnNqiSrC89lcIwXziNHmBppnspsQcMQledIoneV5VZKcx5qeld9P92IQe6PF786WA2LDjVXdcl+
T+XAkvm18oqvsphi4QdzI0P/ppQcw+NuY0l1L6z4b+z62Qr432aEw4b6BYyctU+k5fwaHrGuzDMv
izI29SuP8tkjx2VxymsxZF2ky/E4lMog9EwTDTv1KgLSMwiPAOHHJyjuqNWaE3CidlCZh7lFuhW1
ZxK4uiugIYrsDyiUsiB3LOOY6ZM7L5nLQ6xiYZzDVGlIeJzSzswy04Cu/dVairWaipuf3JnvYMoU
jwa+tfiBQ/P08ldPHtTUpvIlXnHMMcfSa4braya5xM1UieTlhpIlU6+lTpf9WRBFEwR7rnZ2tnHS
jutgtbIZ3IydWyI5cbyKXdPnv5SBBrmT6V3WgmTCT/ziRe6mKauj0oa5uujn5OlzZUfFkvvn0ZB1
CdV1BrtHlYxWW7P2YGGZCzThphO4k03eoXOmwz65tcCQoLbhbBYnSQcQvJm/TMC7Gp/8QuF26+Wg
0NXEtAnZdNtL/iUK5VcQe+A6Gx5ZyFBRJOCUNOGQ1TI2efBWm5cik/P76vuADjkSP7pDZXj3Mm+i
+BrXYEZrx0gXWGm2vSADGlCsB8/9tspXcsr/SrfhoqXvldhz4y0yjTZTNW/9p7nxOAgm/SFO+C72
oHUlEHQyUux1/v8PMhl/Ps8a5oPhq3XkDsWROqXV7ShcMLf0CkUBR5CQY8MaV04N35hgiqERyDWe
q5m2JRLCkWpy9vqMd9hYRISenI8NsVYXyqnCwONe2vvlHpoX9ZmIDW+qXFSYbuBnmtQ+WE69Nejd
Fs2vfS9ZQi7/3kuAemrJgGsVraWxu3A7tWuZEge4GapAfhhn7s2BsHB9+GE1l1J8zKLEs4O9s7Rd
HYFTUeMWKQnHjzxkKVWYhCy86XhSGozT2E7o9YhwNb9bUpDyWVZezAD9JC1llDuZ6dPuwltQhc6R
BiOX7UdnAzZTguMqGreM1ioexWQwAv5OVfjzcZhBWaKAckfB4GzAnprhAOiD2OizoMUzhLwaGkkC
pVyFGTqSSb9UWV0BwE1FuThJHGDoQZm8LAimZt1UeeDZolYUFwS0vJR8aSaAzjjtxavIbcqtKDBZ
oa92WvgYlj2XQgpnbHGNGL0+W5jh7PRbsAqZL6pPBNn0a0HDqI6H20ndjRCXupFudVmXNY7GL4G9
L9zoOeopmqUHfefgr0ATkAizdye/wa/LN6WLF592g3TYdI2lqnLQQ+ofB1P3+f41EOv6QLRiQ6Qx
B0VaTNKa1wZkUDeVhfrlygYxOkcLjsG1EkA+mtOEui5uGI2Sgr2I0sAAdoRKbHW9c1OdkVwhrIbO
QSuCp1Nrbmqz40fQoTKAg/vd06zrdPAoxAulyu2I+kuvWWgCL4sykBqtZHvakWqCXzVWfFMVoSX1
t4Ufg+QiOoMkgX3yn0+Cd/nU0ifwLUR5A8LHBHT5wbUslPVM1ZTow3+cKVtnE8T0ZL9a5+EyfLHb
YLJw5oIU31w8yr+l+xajYMe9RX7GCtyWjB0wFW3JyQHQetgNQ+HreFquLS9SGe8TnT+WnitmY8U3
LUFQd+H8+0bdYn/hayB/a9y3quO2QWO0//CAytq2ZfHdrFPMRTisQ0YSu7sFZwQNtWy4xukYWsbU
6oJ3vyggwpn8ni7M50Tn7HXzLgr/Ag2pE6WbH2o5R6g9dUCT0CtircBWJ9o3IzQOg/HPekRs61kA
mCsyEsm5y8r8waCg8e3rDaqV+B+SQj0O0sRnt15uySWaM5repKJbllQr8liN5YACgyv8ynbm4Na9
N5pb71sUl1pCLMiZWWKa5ur5nE/AViUNkt5lzikPPFN+AG6i+pEVOULbKQIcUsV4Ngg7Gig8k2w7
hWLiuKc+rWMLQZ2Eby02BCytMX3DPs5LyoOGruTXtuCSQ9HuW04fmPeGoAdIQXlkMKBDPjrJDtUY
F6ad+NHeQwnC5JQvP+HVNL5kj7M8sree3z925+W4p6g206mLrjfonWnyux5sfmL29j2Rr3YpRO6m
8ODqFmQTBzQohTptpcdvfcM2iYHCbs004RGH2nscWAPQ/FOvpu7uX3rdEKWU9uHk6H6TezW8+3Sx
uT5BrS6ffSV3CNU/e3r0hiOg5qVL3MUaMzTLeBMxxcKEBUT+eKDIoHRVLte+n0ZGgMJE7voGsdm+
4IWaE8bTExwwOuD9qP89RotNbd6IL+v6jXKedyIwOmD+D4+sljWVOLuwu25j3LLmy4VVhWpJrI3N
ylLFJLMsSRdrEUO9jSxHgC+8o69pRKERX1MI1c037PHLK/CQltSwV+u01pddXPkD/oW0kH9JWuTT
74Fk21D7wtgThpqBBOHJJ40VhrQ3vsRbHC4FVfydM7DWR43vJ2KrpTMOBZUg+AMqbxWZ/e6TJ5AE
uCAss8kpsjPE9CDkIsPB5sYzS853OltocRn4VLV0/ipVUo0JsV4ZLnCi8qDvqxwbPllsWlZHG8S4
xhwE3qu7Pt4X6NDs1nBus9CNexXKQeorH2Y2AytHH1TgNaKH2AWOe7sdQzsHZTEoFJgjPhnb6YdV
XK3/d50MXEObnfJRNb3kFxhBXJGvs9AK+7u6m+vcHMJj5j4ykZ55QsGAm6NmjSzWJREMdarb8bij
wwTFdpfOpieI2JA14nqdLvNb5bXeiicFuykTJc96o/x+BUp6CgXj1hCPI0LScJhtorRDaXqXQey9
xOEZjN5GIK8j6KXKRkht3MUTl5PzU/yJt+ZyCDE3X+LtX5Ia+tRUTbXjbFw9TsCgZDWsPEqENJ9w
UsYrXp+4I2z6OR0G3mgSVSRCGzvUKV2ZH8knRSlPRRQMU1IbCyLzD3KcMZBjw9sH0XN2frnocnZM
YtsMQPSLK5dhQcuJk0+N41r6KHMUa+biIChXdLgspFs6AXaCKtAnoeaYW1EOonplpr33dimLD4a3
i2fWvFEoggb/YC7NtBJaNCOnFg1NP0bNUl+9+wHsg3wtyagP5R/ioPuJ+0XpRob4RJIUKUXpYAU7
18MZFR7/BWFYT9rCy6BZ7lFgCPeiJ30DARQS/gvSMDNb5wecEvxzwBthvzNuG3MXudBEH3k8FrKk
QLjPwTBI5+pfWsljmQeBkvE8dYJ8MX5RaCbplI9wGo9E6fLZgT76JYfP9ULldPcYzvS1g9OBgz51
CNVwfhfGjSfTynhzyDNmCTO5R8LzSa7jR/duEa3aySVG9q+e49rbPrrEHRFfNgKbTuXX7fH4Xw1W
t0N3YyGDMv8jEg8VpbYF3ylVixDGTksTqM2qg8q6asoX9BNQUaFvcl7sXvOoeptc44oVBAOgWRCO
mtldAX6ohvG/Cn9vfnpVubS4lAAt7tqehJg7eoQjCQ6r7lVX/4a6Lq4s+0NpIPIOi8hCDRQTdNr6
TSEmryBqSNgUlks4xUy26fqcZOt2ep4C8gbcPIMet+OOBVincHYYRD/2jWbsrWW5Lamwj37SMr1x
VQalhi+wohk6clrTUjwMrgE96O914Y2ZCyEW3YNb0W/+tuc/WuKi8Ni0ULJma89lrXjO6FTc2v8x
ZLqefTz03FBhSwZIYV9MZp5KouWHgThm9A2NPIHvBCpvUKbNbxqsNvsftLPImNYOQPxy4nfBkW3z
80uEnKWdp48GIJh1HhibQ8GJ5pZH6+b2c2sXKuPD8U/PDjitaiNhfCIngxaDyUvrpjG4/6158aGF
6eRUDkTqCyMhXPPt0ZecYLvS6nL666xLftQK9ryd4DuxQwEn1KMtiFFwdg1eSzMWyZeYEIuiUwNT
05/J7mHNRD+W1Y63A/J8iLy3BEZeWLEF/qm89GvBXRZS2hGcVLXrZ1HGktzRvjJI1Zzbl9PZi7CM
omVtkv4fjS3GMLNtPn4OE9fNkjWOp694OZyb+gxEp8bZf7jyVCjMyJuEAMXjbU2kHDfEvwY1jZpj
cAF6o7O9ijQAgUtB0M39DBWQSDOvzBe+uyk8pcsn6eIK42IhGfhUrrPw3xG9Y/6Yhm49whTNsHqY
914itPwVaRHlVYrYxPowVQza71L77leoZWMh5rfu+5tMEYTuyUUKYW5tuPs9nDTUJKQukZvk8VB/
gBf7VuKQJXcZYDVSJVATWC3A0E67s1t/5pEQRfZ+fi9o3vJjwdaTgCNtAgiO8D4n9YzE2U6tH7nG
/IkxzbilIN1wPqM2OR3BtNnEeHhYa95h7/0nr3/vxTVJ/L0SoGYE/foNKzc4pLFtlSioF4AiMUyZ
/ifwcmTAcymd9Om92FO4J8cvzkwaPGizgHloNkgqE1w5S2NTIkT8k2/n/T0zNVZfg9acHIa8/Ykk
7nx+WqfCkDB3k76Hkikd0csLraPxTf6ZU0RKlwD5L5+mtUwehcfzgphPsLgku74nh/DC8GOU/cTJ
7lj9KkaINk4NUq2pbRc9Cunp3dlT7uDGYwazIejCeXdjlBXxXOPwJzWY3HFApBu9mrVpdyaDZlma
LGzNUJG01X+nYwas+q28fWGqg/xOhv+aDKy1EX9sgRd5DlJxvvaXRMhPFWs5EWfGzzpxfymAqsrK
FuQD9GMNAu5D4Ao3PAY1T9VxUHVNf6YaSL5SKLzGM4wEEwzYvmgqPN3YMB8S2CJDS5lhDX5XC3S9
GViQtzodSc01hL31soZq6g6lRttHjyZUrBX/Vvv5X25+QjNhAgTzX+rMbFBnTAjDdZMb7yJIdkOT
W07XRCfepfhS9Nh7Ki4uSuxxY7LpK914jZqNPxK0C5KDh44feraIrD5z52o+aBHUPRF5mTEkvfsc
l8hjQiJ3L17D2OVMf05H+ovY0IAncE8dkaa4mkjTCe91nh0V/zMn/L86gjq1HsBTiPXjm5U2kX1u
wTKTB9fUjKRL9epTgacbi95akTWaxL7DiHgGQIBWvHjXBr40t5A6D3bpzuKPD/TMuhQs7V8HxZDL
EDJ//8YTLCn7RexzL2g3MuzUoHn50f3RnwkATkVGWMQ8LjUt2dG/F+qCEeTfI8rrhGdw8A2jArow
UVGCm/10ECfUEty8uuP7vFROg73/IOlX7kX7lPO+mmAoD57bj7q6rklG7gS8mJX4ZgrYzEDFA1qf
XEFOZeKm09v7375GOqniEctSmry1mpHztuUzRKNdSE/gSstB2Tm+gR29YRfZhGNVkwYx8CDZsS3V
Sg2pbEnxa+ItrSnkDBpcC9sRMZg8Abkr+CTy2Ef1Vx/SQGVfKOdyvsNYpkZLESxnP8gFEEFOk/rc
WCZU5h29YTILb3fCRWRflaJGLc1JE9leWH3S0eu+rEyggtJC8VA8wLcuVP5OWAYmsZeu9uY1kKSl
yxN+vHIJW2iUVWlwKW4q4LuqMuptRGjbN0k16peuKb77AVwjaIRiw3GK3ktaqjSIkEqE5dny8ubF
yMhdUdxbuPVxBXlZZdQ3NJyC/M3UXBv92u1JtywzuvbTm1pBFbigy3UwUfBsw5snAuz9pExHQsXW
faa3uLaOnoAgvVvLgrzzf3X7hFjdqX7ELO68aE4OiGc3TxuwkwoPMgq7HbiIprti3SOJ5IAH1bd7
Zc+MUSbkjYtLmiDVWsjD/Pj+zBEB9DjAVKlDQtPDH4Tv9ddNqUIvkrGq1KhvWtR5QnVYo5QS8pTC
AM3/pf7qKvPNkd7oaHf6V6MfTcp2baGpFqN27JY8kQZlxGi2q6sS7KTuFf6fjqKVtU1il4fpD14H
KK3wFo0rrKPSRHAvc4HkY4qJ9p2Qy0t9lJVrZNw669IoDoq72xwBHY+V/FATbqHW8r1QOEKisf+y
HzNwaqozZNbE5TtVQK9Ioe3zMVZcfsgOKd6dhpaEnjhHM65eq9qu4i5uPo3Tn0KZsV7kgLkE3tdw
Pq6jm0aaNqTsPEKrA+GRL7zPJCigdFS1CdZuD6o1o4EOStWZfe9xx8Ee8wOdKNbtNi5O19Pf3UgK
pbXpy9q/7/pNKvv4gqN2SuGgl+Kus8UG1sziweElBxVpZIHd2gMvjL9wvuCVVHBx5Kf4dvlrARrg
wBKGTtahGVe8GjkutOEDjrq8C4Qfnv5blLjfA/hOMRjaFOmsREfZAkZ+I+XklFUMXS80UKrtbxu/
5Pom9hdT6ke9J8o8bcF8xM74z8Yp+3rcKFKfh7xxRV54q2v0ID4jQxflvuP5i9OA+XUrAFFE7bEB
EXN5KymyZ8ymH7OYquqbAecrKjLZQ4BiFrIrjdglaQuTEwzr9PSlkSOUzZwJE9i38pBr+g+Mp2qK
WsKib/4LaF7pxHUZqHO18HR2nPvQTV7GuJ1W4PmL7qqRbzTmJWeAHoP8lEPdsqq4Zf/0zxWZmfcB
ESsNlhaot33Fk2jGa/uij7eZO9ifandT4g1lTgJhRFTAGf83Bb/OG3OVot7sSlm2aunoBzNn2Hx6
m4r3j94frodFWn5FJb28uDkuVMNCY4BUfaHwXoT6wDpJUalzMYvImmU5juym3ZrV6upQ+MlBwndy
4RdRpW57eRp3eonO73qH+hx/CQtlT2H4jdZuF4Tz/3YtRKKaDLpinK/b9wVb7CE/R0s+t3iTBYU9
feK2t68IcxSPwuTLgVBvA5zFJHokwkxCi5JFP0HYo2P8iNE3SyeeLyhk3SIbZ5TFvE/UViJL2NrX
lpoXAk6vQlZHXc/lan1CGlgbhFSCYaz+VKWcw2tyRsuSsu8zQOW80cjAbeQEmmtYPXq2yf69UXIL
XZALDOyf/OYAX3NjqYW9DC77WHA3g4ioTn/DRS8zrw36V3YE8yWFN8Wy5tEZ+WvkOjMQxElP9Amp
IRmKcNtFag4aQqt01MeacmmvFQcEj/xeLa8qr+Ip7ZdTaxLG4m3RCPDLab09fY/CVSm9ViA0lp3k
NqpqlZk4vO8amWd4rDhQdSUEJFLSFqEmguh2EugO7PjEz7koQi+R27M5glIiNvV+Ie/pp0uS1Pra
dcMX7SK2zWhL061tAq1QymVheAv7YHA9T1DixQ90xVzmMhWCwP9gcArFWVp42LXtljCYY08yN441
OIFrO6ycwy+gmRniaantmXwsC4/T4axxuAD2F50wVbbW1GGTc+h2sPjBe6QyxxrxmHG+yBB9hxw4
bxQBU7WfK8Tq+RCOZMsfgBONqwhtUd/a6UKofpPed87qH5Mn8ZJYQXlPspGOgT46ltkUGH8pEzbo
r4FmrqnAVchHIOsYs8MQWtWqNOUhVZOq6sIn2gM7zjQt5H2wCG3T229/DvdEV8Ch+IGVSm7veqfY
eNwpltHlK16cTFnTNKrTHaBh5hxbLhyBy/oY5XW/eDsy+PGv+DODRT8SKn5HBM9aSgwAWgyNu7BB
MeX2GqAqTIpSd7sQNz/jdTojcsZT3Cyf/fmiwrHqe8t2aBlrDuJEbPrZT07qangFodMurYQoD9l+
77zstjpZFZoQuvR/nefUVCCU6/gVSUHFwkj+MbmxJvTmPv3k/SSneZddbAynsVqGWW3eYU25UZux
t561KXDUYLEqXrQ51P79Z+V9ozBwQ0Ho9r6tLzHZLq9DvaZ7mzr5RLR8HK9xxZe8JVLso7qecUe2
WY4cx5UYmfn48VSMZm6UWwYl4bWXkSI1RdYcbmtJ/G8PLaS7g1XsbPh0oLLCqTfKQBqvzhrAbbAM
tdbp4izKUnAiT/GDhFTAHIGbpxAE4JpSyryiXYQGn+IOTfl+PhYCkTlzio584ZpuU0gXxceu/iEA
ZSV3qhA9Xcz9riXVcbPyUnb6+kHu6aVdzgK7QGqcOhxQgs1fj43cqu8vY4Rfc02jssrC8/hy8fuT
PWB1qLc1TZVWM6Se2d+/yqsmkUxcI7VHp5UVM3MZ5RiHLu9QyqV2ukbGc0OmDAVVovtlaXqd5RK2
HqUWTsddnR4Oq6QSslX/HDTU0YNPluIqRjK9JtyemoNAZ69KsZoaGPD4ChfIi98otUkUdNmLzdra
PkRgiMUI81H6yIHlv6iO436vE3UDqKVlJjky4C9XJRBMSCp4A7XHO9DgqNZ1C3AF8MDCb5mlJclv
3Uh3LZh+TCFKMy98chAyjWMpACO6Gv5Fn/O4sAu+qpkRA3fKeThB4jGQM3U9+gkihyxN50b1NFIK
qJjgEVlFXWtoN/7c5kaA7kVsNjImbMPISuckKIGTGzRyT5PhUZj3z6OSLtyqR7NPqFmo9ry81/YV
pV04dZRlowNa+e4x0/IErBzC/NvoHGK7beLJ2vy9G9okVaU9DBcpmMr1AwZty4GM6eFSVBIk6keD
MRfGnyTdwt22SdWiLod9JNKhLok1idzMJcihvB7BudfoeknNY7It5ggDsIDadXN6vlF9raKF9fY9
HIQ0UyiGXHfnpYT4SBoshce5OhYV/KNX8oAMk5IeBHBn3qXMiY5gOrD5g1uv8bOSMWcSFw485lx+
iMKaG1qyNHO2zYiU8+B+sqOhQCph/lfFlcrFOJ1dW4rhkWj3JJoqwk+P/QJq5didv8gpTU0KYFFX
MY16rK/+B6FzgZNjxg1gnDz7MKQ4sn4dW/Hpa7e/1KupU6MUjTdFU6e1w6zBDwip+KKvtId4Ned1
aNbAM6It16uVGP+cIuw0nqkcqQtbNdatcByzIjxVGvEKKpe5J5N9MyXRTwraOJi9tt1F0M5uNh6l
l5eZZ6/FQzq5ylfKmaU7nWI4gH6d0SmLcyw1+LYBiiZKEYZ1lkcrV1B9KJKnQTEXZ30d5igd+2x0
c3jTQgcARpFAfAsXtsOhUI0IKPR7fZGjAOuVpas8LUF5tpmhJbfFXH4U7StyU5qJ/yxm2GyRjZ9P
dQEFWUuixpbyJI3qMX6pF1ldJBBRz9xJcsp6deUamSJpJ7m3fl+sI7j7eE0s/vTuNwnCVLEy427h
8U5lJPPRBpNxY9wPmq433DyxsLDPLTPoYc/HKdKHz2lJepbLvXDON4QjsCt024+oVaE2VgFFt0jj
VinqJmc7e7xZ3rZfll0V+WMaGqpDdInmfNzQwqOBMI5ZXvKlmhhh+8SLqfvJO9SbR24f6IwRICyc
J0X9EQE0yxqTI+aDn0kWcizN/4GBKXKTiYAyLr3Cbz8f8KgaOt/c/4+VQe/s29qpnH2fA88l5vbe
zTRybcZyMEZJ6FmqpWAqtremfre6JkHlIs/0I0hrcdFIR8787eR/9/uY8zkVKqIDvDSFhYAw0Ry+
vK2YhU5xwmCtwHHo5DUv0J7L2kk4IF74ve9n+Vg5uFQZskFVxl6jD7jPxSbaTmDhVttwdlcrdSsP
DVmfqFZ11fDC4sXENkqcmxGJlyYmyu/t3zntGb/mm7JbUiKDVDpVQWbcIlkIHJB20FI+K/k+aTq1
WEAADZNcbZ1J1nbiA3VHIA4Z+XRrDwDi3qetWXNtezthtfcedi+iZ+6b54qGbCJ6BzrMyWF1Zt9E
mOLu6kxf/mjbTkmuz4TiPhu0TTwY84veN9hRNrlMGjYym3HyQEK0lXIbUVy6Wy++sdUECzG9ckd4
UhTfDM4bO5pyn/ev4qXQ3+GxKxZvQPOH047JFfXHru08yQ8TIw34BecKJK7skstlhfv75QfrJC/l
xxXuqi6Z3xykwxLLkEy92cZ2XoZ6B6KYasxBE4VjNRzKUm56GyoYElMQ46iCx+UvP6WqNXUMSFWH
sEwgOmvjRYJ9DZqsYs8FUGAemHgYDZZMG6cwwr5uZ8+pmqIlP5AKPOXJw68IeZH5oVtqMUBWXDDE
cbGNmLfYWEr7/IOTgELaPRa5KiZjzFJY/JWYmQjdF4UKwvoGeVpcC0HFdPt/4WQ2UI1LoqABxQzw
2j5bHrIG9INWELZBdkk4n4zDy4UccmJmRXmKPK38us7/zo7PDhLlEoBQEeSMYFcA9HxPkAwW94hq
rAmqwW23jT27LWr9bXyvHVM5Aanws/rjHNHoEEYdsyfYaxHXVcSJo951KzfsWIGWDR4JxWHOHoJh
KjcF+pyQnHp6J1TLwkML5Kl/9CqOYqjNGXN9tL0HAtAp2ATxvDplQ29ApGQTgbi/1TtiUXUIy0pu
NdFubGkQA6eYJhPnxWnlfkftGqPR4WJR4B/p6TiLqEWYEBszmj7QcQv23pzpyBr+9CVkT8wncvFH
Mxfh7RKLXKwJ9fozvl8mA6W78W2keSCBtZ5DdZ8WQSxU5F1R9I+UeFJWbOSBIU8baOYnEnI/pZgw
yF5yFUatC6QF2XTrZoNzaWzeazAXKa97uAiB6itCLplo3/ALfLhuY42oQc8NFtTLbGEFVJV4DUw5
h/XvFpD6Y13xOjPl1X1Ff0XyhEp0QMQ2JrZOXClfYaF8RpB+eZOMe2/nCOFgYdLBwDFZNhE8FVyJ
hRiMIPKnMA8+rZY5NbQ7YsLHjQjSia8t0pMo//8aGlQ3rJzIqTCRjKBIYZ1B3B9Kjikua97GWR5C
szJIIBwkLk32k+YgXSDxeeT7uVZO9gqDcmCpsPytXoTjlZun30lOeOPQE7NDNvDbwcqr5soErbdK
bV/VI9xEFhTtiZYzqq+1cicYA7kH02tFMYDVtP3cclR8i7p2+SzPI4E8/QSKCqMce/figB/JqqlK
u8tz6pBdwzO2yuJ8+PwoD16efAZsInbsE73erpgOKPFncA94rpzm93RZ+j5XOsumwUYFmlI8LXql
bEJjm/GPVz9QuP0FfOsvSvUVmTXFZKdJLze2fqy4Jr1kkM6u+hIn/aMGONpJUs40BrgFSlUvP1cS
U1b0QqvDdLOdwxS29b2acUb68WuodGxgDjcbzRK8U8Ok2WfoDe+mEvWc+vAYiQmVjo0WPIBi/TCO
CFhd0InbaQ6PlpNoqm39q1mRyhXGONliF5TIkITkLeHYYFolY3lGEIAs+jkoGwQsALznJbD/bBj/
7aITfrdnxIg8WwrmPEZzWBmkR+xdn8Z71/mTjdmrn9mxZ0u8xAhpYYVsW0Ysi6H/XXNBiI425Ht1
8UNOFVkWzsIwEwRK3j1Nrwuk4hU0zL/nuJyBE5Jc1JshU4JzsXllBIFzCjp9Tqs94NvUEL7qnbA4
T2wu1ivbYevlkUPuPskr+llztLmt79Nfxu2jBlD+eIbGF2XYr6vCDh+BbpbLRtZpaLbFHww78v6O
CHLZLFY1OOiBIQawMqAzBsmPFOG5mdviwCiU0Pk7mndJgGCnp8DPE4G7CMCtcFZq+axc6Lgc58mv
xDF46gB0YkBKn7BOHX83qktCxN/30gqml5p1ggFH/rDtmmMscXLk0y9FKpghdqj+PqecVcH1pWvW
ZZz6B8vRHR09Ca0Wjqz5SiYRptGvUCArJXVcPWunLSzxa3z2zEuPFCUfZuVM1qE0WehyHKrzIDbt
E3lry0+mPt0/mV0JmuCpeQJB3GYsgx9Cc9h3rUfJe6Q0BM1Z5qd8F9hUwPYnZsn1xZ7YAd2heO00
KioOA9MaREl56JiR3a9ylXqsyQzUiD3He1Gj6MNXgq+rUHDF1DxGxUhar4ejV68s8DAZgNHmg30a
RlLebUkuDRvgFUCUfwc9dh54MkxWi7lDibEqznog/aQR80v2MEOd1/KU0ZHxBSN7HjWeuGY2ZE4p
TuaCM414bCb5dpbpJJDUQM0sH4inomg0qc3kZUNKqSXEeKkvbH0pTXy9LjtnZwc5D47gBIIkMOJm
8JA4QqcZNmqEvoICTvxnIKK2/vAvPlAutkWmJjtVaxI3SWpmUmBBSaEOei7cVD4ZeLKE0XhJNJ7N
xTfRFjgEKb2s70GcTZMFYYdozKUBK7zr+yvYtciKD1HgeIn2YN/BDv5qio3n6TpCjkPOpIMSsP5n
LjZ2yQDwc9W/39ZHgPVGxKpbHp1Stkx7lCMuELymdbXno2CU/I9rruwSvI9hO3rvaeCoIllkYjhg
911djnSHpFEwApOv2iLvtnUxiMttGQ8a2nWUsGSklgGrZg8j6rEqWy1vpmWJ2bzotGvjTPZ5TqUN
fy36YcM78T1BiRYglPy44zUDXXkZfqhsvVLUM6iRpU4q3dkp4vxZHTdM3JuYFol8IKXVYshgjALJ
Kb7cxo52kDLWnHvBH41vMI2Z0eAICx7584Q6dsN/wZ+iwE+RnmR1dHKL3QJZX2sslT0J5hMgrBW3
x7iXs3F6tFBMd2fqf6klYjaS2c24Wqnmht31ZDJMfNmMlcBUridQPLh9tMo0JoWUgakcs83ZXQWU
HsgxZxFsJKl4DmBGF2bXhs93+/4yhOkvF25JNFrjUrxCHCEEBD2MEfI3F+VLwoit/xSyP0EpI2jP
w3hr6s6+6hv23vxCX5tsiUpn8d/ZSDyKxnw8VAoY8ypLl2Ebdc+K8FSnEjkAaCN/16YyMZxhHxWW
3syXYe8cmToAwJzl9P2rySPr/S6iZN26KpNkjHnDX+yY0WCcMx7AxBcP6Lcs0S1zFjZDRxa0a+Jo
QuPa0ifofyFWMQAWMHvCUuNJ6SHObKwRGvmlVQy5lZsTxo5QcqMUZxN1JvKlGZThDhQhOQI0BJP4
4i/TPRfezG43dd6y054OoOwJhd2ARwOf4jwv1Ipkq6SfPa0eKnCca1i9YJTagIXTSNE4WzNlP0Qe
dZ2bqoyOY5J50qJKsct5uttBH6SvhGgd7u55ZwioS3ArpuIFToBr/0hA6Arosta260Ow96uukA0d
pz2JBAU0W6LRmzZ6JgV3zjW7SSzoMCrnziIAgbKM4ZDWjFk0UGoDxA5+XRuAr+l3MKASM1j9umjX
OaWb0EQoiLb0CckmW4IzYz5tJfJFqQf9J+u7tgrO4mchw5tf3VbJQ7khWY4Z++VUslxbeE57s3Vc
1GAS/RgySuLvKZKdi6yxdDz/HrGqR+Sc8FKiQk5qltXIw6Ijl+Z3S9lbpvcTs+S1Z16aJAxcxAiW
HI3d0AsIUVBHpUogICLwOy96VqPLn7ADs4SIFWsNz6raOxVKd2vHAH6VK5kaqrwACHK2E/lnSRoN
bBFJv/knigrPFKx51hgDTEp3OOfWTV2DcVNUekzf3vc+KiLJE3hAhZ1hS1x/dn/xkoHe0t+eTuvL
wQ2QnhKVNJmZrIP2n9K+5sz/0R50HlCxYizac/YDzl8Aaz9UvTX5xyQ3muQ8ZOXKA9tFW4eTqucg
EGOTR3WvsM4aSVJrwztHwdwPwV2isr/4FyaIXedfIGoROPmyi3iEH1uCpCY+BAK4O2aTecvD+hol
uZCrNVjCDhVmx50q4Tx5Egd0WhzvmfjbJbDrU3C6OeIQ+TdfSiFxMLxzrb/lbXRMbhMXrQIm+I87
Szvfs2KgVF/AzSesnEtZ5Dn22/WNKaq88RfH+h8N9h0PTpK5RZQiaa7W1LaW9b/MWl341rQAXXP6
h3EguKcqMsuoq1cCRVOuwmCZoezWSlzUNTEVWcFBH1fXhqwSjpXdRrW9Be21wtPcLpgFn67VVyq3
AVkH3l1u+zj1KwX4+QDb5lqCzcTNVt06enxlnRCu6muMqgMTi20MEz78UIIVHGmQXeiQgPXQ0gQd
lRGGKreV61rPbuRKLZ//G1iyn3fXeT2ZRIVRV2GW7+BhWHsJoUukCC/LeyiVvoOEgxSgYlis+ZV1
qC+YOFhJtWkN1yFJ3NBEhOZw8Ilfe2or7+BmE3A1XOmEe/dERnxn2SmmJ5tk2QuNEdfM0O2TkOa9
PCFvBIpa8O2fErr1CM2I0oitE7HymvWD9QX0IqRhTDC/g419nl/BwAC5P2kouvumrRueWprCDD2n
W3nc2xEbnsgg95CHitikAdlX0xyZ+IS2q2DuJfB4W9ChewDYtespUhEnEAalNFgWbvjFQNAB9O/p
u5QsLic6/vg2gWzpn3OLKJpxC8v2/FXbZSOGlecmVHoNKluIDgpbm03R2G89qQvcQ3eO2tEzDSjA
g4NIWVYUb8lQ4OZ+xmnspJ39FzTAPZWDWOSDLWIiK6sGytGvf8erpa2QSFp79M9hlHwLt+fnlZzP
4fMSP3vyAxMBy1UenqyyvQhcrVqoXDTf1/8LGcBmWZN12IG/BGZBEBZT9/XqtB0hEojfR+ZGeYOx
qecsBbZDSfn5XolTJ39ZWgPEYHMkTNNvuQ76yB7HYFkTuFwopTN98xOnZ4rdxUtL8CJU5BhqJ2PU
XW4uezlWCYRk5EaglVdjaZq1LCvJemBH4nCIgW3fjUk7nrrThNaxUC3iZZXx3hIrGgUTWx9OsKd1
jbrEqnd78+23q/TWhljU64vHIbyT4DzP47aSN488guQs9jFJ8+ZYHvRjGJIfaVEjzh0057DSYx6U
+WKdyJk5qasLCXLS9xAxs3k4cDAHdV+f6Yy7H6oGhGecC+vkLKqk/3Qh8YwJ6BWJCmG62P9x3wWl
5JiXB7u7QE7Bh+vtxp7gZ9+WVIoD2rkRQneZGyrmkH8ldyG7ZUfuea36UqD9CoKHz72gfryH1AWZ
8DDi7j0axkQPl8W1Ld2bZNwdYyzEdii+IRlNMEf+Z83PRhWJyOZZNnFHAVnpeaz01aYZe38s0pUm
g1usXpbSehbE+Se1KEw1o1xz1p7U9xD4c4+YwQfuQBDSWh4pwZ9VrjVjY4NdP4366p/fyUSzK8IN
tUxR1Jvxn6pMLcBwS5mlJPQdHrgCF658fbr2VyFQVkkXNXqGAa/I6oxDV7DirBgEnOpCOVgdz+Ze
EG81faQcJmlcEWv2/52x6P1bnBMP3UD/5eKPm59R2zDojL5mfo5RrVcjeMEnybadZhL6Rx+fOBfz
s4fv2j8DEoZ29ve0f5/Kq7UI28aiawDZuPhiq+1FO6F60brEAneuGXmeTlCnj01SZQHO6d5+0ns8
XHkh3WR4P2Vhrw48wgmW7OI6bTXpaNEG8HFytpxozFXk4iwOl28yvYqEBbFy7FOP3w6EMmlMhnMm
Lh/uRiEKFXuTKeY4sDOsBK7tEmSKPWVgZ/StTNdLJrjPEUsh0LvMQrVv1Wog4QBG0n9zUPNq4Y6t
j6DA+xuI2cCAeQpgT9ybJSdpjA7ua8WA2wemYv4Thgj7m8ynNzE0S71d76cPN3IYRAjlZjSGFVVX
2TSSmCfKs2onZyTP0rHM9I67Ppgz1+HtivA1BznqWQqhqJZV4p7DkBUxqu1lSuB0pBVhsyPJOA4h
F0pSQ4p3Bvyf7KsvhxMhZyUa+pysLT4uh1vNI+0VWf58DjClDh4yG2qSe0nPGYzEu9+QthwFEJc2
zyy2KgDaEaCNUI3eO4LD1nXHZUEXv4u4QIQTO8q+lOR2FcOxKPoH84mARZ3PyV0YY7dUGoqayJZS
jW7YRy9vwakCXFSq8TG2BYo1VeZWgYa12OEOhp4bG0usm6BmmyhUrjUGtYg2x3omVIVrZ9wYDQ5j
Lyj8Mer9/XvMWLPMpho/eYYmV4soyZQvkhKvF1OJ/yH4N/pbta1BzMREdxJuTud9M1p7Uo+YQ6iK
kSo0DAuqZX0D+4DC5fcXa/k+R2IU8dWC1irZH7S45NDFiiQPsYyxRGeUbcO2j9Q52QURJCSj3rBN
OM7EgMlPlwHvdVoE6ZB72vsxMQzyTUv5EQUkhXRV9FXzNb3j8GoC5yty08hghKdr3eM3PpLA5NmO
CZMQznpJ/nydUxoM20TMqhNemxOetfxzvGWfH7jSxHAcr+aEd8exDrX//9xn5MFQdR4kApJE0R4d
6iRqqNhT/8MOZkRmnq/KRD7YVq8CHeqREzG2vpnk2O+/HxBzkjCBuKSOx1EL4uj/KMRdUvJG8WQG
tGiCHRK4+KkeAAlS1pvGdu93nefcWCuBRNAHPTBbW8YXF01ZnJzKDTLyfw3h3+vNZMagn072R9kd
nAr59Ep68SRtWFH3+YDjv/2CETnYAbi7UMsmuzf4CpR2VBrCtlIEh4mTtgb4bDoKkXSWFiLgxwuw
v46PFLn+sFhsevvIFxSecdghWsLTik4Hezl7SpzXhEGft0XbPrX972RPt9vkLedfAdfUKa1LoVv/
A/+4l3YOGNALK2tdJy1sGtmNNFrMuAFt7zs0ndVhSI0+8jSNmS6CHaW7FLXww/HEM3dpJ5lbqxFG
FvWigloL8Jn/NbcYBE/hfDlYpvcAZny3WAcRF9LJ0/SDK1CmJdFPVDXC4W3lMwLDGacH7e2/tlqB
KSioNht6jKoO3iOuwZ/9mUQK6qyp25NEDkE8OcSnCklaVijp1jkmdVHIAjBRpwP0yA+wrEqvwZzj
CbtHgpdIBFHdm1gRY4Nmx3bv6IqKVvfdw8kBYEvGPJKjIHb1BqDBDAwIQYti/Z4V3udXeietmXBQ
zftnxOONxHfQg07PgXkSF2ttoLBoOlQEWJmWkpFIK0zi7qV6PK+oeWyVyx6+5MmS+yntbt3auFRq
mK92lQbi5P55dMuvwPdLwIxaxy6Vf8H3RK4+FrhEPxrAd30cXMbxXSskjJq/pHi79UYctgbxb80M
sPoEFDxifY4fZHH+Ms7vIhG3mQ8LE0PmsC2TDkIbM5uu8+ZLv8dScOlfUyA0KGtify2h4RTg4zBt
M8CsLIZil8o1kGNOKYdTO7uUirG289VZqYTuozYhRO814CiRgfoxJ8hxZl2BFS+nwfuWkQZamv+F
dlfmxZcxKuUrPas8E9ULpN0ODNJOf1lmhOCHa+BTiWCk7i0f3m5avNNe5vn0M3pqQ6u62FIO2ppH
X6XVwTsM2lFGYADuAtXE7AfR27Jl2wlfIpjFt+C5T7d0Ah8oimdgx8UZVsi9wfJnMEsYzJBwiZX7
ClTitZMmcevbKyHk6SOR/8wlB78LR3AeSBoYOQOkxiX+6+GOe53yy+P4wT8bat+QkapOmLDY5HXv
wF4YCqwiWBourQ/Ggb+Xn8D6qODRzEy4KPJrxHzPw5bIjkV72VcYB52brHIoXm6JOIL5HGC2B0hF
xee/nI7esS6ju5VDR10hI0qVFtPFlNNakrKsLAsy3xV3H5xRLlMfmRZZcWlfZCHbQZonmOcg6nb/
JXWorrQx3QYwJkRmqR4LPlSKmNkGc8mV+Um7j/611lr8f+nOGoc7PY4qkRsuva6fOoK8E4g8sY3T
9GtJcK/K8V5TZSl39MtxVPfWYZzzaVpQk86cwtWUFxHqzin5DkK5JEgiD7hnTYtoYUPyPaVqcy1g
A0w9Viq0IXYHQAlyXqNCxua/ccxq51dHBuc3SU8DLSha9MBKTO/OjIx8L9OdpNdFbu1Gjn8pqLc9
mKV8G2oTy5X3tOTyJpvtlEUEtj5mIYZP9xqxKy6nrtOdFFXRkCnx6uLo4BsphXG4ABeM/YqEPd7l
kjaIQfKXZ3Wp46/Jd3Ial9uanUuL4lWoP3fZIivry9cWEHCVHFbtcSG88oKRf8v+0vvMrIEZIiYz
ZBwqw6BZXKuqyd+9B0v/jHqSEnN6wWZh5nMzpwh4drTd9XzlniwRW/2cl693Tjbpp7P5m/pXIend
Q3QQj1EHxzgD0Yxy6KKVsPghtgWZDLdZ3Rae75CQFFkgNuUMwOh5b+UOs6owslpmI8SpXg2rFj8f
i1hCPzcudLx7wQEOVougA1wL+zcqhmLR5eZ3GgP99Q8GcqaKy46czk1SPpLMpOe285ekkj15oxAl
Ysgd6NyQfSAxijnqMqnvVKdFaxAREFwV5prAaIMQ5QJJx96vWG2e/BkieACGXfYzsU91GlLpq8/M
V+JyE4z4HYTCi1zkebxNH7gj59316ZnxnqHOwVujXnJctgsanLU+geeWxK63plQCiuGqVgwJONCG
9v8CheMSxUyMn+iBYgrJNJVQUPV2cY240m3EJfNmtZftonxD+V4PrCGWPHbt56l2S4Xq6nCOSg/y
sr7hndS/q+ijUvEZxsbAIyht2di7NPOAQ05e4D+ZAtxaNa43tClaSnPkeP+Ru+XGdD0NLHO5whLW
3zXTAwXZDod0/c9WUlux3Lpj1mACtwdgE60Vc54O8MCQPaPG1kSdX8dxolFjzxAtW/ilv4UEtiAG
O09/29n7WYtnRc1ynWoOfNL5SbzNsBN1UGJ5BoMd7sck+Wi68FMFksOodZPplpn7tUc5LSf+3AAe
hRqcbbgfhCLMWaibjyS2iIyIBf4zB/Qfs6QDu5H3BIo6G/vlOIdSjWasE5MSzpSsiIqXyFDwj9T8
6vDQ4+h1lEaLjxks+J21i++2USpz1ZvsAjNkbygxOEj1G9zLEhKUxzJJU3eTgoLYAN48mychG3Lr
GKxmHW2VLHGC+tkAxmn3/P5DbovROnlrcGP0QjZ/I4/5XT/xh2Pr2NXMTN34K9doH5H5EFaP9sfb
g5FBlRN4IQpFDA6lFOp+TBsVVMJ4QVFwSEU7JsC2VbYm1g8OMFwUaW+ONoJSzozr+fMUkLqcyYrH
5k2PZZo/VADNAvfKJRbfTPXkRUGIqMnoozkVfaKrBkrvI73GPUSJ+IkOW1R5aFAbJAPcnh3+mMZ3
VfwTz7T4r9CKAsIZlmj4JnBoUQwNX/OW8pvag13yFo+hutRj2LrcR2qJxtR9Gz4NWfhbyLyWf6eP
SoGmqiURN5huZhogyYJdmi2dUPJ+RWK3FcnlNSQ+42t/Yz65ZQAIyfJFI4HnuMEmTvplXnve2UZO
XkL623p+HjC/MGwA9cGvaGtV/BzKQ5w7SzQrpELQSqkrvEnFgLjhs53HssnKKbV/mr2rrmb4iVBN
VSyIZnKjuyvN4tCyhVvyHXtg7MSelDIzu3Mmywm2u0dBfYCn+Ps45M53D/QsP1NyCsA58rMXHsnZ
yUg4gAq6LNXkI13S6PLxynBbV7RBbcxqht+85v49MavnnSWfqrrhkNAkSCmKtjeHBu2e0tJhCZtl
m8omIad4hTErfKeoT7NqcwraeZvca3tuYfw561EXAceJ3n13ICqXwq+UX4+YT0ScCfCAQbuV91xj
pw0W/BZ54SPuvZuE11+6TOUIdRHFbqnKnVy2GCxdWrhK1CAmvKeu9hw3yGbRlIiaeTB2qiFAcc+v
MfU5pOb5PNWXypxXysN/jnC1bWLIvJt3iDE5YFxvQ2SoOnXmlSobGL6w5clMRd9V9AP9DnFrYtT3
AtW51dBhBeFEj1GBoavTo83dWEAetZ+BMuVr873QhGvzXkikXQuIB6lQkqXyuUj5EqjcZ1qu2mbY
1f3IXzsjlv6U9lPKi8WBir85jUvXO/ILdiyeU6M52Onoa2uKQqOdPE4YFnOPCuCtFkePxyCIQwJ+
oi74Hcw0KaeqQbwFkaFOICDKRsLu0mDUQ657TqlzHZGCi6ZvV4PTUdGYt6zXVURU6mkEeZPHR9jO
Jrcy8G71YTStGKJnDDu1IN5+eH79iDhfcuZk5YAZzErtzZ4iVfBdDl+kRjJQV8ZykDcB3RSaw6/u
HtKbt/Wc8Z0N/WTQmJCMw12x4FvrPwlTCme22fRFIroWjpDm4LgHzL93AnW1dJPF+pHHqRC9TSH3
szYsB5y/zYgC1jj5QX7mSbxdHElh6ZQbj6FpPK0mPnSO02x5zIyeE02o/dhzygYkRUaSjpOjVKAi
HOvE8u8Hwp/xkM0tu6srS+T+ErXh5WCwxpzIbtgMyVVDnQK0hcAGQUEaN7kiGOzoveF5VfNksntE
G8HfVAIq2d/FK7dTkuE/RREe8yVOmZ3aL27ErJk55Ap/y86tGuNbQ4N280NOyQCqAKli35w0AHeL
KGh/SH+wx45h13q6xQjmhbtSjPRgDamH9wWRcHO3yicI81IdKJMoD+Cgs7Pjv2uQsH5vRr+GbdQO
h8tTIckFHhJwdyHmrgvQNexAgShbHffuQw0tk/pNQekD74pqrwo0mT/a24U6SyQ2mIq4haqRaJBS
rCjSGnKuQW0UIL5aDxNskIcYDj5gpa3LAhHuKsv1kUYCh2FKRS6KR5by057sRh5gpZX+BojcfACG
PPx/jqxRu3QA8JZzVv+i5wiIFopdWOgpEG6fBtS59le7nH+upAUO52Lc1vig7O/tLQWgAuj5CgGX
hUFyXfY3/8CmlcbcEQhjtwQ1KjTou/cVrU/4taMnLhKBBxNSnedKXbnQTQ9TwUA0CdLZ9afhl0w0
DCwD+7WxEsghgWwwi3J2nTRR6ui4PN6ZDeN3fv7qBZ30mMxW2pszZkRw9YOzBQEftsdRjGOIohys
AokvhFtcROQN92Jwg71W00eEnydnjPgZbEMavfGDNhxclbE9/AbqZS+Xk7A7z6PT/4VqLZqsdlq4
Mh0uRSOBjFOQJPIdwQnDWqB219nQiuQBb8u4yFO2qGRXl3TsC66hZAR2zBg6oNf7Mh4asA76iGWx
ymUPNMsQnsuWlSiidvnd9rxBRgeMcTf8uc8G885aXZFyw7NkDcKtlJFpQsgcelCBwrYiyxDIx7nq
dGM9L5q/jC/7XQVGjztFqsHhiAEC8/sOeFbr7S9dle2uZfk/H6uUH+PS1O6NFWAK5Ot077xUCZg3
+VqcmqRiYcaCzsKwKp+Es9Ufhv3m9xiB3Lt7iOxcloHqikcjd/+ycEn31aw59sXY6b99Ml/478Um
1Ac0J212LbsfbJ9ddSDu7rTTAkQITrsPcog4jvhB3qCRVow6XsjAxMxQLzrSt0K/WGVgeBj/evlK
zLbuO7P4ES/bLdYUebEl9m45tAELp3obc71y2PhrLX24rngkyPzYpYvC0AxXNIiVtSrObyAxU6jI
jJploXjSswpymysukJSdbNiuyENO6ChrYkezsDEKulbxDk8YkYKsMKVYl39ZseW1y9e45Hm9fKpm
1ZCoX8hFOul+NDN4t0dmx7pUNVb1tMxa9o7hEfXCjVV41MaIjfU0YBvXizh0srLdcW7qNXNdPIY+
nMJ3pAkM7aIBRoBOoK7DVdDrjO2MSlpNzNzq82SweRv3Nj4LEY5+AVzqdauShbvw7cmyLuhl7VhH
t8qIvSJIY8YSolJOxJ87sahqVWLiYTSHmT2ALrXtz2OJ1LfoloKs/k7CgqSXfpIOzCOy2rvhIQS8
hW4q49fS9SiNbhUpZgwCWKTqgIX/QbguPrf97iixmSgR1NTVXWxf5B6ceLZKCL6HXKQV48cvnZPj
jWCbVVsPGBnhIv0E6At1O+X+ubD94BY7l0D3OBz6WlPL+wHFvOycgOnZ+Etk9qrTNAN4/8VrLhku
fSHKxdLZR2r20qy2vUodSNXRPLnL92at3GCNbVCxns4MC7mbvlGQsFp6dRaFQr17U+gL2XVZL5jQ
bkXlrBPInmEycqJf9CXOcm5QsYD3FeKwDX6NDmcu4rN+9PfUqUiWSV5oAxRqfIR2lxSPZY3tyBu+
p8o+bRv+3JTRrAxlQ2O4ZO3BYO3ToDmGUAmq182q+YhgJlMlhbYwly3FzwW2bs6DfMTlRTBG64n0
Ne5CmtJeGZxCKc7Qly8lZlj/E/++fN68QUYP6VYASPRMJYjo5FbYHEfAJRQPTBoDM4OIrAO4H4uS
dLKOmIBFytIlHx8agwC4HM8XUvZSmWoxoWw5fiaN97LO4lKroxRh2m/0vMiZEELE1GE21WRN39zt
3jVO/dnxILGyNrgMnaka+ezPMPmu4nswhD/qlXF6Ojiffi6vzmJ5g0wNlRt+5vznzufWevO8yved
gKSlhQx8pRvUuQwoTPVU7VA8VZTuNL9w/LE4+qb+haPP+1GH/Ilgq2b5xti09yPpk2K2r6wqTDW4
Bnr//gqtREwCi9EcglxHbDJnQ29mKAD4TR77nxtRA2Y4qUmdCs2taX1wEtwLoY88EJ9BmtFjsFg9
cOUCV6yXLkJGwRZ0wug8vZVIYohXp70uKtv9Lt+KiZvrPuezqUlnpBrl/BCacUkD2cb6NVkEq21I
rvFD8r0t+uqixQ5yxSLU6TraX2VPQxIkfIrhXZp6+ulvFk++leXfpVdsmaosFEmHK3R0lKs23y3g
Iz9Yb7MKpwW9FFp5m/dbBf+gq5GYPhEK+shvK3ShT3xyC8L+YzyaXHXKv1l2RuOwjtKmcz0loqFj
YGtVtAYuvk/AoG1x+yuA9aUzeOov/Ae8RikFJ372HdR4Jz+5fOfqas9CMasWdSqX0TQNJYguRvYV
hhKqDAuKTz+3+AhxtlWg48qbo3WkHppln64FYNf8sDf76zHbxz9gUeOmc6PsN3o0bVRply+oX68u
9qUlFJryzEcqwq+h1pJyJOJVEV/cBlkC1xkBTUrWtN+DeI9KJVnuF4s9U31cKYqWDEiySmpbto1I
MI2D7bfEyLbsKYRZfBSxILNpe3VeFDuOG1bzhxL5eraHtsHo2DFLDc1VBzz3tuKgRgkukwBp/bsP
EzSsmiwDsXPvHjXgb6pP6DKoaRNKReMTNEo4bbQtun6AU6hPhpVNb1YSDZBDcpz9QxkclaO7rgc2
kTQL2yHqDLhmjrNmWk+UaIPJNyM/GVmX4A7mc/5A6xC0rsn9/xZwUCE8Wg9Z1iqtKnY4MbPn90Sm
VApGfhttW9O7DNBl+yVDqdphclUvqlMMQSnofAtZLeMPlWM2jd7GteK+3yYAy1e7hiGkIarfHjuO
7v5aHZi73VRgEWE5F/3FeXRR5c3zjbjujH4sVBjvwLRwpvScIPmw28HswJmpyAlZEL7GpyvrXHjn
S7GIW9xLsFKWLRtqXuUdZo1hgZrZAXSC0pINF72Tje0sxhlVlrzrBeH929zXOZhHXijsqPvNhXZ/
4QIsP6Hx7KIsiwHVIxkXsmI9+ws7+y57fYm4LksxPDMLTpHrbo0teyh1FlibwlDJjdMf/6/tXN38
eHYN/F876y5MeMY8otGOr1ZT93kEiORgO6kmeAx8My3+mhdv46a0c5Ul+l4qws3UloS2JzM59YsF
d4s0rtQYeKRVeNAs7nHYm79U85mEf1unDkT3yEk8oxkD+3YHX9HrsHv4dh95BPS2BEaAHZlgUk6q
BliNnD0blJlb6eTmCeJJB3jlnrkuhZjJXnYJstaAf0cp/fM8IVTsluLCFCYrBOMwf7gg/07mjFO6
RoP0LVYNq3HhQqv6KAL8w+TW0BzLE5vjFWtbz8vGFtlQlL3LQQqQU8KKMgXrwR17XLpU64vXLVQP
3fF/Pc1g7i46Yqi/kZLwTRT2WWrX15b20HNKdDNFl9fcml4bqdfDrq50CfcwNf1w1NHOrprRXlYc
7MK0Br6DgaeJ0x4hi5nFSZZa//k2ykcqzCwhCgec9J8ljsgkUr1Ln6wEdG3ebibPhA1m0/Lr3bPs
jF8BEeGhTwOqAH6ReqEh8YEo6ckDn3ZgRlPjW5ZDV/l8gHHb/TSFb0btwnEwyVzMSabRZG2QKqwh
7OghO4hbMomD8KBwyBSKf1G4PVwAsuSn2rVNrH5TNO18+pNahXcyxJpmJGJbEwP3/Zo+6GqSX7JW
PVeF/LAmSKug1LlPg1i+HOXB3kyGcMLKTmQ63CJLUi2ghjZaoaGu9VnPfIrsuR+1XJskTquS7Pdd
aVZZ5fqn6IWkiBAcfF9XIP0A2ClQTAn+1wPWeil+zCvT5vO6CuHtHZJREbsLcUXW5JQDk+vTWspM
MpuyQgU+uKWFphrtxBb2ue8TtJV+CRpl074dzEmNFEhbLjwEybBj78a427lUPpmu6Ee+yh9Bwj3b
sTvIXRG+SLmPvVFSU142tIZ72TlBP+nX60nnw1hHfZKmhxz2G9gjdhVgUL8duTRQ8LQarnsoqrSB
iq7EkZi/O07+g7fzW8iaCyPAQJTH+LQOOKWHSDjxiMV81nA63757NO01wqwUKIwlqnC1Xedc9+DW
VHNF5gxalcSfVXYJHzmEj9Xm58mDNwqUb85G796BFxU6LUXeSFwwmMsZVg8tmvf+/mUG9rvq+W9q
GWygROr2WW0dPAGLfZFeI+kfdU9VqveM6yyf+fQzc9E6u0VyXOjf0oqnVyCy1T3tjqE6ACDWOMLt
ApLVB0ny8jWMADu+TAZFOU/C+DLqq1RkEJKn8aMPfotP1MUT3RlVIEDDRpm3h6krJ7aEsXz4CcT3
8jOQP5EQmCmw4NXtQCGq+vnk0emlAngMVqhhoBemTwL8NAiMB07fehWXJKWChbYWnPRvd4IfPe0v
HTlYyh+6ZkdVyTUc2xi7V6pRA1zdI4smnuPnSwNguj0F8vtmYTbqY3C5Mf2O87aJhv8IOMMOeEUh
CBow4C07WwgqR8MLE74/0ftlipAhvUKEtQ6rQFl3H9U/OUUHYP+W+Ra6dQnJ+3v4Zkr0aytGLuOt
7U7473vZfgJhFoqSNVV8jQLB2zl+XMiTIG3L7u02JGRUNjgsKxp0xHbJzNLrJjoWUif0MSWGVXKW
Y8uiGtN2WTIcGsMw0Y26m/Hw7rI3/Qu3llinFWZ+XHnDYMJy4EpnymrfK0AMHJ7wqydWQ+Mpo/xB
A2UBEKEN4bEKFo96r+AmT/ylOZ45jxlvg0RorQo/SkEtnPs0gALuoSfb/l5ZJADSC0uzd4zL46ou
HY5AVS6njmWy/uvPOdp2gawU38POwq8GmBpMDbdnYQaVqgaz/i9NSE/ImZ92ShZG0llNSkrFkai2
5b7kYv0btZdOt4xtnXnAhsxMlp3uQtEG4GuWwus80CsS5iyEdvoFK5znM56lYzHGKItnQFUwjxCX
fdNLz0lYRSjXir3EOOlufvZWFzo3p0MVfxELyqzauRSXk56jPIbGOkNdnAuzo5S4orbn5rYDkRfo
23XuJ8pNORCc6gSNLRqyjnv0pC4gAOWxeP/ukyXoNEU3dCu7m20z8wkGxrvaZwcvC+G+YS0TO1it
YY/RVB/jLVfKHHgJG3y+UpzJ3DixiI9o+FdM6ebj9TJPK3bO1Js1HrCgJHb3QARIJvCXJ0IWC2dt
qFRrpijv4LhekVPsFHmwPT9sFgz7byIqtUhtQtDhZLWd0+2VNK7mxe4WdozYkkDLoFgGDXRzD+0S
WweIHggGjSnLOZ4jcj9e6meND5dO6T+YkoCOMRvgmA7Bl0HzXvYa8Zd9AdR7D8/t0TSPCOdLunjW
RbHTWurmK/EmtWUMy+/hKN8VSk65aHszG/gCDj7QLCKeYKTrviaxlMnGdZVr6J0qwramdIDFWNY7
a3aj5IMCo1F0xyQvcv33eTy3Rsu7mgmYriI+x34mQhP1At5erPSS2NBULL1xwmLdx5MEZRMUBivm
S0gbiluSPaspINT8o9O/k+cln/kiraNq8LkoSohj7+minyKNVvA80d6Juksqvcj3Xp+UjPH9MkRp
7i/aL0fODMM7FEUVaWMKXQMi7ntBs7ZWrAH7GGMEtSWSiBxaDeWvrDJ6KVOjNdLIpzITGim16S3g
FaAqvJc7TITKjOI9BxomUr6egn6tZyrA3y05SdL4g77n+vv7aKfSCNDy3Ubk2Tao/dS8NuUGgadi
aCv/79kQfZkUgcCtGPrf9b45Km+OreVFZ+NCQHz2GrtFXt7BIK/AGaHuzjRrTD7DYi08DYJZLBbv
zQCP6JS7pDBDHiDvcckbjtSusc+kzG7H5QJsaUrh2IRabNNO1PCIaTKZ0rK2rfcwliy2wct5s+Qb
rQ9Y+haWGvWpEAcUGwg+K5AKnLHw8M7DaBiR0DCmqMmvPjfByrdR4BNxnWH+RjsKJUgptrDF2JUl
kb59X1NTQAWgJr9ilsmXVoQIAARLZZ5ObQqt8Etn4G9DVx1E8Z4Lv1krv5Nx3bfVlNRCLqh8tRJA
svbA3ThDmg27st5iXg5Zy/QYChtfnrXF6yP86lmduEdnDoB7oWFHghpUIp9P4Owj4xV6HJtKebQu
lbjHbXExYdtUf4avrPpsDpDsfsYmHdW+dFuqhkdAL71YHYrx4qn5R/WQyItWZTkSTwI3KdQPYSKG
GkozvGohfFccfV+WSD++ePjOeQuoFgkg+RgrPYPXt6yyA3DMXVBQ7eCGs+f+kI3HamkM6KmjvbDC
+wBAEcGqmshq8vtYTvODshqiUG8Rd9nTWETQ6UXDsygKF83PnysyThALGOdRUPdy0sds/GH4FgWB
qLa9OrZuz/Lp68WP93hyFk9dT6ckdiWP86huctLeKZTpmhT8TQm9xrBSpkarQ29Kbojr/MPvtHaa
2z7dnTdap5JNpITwW/OyW3NXRMlqelt18iNYVSqq7bnb4Y878Fzb0ONtginCwoFcVyF3ZteNlScc
a3oxSgDGu1Dj+//6J0Co/j+/L0XovBy1VBqXiBe8Yu1JIQn+l1c7lyobz9oycpgNJzfKenVMmWgW
mhYVV4Y1q//svKqfdbPLV5WR5yrEcrMZC5fehF0CX7KFnPWncICnWq5ApbOILIbd1gPF8nsYZnx2
Z3wWaWhJJWA362Fw7jPGchiWTR3mz0D3pxzVGdg1mCnjezuB5xDoD4irSZtgNzGvVaSHy7XS6xpx
P2S8s1nBMwZE1GpCV555aWwT8WLgwwfgEy4bGWeeaCj8FvXvVSsCGizDCBoDlqTliWDeIj+MKTAW
n2K3DSRz0DvwIcG/4nzKgnv9AiaRTnKi9YqSQRIYUz74CurBa4J9huaO774kJ7vDz9VxxW1GWA9n
SEEEhupdUFzw/W0YFFscpzffvIwQFOlo4/l7r4nt2Tsdb1V6pa/FkenZmKbOvgYMHriCPfPPc1Dz
MyFhVsrFJljY1GaE8mXC4DnZtdWl4Z499Vd1kX5Fsf9i303nlCz7defPat9V1zERFStXc36nOap7
llz8BWgTdkD7X+2Rby8u3MdjDWphr9adm8figpJTSXSCHf5tl4OytSY+JkMoABll+uqQyI3LEHBA
azjv1MmixAh2gX/loeBNKOsuRN3Kv97jOFUsF4AI5OwPlVKnNGLo/eyvmgrWFm1CityktlMlj9RV
4IcFdyTBo6jzzzZxfzTadRuJtBfFAiUB24K3LpDHRyNGuY2K4DE/QhYTxPXdtc1dKQ33AYR8vY28
Jz5pAl2wwxP2EC8wsW3VgoQizB1h/24T8EOCKsJFGZcVpImVzvY5g/mx1rsVgRURWrlpdKjt/smQ
WXbvSe0VFhZTRm3ltWhfoa6Nhoa2xi7NzwQpFS6dQNPGQJe31swuEbxLlX6LhvZa9086sXM23ieU
R3zVrWZehIRLWeSHw0S5g25BNosHOkv0HFcCfLTvSW9Vf49yVgeACZcZAsSlo3acCCh6ou/KRHaA
dIKiNX4uyr2bYZRf1dpIv00NDxTqENo3v0sAWxQ9ROzfqzZ5hO21Ke3ddTxK2AKuuj7Ku2SGVNoo
QzyPkcGWQJch1OwC93fvxbjjfVS0SrDiNv2eLFaU5uXXdDzyU1Q5TYyLRXN3Vd1v9CD1ftzfC6Y+
iN1Qin2ctujqWNV2YxpCApsdh1tj/D77DmVHHCoFpwqMtl92QUt3dL30N8sMhrw/OcG4uVK8PZcG
hnB4Y+bNUbEkhUm1exqaZNIb05QDL1Jza28HkcNS8u7LAFr45JLvTb4ZJmV4fsyH8mSrEaPZmk3r
hnZKuH9RrfjcpXLGoYVFrssv4ss7LkNtXHoArggfoyrMklA1kZeRAH7T08OAcgkk2X7bGIyMz0D0
eHLfuHy9dXblW+2Y+pRtY9HK3cOY9IVDaOL8LZGwlWy6xndie3punQb4caXNwIf5ZihbU3n03EGW
7sHPq0Sl5JSdBNHRBUV/GI+zis2z999YqCsK7cCJczXnpP+hYImZrRQkr1nmVoxplI4I03AIfIod
ebWgS9V5vWqeLSaIwyuMDNReL5mGFFv/KuCf5ZPhu69t3WJX4GMs7kyVNzMUsp7K0PHWVjoyPTln
KQcphj2ulRsnguXUc0dK5HR7csfwFtIe0lOUedcXdcpOKAcFMxZpr92kBo4CHZcIKTQ4qZ9K412a
14jmhGJYpmR7ebvr1vaRS6SXsDtnysOF3MtH80K0QLbV4F4ULWUvlk+HWodMm9/NJDnC8c6IipT9
J14Xwn5zd8eEUtjxhc/I8EZnKJ2xPOM8IisvueCL8Nyzb+sS7qRb9pxBSa1jYn9vv5LxYzByJSq/
PBTdwJ1pEeX1CiLtsJPhV9rz3k2yb3Bg4BoNXS33ecwVNuQs5c45jwycdOT7nlLDFycEE0S2E+Kn
Vf7qEubgXKxdtK59YYJ6LKyMYXLWERW2XJ2CoqjfvacuqcaLC8rMWAdZvtEWfKH6u7RSVqXGv9Pe
BUvzcSgRnkkyMfabF0SmNdWa9T2PUptndiCQ4lVd4V5ui40iJQt5AU+EZnGXxMSFeIorWY2KNfOu
a/mkP9ishmYlP+PjOOu+njVy8GXHK/U1gl9skCN7qcbPKK3Zws/yao08FnCTXAwbwPxuqm5USE2L
NsLC2iqlXtRAutMdrJ8IPSho6e8k8VwS/szn/JLxlJFOLiN5CRLnBjmctB2a2Mi9uVc6lLeWD96j
oMIAXButcgiwwpw1E8rGdMq5WgEF/ta3jaEk8eVp31gmxu2XgMYX00C/9ka3Z59k8NiKFmcY+QlX
vGYXVvS6J1yg5AHbA1KBW51eyHxPYv2Ay+aeFNcSBQQvukcMeCcjJdeYU9UvDNKt9Zi/Z9TA8ikI
kc9SxuHCuLWaoTuatnYxoc+GulrDX8CUpq42/HapMmjJhonNhJv5ASR9oytfqgMzNapAQE0VI87s
iTyAzFTdz3maU5qsiVr3IRx/a8WxLgR2IXUYe+nETCTWcbSXgfMdwB4bDNSDdjIyicLCu2TEfq9f
gLWQYP97/U5eVU0UczBLcD/cXbTxtXGr3k+PkDRiaEvudMbcR8B+vqN8+/hFrMW267GEXEGqZced
K0ItDS099xVeSaDFiQVKvtmVJoMTsnj9lbqwoKrF28h1sgNAg61RZSTiJdvn2PNa6WLthN0Xp6ep
VYQ+HI9GJvBw47IExdUQIBUII+xtx+3SOskJfT+FvtSoo8mek6gkNLfzjcwWMavgQGHHYYCNifil
FUbQuyMb2rgHt/pdGTCI8n7+NFqZn98J/Ayhj4Ym06VuGUC6xPVYXSVyTFLSWH3ByKZhEhGlOfSS
RlvyE2c8RxMlGkk3zuGhkb2TU3ByvfnyWqEkRmZSp/v7QHCrR9oKQdcHZP3+Jrp+WEnkVAJJW5GG
dF1DD5fwx8hOu4yTcB24ZqtW5SDKUwyny+fXneDBOG+iYhJ3ar/rL9E6PwQ/QHhvgWrPpPqtZSdT
TITQmg5plRg652pejIf7/xB2Dix0K33Qa+lPMSlzN+2pc+VH9Fv9SaXjAEUKgpZugIm4DTOG+prM
KQHFXJkogEktX3EvygbkBJCHr3boIROAC2G6MvClpkmtSvUNiKHEsh+cck4JmYIWoE7vRaQZiBho
WAwyhhkD2B5PP2OXScxI75UbyUxC4Lna2tmgS0fUsqv5e6du3nPjjZaQmCnZAYQSpJNEqi5GLDB7
dr+rtq2vDHnk8h6Wsh5J/BGpAJw2p0j6UqcjXn/UDDEJLV8V5PxGCK3pDXVaBA4mcNh3ugI63CIP
pWrQAlOdnSJc+pL9W0FCkDL1xBHlFF+LnfuxrzltBV7NoZWkA3/Ebj29vv/xCAJPoGSbzPF8xhXr
knfdtYFmL9yXwTbgWykpDsbOWE65z86lVo3PIBMtAPConZW94+nqiXbkmWKTB/TAH7Dng8PykC7c
il13s5yzepztvJtR943miwg9miLMN1c9gcKAAD4zj0/FHQGhirRIP0pbqsZqr3+waLhRV+Wjdmhy
JpPizWZrXoAm5fMhgoJ7CnVbeklwhQTLeM5+kr9Bt+TuHMS0JkgG2h520eZH0i5UAYuUskegFn7x
o70Y0+AGpqcZ1763tCFdhlKZWRLdarlYPcBKy1edO7ChgKQ5ScHRJ7l09+7YoTCX0NWvWGmvvaKh
M+CEDnoOdet4iK6Iw932pWsGnexHIcyAe0IbeCTx9qLGxe4dq+n6zR09g4JGyj20dcdsQi0RFLLH
z/Ui/hf9CZMAFQ7BEQxrTb5DOXRpjrcRtzRJqibndxPaRHVZt/2kzdoFF4cMFRgEcsoq9Wesk1Od
+/QsWtjUxl92aSh8Ki2D/QFzk4UA2wzEAAPUg4MyXfpPu3+IraztDeRf8ma2sJRPmkPV/U9Hqoe6
6Nghq09korWkMv9WOerw7oRBr+YjLv1iiJELkhvwIwbD8/7KiAImaVqeiPGnqqlUWhwIGd6iIyuu
7WCDB3fZ5iOGrJsuWHo0xogNi/HELfVNfLEcEM/0tRQGQEk9J1LVId0rdKZJ2UEpBRP9EiXDtuNY
9eTfQ1tG1/JYn5CYSdIk4eN0Z/n1uYgnU+YGeyRJXQU4EiRFe3FmbgoPhBm+stPeSYmELWS3wjFv
uo3MRAZDkobMR/whdKFi8reaKRHroAPE969yo8MkFqrk1qDdXzmWdJyWBru3Zo0JIjqJjw3Pg1Al
JS6waUccSYll2jj8yrzVq+KpcSiwH/zifcYozcCSJ6ljhsJYjg+3g5ChmLQkvwlm1twTyhQf5OoC
yhpIAkudYxQx6eCLyyQuf/vdUrBMwSS8nUX5rPC6JN7NB3V2E8DcFewUFBj0NwotzukXkOdiqY1q
O0ftFpeMRmNgasP186TaXYWOd6p6t0yXefel7+WULUXCip9s8ZYUX9UsoeFd3hrOODC3IKWTXT6T
zj+zlq5IvoBbVbuBgpk/9LkqMzlu4uf4cuglAr485AwzwSaffxGy7f8niEKbtNoihjBpO5aSEXoR
a2pMvkIJXZ4rF12cQYLzahqTnPGasUdC5clsQB/wBnINW3uE3FfEDz7jFWAA8QqVDfPViMIrLpmt
b3QOOQzta9ZO3MnWzXZKUZmdRQ1xK0+JhShW4pCdk5nR11TknR3MU8T1ZlZFqgQ/Lk2YJS8QEwA5
G4WzGGNPegSNXexdc8FOSZT2Zt2ifYhUYDSVmqspaGr6i8bI29dWIVfbHIdJQwtaDXr5M4zUTDFZ
TH/bK2KPwyAWx/QBgi+nVOUes6j6Fdn2KWiFh72X1saLKpx+KaqV50E+j4v3DYUKQPn64/BEe+EP
ibBsOcEPt6NxpgLPcHUwkgzJ/NJVO+ScHRpBpAnjMCdLGDUZLXzJmDkL7UAGVnusc+cVoqXm+gU4
MOS/w93/fmjNT5VM2Is3cBwnzy8sYwymJUK8EN3IttiCg/XoL0bkGZG+9qEDhDVgj50yh7lczWhS
RRq6DbK/+uNoY8kptCxmXAvoGH3I0Rx/ARFmFnnIEV1MzKa6Kh6+HOJXUChKEmLmnQmZ2X2JJt7p
22KtTUdAtpZP1oOPsKitQNAxr/6fqdERwZYCjBD0VREBilDE6lb8jNjS9KFcXtOXujc3gV9U9yx6
m4yOMA8dLBJ1cv1DVXSCVaerey30tKJR3X15SYXu8GQnbUaXqn+yQxTerEr81kyTyN6t1JaN/GoT
zGJFsyO0q2tCoyGgnpHgYspbLp+XaDRBwv5p8dMeZBxe8kCU0jWTOfldEz4OK5No7tPw74wpc8Tx
kJS8wAL+UHmZjwHHcLzBFC/c8G5oXiUlJC/k+oPPDOOL9/dhraFDYZk5Vk9+6YTyUIAPETtY3vmM
GRloFWT/paK2PdSx/tfaNbHOrDTecWo7AFu93bkWCy8dGFc7/7IqCnCgiwdpIjuK3V2coQOz+vYr
t8JtTo1g0DWwStMpczPDrbA7HyEgeFst6dllis7c2PEd4G5VqKdhRjy/tCk9TMh9bFrCSKdsRM5Q
ACs79bwdrZ32CJc3nsWrzIBn3uS7F08lJxbtxbP1jB805/lihTXbX8yGSvSjUQkrtAeJKDyVN5Rg
CMteuGGZtqvA4OWdYhQ/7Hs6pjHkTwTulpqj+mJVFT976lSB5mv/OgKELbyaOjRdjryDc0BPXj08
/KzanYdyDtexiyBpbCtlWWqgXIVRrdBhhbOJlvjJy7mcRC0tOcZsybCCOSw6P+RRYDmbR8XDe4BA
Kza/j+A40PT/mNkeri2T1OiKZrS/YCbjuvVixO366tlH4JRfiXbp2xkLuusGOeCOYls+0HBAzvab
C+JYFbnZbQsAkQOn7FucCsx3wrvgcl1Sd77VIcIEMiX/XnisYNqh5gyN9Q47xGTuQufBYkRu8dk7
ejtvc86JQJAnpGWl+uHZeB1aq1+8kaBIFeWmOb91aEUsNSLLrjEViK8hWRFR/4bS4trTsfZ4UhNK
Qe1VGJ8KgaP5yAlRuAiYzKeUP3w9AzN7KkoZWFBhs6LcI6CIhrFVr/RUcQ2rewn3gw9XC97r4gOC
7eW0RT8EASL/qA0WZvHv2i4g4x7UwqUgoWTu1KSu7t7kDipecsiDa+h2A4+ncO+u3CaCKbYj1NF1
wK6TB+If2i5zCoB/dL3RB3JNEgtsdAbIwXHX8xW4pm4DivJ7By3XtA6Bomf7CqnqFVWu/ttDB488
tngK4qwrzj8fx9D0urtgARjm4hbhrcLJl5kEVZhJQRwkpO5q3zpRA8NhlL76rHyDBWD9TlHuT3cn
N4wXM9WOhC6ZjNa53G7CT404zkQKd3WlVgSNJ44KvJDHxs3YFlRL0U+pR0j8IT66BoxqNamu/Fk+
U3v0XtMOAf3ZacEgnEKInOa0KfKD56MbGg/uIKNBrH1U1CaMJZXjb02U4Sg3xgs5cHenssCvpzY7
tBTx5o6Q13Y1NBqCTjiYp5ehwsOSDLv60FpjukxKmw7Xp8tQ1VAsdoSvwNAfwyPtSiSf5kNMhyt6
9du7jwqd0eGww+cZNYLBUVqdxqT7V4t1NJt2wLWZZc81JPrDR4YYcsXJFWPWs680cqtIqf9fAO0J
6Se7rfbzRNc0X9ZJnrfLdWOrMGPI2ukZkHSU2juMuAJxxFLTyOIN1xbK3iLDqNYipsTJ762HkJWV
AlQTqaSIsyukmJ9G07A/lmienUKyetXFz6pif/mOdt+e1zRwRQHVsqXYlqL4XQYizeOS0A+7NukM
PXflqnn0Zf6CjvkCGYSiTDcwsgjLUUyWOukU5+enFNvvvt/ER30lUGvGX6GFOx8ZIk8IfbdkKJmt
5NobxQbsf+kREhKnpbfOAs08WxwGNO8ltVt4+GXAGLS656+oQpUqd5zg+eALCNkrM9MSmIOq7h/W
RxhTaGxH3zgBC/C8guoUpmeIxc/6eYTI8FyN0oDD0ixeSRyNcLQWYEfIrPG4GPPBwzM5foguOl1H
rJpxSlKzHykb8iJmlgI6ajtKgR4/aMzOopX5kUxdTbm3qiCIzg+scbMT6QGTEYBpeyNQFuRhjGBK
eItbBWbqoBlpGklOI50+S6+/Tle1wl4cGNpWYUlzQ3F/tRenNyLOdWYXDJJpni0LjdTBlFEPZhOh
78s7RDzBSmMg6CLgYBL74M3A2Mo04PKbITAywheQvOSBMVv8LrTdVCRoLcCpxHOVFPn0RFz7WnF1
EvtgG5q5rV/m8W35a0jEBpsh/D2EkR/HzBjXjSFjWV73+fAEk/py9ThiY+v4lGmr66ufZu26VPXQ
k1Dj0LSe4IfxolvPteaplksLTKPAobB+neGFxIjZhYJLEqhiu3dOrbAtIefJ62yr9/b400K5xfvL
qnCiP1NKZVtMvE921kHOQRdazPH0yJYtC8eOWNYHYJ/ddHDodObTVg6Wuty5q1K4uwv8tUTCkJto
GAPvSaLfgIew9OoyM4FrfvaAMDEHbtfr6e0pBo9J8xuJzoML4cWKqGvdA46lqdXM6up0vaBIPfqG
6fkipakTt7+Ibx23aaZKpCBlhVLkbsXOKhTqyU+JxLM7A6wqK3sIrj12qHiV9lPJCCzcoakbYlIL
Yyr/xfr742cK8n/L3wehtOmHj5c0yItXXEt2A2IXCze1org4MQ5EtxoaDKLXXxXG7Sw+2PkDGS9q
4//j29rfeRdnw00lC0foL67XKpMg6IdJcPsDhAbi4r33BZ/pFJDqz0I3zPYUuygP6i6LSSxUW3f7
QeJbraQLGt9zKuoxXI/MI29QJL1PDB8XCC0yMYNApadfa0+ZNq9G8x9C11BvnjmseiEWyJ0a+p1Y
cOBZXZVn8gFcLgAxUi2x51WB452CMS0GtpZ4T4c8b3pYFaOcjw1SYmpflMPpdS/DWhiubFBoQj8k
MfuvT0ui8Xp4sj6hOxzVrKW48FNR7tnzWvNgzulS/5NSmRNEUS9GFdIRfQk8Z/lYZTjI/HWqZiua
70Psy9R3HPQZ38wk66Z3/mfSe+iIiycWHVffjrnkBXcJuMjpGh1MB3awgFrIur4RXPPTJPGf8gwU
5EetQK0/sCsxdgywY2ZMtAysHD9LNKZWhszEVuYzeRUZw05s+5gFw895qLAby/j5GDVqIn61kae4
cz5Zz5nTX/wHOh1AH63Hj87RoE3DLLCBFK/PqR3mGPFieAmdIUlx8lGS2mYe70MikKB37vR/vJBf
8a/DEy67Rz3+xMVpg0E2hVpj/ld1CSyvrIf08g6VGud0AohD0cEpQ8J1zSnMEARump0XHxRKcTu8
axqKFzRJE3Z8R3HIjV01OEAm1YlEnQ5JpmZ3Z3EAiH9FmnALGHnwPty/9Gx/uXuhqZnT3Q2bzQBT
ugUlq+pu5nkRGo2OBFVO+0EI7rZbbN+bOWLZuoiQbEcdrdQU1AfbSSBVgiZ8OYh9IWa2GaNRdHfx
QdS+Q3Bn+/H3nEvCMuLUqYeBcJ1ISXhBTRUy024k1Og6GR4NFvzYxwog5VN0QESO+XsVzGeNnlRo
FaIv4zI04SGYTwNSzp2iA7emICVaMz9hl3z3YTjwNx376T2afkNRQwicIngQ52EdgcN4WV4wGjx7
gvKeOyAZxTE9H0ssbnAPapwjDuBB9fei2xzQ7dSSa8mdnLVcZJoyaPJ3gLGPDc+Xl2F6aQvvNYtx
g65CUoUerbzFh1l0HIOdj4XyDk4Zv59XnRfX0tmcs2zORzz2IfT5eziUTzP05CbUvDVuX9XO5mHh
CggaH9nz/R61DFfaR42wd+v9TH99xCaizk0sTzQKcHln7Ak+LXQz9ceiDx+Fu9+TRRn/O1T+B1+3
h0OYFeLV5f/HiYQnihrjb5zJdBU4RXJ+K9BuHTQxmJh0F4j5hB8y7l3mP4TV9EUz+h9wr/0kWVGT
P+gSqlWUOG3s+fKmaMS5QeorHSbeADGzmUEnseceBGLC3majZ32N3z+tisLCn5iRVQmIiJ6c5HbJ
YQDyLk16NCIXirzq/5u7k0XLIwRpyW0YX3hFwWrCjJDPgMjOnksORnue+135xcDVP1VWIH790Cyg
xfgzck3nwpjuteD6XF/XXq0n6IkLk5eUAP7AhwZ1j41CP4++OwPlr3mddVByNEq5yK36js8I6oEb
DvC5Mlq5lvgCqjmyVIkPoTAhUJ07Dvdw+U9NNLEcza4OjBPVk8IYl/tyum1tD/QmDLgAtQY3wI2J
XGxHQPzD1JAgcl8jGbwok3kcFW+h/cd/iJ015j14tfYMz8uWXO8Eeo2HVsm1d1YzZl2YcCEhVS9j
nI4jZPFPZR6dPlsS5yfZsTh8VaiB1/fCofTpD7eRdTq6Ez5FwQA1I069YoxbfkQh+4dSvXUfUrsg
XstBPC/SxML5zmqtkDaEVt0eAssVo+qNfoWHuW2AlFJVYu0DmFOYjlV8lT73oaaz8Mhq6+YhbhdJ
bBu6lfnYyCY/GGoK6hJCsDvXrBv8IVTQY310oxAevQOeV0YUgQ8P5WnQnksBxfNkwvuPpuYIb/Nv
uoJdpVbMz+VTCc5TH5Iyzf0QLcAx1S9rF9iS4pLSQr0/jX4n2KYS28ZF2GVJffK+K3fNolzrEkTX
NfjjZHjMGlribvUHDuLX9IO5uoc6CysYutGi1/CT5/pFVVpfogn/TEF7P4yR6kznWIJ7U0NCuU/c
i+vrU8U6m18dbyWAOUGokGegXoU+EP9JuCQRhLZ/IIeNRfUCkgpAA0ljFGlxaQlNXgn1wH36DP4Z
rjMzYAaJzeLd5iJ9KJ7yRnVfGEQ5r5dDSasSQ2hubr1yY0drlcEcgVD1UPFv83amkv9xgJbIR/hz
Mm38pHHN//SF4T5y+2ZDa85CakDPrf46p4HhohEDy7UYsxQrt2i9c9Bg8lVWJUCkCEG7XqILhLv+
kIN8ySPjr2FxI8dbjTLQHgZ5PBgzx+k45GKsahytxmYdaubx5bl+wNpeD5KoDbhiqQl3ovefDYD2
1zxqSuaGsKCsKGmC3WT1GZuNM4upbitVCP5eHDERVb9XjhSIPBO6ccfyOjiNk2jV4pedaTpp3g8L
dTAcB1owqWo1POFWm7dJ4OgLTMfvSypanU2yjNPdSGW9kGJyrXDajJTnnvk0n/6Zw82v1jcq4U/9
XB3z+2dQRuaiwCf3Un3OBg23jFgmTaT/6g7HIjGCcsv3aJCh4e59kQS0vZeHn1EFCxPFTwAOBQM0
VMRK6raiBpzfzu0RmR65+25mfi2XK9kfMdiqdxr02x+JqzMYKZlgnYdAdz4jXglITVM/h2nUsnTJ
WownW0MoRUerkTUk7EfsulXzkFgr4kMzoZjs64ETkFdWbVrgYXaUBU9KfWqSNR8KlNP6pNOkPH3N
Y8dkgpmawa/frSa4WrjniZNhsAE2ZY/ytwsQUf2I4btM19lVnzsZGlJCgy75ViowEOrRr2jdmK2g
WP7Vkt7odMcBxoNHs4YVv3NuU4TjduSZjqEg4gnlDhK2D1OQ/yXHZJdvyaqBGr9/k0li960vEknI
dbqU9rRlCHWVnReT8sMFa+DSMFD137cT44gQmOCnUFrii76Z072tqQ+TdGqBSynKXqxRc7NaKtCn
UThKNmZG1mqRBiLE2GbXY+3kzFjVT8uYaRYtY6gmwiMyEM61oCVIqEyndg/PhmYIEkqOTIJ8xbDX
e3Iv2O1SYk32wx/YMt2rHbjaQLshBPAcKLlCNTnW/mQFpuKbcR9B4TgYZ+8FO+xhmUAy0/uH5SyG
quO/mbPjuoxHzhLdE9aHMBFV3CcjiYQstRBTUhbjBxYiERrdd7wzOPuCDbisf/Dwdq0XFTCJJI8V
/fw+OSlOEvUb6KQIwWcKpvudSNXf5OoRTNpm7lo7yrtZk2AqdFMJuxq+HA9IBRm2tlCdoFv0rOGr
jMMg7eKsKcNZ9bu+8Jd5biwWYQSl72A1nFOw01pKcW/79/iQVsCX0p2GOKFV/AelZSehpLkUYJLS
dxYVPq0VcJXgMcLamJHBJES6l7r/Xygt8kBtv6Z8BjLUgxZBBHTLmAOEv3BPEWFvAaP/b436AxG/
jPmVRXsUxqMfW6lArvMTLyxjdLXwDnybTtSk9JLH/Ds01R7tWB4pp/fqDhkVwKkzcKg8u+fV/Jv7
Xeq9jasQ8PLqzlIm7deX6bZROrbsL6f8r+T0e+B+6wQBdJYhh6WpuOrb7ynpVKy7qTgC1RY0fH6/
cfOe2rKfLyHNQtLKZ6ZgsSz685VvzIIGwdN2KqQZjvzXW4AB8rHqUmtIeMGJqBXyQSD1kLxWlYod
kj4Szk6/PXMhngGtnV89tMO1rY9sSMwjoH8YD1bjumvfZgRYXSGVITU/DF9x1PAitQKKFdl4lNRL
Md0/WvdSdX1jxN9kD5q73PHIfiUdlXTYDwY3Z7EYrNtUBNEVEOOJZ5MlHnMD9jJsuK7LqTmcVozA
bDhtqs07AJKGVxk0Evmm9pIIBQ36pzYROSMilsLogqydOL5ljvejUfCQy+F+jDnsYy2c0t+kyeAJ
gGPBj6UxMosnENgQhbZ0zhvOEnVzMPvUbq37nkWoW/m/oq16m3J68vH+TJVbVuaIrt011q44tpPs
5rLdztmtT0RjmF3ACH6pHnVHhP5xm+brVUvGMPjvZJMDsqpFDEmnddOHfnp/ktJQsHPR8cPV6JGu
XlIZDRgOF0Mq5Rkhly5Dwwggzyx/t34r4MxWu9+TqBkEmx6iCguA3q7UwF3rnYfqYi//YV4x6f5l
PCz8ynD81GIr615hUugqXxnx3nMlqs29m3JXTwGhwZ+8Zgk9HIrfr6NyIzXAoIWdlZ1UNrRZZA9I
MosTrrXnU3qY4lcyNW6k7FwItdXs1qHh+D0i244fLd81f5HCSrC2AtXZbaPBc0422cHGOJY8aU8S
YYGMe8YLO7+jTcOUQuoOFVIMLedy586WPpB+RTD6pT/LMVwT1+xYa/+PZJuvz+XIIp3Vc1Jn8m2w
fYfMGgIHYMmTfUObVrMqnzIberRZvVvM3JhQzc7UaEomAvLOLt+T2ePPa/bVoVOg9Hpd4EokUnhf
5JpsVY4YEl/IYsUluBKQUzjlcQwcF9gWHD6JPNHrEzzs/Xb7rjzfqbJGuK4eAgFfTtjXOOdD+n5u
3/dr4OaIaIGCjzA+nE8dI6GDltB11xNizysXLs496V7wnO1KVlsnZMY+fuiQiuivo2QNqWUOtMgp
YmeED9+h/Y3NJAteqx/2rgOggMv96WDpGkAU1guKEMGkzcKZjtG4+p8MiInYMMqaRxKHGkfs2gdV
zbYyfTWd+iGFxnnWFUBhBD4YAzh60TzFOi+stM5kuF/fzIbjWTEGl6FNvhPpe718HJxBK8De+GWZ
qud7SCvXC0oRiFj7I7UDZTeFNZeRULnmSZLZb/yrkDnRVhRqE8zSiGJIKVEBWRedgRRlyMfBvbuZ
RYc8/l8rJ4IqVuxfaSL8+gHqRaqTMTm9jz6UkFZ6sgGir672s/w0+MynNQiOqA+Clk127PHQgHYd
FNlMQ3oZgoA6FBzFWR3QYxZWiCrbEVoNpKjLxgvW/kbL4syYlvVdUyC81eibwbGJuf8+EYefKXV3
9wXTeDPNNfGmvQqguHmptKA53JFpAg526GRqXStYjJcHI8AFYQLVYxoDur3D8Kl5YUCJ6h8A+O3I
EGYpYwuw+Ud/nHhPTVfWUcpJesxxEaz4jRvYukG4mwto5gP7zHA05Ubjq7te8haH16dHLGanZa0r
eb07UuJunrhNdjGFW2JTq8dKPrivU9FJJqopZgh8ws9BsUvgPQNfTW7sox6MSWGY2mZuDXXwhSV6
QTLJIXQCWa8fXFljKka7tYVr8Nt9n2Kt+ZdqR2MdatymFpwJT4FjVUJ6vo/GdeIuHXMBAeWw1aFV
VMR+tTsfMFI28/aWCkbt2nB785ZmHJjPdeQxagzjqRflV9SWm4RhQ73nsXCaJzqw/BLKNKWI0C1G
CGghd/zVuFBtYu115Q60UiyYwxbLMmR+GuWI+5Aq4n6W6Cd+EH7JYOdyxi1VasGWaM+74EnhfkMv
Ep7JIjW5WqvlVmxsEhrqXnN907gNqZ0eV+1FHZVlBVVHO2RPlhGbV/naHexAYWc27YfLYyVLd6lQ
O0Kp6eS0uHkVo7mfSDo1/usZWTHfQsW6KPRGrNgZZVtgY3Tr6tsXJrclTa65VyTR8wu7wV2m5UaP
pO+37LVEVNG9f1GsXd7J/l7441ED+IvCQ2bFiYH/lKqNx0ZVbEOhLhkelBXCygnXnHoRKkXTTv3i
AN0r1VKdsdGo2OWglIa9OaMLg05ZEAk8rVTVuY4fNbAdL8Iil7H8fFt9hoTT0Bk2RBiyOh7XJR3h
9YlNdGFxNU0N4+SU2EoviMaL9kGGWqIIIScFhebYGIQVGL6zyQxH8kaET1OPSAI1reeQuka6mIKV
m6EVeCmbm1kPLRjzQVyfjKxci3IdlzcFFUR/BQLUSNDIgAshyz5tlavC89LDvZ94xqZLn4iwYCVL
MMRnqeC29xC1QfcWtCRtxcunvvL53aTSHVr/79qhdmRQn5ngGhz+sGxvhcaJoR9WoCS+dlrLTpdS
JZTSA/WqIGTO85PfJr5sl12hgRP42C8PtjelTrFBP9tDKP8OlvqkWb5UJ55iTztgl9qk/0/XSk00
akwUtxVcR9X+xfgqzGh6myLTUYKLZh8rOPLSBsW8EUSQT+gwv/0UBoHPuc9l2lyiplyPvRJ7QlLP
s4YrmwQXxyYjrRwCAHwkFUJ6ClcVyMiTRJC0iU5cJ49VBlEON/XQnDbCjVDVUDSiWrhuLYmgr0p+
Gke7tHwCBOb8zPR5n6lOgAg3yxgdfgSglbgtBDymk14nJT9TUW/Bt5Eb9OCeK7CUmPT0X2qyjr/9
aE8ETc+qd/nLMEtJ+xc8XZc3xAoJZVy81Rj81eAEj1RSUz3pqFyA9CDlO6jRbBMo579MubK8LU7Y
yH6xgDComn+d7Jj65pBpgjgPJIaNa6SxrhAbJot6MD9TphYP8BRryWn9zoq3eZXL6O4panIU4Vr+
M5ZLRe6KbNVXgwEQt4G+r/hyoaTIRVRUcyu2nk/Ua8fEHybKdeNJzLBiX14NIZwsnCoLlvdg6res
lcXnhQa2bQBL2It5GuS0zvmmVk8cMM8SBrt/CTEA9DYI6UnSi3TbNr5Zy4Pt1TY5UmgIoiRYfFxY
/IxhrPs1k6kHBH8NAv+mKp2PRy+oX/h0120/hNz4CS31vYiqU8jEADoN7R55SxEl8m9ds16gR6Ev
BHdp+DYNYMTzhe3bQQWupYN+z0m6L3un3QU7YPFPnXPsWrBkgSHWIz4WePBUcGvRJaPT7Fn4vIrb
KbCPVoONzNtrWZ3bBvnQ21M4IklgZ7zQdvudRIPlpARPSKAFNskExTy64sBR33R/5yuvFiU+2T/H
8S28qhFuMag6IHrvnJqPwrXg32y7VCcRJbLAWGyUWeQY6TIpNT2T9O/rLxOz4DuKD21wPnp90qDR
1nZWvAtfRWEYdUVwbezrvRXP8BruF/HDzIH4zVXArSmuespcM1srpeM4GhEjg2mpjkcJ11erFY0x
YL0pYx7OzdtfX66QoOHQ33KtStvRWQzrEW+LzfNPrWGJvwShNssSAhprKkpoLmq7harbdrfVMJ18
ycPniqxHCAjTvIRXHsnnxEhQmWyAE/VPYLkeNAu8oWooza60j3+x3dNAv647aqLu/GsjZIJ0BDhH
3nXkZxGYWScuCTIaLyj3mCFSxQZm9SnftLFun2jR13+8ZeJQt/jRHypOwbw8s3ETqEkmhcdGrGGI
4TUgzWbZZ5ZVeg3H6KhOmuul2H8W44ksPpn6PLtpH8ccGTYTgOu7CJPEnvDu6uqHD978Gm7u6UpA
iLfh4CqjRzKF4bOhGDlVyDLykMhpanMOk+yha/HfRFCIBsDcRMwX2LQj29jI8JivEE9e6wDy6+n/
66LR9Dpt2uwORiWymdPXvkCzJ9RgWxaf8vxcZnHxp/E/ClCcrEgEDDZGzoT1uMm1rU0HcNrHJnMm
5/qkpWoKMBv48OXbur1tBmsdub0JrrM91RLd22MhYg6IfqTlJcAXHH6dc7Pth7GOI+FSTqf/CZEc
tZKESUKD2vYZ8jX31PSgzVOBqQI59W47FmbQkQUFuqgjoNTrTVaNT3Sehu9ujzRdmPVTJwXKrPtg
7kB334HJyxtuJTpsskpJEGha0PiXfNnvCEACsTH7F+Y4WBA7/ultt6wKfSJTyZcyRKN6gJdDBrx5
GcwWQNG3Nysxw47v1t4rJNQ9DVjgmrzlLCmTtm3t/FC1oPrUKeid/hVxSDqFQh7wl7ttGhiIZa3R
YF2CdjPCDb2yyzgZ5RmLHdYsyv9kMOSk1X1Wv0IHy4dOktoTdr6be3F5qtDAoWvGI3mk5ABXbgWA
iitHOCjo6sZkwKS43UktHDMGPyTNVhqj1XFa5Kyn9GEsals/LGMqreOf5WFrxxgVVk8AYTcYG37K
Wk/WQqh+z8kpq0ZVy60iIwjv+dvZu7t2gZCIAKaLABX5x/VIIbn4JlJfOkztUip2Ah86J9tmDDlH
dCF8ve3oKosY43jnM6q69t1mZBg59iTE87FUjAoEOCMbqCzaueKsR2Omi9pmJUF9OLQbi7jK8ZQJ
loTx9WfxN/QGvNVjtLA7qnsGVSZRidJ3RADnTG0Ztzp8RAMME7EsIumBA1wIX43rnMAC+ONZahLC
VIzYLzx5zg/1kB5Cn/he7woVR5azCZZiKe8/5nNOwkS9gcgZ7V7PZG7WSWZGSEnbq1l0hnedCERV
/LwXKTJFwzDcbIH97YRHoxMOwXI6DeDrlnl+AH5/uNxnayBvxOIwPFBQeA91mMd9KFbD23RVpUM7
5hJG/2bFQzIiPRLG+rfUf7hahSa6+VNhfo3cSigxNHpWyo99uPgobFj7hUv65+dDXHbyjQo8zWfA
7vhII8lW3mMpm4dApelO3IieNUpkCIOAfGnw0cxVq0/WuVDRLc0RWtYjQAeBhGpR8Y17Cj2Sugoh
aqOaEmHz1ZebqDz6GM+Q98ZyB0ZFNjlMB87s6SFw5EeuDMDAVeFj7OaV9FKl60F9D6/SLkc0S6Ku
afmJTy4AduawNRphh/4E7bCuKyyg1lhbyODqqJa1FHXHI4QOu1ASTKXjW36+plPoI4lxkLMr5zTJ
7vqq8c2U5BBwin+c+PTrUH6fYoarXpoyzvl1vlXliyOt+fNNupkmdPN6X9RSs2ueJFbhGfbDEag3
M+b5Uf43AiwSm6N5PX7TTMhMW459m/ZmTGboetT4XI5584rD2DOGzjbIaWVef0IHVq0pwvLiKhhD
CDoFL9s3XdzHZ57epjsk7xMw1ko0NW9icRct2lYEK3GQtMbBOCDs2nZRupSfKjcJFSTFsNq3PQAx
Vruk0ZnXsqSoO8s8Tu0Yzwku1Ty5DsCjOhcb2tkR70eHt0ZVSSCDIXCiFr6wLk1TjrtuCtb128ek
D4CMkzD0YCmIj5RTz+QAmMwkUnh+J8w1zg/a0Vp7CAPC4pZ6h1yf5ELw3rSkxve4qOr8mN8e+8yj
QVH1X+PbyA2WY86vgiCtga2s3tJQzWrN3Jts1pSEYs6AOC0644vLNpicv0l/yNpWQ/4ZyAfVzK4J
71vpbYRRytc4QHocXggS0DsxPWJvXE9ctIaj/XpPdcX6A52yIpF3kSuHIMLm0cR7UUYlf0H/8G5u
EqWnVptflsbPFjmNPd5JGQjgIZHD1BDoQxIRhNnUtkvXSkeHg2Hp5kBqwy6X07XLY+FwyHb+zxHi
NW9VcX490sVBdKnrZfO6IUknlWcNwtJ0ucC2MbyMPxYf5HMuUkUaOL5Zpiw+/3thrlXe6TMQUYMX
3u6vnlf4KbqM335zca3wuvnr+eA3T8YcbvKuoiKdjdzoV3YR3f7LmKhm0yxj40g10PGIyDF5rJnJ
R6TS5He+j41ieCFbOfHzpLQWZicUQA5qsXN4vfc/+A2dqa+i8Ta5H6AMRd1/dKfzZPDUYiTp2/PB
Mi+Xvw2xLgBkQdn1BkUdXLVAZH6xlZzf7SYF/ZROBLiqITfbBxacfNbxkHxqPxDC4CyDZVpEiVl0
ZsfD17jwhidGjsuM+mb4awwG3Y6M7UiTxb/r1VAZweXwqFlgEuLy3Dwbf9SbDJburczu4SRMwMWs
IiqWOk5qL0u9GeNwsuq4u3bXT+2iMPM/pfRj/S9z504W3fvlbQ8meKepndinWiePSzJFQ67gt8kc
njDSE/09eWSLALMqcHzSCt0hk1Q4HMEsUPSWtvXKR70Xd7J6o32Og8+jS18vt6s9goLvpr4AXPez
mwZutiHRyEFp0MhP2mb/3/eduT2cogJ+vW3VWgKfSkJBzz/DdHiRMdhjSH9L7qaUJsCrKvCgG55A
PCjZtiz/0xFsctagn8m5EwMYIE7eqmUHAKdIiGYhQM+N80FGANy5xlvASsgfVZoqPsAXecpx7KRz
elI+8U86gduIvyfba9hr5ln0Cac14g7bz0NuCvNG0BJqxgkH8IxnlxDNSiVnLyMiQv3TOsLR0054
vZZOrlh2aril42Tx5wXOqd2wOexodNHSX8/OO/mVXm3MQryrZK/XkrfA45U1wABWn4qqqcnYPoUj
LOIT7gjnzWU3hvrV/YBgrEDWWOhnESXvoAp6iFtPkIE0zPnm34n21fbje8WR8o5PCdcq7xomcI1V
aZ0rQWt2lscRgxWJoBKrjEj7F0Et094TsZwUXVgdM+MLSlOqSXLvgjb2RI5p69B6bkO9TPObmfEp
1PsVGl7ItLpHsFoWxce9QlCBJs5HLaj0Q0PXG9XPyk+v8bu9eJvLbDbvxTf4ik2QBCYRygQqCXXn
gHULF0aWVvtEW1iY2+JiQQMhKN5N1T/0BrO0c2KYesnNbLGG3tLCsEMnbFCU7bs6NMceRGx8xjPB
5/2jZkzwU05goY5pKMb3ExfcMiS7DCFZP8Fzf6OnzLlU3L9G0fp1uML4QSmJeYkp45VSSf2aEVsi
YPl97fkWrjDq4gqQiSaAiF4H5llqQk8CVmXSgVCxzlNMG95nwGju4IoRqEiU12Bar1+if18VBKsZ
50+ZcQDC+t9xQe51Qo/u7unAyP4H358fG+ZCHQemyE/1MZKB/Y//zA6OMuygEIBYPQQKNWv3HYLY
xu2oj/Vs4NrTCrnzpsfAbUDsNwIg8+Hc+MuhhPCLMXSD6IQitWOWi0Nv+7DoWbjzkYUSOXlinng/
7W6Zkg1srr34cAz3xmd1d8s/QM778i4NUfk4IVTsz2vDgK+3+v1DdT9qayLBWST7VcjHeAf99qrG
liBHFl2+T8IkUgWJfHYm/Bv3DZIXpXuVj3fhEUe5Lndh7+DMwpHnPoXo3at6G4Z9ZLgcCraMh+0c
WmHom/Yhlm4TePORzMWGMDAqwkvIh415zhfMaIEVGSRN1AU7u/q0YpbWCN4DSbeILIU91ZxnbQsO
pkNVeTg7gF54WgiGuYEZtd0m6BCBUM4ltX5eFidqJy2sb34NWx8HeDvee5AUXopzASucAIgWqXS8
Twrrd7lrkcOnyCcNJNetQxO+ue05TErGNj/nlExa4A2NrD85QBr+NSSd2jSdMjQDiHJTfTUCv9R5
v3tPr9x6+8D2UrHgQCurUhrHBGhvuvgE1rYz8r3uAfWSgBkVDkjHgx5e0tE52sM1lMGKegNgU4Zz
XsJGqBnaDpuxsUYipomlfbmMIgREv5BsoHAvEljb8Vcr8Nj0xIrwFItjSrpU0j/iiiuilpE4ynNm
oYqNlRy5S8GuiNEr2ETuqXeakyOA5KTI8V61govqU/gA8vphTXD0qHcj9A1ajwEF7wShmj6BNeWq
Zt9MI2sSFTxh0IjqIIwGAT4VYWfVeGraK9kVN+7M8otQfxvv5o1bioxZDrleBG5OcdgNqNiukM60
+gGwD4YmPsfojj6YK9qC4SvedHVabfdLn8vDkZ02o2D36APQuseIpaK7NVUXJIjZO8el1rPpZ1Dq
GAJfPiZZfNoVDw+iZBSeZ8u0MepH0TDlThR8Zsig5RKWby6kHkgIqMUTSBk+Q85KV4T/PcJZZUvI
5oxD9jpMJBU5Snl+qBRrCBo2PLv/G1TX99448L7t1KYt6Xoy9J27CF80MICGb/DXfpq/Z3IEnvcu
U/dIui2NYxNRNOEu8xnr7cBYfW0luZ3qQRJugd5F+Vu0ENz2T2eB95woxZZSCGnRFKfusGPs4mOv
lsBj9Rfl7x+m6ETPOdRnO4+CsVBIWOP1it/t3FvIzBSGDD9dHiSynsBwBu2p3h1+m/abZSeI6/SF
hP8hNNscz3Rkr2vDQKbFuIY3qAQilMsw/McdUEan4wTtCnBCGL9Zk7jCDl0nedHRAxlJtqxHzHdI
MCxc44/FTXEQv+XX0Vflonbq8vbbezw4quVrKRf/uLmZzsCpm6YJ6ZJteDC5ZS06l/Wg7wkXt/6t
6+bLblxjNVPP/5+JPirhHuuUguRf5D1/85xF6v1jwjGTfxIZOdfZ4+5vpbDEKuxrDFLuPA2MwcOv
y5moeu4JII0S1D8oN9xEOaqKpqaRHTUOp2XbLoOmS11Dv3haygAh5RpBC+1NZyJ98gzdroR2BonO
mpxDoVglWzgVZWMFmeuTGAVa4Zml1BLx0+5EP8yerbHlIPcdcusXu3GymFXJRP93eLQ6qz92BfBw
1e782zBx0qpX7ISfhTsoS9ndZXVFN4px6HP27Bl2xo8W5KLm0trNhiG7K18L5COM4Fk2Oa0gqUzl
dAQJ1OVzKVHVFi30clNpq3MJP2+bVgusnRyEr+kvO2WcvjijZsA1L3K3kcENyImW190qTQ/k5BFC
ic/02Isiknfk6bYmZE2dmq6jjQgT4prfgEkXRdRy9FQHd3GztTivEsnG8JLBsCHDe6sWyANlnfTB
bfzZ2gZtEuM6EuU53o5PHnxjq3+6uIfVJiDbRZS1YhhkkqPrMcmNAnznWsj93IyHs6hDFrnd+MaW
1bSpNhQAsM7nccT0TwweB2hgIkvmWPpPybJbTjKlRRP+nskOl32yTygB8PL1XJ3XNyYUj8I6L3KR
s0hIO+Z7cHbTPmYod6VruCpYcgKjyjWx1ZdArTfp+BZAZIMnDk5wjuiccUsW+gFz7NQ2xxiWlAvM
cSwQdAoo6y4rffnX7TB2zDmxEAJdJcTHnGAsnNnSNYOH7Z1jGUyTomz+lS50Cfy/EBmfjwiVX1OY
tTw+t9mBQJDXANAmNNvWVmcr4kIjreJSTX5Gof9zp+vpiRZBCeERteddf2tdpvIPZdvh4QdqESwi
CZyzsvhnACJditr9MjCFaiTP+jM1nOONhxkWNi/qNaBxBd+0ag7Gmh+4XN43QPwz5ywVRKkCZnTO
+xiSRk5r/sp/4nAWSWXfKKGDGyOoromv0gQlF20Avv5ypcWkNyfqRxO1rkpoHmDUTCrpJxZ6LSmK
nda3lfsFYPIc5zim3AnQEbWNRdNlTKkYCeklFfKmdZQrp80kB34z3hcyCr/m1DPrFjwXa4A51i9h
8XUhRT6wDxHhbbDBDJ+nUoZQc17CBxSCUoAZ6eYj+H3ikayIGknymi6PHQrNuGNFKssEGMfklQ8M
1rEgfP6U65WEeRuOdNpN0nSrlX9I41/jT6xJnrNlwmvcHDeFqsL5Lb5UYWa/mrehdfWE6wCaHYjd
79OV0sZpEP0ALV/D07HQzfdmxWqxckXCD+d5UZ6k0N6JGeX1YMBYn12m7PY/7azfa9M0GdF4ruZ8
lEiBkx/2HKpM6awO2N7Twggi+hNhKXYOKFgt7SlJFSY54cAL/GqoTG6Xjet+cGBI92fQq41TeL7r
e+RGsbxIBwnDIyaStYWkcblVE448sUaG+Z5b1MaO1J3j7u/4TmTYCZYekonjptwodQ1J1nbXdXiD
lW4Rc4DCw8QeWLWgswjNJlUxN/MGzLIQsV8pLOGrAnuHLpnb4nf+FmM6WM25ezFAjrFwqyEmk9CS
ecih4wZiWF0QA72GqGhHUDQCuBud/uyrTpkCiLvVBZNyIskYnJjBIhSlXmAK27OXHyR1L2YLbRxl
QcEQZKrNsLojzptZv3AFY37h12SENgYEJNIlEl3Pev70rdefT7rRJjGI4Hq09Kv/+MceKFBcLWct
vmHCyIxR8Jc7UPjKHtGTPqzcPa+nuOQpgEYVY2tlG6OY/kon/cxr+67lMGvnY2jnWLxx+08G9En4
tjAMWcD2RDP92eWE6bX2QcjUchxuCifdtLBuHTicOm+yUwixpO1ejUiAByP8lmTC0q1Q8Ko5h/IQ
VLc8qCmM8WcUa89Kuzu5t9bEUa16kpZG9mZWNYd+sHq8SiRAihpAf1zB6jiMUuknoe+GGJ43t5hm
CyAMvvGhWiIXyAyC/0jlu7Rb3IWlepaxCNvUYdM7q/bNj1qOHel8jWuWTbLBMlsogFBGI61ScUty
N+JT40mhC5EBPXTvicrITBwa+OqozlyEjilQt4fG/RzyoGqYVEQ4LRXFEoljX9nJlR+DKu8SKUJz
mwb3OoNWWyTFp6atbB9wcwjfjwrS8gpOtnsz+pGSi/lFRvGOAtIR0Pbl8EnMI95ApPifxXiapMaE
ou7aZW3vdiSQynkLDyIYJkShkaxm1ghb/odHtj6crXpJHLwHdfVqnoHThOonfIVCCRLHmhEbycRm
ZChvobfQQnBi/XQjPR5Zrx0qsMOG/VsTTIQHU090h9NrBYhmgi2er5Qvgoza4Aq04DHzPs2uKvXy
2oQPAoGF3VaZlGvDbNtxthRtZ7iLOC3MsZJ8k7qL50+HfShI/09LcPNioqn094bDwlLG3iW4DdX4
J9fO0tqEGHy/OgE9lkS4lfDuPtX3tiG2ThdmkSZZ1cWOpgvTzfFqq3pMYyfBvIZb5c4h21mISTdM
vim5e7xEsc4SG760DJzdUILhvce+OT+rQXbkdFRdXy90Hjwydzsjbv1DjNhHst9JqaR6NhVS3lJ2
Se+yypQeYIIy+n3FjXJHytA+XPMuGZxuQXbf8O12EZk7mgdce1O8f8CoMoWt89BQ93Qtg/fd2Wg6
cLoDEXpcyucJgUkRMoJBAKBjw3ajEl7SHB1u5vhtVvdPZv3dV4Tis4ziWnbFDbMyzSAuv9GucZme
057r/TceO/i/e+HOnmt6z6ucJ/Dk/9MbDsAyPkOaNtZKbWBhRdLbU1af2xIuw0zjwK/0iHVOXdCx
hwlSCCpmf0E6TMtx3vO7L9kpDP6CPvlDESvCCtoPEfXrX52w1fgBiSKOUACc56G7i04bGGIFW50Y
QfWflFArVQ+LOrh7eeLDHv0fs1f0vT+5OFNm194Q3nG9RS8nADyZG+8TGllWv8DRKOSpagZkYBLk
Or0PRJsZqPJLwpmE7l9gtqOgZLGVrlI+HZF2zWukY/lmqBIbf7Fz5HranwAg2rz9Ox6b0p8O9az7
b7XNebmnfogNSyPNbyFvwWwWs+VdHFXqXSDNzonYMNo/SPEE0GIdpg+slIJ6Sk2xXysBvybIWQHW
LuOtu3s6AT0LAlAcbnwaP5TIpQZe6tmtq27KX4V3w2dg7oRdNr5ue7F8bgjFXJaVQwqmJYXx9tgW
6rXh4hXNr6hvARamjEemW9Yd84P0IrRkJ9Fve77ukbC5GOpfBoNcP6NtKTd8pjA3fwde3PKqfHmb
XDOkJfDeyLlnwL8XN1ie1s3lUY3PxhVMBsTnhFiEggRMbWjtA2tIFqKo1BTA7o35yQ/SuDE2PXwS
e/5w5Zl1YFAnV5vS2HBVeORyR8ZuvYvipHAjOsKSrgfgMBLCNJ+m1AMbUPFMdPVbaOaqjS3dcxhK
oMcd2LXpLUXAvWMv6cQCeaB9/w0n7lPXNhGSyUsveTtfnAMC597Ilti78b/8K/A5c1mwNThpeOhb
M3CfOCUt5nJ7NAwnn/wftITWOFR/GPR+jHpaUQxiVnELRaO1WUEPUoV2Tw94z6R6iWP/3y5px506
dNgJVuT6/cJoYQMuo8laYZF5A/D6doS0QsuV0doSPYT6AmOBFp0GhqrfKTivl3KzoPVLPZ+3cfsz
iD6AoCsrMB7/QUWhyRT3GECa/2JFIC/b5d+mU/1r4QEYl4Gsedv1QmFMV6/AYysmc6+BDEruwWM9
vUb4+SsRX7JyEOfFROqPv8L7HTW6SOk5mc1zgnIIIXx+h/jL2PWp2LgY2ubV30JCi8ccDOu08Uok
xT58y3xUv1G5h1YhnBAADJ1YEAEUe3lmPGZ/p9lnokpLGyVoZ790oG+dQWKdCTu8f8BNzJMVbltG
qTHbmFModXt9S2+3SQqQdg1ZwlbRusK34eRPC6QGn2mWGfUmSquK1xqwtlP6b9zaH4AX10Mulcfz
u/fsrD9BhIOp5JWkwHn8uaJjTDrXvgh1PqmA+XhLvqoak6RVwnbQqAZMcuxj1jioX/bZFgSdKuZN
jLDx3KlgIV3iOhlcUCGTICg4cDgs0AwahGPD9RyR0JH5Mz0Lmrq9PMULPGmc+ZKDomtQKMyOV269
QkH9hneEud/97yGZchfrzfn8aqIZgaZdpnbcV4Z9QwLAIAP81I9X/uHx0zwdwVlTIDAAmbcSsrSb
CpHv23QS9MpMlKt/cVmxCdhWwQj4sZzgt8kxLB/jw0Xr4sb7fj5+FnGW4JV89XQeE2A5iXAWSshk
XSI30aEWrRGGnamwWtq4Blk9bSfvQ0eN/q0uPSoF8bk3/D+A080KHXNJexETTiaJKt07AN9wxAyz
poedBrLsdjWBlzsscY5IfK7dR3LA/2IqgKTZETZS4yCeULR9fQiH8xRTkKBnxHXDHjiMx5IoQgSY
Cxe5oSRYVvqJEAY0Ead1TTEkPuSKA+C1yU/yhy9cEjSYqnS8oFiNW4FfozZ8Nm0KEE4GUqJtIHw+
85YLeAJT1YfFuyTrxWAJMGSPrmETCFD+tJEWz33qbahly9hQtrziMsGz+9dMl8vUQAKg3h5AhrMT
u6oX21lG8DPYC2PuLtxM374/cKSAREUJYY3zVHX1MfnvMnoiYtkDc5U3Fn+tPmJijiDHfn59WfM5
PwH+5ZDdS9x9U54nvRgVAhTbeq/FhjeGjjThTnxKR198V5YcdWxpXba2ui6GAVDe/9VeWFMKgn+f
cBn2DjmEKlpcp01qEzRQhCG6NdTDif/elhsJSUh7mdhxAQTduq2K72zIvULjYW+PhSIEwdSuFteO
lcDy97Qud0Q0cokVrmOOpfWmCMMFUicUnFBI4pZDl39j5D5XN3dEL7BOk5WZ2LOLbj8ZXdDz6BmC
O5t60gwk7y0TLhOr2BjXB96QKWKQ9YyF1Y566KIJlg3SvGgij3/Kl993/gVfgwS+IijSbguig1mL
IN9OYw+qKl+MviKDoWutvQ/9XsnSkhrVcYQX7XTboq8Z3jv6ZxLDYGW0XkNq/HOi1jL+kKwSjTi0
VOX19Uk7clYyb3tWx5cqsx3GE7NAOvZDWEkma58jFr/+9yQem4EsM493qCj00mT6Pc/2beAFn0C3
VS41PWyQaAM//bMaokkaGiDiyTQSHVYP9tkvwg1hSVjpdSIj/jtlk/HUPuuUAFt99V4ZIwovyMHa
pcmEbjDCfwwn/vxcyEz0XtbTEqr/OsLpoBj5nElsZoWJ0DxQXES+cnGC7RQHKaTdSafYZdcDFpiP
lL4Zycl45agNhJDuh+zvLTXepapEdr3UwfBQYpHeyxCPWu4AgZEEFnOCcOzcXjA6sSlMFMfKwzqY
mW0cV4dK1d6TSWsHtMl0U0z3n1AOIQ8hrJSuUwp1bgjPkEY+j0ZKCQxSjBiSfgUVa/AAFYFMrNBd
ZXoG43zJLhrsRUzMPaTj1YB5PBjsQNshRkj5wLAWFLzCtXPzAhcdnOot+asDwpy6naUABbbS79nh
MYZl588nAPtsIT5yofga5UL3Qj2FITWa2qgYbxyWIxyAI6eZ7H4OxrnHLayn1cxw9I+771VFFV9r
TaV+BfB7m5WMsx52zmPw8b2eWmnkc5pNd/WLIruMkZUaJfa1yVQ//4uJGDT1RKcF4NxX37G1td3d
5bjY3Mo7oihk2l8UpHNdSU5vEzE4kZYmF7SJmYhhG+syW/YKVMOtZPSZmhWhE790YTayAgP1ANty
uayb0KhSo+qNTXnVpiDuZjI7PC51QcbpZZpQDRNwCQnmTsRb98dQl+vrv+bkWGg4C47OYyMbv0E5
Nf6V79fmkAru2xQvqTkwOnB9bi9XyhVO9Cek2dLiN9lNT8Dnyb/ctmSeh9w+rHKH2Aj9+zwEsMIe
TH4cQwl0JSBDVlV1BTW59Mx7yvNzxVDkVVrFJyMHdtigONEWGIIsOj9vKDOG17cBZVj7wzh0DYir
plx17V+tKK+KwhK6B234fBTnkPIa7Vzop8UjL4/+2Kj0jNPlU4aP6idAfKQn3h1md0oTN/zxDRmV
8g2D1iRyEnR/lzTb6sdRDVxQLaza+XX85frrRlU5jQ5acC85dDwIMiFQGBEEsJZxbh1sTS3vRamF
m7QCgevjnkdlWdq96OUfILkcjXOe3Ixp4579JjCRHTfmyaUMh2bjvGZ+UjrTaq0ZvahtWyUwYc33
sOOHe1ZnF7F68a2eZGV0oYPXpz98ujt3Rh7XA/t3Dtrx051bd5NHC1d/bJOTpev3D3lxOojbXy4j
MHl6kcNEV42NJUXKN06fs7fb4OJPkQnqgxszWCpmZ6A/7Vl/oqS2ARHLYNV81M7UWjPkpoBnWsoS
xiqKDxnbS6QnLyUYjt406230xodVPygo4Ld6PttzLZQkmjdnO7v5DEz26XERG0ywCQsHglat/K5A
1Ef5wIr52zpXwahuix+ihIaMHKt+YMC2wJr8EMEhhbDh+0Nlu/Y/iUGfAEVo8z+4xW4ByG091dWi
kGY1ni3Kj6x3TQUq6SVHd29It8koTCXFsMiDzKv9S97gy3zXnZIPW4XOL0oJI6dCecGdVtBk1CfC
ke/DKnwzPeJ4qoMSF6PedDBmI5gnH5dQfDb5wZCP5umEVuuvcq5u2UZ11KxTIIN54UCe146RQo64
I4aaIPGZSfIoKN6qcQvAXUjFpK1YVcJ+2cXAhNBbGVsVwWoveNITALrdu13Lw7vEZJeZSeGxvrq0
XVZbcR1veXzcekHYh1QFyPjfsZtKdZW8IHNcKd1fY0TXWKtzk6H98Zg/RhgUk8sR+CUCqbrVId67
MvXatYN1e7O5+voiKw3hFT/n5ZCNPzaRcNQ/eV2ckPndC0qnTIx8HT1U4675H6DybB6OrWyv7S0M
JElG0vcfrdrxPrVbkoEIqqDQVvv6HSVwjsWmQfO4avDjlp4iXsrF+y1n/wpJF3vkUvW9cVdY3dVD
QCOyG6P+DD1cP3jb/1CbP3SxOb1ls3tA3U8aMjCY2M3hoE3JixeGjsJKH7myuZ1vsu0upHcrCMw+
pS/6EOYCSf+kWk2QN1mQF/SXuxQboU2qdgjMicK7bbTWrjD/Y2sL00aJB0RPrbCLfgoffvTy6RP4
KqsDBifRJKWWu0zSi4Koses1ALPNZhSgEz0DAlELn2SzRhtd33qOFmMNR//juZX/d/N/+kVX8N26
FwvLHsB3AQQ4bS03qROzQ5hmxvpUxn5FMWaeEzUmGtZIaeuD2DW1qQmSMxggOgDappB2k7y46Q+E
qLxA+HCBvj/m8ismLlF6UGb0HIIuE6raC7roEefGuxbmJ1ptsTCkNvRPchmnjbnhqMP1cCBtQ3dp
acE0keeaPxej8CtHGesHJvoVUW4TUSgrQSyLvaDxNq1hkVy270ETUVsQkFs/ELG6X6DSPSZYk94b
197k78CB2uL7ee77M1KaluHYEM9XXUYSLIQFO8SbMniaCmwtKqGEhbm1aauZ6Qjd2qI92ThItESg
u7ksMJQXiPole9ofeN3CQVqmYPDpnFesj6xfogoMW3NtlOIg+P/iV3lvr3xLztwSGLQZPbzpvYnQ
YCKzXayYR7wsIOc4JEZGwMlfmn2oYosaXEwP96HOpsEFID3kzrDBeuclkLiFXpLG3MkQA+zkHGvY
cInaTL/VnCFkEppnXBenyWKBahiDN6Uwu11mpzmvPk8YhyaokfLVhfkeAVBKMCNVcV2EgUKrnbTo
O8kZ7AhT9jP6QPZXKevPNcTSzqk7BxHVneCJTwD+1FaldCePlcOCtMCuCgwgj2Dehc0elZuqp33Q
BUlPhvLGiXHI9WBX80r+9I1E4wuNLlEKDYxp2IE/kpXpMoqtFETdcn8FjMb2eKRQdeYCnJCsqn2H
vkjTUKU1O6oLVE1fcIELhBnubcS62le/S6DoyagbQVa15QrSvwFZPxfmSbctk5fHFnHUakMMlxbn
ib18Kpgozw41tPfDf0YKGh/l3aKwjTJYvP5REFyIJ7RpGgWW/QNEHi/TEujy+0uFtlVD5BHxXoY8
WCNEY1rNAA4Tsz3nifhwheJP2J8HTTnQQzMLTJYA4MSb+BIhjla+VwnvbpgEE0oZ/NlUVxMPAJeS
fqrjAPIKG42rjWelsrIL7KiNdxkfHfG8b6YzpN14ZFUiYhuh8k54f+jKdNUD9UHM3PLfvE78NSa3
l3ubvU6HkFo84uAOBXSzHDVUDxq4wUcJ/lu/+tGlRChwDNNdzcNUaExKv2KlwoXPpaGlP4sv+ojc
YGDB0lbMsM9l6XwcR0hxTArwahI+SLpf/bDjzEU22ZMvSaWTg5MM+XK5l7M5u60/cOMprdagudSY
4jWtI4Qtdg9QB47reNNfrheglYYYTu91xMxlinf6116Ov5htj2Y2VAPTkajmPD+6Lrq/9ByHy8TD
Pn+SfEl/4VFsXkdi32rCbXcrP6NgTab4vZbYKbbTWrrIj5WXfrhJ+0taVc76Vt+Ifv1KaGQxpaY1
QN9QSTMChXUTaktLtPijUrfkYc/7DD1I4mlIZG+2NQ5P5Mxzij/QxebzOtKEC2gYUTT1bRwCyoKi
9Cz7f2fHsrgZtQVsVKkG1mdvEb0xuglFYgG5bP8y7kWxZjL2izn0GdVz9qcxE1OLU4yQThZR6PYy
8cOR5b0sbHuAXpr5fSVM5YvmCzkzd1ZRdA365pYhGjNmJ2fdBmm0nCCq2WocEixgZUcIm5pKMWm/
kRYS1qK6gr92Z/AGoeju5W7eA1HfM5hRU2pLx+/EBNii5Q/Okf3Qry9Z03//yxiyJDLKBSS95hXq
5d1vW9XMRIoce/z/wSlquFEYKY8gvr1kkf/tG2FU2MCw84H5Z4zuzyKqU9f95uxKOyh3B1dsKuak
h6qbECF3hVwN0o/AlrE5TjmtLe/+HnI0qFdwyydGDmKtThPUZYnKffqMsqS/KhhgDnaQpvqverab
rPK72jS9gxOzehq9bVNkS+9mHwLx2Me9KdjqPmz5/FNVkb+VAf8f4O9oQvAkXPDh+GjeXwoai2y1
pEBpdaLz2Qw606adLuT7Yp8joDJ5ZAYkiYF7eCyiCY81svp1kOeuY1F4T1E+Sz7Tl0u+qOVMnyWM
YLhe8+KyIYBcx48Bo4HPc5ilJi0qHLzQ++gwsNRTig1LfitUmCQdfXrT83Id9zx4ULusDqIG4TBU
bVtHGnSgp7X/Qfr4A13b5UqeBAsLy7n8tbPrvx+5YOf9EKtva6zMpjuVawKPZCLTX1I/gYEmSqFk
bMhprjwYmpep1jlnsCT4iNnPoFhGt1RMaweTF5lt2+Y+LW01Fdbzu2h6/E8fbF8/4MDtv6isbuev
F0fTfNeOke93/lsNXHf3OqytZq8tSXn9nOQalh6tCvKrPPJTmqJtw/ugmNIuVGpnA1AmgpIQu+wr
sHwEZdGWK9BbH00nQgnltxaSqOBg4SHHdUEj9c6E9ZKq9LBPRIM1mWmiTJt7Q5YbnvmmkIXJGsHw
euCl4/5F1boBAOXc8lwwW7UHudi/y+tqKSGPaO3/Fn3ydiBp5SKm0mWeUIV0KUGTnIWx4kA2JL+I
AaTWOoG2tVFUws/J2DFXKW6OA+vrS7fpsHWSXJq11wy8sNrH6dAHp7wS/M9xq/Ke5081+lnWY4oY
1fxgUzrouiHc8XiIhoR8uwgJ7hJmVFT5dG5A2QCDfz1fZagj4qrpQxCezw+JXHqJyvZdb1nWdaFJ
t4EKvEgZp3jktvwfsWzzorxr8O5xhuNL8caxnQflDspceTN+XWVhu7J9L5lkmUBIvxUwvi1a6wCt
3+zNUyAYxcFvClIlPI1Hob+SsA7KDvRxJmTjeUsDjAS6lbZKpwcJwPgZFh1P4p+K7Mc4sgSH41E3
DFdvQIK0rcGss0PBDeV5xZs9k6/Y898HXlkWy8pL604X4rTRGGP3ZjRKhnWNAJ1ioRfxBDPtjOrC
R4SEDW5FmqhADIzdSN2q1dNubijHcjrXmJNnJnQT4YXE6kEKsdH757BuR9rEW24SyGgmJcFNHj5N
X03U2DcQNjxz2ePxDRQGP8goO9ANZ1nODsTHOmi7+mul6CTLq4hycXYchD2S2rz1YpOgKmWHFikt
E0mt5n0cPfVPWqJHXdLvaQmGe4LJBQjZIHRp3UnawdAMxOwAYOuKvHHsZx3QcG98W70eoZ5O7/Jd
WL/Ful7qXu4MIFwYSUWqTPxB7iMfFj1VLEeQpXokZcXqEU5I/p/nJ50FA76deuVX1EdRwvYK++M6
uz2JWYNRK1hqeKT8tNakDSgJrFwcXnurZnn42aoRQVJpR+W3wRbltczohj4DMi3r5jSsDlmh8BRT
H9CxFIz469awy8F8ldL08AW25uv7jfan5c24/Ja2zoHqJKi0Vf5amvACv4mu7rc0UxRNGemU1V++
HwSQj26L7qqCctDX9ePT5f9qI1VBMUCcHp3McOmVkP5MvFwWVYH5GwUftDll7l9eKBY8AdmjHzac
y5e2lYsLzeGleVyJOdtFctTzZiiy/sBLOv+Xkk3c7ibTRn8FVpm4e9/EpO7ducpfcE/aamiu9Mcv
+AWQF03lcajg6Eg4Y1l7/837xo4njT2gAaAYp7laRWlU7tTTaJEu7b1Qs2ZblPI9+0AzQc35LlUq
rpgcDaWrWF1EDfEkKa94CjAZWZWkDkGMCFuRZeShGe9FSbJNf1RszyK8+beqOlx8uCUaETdHdod6
GkX5YOjH2gk+pOVGknbq/XZfzMM0R41le0h4ZLmF1XSM2IU9pECHl8hpleFZrAUt04j5GZxQjqP/
2R3RJmzNfpuymtUGHYYUBh8hx+1DbUtKTALJqGc9uAioP+y63ufimUS5s8mQ67lmp6NSn2YsJq9N
/oep9bu09LJpa1xZyazXI86BjAIxFHJz76xpAWsN9SRLAhAk1FVvccwW6KmlCmlYDBBUppmEjt7S
L8XuvNBSy2G8WdSaXLOSO3Fl6cNYy7nR1X9OhDvEssCW2VmajdHt1VD4XIZNGA95vVc66K3+mSZW
5cPg4ly69nj1hyya5e9mDKP1dBMcuSv32uFyHtSXvAYbzBRF1S8+P3uniXDmwGhMAkYptfQE4VI/
3M78mU6egTqe0832SwigUZpDiofVV/YAwxM/yhfbAdHFkuoKC8prx7UBk7nEw7cirUEgsUcxXQQC
Ssshd0skl8WdcX/eZCb6Q9FUNj2A3O2nooL3AnabJsxSeDlqMnKYGoJet3NL32f4MjgBG5UmbQVr
9koCXdyOjHIqTAqZQ6H6sPLrWUwc45RnlGznT7rmH3wEB05TgfFD1WYx29dlQ98/o4FOzn8k03XR
utteADXdVbX9ob3HYKf+h0l1uWlrD3CMgK/f0X94O5VENJ0cF0ng7xa8w2gPoJHWRZYIoPDJJbPI
2+KB7X9eUGRW0zmPwLqk/YsKRYyOBZUoYlYIxI8307p9MMwRkOGw0QLuLI1f4LzOeybRDstTbnkc
nKXCOErqitHU6JpRrrEHNxh/VSRsBAWR7X/4CYgaaldSDb3yZGC4pn3sN7HvdGcEIVLqvLdwab6d
p06ofbtrPmZk/PAVLxNea9c4X7eTKHHptoIkp2foLSc8B1R27It37afjv+KGS9yNGxrRyvp11I7S
Lb2LkfEw3RvxPYXbfNxxddVZNBqwWLTDx2n/1dLtjxUAII1oit9d2R5yIx2Cr2UMKoV17w2uhELU
axNbE+s4fTL2LOwKp1PNlWR/nq9qKIL33gEzocnoZK31lpXOXlvju1e258fK1sMbHvdSw7WmL9NU
aFhA9S1hLYtInB+pwT5b1aWKDOLPPy920nOURQKPGIk24yoRKCPhkoTZySPy2vhR05DuuHISfYTi
DTGTD8sF6OhqKUw3O5qhqQa7Ohw0vtgUnvn12OH96oCvmQOB3xAcoN4ghrJyFSbSlEoGuM+Ielyb
/cqEJd6KuTTsrFYpvQuppV6W6M4VQyF2ydtCXOlaQw8wFQeB+arddL0gG75xTLPPPJzcNOOn+1JM
W5uiEQp9QeF8x6s4YEf30MMvF4zX5lD5O4yCxVNBVJ+1gV1i/Y4MPlzFJOGcoQFYyQ3xMZjdM+2+
FYfxKIggQ0z40QJLB9vOW4Ihf4eNB/T/Vq6tDRnJX9RYnHmHxauw54szs3OsZ8kZaK+d3VEwuuWJ
UVp+iq1XaN6pIQLvgztkY8oUUvR7teyc58i2q1Rw9qZRALq/qHQ+cKnh6tH5tGD1/aWaE00liCym
UhBCWR+HwduqVG+so+BqFMcvKtBMtFEetHEJw8Um/8BZ7cC+DdvlyaLm7+X7enGjutNflnso8Blh
xrwwtN9/pzpFOthT0rPXGsMDOTO3PrP+eycXUTQtj/jlS7Lcy4XaIEGIiq+QNwBrSpehBQeDQz7m
g8Wl3cCsD1dXTOpqn9tVXuiH8RhKbBJUlC0YuCw3mWmKV4kNPwunT+t9mxgeHTZEdT0nNEjIiNv4
cYGFIyCBQfYeUfVI0klYm6RYkDj/JMJ35CkSXQ2ogwSGPdaUU7ndRzUW9wN8oJws3QYCB7em+RYN
sBfJk/M4hrxLC8DWJ8BD9d4MOWXdQp7PRKMf6/6lkEzh0aUm7L8BjodVuRT/wDoi2vN+CO+fyqL6
R2TtoIA/zDgQaNAFhPCOnKq4k4ok/G3z8n77ognbOEyXaNyCD8d86Aa4yXYYcUEHIbIvyOSK3irt
vc1KPKIKrrMmY1Nra1oLvNTq55ujwzhZsVbmZrL7x+Mv3L7YcQR5qDtnJwVWKl7rUZseq8uuIfCm
BTOHk1iUhPGnY6bAkedIQGYJuOWs6tTkVR0+18i/Ed2ezNmwifwWQt0jXxsSlzrM9f8xVWOUI6dq
3MFrVtRT2Mqfz4swogSJAP1igzOrp5mrS8kNEKi+thQPPzgaIJlXOOzbHQ9AUQ4qrY4i8XuxSSWG
k3UkG3m96oZm7fpeHqGTlQuXtIrY+MkOpHzbEfwKF92v12yY6R03u7xwIf/pX9RQLlGUdJ2EsIfS
v1MPRHKejjFH5LwBy8j33cbcml0iO539DOTpdQET4VKEzuyYHTv0eRQ5Imjc5Bv0aH1UGTgSYeEx
e+HcIg76NiN3U3hlOkFrfe0DIOhb1VUKwfmHOwTKgIo2Oy11OWn3cMiNVuF/+qpGzMv0aw8ntzMx
xD5ANEYHZQ5VNeB6bH6GME6liZMd+81YY0vQQKZ4AcRy9iWWHJnes7Gh375AQ+fX7BgKgWKPKEXd
pKZs3O2WPPCpn8aHSQWZILWa3ceac0a2EDqZScnWSv8nBiaMuF/eAqfp0HXYYR6ioKxQ0iyPdZB0
/kNREH3+ww6Er09Ibw9SacQqrnAD70JlIjXz07dcC+ug0PC9oT5onVtR7U0eTh+++4vsmhAYJw/t
dsE48qrmG78KV51a9PYw2iOc1ctyrkrq3OZ0zG7uQ4g1Zvi6hMtB1qvphWl6VNvN5cJE9/pu5ZQU
Y12W0WWaikL85whf19hJBzUlu7u9J9BMYQDtgF81nMFwYAg2pDBPnK43ugPy6F8QWEy3r9rdF3U5
5C5DE1JWd+El8hFbBBn5Wl+I0HQeQ7MhAuI3SCZXnEx0uf5YujTX8zbp5VyJW8/n2Cd0RNbmK4xV
oYw424HRczzdoEzmckxZbHB4RBCRTbCVMbxWZD4DT7ddPXJ3RONVDUpYSoReRECbe0ldxEywYKyD
FkvyAUiwsZc6Xi9WWwRH0jMnYqTjVKGVL6Ko9VWrLSbWjW3MkONVcADL4LH55242KvKha+EPdLu5
Nh4WgEMYyoz9FCfPQbiByzH6zptovEsjapOGJfpjrMqD90ihZ65eJWM7XSmc2FK5QnUfyOd/KZjO
4rVvWL0QKtplosfs28PTSFb1oy6eBgC6gnMk3FoEB4z59RvU3dxg/Y41DfYLajsF9KwbjtFlJrXL
RnGll5dJuCQKufXo01YvQhAURTXYEKsOpJf9X4klpJ72OIJcq/ub0FPpZif2AM8zpx7u7LWXn5ft
F7FSDnYj/sSp6Qlew6DbL+Mu/ARo1/34Fp12lljAKtUUv3g4flMxTWP3JYroTPpHiHtIj6LYQs7c
CGwwmFfGrvsRLfwdOT+h0j1X7O+E6v4CKibsacNIGrYYle8Ki4bRS4lLdSF29ZYs4TnEnG6tWF5s
9W9Wa71TEI8brpd0gEKd/Y3UHHObQnKlJP3qiTs0tCpbQKgtQJhJbweEXtzzR+Z6U4BX8GJtQiIP
D+8XP7mjp9YIDXvycjlL5zyJo0PHCesl2W04QcSh3oYwolTzAdQy4iA5P8oIb90Vd+CEBlpzLigE
JiBw9CGTOZWOgH2uJJod2ifNQVJdsDtO/kGAIcwbkpLDNea0GjIsDSObSb3HeKmDDTm/q2oBV+PZ
dIwrWXzmUmpB0kOZY25s/VRile33KtVX8VFOOPxQ0F9kDHDVYASjbMwPHEvDclgiUVBwxJ1AlRE5
xjnLnxkYR61tq8prWzN+TCl8fWYghtg/pBNN3AuDK0QoKlS7uk6w+d47oORzyN0vqFG23uPlWo2S
uxdHE61MOLsxR2x9cG33hCS/eItGD4SWke/J6E2g9rAZOowX2NoFVRnGbMnuwRM7cNacOdDaI+mh
HaDXgX3w+jlHQIfVJE4amf/cbpkTYY8BqwwDxb/xkeouJqOA/0OvzPJM9QxMGI+czVrL7UCeqRYn
ox8X9csFklbj71opSJRy+bObFcFampmqorV/eT79wO1TVi/oYs4/puiS6lvf+Nt3u/9lLH4W8Wpp
uPOLQTjgJer3kgoXoXU2VU7Z+hxwbGqCF//JgHjZ0YGsAEK7XIzVGZlNnXfLO2/BNTkoCcZAb/UX
nqW3E0u1+Fc74lJ+HCJiabKOc4xq70Z29hOUQiHjnlys1hqPNoDAt4FKr8SDWjIRkW5+J2VGqYmV
+pRqr3veXy4tjbS2Tx7yec1+IHp7r+QIEZynSkS0Gk8x+Kelf9MlpaT9d5ib4lPWLblQnnXQJLp/
2t3c8U9GBpgWI/uPmf6IrE1Cd5dV1ACjXyIZkIz0qjSBbihkZ+5t3lZQV5IssGrAZ4W9OhS+G39a
eMs0pEtRpgQQ4+ZwxHTK6iWZoC7sDE4jGTWftxQM8Oy2SkQU2loLi+nf3+k4ZD2Ba+akKim/7c0w
cyJEYWwr8UTtfjVrEm0S/gDEdWgztZYOBEluvcnCyBUb1m3n3LJMxYxXjEw5pCFIGNgRK7H/ttYT
3/cR4rNYpGViv5SW1ifTrbjfSWJgDDteOlpAGYRa8OMo7CYaztPrQSRnNNASa3QlXDvnPLCv9kSA
7uQORbXnNXMTh6+EjAyN1TIPTDrKzmuf59eQ6ToV60FZGOLjXGNw1bpvJ9GZzE7cXfp4qp49cWMq
j8P88WykzhyyLRtbOPkLTXVR3Tx3QYM9xGpaQlGB6k/JTbNLwzRgaupvQuCfOYP6mAtBAAhg6eXM
mGx2hoDlNWjWCDQdf9fY0gJTqFDX7PAUi6j4tVPDqeS+ct8zGLZw1NY/ZiBwEW5/8ynwL/aqqmMh
UbCW6Y2+9evq+BaEAg4Zto5ivMvAMRcmwVv/oAt2th7/ppuCqVKPyPOYEyIDYV512NmUlFAhwXYO
mjf9zeB/UTDa0n8J/ecnZozCaqVrEhYK7Z+x4EhUdbgrh6KerYuDvwoucbelJrhMDaZ8dTpQBQnq
pFRSMZPDo5HV27urFVXc7vJD25qxKRPiXWLr7364FgUY9Uebqe4MjTtFMZlcDa7zKcVUbKR6mK8D
5d6SnZrHaGCto5vJY7Mlh40+Kg0pMLTUFgacqkYP8yLWKzIJ74icOXEPFLc1rdfZywkSrr9/R8FA
tQL9MY/m3GfOr7nJJQVovnhgSs45e9zoFyLdc4LcGWoqL9/9gNa3epWudUD4up10uM8p3yicfAkZ
DdrTFxhSy5lo1KRIJvYA5KERUUT83U0rxVxFP/ZHFktkPaF85dLKZOspGvzlzn/k9R/dQc8kLeGb
xL0SGOyv69fg87obDHTvgSGEt1QaF/rJedRGJtBUCSX7hq4cIZ+FxMqqOOh7adl3Mq3RyONYnAgM
zjAhJc6b63srwo5/JK80IdK/WSOZtKqtRuregee6ViqB08nZgSfXwY+be2TN2KpYFsRmpiegSfEO
YjMcWxjeoM0NUwONoK7MiIlde3q0EWMo5h6TDNBSaoCREXegCGF5nMR2ZMHfCbq0lxWJLTujQWIJ
G3QjvwAFgZhNrf7OxqSZhkaiOJ4a+0u3PvQY7nQXaWnYs9LVMOWObK0iPRhNF+LP5NnT/GVOJAu3
F5GAbvvzD2h4DgFg0HiHNn/hJ3IOvv4jI7jXsrGaKpGH76VJRTeVKjvA1TUR/eOISwgEuHtFlqFv
uI3VIlxhvBc+bAq9X9ZzVIp3RyczDDOaEAXG+4B1hbBqbLPvZ8RJwQSeJP1/jwceAVzRsuvHsQZw
uiZgzVlU+T3sEuvP0au9Ou++6Ol4O/R6l6atoTTBIW89uT1c1yjbVzPOatmhkN0z92d+84CS2pg7
zfqlPL0WJcebM7TetB5ZDyFVIu5c4H6Z3j/bCu7gEe10POsJFhOfYKboZP0QIQ8bSPSrzTPalzoH
Hg8kozZAfbLwKN4e4W7k1TAmBQh8iXf/3CcruYCMhxQDVWh8F2tEF7A2JcgrINrZ1Ykap5RO3T7P
RKNDNn/sabQH/M5Ltu7bAGierKBDCZX+yW0cQOskltylE8W/CwX/jZxyanQDhNBPKwlhQ8crSJ0q
kGEcl55AZ0c2NNikMxo0TQzZpxidtShmDTAJb8YLZTZTpS7To4KVyLPAxlgYXAmyFw9RDdEgphHX
RbzHldZFr8wf9gi1N9JuOmF50N8kJsL4JH5pbmgZUeYaJPcjf3LlOjTQe6z9BY7AX+1D6Kdwcaqq
BQrnKSBacNSkduVnBzjen3BJTBMrkUP4DHrls8so8AUG4G+jvyI2PwtVc79TpFx/Wp7iTWatgzd0
5jogVOUJwiYEoU6ZrahEXYbdfOUBhckx8autUlwa0dziGsyzZCliJchesnV4tF5R8A11oI4mo7AS
HpjN26sSIR+0mmrXoKhJuJwDDDJa+qHYsTOwjm75KL4t8WO4+k46GVv4FakbRTALOYNLYg1/PWrN
HHgTwVRmcgWz41v9q2uH4zyZstJEBdcUvIFw4OFKPizy8mD/+6aNORqDQSy0dfoeeeOWGB4wtBDG
0sQ5a86pczhCBr24d/JHximN4d8EZLmSEAvcbx4fEKUMliaGchkBhGIBp3qSE1Ld9cqn6LY/Hsos
RB3k67BdskOnFiBFjc8PfjUpSw9MKIc5bkkpiFPZXI7Q37++qZOnG28eu3fHf7d3CdYJDj1qrcnd
vc9BoJC5ZJ98DU5w5o6F0iQyaFvuMFZbzXiHowAqVtvYGMYYuln5tcE/+DuFs9S95cE1JTEM08ra
J+Es1oD/zRPvu36JN8aYksYKDKRa9hIfZF07oKMPxiGyNgbtIChfHIhX7g5zVVJohpfkP4rrAYzQ
0nxsjx52z3vCdp0oRnPxgrR/diAYdOUifhAcZID+Lheiqk8trM+8Dwo6Df+SFLhR5S/KMSFTjtgF
or/SbEp89Db4DREeFzHVkv4opUwe/OowxS0QIjSB8gVxP6nVbNPT+0dBlycsN6Uk6qdrhH8NabMl
DfJYSs+jfxHacbCaejLz41KswXDVqRY6LRWJDOq6wKwHCo7t1Z8vQDdyidu/DyxeeE7vdT8w2nvJ
pr3vc0teuS9QsRoEmWrAHsJwvvWxU+dXZ7iiJms2rSVSLSLHIavfV4HT2IQ3YyJPSTmhprVnq2lN
73QM2P85Kiu+RbDaMzJe0F3/AtyHhfRoBY04wqCxuK+on7S6JREXfnQoAs6yraHK7rEJgWqVpV8/
okCNAujnVupg5kTGSa3fEJ3KzZ9i09KAVVZNz0Ezvh+esZqYdKP2jSnB++uWPwaRBlLGke9vm/h5
uoksgz+mzxulslddCq1hh2uSAFWvbCfds688XfMqqEjssa1yN/fvqGCQ1gtN0Uw+jnEEECTho91y
rkEAQao4Qfll5SSiqMmH0P4FcyVQ9AM4vjj3/ljJv8bGeRWeZ8571RT1807WDHLu93pFFa/1jfEt
OGSsbOnW1U9OCHXcGw3x04jcG+fmLOuKXC71P3epzY25Co1g+A+zSo+cWiYDlYtrzLBuHqwvzVZ2
D+bj5oRXBdDcZZNnHDNB4z5tHjmaC0vyEFmLOcPB7iSr8Pi6FA30Kgj13/VdnaRgq+3hJScwIk/X
LYdkFiTgXOjIZOeh53yyavy7c/gO/hWbWrzbpNAC5i9g9wZu7YQTVMQIkqFTUYRUPSZxXuZEOPCA
nJYOVUKtpgI/9SwYRuCV71WoxynR9uwaQ0woqG6X501VGnVX+ymQywdN/YLx1qbJmqgVCd/GjMX9
LgfRvZAEW/KB3ILZ2isjqv3jgksReIhSpSiJVd1/koltTrDvT3o/FVHC0aRhDcvNvK7IgnNP5Fdz
TrLXBfx/IjfDW7/gZaUUVz9OJdsp3RZa9abr87HQpFq5kBQ5w/hM9L1D60cJq9InfDZNVCVUceYm
AA23IPQ3TWAo3AOpUcedGcy+628d70UmPVRNlzUhx3ZLZCnLGsSYgWmDNFMB961AMcXD00Zbx6Ak
jFARERo6IE2zDS7Y/wfcSdhz37EWQYqxWhCRbnBVjPgqZSXw3di0oBMJbKStvbO4VPFjESpVJo4m
q8BLZXtLR/4tPjGkX2WesEKk+63ao7mFO9Vnm5Ebp9PhgfAsOxaXAAOrpeIEU/ba9D3rPXf24uqc
sKz7BUIBuTaZYJ5Gk1zDzk15JrL4tSOrjH9N6hka6Z/oFnGEdiFVJ7eHgAJsRJJimrJcru0Tt4ic
HFWl2gDnsuAYm/2W6ebDK3IgHvh/Nuk2AiyP/Pd/oSsNeRkJNrtLTDEMuZfWJxREMlk2ZPv7qMLZ
XHaa4eEXkm+BMxn60H5eCJRiMQlwCKpPSUAdikZQJzOv9g82j6qvCv4K1aMPU4NSOQc+Rocfm5T9
O986KF/VIQ+tXRqqRhBXzJoogf4lySDZy3JacLo5jW9G9tLvnrMMouiirMhBnZioqd8cdgFiBpZD
q79TYqiAfVpCMqs+RsHcsHOcijaR875W8xSN7ptBdZ4qbgSzv+MURBf/rnHH5FlrUGus5eJbGOmT
7iEHXub4szu4miMR5cfGRfUTtbna46ffyd4GcioJg3L6F2Dlw3o7LpOGKO+Q9DCtqOs+I5TBnf95
7jrWKQlJkwjcWaSiwiYAqENmkd6SBoys+D1oUitaKT0XOTp6gPWKXKuPG3btpUxNGr87cwdNSddP
ah8sy5RT9xBQVdPEio7P9X6GDH01C1LTvqKvka9tqGTyHyNTdS3hHTPxn4VkzlXd1EjEBn2GmZ7J
KwUAnknDgucLVedru3UtNGnFBbsWMgbPrEyNGyZDLIp98Cz/eDSpwYoMcWF1sVZB3ysZ6+/RuAK+
3J9VGZDnNZjq4d67PR7prIQBB3VTs9Wt9kF9QEAzITfFJ9i6ueJPDM4shaspAfeZT6grBH8qNUmp
SSXW0CosYpI8Z+p6UMWY+Eu3TXapxhIDAGJCT5bMgSW6rVGIBBZADmsZs/iDZcgrdyRf9g7pujTj
SDrUvEXPjxIRH5BMGCiBZ5s+zy9CqvrsZhCXqJKWXZTsygsi1b9MpODkRPYg53apJivugNFqkoWk
VpBZzxjJ0ifwwGSKsN8TvoSSRQbHodzlo6/PpdUy552Vx/gUPVhfHxZQLlGQX/9Wtu5x/ALvWvhm
an5Xj3hfAHnEygZtDLIPfOO0WLkEPG24dVN9OPoDu7K2h/KVFxmhQkGRXKNhq3V70jlj6TYn+1Vo
0lgKg8O8fc8BSdjiBoHwpYO4iTFgE0YhmGmCKo10r65e+WG/TyKPD/pWwXni0fw+gDkN4ohOohvZ
609BRUm/8xT5Uc4RU+81JDaHAjBK0q1MUUbSW3JasvrLsVzp1n0oIGKHHERADxNFhWHHwC9TJSmg
fJ9fytowyMhJeFYrpw71rxkP4jgypBUoNUfbYASgdiUGdT7EjNYEj6avUAfmEm72GIC6HtfWerOK
KN2eMO2Qj9KpeyRcqJvYMa3tC89eOPXM2D+ls8WqP4GyMpfthgtDAJps4KHs1i6vcCzH2rM8RjZv
1M+yQrZ7bE31RNdU76eZ72MmqnkpSEAs9UzKFr2OtvEvuU7wj5U4c4pwWM1lPlyCZTrGOwZ2uCJR
hiTJ71/38KFVxNWmIo6ZT37BFu+JPAZ0AcXAEYe4V/SYwGmPiY1ZcLTPxifKQxCiaUJmbLUddmou
zy9lHkpa8JA/Cof5U+I9feWy9jJJ1iVFFmZtrHFSuloFnFaf1ChApczkDMLcozZCALyaknNnJiiG
lNg0b7IbaFg36MUoopA2LYnr6NvmNsCKd8dbFhW1RELPXc95EOOeea//WoBsuy4/b8u5CU95lwUC
AvYUY3gNi2E7EcTMrRmVagYz2xSmgDzp4oRTHAw+viw72FnYLx5T3WM+nIvI+1zFbA0sTc9SnYVU
/GHPbXfvefurOxtpNBEFutYHo6tmgv75qBASYvfOL6StnzZrlizU460LKzEssCvSRNutQITs51xa
0RQS/PHmNnnmTPTP4g/V1E4rLRlUp8PZ2kYte/mlLw0sQL3kknICqDbwFXltHSxNSyY9mn6YSTHr
wNjuKASh+dZQhUtS0cGGoK20bdLM+7g33KdIcAOvFeT+BaRYNs2I3Lx0UCxIDxufLZjlS3CAwYjX
giqStAmSkpjOgE5DPpgfyXnRnuEnOJwZXFloventzlNbzO9j+YAmvmYYUTLFaniisU7e4x06lG63
NPtX2ptP5iFjMKwoGEMK85LGH5f7UkcQBQapW+D4QkrTtM2ApD7idGY2ZGo256rspA9X3tK9kdm2
K5JFzy2dR5FRkLMsdIDlowEHnjYMnTSjYKiJL3bq247yPqQvCzu21ObV0K2UdE3quCClbJMTATTU
5XQhGB8kI49okfX0/swjUt7njBhjBdc/8KAhxclY5xP+yhxjTyIy+tKNOyzYHJdjy/TP3hKI43Zg
B7GShY9Js1sKiYzhmqhtKu9CPeUxFgVahhhAnqPtYnpdZW56Puz0tlfSaWpc0VgrPxCGSXpMoHYS
09PvfvGsy67waCZQWr0pwDQ7QM/8zjYuHBGW9Ia1jhtmcoTRJXn034PDJTtA/k46sJhLWgzuMFQH
1dURkmbFB2QD/odfPRhR2G+d1FTbTUZ1fNIAi1HWqh2/sGB3avksDIYcoYfn6tI9M8dadZeARtku
Kf9RyZBlhp2PxRJF5dvftVDrUZIofKUV6OmmhGSQh+bYWI1cc6HpoWdexCKrkA3wjSlGUPvRkuBi
AjD4z/SeOqrRIYyT99q0gXm9T94XgnDpDYJ2X7YXVst7XOC5okMfh6f/ktEoF0BIA2J7FRzPh/Of
TIW9ZfitK7/iJPz3Ah84yzcURBiYjXoWUcleV75TBGvL1/zRueZ+adPyibCjYIHfcPAb4zgIQdMC
aN7aeXu+hhGhQk65esa8Y1y6tR9ouPaDcyXAc4WD6JjlELkvUFZNWlgaMlxizE6YhKoNHJjiQUFT
ETx3S+iaWDoXRz0BZm+bRTKG71niRjdmYONt/dj68bMWO74H1tTSFGMkEi5jI2uuSTwVHU2zpSxf
1moE1W9m7/CvE7onSIxY6OMdwEg4H2+BJkkSLbFYgYL0l2wt1eT9TRxy+iqViq/7mcPCjmROb1kh
AExyUBy1j1x7+f7NKZPlZjYR8YBTVApaAmZ5tYIlKRolxBt54rW4+LlYMOC01awQP2mCPa8JCCom
/kqHzj4SkHKeELnDPG6mzGE7HA+AUKWRQ36NHt5JTTC+0Q9O3vQ6XCxWqX2O+1hlJhX/f6074FQ1
Nr19ipwsUNV/+Q828pnOVsUd/rqYzOgQcRRRf1Jl8wl0cFDvKceMbSdWUeExXdY9OV1wpbCDQGwa
XR1HcggwTrzqEo403BCsklP/68XSTlavk1aqm9GRVYw9fAdbaHZbyg3oA87ixvcYyOZcj6DjNVQG
UmBMr5Zx47aTI7NCn2E9OUY90D70PJ0M/amKqaPtrsxs+P0iuyv5yVmkMPQr9t4E1YiFHLq0F6u6
W0pY9rvathS+qbQTHh7Gg7p7f6fr08XGEJaWbaiK82WwQoZlsuNhGX2AWMv7lXZRUZrJyaLQnkYa
w3UQvAPvwFxxpjQfdSza+odZdNtWYJ1pcO2oAVur8E65HCv5tXxGXJUbtEIeAGqB+y7R9vO0vA70
7z6wCnaigBPO7PAwDbMJTBtjOHbrNzsPEg7j+orB9dEqeNNSJM92+vNo0dqsBn7EhxhpuDQVKXyO
6Py8AUtd1gkywDtm+PmBUvow2rIuMGN+cmM805K/yIO8G7bkoKQLUmIo03CwRm3k6jftm7kgEfLF
9Fa6OlK+ulZJk6XP7ESGri/8xz9IZKrcRku9T9S7Fj6/8rwH7QnO/oE5h4c4YKEtt1fCAsmj368p
zziwhNYr5N7+P4SMjEfPA9uuQEDSIJJtihyWtUnDweZk4Zh0vK7L8AiZ17YELN39ki8nMHel+oko
tNc6GKOgaHIfLLIq101ijP/LCPuXsZH5pZnCIPCRjmvCO/R5WgODFhjfSD1GUzp1IlpU5Dx84OZC
pSqUhUtfytQYCch/yXniiKEYoLNMfixBwf5Qjs4orWZp1H6vrRihv66XP3t0JyviA8z2cIeGUrxn
1F7wbTL7ocULptn56yzcgWMW6OBnP4K1qbtxuSsSWymPYi+7X+feQk4ZjyK8HZMOHAitgHRz0ERA
DHJBSdYZg3YCVVZt0ZBqxwEbEFTrJSMSA9r5YeKgLTZocgp7mZL8V06dTSpt4kAc8YlHBdHZtLlC
O3Po/JBZUW7O3kSLiMqIqpQShQZVsItRT/2sZfwYmJ53R5vJUiYtbV4G9WRb+tYxKxrMwVaYLPzm
A+Bgg3Vdqr2rJyDDPjTFFYFDMod2G5gTXSQTsx9UCIE09HfE7/KuJbwR4aQajhSJCOJDmQbrkTyl
nfY85o12ZSF1xsjOa0aAFqMneoXaepdMik36WoN6UA2QyPHQH3l8Agt82we26GK4q7XaHPN7k4fX
oNIVRiybkL/yDia61QsZ10RZYBbc7udw2EbufUnpop6Nl/nlNsRF3RHCh/w3dBBza+QzwwHdnj4D
Wu0Xk8gmCc4h4U+EM+pix4hoXJVS9qvwDpUwW9q+OYumqJEK5UFoq69fva7KAens/d0GljBt8ab0
NBaz0mKFTqDKH6rRLim+TVGvONCvgbr8hEhfbh9G9gZRI/lXM5VT2LA7+YSxtblApYI8QM6xTNcU
/9UDJW3NjoC/CJbPSKOSXgrVBbsk2zr4XxMhkzE+KJsuPLslAjA8rZTRi8D26kO9HznT3/ZP04jG
5PW3D6FM5E9X80Bcuzy+ayH664IFlTXguPzB6Dswa+ScaaVicxTldb6qnRdszzX0lqTk0j5AEW6Z
QQqhTdmUzan2NaTqVhM1b1FMZAEOBIr26qtdOKAlqr/SVEeJJmtom2gCx9SJ8ZBY+UaIK0eG0oKR
3H6z87rcBQi4D+21E/IuQLxLNxdwfd9DVkoA0/MI7EUmKXSVXSp9my66j6Os14N9ClEQ9myafuNC
4VGjfBpY1OQ214IIsdbA8QN4bhK+xnD2kmtkbs+CsHMat6WvjRNpcSA1gVkHcIHW3PdSZGvbJM2R
eSMZHkRN1l2Z+ePchOAnzkAR3TsUFd3WS5hnNP/e99XYKJfsVTKjnAXtNWlNOGT9GR6KJms7j635
n+xPTowPKVipPrNsg38Xy+IMwC4W2GnA3o8N9Js4+5UoAJPsRwZnwTXLQqxTV6YP9lYB1+WyIC1f
QgMwyVwXhkLf//GqqlMWaTyN/JfMjdKV7HZIYRztoYad/0JN3LhgtRGPddtvRlrj4q0278zg2GGx
5d7GJsk7aPbz2v47d0ByAlGHfOWKHuLt6dXIryTVL1qdU7ZXUMw5KqfTkrZCC5DGWuk9VaY/ptki
IvaPo+HI5JQfmtToH4RInGzS6Cyfzj/3GH4cKAjRsm7QleO8ETPE0+3b1KVWAqGsll3v7TBrL29n
Vt+4cLDhIvVhVXrZb3YjfqV5POMTlS+7TBmwkDik/uF/cHHS4aKJPaWeyjFVEsVvQfHmaSEwAt3D
rIJS9S7DV5aMX4nwsKDVuPU/742MMgdXzDNF8L3Yz2tEFF46fsbbarE7wHkXir9oFbJDPNLJer/g
AbdOn3wPUJagJOlFY43iBE1UuXQp14fNpj6c7nlOwd6X/Dv4nhmXnSMkmRSfloUAFLZxFsUJ85Ab
IglH757e1dcyJnQnqZvgesFgEqdKz5Q4yB6pXAq+31TDsINi3WWCDH0yIWdtVLJIy7uNpEt+OTr7
Axbw97M3riKyDuyhQ/X1rw11yPMxXTndIfXzy2GgfB+1lMAv7sN4FiHFiEbmcTmGy7IOcFSszAmj
azqwhmTdx6l5x6cH1Z2Gc9TeyEtC7vcxDjbgzvds8UfHc86N0I+C4nKZLbV1XzUbUU/xvh84JMSw
uIMZykCXKRd9D92zw4u5BsxWBL0PGhWkuRLI7yRINXoVsN7G04Ptg4V9dcbyr5zSIaJ//dqqML9g
iVMpy8oGUJsvngedKeZ7hrL4ndUltxqcaOdSzCnnxWSxIVcmCjtPAon+EvA7Thvhet6DVgkLq8t8
g99svKjEiwO5fbdko33wWWnbFELb+so/yV4j6jsRBanU3IF+Vlej5g0xVCZ3DuWBF5sw2vVOxA1J
7Kx1jwl20zHU/iuyRTmJ7ZpF5b8DujNByNZuWDlJX9ZtqKWCRha9X+orhdMUc6+j/VacpgA7uxJH
g3l1R8PCQd020wfBm7KCBwLE5f9uh5uWguSaV8vmoAfR9reg9m3fFclm1kGqOgHEd8vxR2fMnFay
ANOY90aWLgP8T3yldnu61Lr/1q+Ap85bMor1mdZKzPCMuXokPAf4k+TUZ1e0QxduKr18vBWsSBNg
VEm7L5KRuqSmtwxtF6UQzI3hTXkiGjUHTw+zhA3fn3hwNRdKeIjPWv1x8hQWGv82MCBVBPwbkTvJ
qx4k4swWH7r4L9EH3xNDB1Lp/RSKqOneaT4VkJQ6z0Zm4kH3+JGY7l9egDoFtw6LR5i+C2ebw8qO
A1mvjyXieCPE8Vp19W76zBfm/NtOA7ZqV+TB2bNHNt6RolBTnxQMv7vnQWkUjjuwyQlf/Zs4yhWd
wWvFVs+iivkHX2MuBuk/sfYKXfd5VC+ZxLYR7iR9YvuVkjFIHMyunMiuQk32Z3nr3VgGdrLop7C6
ozC65P2trhOxp5Iu7k3ZFdJ6Y3NkN5/1CoSBW9NdBDnqgQga4EO6BOzkPk0AKo42nyM8+SayIjCi
/oBH8UMd2h+DSqk/VUerABTOhTgd/bhx2xR5OtHbHtzvGLCG/tHeI4jKHkImjn0/o29PPbfDJVSW
yMON+t48/8KrQmmKAsnW6lpkb8DboLLA+sDH0eWGrmNzZfkVCZkL5GDjHdu45I8Acww2fZHs/8vm
XhIb0lOihsU3KMxOSrublD3prTU6XeGKcgNvtFwBvIlCELuXMFCkh7inGI/FhZCjeqbeb7835Sy0
F2dUtb97LTGak34po8XJ8f2xjBwYWr4/I6nQoiY4BNh2YOV1b3EGR1t/0dDOqcE1r0VWHfJ2j3b5
uUeGwVKiwMLIY8ZTcfyxG1eIGXfO9jGm7OJejTMkHG+m73f2YJmhP2xh4lEGrYQLikYTYmPHsl+e
2Oq+3LRwimM3ZFKqQ7cAeEw5653/+bTMhDMIKbdkaaQi//RHr75EBJN7vSQi3froC4s/eTykUQSg
Q7asRAMDGRJyR45pI917NnLekCYfY0EohB1xowylsHJuTPt0MrHirWZdOeO/bhtcX9ZSPrFFzgqv
hlVPxEg13JFqfZ8gww20oho7FNV7W8hzBicgggx4AU2uKpOmMQ8EwCNgaI74bCqN2NmR7+yKhypA
Z/Z6+J3Os2elDFpLCHegyoDAEwvRass4EM+lG+LzeeoLzalfj40odCCQ5cMb4s8vJYPsTv4so3Ay
PFgAwLj+5WUwAEiR3f5+Fnk89CF3xCsE8Of9k5IrpISOoKccFaPUoGba6+7RqYYUjDQDNAFvRgd1
QAEeSZzYWiIT6JOlFowmXguLCpCsY0QY10XPAMuUtOVpc/rK5V4mOvsQJcS50E3dKGWuLgS7i+xa
2wrbvE/HmG6OxpMcglJyW5ShgxGKyEDeSs6OPz2PynY93cYtK8MK0gT0e5tl0CzuAAVX7W+oxp2L
J8+QD88L/68kB8cCQjYNgdvzQurTe6Haqwln9pAp3sP6Aar9wDIb1sg7aCBibztSIzHhuORBcg69
otIXX1h2gXTDlxxZWvIMd0le8r4sR7jyM9Lu9v8dLpZMXCCCG9XnvlFBWezEWzwSwJwBjoGGsZ8g
7lAquV+NKq/grCpl1BuAK7c9sB2fjzT2MZBVf5dc/0Ejc8aFR3C2lYhjocsjeJwJSRLYYg0YgCCh
c907J6K9T375SpE0A2usdcEAv5Y7aaC3GLALv3xKHnLf20yRKnLSYF67pzvtcnTgj+6e/6tF6afk
Jt3qRzYenRXqPjsm9PBD0aC28ODejcoSgm7+ZvZJnkhRsGv6XAk9amuxTuTJ91mZldFrx7QsSOhH
3yXHr7Zw7jet0SOSRRc/YEBOGwZOqFbrdeShFGkeJsQdh6n3wN29SX4K5aGbdfdshhXjNE0lfPCO
WN30kXnInXp1gjJ4KBCBj15jkoxM9qqLo4BOwz571famIksRQvRwUGO5yx/zI+GX3uzecaocZ493
CGwLVa/fw6gDGGb6IJbGPcRxgbvS9CNUiHNCx161PoOlR3mf3EpT8fxaLtjC0VZEH+SS2LykuUlb
2s95mQ27lS/sYzegJV387jzMyHPkbB9ql8aihwPhoKnD2Lgc+MKDAGrUxgU1P4JYD3/zHuHUnVhj
loYMn7DdkYTgpxRGdNJUQHz+FZgvD4UVOV/sNnxZTdivwOnCv2T3tA8QIEVMcR8TL4LMzv4o1MZI
QYKYzWkh6UqIwb5p/2MLzVQLnIR9SfRi+ndWo74M/lWh5yDGAWik5dzi0Y/1dLHMJxjvaEVTkVDM
x+SxlGSAAQfxQtgk94Jj86nrSVMpuw39LejE7FV/k02MGRU3n0OVq64+C1s8CWIlYbfLuSX43NKY
O+7aGE0cwIzCN/RLC51z43r89lzszD5Yk9LM7XRnr0ThVv2nuz7/gSoW7mZiSdJo0TWCOO+WBB8P
Flli7v58UymvT6qQG55C643V4tjh2s5zRuXDVPJyyd/M479QlZH3w+MTZ9XwYxWbFW+NC6KN1QaV
YFuyGwwfE/PnYVkYGEg8AWbKu6j7Az5lcr0fMUqPJqWYqiXgUhJbhoLg0SVjMY9MrL7sKEXeySuh
26eNOvm1rtYAZe2YwVowVqsLeUqaVd5rVOx+j2sOwC9BRUjp2ufv02YMMc1+8RIO/qOM/9//O9hl
cHUCnjkf/LmwPb7zRq96IyJZNU4wram+8gmwZEUFjVEEMQtO9TLVKRWVEBzJ2lUF/dUYeu6MRdjb
otUYQ8vjCPwOju1ZR4a1/j99+bJV/LNoY2pF560TDR3jrvXCqkZUrIOmDPZVKqq5I2FAQlNtNqSw
idsnMo1tMjQU6KAM1EQEKjoc7uYx7GTpNwC/Zq0XuuIoK2xpkyFlBU4VDY7gM9A+CrKlmChY/gii
ZDRuKeuNzBkYPUbQ01MCCClu71qKTAC4uZctEgxsyudOFHDWuNbaogNqjp9KU1fAnmoxhc3uT64P
EoIaw++DEjvwPADjjoxkpiueo7r/uwfIOZtwTYDEHjZY4jMW6btYRFkpGCOwiQsulNVJbOaH1OaE
llS8r74vp6VdmHphckyb+rre3zvmqk5fDZds3PgudKQAZGdiEHl3JMXoUGYQ3HvKBL7H6m42GzEH
rL2WmVs65sEIL2buXng2B5j/C1l/GjvXOtRxGMiwXQ7G813G++XmaQX3JC08IWpyl8nPu5IVyN3c
WkI/anglK+SXnbm3tKmCOZMdTJL6f7iP9B99wY6UR2EESUflEHq+LwoIjyT96IxMtYdms2Nj5qXS
KPm4cDKVkU6OgVHRbZL32P2+Px0YXgFYjHOQPAWbcEqsqho/L1hXWn6JVLLkZfHeZTrBaxfXQOTj
C6k6oT30hAb36ejOQp+TiK4BR6qpFbldKGbjaFX1fk5JSURX+Ty1Gcdz4xmx4liWSI1Z3M3NktR2
aJfmQC7FcPRnocqcxr9FxGMsymSePF+GLnTaR1O0XgxXd5dZIFqH8EjQi65u77cdY1HFp3FospDE
MPmUUTp+emNsrVaekjjQ3aQWfl5i7gbJs9slS9VKyR8ulY+aMQdC5CIUouZ93JIVHj0CCdpYMs6H
wCv1ZE0Ky054nCjata/UtbLuRKlOZeX/Jwom+GG8krJ6vbamoKDjX/3rGXX/up7BGu2muDmljfRK
zfzzWMSJ8yDFyuPcJCLTde+7GGZozsIM39hWUAMBwDGYeMhu8dL2A3ZzUpphs18t4tHBiQjjxQHK
IZwhBBjeqc9eqtw632InudVslKnRqi3DqeuVd6vGVPiY5Vwnzcbsi6a8fkEkqDXmTPc4P2w3Rgob
VYF+cn+6H7Z7AJi7F4lQJOPw6fMKWlmve3/1xy/VgGClorOyEHZzseebz3t4gGVnqb70sZUps6wq
4aenbOhxiyN/j1py6lI5fS66m6oQWZWEqsh9x7uj3d0VbJ4ntTabOI8ROkvUHQ9hwiiPdRjcB3ZU
EtmlwrvLbiZuocEGU3pBJ3IiyanUt46rUndZ1o78ujIDFerZ4+P8BRgHqvfLgrd0Un9o7KUsO4Mj
wwOBW9DZK6batKqga+fuaYKrhMF950Os9aMAWPbmzN476pKtc+tBWWjPR5LrUfu3FqBjp+uXu+mU
9GJTHBYYXdvPv31Re3K09yh2oNM63f1S10VEiTztbH3weT4oon19xzZ9FDhSMM0C7kJpOLGZdhUo
fcDNIGceb+RRK9g1BzsZbNRTvkuID+c2AktPx5OmBbp1n3AMnrZYeeHagu9lwitwWg5fjy8h5YT1
oqfELRuyVR3r1JFHDBGRjm1OzEc4jEg7l76GRmV++38i6xLtR43D/PHaaYHqBjKPgi6tpvpsiGPp
67QAidzx0IyodxMM1jYPbXEDWANq+VVZvQHa+ZXdb7opF6e3Po2gPgQbI8deoQJck4ib/K6OzAqQ
RNTA8ba9OVwrJhZ6wVtO+NbI1dS90gBzpwfQcJP8yVnIjjjkqyiqRzFq8n99GkL4hPV5R20fFaPA
PnYMoDYe8y58lRsWzQj91CX6NblqF2NzdQvPuw2CtV0b67G2njrv1rotINpezrQuZKWsEIjA1pcJ
GjrrXFb1m2I05BhNu/rvPHFPh/fiIVDWRdbRhJ9h5cP83st5XHU4IHdieF+uhXIHVefTrB/mI9Lo
kd6kNqrVreeac3iFb1D7RoQhe83wbC3JgEMerGliNFJrm7P34LeEr5eKntdNzxbuuTiAapmeieNu
tlPWgS9Lne41FBFWTa6lvO2p8PqXaZYllBR80r+rYR+DsPDvGAcAkTRr6xpKNL6lDnDXZjglX2Aw
jLYIKM2ZDp28lGCgcAgYmG0OYnsxgUFE2kWyHnMYYKO8GogqVC2xAidX0+Dx6GrHa+hd4PGs39PK
FZAAz8lK/lp7vPTBwgKIWCWVw4RUAwjctMyKs4ObBOO23HJvZ/LK3PrP2xwgVbB6VO44V7e1BY68
jgmowQOE5EarE3ESWsdDbYGAo7tlwjYmzE0qbe6f/5j8O8E+k+HWy5RbsJDBPNX9ETT+anKdKRxY
THn3W1KYSpms5Xk65SzRgkD0E1RCZ8MoZ/VqVuh78490Wp4d2zy/NGnXckntP9YcjjnJ4O9JOfv1
VzOTeJNV3DqMizZOgm9iOxb+1VApQ8j0Zym62ESJkDz0SWpkxZMLUX91ITqNK7p0BRQcdJcmXvAy
xvXilT81MJ8b8T3ayz7IuBiRk5v6bwb5qD0ib9swlLczx/5CYiDxfFgO9gC/cyCS1965gh2BxB6Y
iLia/3SV7C9KXJjIXQlsn3g9IEYJdFEn79lQ1BKFSlpxMCX/t1o8BYDZWfzJl3yQEFYeLLzJUc7I
kcMdlWrCpPDFEhkBlZH8v/rve6LZV2MftThocD42kiJNRIB/rnWSRhbsnjyWOyxwJ4AEJMBqTSar
qb+KFD5+2qrhDwHgCD7eN2xlSJM45y+j4xmF+FJCPuPDKv7A5M+tj+9q6JPfgBRc7EPapZ/qr1wY
zOfdOuVjiSQl6Cq/fn3ieO567KuqJRy8x8Vqq+mZQLXECK3+Z9S0otGNBNMedNccIqIiEQjTr/78
k95xAtJP2tI7XFkaeyVaySh7I7LCb2DQM12QX075Dn+bj3q6OfaY0absZfILZLgg7xN1JITlw/9j
oQ3B5xk+lbh6Ps3DPSLVUBylQcYAhaGAKQhkl/+7/DFrxIaN1NbFejK1NW+w1aqtYUzngzTMA4gr
4LQSOyNuVRbT84JozTjmbpbH7WtD2/WVvwOfsWd6i5EPLIMXwtAJcgSHHpriZMOTZje9cem6Tk8/
IwkHwcLjA6V7NB4TP8EDuh2iEWYqmubOBETFSFmZ2E1vxgJwdsPvF+uXzTsTCjFMi5pYlJUTAY6J
vBby/76lod4jEwSWfPmOCPW36wQ4S2godBnBFvOaY7vcILWky+R4nbo5jI3Qu4aH3kkej1UrGqRl
cXlv7FkN+1flWjHzuVHJJQcERPzDEG2jb3noE9FkGmFJcWw7ROBe75Z9Y/GKy2KFjr9hg00FJaZ6
y5dRHlboVC5Pk6zPD537HTVCPZxaEdQKAOX2BB/10BezT4zVxbjtL7ZGhH1DHQtRdKveotlcAF6H
Wn4VulpnEbvD3o/OXbR0vOvupmAMgoT6gcOoZVBJeuxxOPPcaFIW4iFpRuDtBvO63du2M46A/ZzP
s2PbHg3IjuDD+xtBDYLg3LRWm4rz/HYHQkQ1UrTwN7OUCm0E7IrV7wQ3faksr3JWnTuItq47KtV0
fpK+Ed1xid6qhiCyn4nfFgsz8mJLISb5FiApY2Je9fEbENiBWiW9ftEL2Js8eagTyjHA2Mw2o+7e
GYaj7VrB9YYgez3/9t1pW696mhSQD+CQwjLnGP+88L8aHbrtCYdcFFGFAnjKBi+0V/l8oVEsHANN
AgBDm3zWRwoogo/D52+O2zkltxN2Bb+7/DbkvMpW1jJQTsOvNQ60D0CO6xjzsjjhwu9wvDALEx8H
/pHYO8rweKqW3pZZk2vzPIvJaPSF/Hi+janXEPMsQrzUfPv6H/r+IFOnHer1+WBNlJyDqbgitLfa
rIOWMlR7T83U53IKgxMbvVjiAEy3ImnVNX6T7OMXbOICKwjx89sgr/NM/wFYOfnwUZGLDoVLpmBV
KIB6HIjE1rTgXD/Kvryqoqoml80xm1XF1C/7fnNzamolfNU1E7k/1UmqvGxqr8CdFaJjuC6mNVRS
E758G3SBRMIzP9g29e3/EGYKynCjaPjYLkcNESASWtfjTvT0bKRdRdMSj535I5tS3f7N4ycF/b3H
JqduO8VmCFavfi9nQ+UoIzTCP9vs9+llKg+ZYZG5kaO+5r6kFZI0Y+G9n1YIvSAe8ZnVvn1PUsnr
pSn8I8I2msU0bLymnS+4nqweK4ueWX5SbNaaxXe8ioYqX+hO2ESjN0kyp+o2FeanSTySgmu+iaaa
B9URIjTFu0cwpts7tHhgmpQ/cVfraeCFXDXjz+yYWNcevif61HrF7iLGjy33ZYssxS9Z4TM9TD4J
5nMoCZdzTFcmGq5WyKMaQmlA5MjtPBuJH+Ywf/LyhIOfnks3kgcEid/p+H17Q0J+pWpwR5Y3gOVt
66zrqi6TMpIVa5YJP6aWDmtXMxqkNjRuxtSKhMMf/Kz2PTRWJadxRq2fW2+m/y4yzeRmUWXP+D4a
wYKSPyU/d0+jIDBjw4uJIQ17Y1B3aOMk3gGTyOnx+4cuInnlpqa6UBWpwkRS82iQPPLMXdZpwd9c
JqUhJ4oKVOTAcAG/r18L4H69Vw83uajmSLoRQuYhJuIJB5S4PoJ6fWMWzmMntX3B+74MEDovmBZd
2In/7LQS8UgIykAkcCwmR8lhCpIOH2dfjkF/5gnhnOMpHO0LeBpSWcaoE50LlBID7wvc59GmN5IF
i+3HrD7Q7jfK9LNV/To6owADGgm7VmH/MDHxafZJSQBkwFRD3M8TH19x3nQGjrLu0AchUekbn5vK
Zn1xFJgIZosF4rTk6GAjDhpdaThHnr8cT/BrZk+91B8K8gs3B38LhQnD1iExHW7+9YFw25rrnu4w
0dPZtCOmc5xfjYvW9NRzZN9dzmqQBxx7w/ewL3m3HmNLErJwhEq4s9Iz6Pt+VNMVjoF1yoOUUEC/
9hWs+YXzEonPHgFo5AM7BldBpwDfsOUpMONgrnxhU7yw0L+q5xlazg68fc3bxq9oJvtiOCC/Q0dS
pUTNZdRZtkJsAVoQRoUkxWgBtsUr5ponxcFzdQ1YtY8Zl8RHd0K9CxBKO9elo62KERTCaGgE3uxl
YGkyxg+ilNP6EEFvOhKVIW9i6qOS5uHV4GB9ZoAB64TpT1/bTIhTfTSKEIAHUSvAgvcoYYLDpxmo
JZR2erP6+Swm2jtmFPxYlzImpDuNyq38bzlxoO5C9aLHtPUIp9plHeitlQ1Df3j8AbwO29OSLB5T
+XwE4GhrSYjHWMGTRWDrnphuoOqbRxOC1rirfApA/5+2SftvAnhRdGso616JhT1MHVph3EAsITeM
K5YbebxeMgW0EbxPKi0PE9538KTf8EcOo40tUkIA0OtbXp5M563Z9IvOseFfqNujOPIHaX+X58Uh
tbo+9o99IXwzzwxe1s3ya20TKdo953EvMFpvhhptxC7a3D1cVcPxXSqFvmzh64piJ9/Xb26SuMww
k59jaYlLIdTXQEWbMTFAZhpTd8nhM6zJuKL9BNmidjNbCcGuI/dmv2JSdw14bp4/aCEWQaUfNDft
zEYHpcTnUWM0/imQWsmSQv7P71r95BkkoWVLEl5Gqx2Yy5dsaAlQMBjyOObpEx9snSXhj3+WFQV0
eSBehrLLr3J7VwHktAB3SUoMWFhqYkP6JHHOfh7wQ6FKbEz3r1ggVOu24LFovJ8MLboW4TS9z6Go
t+1rBZbzqmHkIaHQgWo7/AiIQCWxbzAeLwhLsNo3f4Irp5ibJ7PZpbO8cChyzznlHsVuBEh387tB
WwhkziHeU9OR6SvpNo/7GY0h3yCoA6WFBs7X+0k7EvMPmS6uhP/SSW0m7LZVpOg3cjIN5u0GXNAM
ZmyXyngiZ+68p569t1r+vky18nvTBc34VMxC1KHLzprgQie4Rr1Jy7A4dWQ3TVQrEB0rFBETswaH
ufEPYCvERKRIRMEUcUI1O5sEG3nED9zoYwQ3UB/XJvyHt+jhd9arMoLqHCxczc5Nq0ikxidOxRFW
LavoNy6Oi7/UtkZLtnB9atkZBquRJLql2WXq4xA2ojrIFgpCpiwAHePfjrgkryyf5qNsBiQX633V
OmkYjAFqp6clets/QNUxl8YelA/MZOv1ZuL94k2hqADpO7mGEcv6GX/X0MQ7yBh22XkaSLJl0F0Z
MONS/wgiY7GmM2Lhl9Ehx5nKs0GddmEkOJNmnN+OkMy+Hi+Vof2k93a/Ldt2O6nA/blJePj9ETjS
arXgVGkFdVmPl2qrhWbyVJ+JSrbI/VmwDT1HB4NLfmwqMnlZG+SjHD4KNRsqWbNQSEv101lYNk9A
Q4wcjiuRVQAP9r1iuwKyDaUpr0F25QWDlynow08H9blSOluPw8OC8U/bRx5A17syV7Vnwm9W7XH0
I+9m4khSAMgIlVETPO1d8z5pAIhP1Rh77cPp2bHU3W7HyHCqI6SKszNw4fRvaKZZde+SWegq3xp9
P2P/7fMp00quV21ow3yDAx8ZjUrXITn7QV1vp/bWGxUGBm3cvp2uzmwhYR8DDHI0iHu1woZcoNGs
j7HDkzpsWu61IstDe3LwtUOzLZHiaeOHJr9gI/fbZ1EHapa2sLNI0akrB5YDEIrWpkQ/bm3orraS
4+IcZmsM3m1Y3JgiAlmKjuhYnONu2JHKf/eRTrgQ300G17GNKBiY6zTLDIfhnNozEgwB5o5Fo4bA
Lez4kdi1pY01ZV3aftpEQOkCcO6aRayaVqTRgWTVWuevul/8Zq0aHcq00QUF+1jHDpnmGMs2LhtD
ahzokAeldUA8R6LJW1Y7585sxaXAIz/RpjrfcF2DM/A5Vr+p/JLapMXDTPk6iTchyUv47oiitbtP
VNBUSUTc9TnQUbVUC7xM+Pqk7PfBZ0E1Nkmvp07tK8t9n4rUKhM8khzfldgjmIOyNqFqdzBz4QLS
7PvtKAwovvZyQY/tcWDHmsCUiNK59vHYzF+EHLiZxuhYzBA0RWdjjs+aWu7LAquixJNWhYsNTkT+
vLG/48sLoRwRT8R6wGR8pBOX0kpeqMiDirmJlqHwoc3NDUP5FuVnFxcnZbM+jJCudN5tRzRiNEIk
s5m1ghO+oRaIomdBNGw6TFtL9zG5QvZ+7zmtlOSPW6R1xvL3aUlSDwAkdoKAUOXQhw84+Ev1wogS
7oNoQJify0mo+ipQCMaUXgJcm7/islfm44Re8hc23+6QRlmUQY26P85lTSmYW2LVcMclfcLjfKDl
lXac940icWJ7Z8AFcjxTba9A+21v7s30QZPYXCagxC69M1UFU6Z18SPdyN4b7ymYsKQxqjMW5TsR
SFBreyd8nbkdJZcMJVVp3L+hQB1M14QF2VAAiQfdHHpl2qWt+K0yAbJkRQezAw2R6klI5nFvRvfd
3plpIh/TCbyvZomvLc0BPw1jU3T9DuCp8M4oB+AF9sB25PJYkp3c2oRmFLwAg/9HKiUUwJgkPS8z
8W/BjFl2gPhGbDWuLMZ0+Ej8OApEyluVQCW4bz+c4UuyBmU4JfSgX1VWVsa4h98W7z4zyOpcyo+j
xCOzoVVneL4jPXxzNEWs/WyUxdnXOLWUwcEltt21nRKFnHZkM+uz0KHhO/OnZIcBZrKiVA1bpDvG
0qTDR6ikHDtqOhGeJSsWKKMaaY3AHAzyWtunY2zRxBw8Zy5hNCyIoxvDq9BpcLDBePa/pRLUplxc
mvek25EHs1B2Lv3aks1EnK22U0EPNv0v2jb81PCb5yQduun96BEpWxx/Y8FV9mJ+b4sLCR80AT2h
KKn2fpXNkyLY/zehZNdOqwQyQD80+Ug3nrK2ovO8Qdm+vHtHr45VXra9pB3nanxUcIPY90MDd7+s
JQ70gUsRCAv1E9KTbRiyyHed73DdTEt3qVCUeV6rkPLH6aHzW9RwUtMKEG8yqoLPGCACY8t7cTBA
eeATl//n0PpTPLMI5CoDWT9J5qlkNdq3Ns8MHRpSBHu3dzO1Xl7HeE2lkYJkbJ28plaHJnLjKGGL
e/ao1KzdH1WNDfVF97gG4xkBo0wWDuJNhiJ0jLFzbYknaJoNSM5WZ13/yQsbqTqh8XczEvSCOr8A
NjYWcptM/3sX1eSCAo3kpnaTeb7TSqn7YlmasGXwQYHgIbRclub3RgoPOBy9jI++GQ6k4WhVdiFQ
dkbn8W2H4mr+fPFLuJ/+G6Dhjk72QCgL/VDFBhcQkVZLpzO9OmyD3lE9tzGzW2uXPgj3+yylaBGU
v0Ys/txw4MxndE26iVwD9RIhGhzvTngHfGjq4Fs+CqlI3G5q+NiV6VCpdxPwxa8hlA2/xfu0tZzK
A1db5sVtAIw6RT+bBqR+P/RawwHxeErBOUSsl5Qp/xY0TVSc25SBVCFP/vWCFKwLav4f1Fgv2wfX
0gAUA3utWtAM9gKYMi+fNNjmlUKkqIoYtew+VlhcJYOxscZLTDNY2EHfF44fRmnzCJKWxoY70+/2
eKNuiUwuX6dbl0arnXNRn9YaZt10TN6MIMjvuBFbqgTBKKlcpSQH5ofXUZ2tQ34m6Xfqe8Ck1y1Q
79+Mbibi5A/Bo05keeflahb6Kz6qbYdmyNSVdYZVmFoypVMUHw09Vges+vE4gxj2U72L6X/Nzu6c
7ztt1rpg/zO0Hfy4QLyRfgfZ0GCkpcP1YTlH6QTdR0mkHLQaj1lGlmSb82eCNKWAfBX95gi96OER
xQB3PZbZVllPlfUyVrcOQtPEmceHNF9GvIVxZOW+czEvqNuFNvHWJG8/Q80edbWgD4o0dDHIh2sG
O4pA+r1L9xXzL4GA+8v7DfNCQBKEn4IPFv2DZ4ctISHItNzLHISqZz8Ua+JO0XcUsflpVUjtYZwx
8vuVUU0dYkWotibk4ei55IyLAUZRQrfJfvq4E6VP+QFPPCajq5sfuTNR3PRN0Sh/rWrBqrZY42pu
D4uOKuxsgLIH0OHBqV3zfCLYKuIpzvMKzZHCQLdxWIG0U0udYNdGuUHGmVMPr4aJ62kN2/WwTsbl
lrGNlk9eoduGwazXQRE4lELL5X3MX6gLi6pd27lHKcpae/j6OLGR7M+B/e35KWSAdDZIfWxfNvP/
0Bk+9ZIPl1yI0M/wh7Q7iiWixDoCxVWu4YowpU1uFwb4/HuHv3lzwbrXkZF7mmy0pcKA/dCo6Jfj
ftC14b0lGpe+Xr3h0uZfRllLaG9mo35gq5UMI6lyHfhpxcChLxiBLEkiOvNw1QPXnIu5NpFhTSce
mPkjvVwgQDlQxGFEEX0HkQ3lGm093KwhP1cp7cybxEQnyjPnBf1JhIqKE1tIrfJuokmnmr+4A4qK
+Rl16XaQtqC+5tq6mBwkIRAEP2BpCkp91d2EqlOCJjx6qapBSNK4x5ZiXBMLekqPyHWDxZyZZgV1
h708HSh+Z/EVKRT4q4Lje+HvldyZ7hc4aYb3pvQazSLJglSsOgb5VuFGhrAsosPx6GjjOllSfp+C
tPa6SKRmAmVM78gC6YC+UQFHUB7D3YzrEDiLtaHA82E5LicchQ45o6kbtLdHgCEaj0ALo5L2GSfS
A0qTC5iamjfN891G70Wd9WOyx9RGpzNcEhMiUC+jI8laOEYtrOpl+1JEm1GZSWqCZ5xp9EjA/5T5
vbt5emkmRhp/oSwxbwO1OjCmPvgfty7j6REO789NjeM10LcX9yRd/s8ofYzu78d6A+w5D342GeS3
6km6MDfYmg3dQFj0kgFIsRalxKvBHZeeLiTVowl0kgEIzFycWEk3xF8kEV9qq6G5uAMzgvLndvR9
A9vvBOGTW+1xLYk+fx85ombxZZ2s5rxVCl3VaL5KWvDYgbE3XI7HRUsDbU+wui51udinGHbhmK28
bFezAUhCf1PMm/43LU/X03bl/Yk/fBX6bMsWT85Cs5Fya+wxH50RuTO1lHrybMPd8U1Ske6Trz46
R0X62IUqgFGYILzkMnFWnPJcyP3e2WE5jHxxsH+AiTJeeYU8c1HE5yWV4TBy76VQ5gGLvjD6Qt9t
UnahtY4mvswbulHFePqHHYj9qASMjBTc3Sohg79C8sPIJvPk5hrqE+r2x/BCx/nmZ7+IqoGQVvNL
IEFpIPEeOkQbDP3Hrbizq/y01D+X7DA67jF4c4YkKTdAdjD0LvE5CNbdhrGbybUIuiLqOEG7aMh3
3kiTSG3peVPrhvrcSHL+xp306aBY4SUE50sj/b6Y71hYdVBtastbSygRE96WDnSGkAuBXk76PsG1
GPAiUObmQrOg5ywJ2JmAAdCx6PUSWiatqe1CzHw9igsHtl4MOkYN5bQqcwZMW5/6rVjPs9us8t8c
O/W+AAsGe2vn8glM4jWzsXTuGjQ4fPW6CwsrXCnUon+sBOeux7YJK0cehc+3ARLdC2hxhsQnASaU
TaA4Nbepd5QGqjy0gzGJbTTTvUe/AwmEKklasT9YJyScM7Mz3mRoijC6KC6yvYlkY4eCS0/6Scka
zKlue4C3pUokKH/qrUStrV0DPJDOlZo0jQzqjfRcDy5Bmcr2gzfh2XajQo9e/4Hx8HsG1RorB99S
OAGC5c4+ha1J4u4QOCIOBlMDgAjGH2nO+p+w6RRDTErn22+1RJoOX0i+Dq4kHYrtTaRpEOhqFW3T
aZhWjZLznlK3Ft4I91ClxO/b8+xeyorQnT7+DjiAQV51HHsZB3N521cn4mYLemPTH349l7kOvWkF
QtRYDncCU1oHfNdER/owLOz7WWiLyWT4TRfjlrZZ/FBCSMsAXay9AgxOL63mRQAyM7Oagd4JRoeZ
rlAsw+/PoVS8phhjYmArxdNk4Cl4t08Mo5hZ8OcmxPsTS9DTj9aPkvVtb0ECv0up6dgb23zpCOz+
cFMhubp5f8bbP4JeysprVMYU2EjH8ouRppiKMfzRTtuE69GCX9AWKuEzvjmvcqf0ncw+5BNWziDi
3K31ilGmd1YLtx79/4VJZRYdxmovgKo1O8TKA5zgLCGQBi9//Q/JJripWbldD9EfI+OVtZWNVcE5
cRRb0Vwlci/x9MgwQ8P2Eko/VW0slwjbldFMp3FYHKxl4pHtxcqpv3atvBK62kthaU368dJkzQ9a
gtGoHdpgpPbnPnsD2nEh/JoaC7fwGmMAMrwHYiuOszWt93nPIl2vg3Daf+7pgT2a8v1fOj4yZlzO
brfVM93IaOJd98oFyqL9O2bbS64EExdblA7VS625dIZ8jvvmhT0HHIhuCSctwV2BNHygEyBMIqfD
fPp40SjbY7IatfzEeXPHm5SLHJpuCSoYCd7H69aRy0LSq2QPU5+kPOt9Uey2h72dZrijxHYSHfVE
t6H3UAn92+DhxBYhTHYAI+xWyBvOVxjtLEhg/+Tg0lNRAGwOQtkc37jSLI40/fPvXPU6ApV/H4ZV
SBp8SvRsFHYS5nIe03AzFP8QwYzS2AfVlOveR5MSnIuwnI8JuNRLEgF67WdmZJYVB9nZVofpcm1D
uTFSEjqWnnAafp3nq5j40bhooodiJxTnp4T7n3SRgoBhw5x82OYLWJk7Hn0Q9UQFC6P3HITzy0b8
yD/bzBwm9q7k9z/BbabSH+mpbL5recFZP90NssFnZI1PV/chgnc3nXbeFy10uCI3Kyo2+3b5M4SE
ij0oItE9g9cwDpAyoeEtzs+DkE6p+x8+uK5XhHVROwFNWd/8wJKcuacpvKW4FP8bJQMPuv11C9bS
ujLQaElFG5MVm3DYlnB42+51H4MGDEQB/6TL8tKaaEW+DprSTgMY6CDSV8MorgwIck3kgIW5o0QH
SRlnusCC1S9CvB7Sru03XlPb+pCkDmNV/bOSJe2Hd0HOc6aQ7NRknbwxQHWxpxCcC7DjNKeTpNqq
gz8LRGQR1WkXt8EIQDKW3oImudX/jgX4AuBbLQlE43og5ZVClCoxbckWI492+YGA59LjIKLVhmBB
WZbNQGfwadynQh44fYPYnOr/Z0fKYdfmDe9Y6X+QkK45X2IshCnYz8jc8c4ltTqXWJCvZUuBQBCW
k0IzxL1x3Qqm2KE+5JVdtnk+DGHGi7FqJp2asL45PE2oVYbYpwG4cleNRk0UJY0GaCk2DLVWTsEL
0o42Aa6dJamHXkF81velBm9b/Q4E96xq3WmjpF2SI7qFT6GMMx+uWdcS+eObBnvmnKNOVErpMnZ6
RsTgq3KIOMZ5ZMBZe/bghOrYl8oNd54tWbjZBYQqdtqIEb8Lxjwn9k7BhTT0FZbiBi5F8VvaR4cS
ID39T22ALPQ+5kRdRN7GLbZU6Br038r9P+PQ497fPQedP0D1o1itEPczxLcvFFJA2DXVQ7NBmmCE
0MXjlBCjxWa9d9aSbAZp9m4R8ei99o1Ybp+8M508Jo4fWTv2x+xiYj+rrv/aQv2rUSpFsrM6fgJo
7ce9RToUm0tWah8j+qSPvQjCnxZi+koGH5IFE1dVb2DKG7U8c2bt1fyqMlxwwR0qVwQVmRK25UCI
hPMXPYHOFiO6/VoJNlJI5iJXmVV+VXE/ZfLEHaDhCxlaOdUBXZRhG3XlusYro0wqNKMseCGx4omC
fKxOe6871HcnVbaYwCjG4TUBSedC6jk7ySb8w2mhoRbhWdFloVsEudca3tek0Qqmc6wUVdhF/aDE
AKoAkoBdyhJJ+ix5XDURsB/LVJnxjbiSTyXBVCaRXVP78J0HSPhABDxONa3gxvwvOK8hiTI/kos9
9qjNto/rJfJhFM8pgtkxl5a5azDjX4VHKjbuvetpYZPgo/w34z/TpRGV0DAjn4G3TI/YIGMGPQjt
S39QMWdEWVPFTvMfIWMmclQmB15xIvXNqBW8aJxPqU7GP7Oty90nXBTBxNUTU0pcZo21F0inaoYZ
kI1/l29C0u2UEtikMhW4OPAFT91BhrALD+E6rx0ky2K0R6W95CmmUvhDTucJ8pQPc4hNxH6Qzlfa
wdZywi9I1/0xirRvRZWgg3ovJQnMtg2h9NTtAy8HbHC/5+a4uvjPqonhYfQj9h0aFGNpkT6yaotm
6f9QdSBUWpcxr/LQNbQqE6jRGDvuvDo7cMqJHactUGX4BgvcnAlEh2xo4mvG+kmHgZEm8WX2avN2
UZdje4cKXGmpq2o52lNsI/5glJK3obnhKxjof+KvK/EmAj2S9iwx440utJF8tZozIKVITXpBRumZ
+O/N4EZ2Li3Yz8phFK+WxEpb95IkA27JfYZd5JMN6J/onMaamHSQ1/0s/Hg/LJOrguodMpAiT03i
9x69kwc/IkYZojwtuMmCz1ij0YeInk2iPk+bylni/5gbWw91tDJH8IZQ+zuXL+x6ikEae5qTyqhv
fGCEyWY/l5BgqPs201jBYJoNu8/8njUHjrrXJ6K1npSyYjODOVqjSFFZiLFGiazTNycioLO/7HHb
qNqbScIN7J3OyC5Y5Sf2bH0A9TWwZxqgIbSeXFSR4XPaPzhGtdB81Rszee1w4ic7Y6P22G0BxhA+
5XNug1SLbGPvy3FBzbNQE1vft4S0o2ZAbmeC/9BerzsPXsIue7+N91vWPZC34CNcCcgIV1RHjLjg
yNOElS7/9zLoYo/1K0f8+GdVf9pZji5vI8IxnBBwiUaH/GN8Ht0f8WeaP1Ia/CtA8FPscW32UPvq
n4huHTrrx7i1QbO22pSAnhoOF7ysIhSdsysPqFtXS+dvISu1BzoIb491MNn5SNdBE1fjzy0O28fL
pGcCKY5t832AK6oPDop+4562OAgGJv1OIULI3hvNdoGhlPoISjln/6u9NPOucf5uGB7xYiV46p0J
LFiKDKDdaD/+cA5+APEgX4n9EWaikZ8nEpOwe3DjAaiMqLWqKbo+wbl9Ue5mh+g3XBDevO7zAfR1
M+KES9m60PVY/4DbJacbk3Cr1zTo7tVNTS6+mARBs6UoFoy32iQh3dcU2Gw6MzfGeK8sGrN/NmAy
8T7btUNLLC4tTsm3LLaAdrrV4jdFNlYgv9dgszQNmOZJshYDSvdqkT4fla/TiyJ5FzhwCtz4CxdU
Tp3g6KAWf/EQa2a0H7J2yVPR0/YFJxxfk14nKeTogAGwf+ncTo87HH89bcfU2OVETC3S0gF/R/nl
wadmmkp/Fwh5GcXfql03jjY9ZWF/bs81JhfiE5IfZAP18YWDSb3Io1HbP5ZHxrhjVwqq9R63RY8M
2jeqjovUheL39TWsDrkJgaJNJ2LtfFiBXAFanuA8u7bqqHzPnufirxlHHVAvPdJMkE/Tfh+3mIgs
dtF0dib+vfRvtK3G+migaE0kSJ6ado/NsDYPT7yPmVYzEU/nW6Uh9nYrBttIHNycUTDMwdbJ74IG
FCw0Iqx4jcFBTPZKFeuJ8WCr/YlQiZDk0GNDY8mudhfVhTilFMrBBrIzpm720Zfaj1BgBIOzeNFK
FjptJ7/DJRy8f8JhtswEOVGW4OlzASHqR5d1dt7K+mCUgAizOiIXC3dKsgxEQgSQD8HRCZZN0ckO
LkSVIrj7U+ArudOmZQaX8TO7SKc5QwzwmGdqWsdXwkY8EbnrQtvpyZwQieMdoVXQmv/f1l1iC+nX
DPX60lx7quALTZFqPsgcSet/Pm5mqgIn+qQEVgOkKYVgEagyZrpqurky37yvr2+WY9qNBndmbmlp
FPE0D8EojAhyTd8mPdASvztYQOECnW2cAcsPCEFgWIVOjumRiRI4Df5g0AXq6onsjMnJ0z34jd9W
YSsYNkaBZYjS3I1Ft+mKqG+B4yB9KKo1wgX/dfJUv4An4Q2W+rQq4U4D8RE0rsmLnU0S8oToY3UV
dZnOkulRZDdAb1x1VXcV+3JL3U1FjGIdhajTinnUh1MBV0zg9vLntBOi0NHVvD6HxAn/a7hhj7Ni
IMtGr1J6II9FdqhXd1iCKIqAbIWve6/w+2yzjd7RMCS5c/cZihwpducjUxiMjPcBMXIGrYRpVTCA
5fw392hyo3DqHDyA87gwH64oP8hCRBoIY8YbeC3Tc5qQldFnYlnNBd96QwjUec9azdLsv7ffyBy7
Sn3d6zBzgmueglX/jxlIRJGcMf9jZXDfBLgTCPh7ipSnt+ll9VQf9i8TRMd+ArIHVjC3z9PDJ8Vn
Ck5BUO+4UxAEeHFBf4uosSA4jZVD7nVC5AA9H6yTOH3GKnNWzRrA5b6MyRWe09TEoXuobP1Kyuwm
Y3clL7xrU6HClOvNU9k0450d+1t9172Qbye4sa6Dn6ibHUbZXX4A7sjoL/Fkw+o4y/yizqRnFvIN
3I2SyvoLNdIPXfS6MHPkaQ+3Vk7AnjHfM9zBPPzbKjGYonyUQzwiSK+4Te4V+PhInlubkO9xbAXp
c5jVkYq9AlhrRvSKaDGmoJqowBGkh4dXCxH+i0poG4rCzGybr7zHCVY6/AKepKtKVBML2ndh1BEi
yZ9AlavJiq+d5d7nlAOzbP9l88OuczD6vP3oY60EIKad4OEXareyH911QJJ2afR4bIGqczh1NAN2
T2iQcczCcFubBVDPVGcCQr26rLH/kGGK4/3d23Tx0I/464ySWIc02fva3PlDpAA7D66hK3BG6TWs
g+7Ip995A3IFcFog6Mim2Dj7XV49kDDQrY+ipCKCWQh/TqZ+qDesOe/P7fq77uDw+xGLYCx3Ysa2
g1lr0/QFpMUUwRAms51YBj0ypa7de0MPcU/Hg9QKIwpe0SPSwa/9Q8M2FW0D8u2dwJmYZAPRMpbo
mAOdIZ8GjkKgmztmfkYyTrNePWwcg4oQqVnQic7MjLGAumf4a7XSaZ2zolR5GyzJHqu/yTOLh+Ci
QDHiGlMceV88/8k7qoLDH7KCv77lIllioNQq6K9oBcfurb4LaPr1sEERmzyc8+gDFHFip6xOgu2u
dqau1xRuzsUht09ePLQKQDde+se2cz6yGGPV82kpBzkUz1jGqzAfU51prMR/HuUm/wAHcjf3MpVj
uhK1GKsjosPa7wi++uZ6TFcmtlLvac4+QZaCaaW+H17E7Yucmm5rJzTd0DNwZogyz2BuS1/tre5p
OQsm8zEijiQZdJ8kNI3/KZhsb2sTBY8+G48J5DQe5iSWjtspsD1X2/TvACWQzEmIfX3Z/yaR/7oD
QGr9mFwPFag/xIyMIXXaYtPA6mD8W/y5nIRew1hBx/6IEUeZellobHx6RQw2Az+g3MUQXxHJSK+1
3GkVBT7BzNnGnLk3DsvPtXSZ+NktHt0oVRNUr4+UAYl9S+v9YAwzDnUhdKJ5fBqdcWEOxyK6F+MM
x4CAV4swkX/531nVUoFz+ywiy1XgGfREMUQM4cJXSDJyh7z21lJ0+RAkNVvKq5W8n4YhQb5sasLX
vM0kz294eah2pfkuUvldcoob6oMvHdIXWlHtaLRNKnBgLMpg9mErT/jdx6bSNSDz/SaOhoChTrbj
Sn+aMrdCHMAt9oTXLHH2L/5y5LCOlEGJV1BbIw7G4PtgXRy9mKET5QZBmCk5MA+tLN4E4v8n+zFG
Ycb3FGm1k3bZIezMWA4ty00V2eX3u4x+/jjffPQSbcBTIunJ/JWFBzZBF3rc3zocDcm4qzXADM8w
woAOj9alSTl7pJDiEITu/Hak4+Kmik/9tmuhFj5tjXLNEQRkWYSyls1xG4GR314f7pYnuc7mxYtf
iLn3NhFE5MIxFWf+fiHXXoau1PWkLFxUalv/qAvHLTnULWMMUzs6d72kENxbyHXTxQITcI0pywoi
EXrK93fljZW0aUFNd0586wBpuCOAYSD7c/JCtpk0KsnFy3+HSV+pRJYfIlCjRfLXvloQ48UmodR7
QCF509dwVTf8Qo7g09oWrJxcjTJnpN+OZW68gslADw6OD9131gXFZilQ96YojJCe9wEEiMMKOuS7
3/lftduJ8FRNknpyofRPdE3w+p7PrSljrwfC99XJDle99b63oSLR/6o4XNhpnd36FXAVJa4YijBQ
hNVNzOtYdjLQ9LqUYmg75yyPvJHuT6x9hH/PLePL1JaqRyTBLLopY6TIv18Y63wpvjRmimbULA/b
F+IanSN98IHE0PV+9beNzoN7a8nWg1tE4c0L0FAUXhMhjn8b6lZhjeaaOpkrQaWqtsxu8Gy2jXjW
ktGWHBvW24v8rR3dyeDRO+f1DkZ259mSdVjf2/jTokPSxd7eZD1wAzq4SrlzVHfkFBfWNdHFrjbz
HCWqu+93GZxmbWk+xJDYgfXLbwOtgt9PGQx2zbXrUd4r0tbmfb1/bD0MKsB0MRaMyqc6F6JFoC/m
7tVLb7EvYIyOlt06t7tPczQp/cvFiesMEquce3YJwzrCXDLWQemn72lbv091SZB04Va5UiiO8T29
rOrnZEeA+G2Fa/c/KaICO/xXfGiUpQGPiit32xDK7OFsXVdqdbL/scqf9yPKuihS1zrSu5459L1J
Vt5zXZK9J5IkCPJ6KtSo/9lx2wA7ePTwywyBzdlGJWA7q9CQucixUXK3+tCQJQ6337n9yfBi6T/J
3YsDSc3blMKJhHP6gmdWbAzpsd+fdCpqCYE5U887ZBm1UOaM+bMHzTclUuaZfYRnDkuFFkjSfJqK
oKdZu3JGMD3N8vujs4Ablfv3XaYXGeuC7vAh6P2HE8RHZm2ZFGHioSlJxIwWibWDCCWPeci93Akr
B0WQDZ5JImycEKMXBelPWhv1avyCCHL8FjYRpzCRyMHKCIwqtwv+FQvkk/5R/HC3lM6z9D+5owXn
An9nWGsOENHycIMmOuf8WFQudNofDw4ygsp3EtKF5Qs4YE6OcfB6gSOiM/G/tU9TCd40nskY20ut
bkQhiY6lZDiwqPDe28dCT1T17wtYYJ7xWxbnvRjZV73uHEY4jD43kkCPxdplsh45MaLNogWOOyEU
i+4s/MqhFbhCsfmY3fv3LtE+QZ2tZHU+YwgDlnegtbb0PPEWSjjFLfz5B/HZzl/f/qi6OgEljKbm
53i99HrSTxKNbgJD/mFqOs1zLQbyUGy/geWP7jsyCI8BD2gScEetPcqUb0Nx5pGwovbx9yIcVdW4
QJ7cGJHVOJ958nGGWhT46bxjq5BAzLJR3c6LHPkwg1hhbaLkT2vTtqvjXjN2BBWWZum9COlAKiA1
wLggkicM4w7B9O4sPtUIjQ7D8a2Ad6A5/lH9XILynnhWBWzbX+fmX7+14LC9Demcxo5M+561ENKg
9sY+0RoctVhOHlfIRuDsC5PdOzdTN1w+5ynaOUBuZHD+v4JspofU4SxGSepQYvB3/jW5XpPQTl6o
aShZnzwUmR9mOF8eoCWxn+3RBrrE2GJy5suJ45cADc0zyED5PIqe0JpBCNe5K1pADsgXPDd28Ajz
VzEWwv0B74z7TpFUUWvfycEhR54u9G/3HBLhtUk5RQMpa5MmvVhtu9NFgvLiOcixN1tlAPYQWJTQ
XiQMr/LWYoQwh3U+IFijVRhgK8qZwRQfgtNPQsU9zQee9O7OOs67Hai2ei3GE1CThnmJ2yQrw2lH
HbuQjqPV0t5iIeAn5NRCmFpuuJXjuheoZlxF5MvNlpnME9bq2Vq2Yq2bCm9jyVaIe7h9uskvDlGd
OXDa7Pguxp/PWMXg355JH1n/QuGRQfugX5wEcpaSo6WYYZWIXPssEELbucGmVDUm4gGSxsqbNSiN
6oYnquUEHGM+eDr1UH4bCFbFv492crHQPjYA/fhj9DT9lWqVCdRf5XZ3J9jn2iANvWofnzwBgVWK
+vVlzCuhayRryqw8WKxdkHuI3Y5AGAzoqwDQd2/GGM/MbHLsP1q6Lb0vFupSM2vns019sfLx26sB
TKIdHAywXnoNOXIJh4YuSYjsZYlGllP6yJ7E3B0fyvzvMnFBvgE5tlBx922lB21ysQC1sMk+oSza
KGXIJDOPlJ1yJoaXar/d6udL8Nfa96rPXk4jfj0bwccqiqoWrzEAhMRpzkz+QCe3RvfuvI1DaNZ1
srC8ouYjdpyTeJc5oOl7Lhtl1vm6iKDi2XueoFwORiCyqbV9gE5M60yRZSvV1Dau0l5jPFl5hNz2
dItXw1gN/FdbnqXPlt0G06dnsNUq5b5B/NHiAxIoV9733LSj1zZ3cDeI98NaRRbpNCfgj4BWl7GU
L/pGfRm3zUXN5gtuxr2XxA2GGyfUojTp71U+7NRPitEODPzNdhrZT66yGb2ExqC69zwXvIicrNGz
XseJ5cvAdTPoG3Q31pphplwyj/qDbNDNtXs204AM1F7mtFOVqLH0UW0kFqC5CNG7vUSpppnTTKUQ
WM1hte2i/YNaaSBxdpKBsSwtfCdqNvOGiV5sU641qqeLvl90OO27RQIPzqriOnZ9Rrz7YDbJnGJ+
E2Ksz0rK67ffL4CGk3HezvG0CpmPQtQxm3MQ8SIhZ8BGSzqgNF+dNqzj+wyaLsG8a+hHkIFI35VN
grYBLccyzGj8JNs2JCeChr9h6Yb77S7RAjr/BSJRXhA8/qExtPWtWhhP9YAMi2UMPu0WcXyDThz2
kKtc/0IBbcVS5rwvNeULXI9S19hoZJqS4Fy6/F4DDMmRU4QkG97M5jFK19AdWFxWGNiZkR1afZCW
QNOs7r7dhcjvOzj/UqaeqgoW4eY1v9yE3uu2A9DDhrHJIjTEGWd/9hAAPU7xi7eeAF59fO2fbcYZ
ersUM/VED68nwjDNmxCnMXR6/o+HH65oCIM9PSHJ8itNu2OLs9gav86ZlpAvjRRvSVJeT56q8Ioz
byKB8bnT5EGUqZ3HBEGU9e1H3miGHdnGp+RLJlSjQ6l6bKLMcomxlvYijewmcttrGGiO8nZ4a5o6
8bzjyMAOjaunAsFstaD5z68OZ6rn+AjJd+0claML/QQPmw4hPWh+0x8SwPLnSEUR0mK05nYVEvwG
xRIV5stTPqDjSEKUdO52c5BU/q0sDrOYkN8ojFAZ9Se/b04JyPP4v4hZRR1veVdCcRR+V9nqIuiD
X5sh4LYXOMCiSsf50lsop4Jmc7c3jZRNkhi6y3Zccmd12sQ0kntyD6wiA3cf42RAi+TV58zhvBQI
o8WyoFmJSokbFy+R+kRNHmyq0go5rzB5msekzM6PUwlZleoX7kvpiuSBheT0cjFTFq86nGkVqZ7n
CJ9DrmaSxIbtYLw+CiBjKMECElf1A0YpCcYOWggxb2sS7wEX1WmBrweKXSbZZcEUCc1SGn2JX2kz
wRIbmUBFFEiMQAUnO25ZD2rkayenyyWQ5TqiHhKgyK/eiWF/yRkBsQ9ha7SZ5S8Bb5wJiaeGGbnM
L+Xd1d76yVonytOrs2E3P+1rxLiqV3GfqoaMZ/0q7AZNoRl44Ax+K1vDM88WJ+Bs7xFRLaI3axtH
7G/TMOmWTG1qGwNTX/rx3WbmVQuLUoTeOc11CjY3g3nQ97CHSAqe+rpSs0WS0EUMw7WG5yR7m7gd
d3Zj+yTCxcGppPCDTo3oHUEX6wAxGzvIsy1IcQ8i1WYPgWzH6soItOfRTf8c6M1OrjfcR2+7TVMm
gG0H8BgH09CWdVMUdctLSTEg7sMa6pvU6Xl03qHt2YAZPHc32RPhZta5Cnz1ZFb3iNeErsH9Xwxb
KAlC5VX6FACmka2MVkEUPxwCaLVRybxVuddkATx7pJ2QibbGcxBvHOYo0M8HWCmul/GAdvLjLNaV
P3rMNoziLjTk2UCu3edvIvrMdnzKi/pjDhBibXBvATmmyPE1lvQqzTmGEf484YQ91jq/nHf2SR2h
j66U4fAvDcl9K9DGQnobRkloR1SfA8BIwEIPiSKVxnK5YtKLvZg4Bm3hgTXNxNTHFkZBDxW/Ozm0
qAYk1cLiln/En9zVLx3qSGgOlS3FzjKFTFdSvTAuYwjIdaCHmiuQXeK4d02xbkhXaanc46/3kmX6
JD42NkGwVI4tG6jUM1/l2axl+9mzhw6GG7TspA5uURrsn4sihYgfzVn+dayfxFXYOHCSmanakNUS
//rNUn8s6Q6F7xE4JzRachCYQdUnR+jbaVzpO1p6JQZpArxKLt9POOWgLqE+h2ijeO3AauesMTvS
oHfZ4o8hSTDKCv9qYDi/hz5DbPkxnoMRcwNH5Bf4RAR2oKALlR0Cx0lCRscCTQhPC6SO/Xwid6dL
TCACHPWpxbuNp30DIulLi2jwRPQRpUksjV0PqhZd/oV5ddAEk1pSUl9nfKjK1EO99Owk+U4G3yBU
6kBm/Q6FogfnTX8C0UjcqdSz4D3ax7vI4tV2dsDDLqciaKm4Q/KT2YZF83AnY15I+hkeOYNvM6pN
QGiJvvp2HXaXgOoLswy80hI6jPGy/OYclNPlRKO0rrrxd8Zc2KH+JiWoDgXba8bi9DrptJxJRKDP
wzJb/tN1OIDIgG6C1WGpJF7cpPCAFSeYKlO+a7gLLQqWWd1lEHJeow75A0qfSP7bV7yKq7Y3+WCi
KzOvE6qE3NppTCnHx3FnsPwCjFpvezodu6JF23XRi42HVxqLyy0p3Ftf+VnV2vnGEyE+Q6vmnDra
O1McQaLqwK+dE4UBYrpUf24GpyhPtWLwvwyKq5eudVHDYXSstdD0P799fKY07TGLLGlKp++i8ehz
+eYQ2ilYFVwpWRcBghTH6jclAse+Az2eJNuIZ2u3ZlpRwucd5NieRQWXhAwIGUBfPqGjP/Wiz8w7
BHWr5zCXVZnMSqery9QKBGKmoHnzPRhy1l8uzSLNClYzSTBZxQin/8IKtSJrNaUhLgah2GUX9VoE
jytaNCE4uDuBArfbZyPdgZIeFZ+2Rnpm8Lyg5ZACImAESoW3m1VLEiqp0fTjprM5hqQV1rl749Kn
GcYxkInbPMNAqMcFMCsWIEoFaCSotmSK2+UK3mfuZpY+6FZxUgSPmrTIAUD11btQtb2x5RucVrDs
hHvwuurcj2oZKV6apI0zxTZGC3Nu/QJ2weFDxs+7kfp3fEiSmfPg9dB5q3y5xKdfHpzs0+Ri6xkW
YC4Z7qxFZMOYR3dpbTbDXxcseMblqH4lrHWmN5UB1FNuKIy9XCv+g2UzYZjJ3yPnX2i1sV4EDj5U
2ln6ZJCDpF8X5/mCX7mwW5zOYJdSlU0iQmSQXzbQCGsXH6T+L3Cse/27GiVUnrceN+fgNnbQuwvs
nrCmY5jVsx/moTJct8Cl/iAtO1JHMFEIlz4c2enlcpAQRiFOpx1DMbWU68aYcHoq2XClMn5/REM1
jn8EGOPiH9lM6A1FGaypFVlV6aCw1omYKbfS4eOng4ubMi7yKzHgIH9ORzWrfgS+MGsJZimC9PFv
cJIjub+qWQ4pSS9WES3R4+zn6+KzAq3sj08DouEEp1+tQsghTgLBGuhS/DuAcSSt3whEltozzPg9
iYrYdSCB5XBzhyZpV4A3WBNY1BggS1yyVk7xeHpd775/jkIHuKRSyaBMJ4sJJPBoF0y3QiB2dsVD
6V3UbYwLop3xOVKEIFTxCC+1AXQcVqMSC8TrVzAv2EiEND9BgFtgcP0tRS4qxCklHOBL03+psMxZ
yR5hUpcG5AfRO0IaGtfWerECMg75XtcTn7xjKR0hSzrYMOtR2emGT/L3bvfwIRsqpAVuNW1HkA59
tszb/aZIlcEeS40MqRK3OJW1Aw50XH8lghnYq3RLH70G0wnFxzuVnfjRx3lx09b5ToR44VMdyKQP
pk0CMpe0K3eVUx2/H78aay7Ia+vlnwirROQ/352KXuadKJvYIy4Mb9yGcBT+bYWihWBlXnvwp/YS
cdQreVvGUdkuXY6GNtQk7We/GkIuouEUpQTXm2D4eR7mY3HlL02s9Ygjkn8RTeAGn8ntKZ1tDaAS
IZmtl2JQxwKmZpAxMOKSZYnXCJ8hciEZu9bX2h1tJeSkE9BDurrzfnLXgOsmgaLkES1CORmpIatK
iJom6g80KRYi1htpR2GJQp6fVsmSCCclJ1Jyojhyxkooh40trBWmkFvOl/1U6gXfwO5ztbY+IkFA
41vw0ZFsH53+a3FykgyXKqhrU91znf8j4DG2+EIURZNczDyXKa8eVxeDhpZqqF2drJdzmLigAsOK
OPr+2IIZKfyP/ObTW1VmMOBWRBpmblmwgbMivdvrbEDUqBXVFKzb7UboCX7Gk27/VJiR6/TPcjKB
1AuiS69Q+Fl+aVqSfjolYnz7Fu9zTwSRaGIY3ch7u1n+VLBp9a5trlyaLq54fu3TICjWo4QPxlBi
0E+3+LsXwvBCUxy0Y4banpuLUXRugefLx7yFvTUrs6wdYD/6+4djdHWXqanY7L/tkNrFRvxfL0CE
HtlXqYmf40rQvYHKSXdu20dfSy4tL8Azyj8+VpGVxDoCxtXsXTTg07P1V4OZzZtA+ZoxWL5xKRV5
+Tg2giOgKOfoL6jgqq87YlcFYmvwHMV8qv+3lwS2xgCJ4/P3/VHogbGZP5xlSbVWVykuLolWwDsZ
ruNiguy4pTRDnDN0DS0XmPxohY7KaqVxyj9tAKval0ebABWCMhOph3vY+l1YbLbSl3mST147W4of
SpwM98V0PVKzkJNsB2C3guJat8/k5nzO8RlM2yphMpV8EnHQnQ9+cD2OvIKoFNutJ85QHztxR3E2
KsgvjCkDEZ8hSa/rgw8DG1jagQ8Tm6DmMZhV6x2xzPTTxZ0jZsFBqh/0yKjhI/D5aXL5M4QoWwnK
ShQrXrfZK0PF0XdSzoJHnSQ5gdrxu3JMeaCczfjn1pQSDZNHnYt2xbrR4rbuWNMwyh56vcRX5RRR
zDKnsy3b4VAvE5hvmRUJdKemLPA/GlwKKJqzvMdDIBp1amdSTaLA7GvQ7cfW1r5jxIPB+BPXNnwn
EQsW74gbMJG6Oc7sxiqifQWxFzo8lUdrSU3//WBu9jP2izzBWXZjeJAQ6whKOMP3ufdWlnhBlYv4
OqqRw45SFZz6A8N2rU9nGA+atbHrlZOimYxh6MyEMW9jV5Pcv2AfMJSM3iqnjC7qtxOYzhi45Vt6
WspLQ+lNF80dk2fCDox5UD8Xb6aad4lw2Gye/630ew/QNBp5A5ZOumRTRLwzJI7CFB/y3CQyTnuq
wHomGCI3TWZJuk4G3T1qFPB+Yy0QOW5duWSRI0GbdZghRSIDzHrcfLP3aUfsVQzSx4E4InSqQF7f
l5Y0Z5XAaTrJ3XGqICnpQvxXZ/deVBI3LQirqSxJW0pea/wdIeSbDrUFBn25mZ71fOBZ0K0hb8Wo
x4Mti+meWI1v/x6c9ZiEwaU5p7hLjJvqzyhgqqszuiiooi7g9SRX3hETR2gIVsY5N8jwQjTfCc5m
4MqK3yZLpLYshdlchgdAobMezyUM65euQO1MLbbh4o9S99FawfPUeercPuewCWchL8mYsgu2tcrk
/iBpquepkIKU2rRPog6+kGcoF0WGVrYXv0htNLRMueKIxSkhH8MFi18sQYhMWYMo88OdSJlHU8rz
RCoNnDukDQghq4MAl4PFvF7Fo64nVfbJ2yAs+v5SbIIf/X0vofqMviuM3HEum2hguQtiXtkoaWCU
0uyrb+bx5RLOjDnhArzpE+ac+NKtMe0jQFEgyMajA4HnuTeUR2yZdIt4uYbW3CeB2vUcroFyPbaZ
VVFOVwh1OSXYm1DNhxirhWVmVbEqNU8F0BeLZLYRMYjz6fqNodr5txz/quDeFTaKzWpVMgqe8Gy3
pY/gNd3QO7HORArVsm7xwrYqNahA8AKikdfM3K5l3ryUn/cy1wKxC7H31z5icVrPV4EN+eObz1Gn
5LSN2Ghe+VrO8RIA0nMEDYotjuRyEBODwZEi8PR/jRrNJ9iCZyhDllGQc+6q1rI60lWqz4bBvLUz
fQ/QCXrUijJyvQ1vUqywuZUJktwrKojPAXET7VHqiUqYuvaGGjZlOSuqBXWWczULqWoIDeaFP7Yb
AopPKqAxZXGOjTFU2H0s1j0YRXvWb6zszkQHdhacLPe821p5VYztvQaraNipg6fh4YoVt0wYI/uB
iKYCuI9G5+RUpeIrtCewwOLyzAZa8rLyRJJTV+8BhudcXeFE6yaPOdsZliLcMxfSruccFDxDGnOG
W/zEsMMS8ZRpuP0vtY6kVszN/5cI0RrBMBXxIKRjwB83uEuTCgSYOJoffqtuTxcClYDH6j1BYUWS
6te7YljqwPJEpmROOdLLYjpf2RRgP4NELwY7AqoTnnklS+BMW7f6VX2d4nPkJwAS3cGXYwqMUhQv
fMIyqNQmrKUSfzEpZCB/3VhmVGf3L2QGEwWpx1SyBCC8QtSs4hA4/eMbkgPc7caiuPGO/gtnnSPX
hQ5jzzkXmVa5tmqRJwSuDXlMtx2Om7JLKKMoTu3MOnaBhdM+gcSSfI6lxyQsTaIK6V+3jkkVqpgh
BSY+ntE+/ZW/bjRfpf5M8TMJaZ6CHlNvO1rePbm5mqNyNIpvBH2ldeQam4RXWsyKSAYqKI75TN6X
Hz3Qm4p1fOpC2AQpzgvrskG8BDM3J0yy49jnr0vpfmvNqJlovCW4n1poI4ACs8VJ1o8i9iEGXxTH
Dv+YrpqZHqUmLCc6e/fP+hvHmDOTnRcMFJy7CXhxsyTCFhuJ76AOuBkcIpLaovhcqrbE26C1BSUT
xpic82GrF7MufruD/PQMNQI2AZVBi9g+ayvoTJFD8fEZJtGbM6eqkOH4syA5j8e+yMtRmmgKuAIE
zk0FFPtEI9sI/zdzZpprC/7dU4qjLjnUmkqqawjG23EBOWfjxhxv0dW8v+EICubqX0v7Lff4qlIo
nC0wLZUwh0iPmCqKex+prPvNbOsLun+5SixXgvWFANDY/S8ENHPULbJy5PU3KuttenIvBVe/6FAY
MlRLoh1xcdEkT+Nzjydm77Dv0nVnKravpyy7UzgcWIHJ5omsEuW4VhfyHc5K295+C1xYDY2GZJk1
Wu1fzsWnw3hdaIcuoFE2HHnZZ+cq6JAFkEBo05pR/a/QFiu6bFIjfFAspMG2VnUjSQF0Ha7gHkPR
roouOwLse7eeHNiyHGQ1hDJXHJmU7zDMmI2fOskkn2V1HavS4W0lLU3wHG/OtZQRW3ZIg2FkX46C
phFqOXTcuEvz4S6gpsPfMYt5s/9QfT/QYbGfunf2qNE6TvLGCowQxXCl34+dTtoYaNmI3MQubZMx
z/fbFbTEUIY4lWRrazO3wTbh6rH85jQ5e0kAphhERWcPJZZnHm2DhvojDATscSbxJhzvb0vU5cP3
NaTO2v59KcnhRtnwGELMOQI9Vu0Xez6vcqgSh6nGJX9jzcAaQCh8gfTI61Gg2omk5i/ia/i5vmtQ
aKF/v9qz+UPhAqshAf522O59ZySaS83dhkwgwpHFLJImqIv2IYjyuraYu5sEUqpGyH2tDW2UhxhN
8VFFXRJAHA8DpDAFoT+nHPLk4tZVBS5LI24S/E8cCHxWknvU4C47eCjOPjwT1OlBSKftvNvm0XKW
5nqNkxDUT7aKgyHWaqXHFxzYD5B9yfqKxok1CbmYmHNQXPNvhc6AtECugb7laKNKQj3k8ZVxyvcY
EuQce4FK/qYT/ul4E8Xi49rIDiAUV/rtO6fzvMLm4MjSs2I+GF4piGN3eXZJjAubiO5sJnd+YwQy
1gOs6tbhPPjoSWllwuLcqg4UKpqgprEjSnl/qNU0cfHTpBs53/8zprQTx5GE1zuxKEOKQN8Rcd7e
AJqbTrqZUCCGBjUdM/+4z4WlkY3y3aSc0hH97CDBvmWQ6n8fT/Zq1TJezo2OnXOTVaBDTcXNiW1e
6EG+6nrwtzq3ieOO1ZK2Bi/CIgRamA4DKIwCInm7ID9zriw3i5yTufjzn4mYjjHEBr8p+qjXSvQ1
jdu83dfkSt7BtDH6v4vuOVEGGvOSzIycfsOaQJQF86dGKe1PwVo2vwXavlp2PyelgqknU2SeKXFn
Zrk8qfkj6ag+oIF0llO8dq4Q/oL4Y1EJkH8fcdU9g4VAow2k8oLPwk6G4N0nBP/Cqq+oSmPsFf4T
ZOA0dqUr5tM4X4w49afX2LwtIvbwpLyqHyvj2lLyJ31zMmjT83k2MlMTiOhVVPoxuVBnuRDoXqM8
l0IjYIRxyetB9+KYY/mXWQGICBb6o8dG7+2vI+V5lxVTICOd+Stl21cDFaFwL1HqHq8xhuB/m6RJ
Fq0/SaltTfpCh81l3XS8y6BNIonzZ/px9g5XRnBSKfrSy68W4FZdz4a0KEY6tNXulnZEhihNSfhM
cu4oj2YGftyWM5LXXeJ+5SwRB8idCNh2PJpmCvWgfe8h3y5bXAwYHaE/GVfpaDO/GpS+upLxREGN
Bcbz/dMqk+IrXV3PK4XToKrFijemVXHpu137XGriXemev/eSUseo2a07VcCh0m0/QbjVFMkWlKcu
Hg706kzm36opQDVP95WrqS4ScGcxX7qv5St5BeS9zq0MgjkfdqpjgZLFuwzQutrOOaPFFWsyWTJp
8fat9Rvg2d96SDQVvQ6RpuFStdYEi11s4TGz8B4cHzq8NTOLfqTIvRGe4ONifpL5HklcEgAmrDWl
hPQNzKgPUGz1JQXx2CurSz/MG9KAEPaxFE1gDHg0c5D5OFWc6nmlZ6sCkYgFcJKTr7ElxVyuyMOs
TIeLksdNqMObjvF7XJf43pakh4mW0PIoRhbh/F7yLjLMHr+bFmygPNK2fOOSdG9eDikN75J0VJC3
REWQXOhHDO6LajjGQX6o1qdjIx8QOwWdWW1W+Gg91OyBCT1nhwlB2rUwwDFYPI5TGe7S9O1uVI4O
i7vOGmdZbRPURPPbOyYX+PJUoaHIJaqervP4V5qIrdBTQyWFJEVfH2BDiCLoJYCgeNQ5Ekl+6ikF
IEnyfrr6uMCgwP1tf04HKlp/XZ8Q8g0IuosCzRpE8pyBqJMtrH/q98RM+BfxkfgUTk0xhFGQavk3
r8ZeDnaMQ4sHtquksDJCzkh6G0F4tNJSNuksvlJgBYH0GJ0IDBksYdPL4RvAKYseFuEL+2TSJboM
EYPD01dp8z+kUji9KFfnaq40LX/NZVcKRL12a9kKzI7aOAgbW04vbiVRzPgjm81uifL06X4egsic
aFEeiOrTL3qDXQJHAOIfqNSh/ufd4aCX7HtnLQ22ticivA3N/MvR7MggCy+0uxZJlCjipComcsc1
SJBrxVwu8pBz2awzMXDP7rktpDiOP3sTraCPBFd/h5KBq1+HFZM5ufo8N4n991GjNToh+vhKCgKD
Zs8RKj+TG9N0WthVliX3gRUpe5fyb5L3mDvKLef1ltsh9pM03abvsXWL1aYL68/zUXvhEImeONAv
/FJeERs5th+TWLvHQfu0mGjBxJfCq/0SXyjZAeZUfnHwkD8kdrTKUVS2euijXTgWBsV/JI9v6bjr
QuBGzAZgR6ElZFoN978wo+INnxmIjeERQgDQKMF8LTEshhPCgwJKErIqWmHEcWIuxbhyAJsbbmSt
Fy+jnNC/yPEjLCocmhxNUia/PMM9NdydN6eErwYmQbW0hQlwmMLV/7Q8B0qYKSpDWnW7ZmGB3Bqc
S+SSiOWeYs/U8uqENEq/c4JWR3jpdXFXYQHTrVIAHzqZQ+W3TqFM+UfixY4Fz3IjvCDknXOml5Zz
XB92N/bbVSJEWgAoeqytIAOv+dpfjzDVEEpuImIBnBvzXM6rV/kG0G0BJIuR0D0V0iWh6rSBHQ3t
oddtVEyHN7Tk4J23QHnvCIJ+9o2oYvl6OtXq1T0pHJZOdS57Pn8x60mavzr1sEJ9NP7CtMIP6Hay
kERH12AsCt+qEKe9xJQEVCUSiEOuUFBdzUZAZQHzldxbC2fMxhghI3z3OqhuKoE9dh8PG6T5QbjD
6uxRmSn/UtKFKClqx93MnWBm+PNJbkDN0J1cBov+4UxGtU3mAHW5VAbqVq6THbryw3ctvPld083x
eNUU63rrj1hTEXeBD5UyuZXOm2XuHel5tFC1dAe0QQqiy3CK7LMp1U7uTHMAwEo3BZvFH6I74QsR
WvIm9QIdFQ1h/OgdJIlyIeC7TgKeBKAV8//quyTxY8xV4eGp6DgsiAqzYuNbRx4O6Udr4ecSdZHM
TdQRGTiHKkS8qgJNKIX+vSzctnuEANueLpElwuMmxN+RUgVck74nkPIhxIdNNJgBDeb9JbVPnodY
ZBugTUWLpNi802U04XyJuogGlpRbJU3pRUE+nErQ95iodtK1Q44k6uEiEWj0ghOatYg0LjdMr6YM
UcOldWZrWp79h8YkS8Bukl4jao7XflwfVfa5uFUTq/t5guCUTXPY6+BR4G1LB4HxY4EM3YT4/Ekm
H4B+0yzgte+RQfg3B0RPVjUhostPmu/7arZh0Os/x+2j43/wnKszVuYiBHNMamMJQQ17x0UQtKki
Lun2k42Alb2YGvInr/7mAoQj2yhguY2CA2BJqNLpobVxejh7SvvMaai0Fh6lUw6VCflaucXFyhHb
f3D0TVWWaz+vlF1I3qv453mQM3ug7uG1BAJNr3hBVwWIe0m6YdKroiU/i89Nh2aAyPw1Lb7T7EB5
21ri8w0uLw1gGV4wNaBQag8515o0Asewxe3V9hSTn9jEIYGSZtuK9+Bt2EKMQUaLC3r20cHe6hbL
oxXaCsPgQsDTxVfsBD7kwk28nwDFQgg7VTVeB/aQE+Q2WfkjTkLQc88rKmv+Rs1UQcPhXz+VL0uP
qHIBAE1DtPcBGL2lgcq3i2Vxnhs+wG+BpxRHx+o5e1rPijxtMw4wru/1IKzqaKvdAPAPnbqd92zJ
x4N9HrvOdM9VEiwIqFwj1DRHHQj1Bty7CZHOyDQWctI370pPZrXQCS+/itHhOclDn7bC5PbpA1b5
p3t/WC+iJwjIBdrOZONW+CzD6SwTYfemUR+92QGi1YKzbPh92HZEcZjoEzX5FRh1uF7mDciPpJVj
JIbv8bwquTiKclqlmgBY4xh3q0mBJkKa6xjLYoTh7LT08Ttu7bC8ylizmrD7mZ7BkeTcyzXYeXOu
klwxnIlZbnJSuq3dRi8madis66T9TZ/otsC7EhPbFf01yqG8Ic0hDwhk7Y1DsHxIxKPKpQYeAusa
Im9U+DlpFw5Dl74vRtmWpn3IHLcjVNNHOlMzPNIGj0gzads7HCuvsdxcwfEXAp8Jgi9hADDtYHuK
DdeBq+xzCYPk+B/WW//mAUewZABFbqxEME/7khOH/3gEd/yBzmMfT/R3REx7t9uyAQZhH27p7H+Z
lwAtoNmK7+7FyYdb9GxeNwpboMp5nWb7PoSpBvAukvI9BVIvKs4nW+YbWKuv0w2oPaTjGFTqroCY
+ci6p9QgF6+rV0SCPDAWat73/06vBllKgoqs8Yi4CNBhcnpu9IHga/kHmtXzXJGyKxD5iK1BhFOi
gyMXxMlhlBoN8jjCWl37z7p39cb7pfQo+YPrXImnmUcKB6XwI38OHQq0iMIoIoigu/RSWQl8B5bM
UbX0h1dyTTp+u9b5l8sLAqkaRzuIyiV4Gj/Pin/2Lr9O0XkLwtHd81JGxygEb5SOAyMMSTQuEr1D
EDloDt0GCd7DKcDSFiNT+9+05xPQSixWb/2yvWDxKsXLP68nbYO/yVglyQEDaW+YOzN+xtJcnNTC
bfbnrUiIIOZWTXf4XjOr9pCpdlhPFF7ZMZPqgKKwLzuxS0if8aP8IWuF3Z7k6eIPwXCP/jwEbbau
XigNsZzKzAMAfEAQ1V2CRe2B4n6la8bivpdxA3YwuA3knF4JYee2zSL5nqOYNk4FfLmU+jVYShRP
QPYH6x3kife+/7+yTiEA5+d9zWTzeZ/73zkEDnUm8xlT88+mKWPkmC5fmLM1VGL4ko31dxy4dXUo
qqB7GMyGMh8FzpGUMB4l47v9oZJGIncetPl3AeMFMswqCMOGv9SCskuw/dKkLF7u6qJxHSUJk6Ax
VF+yADf+bHjcvg4pQBnN6CtsfuFapSdXENHDh4iCl6pLQ6J7lc9ZGnCDEiMFiRW5j5lUHke+1FJW
b3sNTpI2J3QGKoN4cQXbO+mNRTw+Emqai3OZdEFdYvdwchDahtO+mmx9X44e3sxY5VTw8P5GMl5N
EyX3FA9qCKaTl0rKDoyQ3ftxifOofheyU+6w404hxgOo5+pT8sTDQ2nVJ5V4z6EfFq4SPfFMWtS+
B7ZnXXlAX7z81H17x/vvtE9qReDIj1LMOGykvo204ZH9hY4QrBglh57WlabXN0o3FOrdZ2sA6XsT
OeNWY14kpNZp3xPbXwk7KxzM1w2usjS+phnl9M4ckzHoj3KeMbkZmTKH4z/SEs7aY5WWXvKSw3AA
gcRJWxljT+4ZBcUvEkkDnSm5N4GlC7xG626w3b1H5csuopKIRozXJB+m45HYoyZffSmBidd8J12Y
VOd0ArW7EgYa3nBs0kpN9SyLzfs7PKKZKkwD3iO08srx7iwv70Nkbq8LF3nUWs7CAnhV8LV30G4G
Gn7XI2IcTa1fypbErEpIHYJCfLMnhKNUJ26Ks1OvjaqyO96XeYZtn5ci/vBjzuEHZI05SBP20BnP
ol1VjLAeJS8bTHRbO4yS7optYUJDQJyEZ4G6MwrB3f8z1GJkvTOGn/Q/VvAFvzdChI2M0hRvlc+R
hSixlmx31ncStXZnDrwLVCo56+l9pf0KtwlCCHbR7bv4ql1LWCq8OuXGtRB4UJ9zKFIjpIXvW1cM
JDAoQ85c6zMialDgGA4jPLxG6d7w/DtxAi9lVP3LWRFiBQEnSAbuqDhxpt4Y+XEE6EUG5N0mjTj6
y9RtHwIE7ugXHccueRF0EnxPTwNVmzE4H/1lTWlCfAMFhGEbYHsidfYc37RPe/r8B6jyCiklDDir
Ckhm3yKWV1g8RgY5hWr89xlenDBNFQF3J1NgRaBa8N9KM98fkYu0kuYYwQyb8MK2+fqCGu4cxlA5
c4684fMsAxQOcaJKlnoiCgAYLXeYA/IGwYVd2YZraLZvwoT7WxU1rRW698HK/v4EXFKLcEkS1ffr
jSQqVf0vvCoxGIwVagd5hK6T3VkLp6mo0UDbxJxpE9bQ6umXYPnvAVw0UkhE0R7nMkABNBkcgN4c
CDUjDz/aX+mtoSPVQtZ9d9HMatRc2IpolCVrraHSzVV23/QBgPwmaMWXoTa/HM2ccdwHhFeqE39Q
bVo4ciOddGeQCdBHe+D5bhDazwc/fcO6zSgAKfrl5oZWgUpd2uk9MJW9unfDVe95ySMQn9ExmTSC
HT6PBZ+o1G03WSd0pLKERD6lc4nWn/9g+P/0K7OqlXw8mHr8MHmLO2CJLEXF6phtoIz3bZAdzFGs
0qG57mqFI94DPvD5LlpJswrQZg6ZLUA+AXPfUURV1aggmXKvYNPHl961Ms8v6z0pqQGG4EKX27je
NdCwdGNaxv/x2I6w05BfJl5Zbk7ZSnxRla6wPAqc5Q6+aPPbIB3B9yHC5rSHtgaaSoslMe1VQHqH
gEOTSN3bUy+wBhGR5RpzbLgVnYaHrOd+/6zKXpJbDmcATSiHRR49zsHSCn6mpw91tfpCSEP8RanN
XusALzexn+wzlGGZrh+8Pg6E/d9HMZv9VKBvVH9I5lezD9I34AdEY1CnFKi2x58qWrhIsEIbWGWV
99HYF6BAZrEg1Y+4zbXda3ZJ1j6H2/JQhqJ2eFG/x8uw4N4kynOj2D02aLQ+a/Cucy08KJUlcrQp
yjzt9+Q2Zd2/Q5D02DbeNjcxlAsYdaDsKJsOsngvskbtVy7kL8mrfoAXkpffCLxu3IJpApAP7OY4
mdqo0hmj/Zjxz1fA2XfZB7Rs43IxdqiQn62mryUTX4QbJQjhx29W2J1PBNKH5/8nkvVe+u7SmWEN
lQM21T4/GgRcbjq908FJDaOLlBGXsxsDjVng5b8z6njH0GPyF6OenEK9xTiLWs7reBvymftZIewa
gUPdHtDWw++Wm/lXJ+ZCXi/ZTBYjD4+yKBQGhzzP+c5bUHFeDNndCgS/5L0nmS1W4J17Lfz7CJZw
A2wiucpnuFtR1BgmuIJyM2jpmN18puu8PDfcMKnmP1oF/0faeWa1KNYDA6FuBpfXWqwwm7Eaj2GT
56WsZ2tw3F+w+p/zF/HfylLu9/bGu0iRaZH/IvHoGpi9VF4rCqKE11kZLar6ADYj5pQJpMmNn/Ks
1iMi9c+1l7SWPpDWsH5MojZdXHiNRoaIMUaMAy8V9rZy2u36Ap7b5vQ9C09/HqYvPbVZzeFjbaHB
9iqZtfuS99bBVvdF3zfKN9j0sgXNV4Ruwd6nsYnAtudOAuy/CBbKV7KxxIMXY8Wq9ZnbG6w1ZzzA
x/aTG2ZlPl/chXWh0V3dTfc1bRKdf+4732Kx5b+CZSvRKInOyFuwP87/1ucdzRV2FdjbgaPEmsxa
vysVBimWjYDci4nvrxwbMxhX8OPPEyLIKlQO8Ee4YCtkSr/fZFkK6nvo22nvfaPQlSWB10FBK45O
9qMaGT56xjRJ0SfLb/nnnlHpul+9yy56cfxMbUQFE2vjbIIjOwzT/+TKUH/Dn/bANibUm6X28hsC
w9zkjNj9/swlx2YhhhdvogT4WQi3sRgf4ZadFzWCZcCRKNr58sP0+AjL7eR7doyz6iuwvLHFF3OP
AyS4XnrN02xE6OGc9a3WYnPnVrgZDefNq1t9JX6AgHFDflojCrPXocgjOTjPhtVgodRljHPrN774
PNcJmefB5pHWSDay61wLrUt3OVoFofUKGOOG6maOcbMOob5gjZy8sFkO5schZ7xGM64wlIqJczoa
phGjemtsxbmlgo4G/b84ftw8Zk+SaaEFpG2Hq+zQubpyvU+wgNIbkT/h2+2satHFxzWCW1LmuddA
nia+FQsGEbADLNVfmFrL+oBeMSLeqCKBdzbH32bZDC7ctVUhUI5rxHzqk4yVfBkTugim6WRNUc2W
/sGyItcT+gqnH7E8159zbCJMMWtW37dTOfemIfKUZxN5+/MJTKHn9RzZvIpZSzr+OJrd9gjJJTlQ
292xfcLz4fsIIWyM94XNpIwpDQOuNOk389JzETVqWUwtFrFJw9NL39QDBSmvSbgB+peh5qgN7TkF
h2LMSQ17NQpnFZaNqmc1kuK1fuNOiVXASdl7PZq4LeXfIVKoxloebBMY/HztdQYhjpTdrbmaR2c4
MQI8p4aVGwzJ/w5ZEDsK0Q6xrsV62wovw8gBtqCqD1lMy9lhImgdYwbS2Hup5af/hwUj/CfYuwdq
DX73Yd6BAvAYxCghLzAWdwx0JJ//PwkB5cpPu1veCCN9QNJoEvkO2c8sXvo/2i5fNUqozfbZivry
dmZSChOeJt1KcDlX7JPGWxv1H+akkIqLa7uROjoLZ3/UgRsuC/2jA0S/o9pZTqc+rkLm1Stz1dSL
rJaXmazlN5GalRStiirt5jYMZ31L8dUsPDBhQ3OB09S1/ySagIRTBH6Zx7XyrKyUtSzgzPpEbxQ9
rG6rLeDEzJL22jqRuQ/7GC+wk3h88alYxx3Tdl0x1zRNfBMCWrk+yZ3PWGiwZrBtOZ42deGmSxOz
A34mDRgLqo6tZcCT70cHEIWE0R+HQI0SbVJpuQj4x+YREsiegUpHe9t/19quYqDTHwaphPnHEypM
9a3rgFP5+h/0Psk0MkNv519OZj5s6+BzfLvwAhzTDHCZAoZqwmhKI5KDAVSzbgtWoiGyg8QIpXwj
8ZfzIdUqPaIh83VyJH7nb4HxT6L7KzMGlHnLftdq4rTCbtBXzAWFw8PYOgr11iHAFqKgammVzbtL
NRwY36IecYKYTH1L75VHqPKT0hwzSFMkgZdzE09XjCcuWHFfbPtPJk6OxAtCTVWzTrJ6Wrt6vwMc
vSj4ayo81h2RrlvDhoTdeqZI60VQPAaHqWuWxJRR1jBdbE8fO7G/DYPwSdc+WI6k++ZLzXLQoUVD
l9HbU8NU4lyWAG+5Dw6IQIbWKotFR1I2DDEW6zhKTBLvkt7iCsknztnq8Q8DtmQ3SCbQQOeRZ/iM
YSDEucuGfcGHSj0VwjNY9eR1z0FXpr+v+EyZ5qkU+rDcL1nn6NY0SQSQP7U10WLSxtg/xzy8s8rr
3ql/eafiXuR3Qs8txHsuYYHDDlUPPV3k1bnOkd5l22n4Y5C4cNIgMSPMFMkanjqd1wOWWQqjZsNN
ZE6+iCG4+8gyzZkAWTwRiNQ0oGnP1E5Rf5C6mSWLKeExMj3XkN29JB6rMv0ey1rof2f1VjDHACAq
58NDGu/5MDzeDZcqZI0zeClMPvci516nWmrunhw8phrpeY9ENnrf3gSOPpwrjQpf87Y+ZQs5tPLZ
beAR19G4N990TJOmuOZ69JVR2giiyzzBTu7c7iGQ5NL5lPHWcl+dWq+70/Micw6gii0c5xwZLsy6
DM28AaTc/1dMDwSQgI5WNAD+H30Rg+RpKi+MxvTZrZDVT7qEVCo5HuFU/jw6LXKCdYViFzQGLJSR
MeosWDSBMtMT4dM3K1XgiLHuK/Q/E5+BX0Z80DprIwIbqpm6cRLExtRet2xf8XqXjtPKzCt8Gufu
HRm3/bKKeLo5XWGCUifPckoHEuwjiPwuFZSULoqGH302O4sEO3P3yVr0vZ10bmVf2t+E3pseZLAB
XgrKFUWrkKVy+2v4WxaugQjaZIZcJCVeXHgbE87YbdQ3fdCQ2WOS3lpSJYUFmTuDRn7nCpXgUi54
2hhDiLVjQxTWnx+XZVuZStIF3kJFyO3/0JiP2ZdgJcU0J1wt8ewKbtcq7AnatJnxxFb1lrgdYMoz
h2TwTMqxBQpF5eT763kyWbd5pCrnOWo5Rq0Sd205poPWiwohQdGdFwiIgUsY/fIUCHRpCYgjdMGX
P+eRSfQS4yWsVHbjZPMcNna1ISyt6dtuuC98qM+nAbMCnQwlK5uMJlYzHC7lK8/yOUCkx2NVtciY
66VR05dn3XDLVhfhaUeD3Wi5C6dqr34N19dSaN5gIiakIt6JQSYOcHbX+Ne5AU78CUZT5KxwnEHh
aAyfEBYLxA4O3LRRcZsR1kh+EYier1oyobgU25OtorK+k/Yv3jzMWJdmrkBEuGupfYYoKfQl6f68
hKf/WHlaedMQoHA00VK/2BEE16zTW6QIHopFEpkWn5bvsz+1x4KITVLzfS0OqIrhQoilbWMn0rFw
MUHv4LHZIELuhuKC154mw6joycV6NoDVFRHgM7lXdduKTaF18XfGEfxdfgAA/lpQgkeaq4wBemEn
9uxqia0gFvXBqnql5055OTNPEpoEc7nw9tDOEt9Uf0PKv7woS/rUPr/XpSJO2vqsZvT34JXxhphq
vnxPjrzGKNo7Z3H6oGCa40Vty0cNw1+2JN1ttkPB5l21ts8KNZ3rTbwMIPumuIjUI7y1kJELSzKK
vW0deP+yxX3XJWWE/n7OurwQmpppNLvWtDPZ9dyMH05GzjtOFsQrSrnEZnSe6Yuf5eTD0h2WO4Nq
P2a9NiN2HJaCJOxMv2M40bFza6Q03y/QYdP9OOHq1EqLFMwU3Mm20XFEzwq5Lv4MS2cRmAbd008D
Nl9GQ+EZlSOFTFO8Q3mh9ukCGLrh+PwcOx0A3Mz45ivZVsZizxc/aex77UH31cmRjaC0J65C47bF
hTtKMxglNB3GwR2114Xe2jIugPtT0Iq/RRLNSYh6nx4RE5V+/360cLyKaOGUqftqsgqqo31qejjb
8Bxp0iLIuZ4tl+2oF0GwOncHaBrJMA1NbXrjxK8wg9AwNdUllwklLZWns5SMWHgoXEvCffS/oN0o
klQ0Whn5SxCu8M1FeZI5NnH/xlzeqJQ+guOOemv3G1CHX7wxLy3deiSkMvcflBttKmvUXmyBXg80
wjYaGLJUONd73460T2e8mG7GaIQzfZYT7rHQZ/tE8+7e08nkpfGDRNnEhwFgle6Vr4ZroEQtHJcn
ZtoD7apD8xsEsAM7/mRLwL1dkY9WzGzyTTsI+awLdX7PruL4JQ1eWauJH4BjJSsSGooIV/F9IsZ1
STOHR2aoWTYDJkMUH/plShQmXAhOpEjSI0ID4mCfU5X7C3bhVPeUuJqTXhF2FK1BQszCVjEQDfnT
0xbNxo6Ig9fsr+v2cUHgZlGx9vD2eItOHUqylITA/N9vLcSemNwCv+Khweble29G4GH3mnGfaSfA
te+dUTORN0340DRLBPqzZddjyfYuZDLqRlTdeqCvAjjwZYUj/Q0pUQFmre+Im386zQZirmurYh9W
1j3V1sFQQXMkQ0dbKJ3tBQSnGCnZFeemoMsckXv2aZGX4W7A3fxPI3j0MWz6EHNh34xVxhg2xvgb
rJVzDXC+28uoOWY7KCX+xA5INBkfUO4edNBPsAowSNdD8Ay3VVoqNn3G18z450M+Or/2emNrGCgZ
PYzHZLderFmpGz7RqfIyqfG43tp7z+G6yWNpDZkpc5VSp41p+qQA5iBA2j44JgxoBjAlXBTWGEA4
0Cz45LMnvm56kKLl0O1uSbnDglc34XPsvjOgwWmZohYH+3fLslvIril4hcFZ3mdunHFRlwkR3isB
SpHqba7ytgU3Xag2sSZiGFerh+znUm8+J+HcstOx6ZXH0bMTqtK3ODiaXhQtWX8LnoWXQujeeupq
GCcGsRGe1y1Ow4QaqPaArbLY0H4jenHJzVnaq+XGnAzphK2hxSkuJVfvU6yI+jsefcQi8NjxG3YO
W7IEbxOG6BdGMu3BvKETXQ2jFmQpUjDAirBdLUoSwiyt9hhOK1kFU8kTT2/fh2VeEbnh1YKNP1Av
HLdDF/I6x4TC57U2afWFVBfcdACE2gcwSnKeTWPiXV0zrVmxKQN31MXDwl5kA09WhjTVDN0YE2AA
keNYDmYwdcHljjPjgv7lC9tZ8csN60tQKLhSAEUZyWHybRiRkR4wyBPK4CBxJ4vOpIwOLdy3DOgf
+dQc5ERPu+ZtUedhr7jm2r6ZLwi3dV6iMAx8ewxf35KgEnPwksjn/51WdgjArf+33mYGTrH+zpQA
k0jHaz8x+a3vpDmYzZmE1ia9fcI6HLGSUQ52Tui+uyLHaell2rkw88M3BAVZZ4MZw4vIxk33x/Ot
JXX34xyraIs52eZHSXsu58GJOwaybomI4UQgjRSlkY5wayVv3cdvSrBL1UtjfJObKUDTodIXGD8y
qj6omGu2NJvaIqSkyXuqbhvF5F/UAdgTL1ZelvCxk5vgfJMjIf5VoHtmL0UlQ+InJYF9AUE5hddv
KkYUxyR5ttWxI5thJiKYhtuL+pDSkpv6mpwRhs+ecM0eLzpBuT9ANE+X1bkwSeoVw6b6osus4z4o
AUMq+HiCWawIvBnGGVm9hKFPocjxPZaGd1XFG4NFC0iCAdyq08ySjR9N9WoMvpQNbC7dYremmALd
jkQ+yae8ffblguy+OQf2xtNveEltGD3tLH3kK42OAGWOj9ONQ/30vR4SFU97ZKpAb1WuK+pHvRMJ
fdXvv8mAL+pUxWN3jcP+S3dqYJlOMUtpeQ6EoovhLMg+TKhAtqJgGtMQdxVr+fto+cv8HRcP6raO
/XyKIdEtjgThYxH9VIGNbj73PAs5m4DdGSwBNhOBAVr26uZWMIP0Is9QAz0DEG3NcFnqMNEqt2ba
iZWvId9kNlogyrW+PKJgX3K1AUAz7Sxbg2f03yVqnmwj+hyF6x/QozScPn9uWGloedl8Yyoek1EF
qAUx06MMda+mDV9LDriG4wAbLchq8wNGJOY19q4MkRSWoPWmFOX+9ftgQ/2YIdaFAUhmpP5zHAUl
mxsxOy/AiqbxUtm2mb4W3eSPqfGZsj+fpOGXiNA9xWPxMwvJqotNzejR30FloWZ9F/jki5h8g+zk
hV+iIhZMlTb59C9+gGinSP9k31l6T/6cuTJbkHdP1eHvCyucKELPNufNetw69RMVzy/QzhocKO80
9iWcgP1+uiQixcB+3hAPCH9jspuyHoxhDWr/VhQFARczYU5xX29DbbtSQYWmTsi15zHZUZuKbfxh
d6C5Gk+bmVIscG+IhMW+VJO0/pBCl61CupcBhdbab6zrG8+l2M6cD6duOpJDq7llX18jo4VFsQ96
Y1o9yoekXRkaNipfmcFOBdvY84R61qYSPBuwvOyj7oLpr7JXmQhVEKXuRKTB4NcFFf1IMRHznuSN
Enow3mXpREalEJW76nRVaI6AjZ9YZsrp2RLYfytC24BMew99uI0fedkOOoMdnFwUmkngz89kTT5H
16tKJm5s/Rw7Z0ANdzMQiphC1u0VUKxljl7wc6hLRj4zvaHk3ztcRghr7NF32/jDlp6qQBvoihb/
pm6KRhVen6d/zlW6utP3ihoHVoM9agAFQk8zCQ0+BXrS0Acmot52lGToLtEJcYlyTdSbWv1vViQH
c/rooujf88kbJEGYHt/4KolELVvJIAqGS70sxI+kHyp3z+KKFSNSz+X6OQS05Q77B1U+2j4knDH4
XvFN5F2WWTRB5CUQFc+GiSb1ZwfvVMbt8izKqYVfuNCLJYiHgMcpQK+zDjPoMai1zF1lA/SeagES
5MloYiYmtQg2/QqsvOYQ+/k2hfkChFOCvBjd88Sa/3fSweIG0Jk4b3kBJ4cnCNFH5aMdDzTNEciN
Rcf4lYTbzCxg2LehS+MTrKOYC9M/MrDr1BAFRoxX6VmLNtbcGZH76dgSTmiBXiMuY4gLer4T1m//
ZgLYzl1tE5A9pZDhwTTd8j7N6sjednfUZA7Fz8v06XrjLmoSd2NIShufNtd6Ae7JAu0hSKQzP7Pk
xue1GSKDEJSzY5y/5Y0VYiQbTYIX3yBd2N4FWB31+KuB4+UKs4AjsYVDs7W5PdFpkmUWZYWqiC5U
t+nm0DeicuOJAUjsjSvdo3jGRgmK5isLD27GZHkwtTLCZ9FyQy3zjrcawNkYvV519LqIaemoU3Et
qcO5bCSBAZYlaGmcL/gPfS7AlVwSIYNzSEp/yRrIYKbw5vyebGKdiHnsiL5oa7J8abJZhtx3S3Uz
evf5nXQSRb2p/kZhPg9Hj9EK1Sow/1QI79RA/gLfwM8TM9xjCLwTVV4y2WLeCpjXGGIKpmetz16c
+EI5Zh9l7nT77M5dYJbgIU4BOpuYw9M9XjouwIFDCs3p9kRoYLo+gMVqMsRackVhceilKjXAbW4/
gwPPStHhMqxda+4blDt2jm6caonq0IXgbPqhYJZWUcRqOrRxS/OrICb5Wt8MRFsbLZ+XpuVdIt8y
gnmIV0Klq6SGMSCRR+BCLWLMqsD5Y2E3Jrdh+I8DCXrGW092v0a9Y7qMpbpaQvT4EakjknM4KCiE
Jv+oVZ/X19eJXLVBDJmtlB3emkRw7VhFXrXBCoNqZvnXS8SUh//xUQKPCFv/JF7k64wLFFK9sqtU
huxLneCoJjd4dFb9fCom0hRbRrESufp6dzmbVuuesm7MCavzHl9XeSLpoaAP4OiEDMnfsL9qdg8O
GB4kPRcXueAOvQOjBDsGsGJ20QYXP/H5DuEc4ejtxl2grv6ChPEriTw7c2ussMilyEjbuSBnPTdE
SWCykVbvL9Ta4y2M8NfXzsPmlQTOHFfCPjoOfy1S+7n/FJ9AGAWqFdQO9Qq+L3uI0IGsAu+1pa0G
v5lOfVMz8ENgy8Y/ifOJ5yTAGSlR1XYtVxjWSic0DK+WJwQIDxd2NQui4Su0FbAK8z/dML9tUObs
9ygW4aGgQEQwpmSOdk34i1X9cpTK90XPw5Ykjw5Zju6JRaiFc5ppWDmL+/8NTxK2QV4lorn8pdjS
nOAQ3zi2NM4sKpkatgqKAT2K58MoToj6BGuJv73DnqXP1uCjQwPZmRFn2cl8/D+e3uEl6OyXChcf
xzkAXWGmwvJOnWZJFH3UJJOq8q02qk1zE7Uwywh8sumJlMfKwiVDJk8CWwhN6bDluCFErvvbc0ie
J/jFakrnIKS9iRy2haRQ53eVm4N8QkY1TGrGKNTb/nSKT0hBPgGBRHJIzQhHcW5d+d1adcRzBzwn
VOMgkMn9usHPXmfhRbQgtR8D8Fm3WQYzhp1h8capGV8ow9GhmlGxveu05MJV8jCwQq8yQkwjVP/h
o+NI6/6+Leo84u8M/hGVjOf/X0CLpx48UB4RUOZ50j7aAfN5Gi6mEbiClQwsuzhsbFo4GXgmibeW
uWbs2GHokvk7TsESC9AIwh7RDnA3Mm+fnpu9+q4r1guExFjO34k7uWaREWHB34KQeHMLK1wfb6la
zvy/ZvB6S7E+aMJ0pIKdtAj3ty4FrV4cRJy+mkHimH5BrlSe/wEybvyP0NfVntuP+I1tTLs9ODtZ
qP3mjh9C4wBqgEitkCA9kb+J4OrVhlqx9pm4JhzxZzE6SHXVTVaGjhy0nRqWoYs2BzWxnu9VWmFY
NWeuMI1FPztxt7Hly9Xacf7ESJdcq+umtdhmkjFtVdOQ7StYXBPBqsIRN8lP66x0o4+1yJpwuesH
gA2tvzqAGGIPPHzyptFnwcFdakB7VZarbPQqnN4aXiJ4dQVI4BLqhWA4VmY+Q/IYGGmtJteFcTC+
tQONDATwISUylIs8RFksZH23YPWu5WH2KLAn+Zn7cS1r9+MazlIzBZNqoTzqOMkU1GPdfoQ0e9LS
CS6KYKDOFVyAMuqh9Ujq8u/MpcTn5fTZj1P8ye03z4wQlw4gQY2M6Y07C7G4L/IQ/W+d2Z6vibnB
zDjSrKn77zFgv06ihz0kSm3vO6solDIKG0iF68lUk2jU2aPecHjd0hOXk+i21PWdq9c73E9XIv9t
YZEETijAIzqbBXkNmW1XQTHteYbZLxdkZJLfReH8sDS/Tn2NoTpkHp3tpE9le+LY8+kT7WUYteap
VIKlve0rRtuE+SZokVzMtrTsYVc+UTEcumooo7d5OoznHvy1Cn+2I413ByiEaQAHUAx85QQdIXxb
uXzWFSYPzjRz3t2CdXsMF5fNlV+1EFzzHeIuCbekhWPa0VPc5AEqgZ5+VAytUu/3OXjk3AeNv/5D
mN/qxmjbRjOHPEMHuau9WmCvbct/OIcejwoz+QXt5H+c6mtGMETW3eGtfd06tEadrwBFtQ1IP/aN
FXrjWA/WDSm3GcPBAbJqWhZwgvZofXx15/d4Mjv+XCVsvG8Ir1C2KVm0aZeTZwknqKEGctKFg3Lc
JYKyk24LgLNWAcUABOTWJtqLEfB8pvXuU4YnGec2gdCTHdt5wsk3x2OE+jkM2F1/2m4H+PvRajXL
pRne+Ik52s7br/9unsr8TOphhDA9PZ0qBvBMB7FEFkGSkjNeG4WosIlZF2/x0DJYgPygvKmlaJg2
y8rVQDA1YFpL+QqkfPca2R1iPDZZRiFxpTSdvG1KiUolce9qxyfQbPRCKyquSM4G1mxeI4d7fJsR
QY9EANqAkbt8teLf6JX38ygJlplsRzxh/mld/ZNK5XzRoYBJnZIyU1csRpzCDsOM2SBVqCK/PDGf
2QyRJK2bd4umVRqNjZHNRPvpP1mBiSlR86rYL7moNbg0H2fiIUwEqjJIM3xgn78mZr9jNceRQUVl
oyyORZH9VKIeQDBSyUpVhRNTD3TjGS3KLDFz2uXH7GTuAo8P+OV1MMc0YHm1YbKJQTOQUGDHpulJ
/QhtptuMtTZ50mG1DFJm+M/PDgQ/icAmkEJZDMVmOr9a8s7sjmLf0dQjX3kDbzQGHew/CZgKI01H
y2D57xKUxJTthtLnKmazv0iEdEpwmhKUpubmjN+NDuinpQZ/wEXFR+chJ5p5WjfQOMqrgw4+pe7/
A7DLnunIn1zhqrtFT6JOO/xa/WPTpjK3gZHM0g562BD28FroCx9YlA0ZEe+VV9DJac2OVrs3HlYp
WrMPnVI1GhURhWTQaOapArghG4nh7b5Wtetw9qXC89WFqxLozALkeyMsfRpfM2TxCjFYPERVE2dc
zRSF68J6BfZH7I88W/AxLNSNMw1TYNgzCe8n/DyPHZw1r5NNiCBZQmrc8BYriA/uCznN25LEPyAq
Bs48jzpwls6sctBI2V1r+xcMxtuprWL/ZcT9aIt8cfl1y7Q4nTUA5IMu2XgxycYv84YZHvzsmNE1
2ya5b9qdUxJIIVRuXix/f0bupBWgQBjjL3fKFPXbqemCkzaQJCjPMeovTpyYAucGI+Y+QexQYjJF
Q/JdJ5ei081y2fZ7HgVSYaruLJ/8MP3ulG8jHRCHnnzwPu/WiDrArF74lCv4+EDwdldKM0wwbR1U
VwJeThY4sdxNg4NGn2tfw4wDTfz+uAKjvrT+0m263FpWm05+SpHPFdcdM7N2Zagl7phtTXNnuI1C
61XOmNp2AKRAnVm6VpifJGHVerCcj0pBcI0fK1VvKpomoHBRoF/vBJeR5sqv4zO8O5GfLVTP+UEs
JeNODB9PDun+Sy1F1loa9mVxls9HAERcZlkNVg3FD79wgxujwNcMLshAGWpOJaFJQt7bGjvThEdo
gfsWXrJDh2NORkbBlLaV6tJ93+w+HmUpfBVLnZwiJlV1tBtJUMOlO7Th0r8w/7N7HhUZk0n5Ry1E
C46smxlqoNs5MewJwNQ60wkyxgEtGVgfp6EZhwB1A47fFZaDjpGpMkai2VcqajmqBaZpN4+YLPLK
pCn4jeWtgY1HQszEJy/6emQkJC6XrScKpoZ8UvbDMCiBMTkc17EikhR2ObD92ZL2YH/njvj9Yv5M
+s++APdtA3uDi3vIIzrY2TUdgKRT/GUn3KZbRC0chjYaJSLSpReKHs/gnguakuAhW5GYUGyuZDEA
bmFTERbFQ52hxmeDMepNYuzqbb728wnkAwPcpouUoN7IyG7rWTNoUnB8mldGVCmPOX0sCpbuVBN5
Bk2/ZScMAE51TsCT9KOpO1NAvZviuMZxEo0xo9b9e4iZV7SLObs3fgbSTpfw00ZiVOEShgu7Ca/U
+cyrinTU15RG2rNHkqR6M3+LfvVdUKCwWzsYWEUJ0Hl9YfOqRX+/FDfNc/wDrYXBm5lArASlE9f9
/jEbl5OXxhFgSxaagl+3f5LL1exj+ihDa3UsYkDeE94+qndIotkgtJrOj4kRuzRQanSuQCj88JEi
QOIkT7BYTyXmTc+ag12hagOEyXQh4qulAoT/lbI21yr0U/pi0tr0Xgkx/fGM1rlDASkwlrvbaOjJ
Vj47MffZOl2R7zEA+7z0Py382NSAqrqMlUyeki6z/+zGjdfKB75eJd3g0VMBuUxAqRiwWw1J01ud
0CQwEkBNZMwOvyb8orc3CkDgFS8ny+045ZkoVv9Zl2PVqNfNTmdqSVZgZBFInAjCnAEXm+Ky35Rj
DgCETDZi9CCXJg1UuV7zEKsByqhSDMDeipUvE3JVWAWJNi7380zdVbCNbN2L6KtHf9KbG25C3Wqu
3bSnurnapRFwFq6aaRlUki+brxzIAgFwbz5BelPE1ePvgG5Rwr933A61BGtZPoUGFdkgfbND//T1
0RxUxRS107HlULCupkKjxd8OAKMdJYpjqG7Ll7aeRGJgdgp3++94pS3Dt1rhqwCBH2jYbX8o0ZrO
LBiCxSWutQn4vdVCQnM1DC0UPoH/cwoy1M4uk+SwqOzEUGtF2UKlAAeFhqduAwv1gHfMf2MPIUPR
qi/W2Tl5RRDbiTvryQdkwfO8O6/G6KH1bzL0m7cc79cstyDALp8wMbjeZzugtFnnuTyvMLAfZpR8
HDWCfYRMph6wPJDX201M5dMRJAyBZXTgwexN+0ogRsw5Lm69iOxcIfszUDraSZd2F2YqKaroP4A8
KLX2dALOqDf9SBfnf1/mAk6ZcGcQoGtLP1QQT4kKdjkDJoYq61wepmJ53O4/KhkPNfLbt6M1Cf9v
jttpItfIgJnPaZzIzEIYKIFEzT2fsbYnFQ33ZD1FW7eVy/7RzroogtfgUxBcKojl5HwUVaYdGxGb
ju3dpTlT4hsfgRYi0p/SqayEoGFshHAiiL1p4NoEKRhWnGz2/vso+2i1jbZWMB7CFa2BS9yGahcI
Gp2MsiEh73xVyigbzOMxGZYk5a/wumKNa3AAvA0cSM3ASUf7fF5tloDkcaUmJbf+BzxCJ7q/Gxcj
dupdwNvt0yEY7kUBmQ2rk1a23DDItCzyI/85AHSt1heZ5XHu50zBvSsIEGJB1H6xodAN1WoJbu9W
PLsfLk/9qzRf5cvcqoTT/2yj8CZvudPPrU/M6yLUPRBRXMbLnX+BSfMyQ7/AXa4B6VqsFsNMOZfX
JF3hf5m2f9wNhVO/z4/5CQqX/ObWlH1LMnezo8IlENbm62/NrDKlGwDD4dxzZb7jGT+A/tlOtP72
OtiGwQ//FCGY5JuSnMOIYvUXScRV3BUP6LUfDrBl62AdsiqgGuj8gCqcd6M3hYvzC+862HolULFK
9Qz9Cn9vBXw0p7P51LTmkg4lbqTmvWgukGSnJkqQBuCn2BBH/DfYlUNUJDp6fZnnOTPc0O3qtzLK
8j4Ol9FSkLMe6j2iM6eIBgRz+uarJ+4zijwRp4I2dyXV/jnzDMrrEbHJ2Ag7uLrtzuINdcD7HAvD
q+LKf6QbeFegNiGp3bzZW6IXK2s4jLhkHP+N81/8Xg52vrKbL+G+hLGUz5+Xklx4LZos+Z021BST
uxlYOG41v4s9fDlD/G3WBnyUaGYm0Su1QUTdjKpvIyKEoGHobBEim051zg76Gx78lYNoUnUOrfPk
gbFPZ6f5SvpUZuMUTzRi7VPnx4MjnRboFVDPRZhcRCnMizVYhdK18eNP6pMog9CtQUo+6J+kkQ78
DYf+Fzsgzv9An0kXrZXV30F24FyfcmTq0CYeXTABxcCZ3/5YpJh8bDzWzidb9uD9H057n8CoZlq0
gY0cbw4obSE+0QgbFV5yQ7OZ3og2mIG8IaY10TQDFVPfEhcOiaoTWZ8V3qqc94Fep8Hl3/WXiX88
52C7X0TQa0WSACxl4Z8DJzfKib+umzzC2bUzyIPA4l9wI++MzR5sb4+xz101gA9jckcuj4pfvW3n
q44FDFaxbsLqbGhuTZyGCroDhBswFyYlmUpIJ4eEPMuhv7rTM/w4yMnydvaxgmSiMqB2SoL+50Sr
cinJuFKF72DdXK6bFqxAgmzoJCai6i8cB8nfzM2QxnFjqOnt1anlj/KwE515syj0VvaO6eN+LSTp
pn3erxH5so58PkyScjfLiw0VLTQ6v31IsCy0y8Tkaeeikc0EloZ3m9N3oBExzZt+wG0bSjEKoF5z
69nMAS88BYnZf6W64ODHVhP38zAkKpYQXytQhQdSN49oCQMmbL5k80xa4z1Ei4EuhitgUXDCM4dq
qOccF3LxmlEr6zBjWqotdPN9p92ymhi4vP4niu7tj2VzHwfwpgbGM1+kf7s4ZIxSyiNj6Z+zGfky
sSpRTKEMfpHFTJy92yaO8kDJ42P1UkJC5FRD4UR7aYCWANBZ+sZsngZ1pus6I6DWzx5V02kY2M7a
D0CutvHjewxfwkwI238C4ZkUcATtp129oHbZAiFludh/hpqsazmDuwdiycTQIGJcARSeUlY49WKq
mAhPJKJ9PfE+sCSshyT0u8ZXcL01KG6BTQbxOQx/8JZsbAMEXGYacCNUuoSvAn6e7NLMDULHwf4P
1glZaA23UShlTA4+XF2eEbcKY8uGG3qrrSyZ0AHRCKMUB4p7XW011wKZ5A0qHGMBPLiVG8UCmVe4
fENhWBqTR3LJ8XvupCFhIAkrdCFhu/zGLzb5d/oIz5jUMrJgIPWKjEXxTJos9Ztk4iRchSp0bXuT
7mivkcssUBq2dZceQm4H1GBpPPWaBQMymjn74cLDo4RCPkDh9HUIdNQXEljoELbOyo/BTdvmgo40
V7juYObHpzbLW06cwIt66OzqbKqUIT7gbtYbqWKPE9ehdUiiU2P+UT59it8da1OT0fZlSnYcmmt2
6EW/sPSMgIbNf4M6MeGbfo+9Dawg6FRWtsGhSgaEOC1p87nzobAwsCl36LCNh/eqWTSGxiyrPkaB
yAV3FX9tcM6sIS5/Hyj/+a43p3MFMSZP+fjsI+GyPeHhQjVc7toIDfnY0SESoIdoZv9aKl8Y2Tri
j1MuRoTlAOsbj3e9JIYF+UZ6iwDt3M9SeuB4GhFFU99L+t6bZfguN6F2SFTCAeiIujpHbJcgLcL/
xhUlbu8B0fiSPzfvjKhyZGN9Z254+z5scT3vx96sAQHOz1mMRne9Nma7MtgfkNJOx0GrZrcZM1aj
5e4URSVv16Lfc6TeBMgxBhQ1jlC4Yhj7BgCaZMPbPd5xWt9DI0cuCAA/e9jY6cQOhlZgh+3THYI/
1U1KdDzZW7tzFqOSUEWZxV3v0+LF78l+IRepW6YmZ7lm/1Be3KDo73QmpBCEMCKmkKYalsp0cLGl
oBlWqQNlS5+PFE5CGeX8oV7GWNnym0nBZtDJbFUqgIO1Q+rKg+MbDMNkkRIMfFECk1/sL6+7EZ2h
OwsEl85XMUCvbycpWsTnVEGyrKIgUgjnCpSXQinNWGZe9GoSbxKvWgn6/BSCZrNC4YZOBmV89p1u
8xjRRXoTR1xiBgIVAjbuPfRFghDbAFxtIrLwZBcSEeM6tPUMTVOs/aKPYhpnTbTKRCiocv173imB
clVKq82nXHYDVizx8SRlhyQQlJiyxPX7I2OCIeIPM4lkx+2TUKgX1TWY8shPQMx71KkU6NQAC8T3
MMaXn8V+DPqNSCD3rJVz2DABF07hyw2xq7yUDQeHexa+Gm9YPFkh1CRF47AttWgVlIc3wmqNrm6W
rBpnOl0Nga3NFNGYReJbXZIVQi2Y0h0cxe1v98oMKH/imBbgbqeXIBeAfaJuAn3cq+TkTm00ecTk
CSYlcA3NLF//FeOMJKTEQvGYZBlNXRkd08/UFyGdxMoWqRnCqUMJzIQ53ezwxp3w1JMhIu2TOFZ+
aYi0Gf7gt2wJ5GYboHSOpwPbFQlDa8fa5kJ819EAgoLA+BN8VjXrV62KVFi0mJp9vNDj0DZoN0xC
4XN53ktl6JQo0BDMMgbY5/RKyFD5lqKkg690ELyyXq0IISw/3fVgdlNpscNPD13myAFyiJSImaHU
sSyvFXRTDg0TOFCsQ4Rs0L4EY3Q57Y6bEpMYBGHJ33QhKKK/995N6kDxcNpDnuO6GIWdRdWplOFh
w4LkyRaMczQBM5G0np51ehduFx/7Ys6KEFwjd+X2j9dym/9oZ1GYmCa8E1GIOLaPoiFFSvpFwwZj
7U8EjVogCR3NeNRBX/Kux/AU9U4VYZWlF2J1VMfYSLIPeovq5f4EUVJS6LDnIbC2TZj9siCyik/Q
yaED6fh2Tc+MJBR5M/ZSu/RLhGsUczyEKTRzCI37BxKfR+jPj5BSQS8hefNMaqISudmkM1yXeeNP
V5bL5iDpH3wGXsqa5u88OR5WNblz0FttgmZ1duiMuJ8mzLey8rtcU2ldQxgkmlBc4Sh3SnPGmjkW
t+N+Aj4W65mimwiDFL1rZwa3FQTaI0KxQvG1kn7Q3We9TXQgKK3MX/O36YoNLCX6tFjfwiFovzhd
jPLvFcExRiIfGEFuHh7VG1mmHPs6kdTgiHKjRgkVdCtrIHuYK7SyQGJTn71vNnZGXU6ByxiHcHKJ
OQjF+S/GQbX5m9iAZvFnVy5vDqv3n8MdO23ceomU0dPbx2r1A6p9WJRzWO8ndBwldgNQ1YrK2G+d
Xrm8Zl50SbiAmAIXPPBPgyvLovvjrWSdtN2mSBClvyt9vTuZykwarmY5TADPiv/70G0i174v4S2Q
SgJvzGAZG9O1Q3qUd4Q+z1Xu2h2KI18fRf/RYKGPA5u0e7ignt6mFNvcNSZ6MgSxhKdE8nz0k6+L
G1ri51R5PTOX95ailiqUftrFOf68iLd4jYB2ZPoVlhkn32m4o7T17CZJhyvPlg6uZivbzxhNJdMo
pm1updkkqmquw0fYV5hK8nK3I0LI+bIPfqxxg6upHABVvf8C86lYpaSnZJiDyI9zacnDkvJ6y2so
UxjWDL+Q3rbddF0u+izy9NRRDzppRbKJe0c20J4phI/OAgbbRfyGG2VIaBx7fTIbWSz+DQ7oD28T
SZ3kZ7wT1Im8eQAXkPxLDXTqNETkqahmrk3nWYt9+BDkDeg+cir03V/eWlbXKh47a+dFPRHbWGF6
rQT+Y4SOzCEPulvPF6VXyD+0iq77nMyLJJa+hawPc7Vt9KAuIKFUnJnSIIhR22YWAi/Xh80eWbKI
6MnX9UMWLUfN4jAxSwBHIr1z6mKaj36B59OlRNKBkCjoqmGHCJb2FiCFOK7GuoyKXe5gofbqrF/p
f4Qb+GBlP4H/+8KulvN3s9iFhZ8zGOswqlbFffX6WK7C+Gbm7XCLSGc1EAq7c0YepMXoIAoPnRFG
ZkBvlF5Y2TPl9oMgVEAeI3D/C8wG/OmgtgPgEgN2VGIx0HwdKgrunCmqfxBSeZsqGeXt0QoI7DBD
hcHdhQNtWbHfnEN4kQq6F+WnDC2XHKlSzgzeNanUg7fhUP8r1eI7TH5TGnSho8w6PxJ3uNl1d+hs
Z9azbSraFlDL0VIRPAjuklW0sMznWp0S+bg4fajebaKJuDUeduqmRl3ttjbylRiCaCakzOKIIKq3
R/fBm2vMyeeFSYDp34Wp9kNpIh89IJ6AKpHwgxIt73jEBwoHWL/kfsldzau2ZMn4sr6GntHjubmd
VcQihQoKoEeVBIcXr6eRKxVToBGnkiQUc3HhL0yoUZ3iTa+/k248FB6MKrjnyt+fKXSGtUOhDydJ
For7+4rjGHvJ0+L9YXgDJ2rsLhhWWlYGyCW4PD1i6IxPw9I4fZ2+GJM22RuHVkBTDmnzSJdcp7PK
himY6aojtzndakyAjE8R3MvyEdwYWUVu2kWooRUWLLzjeyO/UrGuo/hAOV0fu5Z8tamvmbGRhGsZ
Mr9yi4pXfdiLp+I2OfKXzpAfp3MLiOKEYZeQoeiHmrq5NWloqJwby4wCD4vQpdskwAUGYQazZjn6
RuX02rA16l6UZb3v4/TyF3VYfWJi1kCP6TjMTm4Gml6vYSC4ImNKCT1TKS9zOowS5+DG29sduQ7f
4wJLfi7cQhHTJNvW4E1BFlLUGodF6GKhH/mUGEuwyFFoeh6KkneturPbTDjGe6V5wykuCqlVg0Y1
JaVZw4Wsvf9doZCA9uS7fZUZ7jAjX00F8jXrMEqOf+BXf6KzBdNucAjiydNFYzFKSgS2i63P6H5c
l4a1uSWgOZZFS/LSxxkkAQaTWPUGvj88tKkLh7WqFIaSOEA/2NcltqC4kchndOE4XIPQGYKfcvOp
sVt8g2ijzWzJhtTuqpFufTPU2/9X8LDQCTMtYImM41kN3gpsMYDg49iiB3WSy5lnKdE//+8VAEuR
VWpokJ0O80hGyi+QNKVAcd874cbd7zzoj9qxIBtYjJL7yR8C7HlE2u8y00zmJp/OoG+AqoDde7l5
LRMpJ29r8Gefm7n6JpkOwef3C7UQ+w2gV/vJMZlxGqwiXk1kSQc9L1AINUvCQRhtQwzs7c/ujhBj
QUOEAFPKqXRlmj1wfnUr9Z4TrTSg0POSlgHuRGcek70kabAMm1yR4bG+hn6zXugqc55i/2mEHt5l
STLeIlCSU/3rqP9oyo1oENtyJOR3gs9DiXMsGby5YYZ3UUkAxZcbv9vja1p+66EFZb64B561HEz8
ceSLBJkKwol2CWwObaFkY/a9RhaKRcyUFZOuXITNh8L9pcEb0eXMtmLjrlASxEgmuSvsD+lpS7Wk
0RrCmByVU5t6lXVwvLpF6maTRepik/cBiSOrKwwUtmLRUz8RBYZe2M4+s9R+sdrLhvvutl5jzoxF
LE+g1eg9briOixMhvmNNM5cYVy4AJjTPRv+STSROMDwmPh5k5ZpyCoBAgx2mAqzp6n3InBK9GCWv
XTm6qi2Oy4Yow6G22/fYSceb6cliR3yUQOteLxAhYOd/ZT/RVQF3YFVshJcfTjQbPr+qwTX6UT1D
3/OI6p012m2d2z6fG7aToq+dAvv4eEAciwMUOma7YsD4gdHTjeYwkEh+R+dV55+NdqVt9hBxXq4B
S4fIFTsOyIW/T3bDfY3OoZcPbToCrA1PlDS5i+/I5IcXK6xky2p5QYNIQWH+5K00sM9JMLgjWzWe
1p5q+NQl9TIPou9xl5Yo2rHsoeolluMFfAKFLzXGcgP6O/H5FP21GdmtAFdeDh87G8iOPVBlILQC
sSzL2XhBR80mjFpnyOnhG1Pp/T8pMkvwuoSbWCQ7Uy/BYQYc+jC/62zSCHh63nZStDf091vHCnr3
KTWSoy+3YRb6cmmDGVRkD94Hy1WetSVg84b59lYSRyNy5MwFhIfl4ig+t/p+r9Q3o7bKOzWXNuQZ
uGIY7WY6k0iHDyYuCAOkjGauFfniAluKu0p1282Ltpymyk0eE/wt0PzMfm5MwsDktNh4X5kcfCx1
VHft32w7VoePBIzuAS6fVvRqOxIdx8f0q2yp0jl6Nfn0dCokALeW3/gVXaplVPsrC+kfwGf03SE7
Ug4c6Cq4s7twZcjqgs9WwBCjUGw6S2aabai4JYvqS2M3Nlqg0DSBfcBZqZYg4jmPscFEZTZZIas2
t0pr+N1qYjOv20Ki+PH17gmXGAe2w78kad4G5c4iDzmWTWeOfcQfl8hEmeQaDwX/0F+k9ayIMOL3
95rQ/biFQr969LaE5TnGW5GHHZXXgS8ve4mB+H5MkWIhTzjikrUEQALXajYSQAfB9ccH3BJoHSrP
d9TRnC08OcCCTXss/+/FUvtbbP+/ZPmB0/OtC1XbN0UviF013tWLV6+D7u/D1eUOddFklma9Kspw
bZXd5cjAQZHAm8caLykUopAfik0pjrJUZT8PfndRekhBB0afV6Ki0EcpibDyMTYBumNz+7erGI+k
2r3qOVLskBYAoERq/FnsRw0VIKpA/VMqoGSGaHljHsXOmGOaDnOWnXRlrb8lhF8+ZH1GFxzyRB+u
LoOajpoZPd5vOhwXWPyDBe28X82eppVKzRqVr1I/geKF2bu6WfEky40sGeBLTOTGp0dohgZxJ26V
D/irz+Qvb51qRc96Bc3Twx5flRxxi+AlfbzZbiI8OPIqt1t6weUZfzKT9g0Nn/+gOMpwk4Q22zd6
fFc83bgUKeHZefFTW2fT2q+HETVP7Qh5t2T7D1CDzrJmEHuVlg2riLiRYZVFmKsid3KZbXSYQv46
CQZOpZGwscfNjF0WkEbABh3nrm5q/optdRlsMVHoN959BKyrD9+XgrG1me9hJPML7Xp5Yai0wH+E
DA2kOTI/GEE5NnTsDCAgS+Y4r4K4gWAP6Tmhdzlno27mjtV4vonVv0n0D/H54l+B8QUsPH7NKVhN
BEJGAYgrQA560G1Z9fMXUkQJr0AVvfOnpkb7hr+YXJiHj9ncG0kJEB0XWcUPiZikRI0F+eBUw0qa
qr1cq11b6hS0703vjZu06O80hvUNu6aMajThsTxvMs59SKQE/nxOdsjWxsGhXZsPhJWIWM9qkvb/
bsiiEE2UwzGcnX9pUIyOP4ZghEPAl77k0sdV+eq5aCdL0SxUebQG3x/0agww9MyCDoQ0QacFdlr+
jtWkebZc600DyasYfq9oD8MpM2oTUceIAdX3m2h3rwIzz+Kcn+6JovwCFneVKz0/5dc3eZsDFvgO
7EExdxYYlMF00p3GwhP4lNN2az3u1Cl61SobISFk+W9m8Iev0OK/Dz23wgiqjLF45z8sPpgwONFU
AN33tVueAg5rHP09XT2anXFXDglwq3/BqvJt6SeB9YEqUi+fkv3m1IUrmx3ZsWfyRhd2OQia1S9E
pQiK0gSqSbHmWUVKhUYL7AlcprUdsW15qtVc3sRnQtYEDzApUpjzJSISRjQHZuqr+B0TDSG3uMQV
E7FsHD9ELN+2NG3z2vkivNFRHDT9FbnHUOISU4yy853PoPt939N0P7KKDzIhr0hy1AQLM443Vn/F
79qx2e9UAsAzZbBXQppJi2oyPvnxW6kij/ggGkkK1eR4n7u9KPh2pCzXeobrJMQJYQd4alsmTDxX
efDLgQBe0RiMlB5n+uzss/AoCzxNCCJ13dBz1J3qMlvU8K//PFweFktKGrphSdf8MYhMXnJHWKqB
HR4WVFEA+j/9I/QwKbhtUMrl7RbJ3Q4v7HP7o0K8DEzqTgBL5q5OwXTswm7624x3fRaiyj77lCPr
lyPRUqywAYEL9pNJQHqyYIVMMFfO4InB5ytgHCp9FOOeXvXlYDnPj9TeQrTaxwpwjFD55bMN1GHP
DZyWTP+u/LJ7/B73oFIoNfuK3swmn9sSnlXxwL3F8axAZ4DWssdyLkKNxiDiHACddTygtV6ttv+g
XFZsLPL00e3u2SmXGTwgfLd4zfqJY43ZKDl/lZeFE62DggtfQcDYC53ZwduACmOZnEd8ZUUDzR7E
M0XJIm4GBDwoCJke7nYUYus5hxEqvtFVEIcVw/xxOka2VTPeTg9rRvlo4NJDrEZVQAVX71u8xmo3
DxwPg51LHGl7r/Y4n2D8O0B+cIr9VrGivwxNUKeM25kUUebzbuqejOtY/roKrzdZusS8YG1ZxVZm
nx5yS3UD1tqztzbrPgybXntuoSY5p34H6FPK9QKHdxSyEvsfyopzEgnoWbyPnYkSmvFnb4/cg/80
0O1Jp7RywpxuTV8TulQe+PltvKHSgKOxxbAiAiFWLC64+q8Xbgp6+I7C1au216laqnarVaTnEbEX
ZrbZgBpEYUjvgy+phZBA5dODvTfQ8Z1cI/Le9xvtkwSbLctaCH+5dzYCSIKRO9+/bLMNoBrfm2h0
7xyDS74zrkWXJduxVHp6/GnHV0vunNfb/mN63l17EEIEoAi8FrvnDe4UeZXhhHHcQxlYYF+qPKgn
6+L/e8qiyKro8j1FpK6jtnRMPfX8HKdWjTA0LTmHhLoSrPJD6AKqSR6tTci2kR9tFso0QGFwEeC6
1GLIR1H+2duLcOjyHa/I6hEm8G52SVGk/UyFAAyXK0p7xH++z4Wh8utfdn+E+6k9N/pxDmftMTlZ
aF108VWzqFU8wBn/UreqrvIGAezA+LWB7S5HD/ZOHzuBOHLEs+B7KSbTgUYXGKBbtCnbQFYEMKRz
sXSXeEv4JAuFoXQRUGY1ls7QZFt/gwBc8g1E8aNK0LaQRFnRr+bjhPAOSl95hA3EmvjfYREqRAEO
RAyeWLJak3DBk9LxP85/Sx4JsBUHB5LZmBawMyTEv44CLPW2WNO9OYmVu98SXcS8q9k7FSkL5+2b
hDycxGbTq9QAqZbn4MrRZW2aCfGjdzOuza9ho2KPc7/BxmamZugnda/qBpimGgTYGLNve0sDTAwm
hf3Dw9+S0JCITQ8S2+ETUMVfhWuSgDQiU/8jP7cbZb2Qg+xZxrM0j+SC+nkxVceiqE4N6AJCZ4D/
VfqFS/bAkOAqBsaFULUCdMEMusT4AvETkNVxktz3o9SJfXpqPXveOoOXmr4Ex2JWq/5+KjV42sUI
5vKL3i+6tX5BA61WQSq3P9E1PZvczmxQSAiyqHXOOcaJGkUzwBme5TSp8JD7sZdgkw8iF1VzWPQ2
NiIfhMUabaxiLX6juy+bW4iMx87IbfMyLUYC2tz7gDf3KRqboJ7h+fR6gTDj3z9635zRwqeGKBsA
j3uGB8zLyQeedfKGrj7nuHHQL5vz85EdB7NMOGYJiOTjEuiXnLoQaT2TBh6Hw248aCK3hYzOpWZA
J7gGp935VLkV4OXooBe170m4EQYU8rv4v9DU6BVAAO/8TYE1/v2DG8uMfp1mVr2IJYMCC8l+3Nu7
hOAkoMvsInwwAtDhhovNH+z2BuwyB99104+atL1qau1CT7Gj81LWq+lka5m/gEhT05cK2tfEtYpF
3TartoI4dODq0I9rEDe5+JR+H4W3Q6mvZwpAKkNxYwo3uMX66bFGc0Vtd3IcYz2IXjlu9KUEnJba
6raSW02McwJvfAFxa0skcuIci4gjffnSPQXqXsB29RKAZf/CS48UCfyzMsASY7HkHFIGFPygMwpb
ZYcxK1CNkiPpaPQ+GyyypTK4Fn30ms+Btp4HopfnuFE2lM0jmLp7Fg638XHsZB17ZUlzOlfymNoC
+C/ZCNgzFZbNrSG69W3DLMmsprUSTSVeGvBbbOf3gYQkDym1F52HhvioHT6QcpTNHKdkutdjvGub
jZAc1/3Yvn4uqEwYZs705h+rfXlwZ1LMy/D52Ij4MsYOtf8DTL8RajxbaHDHDd0pFE3UUSOoAAZc
kUX7PxjtNxdaI9cJ75+rKJ3NiEANyKLfv82Gr3e4RLhEe9Iy92WWqhMWayncxgTPADRzyRBxcsjO
Vpu1pVQwK6UOQBeRS5oH5D3q3jliJroF6bI9oxOdtrEL3u/FMXphzqmOPqpmdCoZerlg6DS4Dgw3
ucyQbPRBRJUNC3YtOcK65PgQEoKfHnOanY6lQqOvlAWmP6LdynT4QmYqFRd5AkptUxxYVSbIMui7
+H43vZTG+blu8+IBz1yjoZ0jRnhtlF66QnG3aGHqnZwezMVBaj2JSAWIvcwS161B8tsVSnvQhbQf
TStErwQ4oiffzfaT+n62tGzSCkkNdqX/hz0RzdSuin+0dcg6BRFHix8N1Eo7t2DRRD9amL37bkph
WoMZc38nqWTS22lFffbc+BllYeb+vmnKeYDGyHFQ4U7WKvJKIOCvCmHVNPZErJCabLtAenuc9b3f
23Krs4G0/+d94G69Y/ZI4SMTCfWdqRDeLwrkWIu8bho/biBFZi5zMBCyZ6heycRP3gCpaV1sQz3t
OAdXayBEGeWggvpqjXMiutWmhpTqPBKx/PA3TOpOEN5lVP6JaDNdezzi0N4+GIGt1lF1vvNKwW9u
Yeroto+sEzKwaHRnwzz95AI76Y9MJuSm+Lwuv078Fhqai1gq3LlBqd3sSeLJw5y86lMFPOl64ieR
unK8Go6F/fwTmL99FOcICamXL43JQiy4Lfl90NKjPQTpviecqiYfHO0teKZdw2q0kNWq+WMIsFW/
OK9wLDlpwoRYon4ZRRfP4Iiugx1zF7lcwTdPYf8uvyXWVkz5CHjwL1zYYgGGJrMhecQTv+1hn4UI
rltUZYZ7yD6AxTnzbwbdoQW8a84p0BdyRodvMcPGY/WiiHoBFTgm48qaROKvJTVkoVcsaEWfHqqE
O0pGPS8PIsaVzT5xNHipssHJdMEIYaJDG4BvmztH8/4HEBP63fQ7bVXEhwlRmVjJeUM93h6tGR2g
0TxhZHYHODkNoyM18TKm4sPkhaa5Ex0TSzQD+linLS1Ty8XnTB/3oNsKJ5LkW9nA85maazb1GQhE
1GFeNCN66W8woQoy3jUO1AHRJ/SGP0Nr4sbwi3hlHzzU88o4pqw8voZNEwqgzaSW9fkXoYvwfyF1
QKdRx6UI/m7LnrN+ctanQg0F6Dg3rW/fcA6GB6RgZ5FcCWZHFyRLvIWd0YXxgf9mAdXdczxpdg6F
Z1qaVasOxwaeHX0hHLPv8NZmb5MgY6rvBBigGPaBD+UuIBC7Un/3VIqML96KFQjuf3vNPpswlgeu
3820sdwR+EHyAmclHAhJBkHXO8+TXjm2xnsZpmL2NYh9pzS3tcZ9psNQne/VOy3SfSon175XFCPQ
4GfnS7pl9iVI78YGY90liEfdEumIetFk7oeTJqEfDJ4pxluRz+SNg8Mv8ic2G9xVD5D6QAdoaTBY
5zD6SP5bkRJ2vB++h4m1RqvMGm07/w887pp9xLwRmv5qQIkzyp/vHSP7SgIjqKSr4T82azY8JR5B
hOShPD2hVExKfb91P/aZs7/Xr9EFlce1/MQUY35EmwR2Tscvp8qZYNdjibsoMV5TCRL8tsBLfQHY
NGqBXLUec5laoeA+G88IS8uXItJZOL9fLc8b3cX2CebT5I+MCzf88Covve0Aig1XJoEpgNWA1CXA
zNjh2U0qWjZMrNwobiCJVgBnRUUZtWi/naqmFOTwhnjvvzFQuHZoXxSscTDhDNOY2lJZ+XqFIq4O
Wo6rx88YeU8v9h1s/wvM3fhpXVgYkFL2B5RB1wffrPXKaq8cxuDK0ccG2FaR0TucqiQwirLkq4ji
ChyRgTp+BR6Enpl5s4zdm6xR6wG3N4WYmIxQGGYQK56YZnW7Pne9cR4UIi1aqWAbcbT8s/32ysul
/sjVovM8LPgrP+jycu22QnvT6tbco3YIkQZ+WQGmE9SJRqcwswQz+rTTF3qin/fMkQF5+pO6doN0
KZcR1IpcTnqZA8v/3VKlCOZf4wF+GXGyRLUfMHtWTde5P8gmJib/JjkCQkz5T8vKLDUKNbBYGhbd
8ORyt6tOvqEMNup2NRxmpwlxJ4i6YJVzW4wuvaRDKfnlmUENa5dTIxPQJvNvQPfILt3FPSlANX6i
3EQfqco+if4pinAt/6suDDgoQXbN6pLCpjtj2INfcBTAURT9q8BW/E5m9NfshOlplActMnulfrtp
k0CFulYK8Jl/UO3WVTXbxs1oER6pemFtKNLLgel/0Gmv4UvCQkQEqQCrzcIuVVwXO6AbPtrT4607
Fx5U9LrMUlUDilVl7cufZ1p/KLMPc4o9UQCXXpvUW7WoaG9rNLszSrQUoLGI2k5ED57difpeWy6M
c7Rtqn/qgVuy2p5KlXIPQ7iT2o21mqX8j4fxKUTKfXbPIPNHbG/+gWOoLMILhG+MbLMauhRo+WGB
jX0+2wcy4YnhE3F9Eku847spx2OV+B57mF6MmlNFxiBc6geJVmTOEPobvQdga68GUcRYejgeExbK
coRjFiZoeCnOhTxAnSnPHvstfxdDWf6cp2AoOmlf0x1bUKUpILORGr6ub4BJwLIqEq/B9/u1d/Bl
tW83I3FtLUm0RR7p3gDCp+/1Bytfs6kLpa0mUnqeKwG8DxZNggdp25TJME6QwmzYZiZBMT57tSEY
8POq1B9TiYJhRUrpLWWjng2GUkZM8E7QeW/HE4sHqo5qlIigO9tExy4GdCeB0i5TZ9mn6iw1c8C/
YgXkrjIaluCQkEkYE4W0hlTGqakcnTVvoHUjTT6MG/oelut1tEoK1YP0aC2RSGunV26MxqQ3f4Yu
sEpylIY7uHcydKEZN92RWFUol3cJS28TTnXot+qn+eDTjhqEkRRjEkthS217SQ71V2JuLbVu7/+w
YBTfwJSm7d9qKSjJLIFKKNXM424/b1oh3a2hMcEqEUvb+NSXXl2jEXYi2DNeZbQPcWiLTQukQtxd
vfInThccruVuFkKYiKuQqZydm6bXUaKickmLkP6URM3oiVRWJ/gAt4vreXd4oKVqGpeut+vuWHYg
haSRdDUQQ7wraNixHefvXgkLii2Y8VBXghsRbBtrLtFt3gCdsaIQ10aAmHDCpwOhVApIK4zmFe4q
l2m6+jY1iGH+Y4vfS3nYszFUQmWG2xYvYi0A6CscUQAjwIBUJztb/tingyZZG+yw05jzAbNBs8eh
C+2lr4iOW6mc5FKbdWKVxKKcjksYMAPJs4JVMTdmBKKRmKlqDcgRJIYqgRZPalOOJDpUHHpajgec
qGKyrjSFBpJ2cVhfbYD506JKx62SU+lXQP0BjrzSky1TEYc+etUP0Lbt7zfFO0bbKlQrNG6iNg/0
4hlLzo8YxuB3YA77pu+BK6Rvfp7h7LYFMgdaW7F7lfqV4YnWx+SC28XxSZhCMZScv0rez2rI6KwQ
bBe2era8hmfWM6kO7IjnBz3PBwbaf/7dikciPyEGw8U4IMwPYSxsn2cKGviNF9Qct68UJFXl0c6B
MPSF+yIHvcoTlSrkRaxxF4zpZLDGpAJvqzXrKlFvGLRHfMnkX3LSu6jKMbr2aMQFbOUtgNcOrfyT
gsgCi8DNGp1KHefFX2HSzx6cIeHQq1TCVNneZMWPTUx6YRDgfMyj1EVug+FU+wfMKmBLpK4pOFS9
HHDa02lykmD1cg1TiHEodskr+r/ljPMsURLeCy95tOlgK09weJsaemhLpjwdP0sRsX/Td8VAKRoh
hTN7mA8e6FXRlNFCMhjiI/xsPq7vACy2J4YbIEbxfhYEsSbJKB37N2ooGjJtzn3zNys619okOcq1
zvRNBfl/FkjIj6xeWR18xjqSaGkK91o1cEc82PCfOUI+5OPO74rtTQXSQob9e2JItYWhGayVFnhG
Vf0pv2iyCNLRqvFen3OYNree53hyMHyIoBdqR6LAKdTbshhy3Ogsxe0hoVZ3dly3l2mhcYs4Q6z+
D+S9/hgLTXEGwnlsnheH6ko5t3/yCi7XQRyfCLb/FwAz0weeBj9Crv8uxW/v9DPqrX5phM+S6KPn
BM0n1EnQr0I7zlLl6iun1iHJFY1WbQSnm8JczLl9awtLxBHWwzuceBjrAHwV5lt3O7kQH7VjLH8M
RSDk7J0FBsX6Q2zu/DJvQkGb8X8PS7aEiYoiarDTBiUf1BjzUyN1T7ADr2C7fxntoRKgr1Q51iRU
J5/PLMZVwTbmeFYc99/iBY2bFaHOpFUy/+i3auUwQ7C9NItbKtpejw0EVpxY0WrcMssLyKjxQMMN
oHtYyazZH/DvgtNWJvtLj+t+qBmOOHhhr4Tl7V0wNQ1+JoTIemkjUXXp3fl5D1ZMZBrOj6HfLzvn
qWt6BYzyF0OkdOcAZJ1H3gI5y3FeFW9CLs9kRTA2GpkvZUmIvULh2QpOFU4ILDQCUqzKx+d8viB4
S5jLy7Cy/RhtjvpDpqoCy4cnSwoo4rCysEuzhw5K6ZVGHYb0XmzWOxi2tiZzAogm8Xtt4jpRhQpF
Si7+HmB6n7ntVdyTXK+dSMIn/5CjLCellCP/MXY086JOKY2jEmDvDAR9XNVyg2dIJH0F/PNe5HPe
Y4VZhJHzjTE4qxttrRZbu7tojNUMRF3yKYuzTPGHVX4Kml3aA0RyLZ2N2Rxt0z+MC3U8XqYS6Yhq
tgRzYZN35v8hK8TfWJJ/L4TP6FokdJ/dzXqHdEo1iGnauAFylGBc5CdKdpP40ZF4UDu+Tb3TiQGI
vvd/KJMF4n7ClyS5rK5FvPodh3yA/j4jBObGBg0+t2ezogRndulPIoDrDsRhavPuSPplFjginHcE
+8PlVaJsjzSs/BODX08jPBkfjy2c7rT5Eph3gbJ1q93p2in7Hud/XM0eTsjL/77mkcfztyPPVDaP
pcJLmWzfykvyNrEZ3ZIDr5HktUk8ucb6FTxMd3vr96WDWyJGNofezefP+ZjTMQfd1sUSjlpR+w0S
3KPXMfS/lMCXoEhfITT28cNpurLDFw4zcn4S+8PlCZ5T6mhqedlKE23UEM/A/L67jLDtYBXec7Q/
oFlSm0KO6vx7qNd2KHxX6wAOpfUMjh3ZzaF8EpJoK3W3/Hsq+hGD4dLrc0Pg2ra5udTvBSUawgHP
sCjX1430uxiJHk2CPDfnmwtTgb8UyD5BiRwYW8jh1spn5/9/NSf6JxVTMk7wIr8gs8ZbG3duO4NS
47zzxwlRqj5h8/+k0vvC6IpHvQZ4fmf2V5HQAeB0zXKxRtlFlHXWFtvdBm3dE0qosP9VQOUvJxbk
ChZljBjDoKwMPfwO3x5ud7XLgm2casf1g3hhAyChAMbR6dm3taizHDSsjlRHSQO4Vx0I0RjioMXF
rVZ8I3LkOKJ8S2H4Y220/wn4BotlwlyJMXB7Yd50TfdVPExImpwAyaniZVZg0bEP9BlT+6p44+JD
Fj9xJSkDPMO46tB2ObS/sG2P0Y+CO8XInr/93BQczkiOCBdgJ4t7Qyq5dePCdjQl2RQQ+youk2Cn
wPJiX9HOmsQ71tW1LnhS7Lulm06y0Qe73Wrci6px+5BAm4yNUbbUkqJ8fkHjaNxG0vhO0cJXjlxs
R5nGiMXtD489153GA5LsAi802U8WYjxnId4OMj1K1b8p+b4QE/3hBDeaozuaisJeEOgeaCXiOlJg
s1/In8wxREclFk++MvFOQ7cUcrK3KLUIElfB+/iRH3IEdN5fEgqDByQDg83Xd7U/gaJCxV4+x5Zz
v24qkSZQdcSsCLgMVwX1Qg5kHqLYVPxi2SVsacy/QbLRM6mg5OQce+uVp0X7QU0lJ2i+46z2U95x
zyBk4BWoFg6PnT4vjKe/YaLV3ROlxTW/hX9LGrWWm3BEA62wREvJqMxoRQev9ke5OLB27YB3GZCn
7w/9Qa8PrNeWLhXu0jfZ+cyVZA7EGHQAJfBS5/17/cpi7IB+sI43mlguLsOdo+laFQmToRHOhpqf
/4xzfpnjTaLgmfVC5MFHioeeiYu8LBj7c9JZpBsNezdcqN2a6FHDBx+8GeQcHemhXWsCUDCC96ah
77smZdXbTh5wXMW06OtTtMIyDbUm9x/BjqtkacDdpKbqSKqQkk5InEkHu4hAr+W8Tb4R2dUTfWxK
3mbuiPHNnMOjaA7gjM+rWfYwLXUtuqVuRYG28nhcCJyYwHfXpMQfe0y9BGN25uOXTme44SUKnw9f
PLxnaXy5BrdTirHClOR+94E8v3X56AbxslbtJAeyth0KrVri/Pn06Csw5bZH0OpyXpUdO5U8lgfP
mNjt1YQmJnGmHuV//AmrQvp0ADHRDpg+PiPWYVn3NIRK8kuGNqbQ4gFj1JjkMwxwrKhEjHMZcwU6
hK5NpTY5s4oIBfsOsT7kiP6+v/z3ta3UM0sI98FCQR78yyVrV4/fq4pk+xm/cn1qEhNvTN1goukZ
0oz182LyPBZV/7MzQYUyWeQsHVDoWx5l8qnRAL88HGfJ1bpkuG5dAgXIqx4G1Iw/gCBXEUtGxCsq
3IQkTeUpdjfa80onTpfVtDljKRKn/QZzJoYdDRF3Bi+8YkEvr8Gpa57+2IkGvc+tIamKHzVCXEQL
XiXS6e0zv+r3k2AcVbUM9ypva/vOUaI0IZBFO+A7JvKMd65mE+UmCpUomDNbVJjZYUvMzz+QClIe
uXtQyvJ1Onz1cVwc8lDKK7VYElUhitEe0bSW2zkXuVIR7dz96xX9U95JtoYQgg0wYSiprB9LJ0Vt
quyLYSnAGLKCegwMjSLxkb8BHLVjmJlw8HKbHxeiqy4eDTsp5BDz72iLw78TOJH9oFRqs+dJ7C33
M+3ePBuJk5s5XV2J2USIDmGjTnN0ONz1hOnxA/WRZeLVv35hZh4jzpQhGTGFCsphtRBs23ftoduC
z/Te3pRb+Wu7+PyuFyVe8krpuepVJvXZ6BPPKOq8csrgxnROsWBfvquhYm0FAVox/Omz9SXL1m+o
Eyh9jlnWMWBppT4/7FesFhmuXDE1YJHvnYqvk7kW5rhNjf3YaSZcKcnjTelVM+DsJG6UB93oMYnY
DFfFKZB46Uv0ItVLXlLqxQ9MgbwMjxDfDWXS7z2sCD+Z+xOwjFtSxVDyuzrVFLtag1Pbqqk8aeSA
/n8CXF9X3RjG8Xo8tRlWvRiu9luGPAqeQcvmQ8m3ep7S8+SxQV8MLFtEVJVFz3nc6oTL+xN6weWj
bQT7DCexXLQFQLbu5zHn8RP+z5K8rejCCXCYKAvz0tRktBtZPgBcmqsXRwX+0qm9+uvAvXkVtWGb
D21faf4bSS2sNy53RDEnKiQTBvLJFNJbn1kJC2ZGcgPhXFteNRmcySGsBNUNoM+daE6BMszcfZpc
Y5145E2yCSU4dVjI5C8ngWYyT2PMbLiEPXbrhQumZQ+8i4XwkA1MyF2QdyiFkl4JYJv+7cPThNQg
Tk/5pRDj2X6ElmtdBu3Dixvv+7K+Jpt/G1J+wpyEqmApPVNdVoBDvknPzOVj+/PmQbQShGjNBVAh
XRi59JE8uxmsR76v2r87vd0oMd4HQQ44drRziKHlh+USy175Kd0R+2LtnEjO62wKwR1aUYgOOzK7
NwL5j88tw3NL08ReNyoBvndcSOnnfsKQMFA8hlbz0QoxGY92Q7fIYddeQd7IB8Uqv47nTXwMOJNT
awZdYGIgjts2elU++mcUp8ZYuBhT/47R4E32RRbGCC9IikO9rZeIICePQu8dn9N2gD8nPdZ8kJxY
aben9VRcaFCZiQB0XHvZikWCWLz/1DG5c2fy3hH3PL6Mg6zTuUvKRTHtR/KaDp6J31dEMynR0Dl9
MwKX/CqeM/RNj6iPwnC13LQIcp5iGle4MYnmOtWL6mgMgFWzySIJn4QE8Pt9U5pjvQl1WXwUKzJQ
fpTawz2LSaucS4m8Ak18JKOQlIyK3Z2hqisWBTU10QfYNQWsDJwUZkz/Z7HHt9smwyl7LoyAwj/B
f/iqgcvogMGafUQli/1og/mVZ89ftA3EZKV1x3ojVbDlqK7Y8sB1mHdUkZBe4SQpcG2kyLUFPPE+
LCzsKCtSo9FZrwjDF++eeOALKMmJVcNncEl0V2nGrazSEV7FyoBFiXTjUNyD9PrE7xWaNunEDPyR
vcnyqkv/9cz06V0kwwTOzytcC0n8fNpJfIo28ivQLPc4e0e6AtOmK34B/CP4/BbqodZhfLbdVFgc
bfRk37ciiXn488T2MRmxobrFCpU3VI0lPB/0XFQTY43925nYENaI+171Iv+DfghsKkyB5g4SbCJF
3jUMJUbsqlH+1TS3KnVgiAdpXwbfN8noQsSAp58OSipZfo8mjWUt3zNAD3yoTnr9zb1h1zJw92/T
VyLPVlXSrnS2xU1V/4JDlv0nXN6KZWNmZGH0E+iA4sCR4RaM82DYJksPKm1fe0EYofqL/EIfRHUS
4/f4R4Q6rhYh5YI9yMjchi0u3Tzcw3qy2InG0Z/MfT9qAy8TfvypVTkJAdzesF/YJkO972lZVO62
yKHnYiUk5pWCoWSSdOjP3cHPYWnatP1DKWdWQW3UBazDX9DEGRuq2CDuNswz3gI/FQYcU9oUCpNC
fihhTaNP1//eGg8fkAUHOyUSGBIpXDJ7cAKVY0bl/9UAk451/VlvUdTy0D+99T8zSTbsUaI/oOgS
bUj3/4zdORtcNDPr9/6TI5vAAA/5MRUTHi7aKdgZprnGzH9GyKrRSB4N1U1Q+JUgxEN2bkGWZCIj
LLBt7dow6xtgtBw1zt1tF7NuLTVs8k9AiWep3B8+mpvlCkDQkd9U03h4A7zBL6JOY1LVopICm9Kg
VjzdykkHUeMjijE4CFvDBAD8sfWUM4Ny8fQSBbYwlwOK68+aJ7XEJakKmIvYHWIiW6rWLZ44SHDO
DusrxxW+ZrOUVJLcsr1sr0gTJaFzW74z+XYxeZaV7S/7l4XDUZUxqDy7dXUKNxBlWlDj7vnn15Ao
TedwWV0IS1QBmSvATlxuv6gvlpb2AY+8z7qySJD/CNHPMWN0ljFO162ytju+5lDbNpU0eGNPUy2p
QS+FkJ3ZeQKCbsu47qqoc4pFLgazh0phmXm4N7jVSXmPBuzBrinU/guXYDOf2edbpj5H9NQ4AfKU
iwurvnUXToeirQ8JvNcJkTrw0SO90OMru9ueSBgJFvNySluWR7S6w0Z0pJMBytPJ95MXW2cSuQ4p
G/1Dh1IoxKdJq7xNAwgxe2uf1ZdnVHHTXLg6G+av04/6X2A/Cb/7rWcwilUgxvmPQOqj8BrzK5aR
kLMYe2Hzxb6IK5APTjY+/ttusiwpeJ2fHlpWDrEe7Q1qWUCF1PbTPcGmErMmczz2QU0MulBtPqBS
SAX76MJACsqWr0+dqGkYCChDuZOBkVgoUG4h5OyrlfXnUiPq5P8ZqgTqI3EkOaQpQAWONrgAwxw9
/BJx+vCK4qYqE4kRI2KWxeAcKocEa58y9P7pbEHUjqjctglwMSHgX7HxaC+UyvvjzMCQPzxCmcOA
d4Zss/Ui1lL62DBJGGULI3CjP1tGapOQThwPcj5FH6uGcyr6sj73dmP62VCLd9rJS1ypiPTmmJ7e
7Ou/EIVblygrvlWqj7GNrIUBtcDugKfr0i6khk9/C1cGkovOuCId1D7vYIGpB1BnxByMIdNB0GKP
Lv+rOBIplFs8Xcx+EvFjz2YHmE7ypbZd7qIyl4SOW+tVnVH6+vs+a5xzGc5UPX12C2PIPpauqBOG
DfBBL8Gmu+Hg5hogOp/FcE/Pa7on9KdW59l/02di7o5ypyX5VHeW1gQPSboBpXaIr93yPOTqViuK
IX+NFnTX6P+YOzbC2+xW6MC0lW3H0TCLa9gLCnrXzNfA81p0V/4vgNS603MzkhuJn2yVlERPgMLK
9ImtlWpGzVwUqbv9EdSIbJLgpORvbNlZ+RzaWBCfch+LnSj5LgPyx69hEFoqwNzJojio39GmtqCf
oEZSu6W8ZABf5oOimLVaE091c8O+xLp1iLAqO9F1NMksS5ca1EAr7dwVRDmTKpZ3Sk4EcnaBaYNV
RJNJg1tVoSv3jumUkt5A6PekpSJO6NpX0iNfzcYVW1hgVRvT87esuSyHBemoTTrH4e2mxNsdvl4d
TQGvks67gD5YAmI5tMOgzwuM0Yd96734I6Gm3f6OKRMQuLr6JXAmh7UZnERFdLRpe38FRzGauBSJ
wU04rxiTul/GwmeQpoQwIvOBNL2Hk03QiEqHqt0cN/HuEcohUgCrjYpvw4HSrPXcW1VTRehlQXKk
5oeJMUA8rBefya365R1JULjgHDHkHJQEInj8FRwRDucD1wqPo9Ejd3EVtoN/pTXqGHhyVN8Em+7X
RVGfHnaduOvXL8UtCOEn5Rlv928HExgoG1NLC25RjHa6CzkparBeOLjIXaF0Q4iwNjVQUIyU7gfY
OQpzlrqkaHJVSVlSujS4l5kzoKzC0Yt6aOW6fagwzOPinucVjUu+JRXUpUQc+IRVi3uE1F/jFX88
Xp78P2ELwS0JwZJUw6VrbLmpUPMAeBnusMu+iCnlAvqBniPAvoeo9zZYjieNt42Y4EWS41J3bcwD
LGWu48q8Uda6sJLddwY8+S6C9pyLmuNntjnSGLfsuXjci4ESMoEjDJaVkswmPZy7jTeSd/YFMzF1
GbcuE1wemS0X1NnAP8FGsWCm2JhaLdOpYnSaZn3BJBSgny9EL6TdrSwelL13r06LfeoZvze5S5Qv
dvGbnx685o/EePQDERhgYx9Dgfk7vsCFzNLb6O4vnF0KfJXh/a/6B9rapO5jXXOt8mAh9gEQkkvG
MOXM+AdRKt5wNDHsaJb3Tc3r5f6cUfRLHzOBMSzgf5kymgB3VPj6kC0JImtOC5Assv1D3bvGBAgJ
utFc0NHZ8zZdUmNcBMS04HPYRwWh21vjA1y83m15a2Zbis8F3esmzFbjqJNVApRNKKuHPqFmfW1O
F2bFuu2oYsuGaPu2d2/hLBtwgp3tvHEyj1FOOqa25x8DRe75d4kMDcxdpMWlTvQq7B8KkBw/j1Y4
5tlxzGqjA7KqTaTpMZyaylYeb2hn/gybpjxVMBreGCedI213HdtnTrOnecPmjVsSYpoSAV/Szjh2
fYmrkSFw3et/OIkz6H5dvbUxsJQq3JTAstSGw7T0rz04XkzTpPH5IPb77l2z9LfSBcRMOcUiGXXs
awCUxHCoUPtSn8XtDoyIt+tDC8vftvydZYb06Zls8k/XA9ROUFHua7WKjTRBY0Xah5gfE4eM18aR
2etyANCkK/bDfAONs7Z9AOZCDl2rRNYAhf2Y6KKTbgTN2UsAaUUvRIVdtzM0f/HVYJSXErXPVIt0
ds79b02xUMipo35cRtzsRLIRbYzwzjrWUalqE423IdeMieb3y9oJ1PNK9qIjBS7prR4WBal3Ufox
gbrCRX28rdSF7l4JiaumKvfZu+bYk5NByFa0kEVnVJChKjGp3fus5/jqXHGyarbxKQfcCEqZy3zt
PXhS64G+qG7P0axSKfYnQNsupidvo3opE8Fc9iOGtPV9ETvu7ifrGU259kmDPrMBFJwmdGmsnMr3
yUc2DSiZwH3K8lkWKZ0YWaM7+WSJe26UJtM5SZ3i7lnEnoONh8NLzML3zH+OrZV7RdfQazhdFBPp
SwF/32oLWpSmZ9m+DVCw9H9PohQcjQuQ+KgvhhJAbmzPmC7K5DxkwOri5C0CRp5XhRynGvRKXyjH
D5uEnxbS/Lk/97xbDitgyQCyTWl50G68vTppAtVel+gVv6gkmc4csVOhsNTvOJRe1uCElbQ10DG0
cMiLskTYrvaw47cCsVijPzFKR4BGK09C1q5E+7OcZ2GgjA7f067PArN18wcPnI9tpDzgy0G+o/D3
Ja6kK/FcX8J5ty1sB5F3zflSAml2gffLzWoyxHyOXRl9vwMo/eh9hRKY8uK6EPf+nzGtP+RH9ONw
UguFSB0YJasUH1IiH6aVps8lIFmSN9jh9p8JV37azZu4MD2Z8MY7w1vGmtoK8ueo1adlLT8kk0cC
teReaRTOUxJ7mAysssLj3vjwQNnpYhVLrSCp00sICspvd4PKMLzRYdG9DV4QG3+f9a1w0Av/ydTF
gzN95jibrmtm7y7RV5OF+RNqJQAfSxIWxMOWFgaYLZg99fmBb0r8brZSPy+0JZycjPkFGhpnC7I3
8o4YnTNX6+v+9KxrQlh6RBQm19kVIp4Ucg0Gq5K5aFVhh5sWgtUzBn52E7LyzTt2mHU/Gwi+5nbD
6+y2C0zxAmZbBd6jsV94oNT6gZ4iaZC75aeTJW2uKYtCkGvgvvk7cYqcraUEMYS/tg0LFrh9d8JV
ByluqiyDjH4hV0fbxDptKA8cZAkuxliXgliGyE9BqER/SGpIZseYFYF851A8G7P+J041bELTCPHa
sG4w2fhpKL0YJs4xYfsFHtbUbljzbYYZriA8dztNc4aXTNMdgoDanjAZT4DfPlkwvXFKy1F86zsO
RrHFItPF+r5h0nFgbmwNK1bVeXPY6vYVf2J7u0KBih18TKmtbQL8o9nfoVb/3AiTlStDa9yAkuAS
RXcIQzHDLphDpCyO5VHnLJP5vbTynhDumCSClP8A/k9Xhx5GKzkMJ4qVgDks9geWBjkZAjsy34AK
es/FVFjyhTNXg+gTy5cvlGdNuxWCTNQJt83Am+CR3qSJJyxu92AL+mtEa4qV7fK6NaxqwdMt+5+w
YkBdwRl7Il9HXELhZeJ3gU7CyXyEL8dz+54qbDHFQDafdg6gyrVAp/rF5euod37nu0PsiKHUUYWZ
NaDaUYHbHfi8Y6y8wpDk8JGurEu8qu3qqyVtIq2rSvBJEHzMc0mi8tPh+XdFRur13V622molGCwf
T1xjzJMiEAm8jqMS5iFoCHkkPZvdXICvq2yJeDkIkonilUzgrAa4YB7g/jM++SsY8d1vi1ooke2K
4KKICu1rhY/c7xpY01tvhoKLlP3qGV6ER6SuOVT5LDcXBYc08Cq7fUbATigUoFQxZdAdOu/AhnZI
pQQY60Ybdbhb7/qQuDoxUlDRDBHZ9wp04mOadjw4rVHEzAVGeQBVmZtKgzn3/1WY5wmADG5QptGn
1fpMCWeJFqeVHne3/H3ftiD23YAm62sEUmuRzEubv2x0TjoHLn7tFFdjhaRlnLB/yepVZehLs/4C
ktxaEvGZw3WuBW7aaSSwArzBJUFcoeOFWIoozm61m69dpNo/tC0i27cnMGUVMCyHlo8u0yT5nuvF
lI2OUpGNEZlIm0xaYS2h6EbWtmvojN5/Jyi0sPGLCGM1cT9m9pnqYqc/9aqmv+CposJUVEsYVlVf
H1scGAnMTkUOW8Hk3yX5UDoGQsbeLjco5MdA8Vdp4DkA/RBMgKKevcZFTrKigRMRMTgv1NXjCJIj
6IWGEG0LZJRoHNSCbDsQ3fJx3/ZLTDHIAQmOG2RzrWR7OqQq64WZIe3iKA9hdRBIdWNGneNckVep
FXtBegkYhOElRKuqPKwizMZP51qGDXkpgihqoMx9oEDM2SXZSQ2WvPKZpTowip3/DgN8DkwCYX1b
XsabRCDEmUDPaJNDjy0eeUCqVYZpfvlTnUqJr7jvp2gF4DpPfxnK9TKzKAmnfggSh/apN80JWhmM
mggw71F0tDN4rmXPLEB2oZ7Ixwl1joz/06kn81X1i/ZDqlLGq2g/7P58I6o4CXJ3qMu7nn5WPIUw
3g25xVmgJ3998ECIo2h+WBAOocNz8GUMTSfwp99VzhgHPKoFFL9ldBiEHFDkeqo25lmRisESMgAa
N9T43gzyyx35af3ejCzdzmSn7i0cYkebDoTUuLqvqFhXMfRser64Cn9y9/qmHP6YTdPUWVIjxR6c
nETP2u+2+93UEelvg4ZHhCiKDIbMOqT/SPM8QmcKmvyM+Bqaqg4U7PooTGj/JLpWBJyPofaWee83
beeiK+FhREBBvp7Cbt+kVeGjLK7WkcTEXRaYB3eSoflSUbb/xFZbwHHsEYc8kHP+yUIGhGuRD/3j
c06Xxq5ol/DxZ/JA9YJyLhjzyzTYVKth+i9up6tnfc1VWUmCzUzfNJXOkZvKKitocx4+zewTvHO8
QW3Kk5/82ZZSp/ElG7+SKKRnTglD2FgFgat8og4NgRaC8t/+a3AO6tlEH/XDpvV8UMOR/QM/yp2B
f1+wfE6tII5R6e+aGe+xgm53/Gxb2upKQO2eySvtO3L2BazFJ9e6e/VjJlfHAYdFFsmyyH4KYrSV
K9dVZkCOtww66CqMN3zcIB7OD7VlTZ/nHZv+7snqlwuUlz1hedJ6No39Kljl32ioG8O9VC96djnz
AB6T4tMNDtTVrvQFA6/GGrC1iw5CGV6QFf5KA7lDjAi69p3MSB4UQZFn74wyY3Op01HAf3gYei7g
i+4FSFZ41RVST/7kWABPV4nAI747vic9NYRmglfijOKLnwUuFVPnUgCg+m6D1CBhBhWBk9Gx2oVP
O9X/3nCJZXeNhcaD80xGvw1nP6NvOcyy949TzsO9AJAHlp+RalX5OmJbZM24lEFsfsNtGZ3zmRIy
cV7Ccf/tyi/9MGjKxqdsu6uUIUNd7IvkixjTfi33V2CkfzpMeWfq65CjMRBLLa6pypqzf07wWCBH
6ZJTvx0063C7SVo210JS/no9SQkgu+dbM0DizPYA4RmB2SeXpnwoNox1WHWju8lXvv4rljqawKjm
y6COgu6Vi7PrRfcQwkuWBlYXav//WQ1Kaylwcz7hSQ63mj2mnlxzYewhSk9Z7WHB4yDEwCBwwyxk
uRce7L9NystaIUyPgVBjh9SPDcODB5pGxJjbOLiExZ7i0g9N5k33k92lXgTvzOswcRhYudFKsh21
4VkF4KxrwzJxEoxhmK8U4ejQ0UhMBM742yz3Uf4b9U+2h1thPUlTdcwC4EkmMQmkJlPeRm9l2EJc
GWr7C2uXLpsOtRnJvd0eKvD8v1hgiEwnfrbQJMUIcJAKZMPOt1SyNWKwH7f7gPdtLoXCOy95VzFa
l8AknR+UJpt8AI98Ygr4cyWgTNcpmPr5f3cr8tLPWstjQVMqhBFoRfCM6BwGgLC0lxISNlCXIJzr
oYis6E1jVWczO2Gd8dD1XruT5aaDissjtO3R9/x8IaJVbn/TphZTabjp6H11czBG7+A629u13m8X
9uD4qd5rxFshFdGNvUO/QB+I3mXjTXA2v81SJw8Nwb76bRkEBA89mOD1NF783yY8TnDscWNeOpmp
TwDg1067Zxu+MFLjMC6Tzhzj1vCWD5y5mAEnfmIqi22MkAosR5pGWmVxBUlvYWxScSjE+g/cObKM
ntICqgD4+nb8WiEjJH6f2eTX60u/bQ8sKO2yTgb+VSeXBbk1Nr+Z1lHvir+Om/fg5kJTXqt/R+ST
GilwUmm9JFiAe1wotUxrR2cDfLP3jhAgUqJ8uSvjmILRj0aDkR04kvl19cRynI80X8zzTbKM1rwB
5Le4INVi31w5iDeTBFCPFMPisRIffs86ZTKQFsafdjdEJkHwj5ZRb+u1L/7D3hOnoecboyArVGAP
CRxyI7IW/yNy/y236dt77VUKSK1eJGgQpB+sYNjeXVB0udc4jouSX6bXAcQzNhqu8NumzqR2CCME
4nNLmD7ZsRbtDvt8qmNcLm2B/6th0oyc0+h8FoVfwz1DDY8BNTP4sX2XCBNdn3n4xpjrf9bXcB4v
nckjDAXIHvausPKkgImavOebAx8thBPVweLFMg70dXfY9uB+eELdqPVN4/bn5xC/n9h+xbUXg/EK
jdUsLLmYKiLUoetpX8Xqsog1VYtnXwkvu9VVsigOHgr63HENunRzWLmBcdR90fKcL7fBKhBrlgho
S8I2NE8welrYavGfcHjiBQojBnbTTjPoiPE8rpwm7MNRCd3ZalgbegWoAjdvrlTZbPXaHtKgL2VR
ehGadIz9LFzvWYiSoWF05NLTFlU3jh4exd2DbCS+ppkjrz5gS9lJu06Ac8cdfjTVOiSenC4LZijG
QokAlnl2bujreVkSPgWH2BnzNi0dwiA1wAaEkrI4iRDkwqhxz2luAiSY196qbpO8dx0PFBIewuWL
ugljPLIZ9KDfutaKpK38dnqLc49CFVzv5Vpo+87Yb/EeoCz8bCSb5ERa24kMxr6AUHXI2bDnYkST
qrQJbXYhU5kCWJRqYe50OQZ8lzbMrmLV6F4RUXFy3Y03ExVsx5gcQANrqGLMd7O/mqOlO56X16W3
RPfVPPp6JMTIVhA7FhtrclFpH7NTThl9fEK38bwIG0QC6FyenCZR3vuv29bMPCo1/j4APtOGzRmL
xICprwQculOhOlibnfqbkAemLJjAg3deGL39NEjJCV7tg2NbOcyw+MKU8eFXCy5mKJlS8YHvj0IN
feLMc9RK2U5muWXDSBr+/eOLm/wDATGp2AKJygRRUD3m8yc5q/tAi+1y8xR9ZYB0HWMMrtBKcj9B
j0YpPd4iZGNG1b6HOlvdcoHGb0XzOLKcJIJeL1Yr7tGpbA5oXMCEW0fNMlejmx7ijBoyR5MRvtKW
IExECqHz1Xu0dId/PulBrpksrWwJa4veTT0TYUpFjAyg5mzv5K0BuHl8godZh84PzxFLIWkYczWW
dx7yBElP+jvwHN7EVQ5rz2+18TBW6HBg34r8Lj+6RPC1gzOSpeOCMqZPYyf1izopHjBe1IgiZ4Ro
/wybIBm+GXRnLLSvnFjtTrl3qOKSmdZykfGWw7BfnnWi975gMSj9SNC8Kger5tgmNu2K+yuSChrB
Pkxazbzzu+sx98AXdX6AreCAF4A/ncgCJ7jh0tyLl/NIP7wURpuVow1bEjKpQiQZPCvqPquJ/K3w
rr5orgDiYRjqbQmmtVTpCtDcgChKgQVdxH4u3o82W9u3ybFTE7ekIDyiqZ6p20Vnxtjwr1ttaI6H
+1zr4yJ/Xf9B/5xmFk5Lz+ZtW4AWeb1EEDqATcTwRoXFt2slhVKn9rmqNUQMmfCO7q+88we7+4kX
MpoE0IIDQRZsOlCXpWY0UxDquMpKn4npSYZPDwUvcWybE1A7BYBP8XuEp2IS1gCAR2+vfowhFq/P
rhrHG/OHHBUBmusU/3dELxDXvq6Q161jNCCdQKu1IC/8NThvHBIPmDzjVnTfsdgEzWQtLHl2a4r+
QphiSXeRyIgnTc8kEg780wxvh7DEKlpv0RW5fPYw4TRbshMM3ZI4qGD4/dMiCl7EJqywBxKtIF69
Q+CP+gprLxzwz9685R1zn6u0yC3uIU1+DH/sBVrBGsWS93KgFTVh9CZaVbSwa/Ktp0wqnWz3IbXm
UM6f7zd1zti3xSeDM+/EvkMPoXVh7HkHv5B73pJUvxMRespBW/Ylc7Q1EQqmMMW5VW8XdS22Ofin
wWySFsbK74BuGgRj09E84/W1Oj+BSYMCj3cJpXJIjvYNdlVaxrhDxomTOU18jDZOczwTbtGKxAow
x5Fn3SilGiOVvLIyTlCu1KwnBQsGnWum14Dl8Z5ZYH/WMYqHWZgv15EX8YFdpBRnVFhmMKgcBJg1
GZ1eJ/iGHSoR90EhYr7Idn0BcnAVglrVzqymcTvx/dZT5SgQkA0bZy8ZybUm1Y/ZRvYLp0XxvxXX
dihwejPfKWvhb7rYfdKbpHoDkkXEhw6VGxjfY+ZNokUQZ0bdmv2jnaLkqsFZmc5+W+6fsSlOLwwI
bbWj609Hezr9rH/LxpPOeAYqthRDPGmoebdCmpApVaZgWhaQEd+JBE6A9oEmtAKvQ/0c6lUx0/4n
ltHSGH+O1C2upbKTa0BKJyJwM1tdGUAUovNMBEHS3Eppqnf4f6cW42z7zI++c3iNTR44bARpALih
iIU3e+TDfQ5ORSMzfZO26mn6kdCYIPACWIprE0C+V1C3BAb/aPlTrzxREfH4rR+xwt+liu3xOoKf
UGgaNCQa04nVlMm86Pa8qfTXbLasnrTVKWrpw6OODqXgLgb4LkZSI+NmALGmlpaUhrnllQoTTvqm
BSvjKylMYr2oE9sFvzyURkJls/ss6sjMW6Tk7hMT1fZ2r9sBuuSJie1LMliPU4zlap0C4rbWPIPi
erbImguOPkdg6wLp1O39ZlutqtiKnvFh7Pn7lohiPGR0l1A55bs6j1s29X7At5+ddZl8b19Bd6YS
9sOAYpTJ5QrvOVWS0zI/VluVFW5O5tCElcqDReUobKUFjTQ9vQnRKuxk6meFMQNUjh/PPsMpmsEC
Mh6u5yoasWWF3ypPw5ENgMdJZmM0LBKXEwZ7lBhi/3v+0vQU0WjE/hXvwSSsVq43r5yP1WArbXYw
Gqnzs/MMtK/8yPivPzupAT4EkH3BcebbhoYblxNu6PbsgS+yn5Wmy6B/ImxfPMMGevl2vfuH7PNV
mKnwDzI26EKbfMeqyOq7D3mcdrBQbx3cKv3ol/3lXU5iA/F3aG8LlyBLK/lx1NN4ynGNuMyZvukU
K0Q7SOukTo5W/TXOMcL1pFZqbolARiyMnKlDeJ1xPi0nFFWDNuxiJdf7niqOQBYhuxGP7kVRSNZF
oQXfxcmrKT1v2ELb1FEV3pPgKSsR7aH3cH4NMS25yqx8zzIU9zvaTiOha72+IwDzj2PpUFxRicbg
vRBEjTO4JNbZcn40efdYjcqu84tO3rS8yPCAgcgKaDuvPx/DAHOEvmRtSzrTkE4j8+S6yCrTROqd
6aLzS5H3C7p8yT48Dch3YE5NzlbGfuqLiF3mrVxghs6hUrmqa3MbGK2W8Kt15juwnoF3KesK3cmL
tiTtCWnAi+o6+ujPCRsoYEkbrJOmt4ji7cfruzflUPNeg2OOrezGLjBFgx6666TabLYmsqoQSzr0
VGKBS6GqqrVBUcKjxT98E4p/CWxUobwxOXSfySI4IP6Z0oYPtLV5qKQCwH2zdPbFb7x6W+2S33mK
wawSq58e2FCEdvpRvlCx509QnzRXSmg5Tmwq1gzhHoP6N9rt3JYdeWFXXfN4LxihS9vAX50bQq7Q
hXOlqG8HVcJpQn4a/ywotYpO2iwXiYMn3p3ijWYwlTfYcNoollaYtWszMi9RNzb9gD8xwhRw3lvy
4qekNyiJVl7L9TltXXpsq5XSeHZ1AWREwJ/vifYrUchnLKZ5JNEAD9Cz2Ts12jxgHBvW0uXx8Qq4
xaDsZc0rQwFNNGE5CTvqL0h3GIWFm4z4ZvU8bLpOjoNkFS0BxFLtXiQzCEHRT3w1VTJy8snuPSaR
7nkOC4t1ihZxiUEEww2W29UYX2g1FFoL2d8LYTCjtBs2ip9/WxetWXvoz73KC3b2H81yYJU0kIEV
9ZLO6v2+OuuXDbKFEhAoz051unolidIeIR2/Ppsp3AnjgMxKOGSsBZYfJnqtetm3OLTxnGB8dNQ+
GMFTg1mMTsCoCNtQQxVyIkAElvDI7l9s98GZguI/bug7XDEKgJ2e06rr420SZBDjlNyO4rwAu38e
owpmgv7qG8DLnvXSLbFZyp5zXoSO+PzDrbVAKVkyaovYyv6FlPSxlBgHokXhWIZ8IqolgJK4lrXG
OAkvGBgWeiZa2ch3Ssb4X1z+qC/AhIw9Nsn4z5xmq60Ce2JpmMq6K3ZJSyGLzfqRvP05cp66oK4R
C1Mt93YDoFQfj0KAX+7cT1XUZfXvsNlAr/ypmkZ/KiiDugd5a8FQSllRaqXLoP8FOc8cpjRCxTCS
QX+AUOavi2aSzf4+OdRKuY845LzI54nM2AD3h1hvjJrt/Qp4nzi3i+n6c5r57MawonQ4QogGUPrI
YqWvzqN2ZciqkNXUtzl2HoGqMeDZ4vCn+aA2QBlzS2yVWs4TphF0R+OIH6dIpk7eK2rq4A5wG4+f
EBSwVmJrlTPV/qTKVZCeknvMsT/FKbJGIvROtRQ67NTybd+8pI+L3A1m2kc6ZBWQ7DbjiZsPQijy
wBrC4A4725F+OHIwSScdYmgkpNU0kNhcjP5Stcsp88tDp1MrJIMOgc3ca/uglx2RTZiUnW9znp5i
rW37AC+jiJl/qAOVOND8orXaCRBpwknjIwHA2a/OBzOk7ispLjo31+IFpvDo61JNNMXFwCPu+TzY
TSErceEgM+2xyo3WEau4g/s9li+iTyR8HBEFfPlQm8tCPDslUFp+9UQjY54FCRmNsFdREvwVBDZz
SXOSQgTppg6omRx8ZhpohNGryfGvJGuOZshc9ftUmkSoWNcKXTaN/FpbOqqCYxQCIxW5UO2TgJYq
NFJzuCx83JXMVIS1AEtadR2T2py2y6PF+HX3zafkK8UQoj+lkyrIikWN7Re8Hud18eZNRDbTQKjk
GYO2PEkt/42e1IMNtp67FZFyy4UOYnVgaUUWDdVYMIkDR6SS7+IlU9/8IYZ+wnxeg97wthBy4VOt
pNbPU95tjlEv1DLqo+czdchWbMYbiF4axNEIwE5CN4qs+FKGFvhpye/rDZITYce6FNP5Wg0WYESS
cMG81+hxONT4pNM1ywhp/+tXJessLitDUjEnKqp/XP1/tDXIGRNSQQNvdHqeJde60w6+ozwCDT6V
j3U2I29BxW2MqSpVoeoBJGXoq73B0bSSki47/g4W+8lNCWbiyDhEq3ePrxtouNMHv4IuIkMC4pG9
NKyZBCIiyFrt3Mv3UnZPe2N6KZ34aDn3M/ZUPCppF8eqnli6TK595lz74flLmRNmkBz/ZzVx9YXR
rh8COmolvXrNjnxbhKnAIIb+lpkyqak9RvXJBjaL1rbJ1EyD5W/vhUFTRsuxZgDbY42B8GJRjVgn
1SC3NjYiUo/Y96yOgxxNHiT9urEhFTmEsaGhmzsbNJBOwLSaRw8H8TX0ZBDj7vOXWcQYL37J07gc
9lpWQgF8+2vto6A+8mQNWZOr25SfE23MgjGLEotr63Jr1yRR9u1FuH5hlqcAt4WUmVtM4I+4S/PE
zTbuTshi/Rgipg/fSLBUJpdAAsHYNvzF2q1I0Ycj4fbrX+kJCp10PDEhGCl60+jthW93o1mYxhku
ahk0zyJFRW42ocnMVG8/JiDHlKOx5hrqd19lyB5BDRJtTQrcYQVuGWjd5XR/zhx/lWNOj2EwX7EL
e1YnF6RuYhz1XsMtrQctkrH1fr5zQhWcJ8loyVpU9+jIUfb7kADLbfMLMf1HyYCjwPJGvNSZ4ATG
aIhUtWXnpb39evrajUXP7ZXd5IKZ5/d5nJ2tHScF1Zd4AzDbVdP/mZlntaJ4pVr6Av+7LSu1mkjq
jPFIyQPDoJG8AXh02SG6Go7MNHw4Jwo0AOGdcFbJ2vn24Kx2uyBIa7XjTpkjNamW7ZKy7+SScyPR
zgqr3prY8S9XijXve6qoSI8eldqejSt2woDBhIev9S7rARSyyyduK50+mcLD1dWuYN4TGZvSx3Lz
rlG6lq3Pr5AAXRKsaHw1SYRncbh4mePqxQUzwI0nCKjTo0JU/b+cr04xyoXafEglWTeiZ79VxUTn
CyrGiakKK94NXACxo3Tq7ZUrEOqxeo4k6EoYz6VyNN+YU8sP9E0K14QKSQC2Sl1NKXySaAnmRXSq
K18z6CetrGZkf4C6l/tC1jAuj4FD0N2EQ72qImPoPZTJBwbLQl9+lKTwOfzY4QLCgk/YIX/TqmfO
rZWrnUyvnfYxLPmE+SfMhTDYxP2aQwIOZXwUbFdRc1BkElXOVT3uFpYNJNm4hd6yqk+ylr1CSLm+
X9ycOMmhbQxbPjHOAaDYAMSRw0qyE7vbt+dTYgOdAAaJlnLQJdJUvaY7h5qirU29ViK2h4zEQ+i2
w0leSQjNJBVhmViFOXjFd/kaOfXyUuXWTbVp8MoMpzBzGKMANuGQcE22vGQiSlc1jRndAElti9Jp
4PXwyEri2g3foyT31xmf0gUIYE3yQ5+BR3EZaVkoNfE8uidBh0pDa64q+0VnPRVHpEQ0wVbApI1O
j3qT10IUpG8WbMZcImVmvzlH+a1j6DYcWyZPUJ9jsRXnA98jBIASWeSbZdULzV0JAOPOPMoAXhGB
gkFmqWSHTVGj73Z8qyCTWF6XAUb3RQgzR0/NMIQn0Js46NXV8N1qzITI/TS0wTkRfKgZfyhLDpKL
tkkymJIKurLyxNAMa8IIq58ANHSMvS25JcxEK8PByKz/UH36RM8Dp7FeHspE4Lks4ARboZbElVvL
GMGHCZTwWpwv4s+pqZt6ZHVXFASxZTxe3cbxUUVW9SU3LGqD0Z3TfOumySEIVa833dOpoyvmcC1p
R9ddvdH+YsX8umlWDh/SiOJIU4YKOFBNYPcS4vqtDx4uggY8xD8smCXuKYa71x6zN3Ez5wv3IFEn
EkMRBo8s3sXRlm6ahdaI8SJ9JZng0TzmmIpAlYlLLNPhiP5Y8/D6Qm8590CwrZpHbgYFucsDJnvl
/rMaOTzTEr+DtpuiQ8YrRwy2hf93EJ8si/AYbw6E/k2hjMRqRMwHWXTI+DJE3rjc6Aklld8xczeI
zT+lS+HzOeUF1aZK0eAud0LKWPacUhRG7av/2clVozTMkd5B4/k6QdFJ7xKx9fyhDdMN8+jEOkag
lzbxDaQqHYjEnBk6G0Qb83J1LDbl1xzGSQccKouyTCS6gyvB21XeWOyeHdVZqsDwzIehAfOV42yc
kDfbitWQ5iKBwmG0Lu6e5LeSBVri4fFvcdsXBr4/3Q3mg70XwCRChgYplDZgMuDJRZVbUvTbNdYI
isJyc1lV6K5MjOxddUTtMS9P3gaHPwyDDqZd+CKaxm3Cg0wZM/ZNSaD7yovhbsasipZS8F6CRm8p
yI1KbGTZzYoczrnXPPJNwTjHwPbjhgHab7j/MHfEs+8ehjfrZtvOLwXNzEP+Ep+8P1jfOfHhF39U
NGhhwNE3fxKyXc5Ghp22pEvGQqgnn1LSaacJ4Bpd6xy1GORx/56yifj6BwRHlOW9HoGTmI9eDicQ
qJsb2SXyfOYOzlV6cjPjPOPG4sqX0WXQRMuvO3+Hvc01fuE2u5TWMTAXz1HJ5OC4ArTIEPBzn91v
kI3lNUdp5CKBQ3yYcnHZg0G9RSPcMLJjWaeFWkmpXQRiNFvVagQh4qsu2f3G9Bh4OJArfu0YKlm5
TeQmmqHoCFX3IXbRoLIJOOaYsTsqD2UbXgOK1+uTSEPX0QDo0zQQbBCSHBKp7HlBot5Y96tDBotM
/hg0zrCq6nmcXzSkxBrlHuR15VGxqSrc3X9Ic0OuJMRetTKnFFkomorl9Y0AquZKFvwoUlkJpGfZ
UGhtqc94ys1voahBqKUOBOg+YL0gEPQtsPOVEXMvWUj4vq2AVN4EhPBqtsxOO7XZCK826pGugUnL
5UhXeQ8irJSgCZw74xfbgmG5LnG5Dp+ZUQmFGWrxvDM4+BGza9pFQFGkPMOHwMAU7e5zIfTuIUnJ
1LPzWsb8JRP1IhLW2OHthQBgw7Ry6hu23NDzDO9dN/ISPVDPaTwVLoVuRNJJGG72cSvWCCQ3O/GL
QFzX8cq608bz3EtiogUlOX6+HBalC101mmd2sRbNwg+CBt4aT6JyJVP52r8SYVc7Xk6cDAplgroq
AJeNiGU+0o8WIdcDVAPPoYf6vVkBkdbzFVjyZpszHrHKk5q4qvuEeNJv7FrXo96QUSyjB0gt/EHN
6OK1SsCwi+KyP/m+45JaTuU2pkCVTjeSUDe0wYOYQYqMgpIpV3sS2x9tTixZG+z7wF3YowP7QvKR
PiUS+FJ9drIJjNeS9Dh2jrDVFl4kcAzlO2YdWhKvuSjJPS5I++K6yD88PrHMPwI0JUazhowhRSD6
f25cdZJTp1wOzj1p7cUGrpqwOa3+StcWGfYGVVc6+3vLlEl/xrKv7ymF8kb/Hhl0AZCjDgfhLXxf
msQjSp71myQgWmUr/5QRXVCPLFytGxm6iHfbcjJ53ecKan5wecmYm2sy83IIYrLgSGhMAqPYtgVH
S/QtEI8N5q44NncqzXV41CqYJ7zCHOjS28YJmjtLZ3FUL1B81nfzkQHEBO75BnLZPxmikKkZutv1
lCk+u/niQN9shzCyrt50yBSUZ/lHWcd4hFfQiSNusQmMf/LnU3ULvi78az14T/uYcLi3tlsRfhcq
gpi1HWmrQQNC5DtfPWsavFxjCNyFLiN/a53kNpDDzX4ScwLVoFaVYGu0uIosJ5J26fWOqHeajX0m
QoAaHrn4eRI/OxYx87d9PVZDsyVDP1Yg66Fh1OiA0pLVsAzLb0HNZ5Slnh1TXE0mBrHXYWGaF5nZ
etwiwjhI0IB1RqxbeCqjx4G4PY6bPEwLuIMVp0kFRPidFqufLdChkwDaCBA4gAIYDRXQxe3xq1wf
qBS1wpEYSSYOuMKwr22DRljskKoxeuuucsGlQ7PdS4zR5VpnsVa7P/VAaaASmFaNU/XZP7KBNosI
krVmG3NuPxkEIqROF8NOnAmJ3ydePp67W1vfWMREwD+tWQQ99PI+vnpKnze8uHf4g9uMhDj6jSGR
eRZq5PEgzqKeF88x0d6AYwc0rtDzFwerdXIw4fI1n9Jlq/qnvz/wYNfoA9Bm+MX+qKu6o489Z7fK
EmWPu2mAM81l4GF//NFi0jihrIjEHei7gnmyGosiDPp4V5i2ffkxJA/lHGwFylEWjpqLp9IpsnZA
gLBsw01msH0ujCqBAsdaQv8fMbYLakIDJykZ3DdTfJOH57tQKHUfDhe5DGNo+lagr6FY7QrrZucR
9qJKLXxBnis/jDWd988/mXEcS5fWfoaT01+BtiEmkWYe8aw5RPhM0S1AC3FOu1YIbNAlgKAEEzyB
GqAvqigc1VKL4KvISGzcDZtOjOTGiRONn/IkjprHoV2t7n2c3bHi0IGpV0EvLCRi4R8mmnYeC+Kz
o8VUFR/Mni7GiSnQbRcQ9Fx+QFWEEETHnYf9nyaWDNcMB2Mc++ZELmyxeOfxClWwDbXrczp+fo7y
rMgp8po4Q1s+3tDdgMVARBpgJip/WXOHM66NokeaZ+PaXEVeMw24RQZSjOJdUSKaDHCBF1l8PAap
EXvVkJA9ksQgiG1oCHb3E83zhcUdcKygeJV4EEq3i3rjEIHphfrdQ4S9J8wr9D1Y8b2Nq/+R0Mxe
h5LN+OKSTV5AQUIIwsaow3h/JwCDmgIuRY1r3f8tjS1oVGnZsDfnoImRNKptmOZ3Dbue3c4ty/5a
URUjaME5hBwY3rJ2zVcgfZqX8+uASLerbYaK+oOzWDPAFSPi55EZFRd4rB1ty/Dt0fts27C6pvEg
3ngjKs82HA9iX/LYtTrGtdQaOyZdcBbe4GJZgPQlDiHPqkzWoREfVCbTENLwCuS5ffj7NdCxHWOF
dTtWmx7ON4pXmJH97xiYN9PaO24bIoYj/v3vNveAByZwDhExd/wf13R1soaO07FIHMranUvjEIm4
PhQX+KK+aXUHYx+d8niczyZUPdJzgx0Xt4g/pkb/Cmo6JGR6VJ/IjFouJiZ5dqRytCd/DKof3+A0
SK3I33sZA7AUB0IO1EL5YgU7+vAUaqIw0lvxZkZlNL0eulX0NTLGneVk+FFuCOzHg8R73uXWRXfp
rooFfcYh9F98S0tUk95Q/yZXCPYJIpRaOUMWaE/S8DAGWwzeTQ6z2yo00jgUt+EOsPuPTZroQ4/d
0ARaOllhjMqhpz/36ZTySSg1/neXTaQknypQ+MEApjCxNElKL93cKZd6dnHRwhvgcq9i6V+Co1Kc
i5tf7VrusYDrqdaE92HbzcP8m5zgVUw4YgGdnD6uGJWM1LNwR/oux9j8mld3K0GRuwgquIdStrxz
Mkb1BiKzTRnS90DW/SOqWM1vA3Ea/DGR0nArW+BC8HIDOGZX6aM1V81S4mf7N6e6HxJK0iGeoWoI
BA5xLH1dlTHh2MF0bJKzN7hxZM2jVKubhUxH5J5Wa8G/oAuhaYbnqUZ0mexkWErVXwMl5UDgNrwm
pBThwzWM3DhTGLt6jdw/KaS5QqCQfutHEwXExkZF+hOpLsbxkU2mDZXW+OQW3jHvsbNmIZQs8udd
9ISTeQrlrfgco1bm4CeJR4u1lvy17jSpadfjAxQbQjJVGy2fXhB15ulskOsYCX4TRZo2vH+ZR8B+
fcHKuTaNP7XeJUsnsZyy+GbedWKcAHJFEaEpqiYtq/nOIR86QloGm0nugdwxG5JLksrnV/3DOY1q
eOoAV+xXDp/MjWn9qoe0Zaeig5orGcrefy3y/MjXZ2t65QzOml2RA6riT1ezMnNkjdKW1dJXz/1f
ZUakNl86BlKJud7rEvH+TyVeKq3cYy6K2JrUMAFAeSXBvsJSpdhenHx39S/cRljzdf5TU/20oTom
FIyyLI2TFgPxJYY0M4FdP91+ifnoK6dzUVlkd7fDebXikKFev9GvhJDfEm9Fz1wVw8m0Sx8Bsm3S
B88Td8V1Pj/ii1WSigIAqAWej5ddzSXPe04eeNxYc5wyC/wr1iecOI/wmWvZctUyV2n6aCNfnptF
eml5ArxO8F1lNN77PymX6/d3sM2QgfCpE8qcJP1ndCOplwCUU2sEstBpn9xHZwe0GfhHBBOeos+1
aUFKZufrXhUobc80O2KLP/hNAz0yjrvcgFDe/Yp0AvRmm8060esmF4L4gjPX7Q+/6RF0/sLrDCqM
xeVKSvs89R9YZF8ohxfUQCGRHX/Nn4mVf/2h60O77kIwUid+KQIeTjUd3MiVw5bvtx5QCrc1hmuW
U0hdut/NiatU6f8WF/JFeBLMDQ8EfhrU6JxJVt+R/k/3QQyxWEKErywznTPJaf2swHRqSco1Xv5D
AJdKJKLENaEwbqnSqdkHieuNmDwlHvSqyPrfF3sRZ5UAhLk8c9INpsEsJv5fFv1JCe7iipqumdCF
qysROeRKJn+HLqtySwIhfArGCYAd8qkwiF8xsyWKS6znEedEr3toUDoOXG/sXs4ZqRsjY7If50GM
FhRhXbOGRq1lBfT6hdSTRMUcuTLbB7NZH46kOOOv7f7B/k0QLjW5MK0Edas7rjxfVmszH+hFmHJK
PqdnYTSyTTjpRV8IMexI8uqdGiZPnL4wzUh5XCODUHkMZdWUWB1JBz5Q/aLdFY5PKRq+hPjqTKyt
cI6iyVgFTDlP0Vjs+OZCW+FnTdtaTXvul9oarHFjfx+zrHqlvcp9U4ViPrlJD8LrpZghlNOSFRWL
iEWrVyWHehbrVfwNjnx/rAgfFAcN4l7v1dLBRy4Ab5fDsT7tDb8TxULdwRaZyQ3IhrJGy1wT4lC1
RyvhXrW0cf9i95KN/1EUlFmo70O9iLEpMfwdolFKVaXqGaqcNY7RgTa4JtoqrXDcoD0naI9fVGrh
ni9HezoT4BDKSKZ1lIg5dDQoO07Xjfr2v7OhEpjMjo9N6E/Z5QC7ozY7u2Esx8zEq0hoMDX4mhCU
XHst5gDyha+PvOZRkv3s8hzRFsHL/nkeQxOKKUQbC/iY3vVKnCKLDfL4AQDwHS1YZxVF9x2xB27U
7ecyhWVhPpe5VjiBjQkvzyJLW7T95/gw2lOlMcbEEdh7Q+/ko+4kpdADp/oaG75W/WL6t/K7yAO8
NQjnIW+GopCqofs0gYq3BzgM+4M9IMiC8e4bdNYnZQLMpOTa1zgmooGC+kf2uE02frzsKz9a5f4q
8Om6zIH9KyPZ6dbdVEWylZNd7Ex94ReVJQgFpsq2Kc56A7zr+Dm8R8uUImZ3OXpFJMm8w/KbOc5q
ZZEigH/ZF8GwRriJCCC3whFScS22KT6IJmRXPesMGqxUCcAqkJlXapEwMB4csgR5W81NikpNhMTk
17OJoIhVEgmOiC5WTNn3qauvcymPmDhFpZuhVKyWnMBnMA9pLDQuaS4sQhqeJX2mn7Zz14rSd4nl
5vNEfRXCIgg9VtFgmH0xpTh5rP9uswsM5f+/KgdAW/owiWGQv1UhcAJqSk2VJVcZehJZm8pSB/Fg
CHzzkIhT4nJTLKxmYWETwczG8U47U0B9FgoHtuzJX6afv42fo3bqjW2r2YJEzPC+xhEm3ebqvK+4
8AOmK/Ly2h2rI5J23wQyJTCkgsAv4Q/YViW+ENIHPeHav4bbMJgfjkrhwsFhN3YI0+nx5sHLekfa
2LTI8lS4/AJO205dkKOfHskuqPijs7KcsKgV9u2iOcOWtTWJAbQJxBd4YpZLW9hLKY7Jw6iHu3qn
nFpAsas6JvqwQicIg/QCuBWdi+kvqYdezy5fgFIRdT8Ph+mqtoq9+TWm5nA9lIGKXRh4WZsk4wi1
rIB7ax6f5fNv5w4VI9Mr8lfyPkMThFA9x3xDlLAzFXyiy2f6Cak1Ogdv4SQOAUedXIxe6Qbbtb+d
yLKDgy7/Roe8Px+cbqjUosCi2VZXh/Nm1yCZxAaBJTWZGbAcx1vUG8oqqK3+/cpDrNx6f1s2hvPC
XuilkrEKFL4SI4K8Ne7JT+ifNBht6/szHMwwwF6Su8Jqt429sEuHYruaQ4bos6jX0xoBAiOoNeUj
dqbMTu0cYKQNlyX9SK8MhicCbxlf2yguknU7PjQVtL8WHHNafi1YR15PwwsxSgA6qqQEm15JaLqy
n3pyp3JRqZs56NQSAAzxhP01m5mhxqO6huEQLBk2H+P9nzVCZnvzn6PNyIqqmZ+LR7v9KXHjvd44
DnZcCibjAs7DUjHmV7KZ7T8aUtOqTFPt+QKZzoNw5PaiJl7EjwxXzHzF+Sh5rGPYrrvBObTjkz4Z
7g2yLrAi2+RWGffMe9OwVQkCoMzwHclGT1nc+xQPVV8lQKYs5ZNbw6dDxbui3O1hGu9mADJXqDf3
BkROlIcMSpMnhC26F5oZcl+rzJ+ZmOmKea5RV2pFV6HJ+O2UixpA7aFr1OOSljxX+9yTnBTcG+LW
pLTyMJWpUKg8CrzjjyWRkZqtcBtgIgKcwfFrbaWDCT/0HBJXevCNaSizqnudtocCudp7CaByNhJO
V2PHA2UnemR50EyhKOwJCaVQTpPtSkWivTvfU+ytweSNvzarJY1xmGSTjzquRk5zXofrW1Tdcl2P
dua+zGh8i8wsTaQuGO59mBJENeqtWu2YTKrnipeo/RgiEImlizD1umh2KvnRwoCnfWXEhHg/GZCA
QXzfiueAQY0vdHbmQpgNK+VrJ1GCN3XMtgoog94ysT7XKFATgmA1A9sYHVPChlf9SbXMFDrPmrlr
gA1w4VPUxmATgB7vgCEIsnMpY1hUj1V3LBBD7RaOlgxHh0NymaeTh8kVmmHXI5/FsgUfgn1sZL4+
cPr/mwN3Nt3SolaXgqkrWMQYIfACby4t/O3mKypTFC848YYC/HqygkKaThT7k3ojaWyhEyhM+/wY
Q3TNMszJkiZFJh/RIN39rWdF7wGNc1tkwQRHAx6e6L7tDXvXNtrx8VPzwviiQFL9y4iDFqxveG0W
LB/dd/ERlwLwpc9Mng7dGC/+O53RkkaExAwajyBJ/wPwwiKdXvgFAKH+D2yiR2NocNbB61lG+0kQ
whRsHkbZ/Ky/IXQBA0LvC5nwMok30dBDvuGcMIYCvwfNMFzdxwRHE184Lyp52ZCNF47hBZ5kdsUT
Z+Blh6BAQRfpm2Z0wo0sJrDQcLN/Y5wyKvlcRoy9EchgkSOqpTedSZ7vduYG0ljRUpSO9P95VVwo
5OgUsphc/6921iAICSfEBVqaX8CICHPnewSxHPk1+w/eVReJQUGpivQCzEiDE5DaSZvqFrR9H8nF
rBe4YvxYjZ8Ou+Zo8zWuiNb95xk0bW68P9zfbtxZLJF+v+DwOHUAOsrxXjJHlUPIZSMvhO3M6dK1
ZALijaAF+fpGIT7Qy9+e/uNLScqbUlvv7bJBKB1bSHp1AYYfTMAbtWoNLmV2TPSW3XjrqnUL+Zeg
hurm2GnQ/yM1aaVquQFG5HfSvkkS6Dvtmffhw2aj49pTqtq3noxdBZLBySZLgDPxgGE0qoHTnUoi
I4w6DI8Xa2QhVeHA8d53DbeivWgDWzzo3mP1XDuz22A1LS8kSgC/mPxGF4TlsAzLnzaGrdr3lOYx
kipCDf7WvDqXF1joTU2FRomRyZFOqI4dK+ApO0k6MZ2JWcx6x1JqXHbAh2KHyxWv2Wx22V7h2daP
455qgEp567H1SEiTriZ0PTZGPBzQ5Sn3Nm7TCErz++jcu2ZrBF3dDh0KwqUPQFuCuE4ju7+ZmhLD
k6MeMDK/CB9C0WoUv3V+xAaV6wxAR3002WKT72GpzeS2p0+MvM8wB6U40IGUe2+Yas8vRo9BSJy8
baGYMXw1YTNZNWZSmQk224tK2lQPio8lVyUBmymSnMbgBqgtr6QCbRAV2z2/l7OANVL6SYNczcyr
jYcm/Z82DE1+zwjNtFQAdd6yVGLchbk9F+K5RZmzOwAecy3YqSDzrDTtESk2yC9R0Y2kKzX+4eIr
PZSSm21RocG11rm4V/UH3+X1DS/JEsAbEyMkRMJfoDb00OchNzhee3eT+0MrDqp5eJcYoqTknCde
KrPzUR30+WL0PZpd2MJDqyO3RDDq/3kc7IDgf1fzz8VE50JU3sNlq6rkSiyFQp6C8fqxWG6hhdBU
HED7yAVU7rGnhVFSgEvpiVFQA/aQ4+17uuk7I5DsOuAt3r72u4jNsxhy87ArzugKEMrf/LgycJKF
Ki/klWt3QTp/nCWs8bj0XjsD8HPTBqHGOH+vusNRhyKP5qAjrjLXlvu7PPDr94Sp4X3WkIRtm29W
0yczznV9GFeRBrMhNl0Ke22vJfsZUqPqs+p2+5zDIJspPjGdH3W7MPObcUs9PrV+yxvsR6Vweree
fVMhQOC1aI85OATWtlTEmzD/sTPho1BTmppY5hvL0Gh0UP/XwZRcSrwXVcVheUmtB2KSfVYxTtNs
K3+MwaMUiPLyaXcFAkiL0vIPMf1sypc20EkNm/lDSUXSxYyPLOBum0IO8Pdf/p3TKug6aP3+cH6z
AMOs/cTXRzJXcFVwZDyoZ1x7Yf6M/ZovsUkBmpHunVE5p0mOh1GoNre3VXZGRzyaoxQ0Doc6lMnJ
a+fRhKwAS/twJnlGtq05msuw+NF8aZ0hTp4FhulMMcUi9votuK2XhEfoT2hWIStLThxwrUPDLMEb
7kVUDnfsTH3Dec9DHvD5Wr+I4p0banqKM/dH9tjMHWr5UgDvuWo8rZdrg/4m1dCGu+2twmUskbVN
H+4XRfGNSFHJBpCvbWJ2Fo8EcEhrFRwlzkWsWmcgnGUTKHGmdrT0LmA29nMqakJGRsQYgbMFA7g9
ZunGNRuSoeuz3O/6+GnxfB2qOZOSMgjYc6RRhvH3kuA0GbQ0eH246Y7TgKHm/n12bQuhPYP4RGct
JbY8SjJR8R1IIAUtmJhBHceZl+gahRKL4Kb0rnhgrr+53fbSqKYOaCyKKUAskF8baUF3VAR7Uzm8
fkRCN27gUbvTYU5hHL+IvYCbRfneWnsF4hXkw38eNEtMlSKYV2wBcYEeJRr/j+chDHryAcgljPym
mkTK8k/1qeZZ2TUJ8DHyv77w+qWzHDVssqINbcmkseFyghr4hWPDQuvmuMiYZjL0YWL1RBH7JqaI
KgO4LyJGMk1T3L9BEtnLY8e4YpTdL8oZXyf0l4YuLolZLAoIZsGTZzR9tNideINI3kFQ1RuT4+7f
xOdvqsy7l+lbfdLn+NRea/8BMIC/wveUOeUyy+viKP5WTvGPU5vWLyK16cweIxPRSPXGZiMtTW/O
iETXvMn7KgiH0osXhHm2wnAVpop+TCyfQx4IkP2Bem85z6R8S0tjITGc5YQJKAQrSb7Rp4Mct6wR
0HU7pH2oiQVNZDy6U+oKvnt66FBovbpX0lsBOwHLAT5SgS24ms6NuwuxsFo8hlp3nxPdi9NAr76R
MhHuexMTXHII3XBFqzHYf3kfIwVemdas1LHpu14rIKgk0CavEUFIwyPJpaJoHy66J7iPznkkrbAR
5CDHa0IWLOszovO+JHa0nQ4+LEUSfymQn/3qsnpbE3chPmXXD0gD8quOXgMfQ7OOTs4IUspVIt/8
bsO1UIFC4OTVr8rCGzQMPTUbLXBYJGgJf5X5PGdlCCcg9Cfm9v1xM76PTANmPPuhRLnzyWwda7Zk
erzhdH9pRn75ghWbSa8W+qHub9dg61muv7L+6c528MG8c2FLWxjjulUy+ecUafYS9xZmCrkvDHpn
JBKND6/ydqc983qV36EWRVfpBFNvFDGB/hWO1goqRpp/pcKGBN6goefF9cYqm1sxW2C6UelR0XKR
2hRybry9TKytiu6MPE5/7tswT6WsCGyQjSKutbqpsz8mheWNVHaku9iDCXzN0wQXx/M8r9GuuCyf
7IoJsOrcEV+4+DktNilTk7ClnOSphIqdmEPS/fc1XI1M3nibaRYd82SxJDRSrwWuUIirMwBBoSVK
9f2xN5g//4SAEQu2bx0GL9rpYSOS8kWSkggamxslWgELhH3h3lFH058PauasNoL60cUr9HxGOKzJ
jeKRLTQEx7P6mX7/9Mo7k33j6H/1F1chhFyLv+SX/HiNqoMtfAPVXaRiJAtkRWqh78j6iIbpk8MB
LKgratouiOt2zCTLhs30ZzUHBTZYZT3f2aRubQPR5DEG79BIrBBG3TtWK1l5lFezfNMFHlOp9plG
P2mLyAbzeQ6GgauDhuTcLRVPPfhg9PuYQfEzFxHN62jysFGcvltsRhegVba9/M3HTct5AaNp72QN
QzpgGrzrV7Xws+WLdJ9qLyRIY4SVSRUtW/HRUDIJsIdFBthABu4dgL2D8TgfrusCefNg0FhzRse3
STzF3RDSyKoHPJzg2J3g3bkQTbwfzgPAbbxTa1ZRhVOaOKi0FGy/5D5PrK3pr19VDUxq/l413L2q
HVd6tpqhJoKXZ8MabXVycBuMwooiHhE5u4bxASEw+HAfjPTE8GjThv4LiqTMRQcC9T9RVyiZfFu/
Nocx51ihiCxufp0jlVTveRS98fR2ZB1Z/zvCT9coX1Hl60FQo+RGFDJvP9XtWC3zqcs3FzToMoeV
P/iwkQ+zz1rKcqF8kUIedtE6T6hdAjWF3NgL0IrQjCiAutNcIQAMSYC0v6ujbIQtwa6oHgQ9ONGC
SWJIPQH/znTfWZrSQKcYo6MQilLiTmjiEdY3tmKTfSqU/35BWH3K7xUbHqQpCmOXh2rqQuuUXUGJ
hUVikeCRmMyd3q+sPgNYz/wdXj59FVzTSmSsv6lc1pflifMeFKDQ7qH34WHQ3e5/Xt3sfqW32R8v
WAC1QBm+deJ1oPQF0oP5SrEG1q4pVt/0bHo0tHBx+8Y6YKUwurYuhx0v4EdEdkXpbI2eqqTar/Ux
DWfYxK4uXZ0L6eeMgzqEQC7SJWvqW4XmWxmZDOiWZgpOov6WJIYL3ykIufYPdz7YeEfdHYXzIxhE
3Aztu24GToyhKaPkNHyhPlKGF9viqfC4pAYB2tywamSUs6xE/svpnIJQD+FRKRE7Eo9RFu9lXapy
ksYbPhQb3kmUrnRZ9M3YSkNyTu9yXosCNat3bj+JrbYAnzMhRb2WftVrIs1+WAwUi3Ne63snbNT4
Y02VS9DQO+iGBJ+8OVB21a0SFdkIq7Ab2KMPWQ3TU0p12yeogV2D5aOe7l1SNSHjM/yTpQXafkv3
26HwdUmMMVqQQ5IpmP+1gpvIpov/m8XDrE5mr9Sj/9qrOjZ2sHU+vyHZTTlgvpId17ciT7uZ+luT
iz+M8VN8Sg7udBCeCmx3Ug6YK/re0Xxn2YtYCEKHNpfHZwsAN411BGxSvwkjVvob294Q9pZDTenS
yU7YjGAcsKP/+HhUtwlpep341ENhJYoWhfSD6pjad+ubQiheXLDWqdqxYDTvLh310Reu/Jib3Or8
0Ag7jJebLmVdQEdCgAjyLcmZ0BS4HFUEESg4oook2z/0av48ukzu4iw8aN3r/ZCH13Yc+jmM32R4
t+PXcQs90ICUraERrR50bR6PHQvlWvSvXACPU63TYS9QruHYGB7wNPkwUG/f0E3/YWtQNPGXS6G3
I963UV/60hkcM2u2BmimCjlhuGUuyty/0EhhB3k8sn0BD89O+prG8n2nVqBTNGIT01F+5QT7xdaf
QjmaDs/iDTd/LG+pBDGWPDvmiAc2i6kV/s1Ugd7AMdM96PS5IjMW5XAPgZmvTpx71uxQ1QBBdIzn
jPc7h0MSVEnvtn7mFT4hXH5UGlIWIr1XgDYNWjz6mxLZ66RcvaEi1BJcZ8D5BCxZWBiP1xot6A4n
l6Cyy7YBX7fMFgdTudFXcedf7ffJ6pkwQXmdP0I3J9gnaQjQSJ6qgPt6DO+1e9FzTBb2l4XSBI6F
zw8OwYiXydLuv3UOhttQcafiMKBh5rtvDi7psGsIvbXQ6XmpRB6dMBV1fSziobWNBo6ioicxSGEf
EguptREeHK02b9mAjn3ghxRNZrhY/GF0u9XeEMoZkfTo2HW9s1+mGjnKr3VMIdIcrHNGrM5TJdsC
quEe06XsXVC3MoTdPE+95Xwvda6+6I/lOtG+4S7DZcDQ4m7YirCfRPeikq5LCdkmpj0nciDJJvNK
3tGLwwlzSuDHqgismdy9ru713uVcS1/f4urtRe58Vb4kzqmQyIf8a39J162C3oRC+ZbveyqtL4o5
738N0y9266grLZWTO/S6Eq4XJn1H/qtENslNtIOCvBn7VKSfqMbsFNsxAEQs1It2jsTT1vWfQoxA
02Q+Rt6N0250TJ9D67sccUtIA/dGEyTvv0dTUFRou6smfEb5ycO7VEQ887EFI3fdhmmFwgkA4syb
zGixgxMw6we/sRWY2hfNwhwubplgLCCLRZeWIzNNYAN5M2/5ChZtw8stkJSKu/lwYNmJUgC9hPq9
41AQXYpyNcj0kFm7oFSVPogMi3hWgoiOiCIvAPxPLhpMNEQixDbXi6Mx+lId4Y9PgA83XxIoLZY5
4DqqJhlnngZr6NprjSAnyMqsAJx7MPIO/DaSXRwyz/20drJQUk+6CAWXNmcxyWQL1YkB3eN1kOze
I93Oyyi+2Y3xJ/lV+pE7CFnqrRYKWggAOntF63VFBcJb/kxggkLiNBdfzKxazzeN0eI+m+Yn2sBf
IhuTby+YmqxtZbFgDbzkn0ZXnZFGOpkX8QFtoiDiW9ZINP1J1REeQ+qeHAoCikguOd6tFRaRxRL7
PZ2FMKxcEq908JdpRDULdR2rT4mZ88rl4YunIkiij2ifMbOX4+D634xHFtd6gCOYhK+NPu6yRmGG
CwHcaPenOKBtbBY06Q+/oozpHZJfkLMD9lIP97H6laNJJg+vdNKLgD/C22l+E35TJF4QYchbGBar
VDtChSNEmKT5J2U3JGxbs+Yn9NRSZ18907ej/C+0RYLcAmYymMzdfH+46BPqUR0bVQLTqcEHeT+i
Q0L6wam1qSUSY2wUNSKMo3Bvb10BDwPhh669QSHQKQm0zNZP2jdRIzn58UtxoTNk0ZaIcWT1pRmf
6AHUc0AZf3LP0CB9gsEFez5cLuO/RCUHtAjLlYwXhezI5kGF8PYaqPbVjLoq1el5Yn4Pqj4K6dQJ
Cn6/e2KkBVNSJKPsEnnU8in4R9+RxNMpfAQYiBYWCkUvWzHoTvk2t65fU/4iWEhQ5Yi4fKSWdh6A
N7i6YvoB8OaYjQMGlhe/p5CgQdEN6Mu/i8quFCntaZqTaNLtBBLNuAZOgJ5J6iTdUFN+Bv3LJy8r
7JqcZsqEj5ei7jOhUCEUuaIv3RuwuIDKeUm3+vFiR5h5e43fRVVu7jIYUayw400QItq8TzslkXK2
Yy1S5V7/Uc2wbvYFb93VpkuFiO2pZdbrzs4Ic3gnSXinPYJX1P63QC9QCDOaYoqimpYenzTpgTkU
1rnerUHKArXDHLz2MWvuZxStPQs8B6NWGIObzrcC9fbYhpPKGWJpNmKzgkLX4hBobyz/j0mwo5vj
knisIpIE86k4CNeUsW3V6gPIUs63ozGsM3x2AgIpA9ECEBIjNhpx3wQ18ueHXmwEeiEiRygt1jnO
cYQtEbj3jcDr4gPiuZLB2bvG5rhKuKhutYoV4/+0Xl75BCqvOGo3OG6vY27W54RF2sSFvm1OfQpT
uosZmi2DFkrSQ1pfVVyu4QpUda16gUrXZRKRNzxQvfw9FEunbPfCg3TgmQdBD7FdNRWb0VzVrxpO
AOc4Vgxw0I5ey4fhyprOpghmIw4s6/+s5Ol75SlHN4d9QSVxoly5NjKE1HtnfDZoRg/OWC7epFb7
32GbrGKs+i6RHrL/qexALYFw7LbQuXsIRfTtnyVFPugMkvXy8ymRgw5Adwaa/v6VdyN2kbQ0RMYk
LsQNiD+vgcJiSYxx1ll8UMIfZvQLG4kdrFAbfp9gA8VkuuP7DGqDcBcI484yQdKa9ChLNMEcWO3u
oEqfXh3WSMBGsE4oTMFyPoQ6fKHJiK5TIQlrzsot3/j/26JgV2cLfG70DShgqQLOqUdpWamblK9t
OH7Hw7EJkiX5TZP/qnZoLpdh5irkJ+79LtmCZZ5XyGLSWQd4wDHKGNN2q/TNFfPWsAwKLsObWEB7
4Z1WeW+XOy2M9+VqBEoCiA90l2tizrNlJ2/4e8GF0f/dJgxlrW/G5H6EuvEyO7QUMRBJwQWS0XOC
EKXCkLy4R0C1G+WX3jPt3WilM5z/EHmKP+Q+022JDqCTCevMyUrKgobTEDHIx+2GQJsl+fFP3N/Y
8LhTIO8c63Z14jmBk+VomP5S5kVbQ8i65vvY8cI4Du97P0M85poOPzY54XIMqHKf/WqOIDnmadQZ
pFRatmvWhmgLnGd0smKkcI9z7hbnO9ISbebXGzRirCgnLtPpPbKdFb10FkaQjRGH3Td2/XkxkG+x
Ac5E6rTqJYiErI67OFgfqsw8O/cxPMEzZfcl4qOdyFGnT26Kuw8vtZhLEZo3nvCPfaPauiBHG46S
7dRQskQcX1xhXGAHYc2QvyGZdLCO5iezET/pCVHtZGymavcELIswZOwR14vGQehVPfzCud6qzLWy
iGYSAN7Feb/itmTo7tO07CCC5Dxa/ro0CB5Soth6ao2+pp1zk52eE6tXGC9bPSfCBT7sUz75rBva
zuFgnARgHK8GJILHeElsp1IDwI91Jqb7FPGW092yAf3PlWBZkg/0ZBmZrsWpLv6OT9VQK27FyfwH
xOEqKCtFERZVtTz5+QuIyS8HU8d7aWegTmvX+8tehgwlzUtl1rHhSyTL4bg7yJV1358OhQFRZF+c
d3YKq19z4FVNhbuX20J6mOsjl+DFer+OZgWh0hTrPJhlaOAQIDkYwM4NbqyulGoV3goOiBbz50J/
+qTwvjvMIheFGTL96AXNHNTUnxXqMygkn8WeDWbqcNNtPDEDTaPiXxQnU93H50Bh/HvHcw3anyoM
DquILDsRBK6m1kn0DCY9O2kKnIvRCAUVdEXY+xppcnsaWZ9YDoA9NIMfQkSNOC4n2mU/n8AfnJ33
aTLoURPi/pqGCDImOXbszEEp//yUIgqW5utF0ZO9fBFefR7/DqO9uopIaT/sPtSAFsAHpD86wqq3
BsUXMKFm9zgh6C7rnWbJkexTGwBpbM4rWA0r+H56vLxvP36MMCcrQA6CSaofTtpx57CfH574q6nG
/dXnSQ5z9a1oY/Zjj8gnv//SPG05PqeYxANqNxdEU9xNWoPea4M+K5EC9OwKVBVDoCW6GHkgDoSJ
Tz5Y31hygNU2s/nVUF3k5gq5Z4XdbdGWcioRYt2ZvCvLerPfmfglsBg2WK2NfqvYHaRYFliyP7CF
YicND/8VrSa4H3FAERN24ZzgnaVjxpXjBq1pZCxPQbf3fPwLX3O/tmnGTFVyA+C8RD8BN2l8FWOO
q6D9qnZ/aAEXbAQODYp86vePAbwwtZM3ZNKH8VLYMacsCvVPMW2SIUYL6XqE1uDSWtyQkcSplzSf
CrKxcEpYRB338vBORN8JTZ5gzRBU4IOWtcncZnLFRHAlAqAphuHGUhMolpTO4UUImCgL79K+Swbe
63Zy6NrVIUHA9AHV668VqCDprlL6qGfdx7/TFyMsM5a45zDva7MEoTI+AftnWcqHfL2KFbQw4ZdW
04o3ggmReGAIlNSsR/sslvtJjU+LmCLKEZG/gpDxpR8MU1AFUsfr9SOC9iJLUfktfo48e2hSGpn/
ZG66+ROmLOKfHcC2eF8GT+ipEnJsVMVm8h910YIuw29l5CIJ2wmkoD7OY3jewxfA70iSSa935rdC
FT9NFWu6GIRT1iI6QLc53ZO46WpNvYM88s5xKu1hZbK8B13NmyZ2tBCTPlGXhVQ5Mx39RYlOWH1F
AKBp/523gZiQ4/fXcIiVFeOZkJy9KvyEC42X9lcvjgiF8Up9K1L5cre0DpoPY/sfOGCAnbA9u00h
8Xrv/NHG7jyk9c9VHzGYy5dbxEvIGLrY0Phq9aWQQe2lygTY3AVBhqk/bzZu43ZYnsbLhRKSbR4j
sQJ4zqXnIImDD+NvfabQdTN32p7wG5CCkLUhN9Tjo8GSAqeN3eiksmillEN6MUZimWVA4y1AaN1X
q42TtYfOCKOX/sSpLvXwSjcSzKUvtpw6sZpKGsd8SBZDSGAYVQJq/gW8O55yZzerFq+fkuiodugs
U4+oup0UxjMrYlYuECvmm4l+qa5v1LAcoUJPUjcIh9JBn5IOrwPFDZpglyFwBKZ2E7jLGTbww6QR
n4aYMTKNZa8al8zDkvpVA7dD2lU1gW5ZHplrLtTeFwyIP3YKQ+nveEQjDBB2YFW+I6NK4RW/oCs9
XWLE5kh5oKxAJ1+uApo8ctTnrySAzFW+m+43aSM93s2Ez9eAqukbneeLi+jSzu7uAfrU874x3Tiz
pCHiuRBpT6BA+sjpewdqzysmV+mHk/4w4wY8NYoMsskIelt6k15yrbQ4H9dc/Erta5wydh/FqTs4
bDz8+DUAiVTTaOnA4cJc7x7Y0mGlZGrYKY8ZVZ6AHsSVeFJCPSKAwldX6iB+Mf0fahlcIhjkcUcO
3PACtTsKKSK5dw0NGm80DqFkd4vttGWTKRdTVuzy5Kaw/xHHZmedsBATxloSjeWxvo7ybMk/Bffo
yKUnoCLz965Ecw0C+2IJ+TfgwyukfPc/3upXJqwPaeeS1emhE7IEoZglXMdpv5q5p3M+3r+Ouobe
z7G3YwPrROAyojOfsfaQiOZIseF0XZs0Xr8qzsQXhL01e7q4VhCjr3gb2WuNpMA5+HLFwuAlNNUx
6pRcZP+7n2ZG6KOa/AjZkeSZgPGvWwVvpbA8xGFei9dfeVckGwKzEiPNyXgql1K4GHMHbcYlyHAY
g/s2yblqwt7AMfclj6Jsg1rD/Z+opnI1s4uEXhM1TMlMqepTDlXdRYBpSU9XKCTXA1jGODLGN3Aq
Ll+T3X7OL9BCB43JnTgrGCVoWLpaf1+gnH66yuyDdbOZLKnaKd6OpgEnzRIIhWfJNnd0zbG1hk5i
Ule9JoKXYFu/tg3n5p42cv8T1o8AZSVcwPdZZ9A23ZJjDqIlF9/9GH++XopUS7oPe8jgRaS53wti
8KuD/hAKF3ORklrvyB+TBx6B1aSVjjxJ3FAfjYFRWKZ0cPRe9yui6AyQirDBF3qVLrZfLJkvjokD
vgx4yU2gkXuJ6k3aldHE7ET9ZIiRtQ5wv3brIBEWKEKvKpf6Vxjtn4Pcfq8tV4r4aUzv3ab4+Z0C
7vhuttbhFJuSP2jeW1XyOceQD2z1gCQAMMwk0SVvOtmRto94KZBGMzmkY6DKjz5vQ8GMmm1nOOOf
nrZ8NcQEqZfTUwGdhsxctG6eUq7U5nnbBJ8XXjcjIxlB3AYKPmDfyQrEAjsm9mWMh0SuX2Ent3Nt
hFCTpZLQ7dkVyfSM5dvBbAThVD1I+C+BSa41psw+wyiAvu0PfbVAr9hTeBdYqKM6VCjmXi6cLFFq
RwRF5OYNIlUMS4TG9JoN10lM3MzT5ZmGXjnTtwqt7cs28PQbzV/Oy1uKx5oCahuWCMkPXsxE8pJ2
ygd2nmdXA76EawucVJwdLpfGPbsuHmY2pscD334EwzzDff+6TheW2QBhiqlQ0eJxWLhXrWNFtDvY
gYq1QgWKozSBSsTDgAQ+vftPh5QnhPvmDryB5I9Xnbh0ekIjs3JPf3BMZy452UXKjf2jS16xr+k6
vxJV58O8kE4/2qHpoKeiWUN7Gw/9tVn00r+BElACGAvDLiSFhRwaoPw35BLowEBjh2Kkod6lz84T
K4qvYzuvEHj4eraP4hgMK60m06S9TTfsSWmnauP5Tles+OMMuNs65zK9yzYL/iVNcTcxPOyhVwFz
QYi7ZJ6b2CoNlFuuOOehr+uAJdtmz1jlxcHPME5vNKhR2co1+kARazMFYtuAoWywIQtwHV1FyP/c
gGodO1oszt9hUsw5ei17agrAvNoVn8PWD56GB03zuo7+UOG0o+xS/w/11aH6H8bd/PonPRvyo/Z+
n5T5H/81B+WHNeOQHlyYVah+TkqxUrTmh4mrZVmDquIWE1HxedS3j4JI1Gecbb1bJfJS+rYmP5+t
6kRg2bv5+V+Fis53/ZCQNDycwVn0y4PE22dzk0aCPSXiiOEVjMqRPsGdyiiZCh1BNZWVaIf4FhbF
h5L5GeEW/n4QqF/daE4Cy4+stozq0GA9ESqBalqVGvrALqIeR2Ouow21gKUA+YhM1iDwbirXXKVx
ZStODnWfC7cyZ6Vv+xXCI93ASpFJjHowe99U4OHiJ6R6MBLLZyCluUESpphkDHsSvr2qemCxEEjA
R2uYKMBFWCkGM5p13Y+KodOy7vKYjW5VLJxzCT1c5kRFB29IilPm7R3+OuQb56XReby1/CmLUFS4
TP3P5kW2VNF9c9k7Y1kk1ZeeSP+RhIPiqDmgabt+3n2iX6zfZWM/K0d9TJmEKtvj6xgTsCKIhYzc
LYzaf4MiZwVX58LgoMCNiU1DIWniTmeGllmiRnbL4z++nFAZqUH3ev/8kOcCYH00k8jRxPlOqW3L
U472DJTtnEnCK4RiNgQ1yOmnGlSyQwfl6NZphwV+EXPoIxa0j/resVZf0Tp2XsS06Q2TkoqtcvUx
pkswYqGLMlmAv0DGIDKxSKzHEu0z1VJXbS3b5KhfLRhRC7PNkvM+rrhl5N5EgZhQ5no04X274UnF
+4OvTmlbuffzOIZ85GyqJUqCIlQ6dLYe8YAhTX2Uw/lytFaYpGW7gsNu+G3lQNNn453FUaUVUSM7
WIfcBkH89O9WqR32XVrJeG5u6nJTp38izjth6rR1r4EJYMxchOEJwVIMXMy/cFgDv/+4fkqfFNVK
sJFB1oVf6dfEHCUVi/xLInbX78xEbtzrK5wx7xRZTqkufpaXcR7obNui7l6NiQitF92qzWzcUe4Z
t7YeTDFZAT/99Np7ZBKYwbMCQR9ojPsQfgmjKQ6glMvzv7hghZOUZPJzGlJe6ZeKto+Od2d1LMur
Uy1Ft0OztrYZQFfFAMyZocbakWZlyDXmgw9GOWIw2/jOmLZ3YpxDtBCfBfWaOwG8t464Af20w9t9
8zqF7ReZ2YVIFnd4S2U/REoD0BTWukPv0LJd1hW26ZMcbpFJUV6gCh7JYqhgaGLr8hO1aGVft6iX
7iCc9dQKYl83UP0LAAyNL6C4mlS3IW0waST5D6e75tH+i2n5mHOAx9M3BBInw00leMVBsSIaN96q
Qea2rwVyV8owhXqEKmD9V4WNhm+3eMkRJ5LWw4rOMq753kDwbGjcMhQsvD0gK672O4A3KZewi9FH
TGrp8Vela4pVByTgqJB86ucXy7lyKRWOW1yrJhuCRDpprvF0Syo8jsP2WThT8Tl/SvR7xOsKDxc/
60yCIBmvoxPJKgCyMr4TlhKFwdKmtv/LA1PpPfecKn63ybsddm1MKyI5M4VuSZcCQoO6HoAqxRBQ
vfDLW3nEjuUaVGeIrFUpaLXPFIQv0j6y/w3AN9m4I2G3ci6kUjRMxPqlufBM3If95LVohD82GCon
QlGieEon1griiatLwvyC6hA08UZfnGcAfOrhPnOv5Iiwm2W0Bj5XhcpZU5l+qSarjhHloea2ZSb2
JdJnL9IKqRnzIcmMnihdOPWnakMxDQCvF6TJ7DcJgii+QFsVN5d5+CulYmyJNubW6aHUF6yvY64s
q+5SWGMUFgUH5IfvMyvbeZAdN+AgOUCByGH4DU9eMSRarar0n02MV0fFwYRwsbRviebOsTA1AvWD
N47H+8hwywTUI78QNPXo43WRxcGUrvRo8j844sRLOItX3YOi5Dt6PfODQ8+rlSMDwpxvsx9ai/aW
BxRYTcbrN2jrSfbjKg153VdfpqksbAgwCSwbChjMo3Ja6ectlKS1hxytUvO6ing5JrMK2tvtvJ5b
ho6vKc+TcDWU5XSsnkQI7LTB/x270rmwDp+Xh3/1uS5mC8gy+Xm/FVJ0ygQ1k6icjWSme3EF8eDD
g9MO7s0kgiLeKaO5NlR3BnrUCU3Aaquy6Srkmn83bJaMEnxU+4I3KLicap4zlXAmCc1eshOREHdz
vMg0kPLwIZMYLbAFfG6XgDeYu/rBpu+NzHX+eIycf8t/mS9Ig3VelADOhC1seAHCwcD4s9yj0O8x
G4r79soqRUDgv7Qj0b+STA1yln8xhJ/OvvaiBBMSISrgDAQ1aPdewrOH67LJooA7TINe+3KRc9yB
W1hgNUQqN1IjwYHGXwkBHMVV+sisFZ7FYKKFdXprZ0kWzv4X6ThR/e2BN9jLaKkSKTcZebFC9S7U
W38hL5Fo9AdCG9NvB9MyceUb0aPKOk+Fkqudlaf07/866hLNoLmtShnr6bU0DaknC1XfvnJWT+UE
poKGPtON/aRVR8LB9IjF+2QmC0vb3aBYXtNPmaHODq02oX5K5Wz7z5LBIZDFY1sX7q+ELGkFer1m
rkPOlenHtrHRreR8kfPGySBPBue482htFceGrfyv6BOfF/DJPi0Hw+CPcqqPfFHJH8FwyaC2Yvgh
MR6yIOwgXQyS0sahryFDBFieq5vc52tc+03MuTS3XTgWPKqe2qhq6N95UUISNENDnwaqT4dpV7PG
wN/lD3HM474fZDVtjD/FpGLszAgQUzfRo3gJzU3iQ/DxawCjDDYTXcRYHzBziNwO6V/g5o0ImSkN
0CGUzC4SGTNmmsm1TIwGrd7tiQ7cGGqcjJGpAB1cE4nPYbu+NAC/bmDOTuRfDGCkcPV9+AuzJsFo
vq3/V+ztLSW44nVXCZaWjtg75cgzBiETBpy3Am3ktqTbI5zrjIy1NLAo4uJSre6gKatTQoFmch+0
qJoXbe1zRtf+0fUMN6fESsrJ1EjC+OU2aXlheq7p/TsBJ9rcGmoX0v9EpsaiPo++qiQTK+Nm1zze
sPeMasxdiNIaZyRTSaFi9gteAXxTcIrdTw2dGhYvmSRO+f4Rf1JNaEOj+Kjvsx+0Bgveoxd6fkcg
gNpOC/K+30Ya1jbQ1dayN2swbJFS/4bOepPMZQUsADkgVKxT/9lV/w+6209/4g46doIVtRZf4h6J
NaIJJvdsJoAtRe4LcmTr+GcoV9jCVElqySTZc5p2VC/5bBTI3OzB7qrrGpRiFdJwHXpFYjuAYJ0M
gLHuSc5kD2qXzZw3zDG/Grz99LrnI3LJ2mR6ZaskhGdn/oZE4yYyDCqy03vYkJ9eujANYjhLk5yP
DQmsaJBEkInmPASpWZtj1U6+7gay4+e4095OfxyJCMGP2kPi7jMq0rzBm5Ca+KFh+4RN/UIvXfb/
897A0C9Jlq36dkl/rms6xAEYDTnNm7JDcaeQcyMOJDhhwViD1uuq5RNBZ28U8/kuOZbIjWyHIke8
1S9nfeKfG+g3pvoZEk3xhTAUxOXiLmNVKL2R1AOYdr3OLwt51HtFz28J2JTchVmDOZ0cVb/sTOXx
MwMggT1vEUHsQZIdYJGUASZBFNp1u17YRyQNAXLukt9pRyJTJ7KsH6B1cYMH21Cup23azDelvFcv
5Qg3EpWomMfWATskDnoWirHRLOnTZ66ZoMKt7pibSA/JExDjlKJ+edjfAi2ETvZfDnzy7atHMOrm
NQ8tNO0uUHXtvh4wzDkq7dOUcow+fPMDA9+TDGrPsSDxjJMR7L11S5Upm+XbHzmGZyXl2zXwHkfh
BocVpiGfAVsiQw6FBRXtynmR/qSzft4JR3IgDLLeRtIbag5621KAoqUQ2OPBOeTYNIy2NqavUSU/
Yv9bCi+EMspYxaAKjpRXg5+zX7asokWmXsc6FtHbgeIm6hq4KpPTeeczVjIJF9IKP4ihasIC3thJ
MD1ZOWnAjnfWIZCqzZMESYDjC5jIOyFRgLjY3+nbiJ8lyQYOgFGefz21JsyORvtbRFvvJuD3boyT
ozcdY5O807v68yqWLtlECHmNeH9eVgv039xJa3yN5VhXXBMFrV8CSmqjNR2moSxuG8PNW76gPavp
dDs/vLs4UYVKPsRlQo212JjR5B3PdSj0deGwU6TjOnPFPGutlk8P+aAUXep91cLYKkuDwL/437q/
xq8gJgk7H0+PSUckKwym7NUkjBJIfSn3vM3GRJjyJQV/GneRpb1A0brjKvR3P/u1DWmREn86bX7D
JLWdagf6BVAiC4Nq5WwoD9GkPXNkjS6DmhYdmtWU1jAxN5Q/SzWP81UOPas0rAn7gm5Ozk/z9rif
ZpAS0Rd7JsV/e29qio0k+hT1PGSnVNxkjvkFJnaCHfGEZQd5Rrb26fl++TU606bEen2wY5/GIMtA
0i8b9grKUpLI+bOFDRVmsExGgDuTkJhz5dRBLBmTS3aMdWD2Hck3h7iG0dUIj3NZ/P/h8VW1yIlC
7e0i7VXNAs97jDNAbR7gfzDZ0z380X282bNDxn/8JE8W4OV9ZhqnunpwVrMWKCefMV+VKBVxi5r7
qjev+On/2CqDfu7aQlth9XDsJNphoplk0DJKF2A+GFQ8Pa3SrcBqDBnUmqBPzVf6K9VKB+ofAXlF
X/aGfvfFw7rp1vL9UQ5ulHun0geZVU1arxBr13VsmrkQfDovmyxYv+NCOADdk8cBjyW+McRqZdDm
nvGdmZeFSkUbfLQ8J6VtfDzPAWovF794ZR07cqpZWFFJQ8FfoPPzC+DJit/E7Nii8aV4lJd12YC8
wQ91sa8ZLgztMmpI2mvbWlcr/wheqgvQRYxaxBQRPZGaiWWqkL+XLkDuqtj0GxGcaEGEsgtLwAFe
18VE5L3jvWslAOpA3PnyBS7mYsItX4q3LJkEKpRJ0SfYiTTxhj9Brhs4T4uiSwbbqbT+6Cficl9k
AjRywkrjn7QZN1dM0VPRniB1R8bkE01a6tBBnC/wxACWqqhqXHKRn5fzL4FVTY0dylfdKk5xfYvq
JmbZI5+3yAjnWHlpw0Y7bCUxGaH2J0P5lCd46SjLLqoZko6MDLbsKZOwzDR0dpCZjhwabf+Pqy00
dJ5HPoQgWBYAUF/geivb4MMdSAog5+fKYNCNu40RkPm0FHjJLoqHIt1q+99zuPjsLa/Hm9YVpUfo
8mvWS5Y/ZyrXnO/QWOwDduU8XjO+eXteLzCm3r25dPtSc5MCtEvjv5EsgslqEy957QZ1kY9K4lkm
C2YKwQCRsaanQUcNwPQ3gqwu8rORxNKu6sp/hVzmkDzDFLgEQc8H/gSsb4qLqd/vTWpSjmx7LIhd
TFZ9o6JV3btjQm/SVEm2Cvz1fHw2YhijutOK+M70xhl/rQjIAQWCSJ8QPs3AaLgLwJRmobUhoZyn
/M3YZXQf1Zlc60RhbMSUhRr2VYzxZqY1IZQdRbd449XCBGamHVEy5Gl4tMIQsdeSRp1uSOGJvLeL
0cgVGw0MgA3yEdX1oy3DVvJaAOD9kH4oGFhK7XNTvbR9MPyjUnO3jrJAOqs4qzjJxNkbeY1gQmJs
O2q2euc7TI1+jawcgcJfL7O9/O29lB39ouRSEdW3SlI5DvKvRGiM2QVF3yuwpHZQs3PFPT7qsyFO
7ysvail2bgGwvrmmQyLbav0sHYakZF3WOUJvAdThcs0Cllrfomz8GBwuN9ruz+zicTeEJ8ZYvreg
LlsEeXW0jqFT+BGurQAV4KqBGBzXqHdPUWZfrWtpgV2Cc1HtG+9oLp2b86TIJaSZsg1BHaNtjr9A
0j/Jg2eEvVF47lu8LxfCcf8RMADxFr8BZrfXDGwGGEug9ZykfhHw2jWUgkvaV4p6QlMqf6wZ2UcS
MMfJCq28o2/BKAJZn6/W8Iw4VfAiqT3oEJt1SebvwHljLJ+wgMh8Dal8lTaE+m44EaR1WpOUKRK3
G7eh1YyWSHb7TAIVSwyktCNt6C5ho2pD5pp3JuzQ4tULSjduaev/ufBuh1U1Un5hU7O19PHqxszr
NdMx3FgtwioF8leGEEUuMHf3YF89m5cxcLAmj2lCZQ2zP52cvsR7QxHV5S+1qxIukgCZCGuLOWB0
1gG47kFWCXkJ5ahQIiHrnV/ofrfAG4etC6MMzkkfmrQdjJ/K5Re/huVYsogXQtXoUS68M3kEvbLI
3LxKEYqv+vf6sFR6JlpyMOAeJpvHqqphtOrho4qQot5nfeREAD3WtArKohXqNK7Yewul/IxERHMj
vqdlIb0nHHAQ7iAGH827p2T8SqxtUSG0whZms23dV2wiX4Mlhxz1R+kQ54s2DqQuVFzLkOgDupFc
2BUm9GLrcNILig52VEQdHJpw6W913CPK9kuyEmbJgPITYPGFgTutQ+jEtN1EJl5BOYzfgMP27gsL
kOZg9kVEfYLW8D3E8fY+tXnQTWIlhSW1UtIAEfU6SmWNzQIIdgKeYuaa+QDKWL0dy4gtg+IR955X
/PvdOApjV8ZqMRH3rA/bVjDtVsErJ9B/3DLEou/Tc/hEpLHbBMc+K4NnAu2oCRXwNEjDahYI2iLu
6GKu+irm8uIrDoLsdoyxWOKALBsyJA+mUksi8TMIeq5AZkgfbUDUWhjAwx4tARILUIcF+0KXVEfb
cXyWE1CV8F+SXzeYtuCP69Thf86jD7aMwaTPnpEGS4GeUG6O9omixe4id6+rdwyFDopoqeQLmbSG
3LQfiGohi48bc3QYQn+PKxL++3XiCR1vxJgzK1bUnTHtogc5fJpEfgTBC4L7wsEB7pf+zp8K0Pen
h0QQVfwyXL/wqm7FkKd65UcLKGYqYLR095Teif1Fs58jwa/mmkuG+DPs25PGs8nhJQ7vBrOW7UFr
D375n/oy4esWR0Tre3ZaIIaOwe27IgJV49cA4mhyDT6TmEm+3SoaaHz8dWc7/LcRdZTytVHNy2Af
P13JfSxLUzmeTPQ3N6fDZ8EQEbiUPf2LT3hSnuq0NpUMuuxdJkl6PW7oWh1rEEerKBJwCca7Ey2C
PMGOAloXAfIb3GqzvJieJrffJbJGd7Nzh0+T318FYC9XKTfPYHI4c5uRvrDgHgx/NWqcSvBHiUFz
7VesJoq2JrXq0bheKhXJEeDVah9hV+4AHN6G5m/Ekxts5Avskx3GSdIjqEGVRDhfAEb8xT/vsFUu
yBWAkNCse/taZNeUrdCPCNXTZV7ZQMznD2hLd2csyLnmOnPOplTYX+9t3mkFxz8XHGKgV019rmq3
9EL+amJW+gkqE67zlaALwlAPFFzY4hpfQenYDuWrDqzEAAwvW+pDxLXb2oiwtHHilP6EH+8YanyA
gSofR5+7I1nMF9GbDCg+P+J9b5yjif3w5xhQJIOG0CDRIB+buKqrlDUSQJglLdV++asIdPmqoyAZ
zlBz3l9e4hdc/8Y72Zbi97W1P3Ryu1nq/bBr/eEoD3MP/4fENljz+MBnEH1vMC8lzTH+bStyyX7E
Raks6cGtL2zUdb2ECpOUwoXArSR3Szs5GVst+H39hVKCQREnQw75aV6FzPFBb3mAorPkU4rpgVkA
9fUGjjPC331U2B3v7bie0wXJ5KQJgB+oa7eCgQ3Z7LcQPDtoXmLsP/v5HB3NVACElWFuWC7bBDib
MsHNrJlBY0G95/k0tejXbv6olOlQHWDIJiF28v9XNyv6lxNZsLpMTVclZ7OYd6zMTRcOYHSho5cl
Rac2ki7SC/plNc+9DLUXjnBCHMjWbw+CXNdrZ6xVvlFD9573R5WJpj2NofFolDMNcokSpOt3I8J4
4FHBHmmHU716trVcNMmpqaa+40qh2qIhAHujD0euonyAxqb4aMWGgmsTjwLxyRurBNPmrGOV7J7G
9SwDDfvxYnjGegMzB9/nYlYRt6kHfHwKt821WECjOwxP7fCX60GC8f/RAa96K3BoOCIAfLmAOKnF
eys+rosozLsSS6qPD+fvzIlkJUTEhbsmN91DfTknH9MrebTgHsoJ7Nizw+3CPRKifIjeV3kThIWq
1v6dI7APikvqGQgWL2IPCwcBSoPt8LXd2atNuPcUNh7V9OBrxgSyGIaqnV0YCemR2AhPb60CspzS
cRgNGDsfFrb6yA5LLgPrkkPwg+06rLGSxqI5FhnXmpJivLOv02TO8jiYJ92zyiuZj6y4UkrIlFfv
+14fTPTPmjY9ehbPV+IV4kpZFb8aRDnh+Q/DoUFngPnmdZUAthk1GI2N3ARSheZ3k7CkCRpXJyMo
GCaUBXaMBor3qaRqHBHAEduDvTrPfa5DUEdyVniZf/HpeBnV8iJHu2sCh4/uYn9JqMFuRNcDsoON
e8OBcQaaduSBbiK7o1r/Bxlo5lWLxbLcDH0EfVTbYcnQHL8XWzOwjoUr6YnoOl1R911CcA/OsvkE
JxQlEQ1UlzNCFMFgJWS28iBmah3LM+hKMAUmaKXgSiL4ZA8Mx4BJDm1f0jhIJNzuKQX5DaHAFdp6
EtsyYwpF8t7ipN3212bUs+ujsdB3HsXbDTC1XuNcWYF+rYwyJyRo6MVDisCU9F9TBWp5M9AB602v
nIXeZ3xTwUOaqVzNAjHvE2DfEtaA/JcU2ws5vGEhcDqsc47XTqZ7JLevuJxpBQOr0tzdq2BPdZfg
HXEIi69Kj+NmNMT6sRFifsymTmegORU8qcNbFdXAluGwX3HM738rXp22U2V/l1w0osTsJI58vNUV
6/JTV6SA8ywoYsBLaBwaHKeS8HxFPLJxUOSfuH2Mr1/o2KaUMYdo1XXi8uJzufO0wYLwlES+kKR0
vbij16WqjJmZqKQWAtoSOmBZi7qI3+Z94NH7XLAkMWvVoX1rP/h/7m4XGgtRKMMQhGaHWWS0v59P
Hdkt8ib/dV0fEm0l+xs9OFo3Heplbn700p71C4LB871KzITAWNwPkOIDvAEIrc7VzXXidYXpYDDN
NNCV3TyJUvy+Y1okuJu5+H5hd5RHweEbBiW/KzLdnsY6NZ07IBG/xf2+4hewMMJeHhl2BeajaXqj
31jCev8G/8VCdsWl4MD4K2KMvLs+mk0AF1LIAWE9lQtDW0iQqEkFskx8LOosF1RncOZx6ZuunsvN
Cb1IfvuqqYgKh3X/uKWpJg3LbJl1ckviRaAtbH9DVgBbZABm2acLynBQUKG8YzHxnoB6tb8b7RtW
95vF4SVIL+RKETeUphCh58HEBBFs/zuvVfzg71l/xEO/2OqJ4Qizyt9Lqzn+NfrOtEJemVxH0kPg
cniZVxdlS7/9EdLNyb4vMKIe100+aX2/1qyz37M082mzjuiuUsz3OTw2Ci7IFork2H3TrmHXRG6k
edK9fEes5oPdwNHPzWBQez9jsILwE2XEKKcrzIg6bBqLmBK14Prt++T8wgZ5dokmiTgTBQbQscbg
/EZ+QCMZQhLl702Ibap9jVSSvtZmaTvYa5pDIw6oNvmqNGLI+gHpMJmAKSkLlXeDy+itZDUfI7/N
aMyk1MQmOpcEFi3rytUSUBQtHwfNV6dPe7dArfcIkbkuOXdgdK2SfGQ7VFgDk6XRfUgq0Ra2XCDy
SAZR0Jy8hAxLE1SYkWc7xgruoXYfqOYofhWeAWkXbffd44ZI/WhOD0G1sbby8n0FoTQ1JdS8wUfH
elkG+ewp8u4EAlRaF1GAMbGsIhFgMFxTFvFF5xxTXsHUXIWuQuT5stm0Du/r5n4ywz9kvAgsz+sK
CyxrPGdu8o7XAMFH1Yz3+lN05gIxHakYepH+BmfY+YV3Ct/iqid5NOqC4ShJh/JIbzqYJ4Q6LMQE
+6Y643TVVt8yGZ+gN8QLPzu629NI0zGY19GjwemPMa71gXiQSL3nMZ/pkqZQhzO+1tYKdziWJp5P
UAhS/XeKrK5e3zZRYBdwHjzFcvWap4FTugRE8+3bu7zwgVVWTB0zhDdrQ4Ri5fcUU8iQtAYZ2te5
xnj01ln2qWIOLKAqXAmdCAIXHTtTgiFhhtGi16XJHKBRvLRl81DxxZ/3ReCnYeBkJqe4C/0a0OYR
jeZ4izTZVT54nP1HK0O6pl6Te8B3htvkWKopBGoaAJjzy8VhBqPmpJn0mBvaK41++gzLbk+BcwFq
/BiwSZogR9vBQmomsnfYctVnYoYtQM8fW8Wy9z70qEoAWnu3Wg+5pFA8a0NI/9XsHR0ckaS7lrB0
F5MMKFg98TKxZKfKi+184B+7FwZ9UmUvidL3XbL0DziJM0ued393JtO895a6RcPCDGOhlRKnTumh
CWPscm1MaPU0W1VJwL2Xn0074wublt5zACZDJ+oS41FmSywMr53SALm8XUQBfqajOqtKF9uAvBrx
o/BuBjELEmuQsC2aSdqzO/nsy6KTpGJv0kgeis7fZ6NZBzVm1KifAX4jUJsEe0IfyHON/tyStFaa
DrVICJLoWfYxSD7GmA8WuDRm3GYvzMgTdmxqHrv5iHfeJ35S65yfJ58YP6iGptuMjOVPCjoB3oEc
sKuv0nmY3FNyoj4a+5BdEbItog81cZGeap75PqMMM9BQLe/mKmNHjooxiLwQvB0jZsZI8cn8xhTI
ms6i++tk7wGddp0+0VIEu3MOaq6hJ15pdvDSVCd1f3fS1WNMRWbKVBBNggzNQ6fUcl6INDdsJaRB
9+oJbR0zbdtIDuQzlGRT8fraS9sgt+iBXxcEIsJmzvR5Et2QIAkcekjo7r3ZwLAsY1mognyGAuJm
HAtz4PfmPzShjVmrI4FBe1PzWGhnSq6jevEdHEldOXGTTNBSTF+UNO9pv59USDd2YzZ8vzcr4PaJ
1/Xl7LaOJJXlrCLmclOwceWGRfr5Qw2+GfGxg45q8ElWLIFo89TP2mA+kSSvpdxTD0wh8tgCRIUx
mqjScVQP8kYJw2MlRx/doU44W+wB/neLaYzGYIVlSzW1jhnxudnRgJvs5juRRr1zTp5KzL7uXjeY
8m9MiBuo5sf/2tpmKnVRShgxrAKrjB8+eH2Bg6OFuwEDh0xlnO4aEL7I7WXBG6LzJwOlx+BOEfg4
HCa+cMcejzrA0OWIEfcBeeZy11WB7ltSDixLb8k8fZ3UecS8rwqDH0kKzMoSsowCpnvbHeXKIUYu
U+7Aj5zrkj/zSJWE+J5MhGtmwAXfVZI8g9pqFJtj7TN1PWTSYiLgfYv4wCOGeLUeJ8l8IgQECltr
G8yWKA+xij+dFYNUrYzayI5dUajnB4AxkIUkw6SXaNmw76VuL16cLMntSGwqPhPj6xL7ACt0rPZp
TU1uQ1WORrkM2COvUnxAqFH/n/DD2W2cjUgKBfPEuef0XYXN3+PpxwDsEaTkbd+aEy6QJwkKDY8n
K+rC6B3vQOgMyHfjCxeKshl66trfjiQlUnw0BimGKPVF6BryMnP7PjqR53nXPxMcFIsRp+FC+KWA
6M7dX6Xgkhl5NmbOYyjC3RYTJuuQYkmgnvtSnabG0yI0L2V04W6WwuuQmD1TMJqwp8hris2C/99e
cUJbwVFMtTbx2zQI+0+LcIpjWS4KGrGOtfFh5XJo3+0IHiCruwTrWGUi5h5Vq7C+c+JZe4eXX8mq
dCBqIrSds+ukBMPCxBwPjTAr/U3qpAtoLVksmz2TGoTDTTFHYswvm+o2iXC00dnxDuoZ3PqbBG60
Kpf2ruzVxCEoz625x1zSwTV0p8yG/1z1HebOyzyFPaeSUX6hg4W+bQLCP0kitQ+ttqFk2+8GP+5V
8GY+LW0tFahh0LaEC12fteAOQl5x7k4EBw+GJ2369cPrkZBcnMLin50/xgdqURfHO7DdAl7aZ4Zj
zzju+GyhMWK818B0nGlHrmHU/QqJyKvBvaMSRnuhC05t3XzhhiATs6NuldGY+n7TV4AVON9jP3j6
1I7uUxVLUB2Mie4k5NtYXSzJciZa71LTSRkzscv44goqI1OzB1GsJV1B2SqJTkF0QTNjzcyV+nIv
zDQXbn9tCtyvbVCjx0vO5EdLz/NnTvUdCuKjh/Za+64z0yhzAvPbx8dEqPaTj/3yi15H8D7GBiX8
6+75p+Obm8EJRL8q55dXnWWTbkRdGfxegSyOPvZ4w1JcXhxgAVEJJjuoVIpgycek68Znrze/M2LY
uhDe0xElHcQNKZl9o7W3mXqCyhlNiaWjfKy9T/julw5qLDBHACfPlqGKrrA22NrxpfgpS760TlXX
ymxz1vHnas5sYTNIjNMKkAW8Pcyx2zVRHEzlfzzByHlAdpfTPhPoWsspwEDA1mWU/joAkoHtVPtt
O5Geus5PwPagTXuE+kaiPFfMKcec7x/8eP6KVtnEalCqpVaXnokEpp0CgtpF4QhpEXqxeyN7YZj7
4nuCzH+pwzWwWHRk+MH/IvGAtN4RtkAfwSOGBX7dZ4WyzJQpWvvsEa7HTW8n+fez7ppW3nGNiep8
ap/YIJLx+O1F6IWL79HUj8pIAoCcfDG+Nce6+v+O8l1x5qjnrR+FZ+8z5xUAg8znEsMXEvwnLqkC
3VBI/E/nfMJKzhVjExMnPDNPnf4FknybH9TnLcDWdHf35uVbD5BzNs73GhJRgBRY701gKbUPOSI3
dW72BECUcnboFw2jLTAEQrUzhG/nqN/gqJAc71UajE/d6EfDXF3Uu4Ld7UaKvCOk6uOkEpyWJNMH
DBT/kR1JpbFISJBMejCmKCi9nYrf8hP+rrYiTWMDvi5Iq8KoPyKBZcJHOEtnitBq4Aj8sODRMNmv
QRlM66WHwkZMT099ZEz2lF1pquSGoLG46+IzP6K6nkYNLqEhjd1RI3Qj2JxvpahVw/uRopmAeR6j
xGzwRX1QofXLfjaDVQjaOlKrBJx4k3uLM3ARjhlS73+jml1WzGRc5akzeeHz8eVjGWLBFdU283ws
uT11IdlcU77nXveLa85pvIrCloW2Rs6V3KkfPmcUdgdjrY+OXB/mPt6lENMjn2R+36NkmvQG0cbF
cqDRrkZ7PUsNhM/miz7+ulGjAns4G2M3VKajK+9DCyqc9FHvtefozcTYq9wIvLsirvA2KqlVGCy8
Dt4VwjIlzBrRlD/0uI6tPjYZSKmnc7LSKvyyj+LnzTDWDwo0Q29/+vgSjee7+LU6c4aUe7uG+ZRY
Ghlt1RlDe3tAW0QjC3ntYtiIobG5c2upR8A1vt5F8fC9s85kzViaOePveOdlSIoWtYX6kpmXZw09
X4FPJQKQKIgXsur2TSqD87Ck/eL3JBKArM39KO7yhzxVMiwgDa+FTJlEJtGPU3xT2uYXDrD0raCE
y6R2Sz0v1kNmAFaPwBKLEm4C4h+pyMeY0jSc1TJBfe8RgutNgObt/y3HKAzHGUdkTPi2HNh1OcIr
gdb3xqQ+gdTPx2W1LpeT4JS0aSaNWbIzDydciasMyaJRRTiec2sqLaTmqQgrbQ7tR4f2mqzW72xT
BzOrMoznkUgTMvVrgihCxvHN2ZEILXsKmAP6BPgXVc1sz/CcummvqMgd7K4nG2QH7vkLIAEq53JV
TdjmjUwUwPsv3gnx/tJrwCWMU9tBhhS1KuKtWtfzX7V4AcEt8dhjg1Gsc1mW/PMaZf/2uncg33q9
1CnJKtCJxD5nsBy9JX2krRejIQ6yu7f2TgXOc3PV9rKjezc3WT1NQ5BZv1+zc2fQ2+9q47lLBqtI
roylNsZUyRYlOGc64SQQZ1wnKErois3vNb/waLEHaulbroiKnDHt6Ok719o5STeZ0vkfe3i/8w8V
sGc3Uj3Euxl8uGK68LvenXCf6jzWqcEG64do1lId1rqRmLY0grYvAiyH8KV8QrKkXOtJGq1npufj
IM1ZK0mXVvchKUPool0Ra2cQjL/pFdqC+16bFtcNxylyZlgxlavSRDUXf2Q0tRYuA47OARDtnRl3
BbOL+MjoD9HLW86kUNVUEHpP7A34+eh0Zps2zY4e0SV0+shRVgK27P1nXv0d0EFFNpnxzc/skyni
hft0FazUHE1dT3IO+vH6js5jlkmCUtSEKbZ6YeqkZnhdanb/ZSWcerEBzU3ZX3Y7j9NnWXiAJTGq
yX1w6CxLmieNuYs4N39i7iJg9HKAC9hNlDhagImuArGhvNW6CiOOMRE7HqaUBBSXUbyfIzpxs4Jw
SVF3EASFu3KQcLZOUzWRmaIuYzVzsCG6UMgvb8hcgWlBBV3DeFC4V6UAlQGFbvDGuLf+lNlN1u5b
sg8fAA/lZnHp1/xGOZQwSoUeQ+d9oIrQ6qP2PMC7v93Ny+95/JgAlMOCH5EwUE0t1qbkBB+TaAAr
luidWBTClFtuc9c97mzEzDTb683j2+iovuE5O8CdYGuoRSHXuaWr+OxeL3h+/O4CuEmFHiNEqL/H
4Q4Jvrpgj4RMxSz73mfCz89sDBZ+kHFbTI6AST0lERLvhSfGeaX17slOk6Rcl/qGSbaKDqUwGlgm
Ajc4H9f8bm2FFSerVbDGix4TNs8DIjvpyn1TTIqDdLd/+zkG3cZQe4R/M6DeEz1V6ZeKmXkGvkaU
+Ye2aq84sEnxCDwDG/69DCwxk8clV+IMZT558oklp68+3UvTgQ9wAjpVCYTVDuTZH3uQqsc8jEUT
YCTgeSOp/y8x9oPmTLOva/+uFuZasA3Sovkq8W6WpRdI5/5kq9qNIBX2F9XXHX7OzjKA0M8bQ/h8
FmrF118gfkg9z+yie/6zcUSNSCpCAc4c/5E/aTyMYD+fNqDrXWLvh/MPOZNiCub6niX3i0uAf1W3
Olan61FDtcxB/CSBlORPE2XNarZO/zLWzdNKmkYAN0s4dBZqmrHnti9aTXI9ETUhJ23LBN0e14ma
HLaLOnNQXryY0XONgi2GAU80wzw3rozEdaqI2ynBIz6LJdaAHe8AtkJhDdBsOLXFCwrJqOwIEObI
+IrVMGYpx3QtF681rxp6k/wi+kGCThHdYv23/sRmCUcCB7gSEMVGOt3oepf1lIYsWGzsagECvC1c
neEYlkljNicTMogPLHmwv2F/W+O/k3MxvRv4qeQIGXU73O9bfBp3MGrIrFAJ8ETa3DcdNNIicY4T
bg6sb3G/QuYIqUUtKS51bfeKNpRICwVzqtaDk6Kz3dH9LKp71KxW1IsfihUOD3EJTgNtnTiNYukX
35AnNZrpr0Mq6+Ovfzl/k4EXKL241UPeoSeJhl63daa2EhfuFISPL2q4b5o83h56YhUcZnIR7Iaz
wU9M7FvZC1iBc1CRr7xCJf70wtt6lGQbBDK4CkSzM650mNWDKeuJLe0e8BX+2N3+dUgZngunA1w6
CqQjD1yubMGqpbtgk4WXGNqsyCxOE/cLqWPWllZXjxVaoJ7u1wTebkUxWZGeUIJD3iWhBvi8BNE2
khwjlrpEMRfCr/5U70W/vHGXgJmY6WcvK0yfnL1xkeM0IBK1fy9g8dRiJbsuIIP684f9AEOYHrve
7Yf3K9kzJUorfhUqCuFSd6CfhuhCyINt0cbjqtCAy2V7RcJK3rfYWMOAIk3sI8bVuhLGu0JTSbyk
ztmH8GPGRLe+sXPxh0J2u3+pgsxticutNeZgvoyigKzvLg9YrJ+kN414LO3FR7CUlCyreZ4WiYgm
7lL2Bx1LuVwbVxNaWyFdgBRRWagG27i2GA/sVDzKMpOFTocAtD048kLtymaEQMP3GjuQlTHaYJWW
/t4enZcMgc/QsWsuGvMLYqks9JNfwbxd8DnXvtrI0kRoBzCDMo6Pb6NFJgEVEQ/ZmeiATpR9RyNG
WFZzCDdCqBgCUe+o40pnDZnjhN7ebNsTsjT77SVrcxTb99mLS/X8jhWzq3QTondngLxzyaMDHOM1
IVeXT/jaKI40eTKiA1UYBxuhWiYOkr1TbxlIAZMWQVdeWCMjUB9ulaM7RjABUh4HGbLlbdEsWiA8
emcwsIgBhzpjAnyNVHyB/kI6jVguV3s5JSwsf/hn/oW08bHsx0vkj9fju1Ha3pFuNL7I0b7Aonjm
wccJFuVmJJUgUrYwSrLV6LWMUAS6ztG0q7ur4Y9+8hETaXVB81lkoPu4+lZ/R8QWBpWnsiD5TgxC
UIbOR21XRKSp+Y6/ynHbRNaJFrYB65xee2fDeDi7jNNI3NQ7UuDGompi/Dm8DXzV/bobxKvHQuhe
96I5iLj7hDRzxtqAId6sKNo3KRmo4TcbqWhcBeaqXWvV4gNVEds6CTYDkUmr61VJSVwDQtG15e4b
J9P27aazq8acgsqbZtO8rEbL4nczzwabXX3lrWFUND1Wzh2dFxZ/Q6sGZcDlFhUdAMJgcKE6aRq/
0i3mlz+70cuglsvxc1ifDjOTSqNMV44rHCH+AnfSgpZ0In+OAKVPXm2iYkEhWLplQw6JqT9EEWw+
8WnwCieIMA5EoqHpH5cLcPHCxZQ8Upx8GfkaR3Eh9ePGOJh2L8PTyR1ePRB+1CXl2Tp5ExYVwJj2
ZMYq3c01rt9vZa2C4BwtAfeRmhFaeb/uyb9TRMN9HfTSSMSu1edsdjyRmoqDByL7SP83A1GmTx2b
TqxOEmUeTOjJsWsvWqy+isISwXdz/EWC6E/1RRUgoh5IDWJVblj7z5hRGyEmRtXGfYvcHs/fwT9h
GXS86HTd+Ls58iE9fjRL8O7erqPiX5bJ1HqY8t3FOzjE/JR6m0j7qtOmuXfUmx5/ZNdrtZNiBvbm
RMRVSQ4DV97LCyopQyih+7WrEzG+e1lxEYyl1TQDlM/uTCq2A0mz/+oOeW1Zfewp0ZqGM4SYEL36
n3SCQjeWRGeXYaQD+RqrRX7PQMBZc41d3nT/A3aJSzvDY0nC5dmeETKZipfzJ4TOm7KAJeZZ7Nww
GwYYOTTLio7L2mB7nyl6CKI/K11wGob9up6vsc/Pp63Zkc6LW+9y1gYj2PtNfzpqsVqLEdkEMBUH
CrebeEPFYaHXI35H86NuPZyjCYiUHEYgBMc7z4Ex8HhL8f44kU8ohPSqkRlaaSdQNLntEEobZfIz
cmRZ07nc9fIZ4QFzMw7nOabuFbz0U/hQkdi8M8aK4uWzOZwmG/friJyVeGJQGzKnedfeFx+y5Vq/
MsuR6ES0ndYRXhToGsVbZ3BfseClHJQUw5T4z46jc5A58brIT8tUyFtpgIQ2O28qeWTl4AniCKAC
Yl856g9lSlFqyMgi5rHG7/mvnzzfsS8ce+IMiI0nIrxpPyvKQ0ViNuiphCQsrB/aXceOCbt2TLW3
yaaSHvxJ+nzSMXFUNKJkvPC+098EQiI989FTJJ4TaiTVszu0jNxMzkt/XWryoavdE+KIOBT26OMY
f4gD5UGFQZlD3lhgqetHGSqT5HyTzhUu2VwE9S5D9c/k8qx1cMrYS7O1+R6QeIj8ZhQ3kTEFoK9k
G4GZ+EdLBP3O0s6Cueg1XkLRxt25iHQ6dd/cuy08pBqNpwQ11J21piiXJs3wgytk3RUZbbTVTtoO
X4rt2Fh7KLjGGa3uzBFtEXzghA3ttG6AZs2FKbJ0CIDotCz/PIsJ4dzdPdQCeTxUJIoiJ/aJGmdt
+mvJKFjQ5AFfucf4hIWpWEp9x7B3z1BeY3RpVkxKX91qUC4gUvPsVtjTuc+eTipDi8zf8Gv/P7Cy
i/26NSqNC61bASufVuVnElFhcsiA9qNpQsxfKa6AgnIxxDqwa25ilR7nZPv0tSi3427eszx0FRW1
74wzfZhZTZ1OO184cZ50YCN4uHmQi4SgpR+yh0daU24IJeI1EMdMdGUsEz3cNdwGzL4RJ0W78XYD
/080aYOKiq2eT2SK8GbCr4lsb9UDmDYs0igmCLmJMzwVnHX2fd3FAxKj2L5bCkJDeOEA/CU1VkRY
05GunOnk6HWl160RyI3muNmNKyZ+la3xyZK8JzsVFgL5SJ2XDvFVUF+nUYKRWP7S/eA6OJYwurLz
+KAhgk31dR5iy3yEdE/CUOxu5ijKKGPibI+cKejq0QZDoHg1cPRM5stHRaiXrt7OagSr3lqjZIkb
goeEIpY9gCv4/CHBBwS7+jwe/RkQsF1bOJy3S8/XrQdmjDpZbEpg19GrS3CyXITWp3hMkNAtYtGd
21OZ/kPwIIGEp/cIi4nC5eQE3Z7N5KBDCdSNV81IjMY4pUtvyd/fD0zkI5haK6L0y+MpaIEo/AG2
CZL0t3AKLSEvwlv6KNAMkoleYn9DLjuPwvGrljc7H0QZ0K7QOjXd013O7jYLoX6tjCeTxA/57N9h
rLgEKdQpqf26BD85puvLDPapq+ArBAIpFvyAjONXtgMEwApkXBR6PrUsd8vt5yTRwhnXZagzc6V/
NQVHdV1miQau5ng1Mlcu+EuxEtr9CEJLOtea3Y1wj8up65ihGCqd/3R6xEohQPsWwMwzXCC+wiXj
WCyJLgqwu0PPXjDcNg/3glDp/HUMyzE6BjA3Fhuq7Ms34N+aN4VJmJ80WwwC6BNpY2q7nJ1E1wtz
AvKJGwj9cvgUfh3SW5d4z+Snw6Qhv7YDmkIwBLqW++YhCdruSXjY9syA0FIQa2M50iVBBoFgemxu
fTDeX/H0//cQMX1S6NoUhCT1Q0Pcu20jGr363Os3eqKbki+HYR2I2fA4WcfEAQ2WH39En/gev+QH
wwKH8GdA/zvaD3LJMPb0l/JPWK05lGRV49eJfi8yoXePiVhvyAjkKhAjcH9tUH62mLi1AjDB2VBJ
OMOaYKYeIxdtC+SCl1S7wzU8NQA6uac8MxMz0zCVhZfq9CIw+qF0FoWZ3qLkOoRYapxn/Qa2lvsi
h7d2GBPutZ3NJFHIyjRX6iu3ehi3MlGys/ztSrx0PZNofJjuZRqUbJ4fb+u8INT2o+v9UrwDL62Y
XCkFpfV5Z5LJ5NG2oDx0cldfBWM9QEyFHWCXhcDQA8y/olRWreU5JTLEWuNDs2J2skFKdkh6JRcZ
CLuQssI23lLtqGLO3KA5daLxw1+SVNR8sTd0u4uofuFRadO0VD7jLn6qsJyin9KeEz8WOkZcox/Z
gWH54AE8dkVHBj9q7yj5fvafsKwgrvkpOHeGJgkhGN9wc0SaLmsdC/AgkcqGuEriuuW75lgUL4pe
gxoGujs839CBDkIGBK8U+Lq4C+p3LtHCQd5d6WyCB1EuVNEBVkQNGvVE7HkkHgE6o17i1c4/jNow
uxONhWr8YivJGrZhuKP261DTMuxRM47axKCJzbGvwxaN8XfY2NBWDAJ4eLVe6z6tKNx8kQvgEk6z
HHecRD4PBGTrbQLq8xeLmWZQAhA5Qr7O9JDw/4K8l6Ad+9dvSBJ6yM2TbymLU7fgNyFgmMcC1ao6
f3GWvVWkXsqpYWGtNSlE8IDOPdzx5AYg5N7W0pgcz7cjTbhw01aHZROGWxiZhwn7tDlURQ0tNapn
HYGQ8mp6YvK9CG1BZ2skXKqCemaGYFp0nY4hCr6GA9JT7waqRgyqIQz7C8WPMmTT61ylPwOize33
JFGM8fn9LU8UxffE3edatDG40s1RyEM2QWeIDNXgwxAabpn3NhQl5r0O8irV4aR2Zhibp/CjX84X
agAPctpki62Xald7HfGkH7a3AjhrBXJviv2ijGJ27w7W/ZdrEmqJBBAMr2bS5Gr9GvH4bihsGY2h
8QN3Jwf4Fi/CvmIdUPlQEMBf+1oUK/F2oO+y7Oc+PeKxArEBJEvcYreqX1t7oQIPsT4tUI324LpS
C0+k+NQtLdqcg+F4V6J6IzQ8sf/gMfICSS5iOAmz4R3cqVRPESwO4jBIh/rJ5iypb9o0Gf17G4VL
szfg853RW2XrrrU+bqYhcFUumGmwKCcjPdv16PhT1xsaVkKgxRF7QBtN9lJtz7P7b5bMfTDcNKTt
2VhLaIQQpA5u//Yq894aBWZasMS97QPcrVgjUAbTJovD0zpfH/ejp1VbwvcHkBgCCCcr/aCgSDPg
9qdOZAiQfUfAugdXDBW1Us8O+23wilOrwQr9qzOtj90I818XTayaAavD9c0PQpv07hSn/103NTed
0LtfsLKgsX6EAcguXOmO9jcQCz4++WrEZHQv0Kc7i6HRxiGDKjRASAIf7B0PWO+eQHyV/3gN0dhE
8qpc37Kxp1EZpSxCoy7D3Lw4qXqwF4gkQQjolbtVyYML7TLgZbc1LpF6eaLsXbJ9+bsKVihn+6BB
3KG5WUht/p5jad2nvdC/bnWJvMUkAhnQnB82vkIcs5FDCVcfSWSFOSv7mgKyeW6aomcPHVAwrCEF
d3rZsJ0yn+sHfk27ApOcsM9YpzA3zB83nHJClr9n2Srhj/kyCoyp55r0rSMLyxd1TMgBTEvPLs4A
AsxjON9Bc5ERh84kE50xHXAB4r09og9oIkRuBZc8h/V6tlziD7FoCW4YMJRNkByMzJqMGBhr4uJG
OynJiyIu47B6fvP4fqcQlMuKvnQIt/H8tnCWUSk+wQaJCxF/9lbshbktG/6VT5Wf3Kvg3Y7eXP3c
tdlwXUL3NqHJAv3GCmwNLoIltOmt6Dn+u2cGM8Uslk6J6YWYfc0YuDIGIAqG8Kijkv/9UYybGY5D
CKbbci5+QkO7tvdUe6hSXOynexWxQW0NzfViuTiTDEqmqz5yuTUHWIkvhZEOQLUEMqv5vvyC6MaB
nmGpVcV5K7Jvf3KgNJUWfrOxjz7Ru+4tZfdVvJYwDqk6J9QcTXR4AFYXKK0Z604WVyPH1YbjCF6x
LagT0yNAxo69s0sdZO0fkzOV4jpbJKlGBwXFzrsc39hGCPWyb2MQq4QMo+IXXkMq3n9RF8g1kP+f
UqU0mH+kRx+EAz3vHkEEwuDSfuMheBy0SpFOeIeWPN/+GrFUJgMFYrx1/FtsZNUiJZxtUrpyvVCj
mj8fzjnvpVQDByN6MmY1drHPKW3Ks2RwfD9MPLoNnabIF88dn/bK/biE9jtEjMqCZltORehbRuPY
AWPomsEfHSqGljo2x+SktX8WgX26Gkj2Iw387ezxIx0w/pzSN6xv00OL/4LOQc21j4Nav4zqW87M
ywsp+8tQ2qiu5DJKQYGQtd1CTFqqqpluD1YtNsSaLSaD4l4quZHOQ8/Ks2hPbligBPzaii8rGwkp
7IZdjnAY+BLYzYXKBxS0A0sTrLW84Y/A0KL4UhuhJL/tkiMMVrC7D+A65JaM7z7SLiNtCpylcvhl
BMsizE0NXywOLPdHaSXN7w6UrZVi3EE2pARrmNtzMMFNkg/IAaH+kDEYfko1d7jl2P6IVipJFYU/
LTGW4paKsl1g7Iw0riB2QlhIxzqH/aRhXcyHFRi5BlC4Eh4JFGlLDDsVBdPm5Iha97jQ3JJc0aHj
QQIg4VSodCOIe/EqpA1d1mtlLc71+DnXHjPAxuHQJ72Uz4d5tS4mWw/kSIs4Fe69fcNjU7SsfFqM
43TGQN7Lj+v9c67rODk7sodOkb2ocjT3zhgotum/9sH51rFPMW1Pap2vtR+BnRMAqODV2ADzQ2uB
iz1AeuTWfHndfXBVjDXP8/NsS7T/BA+YrGzPN/izi0L/GV0Baz4NfelFkU09cdmY0/k9HISGhcK2
64sRxXqG7B1rJBdGQijO9h+sQ38UA6ekGe9eCNa+KQ3ci7DPZc0/pBMsoQCJ1+DCIyIvozf0xg/D
4blrtKuJJlEy+X7AKrOtap0woS06DHf64JK3KlDY1Ht6fdMtUZUrKFpPm/EGKQ3/Edz6Yncakv7m
sAc+U53VhFe9+KfCT/pZ+FAaxztAnxAXIjQCoFhtN89j3+OoGfJQJQjbzNGyZ6bskJhxsKWIhmoy
zzh4eA2tVWUX5OdXu4upBCIY+kYxg/lRdlyx4gn7GdUefVkjC1cBSOci4DWl8vCbMoI2u8xOE7CD
KQ7C57Bm22N44CmGOrOVxZtj92EBALAHcilwLYthdy5ubk7H9K+tFIVfFzdCKbgrrVH5IZ6kK1Il
9ax/NHcTbvxX4rrIxCvpJaQ+GXCiUSAf49PIuH8ea4iRgs9zpAzw3WKNXRIGiZ5CsqqN2V7/bGR7
XhV8jzsHwfV/ZnfsKVZ0tKSm4pvP5wzGC7AK79yh+QOweP1CrhhW6QQg3EHHDvgQiKx0iZ7SdBlX
vsKVsuWaFsT1QLh9b92jN2RLPL/6qTgHAbvdv21EHDLIZfisEqLTl94vy0/enkzrF1gFQa/B4+Nl
pWPa5spYxhrVGyDEzdrf7zMRRcgvjOhBi8LcA2MTPbXnJB1xDa//NHYddl24Z8epN3SMyU5ae+kz
qcybgfHRuwhgUb+Mf6+NSvjkuJQdy6gLvYhaiQ8WTxz4vzyQdxCNkBfr50e/t44guq/686ROGdi5
/IlOxEpvGffLB9jgYe+PZ4BIUUuEDO4T1Ai7lL5KwOX1bvnkOU33881KdPEgo0wP7ZC2mD23n/AR
PfaJ1eSqZo1+9TXT9QHFsrP20s2Jf76aFucr+Hzs+KUsmdqlL1DgHfotY71A8NaORFvu+CYBYess
FlmMuzIdmIJzc4aKKlLSFoknxY3JwKQLVUr7iQw1OuscEyHLBo8/p2RWRgIHqUbnWJra/6afOcLu
kzGY69k4pLNpqLQZ/uniwiNe+60q/r973OTmBQMMH9wv0pNKJ+AKeg2aRSafHDa0Fo3TYfeiccQW
ERK7baLQLU7I0iUZwu9yAc5ko2ThhD6KP2TGP0jgNb6xRFmH7/J5giZEdOD/gOd1FV1HDP8aLcN7
yDZn6qG/uOhy+C2jubfeN9ffVA5eA6nhaUtD7rmHy2Dd3+Zrkr8rHOTv0nnGkzMyx/n7bK49RNnS
4Gs1noD+bj/8hEyBP83wj0RkLRocxm1QmCaNoWFqotB9PAJ0wyNlesFDyoU8/5k0tgAHz682+SBr
tpP6N+CPx92iDvrGOzCKMPhFVAToS44sQP+KUe/OzSP+SAnY0XsnLz9Fh5EexdtCwvaU6ycoYIej
76odP08y7ih01uYoMgR2Qia7S4M+Y6dC9ePdNW6zrIGmYx3RNdshEP1H/ziH7p2WeKIcW31SR4RY
qPQ/GR6cU3Yzkz1Ni47OE2L0iHYrJfiqhQxIjAoRUgzPVzj/XvErmz2WirHH2A34KuwQvoY8KzGt
B5QU1wWIFTeMwrdPaqpDxd6mRlmWE1moMMpJ6VQeoQYNlc4CHSvIcBE7gy7mGXRUYes9ndlrUitS
Sb+iaRkTsQEydyTRfZQyny63hAkm2KpudXeDNqcOjdyWHMA+f9vkGvAEnItJkYQjlwbU2/jxVFRm
Nf6RRSfwR5P5G5QwClrG3JbUds4QnN+u0HxpwuFyum6KZ/6660GRGLgXUT5kC8kw//3PFGJcDWvr
ojf65O46lCAy+7MOg7Yh2Oi69Po079hpkAQZYWPDMLS/yUYFreTK09zvGkdLnnxsgk3gEOg9BN//
h/oO3cXl0A42RWK7jaPXmZmYat8jQkdgkV+31Bb/MnMGibfM63bUvGLAB5lMJBLZ/+QOsLOD7HaH
zPATOJ+/X6WKlnKdc1dzg9aeTHBC2SNlwTygqdujn9rWbCuVQapugv/ws+jbN1QgDF731QMKu9TA
s68Ww6/c8/bE1l2/vVFrp1xPmi5WFYzT2sWCG3/jzz6zktFDXIKYrVb/Xq4Gsc7WrNmKN/uTaISW
M+B/DGyvffRaXTfPYWwylO4XfGIL6b1MMuMUfcEx/imXOqhaE91RgEZ0QJK4YaPKcV29XSODumhw
ewaylKv4kko5/lyBzbRdARDCjro00eQkRPdeoWxgx6zBUT5MMSs0AkjtXpgfLNi5bJje3qgepSMR
QoyJr8QKG6M4vlcBmMVzQfvC0aO7dWSvdZQ0GNhGVJJ5FIS5eb1/UrjpPDmKY/4a7pUOoaE/o/9f
QjzMY/KqKZXS6tlgIj1h+tWMMmU/LIVlDIKZCZY79mb0Rsch5eJVWTdA1bB3AQV5DIGGh5pWalo/
N8qBTGovIKHRttShUEIBR7gwXM861ZayHuq3wudSMwfiXQnkaktEWRfaC8Ui0RJ7EtvwIqohXSfg
DTl3/Wbwd5XLbxdhlDS9HtucfUN9SjsFwu8x8j2b4gghdQC5d7LaUtICyAws98MakwjFaxDBpfIZ
f9LS7QXjptoYJ/3UzeP1rkQFukCSniuEAoFyj9MZ3cuAlfiZxGRXwlhFf+adk8Vwkekz1Bv9eq6Z
fRSIruEBFFSKY9UZqouV+LaTy294BhhGNwfO8sJr66ijlZxhuUWBGfM6WOhpKr9r3N56bq5BE3+v
DDV51yM4nZeyMUan3PvCECOryZqJ3uLGItBHVe2tvvIUdWQK083tzxQCXaUNTmxC1dS9iKVnrp5t
xspd4/LeOSUoJOpF41iFug50m1d5F2k73ef2cr+QeJuFi9rQqaaHpRuxdeeHslSzM3I/ACkIiTCM
2YMeVZpxfjD0jsOMQ1/WNWc5FKrzunzqe0aKPzrP7AfiVUcN7iDXbtkhsEkUUBcyZ75VAltmEyUP
X0ynMMh+OGX9TtJ8lJSjEhncuLJ8g8cpCKZ8DwtrX2ubsnRLAI+yEP+YqdZFEx6tTMhq5ebZIq4+
UMHK/PvqW38J5RbtRcrtdCQuE71EDqY2hggFzSet6F5/Z2NxWG9DAfyPovDEeDv1DYxvU3F+Ibue
3+sstfn3VZxG3bKamy5MujUG9O701p75+aYYbPWquOV7Lx0vLD+kX7pWhhTSFL+PTp6yB0U96itW
359jbxJS43NZ7GprYyLO8BjtVuZap07X8oLvyJp4oASMulBvGD2oS99zED9+AHS/rsi4Rm+IJDmS
3WZhWCau4WHzeAHBXrni6Nke3PR5voyyDSd2gKY22bogX6TSesWrD9qa7IR0wNIxMH7CBIehKEe6
OwbubYBN33tHz7MRC3j4FGMEaEU2IvPVxZye7exO3C8YLFhhb2lbTifrdN+dnF/D4/Q6eRJj27Rr
RHuuTC+DLP022SKu2ENcMyAdi6gUT9rYxAqlGuDRCBpLQd2CVpr51RKA3B0al1RZREb6ZTlEfF8H
iw4Axdo/GPRO37Bh9SUkRkNWp1mTTp6PLuu9WBclWIK3LqcqlXN4z9VGA1tU3vZ99DkNvUSzd78z
wLy6sdt5kBJn/LOz0LBuVgdrZMT/LPmRwKULQQXoFM2Yo0oIuPv+QIX+bXvAtRJJDwQP5SAlhq0k
xHhP6nFJ80GErSVDFox/z4WM8ZdM1AkXVPra1gZg1jmAlkeINu8I4a349RDRtgwXPe+9L0AVPmyv
bgxckzxoJLuDFkd5B7BuMqxX0xK4NjoRin8VGUSyK/Cy4BLqP9VJ2Od3bDwSXOYlaYNOq+xtA1gD
XwgVJQTFiNQ94hPx4QfZl6SiR8Ww4QsE/qs9hhNIekkrCuFgrwLnWIBX6iRUkJocFuw8CQ85DnFj
u2XrRZqAzuXAjPw9HQBR+WosKd7FZnJKCGUSdBRONFqkLWe3Fn6lZzRbJBaMKvVGZ8PfvZv1vT2C
cYZwE8VKoPYKXkaVrmX3rZenwWbXDKYHEtaH4Q/PpvBbGuzPvwzU0E1LYGnT3DGtJy3txqtENkXK
8lLln1Lz9BjVo6J1gFqYnmlhgQZ6sGj0kj/Hol6nKV1sH5sqYImHfxh7lOFFwkHMc9zg5pkK6GF8
pu+zRVe4WAZcWIDgv+4fW3l93UxAqgyHy+MiDHEqFzX7fdclgFooec9yFwRYIWUBmEgwH0hzmzTP
DXxdHvZn6I25STs3Tg76weEUzdxnxfhnWrWgBSD71a9IKVu6P92oLhbu2bl8CJGjbwC79CwEqGA1
yugLSEFYQheVmd0FArVgEGg9fCsC2uaDmNxg/ROh/1Ya3Ez/SI1QnufVYJ1bCrnjDfPSk2XYfI3i
d7CQegz0aF/GVOiWm83yu9x5f4X804X3z/8k1T1LnSYhiou2HKLrUbv5hpYJ/d13F7hJoIUu99/q
NswqzCHeZzphaskSHZZxV8LjES1wZKiibuesIH9BFFQ2nDs2Kj629qarJ8BbwNe4rnkTzZh9Is2c
3FXMvOGuhqAWRWS3SYafkA96UdW3V6mirI79BdkQQ5S65VWuVrOrHbZZuzEJCllcM/lucUesnTvg
3C3Zte7+BTyFJlcLy0W2PjIitZkVNnGDE4ima5vnFecPwR7jtz9AXdUJX2+BblYKXpB+3734S+Ct
VB/pylNFiAWlGI/IzBmNeOC6nj6GEjNbEN2wcGSA0AHiZKijkkC3TBjBClGVbU0GkAnnR0Gz1f1u
8pqfyeXIAslw75IMF0Qv6U878qWLysDYC6qt/6weOoC9hs9/eZ2pDd6FrP99kK3KlYED/o225uXK
Xz77NRfwmZHLYJF8ed66z/iEp4TGjYFeHZl6hfJFybo7iFWVWoVTbDgdRsQrD35lXqAJD8qVxWQe
YM1kJzYl6fZFHAII3fVMFTwbgXDa4hdvQpNZHC65CDNBS4yl5wSUKHs0JiIJJ+yLEKqs4cxes1qM
cLv/6v95cBDxS7jB3iq549277cIdRJDMlNAhwrCRsoY47szO221528ARYO/hH9YmgUoL1RnUGWdW
e9tC35xRChEg5NJW5fsnXrBYSh+/I2BBbFYekezv4bNcw8nX+yRoybxv7iL3z33kQNdARU9ixR+x
B33Cxh+suvmcLnmCOcq7o2opXiVthV8vWmW50eWE0NizgDOzCM+mW+Nz6UxVpMyyolqjBw+yDx2Y
xIfdz/4/7xGuAZqURAaBa/wLXl5+ufbi0FlwZp72WldsOv1/IErCWIacB+joxF9Dvdbek3rosEoD
tqW6SWq8Hv8/w4rRM0M6xYT5eMYiQOmSPn51VLZ2MIEhtkWouDDAoUnvjW1ORJx1LWokrUW8ETwo
I21CT/DZGFjiaWZ4JCm7RUTqPlyV08kcuJLyzVr2L65W1hz66afNqaB2TCB5srvZ1srfIthyghPN
7wh6ytqPTx+g3Wy7eKJ4H/vAjOM2qDU3pY+C/rtCR5ZxTL7Wiq9QDX40sjmlTCty3uVMPxCAb8ZA
aAKcIdRL3NGxbr7Zoa1EX3mSa6kJPnmuoaVK4ADrrzm1dTYwyQU+e18bhaPMPNtxR5R7A/ODyXRz
rT58t8G7ethPOTe72/8Fvd6CcMQ8Rwfx47z9rmO3cz2Ohlnu24Mo8qrZ+zmyB/vgBVnqLn+znaD0
eBHVhLiLQ+1lT4gqZQCOJai98ssplSqwCdVK9BvNFpbN/0wMLYgL0EE+dc7LYkJbbSyHmPFdvL05
sv6ArB83Nh1bGkHSQizoLsd/J431EhwOs66Lj8p/9es2td56klXXlDquxk+wpyRFJYLM5JUdpqIS
YJHEgbrjA/uxlD2hE24N4FdWnwDNXiLPQk7HiTHu0WEL2D2GWFFFV1ytukCgwDhZA3lzZ/lkxbcx
V4JtswcMwQe/hLPzDUmdAqiDrhDESJcr+OzhcF16xfb8L25JmS2y0VDT+ZfFkBphBMZpmG/y9U7o
F25YJTBi+HYSxHZKWZVkqglPs8/oOTj5753Yt4cGE/pScz3/KeMqXFxRvCxBOYOon0HfVCOMsJ9s
Qv/DgWR3FiLW1j/u47syYFsPfJjzXnSSrSGhgzQoReyIOD0ZXsRDzcEWrm+E0V/c9F71iLh7h+be
Ee6oWzWH3sNbJIdqnlumV01dYzItLxQB8liwzrVBorBITgF6Gqpfk4GE4RgVB9tK7QaZ02p3g3HJ
Ky1YpG7Q05Vuc4XDqie/BqevKfG7SZK0Iby2lFELCpp3789/quEi+GeymL8/se9XwDgdUVVRAzK+
N/mK1dbBquzzwzFyzHwWB0xgQ755oVCumvycdxm84yB738Z39iArIkWPIHqB7a7aLy8BTEZPM/9L
PYShTLVhyPOrfEXHioFxyHcDjyzhDTX1ERQvY/ER9oi2AuJxwAPnYYMPR9ZBGjn+0bm9kOPgml0c
6CTpvytFH0BqeI1bRnrmMbcR/mfm1ohYpU5sLScjXEzYLA5DQlfTUeKvlgxVO11XffSKPe+9qPnb
8hzaBg83VlxOc7iDqayUJXTURSczY1b02TKiEiY5X1hYyuuqFeo1MY47ucUySV7bOMsIcQAIAsIJ
FD+sCOw/zqKXzIeQs4RYDEnn0oorGKpph+YnVBAw5t2/9CBY6RLO2DudML4KbyOeM5le5ZZg6p6N
/ba7gVlhfN3c/uaFU3p7i5Y0HTb2TSSmvSFldVtt48ajfVZjmzp2plOVvFFynZxa4SEnriFizk6C
wQ01ho60MXdhAG3l0V9lWHA7VVzWYYZK8bfuHtQEEuVS7SQ6pvA7ZnCHLPemNYwWDqxFgZJMxb2x
tr8mpMjIIuxP32Bkqz1dEmDKGsUNS7a5HkFNA8Jl8JOLukYHm8nRNggaxrG1HsSoVgBTb1JEUs8T
y5kScBsphQ2/JbI7vwT5erGE5rbXFDbiFocMHa9NI4GsNnr3/KFFgCZgIgqjHc0zsI5BnlWW1Gpj
3P5/qtj4//XA8HefwcmGGKml8q27W2/AeMh6Biu5OqpjgqEPVX1iDsN9NCcEGxbTXajVXQi3JeZl
aT29gIzg9d24WKE39JN4Y14kEnfmYWicvCalPE3s4WFwR9GckBC82pdp8vUZXPQ0IQ9DwUcou0rA
yB/65e5doaFPUJVaGh+hfcpcPe5BQcr2zAP2H/xeT9lKZnhGsue3E18/uyzrBM9K1KipOK+diw8z
WFtt7RxQhqYBA4n7A6OP8i4g0zsn2BGz/jJy5PF30cSBuB8ae9FRPoOERlDmXA08yxIOdVTVzZRL
af4/5dQmQVeYl0pBVhCNG7ZSqUxuJL0nDaua0kAo5tm6naaIaMT+yfy6AjJJKB25jowavuhqnCuf
RfUIB+xHxAr1CwzQ61G616bz86ohNXEqYQ7g1Rqhf6Yf3hwCXNgdZ6P+rGYV1as1J0MMEabXd5aN
DW9aHuzsLoHHFXFuAM3j3UzL8DR6Mu6vQbv5/r2uGVIwylhA8EfC8F8rvS//czbwl/7w8btGcxHb
9M+JTmuG6BFzQ6PsKptXnHdzVZ81KFtlzi9RbO+Br6paqhHHV1WzUvvbzM03yWVGqoIb28nKev8X
5g007pGp2peAvOqw1lMc+E8MaUWBnBrX2dBCBLfRE+NkhYh+rpxVV5Gwk9S1pI45YaoiDFTKn+6n
M3mULHnOgR1hXmA30KJDUgAG5rwKSLVDbSNEa3f7+vhrb64KAK9XzHLpMfMajzoXHM3OwJ4AQp0T
P+eDfLGGJ5OUHiVV1DuNo9Qk33GSqLqVax3Rzj32soSg9yaNBvw+B2OyEXAXpebJ5Jf68jTbOEmx
ZSf/X0iyEiOsCizIntswjDuxTeOws2BNYRCjF3TEbcpvyZz8dIY+zhQKV09AXES6L3gKp8TwkezR
SPygTQUzCxLxNuteVo5I7dC6k/dd92O5lxQib5P3d3iRxxoVL8EKCPP85B9v5wrnKKGxwvsVFQkj
lRgRcMRm7eM0pjcJXoM8rHWUglQAAl2kSjYaPbt9da4d0trGrnjRrsD9f+RTYRlTzFJgN2ztbWgH
OLB2ANqE2f4PtRDFUuyfcqBBdgzE4q1WZwFIOUhDRnTYK7/9213UuSAGLYGSewJbn/P4FmCNm1TH
WvKubssi41XrprFTvwF2bHmXvEzdC8QmKz6+8rhrdlGzOXYztduB2wY3rCIUwM2obU89FN15wgfH
/HkxYD9mQrvqSEYwZnruHiEzdgRogf7kqoQ6cHzxpYuLw7jNGwv8rS+wPIWTh4QACWFY6cdIGtzy
mll1W99kUhV6ciU7/cL5j3slbVpmKbNcJBqk10953xH1RqNarotXWDOENQuvtaf4F2rmqJC275+w
QnPCXg1IDLXhBw4bJHsf9U813mp8K9dYGg7dJ0Wpu7fe1LEwRXo7oEjXrX/ZkhulwOyEycxmAMdB
jkrs2LCH+Rnkl8t/8Nc2M3/JyKNmvP7B3uT+HvdTZdV0xwdUOvzEoh53xOmJZpKD1ptTQoDXJ60z
eRaqPv9l7481CIOGxrcUovc3jfUEMNrEJL4KAA0xZbVCKtoQQxLTKbyj85XtF/FrSkFkeyzef5oF
0wlKF4W5MRgHFjHQd8H7IqB3jVmCyUhaF6jURVOfhH5bPtFolHTS2oenp/zPghilwnFQ3gwDiVby
4dpgtmAzzZZ4JD4GvE3tjhB6h08zE0Zkig7/w7iHMmRXr0u51SrUbeiZJfbxtOD5R4MWHROxSu7j
F9AJfpHgnziD6FXSYGLPUilbA5hsWFsllDTr1IQ+pxtJZf7/mgMiuGwjHLYowYBBgfoGqjD65nrM
OKnj/7q4IC2DC4Cj1HVW/Z8hNnOQcuNfuqSN1J48T6CtDcXx4meP+LWsMdAYd2+fgMKPnF+bZqCM
mfgppRjWZOwfBb5uIjS/OtmvyhRZkBSLlAiJC93o9aN6jBXR3TwqPQIYog5ywdTM5C6hSOabpQJf
hIvlg8C229UfcTrF8YotOvFBt3/63OsrRSHB6mL4IdpVHGdSPCAGaID2FHfpUsIMHFOyYiY9Wqi/
flcV1r9EUk6XAM7m1bO5F57OipCqiWDDdy7n8Wd/AV+A4lISqPaziSSH8E8rxEUvbfTWEmCP6Xu8
l9xB0+UDIRq3SkHmcpuEDCLdSRcE3oljNJIAaD1B8ONzXiI2+EndpOUKrx/9yVsg8u8rFPavghgz
Xlucn4rKI/jtsPirVEzLAAr2XamxJMT9/d3/lpFZJr1c8ZWoGPa+zc4i/i/tzyEevJliHWh3EoRe
6P8433UgM8QmFkhjWHYYMKFL8w66NEDiXWVvgBaOyp/JVscuWl7o0Fp9jEl/OGmK8kkUW7cy8d8I
6Z9TDd0BlEEYP2B3kZH99D+Onghh9BIq44xvXzsmEnonohNbRDghZ2QK9v6qSXOqQnUflGFC5Fcz
w7a4eU2h7YpGNX6wLH8YHuVUPux6I7gx9pcnFaxENEjILdtegQC0cfXHt9+fQ+CYxNDewAJnHbor
wiHLZeS5M//yR7cT6r/DOUdIGUWc81fSQbiqLDn1r07l1QFWFvB0ADy5UdK5YkV9e2+fi+jgmuiO
GuE0TrnhAbAecs746WIjMgTdiMYnk64UQJIf6v/4meTJyHHsItMHOUIsPoanGQRo7n4U5jM/faow
wT17r28E+v2MT3CnpRBA1+QwtLYDsXmnnfIaUAiopnABmxlaOWsnJ0YnX4tUdecsnF7J5ZLyYWRB
4eUWtWnJ+dyI81lw1Zq6lkykHZwQFxEHDhPmBc/zsOqKZErJ/a5bkqhIBAlfvE64bNbYq6gVQG3C
i8DondSMGLMOfMHEVV2tRYyvFF3aLCk4qCVDEqR+aC61OEMTuJwCLFQWkq/3aAwQGHErF5nX+5ZU
jWicVfUea48Vk2do5fcUKB0VyTlx6z3BsWMLXNwuRNtkW/3KRrucyuSE5Jd1FKPXRiR0gh78tUFl
klyMgpP1Qm5Krj85hgkqUr1PTb2q+1f7MRKxA3eeazRNuh/E9/ftY1JZSgl/ljyIL24U/zERG+cH
Jh4XOT4Ew7L68W+1adfc6NaVuMFVX24H/ulDcoUDqdhfd3sg9kaUa9H6SidK6ZNmqKcrhlUa8bNI
XB/hzr0A8TYBkROYgSYcU1mK7M0GKhK96dPdJW1IwjiU6Qen/Rx3kE8qvUlLYZiu3G9yjt1LVqjP
pM+CJvtVZHXp/Guu1Vz2dXo+tLnzY8iyxK4o/6gf0buIrvADXI/mzkPTaCQxIuXbCdykL2DVcW7m
L3Jbv+dDdSZESp26QwT9scNckf+Qfj6Ivbb610BVm5gdxoTIcF3U8EgEzdR/boAM/amiPmYSknS0
xefaspwYSoR78JBPhqGdWpBPT3u9VeRHxcBHtBIjqYePNJt63HxA+1HFmXqQR+9eSjt88D58uLdS
x/iYj1Y89qGP3M+jV4brY7F1/fn/sVlG1CcJliKbExbEUDOSX5GOgYugs7fajIjtbg0CdHzemJgS
0UaLR8B0m4M+bJltrFBUvqWN+WIAkp0JxB8aiWVWcAmC8yQpD+gdmisY8PypzTF3HB+rKlvUFJi7
/gd5joZzRVW3G6kIV3qWdtSzT+9PpuswbNfu8nkALl0OwlIfFdKNNUjfdaxZcq4W6dFq5doE+3Th
VnME/2oHp+hZi6js4eWzjbaHgoj35EKWDO2OZ9RWBF44PhKOpeSS95abWISvHwekMn/Nv3tnireI
heQErEVT/mQfJWaxzj4Qk42g6ojkrP6qnfzO9trRJ28oOQE0LcvaWAW6pY82PrRNnLIFcnkUqFqX
mAmcNIoF0hTdpBGE0v0iYjmQH6u3vXw+ciPy81J6iepmU/twmpB7SBV6G9S/V/NMQ8vZruojeN6a
wk4gmEUjjXM540230Ht+4QmlrOq/UbpzHUaCwMiFUnIm2CN0KhMz5xNTFpvY+ewD2ig/oX8SNtZD
5V/B6/F7+frNp63MRhuQwLcxXxXZijG2522Li0/IYPI/rsMYWC8YeyyHWEdOEHe0h1ux9+tbTEC8
aF/ORcR4KAtwt9oTFDi7Hlrr1MhGJcaUPBy0qCLf0TUyv+LnnL/OhQbt1VnSS1dcF5OvXxfbNlR3
Zh3AQGbJFVDy+UeJk008vfxBbEl0JIYVdyN+c3O1PvGkc2sddErioJEV/HXHGaQipnlPTro/c1GW
PLuhJqEuTqeLM5jqaoeFYiro5vVdu/VwzyxYpLFNUMxaGoenysdHTzdWkHOQ4PP60eJ7toOKgSnj
6tvV+RG4nHmLRF+b+FbFWwlc0pyL+aZRdlC6OUajUTD46UI8Hr27Zfo5nOQc5sZlQLSVpHposwhq
ddLCc8P56xo+zbwIuhA57F9n1zn1OHWT/WYpiR2abdHGhkqqwuf4RwOYqCqd7ykN7YoQSHIkHV1n
z/Qcc5ZocFYp8xowOXyOtdW2so9Ob1y2MsnZDWnZ2ips5p8owCP0sdyxsjgDZwknutGYoPd+oJmA
seFGwJ6alRrFQwABh75mqKfSnaXxEsVxrBzwuJayvMcu0hWox/2BulqMGhc/cFj7gfu6NllXz0Js
sQPb43jCiqzGrmiRonFvOw/g5pKqDjt9DJP13JgUZTbQaXEZR0XiifsbxYFUNq2JP+MOXrFRt0V/
81pawEcoxymrK+77pVfrAkl8QLBEfpEOPuUbSrHa8fJSOA7NK2oWrdoHT6CtA3lJ5/5bgdLDCvCY
5npfRPpaToJ+x5JAewo8266d74pemeSduSa2rGPqV+08nEFiYzn4iQdyuUeK7jq0hPWJNtsHq0LV
P1/PzQYUDQrOTL5zoWzv1HLDC8Bd0G4ff2Cki0aV/MoRQyXwZt2RcUjdWs8Ed1w1gynRMSVxFhdV
31OZ2OKT7Srn/BO8ZMSMNdYLAUBlNvDemXTkP+Uk4yanUQPz1Yw+is8TsCm19UsKM+o4H0P/Q/Wo
XU1/sdzdtPoMIcvoDfW4zaE08KH243s8kJlxA29fKR8ActPBT4Tstg2nY4y6JoVUoY4iTkzvcHp3
p35m56nB2Tz2mMsTnLoLflbatMTm4+mQOLjYN2YljBj1bxSHqIYtMTq7NckdbCf5pdWTjjCPK4Lb
4XwnK/SVTqnugxtix0lymv1bURbjTBLg+MLlNX6uSdJLit5y3t8PHwj1czHkAJiNoXSpo6c0bPV8
PHLCHOoHqWRyy1w3R90c+ltAeI5y+ONbAxrR7eFZp68DEmgG/hHiCxTiTECzRWTIwPJ3Atix/gzf
5O0t1t97TmuthkY04W/VeSQMiufMnJl7L4ocEo+K12tJLMYu3vxlzarBL+N6CXmA0KDB/ijbBBCC
5zrLTHZ3dH/u+WflgN+KRQU2jvQCJd2ghxP3x5m/xv8rbZHbPoXMFwMiV173nXNP3T1wS+0Js2A3
i329610vg4STb+3XfNs6E4rwKgiS90buOxt/UbqyyowLHQUh5P8ket4TX2HXFUOFycSNECEeMA9w
z7q4KjjoGOigf2aSWxjLVcKLwwaZjBAm4D1Ly7Rlp5KQHeZbZ02ta42O0Jn5vcK7llwt571hrROS
/SLOe+Gx8NPRakxZgo3oLvrwYaZcpXw9XEblgl08Gcx2sDo5O9dh6OlQBs1avyEs6wmnl1Bj1hAI
xwgrYtE+iITCDB+FsyrLJ4YEx5FPqPTu6fb2/fEHyIjUwPfr0S73hBPFpe7v//h1fSzmcWcWPW8u
T1q6nKd5sVD5dAAQ4s639+LkX6EpqusSYureAXVIvDqmt9FONDaQnfcxePQ2s0P1ALk5V3yyLQd8
lHskx6FbbT666hSVe9tf0x0ES1Kg2r0zOMW9iqyKtqkq/RyQBGRUuNCfnkvSMYOtEuXOc8stdRYn
v+G5qXNdCMbtWMDrdkUCZFgFIRZl9MqPM0KMAfZePavEXotvxlaE0EL7R+8P6yRlH96dQc1O5zeA
MvH+eQmUmdpCAh7+7MIjfEK00RwugsTaZWAcEgTWywND3ONCheu+Q+/ktSjrnc/D/pPzFNV4XEoH
Nq7fGIGUJNU8iHARqQK6jEXBVp/Ztocn+F4l4RMOSJULZk+TCOGirpUDDBTRHz6shuEh+sXCnOBG
TtqieQSZJT8RkVjGzqq+9mDlMxBdfA4LpcCn/5MQ2KbP9UGHuohCj/Ax0uaC7caPivX5aiJrWg+O
zflmMOdu1hu/bft0AoqphPOPF+bZEHb/lZVPw5urKe1vckAj1Z4ois/7+vwvswuK4OmIlSBnywOe
+r+YFkIV6vPNIJVslM4ILqIAk0m24JLEfAA1z5jzIqJNBl8+W/A9ShmCRUUS9au4qhnTwugaIpIn
OmJ15L3IwCSKNgIn/FCCzh+ru7CCOR2tTFHAaD98cMmvuVQSRyRX5UASCghALlrjs8+XRXXPL/rH
axLI2oHORJpBgjdecELt3oMzp5n2DBqpY0sfGy2pg8ocQV0vcf86y5Ajdak3P61pPObKk/Pz/iPM
DREMYyCR48GdCsRLeazkKrIrCoyQjVaJM8+El34s49hANxPlui1MdwxhoUmzYisidhNpZpK2S2MG
7cMgtqWv5CoCTFUrxc0AF2y5c3IbBqwiVpzwFxceQ4ylKVLDft2otKbAYd/P97/Sj9OBF8Nr7lfh
GXbKZmyKZpnF+7XtzR7nW6YkHSNdIKPWUNKUFWQeK0Dy3Pl2u38afQRa4swiblGge/8XR2SZJGRQ
6ZEK1Qomyn7IHjjkJU4EOEfsKbA6leoEZyqaZiER9zK1UhctmJPKSsCKOSryqdA+VbFZNUC+FRX/
KjuSrorCHVMeg3hGTY4knn9mPxIXon8ww4PWZk9UxoBjrAnJh3KXDoC3ZIIkT5a4lspb6esQUuFD
0Tn206qtw2oV/2H7IgdAT2t7gcNcvr5KHd5AiuoH2hF7GUsU/F5iFY+OSj3zWsJ8A6G3tDFTeLCX
/a3CBZzPvDexf9IAr1wb7pqIbyE/HQ7LtZywfZa4S0klq6/gWlN6BVPgS/fmz2Fpiquh+njBN47T
E9uthJTgpGUUDAhsZ4oBSgYJgGjrHFGZ/NyxNd63GUeZ09ujIyBMO+45AWmxzG1yicGLfv8bYjXE
wH3k0/w+8/04DBe5VH/5iAYP0Bet/PJ7Z7s2uQKxXahbdO8F+gfGaBrDz0ZbCRwoxDqXKmaxia5t
FlF048rAx73uPXvQktJIapoESYdu/5b07BmoyXdrACbXFKIN7ePj3hJNI4FRKINHpKy9H0WG9UFR
KLHfarewWLvb5pOYyxGn500auhvaVKqtNAEpuatC7mykkFiEIJQtbNbh6pb6FDPWcYR1u8Qe9ljN
ZtvmI2kEES+RcUI9jTy2m5WC9A8aD6yAUJN1YNgXQ6ip9xz3flMVZxP/zePFOCDn+HYXPI9cm5ld
6z1Udklw7nT7GjXBFqYjJPupf7/7wmFnE/jJgfdY6zuuj/aMhZMT4HIvDLjVt7PPwSdnU2x8Bm5B
+XMa0hw1ZkVMpOHAkAdnSKCtvFDxFBwtP1iULYfLGMZ++esHG4aIy5jFLWcqjTfkdis8ZtwYnYK4
NeBPyr8EEmJqmfLOMQgndap0KdiwtchZCy2mk3vl/30JczU6CfMgLp5pEEyzKw1FiXjYxhk1Vbjj
6+zpRD1hSRVHIhvH/OigDhHq89AFdJQvMH5FedK8ZvigijGmFGjBjqGwYxRw5SDiA1hYmdNMW783
ITxdv0ONp0DoNxjD3A3Fx3qB5eQMp5+qpgQe1y4TrvP0MlMcTdBixGI0Y1ab0NojWERCeNLOAabM
/5ZJC0nml0rvcgVG2qhhZ4BNIpBbJZ8hR/cUmQ1TeTLy96ggAXRHGH6YaI6/i9gAV4P+MzfVkyDd
ofeahz/QGJyTIpIeqA4u1+wZJCGoDKHrkzcLOVsO3f+EbgG2NUdVLBpInR3qfEQbuVviD943luTh
07nxaVnFBbch3ZN3pPlTk+3NsuZ0ntDYp6WkutPkdDw0ESMiuw7TZA/+f9dd77H7FHLyPHD/lS7n
T78mCpZ8BnFjx2Qg6cbsMmZHcRndt1xg+0GKSWguNuGFcueaPfs0GpipXyOUiClt0cs3r0+jP15A
KottRnG8jpMeGtguLrIzQxn2IJTn8XicdS1YbP8jXZuy3/BzQxJBQffhu/ACs6CMDob+vrLRTTWZ
IHzHGFE4/ewuU8tPjKLNQHxsFfKlLVWLD8yVv8bW5Xt9x63tlwNVkeBd/GUHVWwjLs7AoRLbgjeU
cZNJVw7hLGivtqFS60UfrX5Sdmt2/kXZAF66ydya1jlQRIy646REjJuzd8VPx5GeXTWjX/5k0gqL
qllIByZ9zaoRdbhdGaFN7vFySLPgkRvyFjNqPp5jvJTgR5IcWYVFjypyf+6Nd5Pp2aJG6LjAvfRJ
QPRdjkj9z2P7F5L7UQIdJOcwUDXJz3xhy+ec1FU0FxR3ipps39fyWGmU7vp+bIyAf7gtQylJqSRm
zTcySgYjDJMw3AM+axMhWKnrd7EAxaVrCzRP1lOLzkv0Td3+9uuoDCQButTHPD2jfRh7w/3nL5X0
0CqgJfZdJ6RyhwFFup+zqR82nmnmVbglixSWISvjKGbs2prdppJq2QMtS1mEwdtQQQMhy6ssvwwx
W0qbGa57lSRygoWA87D4QrDnEOMa/s15gGdEeJqLoeVEwzSSpJmYp4WHvUWYMcMLg7T7agnMhcS1
JWHWzfgC44eszk17vtijH3uHUgCuXcgrvA86B8W7uOfs2LGESJeHwVHmy4WenhnjUCIpU93Qd7k8
YLRTxwuO0/ciggOELNpDPw5Bq1/lE5JCtVCiFR+prc8XhvNssh+89iv4RTi2VjQuDxmWmzbvlGaz
ix1r6Y/FcafplhMDKmE88c1Q2Yz5XdUe/CR6cNhl0KSwIOe0WWNpB9F71+ntgtyUFUHYh6rm7ZUq
tpLEmvXuRhx9ipau/yGQS5sl4ONT4cDiwHFOpN+ETskuzh1SxEE5PcIidBkwFNh7/QQrQhH+6dY1
djJWXwK96mBxQwvLNxWI1SGgc7XYQHXx+Jy1lPvYuNVwW0s7a4FHztaZkG2hfMmmqF7ReNXE7mAO
TwWHVQmjOSdAkAy00iSBhGp5vhF3rL2F2F8phHjU5O8WHPgUSVibu6aPLBH0JukW+qlh/tGZ44FW
KeQtv+pTXS1WdU0YcPt1L4TfImzVyL0afMy0zYJ1yBJwK6AXxR2L6l/FkYy93hwMr4nAVAvbZDDa
LP9pcufMqC5Gqs95hdgiB3Lu/4P7YVz74799gfFCQUPVNR+WOie8X6wetPhq9KtNX/f5zxeKyu4q
dTePefvo9o5OJNLOw9dS/B1IwyiOU+d13POUxufQBg0HNp3AkEy9VeGcDrIBdrMpYGfLmrB2E5Xy
Qkwq2gUuzR3BhGJ8lCCem4HdRwob0UAMbNZxk4eKfMfarJHEkf4K33yoMdrM6ruqXGZc4/g8cwsR
2orYSk2V1ALsLGdNmyA+aN2PAidV48HrVUMVUq3fpkAZxnLLiVgeb5SDFT2vUl9uthygpMOJ9yGt
u0I00EwAY3TNpQtxDC2mYHkEeEhTynC4kw8yq0vF1Fu+9MceOkkLgd/QTtgBdNGOluz6IkqgjsJM
AnTvSSWemc2mxEfrngN4LN/KgK/Oug+2lD1xmszZicRy1tdsjA+S1bV7tR2CvUTT+mBD4ZhZU5Pv
adN2cg7P7Mpc0X+YM9xxuVx9AgKxJ6Bn6FsZcLS3CP5JpN5/NblLA7ANEwI9hCDWqB6hIBDeFIc5
5rPjx0kfLWKlygVxDLRd/0R0jURB6bguSGKaRqJehTBN5AUAhHbUd/SdEqOcLRV67PY+n5/mPQBM
NWTDkjcKB6BNUMgwkzmcv70QFYFCDjQTKPyKZm9XhcxfPIoREiaHucjJfuE4gIqacAnQAzA72JCe
Ri+YCxsmtcZfgkGd7xBMqwS48G6GsP650nYLRtL2w9eTesnCkp7v3XY8qX7suUXzPXCnbFQSnFrO
SstwS0hdXofeHL1KrHgBt17NyVlbwua061RacYnCYcvRlrpNzfMfednCFNrgLLhoHFpb0vgDFbct
YyCLMjwbzHyK3Ac9SsYC5bX57h0AY2qdsahPiVMUzBk44gzz4OlD9+GNqjF6cPlghfPQSOJHd/u/
OJzFw484+VZwNeEljreJ756HCYcAfoQNW9nvUTtgB1EWxQibI0Y6U+i3xz1dpcQxoLVMzV23jBxq
4i4xcNeI4EalFtaRTslf3T+p9VSlR7R9syLjcoG5/mKW5i4eIE38boz3dajs7ledjZqtffs1etXX
Z1vK74YcTzpAZcAbZqYXXEoy3axJkJlCq5n8M1cy7JjC05AF885frgcxQRh8CxVK/OP0uzB1BuZB
HxtYbYyg5LSGbw/iIhJyI+a0AFQ557uD9dyDM3NRwwLGY6YhgvLWLQBSFwniLj/MOXHW5xNbTDnE
bSOataoJinBEcdISAIISDXVejQQBFrBF+6jNKqTl9TVQuEerm8U+aTGSulaoSwF8NAbLVjaeknwA
llJYmEdi3Q2xAK94NIVNN8y1+6SLMWau9FVGPdAlznrcc677qVVmCwW+4WM/1M0bVKisDM1qUh0E
/1ZKpcmOUkvEV13JX3vNzUBWf/DJORQGaIvWGPWd/hzHSTKBwr/mrR85FgVls44sTrkEVKfRdUdf
TUHrouXjQS/cVAC9xmGddHRxYNYb6NrTf9XY3yvrPMod3bXlzsNYLcrxy4UF8cxrazcG8/PPn1PN
c2txGIQxqx9X9qg/Oh6fxWXPQcCCbxPW/VVpkWfQSMZRvqZ4b/JBoMgOXoMsUGItnjnnmNaghTMj
8JIqqVCLXJeRiCFNONVK0O1qi7mSA5CIqTYqyZUc3DjlDqguiRhgFeYGnFforQkWHFYDf0rb+NOY
M0W2Ct/tF+xGltkqjOofgl4/ENNEbVelUmEsRK5GyqndNRmkiBsV4WJh2mxdvAGGvcuZ+NUUt71C
IVMRtXrU55iaKjdusBNRqck1YIm1uZ+XLqajpIRhSOpOVvp96Hgr7U13HK5NffyZUJZekcJTnWph
oy+Nj7/ZR0Ml7pxRwZPupa+YA/wDtMmRRCSwcXZ2yxgPTfeeZv8AhxNbn3JP5GR62ilSgoujSRdR
0Vq62R23/oiT39d5PYekaQPOE3oZBO9vMuh5kgxKvwb9r539VUv4RFsj9arIGZO+SD3CCsSUmL8q
6dNw9RQTWL+Ao7dK5xkYFIdSpWGBsM/ifSt36B1XQ5E52BVH3NcexGo6v02asKWN0pgFA5hJKo7T
agJRqJ/Logbv8PPU3NA8Lvv8H0+cesNoNRrcFk5NtfXO6Cd00ypuIlkNB5AlmaXJazwOla8FIXNm
Y0T4CgadMnA1IBUaaNwq8Gss/2kAISoUMTc9gKxrCXJRN67LQtJHtGM1YkEvr79TGy/QN7kOAqq4
kn90FwJhxOR5lWK435098WXJ+6mDanDrLIXoq4MPoXy5gx2uxUrGaW1rLvrta5OsXpOiyS+P2JLw
XxPCIMywLH/UGltz5Fj1qxcVLf/KkZmLjD2HM+neJwidiaRjbQKwSMTL8+anbrOSgxKsKNv+Onh+
IzzqHOLuCFIXp7vego+XivWLd7k/J66WQzgpJKhfM7VYsdJzr4x7Oe/rtoQJWgRc2yDNO45fdFMp
bNDuhBeOkl0LYJw0Id3RqIcMoVCF+yHRQV3yRYLw+OSwjZHSVujzwZgXDRvW2UUqHBbGAwZD9fB4
7RTq0X36EO7uQirM1My7iszGiW3ZZ5Qu3Jg4CSNCMHhQKs0dtE0sMm1wf85wfqZMpotQnnt1qpgx
ZFz9rBzscvtbIV151+EyTL+9INCIJpR7EQTkGWal0fzveMlAS+n/cDBtw1nqH10JRWrKKf+j8dgm
+f+zW1460rXxK0YouxoUNjv4E4cU3/JWEEW+1hveiE564WEB19rjJdsIISplBkHTbjcuFsAEYtXu
JQ4fw2bre2au1yrZr75XsJGqVsiTm5R5MrBaQG6VgdXkHFt9qmvdNQvkkKE25q1iUY992i3I6XLs
MQ9vHGvubrRSH2ArQLdhMd8XQnNuAaI4KHdJ+u7GUl14Wcg6RgEJdxdGeWG9mumSVCWK79hhCZJN
dOXGqG/z7RfWYgHxYxper/F6jn97Ca304MRByowaJMowBAU1OVVnynRsNK23CuVgOh0ieKpsAv4Q
7F4D5VTEDPjdnyble8MSHTJZP/2uWai244tdPCsj2WcQ1yb31WlcFK/G8vNTyKy7oUPTe/+dFjzR
XHAs/7vR1KaL4nhIn4vnr3EgWiUm0CyNWN7bkdrxKTn0mRT8bDshX4/rG6DUd3l+6h8QhDgmkaxu
9tXVz8M/S+Kj2EY48DHBsCHVFNDTHzvq+It8Cc/WfQfKRifCsLLsDSnxdWnBAhEGgV5MmMVLaFL7
f9c1fSMV4Iz13bV0jLxfk1P23j988+l01+pyQNsuxwdM1DtLkpCl3Rs0VW+Xid/pB2/1VDU/JkjF
NnLHYB/rZbpGkeIjNt2+Qi2UMoy8qiVRpElSBuSypMVdp+rNO+tznE+PTrA3UMLWPLZqgZ9QPfoR
4m3ZB5Qx6hshuoUesH5BLRgS7pOXbawg8Sd4t8bDYtGhWeX4LTMgCTk9dDeyBbwBNHucETOLoKKx
xnFz+aUjoHY+yHX+38FIHOaiNhBgP6YT8g0bhnkG3vDFud5XpPUTHzSbCltpoUnrmbWirqqXEoM7
kJKlxGU7c+nlCzEHg2aALQFYXrMlsSQXGs3c8YuIiG+bx3PMPbMP3eXH+VReTWtFCtI7JKUx41S6
C0RS9FbirI4P737WSzNp3RmWFu9OlY0hfjmyXVYomOGn2yEC4RHip5AgvzCbu3NkrV8BBylvVtBV
jtx+5rTyFiAoLXdfofrM+9nRuTNNPMJsJ8CMFh2PG7+vUUCsAdekPpQY4p/I9OfTSletD/zEUMZJ
SFBdhqR3hyQ3r3z1WD/NZ39fIt+Vljj0YXNveDYoKQAa/IuNSe0EIpqGbGSZT770swXBsQzxTksf
Otml56/Jl7KXwP8ww0bC/8LWLXjSM6Tt181bpc64ADqjSfJU9hDGc1ARyCUfq9FT7oQRkz0cVePa
W1KE/Tk7jK16YhEoXb0u+v1K72dnQTz0kcuB9hNQOjoTG58u4nli7qzlA+BRnEQLProbFAFoK+9r
BrBX7Kevd81IensZUIKrTLNQBJvltFvvU61vy8OvDW2BU1hH2yOSWeXo1AhX/SgnEmhFMXw13wh3
K2d0FDWsD8pypWz5be2aZorxnxTqPH1VnXLjCV7QIJTdNp20IHdxzb9KmgwYah5sXczlnH6Bwkmu
n+8pkQ2UGDvUjOrfjB64hlbFB1Az2coMPH8pbZHds+MXQquEo/h0N4WaeCPGFFOUYc6BZZF8g0fb
1Vqa/ANZfdbDrRIH9sRW/D9cwVRjSd4W9EkI7cnwOlM+Jim03BvZB5sZlaWmje1UUYYxImQL0cyg
SY6q2AzRED4/AHfaDH+wHq8U7RyhGFZRMBZulCqvqzMCdAiBuyaz+/8X+3WZu6eCYeZrqCeqfqyk
5yahchaAmkPFy8t15tSQ4iz68zwPdn858eA2a0nPc8p16PMn1ktvpHE56RCpmJsl7jtgnkQ60HBd
QJVYNm5cWWcrxcEtXAKVJLBfrF+RcSmUgR0wO5kzludDMy49pO7/qPGYeK2pTGLXPslsJOJnBwFW
EKT8s8zBUBTdoLK3PHAPyIYqCUs4RgfFoBaLJ9n9OSJrtw0eIyGuMPxqZKHwZZHGK7Iav6RumIma
RaUGWaGTNOn2aJvOuVUP96CDdKzrs2SyOt5LQTU3IZfjSJRwo0URfiZQL1BqVMivKvEs6U6mlDfe
zGHpnLWq5co6PF9WGXNhG86iMS4ml8jxMEgYCbWeHNGdOOynfNiioiRunSnyQXcOzzeWWLZcHch3
TP7WSvrlTpOSmS+R77nZNsDyG7JfHVvvQkNCZLLVsk/zuNILb7+LogG99lMG/4PsbOaYdtmD7Ess
w00fEcQSn/04OCEDYTQR2JuXwW1hdSG7LrBODBSPRIoTIna99+veC0zmtlnRZPGG52rEQkayvonL
6xmKR0ixfdy3/Yp3GXLOmzHx1hE6OGBrs7VopgEfiAi60FOHLi5Lih5o6iVSSBnDNLZSzX5q4fut
eqwLyLRo2AJDVNxH9ki1H5+b74VYyNlLBbtR2My6BHJ+hIYtMpKEC+UMUwy9IBvAoVBIFLFrbyV/
lsfF13cVIImsy4xZ1AigoBk7nMemh7Zpu+cdMLxjz65vqq4ewZy38WDCFRhJDsNQ7dHAC2K0hSND
tzAHb9Xg7L8lL8jmyOVmFfiD8rMkaerctu3cGVkesUUr1l+SBYDkX2MvmInRzEUn6Ml6BTCIjplu
LZdVhubix30100jVHSMvkWSEBAHVd1xaVd/Ue5Ii1IwNKk8+4EtsWyFmWKnwbU7t3VTkPc6/wlWo
D0JorUgpYm+6rZ489PXd67rwKh8kTEIy0tb2T2/aITkfA60/k4ekyfk8v2Xr14cpNAaKmrMb51TM
xcYSu4ZVVVrpI/RMXdMAqlXQbRnMGYpnL4Yvy2SneAnxA3LR488tYI1GCjBH5SKDV+Mord+N8lyx
OiluD0EAfRYcIKVTEULSeTJsjN+HDXxjGkBBMZoek+daA6if0yHbElwBTGl+K/jrIFYk0UBtHRZJ
ua+Yt0XCEKWiEgeSIUKlDBNvWIVLA0fPIj1UH1jgBOwgQz9ZUol4AHMRyD9u14Hef9ig7LoJGe8H
V6PFJhPK/MnC7znvCcvgif6c0UJNnNvR4HSvCX06D4FdM4xQ67peYQS5SuLHiEYtT4FiEgSBIT4R
kUFDgJR9ADU5wHqO2IoNpcVJO5oHRKxjkXc4p25x4oz5QNtipJ26md1Ugdvf0D44prrt5RXw/ZLo
6ziMPMydS4rEUuWF+FJyNUGR9f1ZCpHAifAxj2jeYu4q3zpf82lSkMcM646bFLptsKN8f1B8SLEA
EjSsYRUSfbE+5vjJw7/c+2JOWC648StYBr6kNYH9FnWtS867ct1W4rqFr2kcFXGDAVwljVUtvXlf
NoHs3/iUkaUcuVqMGsexRfOj1dd2JhwtTU/mc/ZSTmiOXVYNKs6F4DheI5IYw5TB2CuwC5rUIr40
M6ol8pDHWAcS4BroJBCa6nFXbNO18yiR8Mb/9LE3gNEJtl3V8dT15mkDXJIXNm1sfZijHKg9wJB8
loryp+JX8px9BsXsn1mVYxZvFbrNrXyXiI9Gq/wXKlVNqN18y+wLsNcmwXsf27wWjJYkugcA/9C+
VldfLwYrJ+5de2Y+YUlRhp3aRu6ACUMQhf5vuYO1urA4eDTdn+Lu2NcUViHR9pnZ35dyf/HUj63V
GKxRlC8AfKGENGrEP5PHRKXN7TvzTLrOQeaOF2jWQcfJf6rpj7t9MDn4SrymjJFmmzdM5unzPlfb
FBRwuNuacFJN2E1h5Wkwwyk6Dq/oGErvqqLZW/mzHufR283EGBsuCAhJHbuRzS8TjLBJ7SKE57Fm
3ryDNv52d70IJMNZPH1W/ooB3+PwibBSZPYlnr5u7wq7GvQw2O6mEH0Gg7JvP/JkZzJ9d1DXYGaO
owL5b1OnMWZKrdg5OI548N91k/Q1MeAJ4xmCkeDgrYXl/sSw/QGKDpJRHndyvFtM2xsuXwsmqRmv
fywIYoLXK8gVC5dZQ4Y41uw7WP4zm93gfW+QnioN5tiwYgp79pjOPBbdp1xEWVCQIuBtbnBY/Bab
zijrLKoLkk9WN/M+Hqf61LWW3Rg0hWI1TUcxoA/CcdQX00OikOk1or3Xg0EHZvnTuiF2rzijKGqL
qLYIX99zOukZSRgIjn1wQvx5xD+KJu6n4m8A6z14lsXyeCUKDkg2BwwCzueWjXVaRwfR1dIWRqVd
xxFGQ0KkKLiVc2XOW2WzmRLnDXr6v6WFkxoDw4CevIs6/a+q2jlIFxUpMTq6PVR1PhxoGWucAII+
9gqAjNeV5NOXeaTztjJ1sUv6mfwr4eq3CUjk6THV9E5sSEw5lA4h10OfLQljj48BYcxAVS5MtBg8
eZpC3I2yO+YL0K/Wej6BiaCQXcc7JiNKdNhV2bmBve2I9TjJZY7BWGLuhXRaKNkeAB+LlcZAKSnG
UvMINphlXOzYDmpeIPPgE2+GsQglq4LgM/Q7cBZHUfZsmelUHYeNgR1brnPC6xgNQ5y9gS8n09nV
q4Wb4JtuaLVI6iwq5TFavJdh4uU7qlTol9ChDvQYR78f6xebZ7sM4i9LGja7U+wnwjZd9tMjwrjz
qCdOI/lxkbtvGTxJEaomS+tV3iMYcxq7FuVWluo7OB0q+15FQBcCt8uL4c+NHy0VWdyXamD1BSE2
n43dAIoLeS9Y3R2nTpZhkNDyqlZu4r5AkMmsUyIarXDU+3noSJYKcyL76MLOYFhidolEMQtVJZf/
6hcvCT0jEBxMGA8DOdNJ3eTdYeI3ajuiWgEp2IoGQdY1VVqjqCA9xSDyMa8JRN0QjgtpPciv/Dke
Bm6UlHM+yArEaMYtPFJwM1TB/OVav7x0mx/Iuhxm6GedJhv9p9ZL0hJ9LJFwgTqsiRhuCfQFtJaE
GRQJzw99vErYYMEv4YNorwNaxZJ7THNqpUsqcm8VJlNBNjKg/Vm/m7TWnn8CrtLU/xMaA1FJ4SjC
ODCRIlj0+zkibRe6qTiPkR3MdLca8K2YsEHFQUFtx/waY4DMQSM0q0Zn9lAIc2U1XOAgkEDDd3Wh
/rEatl2wNgA/DPGfGXRZTqSrz2lCu/rUEa/8mWsdSkhtCJVtWyDBT1QJ7zLF//0DhgYB2bjAORqs
PaB/exj4q4kHhoYGwjElWwW18UVVHprI68tkV2EiF8rjS9PzmjVkJkuDL6wH3uPr8JDkuYC9qxt0
wU4nLSS6xfJgG/iKGG4EA99/CmMk88yK+KMRn1TgCIz+xXu2lNQRBpqfMcX7AbmcT/6oBmAuZ4Xf
wRfGtLLrUelsLvPF+aBGIvuwVIGimcKfGwubPLn98I6hCsc/dubd2YDvrmoVHQvESkliLh6QPfbc
Xt+blRGyALlwdnY21A6Ty+ixPs/QABFPTs9lT9+IFTJ1TcG/pxc9Jwf2CeDUbmcTxVgQTYYWcr8j
VIRuqe+hj8sBRam+JJwi5fGgZ7+R8t+zhMRpCop9cFHKu+YJYTtBd/7Ne25lzUlst6sNJWxkyJxI
KKnYPEYpMGqVuc8ZpKc+ebtT/ALPJP4KqMuvRneu6YWTg6QIBFaUi3KQNSIJkZwgWrKbb1J3Ks/g
pOeI78FEh11m1bhMc5u1aKlQSzRG7WLB0c1YeSGwpuo+Sru+aqL6lvYfWl+zS7AGYHxVXvo8ZEET
ZTkCx8QJqwLqmVrovJ1CjigZUIvX/w+ZmHQHOj9QLS2ltEaSYQFkZkvHW23erqp3kRZvHICkLwGZ
MKZ3TzxDcfrY8sOmiY7U9iksWNzGHtPB4K24rRECtkqDuXIL4ktP5FgvxRanSA2UPVGe4VtyFEzf
AULIw+Bj9GY2Nuh9VOSlxWldZEDHblUd1cj03u5UjiTfoaR5QTwgdTIlptyJFV6c9z/1/d4G6lpN
z3/C6fxnAhZ6SgrVa1ncbSOZWbz5t+pF61ScoW1Ywx8J7b+JmvXutga0VK5moYXEoPQAkcaSWM9n
NJ3wT/rz8bN32ftH1htKcY7MUco5zWcDTldhy67fpC69Q7FOrLYiEHNPiqn1goa2F2VJcW+5JiXz
YLqY7RareI/gcMWdVsNaM6QF+FaSZeMe/EpZXTTjWHvROnE8azRfd8bmqxxn7y1CYHw47Hb4M564
wqI0Ljjf5c6K5jRENkFmOjYeCd41DHLoV/y3ayj/0XGzRxGmfN5OLtUp2nKVcjYJ2Jj5UaO8eN1B
HqpoRdq+8rRW1bSJh3AGvVR+0rnjxyIs0T3bCjoGXNuCTGye0IfTAufez5LEP4Zg6RIsrdtGDZ37
e6lulPTEfvWZPmLptntVDpltEql87/vNGI/QKgdax3NPe1f6XPU9qAbnSupsFVTHh5nkcRCm0lfB
cUZ4G6uSxUlEO+TpkCL/XbrP6bBqPKrxTe9gFWBXl5/OziqALYO+zWsqSqMu3IBmkjVEQxtFFjH4
URXkQAniNKNR+3pjatcY8oxOJh5I0xYxr0Mod90wrIjF9618YXqKv33a3OPCVpBiHzktrkFDwe7x
K8Cepw/LyOkDM4DrE9uveiQIXmXC/d0NzJYTigfDeENokiZNwD8qL6itaEnayG0c5IPhz/eKorBf
fqWgI/iFH4dEs3qUF2l8qzxX6LgcaJHmSJpFZZMGi1OO1xJ4+ldzNL2hey7iTMcPpu8dStnWNwkb
irzgzZTyTiuHoAsTB277YnQJykmQtth+ufKWxSntdnTawo7rg0n1BkCEkgmvhqVl82rBzTRmImN7
qU63Kpcw5MToozdYKdeqLZizSWR2yMQJHdDqgkMweWUMf86tlkrIJHIM/c8HZhXFG/tkWzwQg+RI
JG3Ar0amn+NpggyvexAZpSRXXZRNEkLhbpIRU8t+0B1E+7TtOytgy/Uhd+IdyLfsIa0rTb2cXIHn
eiWv7xgmEENTmHY1XvVL4407IbJWTMoSKJY9kbVvECX9HpSk4FGHF3oqvVsN4EgRnwOyNu/OBv7U
i4Za60ZrM+Cxcuga4D0a3qRz1dTYSS4xbvvgKYBChDL9RywzO3yv9SAUehvIMpi3v8RlS+W+sb7n
wFrkAzkSI16sRGMsRGW2QOrwQlKNLuAiLYmLygq44yk+v9R+fzSYMFhoSzwbOVDMglIwYR+p34j2
yBBA++4NmPTGKqf+CeUwJsSFx+Zco0w1IqxjCv1YyiyXRIASz58DfP6U69PtZzwbdBA0sdT/vtQz
VeaFwQ9+WawoXlKppNtZQXprccLSdYngjfYICy48GA1kXm7i2wa+E97zqsLJoCOOHyhDzSSnL9rb
zIXPUItjjfG8/HCftFQAnVtfa6OQukPk0Lana6DkHdEeV2tmt5RfY5pkMCaKmI1VPnFdJFWytxvC
6yqy5Dh6CGTDUpt/gB1HVjqBG88/N5FzBnbkjq3phFfF4VtzQSsnRnFW0i3iZxzfqK1V32PGUpyu
NRMkB8rP35bS418/LvtMmuuI9YqjnAchXLk0Vg+N4hRdYFPkpD/C4Ftrcvtq0AbXMefiBJbzZIen
MLk1tSttawzL05oJnWaznt5FkQANHQMK7MjQpyIiFKRs4da2DncB2zgm75dYQG1wQ5R9w0pgdAxY
5Pn5xayQPMSZgYDLXHNBkNN2YPhv95W+o/QelCD7RhPOsERpcsZVY6MiO7cThk7BHvtB3pg/c3xw
zQ1RDcKzxYvvqSmWHL+OxDg2uvaIOOaaMU/1p6Fq+pidz8dpW7dvmLodetYxRsopl3yzhryqJr2w
bcFdYhwjyXfQz+hvMYy0/ccdXT87m6a5xeMxzWj5sWOahWuRGoZn/Z+FBbXTDqf/V1gLpjesHYZL
yI6BojHup62Pey12zXkHdegc29a7gysL0qYQPDw1BUdtDqP9ysKQHaUsDOhZWX5q3RFAOxeU20Pt
Xro0sL7r5J3SH+D1Hhq0YYeqUFS6eUSuOdW7s3ahvoUAi9S2u/e4XDWHiYndc/IvX0MqgLoU4Yjs
M1VeujaUFO+4RNrhF+I+tUn+cAww+h5uHiEJUndWLtP8BChaD/Z0v70jeNwPxG/VSgOUBMx0DwmW
rm4aec6m4WkSw02hTcEcUBOHWhKGTGkRYJNaKNrU96zlh6E9IQyMSV2xoNlxdfM8tWDf+5Fq+cua
z81ECuRPrROYEbrt4IaewjUb5uC9oEt4KwnELbJmvCM2JffGvTndcuqpm9VLuHkHcyU91jgvhKr/
9RdYMEoeI/oEnSthPc6jtQGTK+JmjpHgtGP7RrYzoBk47jYPaRucYqKZu+1s3OnWwYGp+zUJOjPh
x9+9TG21ZzLN16mGWUHX5v858M6M47cYMdUcn8gZxQjaPRMVTP5VS+fhi+erZc9Wrrk2ApvGkGQ9
RmPJmztJViR7NnxaaROkZWcImuCk9o/qVkDnaI8CZ95nJOe39GNNXvXRyP+YryZCqUR+kRCKZ6ge
/m6sXDTRQTrttNQzbsh/cDUALDwnQNyDd8Mg7vifykST6wsX+jkybGV0WuI48XopnNvTULMoAUEr
RBywwhLK/upwo9MFURE7J37hDW7nWIp16IS19QMq7q7BXsGnHSFCF+FduUnApgxLjpGvCilWu9Zh
FQoFjpmkhFIN1GPX2PsUjVNe9xuCR3DV+1x7As7nQmS1R2Y+v9QF4d6nHkMFh92yLZ5mw7VobKFz
94UKM+zyi9/t69/evFe9P96hQFl/BRyIez507s2PerDOLV2HwmZDnV21UV5Gc3IeciHQ2y5VXQ7e
PlesJUx/HTQOI+BXLDJ7m87Yp8CRWA82W/Zj8TzUbx+46h4hVKLWSeaiSzM+wCm7+fAf/0dTfDk5
RSsNL8qH1B16+4VSEx7cQ7HwftpXw4mhtQhj+A0nIloB+Rn+HTzGg9NFp21q18iOShCjkEFtWhzB
IKsLGbOBLtrpu3cN0Q8cU3aKhS2RllIfT0oyiYK58Yy4vV3wAW8vQzPNj7w8rHNtitcLFHzEsFbt
2flfgZhDbwxBpLA3SzTySK2Id9gv71X7YPsmtmXpJgqF7STeIAFPNRSGnrigRVfNLG+bXHNbZXmO
QnfSOqbosj6FgQVQQycy1imQmXw+AyZd2ScDjMTflm8H6D4fi6xSR295EMplGJc7/G0gNy8Q+Cvv
WFv3/JBrRQqqjRYCzso0cqjPpkgsHIiZ44+ez26K2GF6ZUCnf574hBgEwRERp1sZgbkhxuqjJUvB
eVM4/MoIygQv6i53g0awHxAMf0+IdXvFYsT+VI1Bs9EjA0Rp4OrB+kuuhc3AgLqOldPat3jH0+to
VkGSuy34KpN1EVSM9fFthZccdszCBbX8cG8W+xLnFJCfSLHuC87cTCPiZTB/zFRG//yZwFm3SD4E
KOhJEbbn7jyWd3QMaXYVXV8QVO6ak9oaRhG/8/rna/U5jtag+x67e3cNAzw0U4K5tl0p8XOBOPTg
nzpg/uS9kRzX+uhZoEUVCEe3yv16eJvsek2OX6Jfyq9t1eUXjATHZHS4kfiqYAp0m1OdwyEEG5VK
RLPoMROYP2uZ9NtZO2fx4klwsnp8oFsJ49YsZ5BOnQ68AqRlkt7Ajl9v2ksnv2m6oYA3kzC7ftZx
eXG3lslvp9OkiSoaSbPKr2W3d5eEIZzM1PTDyRUFf5O8f1dVN/VJ2/7fz59coN8h2R4mGZE0GkjQ
QUax3mBTC5XX+BQJ2UkIp5Wv6Nl5D96AjXCoL6tss5kf0O6YE36LKwLUuViNtsNlm89QGH/+D8Qd
UwGwVZrv+oYhuSk3klEiX/9LMvZcyVG4zpSIUQ2nU1j2i+t3ykp+978K/IxpmoW+C9lCv2yvFNlk
Qoe5ZNYpFLJ1OuXN4Cwaz5HpTzNjuIGwhEPh5gDJkvJuL8798cW2HwlWOThxwXKwYmBNILnmV3tI
XxHqILq8/ML9Hwx1ARyrZkug5TSFWRf4SV0x4RK+5tL9ZCjQekqMZPXqwyoYyKmKEO7Yt/lO2kOz
C6A8/HFjo3BtWrO/bhAW+KLiNuYSyEmQcsBAxB1uNUAnJz/H/kg6K2tENMlo6JhUM4LBGwqjq9VP
gTekHUN0ONY86pIdEY9B/YTJJSyYCuCq/HkPBAXnXkSZvAqhvA2ZpBP9OUH3ezyRHI68sDuIYW7D
QW7TVDu5GZXFEw5tk5uQwl14X4pbGdXaOdap45m/oqys/z0OexVCbbct54cQxVenHB8MzudrsOQH
PY8DRyc1DIU+yFeceoGpak07AfCdrc5hQcZwcAhrax+vdO95Gb4QpHmip28tML/7rzQFrjITpZNC
wYc8BxpjSAII0treaKuxTquRmYvK4ZEh0U9CWtFJWig0z1iHB8A1m6L5fcuf2UoTWQMkZmDVrE1c
rEYLv3JSQuJgBGbrBpI3hXSuOonieXdcOHQDJZE0D1u1orTlM+Di2yuQ2z7dgrN8ISxke/o48xtB
zIHSQWhbc5ADhSHRe/TwC45m6ZMk7yv255e/RuI20w9GDwn6dDigQIyyJqEhMySfiH810D/L8Iad
TW4NGsGThFTJKZ8HBCknfAbTg25nJLciRbnvGfbKgcVnneEAoiHWWBboy+PcvlFN1jlye5DqM4HR
4/iKbbyurR1tkrWgWlyZgeuOFcBI/9qKz/2ErQPt9g14DfMK0ZZ6s5B5VS4WLyrODTBXezB0dcNi
kd3zagPZ6EnkJCaJjQW//ihxSqQ+IVjDsSRKkO75mtGxwh5KJZIzAYB6Zkk03KqAUOHZxlGHaDJl
7AjfAQTCLUgUWCR6tjkjokOYbrU66AT3RUW4mQyAAieZM/GC7PmGkxrgMj0GWXypVN8OH3EkKGZl
xRDSYF7BNQOPua7xMFVJ9hAU8+jPAGJ8Ay2gsD/IYQCsi+xy9ilXmaOheA/FBv2WMWYIPmN8S5Bd
XNkYjCjONDwswfHekkZ/ATVqSxZE8cgl3Z4iqtAmp0T6CKUnEKGpLWBJsk5kV7369VO1N8oMgf7l
DRTuQlC4C08lqdkO4AUfdQQZcXKDvUARdehBsd1uhVoULElQu4Z083CiFTuhpJYLaqqrk6Ye2q72
U9LHyOjQc4V2934xVcYid0SQLUi19GVxmOyq3Ym1MRt1sdl56yg9C9NDj2pNGDeZOCSLd7DjCd6J
ErMWRogImAPPLBgM6e/59t0GsTYkQrvvU6hTM97BjMVhdPukszAd4+e9EV+60MVCdfGqaKHpWPmD
0fevKg1EjJi8v/hMaKun+G+ZQDQdYQz3JOHPIj6dLSd1uqr02VDfe3L9JzUanW54Rs9jvJBpEwbw
op3Uj+QsS4KiKlKqpTPLoj0VZ6rkwP3cD1zaMsWFvI5y6S+k5JYAHhuETxzOsKG6p/rHhyb/IFAh
7VoALxcnobDxMJcU3QGZDmvX62Ybt/D5X38wyMlgY/75MnxX6+V4Ht1AsIasvJYXEzemVYI0vfcv
gklKyJMZQFfRJ+OL2DX8STDdTU5Cse6teVkb8ue4cIOxOOSlMN+L48Xn8590SLyu3KTkUe3Oel8T
YXdRgnGX0t15/bcimoUpX3QoRtEJWsg+n7m2Vstz3sfcq/jx+aGfq7Hm3LYmb/WNGa1vEw22A0JD
Doky079uQDJd++Y+T3ZNqY/RiD5phAzT6Q8b/ScapPyIzPiBNtzWJZnJ1VnxOWmMZV0I/vXl1xCX
ajpvKsbRw/2sZI17GFc3+LpTrfdA54QXk7b32GsuZ+nWS0AvBg7BfK0P8tgDuiGjc7aRXmVwIVv5
Y7DnO6+kcKLIzZoEYM7SKHzwUaoZ+0gnTau/y2FYy5j/RmrMtCXxCprYRbOyssTDWkN99JkOH7+y
1G8OZ1j8fxGbQPxvdYmyNZm8zN9itTDBWSca2J6opNPNsfTVgcjx5eMHlHt/RxrxY237pBcfAuwY
hpDSPFZQqHBrLPxxjWfNqMKOxe74AwGNtlVSsHHAwZAf4mc6XFK/uMMNlDY1crJTNPqc6IhWgF4e
Ei/wGGyj6Ysq4u9xMmJPa39Hp8WPdSCbRuiTxd82wwq1lniJjSPx6RB+YPA0HN/OtIkmHoKyh975
/eQZH/tLu0Ia/v0mtfE2YgBjdAyqX6IrG/63AJWSwELpoRUZvoA83Zf2iZ69TyQs85g7tuR6fSli
cZW5OyLoC9PhS2qVFf2yOFs8YO6IBsFTfFizHr1HAufpGgzSDR8wIzG7zFRqFGgxb51i5DHZstl+
yVz7B1OR7Lmiumn+r3C8JlUtVOClj0FXym8gnAOniKdEURdZWTvYrm5HXQbiv68q5gU6MTKF1pcW
8PN6O98zWaEtX5L7D1i3VS/ogr+kFxtpl/g1x6bPdOzhHEBENFzIdbidA3xokFVl+aLHyfHH5lZ4
R0lnm1NhoqLyDYEYYVy2FWZdsTKGxmOEadYcIexgDg/yZvuh0E3ZOzzUDMJp63TJTW6gIJcFdapo
inmgu5vVQRye7xKZx+RxeHMUOrxmhg9nds34CgoW7GMx1xuz47LKHZbUf1mM6rk2ys1JzOj4G4kn
8oISG4aenEe7UAkqdB4cEaZvTLdSTLhVmVJpmFOk0KgtIhREnJM5AwaTFzozkuYmJg6iXYxOEgCF
IFoiNAdmZgbp0F4JmjsTJnOAqu9pR408Wmi2K4KVQt3i3Jiy774sAFrckP906ZjYFn7L5vnXenXD
Fnj5jSTYAzch2K0mRugz4xgPJODmSL9zJMVHWWGWnOyzWWnTGFr2VQmqvspu68oPEMg6AfEe/av3
vmH1te7p+OvmQ/lQoqIli5dPZ+2wBNBC8OqPBQiGgSdfEF2WBOo5c7VQy7yiMuPimCVwYKKq5J1G
yuK2HaeebZivsKRr/EhJUu0YGsI1UYiv4akwy1da4oMsR8aczsfHXdDF7AwAqCCMG5uiRQiQPVYL
/mnngMbfy6+uZl7IGbQMt/3iK5znCMw5NAPBfdGg7HshYqGSAj3KPsZzQgcB/+cU2TkS/cPjnfMg
Al8BIx6MBZb4GwLvlVoi3FjoZ3buX3Hqy7Mg9Yyphnxa0eP/+v96paXAM6MiebOB1V8YTr4Vz97K
KcLzY2/AhtFRTCp41Z6DFWOtcsUpyvTC01idPZUn0zJ0hReoUKIf6Xkv/XP4uTIj9tzJ64m24rEY
KRohEDbuTH6pH4rkJ8OLoqZhUEGo0Tmj/efKQobYjqQqOh/Tl+jC/FknzWJ2+NJCmjkIrPv0D0m2
Ciy8M9mgnvRgvG9xrBlPS8mh71LMm+V47KBRqMOmuNdkGowp9cClgvFxvzL6/KqMMIPyvA76hqnf
3NrdvyOadlQmmsMEpdCeRvlRBEHsVg1Zs+o4HiU+l4+XWUeTAFudqd81O8JXNq4+fqsj6+MHnrvl
xXOU7pB/Jyhe0f53rcOL+79fpM3I3H6u5bUEa1J9qphcBNTmdOEstAXrj8mcZfzYtRdVxOt9w9yE
Fx0BIjMavTS1tDYC5KLgKJwU4KCXNKP4GVRmU1FH+Trh1EXiM8pOGRMzDiSvNnt5yFhkGYNPsE3c
rIMxgaBUoZN2B5VJNviq8nwcxOz95wKYCb+dBPX311fUEk+ug+r23y3KVrbjcyvg93Moa4yjSDFM
UJ51+g02utVg4fT+k0Xip0nexSrAlmPrn9r/mnU2FfrEG1Pe3BZpsRcdF0TjLqA6dmFNs0dAjbGy
AK/Papuc9twVcIqY6utiY0dttwZy2NUo7tpSzgzlTGHuX8V8To1wyVOTrPo2y7TduR10zoVrYc2n
Edbcstn8Z/qgi093z8umq8qwR7Cbun/HyuOhdd1ROX3euv24WiKNMN5Q/aGH2uAzKw023BL9euQ7
DhJhfCe9aPSUObMmth2gn6k8XRm8BszpSfH8dWmAwcxeuNpzxNFs7fInY0q7ka1rEW89VNjn7Jze
2EVc4ckrjfw4noxC1YZSTLyKcp+pHKTsLl0I2HtxjhFVcT3lBd9Ju2ybN5UyjAILoxZDzZj3msmR
GLiWdvkEsp3GH8HCVWdj+sHopE0hZ7KZUCsnfmGF41kxFweIlR6XescyI46R9awt+TcPooYDDSqg
0Hu/FCsY1G+9qTOTTnnx8/ugHY8XrFaFaFugglf9+4C5UlEFa9PZNF2faiu5bga7/NqdaAqFbAq0
go2htOhXz+yeLX0t9S1R+FVdPvIyOJBwOoJ5Mo0cjvxH/Q4A/qS4knYgRGjPNUjSJnu7tPsXdP8d
aSbWuXiz2/oRKZVrKYMFIRFwZRrV6bgIw4fOMfrxvTwQfW8ELVEF5po07PxO4MXha8921hR/ytxU
DLjCku+blk6tonA5l/R6MCySvm/VgYKCVzh4Ne6bqJL5u/WKSZ334DADnZFlUGOUNbAjhVySBLrp
8w8z4YTbOFHmcgQ2wmZ+vBHdayc0YxapjxR8Hp6uRzrF7pl8Y+qt6Fo4GyfaDtucLGGtW7cIkNv+
B24571e1UoBmNsy0d+709gHehmxeiP95JQSNUdS9uP8UcKF7InKlOKWpyOZ1+edvv+N1fgpXpypT
KzIj4AkLo0pszHFEvnbzvwKCFx+z1bhAD/HmNlNAz3eE4xF3n0dkyn/yqJGpkk1kRRLWeC3EMHrA
Xx3RnUx9UCbFS2Q9bf9mQWIjOezN0xlcAt+licItr/RflLDi+f9m/okLa+pMl4l6PJyfFs/MLn49
XCzWLkuQQh4ANBlp5EUxh2mU8qP3dgn1lKh8yHQdCjQQm5zsCeGW6zoMH1GrzHtbEZPZyYXFoRD5
mLyAaiuVqoDf1jZ21ABE9F2PJ2cDwrubiTztpXHb5WbFZedJKza17wtOB5MgAjy4tZKb1eQpPQrv
NhpiOyKTgUcVjGyooP/F9DcDVUROrQKXxZXfZ34DG7W2mPllqlYvekeZYToutgfM6S3zazgS/gcM
htO1wz+6bru9YI/qAQxmXvL0Tad7E/RS1p/gLMCRWwrpdGPRu8yS2+s9R+vkweSFBhRU5DRJRqYS
GF4/VzXkM1PhBL/5fEVTbgnfUU/PLmnkAOuPdQpMEV2Go9CyzRs/pSoZvNfoQES/8koIVaIUVE5Y
6XVzayYXliwW0kFN0GMDuMFT616YNLTLITmQ33B3B7GO+XZwm6EZEpJukbhhQGe3QkPaJy97wbhx
klnSZmvBuQ+/ZqUk5H/+Wj43c+Ados2lIU5mXFwCDACQBCOn3B2F1uhcPGQQM4KIW9kKbu91OcOb
FrV4RJZNTPgYo6gOggInxcUJeAtcmP443VL6hB77sa5ihA8k75lxjljPYuZthr/ruMqTA6XNX9zi
OZpmvkFamrI85sdMyRsPjotsSD4437rvSw6ELpopKnoR7zRa7nXakTiXaEAmY9Zhi/fmqbh3FrH3
nHjnNN+sos5rTrNDvjq6ZT/K7fQTptJgn0aVB99wHH4MmJVTeGQ6JghbNIoW5NQtITBQ0Jf4RL3e
AW/OJL4SqjiN2SJUrvKx9mh5rSzvVlK/jS8yguHxi1NvDCaxHgTuyA99rm8lINSTTHLqYRQPEA1+
6bylgaz4BsXNWmi068NGnvDk1kXJ/YOAcIAyFpAtcQSGu6x0tdKsV+j75Ma92Jhu0wPc1tvBJb93
bHHh0S2skNaUcZPMdLALQC/ECZIgOGhXslQdunLH8xENlvCCwPEjYtLUVc6egncrmqSqx2Z7gX7T
wMdb8HKdj1BhM9G4jvdZXbhf0kAQqDA+iaojz36RNBAtcLRXi+SJ2oDnclsVaGOYm3er5IgZ7vTx
SK8Vdr3AxnwJzJZ7sIoZBp9PFLhzIGEcIor7FtAPY6V8NyeqVwgwAR7cerQna/iWu6xhGIGieosU
yP0++i4+l+Z4YGp1qifuvo5nPzvkPvTWMqIPg8v1vwB9G1OmZifmToeME8eahHnmoeujCPQw8L8A
pRsweVhfP9CL/h5mPf8TeUJiYZu+XgH6BHBUc0F7B0hTP6hZHuhW3otnzrwKfZKHIy6fSF03IGkr
/tVBERpEgRVGH/KLeZQMYE/WYWq1v3gycVhQaQeFK6EqI7UAJ69Iyo3scaMVHro//1k3CDh2qV+C
P46cY7XIgwSkLopwz+fzuDDPu1FC7LH5QKlbRCWDl/GbHO3YwAyIGjmYNyrE6tpKzy1h/sFw4f0X
0xYOxwBokUekl+s6mfVZy0M8NHtFF2R1kgsK4VYKKfJ+kh7axfARnZm36y5dWTOa2p6A6hi4NgEW
In/IRaFX8uiRhaz7aCimzQ56V+A9rdCRy0qHJHMNgDk3YKeFIgq1I//cftAO5oUjDslYA9OzIo4q
aRfxGroG+IvGBuHlscpkiOLTsz8w7+huL/w3Tm9zAZu1MObMsKKZn4WTgXqd4cnhIBYnmAfBVnhS
ARQIwCY4HFrwV9G4hdv4emtILuX35cOJDUsF1POznjsJshpYNlkAiVmYPQLRZI+7nOGfx+YNHE15
y3viIt2SLJ2IodTQ2a8RQz4u3MzgcKG7CTlwZt+bQk1vsjnGMoMaCBykmULqwxXwDoehBPqkQwjB
vazcgN2PNEX87OTNK7ypaNROY2amFpc2XPyy8qH3rkdrMYLL1vNoYWIxfqgZR4WL1bvQVnQ6dpgr
vgn3xwlX9bP4NW7pRgBlcfQltupwQUkxH0WFEuAO6FhuUQkvdV/m3CnQzQq1Ex/4nbks4bwu0Bjr
/798mfflkHbVI2K6FJoLr9jg0x5GB2aGlSPAEDcPd6rVTC9JCJm89VDE/TOtjUMANR8QlMqTYpxf
frsfG+Eor97uW68vsZjCFrK+FKVC5+YeKy9OuvOghaLndnts313DvYxC2Kmv29gXhrFLe09QyYDP
iSR/vglZ2fPhkhJXQ1kkg/xQJ4hVeAgTRxnoywQmWw6Gmk31mUek446XGUAQIHvSUeNXMJ/Ivee2
yt7WLMAuYRfPBp0KQA0EihALwrFs16YJ220VL25T9IGrlMrA6sLycaJNHGxy5yHSEIOWIiEMGBaR
fKTPinrwpvIFVFcLtluhD4ryBH4GYyasQrgogKe7fZbWDEUgflYffIeCnTNrhr+qQPvTj5QbI3ck
nn6krYGoi20amQYS3ksW4UkbH83oGYo1STWD8AM1mBTIMCP5pQ/6h3KitXqtm3JeZw+FgNaBGnnJ
qasPF7zVg8ijCSK/EXsNatuvHQxMbGabCUB5NFjhKpQh8jEqM4qqgIhTPacRMN3gH2DLLeRQlPJI
zQkgTYGFRRYjd7oGxCR2JfTtiIiSme82V3o69mIvgNVJ0jE0V76V7Mi0CAN4bECJTOZOPTWaxsFs
w0Orje6/uS48PzD4Dt/aVDTIo1EeSeXmM/rfJM3YuGJtogVfUmlMNmeMdtQQurU+k7NLul8h3Li0
uyNFI/EUG+Yy999rdVkjKp4Hk+z+96YlxeNWZpWhqg37q/32C7Z2+IE8MT18wwGiiTr5YS/2LOP5
XG+fRyl6nFBw4FkqYrQuVaovE5MEt2LKG377VcWxOIrOKsoVIHMbZoFvsBT5NN15RmIYnEF/rNs4
l5xSe20KF0mG/1fIBIdpiBECPiIGlJHvR8d2R9RZzk7kG1Twgd4ll2OxmQ0uTUdmiBJuTVA+6Q0y
Jp8Q5cGGxgaaAkhxoyVKT5ihpnkiMQmM6gBmjPzTrz7fgEmNEbNQ/3Ocrwjq7HJ+xuZXnuLJ93Lm
zlA6ygeTJFG1m2/Y56Tq8Y5xQT/e40OoTV+eJgzWPEcWxGbMVAPS4ImV3bov236KDAjxambpqfIH
TvkYeY3FeP54muR9qh4MLQtecR7zIi18XSaO5ybMgwLMEdSz78KZzI8UFC2E2G1UOi49oH+b/tDJ
Jnn8WTQoAw9mnOzt0vEqwVlJTyhEka7dFp7qd/IlQJwIp+5+ygzhFe7CE6YbiIwcm8CnGL9tPEp7
zzPcocR1vCMQSWy2w4t35hkeUzNPBgz6q3UIG+RdSjntQONLGF7EAjjs2L/w6GKkCZX36UshJac6
K14niMOqPCPU4iiof1G4JJQInBunAR3/YQ2iGS9T4+8PONZliAGHjuC7cVzS8fcrphgAAHTkawsT
c29Efhp9EQHw9rz865ClFb9er1Lv5Ag1IVraQhamb86vS45ZfKxRcxKF0P+H+esJcrBPV6j1rMuC
bkP//rhZp/M0Efyfrmx8ET/6ylu9In2Whbpb4TexyIzcIcpNQzxDt9ylXZLYDDS6B+ibstr+DOJz
glgdxyg2dbQCRs32ISqbbfbO9k+Mk7qOsWm9xoIZCu5flXd+8uVwdYekxrV10vGGP6bDuMA0eky/
ceiu0SUpIs7yo38PlCU+PnVT9yistzDP4WcQImSKdHFSFS2EXd1d2v0GwyhwhddrZFIvk2ZozTHR
/nVoHIVM27Td8GJnyRRb2kfQkuE+QZZAoS36rTXvPnYfS3Mx9IG91C8CKB+EdO9Lx75pkC/sMxfa
JmZWSlBuzhERg/gqbbLNRvcrJXxbQrJUQVFGR+d06HrCKe1BxkVIfjHpWWvYlLOSPMcG0qPM6Q62
8M9UvUqYDV02SmToifsQh0kZ71M033vPy6cNNqcUE5Oo8zWfkPH2z1IKB9cb6aERyblMJ8bvTV4F
5uJFrxPhwj+ILoyC0aO2NWB1EkGUmr4MfZCpa3fw70Epj8e6LqCjK133Mj9mY1uUP2Cix4eQx3VO
nL6ZbzIPRdL1nfmjEOrbZD+DxCnvzn/j7Qc9YgTq6WmxXoJ6rwX+6kxnlsDbIMRO8kNsRv0MGabf
25Se0nhDIiy4NjJJdosEJymCMZ1zdyBRaNl0Siba8YZmjg8EjcRXGGKpjSb2HWm029GgoazFF6YN
3vrnHfZ4eECBJBTPjqK/TUEbbrjkCEly5E49XVV9WIrftSO+pHAnl7Idqlvrrz1MEOcz8OFkNxJ+
F7ycqLVuzPldKDoYZLkmzdCYnog/8OewNIh9JZ1KOsrq0xa4JlaV4SE91lrNTuH4Wv5nuoFBx6PL
ceoZGwM+rs95YPqTVYO4Sof5umOsQAz1EA26Atdh1ykOKhC5PSfgzERvqSJFrQwSpASM3cMlQIAT
wV8hFCO9DdCeMcw1UvgTkhXXm8T15JhWbNyEjcbsHEUOfwshp1cQzHZpz3XGKpPNKX1GUcLMN0+V
KlCvE7W1yC4sMfW69Am3LYo6/JWwqsvPAGTClaDTOn6yhzUtRPrFC7RZj8b2v4qaew30DQPj3+bv
BwTqNA0aeG7Np+CKrqJQVbMvtlpPZE3f4kxDQr9Vqs/lo7o+hDAX7wovaHkL1o6qFeYkwhEIvPhn
17nSgJPZ15htwft9kDZsmc/YO85gCBDgdiXflaxh0j+sxGm+9SjxuS5FT0nxHSKblU98afZLvMKB
KW/GqbJ9VaQ4uuf0hYH/nvDXInhoUrpolu0XDv4HkYYCJJo71PcDyOzsvmF5QezOhpHlZmfrf6x8
G3pxkUOgq/TLK2tM9mXrTDn+d/aGaCN+RyxWPUYxy9CYlZCisxTD0+1TOCKtbp5VlftKI2pZnJwC
iNHTpLvwUSiRLt3+F/xQcaeQNdIZlMsN6+a2HRhkG+oXmginzhxyWWCu2R976FSdPMP9vBYSL/Wq
uKw6ItRxqd3rtoaa8ouCaaiNpNQPkPgmbNQ4OU4Gj6yF+xkADwNrhB+amDKJxvOICq3m+EwRNkjC
yAoOx2SI3haE3SokAlzo9lvUVm55JNC9520lwky6zJbtpSlxdkF8ol7rv7D6SYE/oi/+V01J58Uj
IfidFPY5xZQ5JIhszA8aYXMz0JxSij3iJHPuS0Z4L3GOI9KkQSzfFPzoHjDe8fJ44tvAJQZQCjLa
ySu3e7u7wUtxmZtv6haATgNSSmVGLgRlUN3dzimdLBRuohHu16xGkjEO5ams+hlVKjLHYscUYyq5
oWPOsKv3hd1DEqH2bStc2G49Aoap2PqyXfgyTH31P/grO3lRTDA67/rAxMNmK2WEcdhwcPj3CGS6
37KujgplRw8byAcUc083jxlCeV/rmlzz5w1+sevmU5M5VKiTpqbXhUnZ2SHKglPKfKDBa4QeJP8b
TzjExeSc00jf2/EmNjANOj5tRnV9iug/dMbMeRIvtP4sLtM4DMCqCto7IuVyj0S7UJ9ZyvRdi17Q
WJLAZtri3f1uwQAIF/DF+50nffvsls44jmASvgZ+h4ePHTTRn9nASfzqMnfdQIcHaAKKYlhMPLvX
MQ/QEsTvIV+6fEMC1phsPn6TpdiTkngXQTgV7SWjPQBJGL19T6jqjrKoXy7xqNOnekJaZdWVClIX
C6o6hiv5v16y9ykHUuFz4T8K8323ctUKUV8snFJVH6bUqwuuXPYX+KWCyropwWesvBqGJou/iS56
F3uCOahO7uU5SVGxMaEVTrDv5lEvoLMnqlT6jf7RE31fbTjr/KxgYzxurgWUfE+YemdceWXuLvjG
ZxnffkEpToaK2BHvbr8AFbPy/mdfdFrCzgpyJlObaTeRjckb7fVZNOqmO6xA48BJmDjWJ+cW19Li
QIhQxqzcZIjgmR0l8pzDZMiHz79U0tSvJOC6bLNhT0RkI4ZVBRgaw0UILRk1K6mhsEizFz0VidB2
GKajxtVnI4Ah2IRmbJeKBGDylXCqP49fjDTf6ie+Joqu91Eo29tLqXk0FEAz1/v8UQ/56hpXLhFD
CbkCJu9LHIzvL0a3psvof4G0cGDNSrSbskZPs2t0/EzewBDZ7wnPhJjwMwVx+MOwjoKT3b8UpRZw
Aoqt3kHRvA4hYXY598yaVycPY0uCcT2rkgTHj2i4sHkiEJ2B4BjOac/RAWOrkYziGuBvkY2B7Aym
X7V0acUkgt4UudQQ5mM739xICL1rAzQ/Ud5EWPoViAbPrgjM50URhkovUOD+iQVLWBbY8aR16a6D
0yvrz/Efy1sztRpRyEJjMVb0Z/ZcYfZL7LUMznhLZNcvSe5q5K0mqWGnlRXJYP70VMMc94fSi+zM
5rrMR3/SWcYyJF/QBA2cl/wy6rQEGuNVPXnUYrpT+11NratwbcgJeuMW+AcNTkdDI22MeFSI+BPS
p4YqavmCjpZD516Q0Owmo1RvJKnPjC9WZcuPzml50uc8m3KusYOd6uYyFWLGoZuR6ofJmseEhBtZ
L1Uzgbz4S7gV77nZ2uDS/20JTVgwc4iTu5uPgJH+I1OkicWutCBbw4Cbcf3ZgiJgYTQGn7OOFBPR
b0XOWFSIxmzChzw1cyN32ZAmXlwxeHBGVHK/hMH8BkDt+/QeT4kwrnrofDqa5C+VYHa8JFeWg9eE
xHp2//qdv4sQeYV9hI9gVKy6GRfQnoxNN54OUcE8S5AidOXkE1SCry4gSbk2wU//BxeyCdLxc+fe
EIr8FPJx49CWyPbwg5pRI34UzKWXb5OUSa14M7ASq7LHU55zfke5PgjDTFCWf3x7PuaQtCt9llp3
k2Po2BRpSdIonukWwZcZsrPkGfd8RgYlZExFcm7mQ0Ukx+cTD9b5MlNHXxlCQZPjUFHyQRE5yr5G
UU9iIXDBE42aUoIidivObDNoEsHLMTi4WlKsJt//2QBKBc/qww666o2HchvL1YaOeMrArz/ggh9H
ismd2Vz1mdolG75WIZvos4Ss7dK0GjROLtX37yUcVk6JvrF6QAzi90+IlP2klN/q8DX7cu5rEgL+
82KNUX0RzFPHX3Y77VNKv75bdmo7O8nGpyONPFBgdA5+6Bk+BoNRyDngnEh9s71mU8PoesX8JsJa
kzHSYvCFbeQ7U8ZQMkRcxDXaVYNf9wA3mjx9QsoWRqxbi0ZmyAV53rhM9DznWY0GEI+pOqnyNdaO
57jqkm7fdCwNFH02k88G3PWNoIW6R7UPMsoI3k2vFf+BdWIsnc8w6giuPxU9DzwrJJ+EVYxP7hNA
lz97bMAYYM6TIIRv088HAFwUaL+ymQqrPnq/LBJ000rL8IdpDxNim0j0vIRHRSAo4NbGIgI0Kr20
8kmqpSBRMAf5prNC0gAZeGz4R9/38VBmAPkYaXCR/2B6sebvoc7igQt1bUuFuMhfLI5TSt61S+pv
jjMP/1IKFbbrTVMag0Vr27OykdWpjb2C97P/mh7VFfnLCONIaQRI1AvhRz+4z2kNpC0H8CceEmNP
UbyC3aXdYWZomRkICq6REN0vYsecAfWu3mluihB8Y4BCypFQqX/ccm+FQHWZSOC24rINmWtD2EK6
03jlHWMyT+XZBvh5W3jWZ6ErPRC7IfBgqez8KEz5CA840nW2nKRTBv5GN2JTdr+3BCnNFjWl6Bjp
pSl2NFTQDPggd3vGVRCoMr1OyDBIZvBegIVkTzTLu0+qxSBczi+TAgxGEHoV9OoNJI8l1EzAeJsc
kXU6J36VzI4YCXaxD5iBzUWkMnoc0xRPjZ7ylBmoI/GDEWCqB26WSegdtEh7PX1GRlDduBA50M4H
qJhdf3tHh+ptNSjDyz4m8VKKlTI9Ik6iDlFAyA4L80joXaBXgva8bzuxUYDtqpkXYdLJrhnhS6b6
JCozDwEft9H6HvOarvRSbSvAmHpy+E+Z1d693OGoYi9ojyGpPFmKH4O0/oGNcMBqdLq95nSJeUbG
+8/+r5Q23FdVWPm3ZsHWG0BZSj6lJk6zJySl86XGun0W9Pb7+aI8XTM4l/4uJTzgtu6JsespR5zZ
KcAa5jgcvDxvvV7DQe3Pmi1HmCBAaoD/q/FbPZziUvkNngs3ofI6Biz1pVjeEA1zoll/qH+EOsp/
veFTFGJ8fN9FWPwgtIZTtDS3AXnL8H5WYoVji22eNhjG790xgZD6Nst/pdGg1Xz9D4zFDmvg9tO+
UvAv5tc+Iy648tbFH8uIGpbpFBv+z5ZDUGGdkS01yOUs4tKMIDj1cnkYQcv7BvBR/tKo8lg03KCU
5Gra+PlS4I1tGjr2Lbxl1ej3rn4BObNUeANMqQbPuEqUqUIDo9sCBqd0ZVUQ6WOXU8cD6GrGShCH
KfEJ4uKoa36czoDwsEXRRSV1eSvCC+DZP/zRBC82xhqlbOKgs5uTsdnOdJl2bFwoAkjeppSZF84U
O3I/yrYjZM/8IltFHi5bMFGKYMy7Z1i4C/4zHYhr8pFLGYFLb3HteV0PoMnBSP64rgeb/RKwB36T
An0YXfUBfXVjnfyF1/8lPUUrbRTCrfNBmikFpWnPsg14bma2AojXyINaAHskObPQG0VEAQNt+emn
mM1xZwS+zJAVkak6fNPP/Q5FAq858rFPL9T/kv+SptZQiOYy1QYGJ1HCxKArz3zuVNnsrPyNR998
TJo0txL8hQtSjlO+9A8Cq6fDOyRbp9a+zFApw/I3+OZVfkD/1fE5J91p765siZfDb9M9nz2Z2/nD
6GRpjm4H9d3ndzf5gFnp47UgpVpBw4CwvnlfKbxrYxegCAf/c+jl5sT9unAvxg2rZkd/vKxIcdmj
H+fLGQnxHZyCqe8HRIt8e315fSTKQiOYU2cEsLqSKliOWlxm5Aadm63mJAx+6KWs//YKeoV93giL
rngDAPmF83XXMeYWueNyq8QSuvmYK/dGcqEQf7MhTotYW8nuMYWSEJmOFf7KmsAbrRGbQbGp+n5i
N1ASGlG+jhiAcQtjZybzA8HNaHRnOv8LTx8sAnTZZBp45kQ5TpORpBk44mkADwmIo0hSXdlcVZ+F
rmjaDcFavYVriMiRCM695weJzi1K4fWKKmOXcH7azn31H0kd1Lvl9BEp4NW0S14oEcqkZptNtYZa
8fch0qiC+HbfBJdP4CK2oWrzBwNY14+wIqP4Q2kHx+4GOj27WZoa6a8RFBnAqfYeM7eBHB+v9ci5
NL1u3XnrGn9wSJo5YAfqHL4CaxdOgl8I6UDP2I6x+0g3Cyld2yJY4CiaOYBbV7PMd/N5rngAOx3s
oIHauZr3t6jeKO4psyQfso0qCO1292+LvciMshPDHZMOg7XZybhys36k+k0SEyQzMw/W11yAEOBF
8C13LfHCljlkk1W7xcT6Zgl1iWSkRbMeyJU2C8gElYZe6hiK8mZ/qpXKL1UtPTP7Z1G2diL94vU8
KWtQKXGnJdZ9xEIM9PoAEo/6wtuOR9LjHIDk0Ds7Bvbt0ecGLPOGbFd77UhzmmRpIe7iCw6tScRo
W0qE92IcZdOeU42t02+w5IRS0V53Va8Fz/9v/oS4c4cchlhUPTz94sV1njyYjrBX+pjskFXkk68K
fazOtkqbf618oGMSFPEIFY7BbDll5O+W9OASWo80P6BYeAbq3oNv5HRlV1KBugZawtGzk/cB4orH
I7q7zIe6NcOAUM8HW0ZzyZciADRWiB5QxEcMI34GBW07O+KLCTNjkmXw7yuogUlJYTxslh0qQ3bi
zr2fwP5H4P6+YmG91Ad7jj2gc+sacvyVRAkaks4MG6TI0TvcoGE0Id6kr4dsuJRjsulzNVYH+pXg
XdviMUuKS2Bd7F68VTrvGpUZfQO7o0EjNC5urNy3IL3005oW5zSW2GuaYNGsFa0hJa68UkH+OL0z
riRYCAPa+VDJs56hl4u/xhHusS7AnMpA/64eueJTwpoljKpn5hHXgYT9X3nlqeqP4Zh1P95n9naf
FtTgCyVdPY82OmS0AkKw6Et/8jnFLJ/KufpQD74qI+wp9UxwIMkUZMLKRnl02AEKUWnGDRzvVIYE
Z1u02jVDqQVs+NgkPDPl8xmgwXkicP/ktWZoGPUVk5EYWYg+pcrCfIp1SySf/vlWF8m/ahDZH+mm
RtU3/QI2MZUhTjvQk5w0SNztvx7UDe1YI/ZS3J+fUEiTBwlIV9L+9zVNfgRU46qCOfYV47dDoLpf
+Z/ZlGUwSOWMTshSyxlyrl9CFuHjQDbolWZu7Uy4wYPMlHTsOR2PRsnCQOAbb502Wc+Wudfm0S4b
90Z1TJ05s7gSdHONu5ehnO/UH0GPJAqdd8nqvoQvREFEMjat7C/UjftPKRd8RolckBQiHT275gCz
GEGFgw9uPph1PjS9YDEgmvwndrXKoJcUMtCAddBrAtvHuma/UhQuyw1Pr/fPiN5qNN8tJ8s7p4h+
lJATZa4HuemElPYfBjJS1wpyPtgGLaQYEwbNfmuQ+R1ftufuWmqUIGK5iZKT4eeU7u5Mh7i8qDUm
IZgxK+OH4JVfopnLrpQoI1oo792U4mWRITnXXIoj5TnR+hnWXu5Rldbb3fmWeAeeIWdZdhceFlzK
v/SwdUpfytxSYk7kKtB8zDnWkdiiXurmnEOZWVpK0edpQp0W4DbPhNieZTNy6Z4Dd/PvGRrpYyXn
hlRNuKEM8H1pAzLtH+Wu3QsrUY43e7FyYYRLd3qNV/VlH2VQWXvMrSYrqtFpaVXrx9Gft5Nanhm+
feBLSk13isEohBZF9BOvyWf8T06a0PQLSKVV48/1ttENPsaJElTGeysdENEv4s/wtBAQiZz9BKfq
e4Bc3QUSloAIg/XLG9QxqW/y3b4d+YWqyJTFEzBw42FgpB2xWTxFQkN7OuPGm80ypdpOdZKayrEu
ItZi3VdrUtuQN9WiAQjz47HH9DR5me4aLhPRJSiG7ozcykorlCRv/ynvC83C3dzgylnELykEziP1
BqB2OLZrlqZq7YBBWfmGovCUm6ZkpvBiwsCctuIy9Ju7fTFUp8CG9pDQD/WC2wPbIe/trgbKYC3I
l44/6rNm7+PHVIIW9SE1Qx43sPPAMBdxFiul78nZC3176tcyErJGt841ocECBPSf94ays0AZnKcN
e/OiJq62LFA+JOQkz5F9jDxv755ZO8P55QYYIcFvgsox3nva+Ytd/e1qeL3vlLOiB8NV7YprwJ67
SUwl4f27r8yZ8xKBvQrUogaO5rjnhWAQX5IeT00RRDzO7UJTXZp1XoAeUJdk94SNSrO47blr6mSt
HA29PWauiCfryBtc0liziF3vALWFHkMzXdFeIBLw9gaMqe6i8skSphkIzmySrhqiLLPgmbSIwNEe
PVUgcJLa+m7ZxRfUCdZqA4foJwg6Ez2P+wlEanDJW/iL8+iqVtf5g1LKSTkKjbiWGNuHY+DYMRYO
25EjQa4+Agpz44j2lDRuv/5BNlrj0e5lx8uEoR9JbrCK1hPPhRx62I+rUflaBS88rCyRRs+VHA8C
WZ+4fmfEhjZdMpInJs+rg4AQhJ1LJFVJJ9lonBFv9cD0kVNX00q5Y4l86b8CMz1iqbLmyf7AH06Z
5KAh6QAkaHfnwfbYm08wLjlAG2sLXXP7Bs382cypHyCZ2lssfDrnOBnE14u9OYp4AGYCowLCetKN
e+UqpYgiwStnFNQP0kgqs5dKyP24kEhI01kWKFFOgZOnpd2FLEteQdeazVRM3G0dUpZKl4Eai1rz
iZ33dbpFjzPbTeT64mAEfSAymQg9M3vIFbuGV+OdHeNickGFa4pc6qUcscwDHytguFtykAfRKGYq
omy6ASxqKNYyAesPokg4VNT3I9zuf/QqPmNfGctCpfgG2H+0hDm4RizouuAWHNlbmq66xIZrOb4G
QlNfDETvSScOqye+j1vyz56MEeNMqbynpbYelT/zYD53H5ruY2oG4gtrIVLECMBQdM6GKZBo+NdQ
cv7JzLQcbgMMUfG4ciMgSGaxfhaVi3qidI0liL34Xr5C39lWQjDDVMcfRzJo49OHR80VL0zxN/qM
lzsOyypb5Nwi5d/hudBHSYQ9vuLmFvY9rPjxbQ7pUb7Irs09Ykk5FdKdi0i+bx4UeXAOKIftk2qr
cuOIwLafooI/IP/O3qiiEMR5JNOBnwH5Fbt99FWsJNfQlf45phNWxv3/kIMxOaKCqgyUs5BlpJkq
gQpcjp3xL8asri0N8q20K6lAQ4zZZeuivcY2mc3XrUANnv8voH6nAxeLroRlMvpIZyhtKIYW+0zO
R+p63El4azP0Z/ikQR4FfzyDh6f9JglzA0XpemISsbkEGfKhXSEVlu0Yfe4CV2S+uiXGg6oe5B6V
GEecROziuZealRVituOkd6hVcVPLiV//2r3+CsdFsBnADFBiyAlYKMtoHga0EMEtYd5m8MiVen7r
uLylz2teiaxTCPWt66QJ76TY9TM0xwjQsBgWmZvtQIQjiRFFv5cXrpLE1NLiV47nGV05YIx5Rgwy
O97fi6Z2tGHhD3vqCgM2tRkQcmtnCvWypSnwO4Op/Q4hfS7lGJtQCui9hR6DHrh+5V6ynkKdrulC
nyMBpQqyMBFpGAUxzcSruPcxhDb7L6zR0FSxJKfEFGDCK/p9uZU03e7bypSkZzhKWKKmvjfF2oRt
1iUOhQc3JxG/bIfM06ekW+dkejvXp0VUyndBLtRgb2i0Ofl5TXnyO1p7jDUJuKUzURmER7mOx0gm
V7sBkStEZbMgqoMEBrhiCHXAdTDjtQehREoymR9X2oqnWnja3JW722YgZu8lW+69HvRtxRsCmeGo
oqzj7w1I5/TOZF/T7OFIcMXYtGYBJSjVDxN72g+1o4sYYbDcwORwqiB34UBUdSELdiuKj3W0DShB
W7dXu56cIM4VvzM+cVdVAz3WMaC41N7AHXlsS7mUKmtswKmFA9nkcGR/zjfY4Zz4+6RAbATpMOSW
0aglnuEm6F55ZOQiPA6cgnEFMsTH+9tu6CdncZW6uEZIyDt4D+lSkTAh+A0VWffmU9AMzjYBttLN
7RI3Eee7NHtywTf5CTyOdMMYbiPnXs5G6D/xq9tWn2lZ7BIK2JwmplTGm+dUeaDHN0uBp2bYGc+t
soECSlxHveyY8eOZwYd/CbuICc5LEO3Islousnfq6JON2R8HvZgs17XvEyGnPWeuXmSxJSoNkxUY
vvwC0poEIEfxP66LitrDC5qgj/Ua70LZEyN4/eooJIJJljV4LXCT9uv0Nj1dBECeMBqhiT5iuNOd
+eKBmkJbd/V0ds1ThlbPAxulJOc9zTefAEkYbML8aIAwScq2BcA/LAM7DM6zvmur8ATnC19FyNEC
rRIrgY5Qj6IA4vYKoYDZmX0lG9W1X4EUtl9SuZnFgqDtH4qsNjCuqgFOOwAQI75gSdsmtODbZHdJ
f17bRGkiMgAtuAEI4geeNnqemS0QeFoZk/o0FePW91lYnvd3dEO6EaS0XGmJHqmSrgjIoydMNQdH
7ASXf8hu7dcN/56u014AiVUec/jIF2x1N+IHykDQaudcAClwQNlqdD/sN2WHvQeBlE/0RIHUEDoO
jWbHIeTE4RF6oPZHQ2XzYn85Kiz9x4A7hkgdRk3HftyMJvphfEIII6R7C5qh8HCBtgD+M4TfBggy
MjdzERwTOE5qILCByBMwvc7RimO1NEFj1xuE66rPWTSz8pCqruaADpLBDw6Dwb7FbFHtVqYN+Ecb
OlBqmB2W19CHNjK/u3QyNFtcFnzv6Rn2fiPUYb04Bp5DrFBqMEmwpR2kRpMO4UflEJVKvnKW8CBr
pY1TYFeN3d8H56hDfgApX6kGLdYva6bQuxXPsaEU2B/OYcxg1jOy85Wwv5xoZ2GQH7TZyJ9Y3xfV
9rePIa3J9s7eePvHm1yRl4O2ZxHQiM2zmqRBvrJgSobE/gRfYMdS2sgl89c8fByzJYa+ffPaSJ4p
+aRl3NFFtvBJlwrtBrm7gmwQZsoKBV424RdBIZzd/yfiWFJhhxxlq7zZ9XaBH4Tc/ICPIQZg1VsE
PODP+7lluPncthq3DDzusMvHAP11JAbQERaOUyn6gApKU4j0OwcLc2RQmVngB491o57lsWO+0wYT
VWMgfc3nEu3DfSwAGG07nhQDlJJfk5RnNGXVOsbKaXMUM+BO1ZvOR/IlzJVx5bljoQGpEClo3fWY
Ed49ZrOjSq2uUpY60cvt5dwQ4dluQFT3uFPZO2OPa/NTPPq+mVKsO3F0Lh6MFe8AHh/+m5eohhxb
LTLTAlqWzwoXil9/FhAfGRAF5M3neH4oYRyEPH2qT96K0Ao/rpsHDDW6ascjeNFbIDui7pNX0ghz
VyWQDBJIR3GwXqzU6q7p7k/FlXuib9jDcc1AjmDrZGD7AVsM1r3F0ILg81veSKSw+4F1iWNg84s6
bzhWIBz4Pn9ca8ddEVpCcrLN2Ev5cXemjK2aSx6kbO8IMhSv9ao5KgZdzOku71lxRIpR+/DByqGm
kZd3FH8VlG9MdCrzI1uoDy69lX2dcVqq/P4+/fVavgMX+Tn8NgmGQZIvdhuGQEP+5MQXIAwFcCUu
cCM24s+/hhC0kSijRdB6Go0wiEw+QKOcCWmzDeb4aXvhyaBjVgVrF2ajiWIQh+QONax2N4/9kjHI
h7vAykRK8RLSEmF6iL6V59QVz9cdwKEQv9+tCQuVt4QOZi9Z0NVrsqkFj8CtQ5vO0u9l/EiOPKah
6r4Ao4D+LKhQuNxDaAIvWK0AZBh9Tu64wqJgTGqJxW8fBRF/ciieobDdJd5Q5Yjc7h6YOoelkIqG
UiltWGngtmW228WD3Lb7q4LCW4a7GtbhnbJ2OViw1yIKBpC4sGWyIPuTVwYpShGqnGH582ZKUSht
7bKpA37EQELzB4uZmG+6Pdmv7TCb9MoPBh5/e0ydP6bONmwrSdYVWE5fIJn98f6LQPhQg890Hv/p
nQDdVqdQKbQ8farb8wCdwQPvJ+cKv/wkAHYVjYXSBUYcF+G6b6Ca2N1O8KNX+mIYs3RNAUwNl07j
WJpQnKUt8rQ3NA4ZRHG6Nfw49Ioi4r2v4WabaDibZkEdCXZIUy6g3H1QMns1XX1l+wvWpRYlqoNL
q3zKsmdcUxqTkOhkQy4wsAW78Ayleq+OQ62c4TuKoCfwZO7awKsHXjZx+vjRyT4o8Mp9Tcbahw3X
B+m+uiCYbRJGnufXoBHs95GAy+y7G7Vh1S82GdTgtA/m1dLJ50RidSIK691xbeUdIJ2DYBHyc3uw
2MEQoIklB2zUt2a/feMDwTi9Zz805I31xUHb/loP26ngwF0Eqh+dSaSxm4qwG/PWp7R8R93fDChH
q4k6uL2ORyYuinQXMZH5CRVAHWHueXBbZQfFwPsroGEgXq1u6MxB4a8RE+qnek75JnSgEAdi0Pw3
m9O5eUU7GNuRqLkwlE7vZiB3Vse0iHdhZ0wa+XHQj5BLrrm2Fkea1XdxTXbj7jGGL8YhZSK90jQ9
JrbOh8fWykJ/E59XtPMpqbKRSCQdngWGvPoEzVXwupkaV40ti6i9S6iHWCCMRbOhEgeD7h7/oPgq
TxDDBVbbkk+mtLL77iOHCdcGCSplmyzEeW0BHxqH72wDU7ZbZNO53AwggITrE5t4MsnA3GUomndF
LRmWkbZVmzWR6Iv+wB0cYu93z2CrA3jtsrDFsxRba2mSsXYZcbbLua/7s+WVQLYZD0vIGXKkhPtf
qIlN9sHHHgU1YXwhs2khu8GCXupCiPVhEPjE02IpRXO5zL4NRuL4JKqbAZTMwjFSJh7lWZ7ghV7P
h3qT8Qz8Qpx8HQmm7fhPmZK2fBKmHNpXXZhgphCAwiuCxLQBxzo/F3bQc5xow7EJvXugTfK05UzY
eoZua1wNeIkbBgOm4O/Q6AGLdgVofQ+lzqxrBapYPLbv5EC5KzyCfQ1xFV8G3+NUgUAFVKSrZVX/
rhaF4geuyj4dhKPDSyAH+NY+foZ+sYJbDDEqmKBBzp+QDhM7nvdJEChkJVodI62IRzYaDk11R9gA
Emd51QriKonDsdJnJ2CBB43fCF9hOgV5kSaZlNfD/utZo8xjY+vvtFXDNaFRA8SKTU20hQsu/YaC
jx/bZzaZZ9We4XsKJRK53pzyIfJEYfd8OIH2MhTowPuQ/xKuph9KenfRx9Vla75Czj0HRfGtP5zk
9Mii0Yn7HzXzvnX+DFAm60Yh2eDuCVgaYKKKNCgOyoRzIzz0hkEmTX2qUb5uDrC2APEuojUhCyzB
Np6dvjaiJsFVnSScJtBqVMv0BhE0aP4D096Zr0fNTvVE91WGmXWsQZts4N8w+8B0+4LyCfgETyrK
q1eGoTUIc0kYg9lzVI/O85yB7mVK82UL0iWqYY5jsOGBdFv0HvACvOO/N9FxiVwsgvaO6j/UsUiq
/f2RV/tQGVpxy4XKYYOCiQXCBF6aagHg5sJoOdUcXh7E2OzOUPmKgcj5s8s1guSBk7xXAOFut9IT
WH/X+kiWpQF0eBYXGdhKCGFnap0z4MpaDnnLtqoh2T9bVHXRdX6wGHg3pf4wrlv5XM5nRxxT5dK+
nx+Umwm561O3ru/zPa77iULfUbY0GYWhMDbt3zTg9A10/IbdGYEQvuwXm2OnZzN+ar6kVEs05tNt
LZQNPZ6af45hjXUXo9tRJ4/RPO0ySnVug5Qrpn/VB035+4THj1FTaY2pWK+Ecq6jezMzS3YEPFhM
e5/FZHW1zT6pu4usJYI5RsBtseaYFSgo2erymhirRwL8ymnRlK8rmjYvCYhy+ZR/0RDMyOIUdKK3
EktnwFxfsKmHb01XFd0kDpy7u7JB1Kzns0jqP6J53SlTL+q41LdtGLL7RGLagHexBby5mbApri4f
yb1nPGUHi2p+KDK0DGac8VdCnBVfKVv0XnubDV5mXJxYADnfjQTcT8HlbsV87D6q1PZYL3cXzSks
Vw7woKCWbjX9YkLjWwzG68A+EQV5T7yiA3CP7mTUjRtUQjNSiz5dzHRSSHZSVC5Uk+SnxdEUVZzS
u90Bm/XX9z2mk/L2pOnYtnSi+n0qu7tuPtfk/pHxM2Xr3gQsByloLTXaCuWwuSUQOTHWI1mojiLY
FlWhaDHCw86AKGJgHX56M22A6CaVxrC0lcBwejbP3SS3vgc/pmhELdjqsCCOGOFTJ1W4JsLB0K//
h1ALN5PoJlJFZOYXzeyfKNpNYPJjsjvenQR4PnrDbQ3lyFyhnzVYl94YhOC0LZ4XOla1535sr7ue
rQEzj4z++G6oOiMCocDXKMBLcRDQJuL5x/RXjdi6hGoNSBZpmQ402f/4QHIRiZbOyVWQgrgez6Tc
nTofoFsdqcJ2/OeudPM6HwGy+d+CjWYm6ffEvLOLRXakj0LRRNt087N52jszN+FVu52NHRnQMMuM
L4/CmRbVIrgcO6jab3iM7ace6DElGKmGwCTXYPA50b9dQ1+nFeOiHx2PYSedEy9vNBibNcj+6B0q
SPwZh+BIjKXniHERn/0xYtriQahsJtWriRuGbQaC6zpUdSKXCvkZtl+9GIRZN74jK6AST9ayvPYC
O5UshK/ncULffARQv2Rblqy14c2GTdel4ONSbsrlBf3UBSDFVBGwuu2LZQ8bdMF6FsmjGsZ0OYkb
YCqS4JeAi2GdB3SIh6BFFaaUvGr4G4JQvklodxvRQs8Erpwf2Xefs17Dk1mTmda5pTf7IfYtMqvz
b4SUf3vUeZicUdXYiLSQwKV5IjdEj3bMiQL6uObj/oXb60PA/Ui9jU/o1vLe6jPYjw98fHv5VotX
+G+h3CisoAJAfBD89PMhNn6ro5F+ExURhCB5T8Pziiyi85A3Dxgr+es4pWfyJOetV07UcAks+mXP
f/2G8ZrnBqdp1hMXVVwLdEZpnXGmFveM/y8exiyp+JyKoUzKPWTkdqwUeNbM/G38oSaiZDh9yzqi
jSZAREjzRWPGsJim5YNYCSZFsKkDJYGZwdXdhinvqI40tG+/dWGJh6Tyy0X47Xdr2c2g6G9/pSGw
Yt7pOApvZww+xdpeR79h4PmIf2Bsc8SFsz34LkHwaZVEAapxdnCIWCiKaUpdH6zqurKk8AB2ued6
DI5oxEHOmp2w/ERELPgyQelYBqbcIq58f7rD4Nm6QI+AoinTjpIGkfA5yDq3oq2xSmFB0L+lPe/U
YwthZ19GuEb8DNqmXKPwlGxj3FPbCOxUhhedQgqkIdHf+AUHJWVrj3K6/5QP6m7rkhyTDDeMhLrn
e0WPBcPXw1HptZTprsBaT3g+foTNJ0h8xJw7pCgq550qyrb3bKW81Gfcgvs1PVobP9440T2xSEGY
a86E1TUD9QfsO/UoZVWkfquMqLvFqXhgPA7NZymHdiFpagFQVFmAIasUEswf40oINaHPScJ9EzGl
aNEAgPNTHsXnvaEcLqYXYjefvnU2aqlaC1FbebqbY4GmRcd1TSAuTkUCnKjZz7XLdwq89e+U4SSR
W12njg2X3DNg/rAz7CgbQnTnLGNsy4082syc9iuWlLser9WQfB/8nhaCsMuQwM7kqY5q342E654D
Ca23wOEHiijBSgR6ZdG+hayNdnCTkt0uWlU2Is196ijhoPeWFM0gfxzWed0ZvB/y74fTUTesseB3
G9gBHUIk+UAkrqOHuXi12QiVRPdrFiKx9LGR1R+nQHnFIajf3QPzXl3PBuS9LuF2NjZDZJxg6Tdo
MFvUMIGNQIgWBMGBuxwiTHCmU1N2n+IWYL7jyBNEX2VQihVCOn7hrgcbiMz0uKSsx901fcr9ghko
c071joZ4mrBcwn5cs+DkWIRTNYq3QgWVq1AkkOnyhgdAZeHDhjwaXpbn4Yl4zldx2IuR7QNdts+H
CO/0ABpRFsISXAb3ya86SON4RQpQFCpnQiWtn5jFmu0oZePXODuYen8qx4nF7K52eTqxb4JgSfzP
PjsGlw50zUwLqH5I7cTDDnVYQRCst+XK+1F+2UXzHzZOWfbw7OyLvOVvRDtwEV1YQb+4lMrWHcRD
aWxubbj82AO6kb4KVHly4a3tNQANH9BV0E8M+j+bLQ1g+rfKo7ZjlWaRwdBYItvbmtJkrAZ1H0Bq
OL8FM0WCJJ+V/RcJJj1h6HYiCSj64MdjnkDz1X2sqgkSjN/1ceKht+Zu/bK+2pAMEKAxQXE2GWGA
klfXN/qsvZnwvYeyli6LUKCcnbedl2mH2plkLmrd0W/LQqprVDkR2ElG7Fab9R/3/6nV0qJ/KSE1
3sjD9lEX5KySaK0oZwbvRa+5hUPKl/Q7lvvUfSCk+wUX4WfZtsWOxRGSiMzGpii2aaOvGTauPwI9
blptf0CDCs+KgVDvA1D7GluDDNSQzOea2cETSSgtAdo7Bnz2wnwpuHas8vgDusklvKfbFpRMluJX
LBX848/o6ECeMiKLzkknr1A0++qjiwgzJlbBjaek2nXGogFaA3c5VTiX4TVOMXQISRHUOqC2Hu1D
Br7+OIpQJ8e8H6mES3ODRJBcqohuW6CVT84W77arbx2FLcxWBi8lFePJHEkeaRlZqMSv0DeCkLHY
j0NeYOLhg4AqwovGrcLnhUe2ddoyIArJt9BbW0dIVeNlhNRl6gI8bp8Jho+WGkgrRnNtIqBXt8Il
a3b5WIJRsfeuF+X8gDEtkGa2HvTerpUJrLwJgTI3q9JLi79EV6EiwYQKSrMN7r9QIroxQvOrQ/Km
0bayKXEkhJTUBrhcjbNTcFIC2c4Kh1tgELaVxbWV2ut7MMWOGj70Z6l0cmYJA9S5O5GtoivF0l92
ovfC6BhIYb76LcUlF5LRZIcTtDeOc0Lkm98RzAPfFRbAryw+AmtTRns3LM3WzmVB09EJO4nABImZ
M2O3iYETnavckQvh6MaUXAKs4LyiVGcw6CuYdhZ+mDY/crcHEV7rvkxaXccuIodiUjZc8b229o6C
kYIfEfkxUNTM9VquTNTJgoGTT3AzBMaNnPstZf9L967sIKXd5VL9+HTjGvQ0JvoQFa3KJhHXsc0F
qSrmGAwNiZxmurfyF9R8Rrx9pDWOGo1vPHuFaafQvusjTszix4YBWEg4jjxDZcSftkPCDYqprSJe
y94BLg1N0XvsW/dSNnzfmDShWAi+KQ3bUJ4stUDpIP5l5zUa/sBntRf7+oOk2lKXoC8V6ZwMklcs
4STQc/5IUW8ScIUEhkRDuWnXWu8r6v9coy1EEPuw0Mu89R/4+rpG8iplwxgp1SL1XpSc6+4H5m3v
oXg4hd9QS7dK4wnCdUOm3M+4sv6RlnsSM5bNsnfgbU+9Mh3+hzT2LUkcx9/y8Hj3RiOnbU/I9mub
S2t6wpNyxRtCN0pogUXDx5XNQu9oYg3oKhPegfwA4R50FYz5bW97a4UvLlZ0bSdxS9HBrRsYPtzM
RcVK8khNlPNTpbdBw3cOY9/eZESIn3meBVAd1WZBh3OYOQJ1hfGiLAEH2WO2zY2ObUDWjGBebzGx
l5ddUDHRMzpxv94jm38xjkhgPUPI3SXcl8/p2NPWq1X/GA14lRqECVjgODbrZWDz7MoUTM7Ifrcu
jFYXYrUO5jZU9onQodaR6KjBmVkf+UFnw5h5Je3J6QiFPut0zJbyTT7JwohWXeStzWivRwy2/TmA
U4vqligJml8p/Ufn0gPsbNmSRWobF4yHfYeSWgvhvboYu4m5yqwIxAH5lmGPfnxPFqnwa9DT1nt7
Ye3vLJjUjZDUhoJTy/A7LqrPFsZb4oN/u8WbMhCk/UIwDoti3db8xhlkRmuF1eGUBP/IkEo3fj0b
CpkrWKSOq/96K1WeAKTRmgc+Cn35Y9i8ccSPt71ULyt6xIfimkmbJKgtPVTIs1n19MtNodNh9oVz
93DYfA9haUYTzREr+6h7zIcbO4lm3pMNNQue2TL6+zs6K2eG8mNY9sA1fJPC8OERHNNQB316Z8Gn
bqWQIsnXcwT5JzcRAey8wRWbfTikVnU3itO3nkqAzk61P1ygSgr+bpQg5NEePBc/D7klQ5rlpIj1
SwzFpH4RaBfCxDstpfOB87JQNzUk1s9K4jM7SujfzfuQWqP6Y9DOyQ0mALw3D3jFxsnm5jfXhzJv
azvjH2Gt4jy3tMEMbne7j3Dk7iTKrNoDvE0POim7sF73j0gn6FgQE9nBVTU0nvI6a9t0VNa0vn12
IJRG4i0fZmTcNZtOX1UTPyxvdDXIyUTbKX9VaGBO2dH61joSdB7NVANMs3F3OLb5IbR9zzAxvtgS
6lUy0nOaE2xU2AbNd5OlI/19vzwYZ6j+0so7mlYtgsX3oADsmxm9U6u3cxk/4OgBvzkHvkkQZ2HK
RSlNjiGQdDJB8RM1m09Q3Zm+wlIqn3jEEsTVykPp+951X+VHwSDhCecmcHVIEXE6Jk184/9N6kdx
LLC8QBwhtSdRdif71rEiqXu2hJj5xGIqN39l3cj4XhtJMpzIkVW9rntho02QVTgIE152/QPnIpPv
wFM9dLfGRQxsWLiX0o/zor9LSNGiGeR0RWVkhqd1g6Pq3bbReZXWZoWshnkmI9uClbEh4Su3S/cL
rE9+HDCHTNUDUB1B5eakOv7NkqYf5mCT4MARs8r9Ht24Q+ebW+PQpyRD+O4ov8kw1mWwMfDLnwJO
JfFHTLB4I8jxzdksB0jBgNX57FgEblepZDbiLhpjTErSumQYeO+rtaMlcEimftjji7nB5FB0Bi3X
dsrT5wC0CAQDpEZxuYuSfQcegT36+VE9MqSuR3xcn8+dsf/Oq7++pT2itnv804mEio3rbYokBblx
CG3En56xwjOg9C9IvX3OmEq4frj2a5Ech91rYIcqTnPYUyQlG+4+CtaOFwlMi22F1Ot2jTscu6gY
nS7bxpI09gdpYhnoW+cXZ09/+C326PTF0/TwOkVAp859NfLnYlqyMEmC1JNEAFh3K9g4MAR2PJa8
nmKwJf730AOgasY2veMVOTLWsZh3wCrOxYk1cPh1Qp4EX/kr0Nft4Iw5H7G8ex8HHP0pkr16IoGc
KIsrnN/EfLrntniF86GhwMq2Fl72izHDd7rztO5HM7hMB0+3rq22xBB8KN97uRfEmCxx06GGC5Tt
kUDMsNinZ9Vf5WZxKyan/cBWOWclBHbb0PfRvecpbyElyxFrzvvohUFZBc8ifzAiZrF8EcJRTmvs
nAPRzxKrLIZMSTUEAHLI1HrikNB9fff8j8hlK9SwOrRkbWD6wdy/gE9xT+CE/xZWefvIrjp3WYRG
7RAD9YY70gz+Ow0I1jJDg27yHCm7mwcYNOdAQkiOJeHQCJmUglzNuxlnQGXM5DtIoKCJB7Ku0u7U
KF5A1CSJwIZSbdSlVKyw6E2u1YdBHxnelfcXwe5hgCXGR0OddsTNxLqzqU2FXEbvhFKW0DIX+zkI
rjHuxjoPbUKwVvQkgSHDqpgA9Qljz3HBhIGxibLM5ENb2h2fvM018uO9f8hIvbLe+wGWKukrwoCY
aMPik5BOSBDNMyRcw9h5zY82+P4HvYWRILM9aW8bouPtcKl+olp3YmQ4amxNZzQvOPCqwYRk37Yh
PHFSfATpNTf/kuEMZE7w+MLTT+May79TynHQpetavrZ/68pJYrEMY+RUUx0JCuEW7pH4hr9MAUr6
Jygqg1ox5Op2tvdDZ4Xa8j6fk2y4bEGqhQabgBtbpI81xatPB3yWqB23Th3erSFfklCXzqMUryG3
+0VrWlzW9ZZbI9s+HyQIfKqM6ZC+c7gNGMPb9GHvHpZbLtc2m4r21oTdHXwOYXPvdKPxPP+69d/X
UhuagSjZQhm9Rq/Vtb6YB4f43uC743zpQ7wWy6C7we/4CYAGJAF7z2xT/PJ6BFN6XA+Ss7WvLqS5
A76X5hcAxIC1obsLPGQ9dzwM0wMSvCSSG9N1fXw8bzHsSfMWgs/3KsJPrcBRvnJSPvGszHHTdKf2
TJTBK4JwhJivxT+sqRsvukdYnb58ULuvUsz9kEOQdv2Bya6bWihFHpKLYllVQ2N/iyW/fyini9WS
fPgX0drSePSZUxnvWKAV0V+rZmnv9RTzAs5SklYaURLHNL1JSS2O0OUqvTRH48haz41JSG1E8psS
2zC0OCDleIRPI1E6iwaf+gQNdMBFjZB3GCZpLme605AlOqg/6w1OtUGVkZkETujceFyfr0dE2rT/
/YPVZs7JNawWan6m00xozqmNQ8mCRVWVaJmgCL72XFXy6nL8AbsjMw//cloLhk/kVEL1XIUhQtYq
kYZK669g/qqRcUzC6Xl4aO4FxxAlOEtBHlSRgGdupr9f3VqsG5P8WJrHZQTzzKpfYz8cf7pWxckO
rpG3Y7t7h4NjsS1ZM3DCNJfsUMN68h5vgvVKXZnbpTEHn/BOFQ0Ro59H2Ly3YBsvSJmCB7coOKzs
oTfPJxcBn97KfmpRGMBZ70C2Ye7mIxpHEd21gF/J3hijPBSH0Bhgi9B45GUKGmXhzQKhG/zbEoMr
v0TIWrdWb5e7F6jXwMzoK3SdaBefXBDYslLUr4ffI5dFZrUjB0FsEHccH/LYvGL4cf2wwAF1i1U/
2kdR1MM9JpvZPquJMejnmSYwTinRg2WVnK0TYdBB6zMf301fJUjDcxZT7dIWLjogiFFGD/5lRgIN
0bx1SJkaGLBo7pvQ7IiG2Qds2Sx6sfqFg0gaxXz0EcqXkpmHGVR6s7YV9uthxarucfTv2n7JnG1+
l+Ig3O3ck2x8ysn80NYick4dViUiiRsXmirMaM+75uSQqwGcxRr3K3c0vrrXpJqXnMhd1MJ+/u0O
qyTEbZlDghd2uDvesWsOoWGzH9YT+z1BOYHEmRQEAi5x/CF4kEbkfUvBKkdmzJCgoriSH2/0asgr
nx+tXFrU2l09ZrIPayCU2e0J2wzqNaWomvY15Q6J6FFHIIJ8XE14yIDF5M4O8QcSaDHMQTxBK6pJ
9a3XkgjtzIPWrQDnxLkxiizot2O0CG6y27zd4PumqUW0cebmkNrmShGKV58mJ/GONFEKGYKxlFaU
1HMZ30RSWEJVYOVBYLTbWyJhlfguQ0TQWuanWlNmc2zngmdge0aBkSDmTrWXVddX7WMGrUXMarZh
Vrpd173nN8Pe8++p/j/uwfxaNbhCCySb9lOJGBxcCdLPzprpr3zu1Q32oXYJ06CGAjGMdtTE9FQV
6Xfv8AhSGiiu7XrYYJzTEVhfzei1PWJGsOWYxKtzTX8eX+xAT4/JlUm/bqbn7Ojy0gTRZ4nr4R7Q
HuwCr2rDym+xe9XcPG2xQqJMe0ijCJEXkctE7gBXVMd0mviqWWbUSLl4uxKL5+DHkLkJZ8tyrOzy
P1M0bkBVqsmjjwHPPyOqfyUfFSbfgU7c5abHeXRUukBZan3amYB+PpCfgMs8AMeNBSiOTvPB0V7F
LWWme97Lc5Nl8xPP1acJsacuDVijMLGFB8f1SdkyGxwCl21fFJJ+01PELV7K88s8PaSA92HQP4In
/EjlH5sY+yeHOx6sscslyeKA1JEHRTyLT1pTGueh1u7BdcvOV2Q72CFYsfGsNckuLNnsPN5wCYB0
QfjtF6JS3YACg3Fk0Yqp5lOGRsJNj0xDAez0n3a/Q8URUaYlyqTG1AEFB1JBb4EXkEAeF9GTpiYQ
kqZYZctv9q/7fqTXOTvEmrPe8qEe3c5E/CnWdnEGnXIovp7MCW8WRQYKtJWcxdk+8rA/BPx4k0kn
3vLo4VRRy8zJCzobvVeJX/oJHtW3RgWzAnYwt4NqbZEAWqj2l7bOEjqbe8MJoZ4hbmxd+S+I8l+3
R3Wy/LKIVPaJNTSfYSFk2G3Q2UCUdQyVZyni7LkF8QVg8eQbbSGuMNlPfBzGeLPnhlPlmK5NFCfO
tTUZ7ySlTUmXqAVCKtc3yGdsy0q7WL2wkIcVIepT6M0+vpzEIesU9Fe8w3G9UJaO/OR59PhHnLUC
YG2zIJEQZvend9NSUaNwawltTGPyDslu0z14s+bp8Yzn/hRbRX2pvi4V9+GevszCc/v3WfZbyxHc
ugJ9sGqNBudK+tS4A2UI8iTX0GXeB1AaiZ3i9UMJuaKz+h/zeEkF0+oIGBRz/YGocKhSaiiR9q5H
1ubGkPxYlRmITKjV6pWkHsja0YfkHT5VDkOaiADXHhG3CEwEs9qX05Zw+nb2h7zOfclYz+msImQt
oXciG6h4mbOhwH5fr3HJZ5VbDq6Ij1+Ar81ZDkqsL+ChFtDm7dLvvuOp+vuwgNYrtLnNNORCZ8We
oYpWlsLsXzoopLS9DveWXwDoFcfh5OVpkamKJwVHfvfGQzcB0LbVOU61xp98D4RuXeMfUldinc2Y
LOjduz2f7l/ihVdBP+m7l6o6nZWZJgXM6aWtc5Ou6aJoyDv7uB3YT8GOxpqxFDC9D2fEhlN+pnRh
IGxBfu+M+N6FC8kAKqagtnv/JHuFvCM+L71e0H39mjarv/VvQO0FLm6YQ1sdSmbFDkf8++41VDmB
MoJ15zaZQ1JYXZyL9nOtIp1qOsVkIpWdnEgnXwWy0f0RHjNC5u5GZcP2S+f5PnHLVuH+o8Je56ko
4FjA5Wlb9zi4guAezQEPo38N8taCiQ+81gl1OGlEL8SXD2F6T53BLOUnliMn1Y/3xDAwQcPu4MbR
pgHAWDuQzqaiWBbzbnxug5S39K6WzZcaLaxrnSyNJMUZmUiTJohTsrQXI3WAS+tJEmFUAvs06YF+
457yO7jezm0cH3GQMaOlSyLRctArDA754ZUmCZbI1VanRsa5LPOvgyxa2k7syRTDyc8e8kgAR6ON
6iAFhaPuEs67p799GuqAtOQDlvNMeF6c+Ja9NHWZ3sqJVyI2NPMgkkGk/4nf0d6xZBr/yuLFOWK6
6W5XLBkhr7GnlupbCOYrFikPsOq3sw9CmQ9tvmJo4+9PYarsIaYkzr9NG1meVJbYn+xRJlRTYxPm
JkwwU2Neqkb/Ok431pSLKDyLuLn02jbS+B7OBx5fOK6s1lkbrbCDPaX/H0NBO7TZ/eB3/AR7px+a
hI73+l5VZl1GiwHFlFPZPU5qERJGrNSF0udl88+R2n2vvSRG28Oa1vuUweAaiQDImJb+qlNHdLK9
uzZz30ckQKRhrwT2brEszNDrS74O0D9MkpHy8+OgGC7hlNjddSSYT0x6Ku7A/agyzdZ8d8TOFyj/
Dcz1bS4W/YjUSghNAFq3xz5dHl8nNrKL75JY11+UreJ3V3UB7akS/qSCUy/UayD+ycm3iRnMvvcG
BrSA5fQNtkuvfoDCBEdvjgr+JNl0mWgxNdZEbbjI2wYudQ3nhjpe+FcwIW/j4++JGggHTDdb1f1k
zIozAiIeVIcN2GrlKbIgwLk03XrSbHzHgTPjRJBXp0XQ40BfGWxaiOk/NIxrpAakewh+SThBJ/bq
aBjTVgr+eiGAVkXcUBSnOQm778IzuNI0lMXi4a75XPZ2va/xfLm0jvPEJM/2NmfdoRYUG7XpGyHv
n6L89YV9PE22uIZwaWa9BqM7nSG0vW3oPbM8Vn7blPZqxO5GShZDZyFVcetKA+ft79FbI9uQwBqj
dWJhWyNJScyqc+X3UWczeJ4B7xAhg4CjPgTNGZ82/GS6L8Ie8ZhC0pcIMvzcOvLf/NodMli97XXe
QMWCjAZOpGLQqI0seZr0woQp3Pk06nit0l32URxS2K1+tBNIHNZfPABqzaDr5zV2wmF+6yPpZo2S
G28hAzRPlXoLAHUv/r5wZ1Z0ptYpkx9C9O2kJ85V0t5xwGSBgEfCNd4AXk020aIVpCLyTAo3Dhye
tiwRzOT6EoEdxpjKU0agq15KdCQAecQ8YDUf3EPsICj3Q4KrBKtu83Dubl8eFNLTGDIWJIGDI8hY
gGkx7BKw67n6xdQG5aWuahRyJCU0KyT0Tfbb4lJk743gvt/nFd22caUKEP1gF83BnmdyllFKnBdK
PX/jQF+4umdFSRADTeiJZZaBq+cXDlQJMB6BKlNux4K2xXawuGxBfgRVAVQencFEsb4V4EVkqm/U
PRf1DjWqMAzJ417UL6H0YLFeW7gDA02lIucob2p7hpKs/c4+imLxttwET96b3GrtHl+mVuGU8KQZ
5al8AlnasEy0vDy1u2//oh0UwC7aqJFEYMrK50OOnFY+Kj/RJFxLbWVQwXTlCVb60uRORQvNkvys
MqZKc4TX0NADmvbTY34Ogq+Uvl/Hl0oLfrlGehLPBdjXOOHupwUw7Kd9BoNU2Ol5netvEAEoqB4Z
QlHwZ7U56Pq33Rh0ZhHT/XftkyDS27ZdNXE4eca6r9qP52bijaISYCXG62v8OvhTcptpEgo+2YkU
5/GC1h9KEQz+TrbX3M3M46hZ7itjtkkS1LDKHLYGZLXFDTX2wtJ6P1zoSZTK6gCYFbH/lOu8Ppc4
Lxi+ok30yyAqT0DD0SoBvIBghucjX2TBgYpInTrQvhdYFyolbJKOoS7Fe8L8XJpaRbLJjFQ5sM6R
VBiGWPsMZEEYu7OCXjoBWxB/ZYvqIySN4mBDQZY2nlR9cyH7QDMMZQzB6uuUnYCQsXejgPBjIWOw
wJGBPi+GFcaWdIO01E1Q6PLevfY3Dp4gVTNZEtW70nOgGEOkDN4m082ZryI5aZ2MfUdLS1MBuC5B
Im26NAi6ka19QG+rs25fULvdAxBxB0wq3h7Mx1r2aTuKnrqHT2yBX0XUIFX1XdFG2RlX7FTOgrLY
wDCCpVwUFD3r7i7w5EucH973piz9rwhOZ0g+g2xRNyS54yeDB+FZRVrUSqdKDn55UqvRmpX96ijX
LzLbclSntbs0Uz8eeo9kPb3DQ2tUpmEQf0VsCrv854YEvpVeu/Y6lu3/7CCugvxDeR+B+EgYJHZm
pqm7eFvXIYeFd0d4mvpN1tO/TVJ8aMEFbQC/18kcveqlFy9ktfc52d53vsKZoBkShUweBlCNveH1
PWROoMlva+4lny6CpmjUm5rpeeWIllHWByi2JiDdkh9aJNmJTc8GApIaN8o8oqbhAY+HxK+vKhI3
lONYRyccc8Gi7/hn4I4fXRPX2eg+Brts9fqja0dw258jnzfiy1e8FpHcEQOFxvx38V51njmtCZPk
QRwQpo1d8zqUTdNyzZtIWgvdgoL6Uj987gAXo96ctqTlvZTS9wqajyDU6aqcIAnddHtwr+X5tIp8
kiNt/HHxMPTjwBGV3guWi8twwB2KJ+V+hloBYOpuUIpc2glBQmhY2OU2dHXlNk+obAXMwRIXboTM
hB6jd/EkVFG1mDueq38E02NcBplIie2NOjFJ4GBD4k48lle0MVcjTunuz72bSwjGexxhq2tMTFvz
RxDfk64NdPFFR2W2BmmpF5ym9kopz7C6DPbNCkqxSCgTdl9fFsETAk7Icur8l/bbnfCqdDUo6xAK
EyFzB+i29roHknHG352olTB2TR6xBbYO5IRTzHzdc1ccVZk0xgJhkifVzQ2bLkZFQgFZ1fyl7JCb
DifI7PQ3X3VaanToBDHur+GoVTQa8GCi1Fa4kIDhoVaBv6q2Gm7kGbv4pSSyc+PNmV6r1Idjv+NM
AKpHwdj8Uyai9DFZ+npg1oPdxcBO949r5dqOZsowhGU9S/Yj//mDQBfMvCZfZgn2p1WewVyI/arE
WNbko0Ut5aHcWUZX3F6sjgbfDWNHvbcBbdMIqWBtrFkDxdgF6o+R2tk7y/SjO4gHJDJ0NDN5i23v
rjl/AS9V82PqBUyM7dFjktk1AOaguHQfY7NhCWzdBcSrCMdtHI6QD+0ltWDBDm8xatn+mbZ2Rs57
8niUX/AY2LL11hxuYrRjZKKO2uQ1JCsr/cOgGbYL2Fsra8OrQi81B/9Jwbo5ficXmXaZF2BVzFv5
XRcWTn/mGzI625igR6/q42Y8O4cPjTCk+h6rkxJ3A7rix9RWseK9RnofQfzctrRYrrK2WhKSFa+B
nqikFJi6ELJZMP/Yq12/X/J9WWIOsqO4XwCYCRm506HsQ4BeyB2QQcr1ccco1+tMdwhk53mqF2GY
bIj8DByywUwbbcVzybj/IJpfyAD02t/JwCWRdW50z41hty1k/8D01YqSQw9YMaEkcGa1C43aiSCR
6C0Cl1tujAkuVlUMl+VERPemowqBppUhBP3hUX9+gTDVXT5XoOojXA+QvJ9L7uBVLhb75rOdyyiJ
qENmQyODNF8cPiIG9bwq6CBEE59Wcs9Zqz+Xg6gpl8lHPeZRakBqYioIXK1CLegwRzzglsPZUK0z
NOFYmUyzaYABKtMbOhBOklQuOLtto1E/0kpNfrIHYZu/ykDigezEnsMwMK+kbpB/iyNaxvNKw697
RBcweQCtzCmFzouXng7RC5DuiRL4DOMOqyWZNEM2f+yT4eN/OjLbPIFSxqnugAo2twT9K5GdePBp
NUVt5YpWGpjwQg/7rzT9cnsnzqUVYZ+Iu7l7X7P43Skuu0YvJbO6tm9xdJCitwL7/BMScjGY8j0m
BlRZ4Fj7KdpVy0psv6ppw+LFALkcqf5PJveyhS79FUUUrCOrQeabKl5xhC4gNmx9amhU374gokY1
2LUo67T9ZiOZK4es9O1X/3HhmuIqFMYMSKmoykmEKiJyq5tK3f5VcoUN5LRCWuje5/QVEiLkVWf2
2VRZC41ou/f0YS8UGvPSbOivCaBUS5pBCzQ9cyBG+aj6hB9o+ilkNgMWar0Qfx60UnDixDhCwh8e
vt3SlvcYPRWHayVa0GTFkAg40KvY1QPqgK+i/uA7LdaLMzxq2/x45n6sRwNSDwd+n4/00Qv8RJCr
foMtw2ZGZhZIkHyMDim31mavD5FjKdJRB6FvyMq6d4Kcvd58uMjo78KRiU68SfPg7EuVUvziqLjc
IdFRQ0+BXcuVt94Hfg8+GHiIetouMO4C6fISKXvueo9WOZlPg4FbUykEXdHNDgbn0v/aPefelUrb
nQajm9Mshe2kLuKLQw6F7UYirceVJ/Q62wsNwJX9lo4E+GXluPoppl3nEpiqgDCkzpaFDGTm1zCx
oFCxTWbPNvp42L+pYjuhYRaTXeeMkSAlWNgvJ96XyTU5ZfgTNKecVAiKdEYd7YeoreBGi/hNjadd
3igqYLBmBf4mgcopNQgu8aH4EBHuWnM4jlb00I2sWE+dL4da3J9UbMc2eIoyvea2lHO5iHMDL8yp
Xe713/V2S8FDqyZgSQUn2Iy/eBSV3a+wdDuoQAf12eATdLvNcOJPS3VU8KTXNcvEiz8dm0YttLXg
dA07TV07rXd2A57L33ecIGyV2U8b3CbqtNCLtE3Han04r/k3O6ojL96AqUNsiMY+J7Ilnq7hy2kY
NruV02eqTDhrq9bTYmw7+5WKvbS/iaJVoWTeoGjhStc7VVvVUFPkDHhmCiiCXfhhvopYO5qzeNYG
cQp8F0br9rfHiz2qmJn4PrzQ5yvila1jJaibXonbllhtTEM4pRCMPNNJlx5LhwXQDnOV6icJ4vbU
aOyRB808ObC6E/8qLhjaqT69X6INF6VTsnm1aouF8KXdT3TmKIbNeyMbHYT5fBKtX9q/+6Fbefx7
zL2Nn60itP+eO1w7FoGco4C2ajq5Mx8UjdqzzUB4oHaLeg49wLHNsdq7mesZ5qaCZWD6eUNqr4Gv
fjvXVtRalWGa5JzITZKxPlLWj65zgBJzaOIcvBXEzOF+R+cQhhq+ZevZGGrcZRf/EK78PmN1mdIL
NQVc0sBpVU1KY6PYwI0Aj7LwV9Z0+e/1qKkmdr/K3KaCxs6pbmWn6+7Zjtylw9KS4kRN69xRY3E6
lsFnp0LqVQQNvCob5TLdWLML88Vbwu60zneVbEjdfseHv1oIoGVZeSaRsDl3Xp0OA9S4hQ2Px+4t
vjLiOMMMolGdJD74O2ZpBoS/aDz92KHLHKtTsAYD22bDzSV5RpdH8RcD8e/xUYlpCsdacbM9iud2
sBQfNO6mnW2Ic4J0Zn0NrZgV/CbARSLMgt3zeVLf1kmYcM6k/dL8rKBSEWGVLv9n6xY8yAFL+E8N
ZJyKKHq9X2ShHPdbgZQhwk32Zyksffi3Lbiime3b6Z9Dpch7lZvWDZGA5sNbARY8Gq2FLyNdWRIY
WYJxe08knF4qLw9/hOyBK8c2q/pzGe9I2aPlNfhA10wLBxkHOL1UhIR/TwtnQolciiPzzXzBWHbl
kJon0sp1gzIVvYgoQwjuL7E4jG65J09lpoUp29AL0YIneZy0DBo6qE4lQ+qTG+ZTsB/PdL8tjmGG
AwcUfsHeKATco9smPVmrMbqMxLi8a1QKzwYWrW7YPiNNrwYS0Ivua8NJUbTVPeEd6CT7APD0kyM0
Ehdm5XPLQQisamgbShLfzF9UZd8Qt37S/e+MZnXmGKpyEU/x/snXHLSRouBAZijk7l5KbA1Bf+2C
kFbLDd6Anyo0pWRpHRw9g5vJ+enahzxLoMs8gQ2jM+b754VDJydDZyB0sEeCesdYnZd+QQCbQp47
pbYxQn3Y82MhP8Ry115XTFx8Tk3rRnsJXk18zG+yGwD0bt/9BbkkAUAitv+o8b4AL9sBBUkfptE3
xgq6jdHl5OzPZAi/hL1cZN88Y91OCbTExG3PJEyEe2JYXdWWh8pnEOK8m10Lij2nX7fO6lXFIOkE
ALHCj3MiQt9Yhol2p6kSu0hqVEstGe0omP0n15bMn9JsaqFEDuUcqrNIBeCFKg81AizFaN6ew+gg
VFCsGzRQuXtk8MSbSgYov5vIQnTFe1CYaWJuGt+GzammCsCDCGaxwKrnzZ+eQEMXMZthtZxv4YPd
5h82A/fXZh1IIirEjZi9Dy2JOQvgXu6EgislI+gXhbJzPsYIh6CGXX65HUjzCpqP9sp9eomQpyXZ
f0FlTMC1gBG76kpqHHzOmlfbweIUzbi4ezLxQigJUZHk0rMZxJHbseq//02im1qe1K/9JTsWok+E
GMdaY21hFU20Q4iHuG/7yRnEpTR5Wi/gvNKoP9+DN7l5myvMCI6MIr2CETfvGNmOkw3lIMZgBLBZ
MhNtlPKNhH4Job44/gUwwk1YGwZ5cIg8w1ds5aLFcAGEP/qsYNgxESHxkFBcZLXvPS0izgvZ+9Fs
/71tzpaa1qLzbEFJOvcHJwUaLSFcXpj8Nn9CYwADIdtVscOxqSDLXGlEjCVW/hDC+VJlx7QelfAn
CvRIG8NeIbi1weegAdiEpLrvkoZ8NTYr+fBINSBg8CoPTafn4Ec8IjRfK+c1KTF2OlG6WwA0kYcT
24KVKd9OPiaXRLZFmGPvvq5+yXbnFQD5wF0pUYWuRshwQORFeakx570pdnXXA/KiSAaggB2Yr1dh
DImyELz2MninmGpAmFOzoGwioeo9OKB6YwjvEbYfdngrGqjFTxdYOqm6GS5+XWudICY1fmkILs32
T2kCNAPM9CzU1r3KHD6arl1WYPcOZrxQQfPN+pJujSDWxH9ysV1VbzM7IshuYZZ9g0Vglko/7B/L
pJWmZoywTMEbLBXJdWWD7LvEMMahT/hOmMimu7ShCy9/vsMzoUIqBgFNxd/LwvMBfxpu+/7t12S5
7XullXbewX8tsd0vbWXr+YCitDejZgBM9nLBNUWuwSlNVmeb6XBo69Wk6vddsnUJ/qG9XO7OKS1p
u4UH1TujfcZQlVlUH562fYizM0CIO5707psMMy+SNNFAJf/f9yqQ397uNyEkCPL12tagWcpPr4Mx
zzZV54e86NTh9gcB+vcw6TWGgxA+R7mvaPGfXRC470aiPhKHjoeyMavyqCvpVSiX6UoyQ9MzOKWT
PZnxKZTdpfiQum5LzGsCMgezeArE0c70aaxMCGzh/Kim9ewTZ4at2FvYdoRQu9104+Y7d9KpV/VF
4VvG472+UBU7XcOkD4l2OBV+xPV9L2Z9Jcu9eooy5OLlr6LQIaLQvsKnCYIpAJulJBt7ZgIrY3J/
jM0/o8OOjFIO3sNtw06hgjkorH6qh2+OZ7LCxy/Oq3QCX2CcI9H1TWrYyNXqE38D0ea+jrngjl1K
QavQ99G6eG0PBHHL3m5OOJKuYIoyFOjdMA0PYOgU2+8UmOr11nqTpTZ9r2toT8SDDKe13mN8wVtq
ulibZvYQs6f+TvWjtoS58T49fgGwVi+uxvws8ret0t71mUSFh9mvBJ8c24Y+UMY4iokEjP1joJfC
EDeICfaWqVzzA+hqKDGKFv+w6/ZZVeKTsBFSv2DXbw1BW6d/P2kb9YIAk59dj95vr65ZxGYHv+3s
RXa5YdQ6LmpAhsD0j3zyq5PlORklcetKfs9AasTgXFGnfLoBkSdfuWS/eMEsgTCy39YeSFMW0LCW
lYtDE+xgRrPmRf3JADx/5VMmS/o4TZ8GKCtDZKweKA3B07H5X7B29AG3oD0No6V0nqTWdKnd6ItI
Upobvtfm+1cv6+/y9uFoTJiYpXX2xeRZ8x1ng+fTloEgcfEx1ad2IiaqwqMUEhqI3xX8d+gk9N4K
s4S7Q/Uo33YH12zcy8YldadMDf4pTXG3QCaDGXUQmYkgBhGYXKZ4m1q0pxfIaLNq+DPq6nxgqgHQ
6see+oMcqqa3CZwJmENvRptOf+DUNq4L5kSErUg6qrXhwauOKiIBIhT0qDOWbZ8cuRo4zPrPkR61
OXoAFA9x2pWR188TpUnyRnnqSJrh+53rXNPx9kEBKVW1RtCN3E2vhE/cS4NInaaIT3kBOfHnRiC9
vq8Zq2DTE4XXdsfimtsCdQDwr5ALrlUYeyx6EJTFhAGLeP0ewmNh1Ay4Or59AEftnKEpv3g8Enh8
rEIRD5TUl+uxXqNp6/I/Fiu6q2aEnKuJry3qEy+puoCyrYhf96r8UJ+N3o+8t51loIPQ4jF+fAgF
J5D+4aopxPAM1wWpDQjySBnJtqMDIg55a4x9P0YlGB8/6Es6cwY2IaYv9Zun4OlXbNnq8od4vQGp
UBPpC1qo28JhYYdGiZJLbgqWceSqcY+uIn2LROfVt6Nd26cPJ4kN9VdzkYDDGCpi6q0daoFnr5Pk
yRkqsyJE7Waf7cfcVJjXbGR4YDSo9PdlQuoyxeABCCoe2TSDK3jg6gorKU9g7CmeLAX4217g1LXC
vpY3y8PqvGulwtE0HOtZ/vPbtkX/B73cwKHVMZ+kruafX2T5Aipj/uA7C7zZ1YesttSfH2eydkxz
KtENn4d60cMv61B5xn5UQ6I6tRqJWrZrAq2A78tRfr5mOrrnneLYU+zBhkQ9CC/NMeM4gswQeQLu
mGKzeYUJdVNmlxlbWYYhNGrkRAt1P0oN66Zs0ccIoWTANTdnhsf+ogPftHfeokxjsCA2BZ+Z/cKy
/bxBGvW4CPF+MR8o9X52cf1518Q/5yb8C7pau1Tk9sZhnVPAbrrYRGQqGjRnLnOVuvZ6rlkZlEwZ
KK0ZpEyRXkwotxFHSgGwxY8AxPZ66DvZdqynIUd0ZGd3l/JjzILTNEKtg199u2udpOKZnljt+JRx
4+U6PvYj4fPGvY0I0501AitJIsuAcOLyGp4sW6HVsDxPMtr5BXE60wu2A3uzDDAmeeP+fVDyD3rX
0KEtUMWisG27S2/1J252nGjIOmJriUTke3DYCMi32s+nzPa4alj/NHM9poW7Y2qxG6/R1BkEM45u
2owM1xcUgMU6W9kvJdQDHoCj3A7HYoy2Qgnv6mMyLWtIEvSQvsPBOOJ6eau4ladk56f4hDE+ZIcb
1ycD1SvOJjmm+ZnmOTa4KBmwxMo1c9YO95tWCvqQAN5XAvkkwK6C2JsQYQhCIqel5iPDDCPWU4V5
TGt9d+DcSSiwxJlcXKjpt6MfV5UB5EbUOJnh61b/IAuM0LWXMWen+hntqLuGHE/TKEt3Spu6z6zg
dkt7USlhjRD5kCcEydsya3wwNWyTu0IjbdpS78ZBWVblkstTcmYFIn3j+nEf65yHPpVKsmtkUBQ7
XVMC2kZJiBn6ZZ/l4+K65pNz98deQghH6FVZonjTzhQigU+Gy+IQ9usySpCnXQQTwljccrebCRA2
bShgQh3dcaWmFuxZ2Y2pqRw9TXDe2xMEB6oWa4r+uJNWPGZVjrYERg1GSTCO3SoVKtzwTyWd6NIN
R1NDHi3WTAUh/BlJCQR10YX9rLuJp9uraprEmSHn+O8hOSUVhI9JtJjui6uRxH6IIRV95/1s1ur1
YyCsOFK9MBDKLxMSiXJ61i6wW4YOq9Zs9rJtB+cuU8YVxlFbSgt9uhfEtRdea0+aV+Iy/H6Qylii
yn8AW2hfovebXkHJNboTTRtIqZJut71vhO2UQAKLNncRK1JT4QmXK7+2UyHCMyyXAgAbjzsHwMnP
xY7MGzH+m5Y0++v+sHZC4Twe1aj7T0iJr9WtaObQcyLgUaSXiGHDBo0Ab6mmBuuzEdviK7XALhlU
agfu97IdhtCbeO+QKgZAkIqaUFgjwltgUz3p6yL0O2xuLCeP3zp+8OGMFRRGmSLnnebvsA3jgAZX
7SmW64lCuzHiWXBcTYD9T9Z/TigNQaeA9h8sbv8OQK0IpPA2NQv6bYuNGrMf01HUopoWlgOzCqTY
HrrGmUusy29pS6LoC3abY8PEZpbfspUQHPPZ6XXGovKKJ5JzHWbm6OVQ2Qt+CC1Z23qD2AyGkXOE
psFQh0D3NaWatpJCXVGVvz9+2xy6D90We5j/LMIKcVA4kx6CkvLo7yRvcTCGYkJVpIDam034gH3I
GI+nTINgp0Lt5hkPfjiYiGszO4LT92bNFge1TCh46EAKuQ5hnayAD6vNVZ4JZLF+hFlJ++a3Q1yC
Q05vf7mP7uKoxWtI9ZSvvJi9Rf2Ux/lL4csdZGAomlNmnMdYmyvaDrOeM1Iz00u5N/zjMWVVKEAG
ybdxqTuElAptUzVbjc6pFA1xcwdUA0DlJgoSKYQO5V++HoH14Vdy708efV3JoROAi3xb+Tw9Fvk4
W9Xve+my49cE7e9bcB+hQx6I0O7Jzx+2/hsvN3bF56o7/fsaPVirB6SOS+sYS+Srts8LFVFpM4SU
d8bioJ2SkBqVHRLoRSee+5G8W6kU7+4GQ1oJtZ5uOJ75no/v984n3u1yrZM8Zzs5eiWPJPQukpQL
hOtNtZ5skUMcjWvsb1PosLEcAzFbbIHJ2dOYQJ51Bij/zHZIfY0Kyu7yaGkzpANk/CQBbZDrO74m
Bbj8mkUpjg2CTwqNiCzJUO2Ndxwp+zdI0sSgzbFtm56637wQYriTqx3J3dkQh5NaZk1YTCaNRUdp
MGmUr25htpTRdXFGJ1B/84+mgOKSsC9jB76hOaqAbotoJsuCJUdqHx8SzmuNrF7Bi95tTkdtefGt
jyWPRnShKkNpXPhMuu2ryWtwqQUeanLrdiZHbchC6xqR7A8d9g4H0cbLApPEuBBWGVd6ErL2pszo
TObZ/cqKdGfCpnIk+29aQy6HaFUt9xs2ISboh1cmaHyTAiLscM07xjR1Epwy/TlhV+5Jk0hf9WLq
hXgp/NpEaiAe9jRFyWfVqGguWK2nUaaYV12CnRtcJ7QLPIKYvZK9EGwURavGqeGbQx4TJAsGRHhN
ol1xyupAtsoSzKeYCiGj09KKx28WTAXPgMJ6ZwYf8ZxVwjCbtn70EqEhiNLxZ/QPM5g3k30tAUxT
JwIpO9bAPfULDkgzflLicBOYTl+ilspnij58469PFFY1za4MSl6OqcsiCVjq4c8dDao2VrfUfAsD
URavz434NNpEToaB1sQKs6TQqIelfW2jx91yAqZDA1GIs17JSZYPGMZ6DOBd0RHRw/QZFGQl3MoX
mByrrS3WfDkXBSQafwfpfysp/m1+CwMeG5GO4bJjQcjTSnpOwVd2uwOJz8ti5Zr20yBKZ5VqVbCa
zruGZi9dcVv7tEgSSOjHeUIwNmAVbS9Mv+PODL2a3MYlFwsumD+5CcxblPgxKN5jyoOAthDJaMoU
dQQZPWxQxjFKz9lhER7fKr7qtmrrhMIGFFfYyGWhfC+XeN4z7RRhFGS4yxIMgqsC74f0daX678Mc
br+9IKpvTgU5KNeHM/btQgTQ0wFgkD3XvEPLA46wN5n6+L7SEgvyJqkB/88TWQRZqDx8Y1tQpCRr
Hu/89Gwab+nIBLRecKF2rur64LTvEX//sWhe3cWOajHbWH7YAE65o2OKYWT4ncWh0QXHYXBOlc+S
WpLUqB/Pb2Uv9KiB2+LdfQXk7UwFtyQnh04eH34eLMjV0OsXIKf6q7+7Cefm87JWf7rHlMM0TOpO
QwxfRa830PNokkUOaWALCTm+Mh4hsRHHH0bQkqVY6UFJA2j2zkIDjJHNbzCRxuuCNX73gkK3czWy
3aX10Dvt0GwBIdAznBFTih6k0eYh5jIKol4AcbBUB/UEWAU4B6q+YNWh5Wfd56TmD3PnwiiHOS3u
MOCdBRqF8ZDbWOnH3j8UIyjvubaaEYkbZEaSlRE0I5efFMHu7jM/WkretmbqsxMV8ym2fa7Fy2SS
N/rmae+L8RzWIcF/JIP7vVsIIMYdM/dY0zV6kaLdmWYDTM0z67Vh7bufXEByKP69FxCborTynszo
Y1z2zz1YFvqpTTliVHdcb7Fz8y28GPjagQVjRR5OAb+EU5pAsBHSdMky5IMRJWvD4EeNXAEkfgx/
gLLpL/T3woQP7CMHqopUClU7aNlmy1EO4GAWwje1wUzzvrt5FFXb6oDKv3kdzjYaX47D1e1rxR8D
WSlXkNQ7zi8leyPcl6snFdDJV7NXeNBnlCrD76LSWjrTm+6Ql+wGc+Z3+hLs5GTA7hblWoffCHMu
f7jUSfP7Un4rhGvwOKGqupZtliSRoY9xjez5vIsmUpzJndlU+WQeFNSuYRLluPLaWWt5J9YDUfsG
M9gns1cDKQdQpA+jgAPfwmM098sB3gya1cU76dxd+5CdcVgLzzgixtiR2wPUpxaKWo3jQcAXMn9k
os/zqBxL+uTrj2MLiSmXkUq456A7+JGAc3+8JBFvGyo8qgzB4OoL5h9TMbZbymNm+YG+o5qhjstf
yclRgdLROs8gyn6Xpj9Pv6WE0+UkJN7Ct7pDhisSyyCoLgXmdT1VLq7bXntmd2yX+AnZ+7ZCGwiw
5a05tV07XVjsusSeq4zG2kEfN8JNtzdrsT9Rajdcv7MnKiAn12sPP5ckduF027i985TH+bQ8b90E
GQtTtqnTQ/bzFXIiCv7DanUE1iajNdREyXKfl8ONXQmPVlub5/0F1tpXEx9nC17T24b/2ToeILJn
gPZeb3f5Y3I9WhNttuFWWuuvQgkqj9/S0Tv7mJuW7ORjltvIegqfQYM63o0zF8w2rFMb8OVNuLDP
CNN3OjqbhkVaXmUfE1dY0xG027Xiz6Lk97Fi2FrDO9MGrHnkRlrMw7DFTJyqohYFPXunE+CpL5wZ
tt/iKe0LYpXiBR9qObqNwz3hZp9JZZWPQ4j9LDIB9RbjCB1OkuypyhgteYCZneqFyN34cNDAseA5
EuMgoczmzhogwDcXaHGZT/Uu1ml1A+yodg3npPmqtskBcyudZmCc3wnk/JB1Oj/SnMJuZj64/63a
rxfL/nITVmpGJP9rOjUtssadkEkYQcn64OOpHhT8+WGGnBZzcPWrNF/EPglPMjcLOSFXF9tp8tux
f1aVvkpKec5N5rkf6Buma6Pz3miIOYWW1oqoR9jfmrmPQdHfKPIekZ90dbzXy1MPta6LMrn/PQ7Y
jqWmViFdQHPnee0G08O36VLYI1FQLZjNmhsAS4aqKuRyeY8oR0HrrPBG0rFv/HRPzTKIEi0uOqz9
dvFUHfq/zYavTs3CtWNnxIIVQFWcDVYuW8oaqp3jPSUwgzq+e0b1kNzxpJ2j8oGEZBoVMa2/INo3
Md7Bu0G3QoSKdyM6+JUOVpgtUPw43aBC7I5tqJECAvcFTOZnh/Q0E5FxBqrc2rOMahUWtutBz0Qm
VsLgOmMXE6HPBhP6bAgrsJVz/dHHNXymZSrhcwgM0rWHjOu+PEYPuQZIVfpQLpKGZwbl/Ak0s/NN
TEkC80QeslKT3yteIbSOL57ixoZn/2zdFLon2MOiIPhwY8OAyIF4G0z/hdnIz4FjjFbH46XKEJmA
mTyF7Sen8rNCTfbZVIx0TI2xDtZmazwuiQFWQM/nQPc9fLojZaSAmfnT7mT2fTiSu5rT9WI1ruX9
QKlrMh1pi4RJ8GG8A7IzmekMhVwHnZeO5mutXRoaLJJNOf5lYyVx/nNCU2bATNFeOPwdLkQ4BwxP
r1T+Q7lKoWZiUxaOsx8FRmarAgDIuX5S/D6o1gHh8K7Ea03mxlJ5sQJx2YPqTPN6Gwql4alCKykw
DhLEUTC/vRywHo43pZHNnqro9LpVTteh1gU9W6iQ0O+KqIGKwK67JDK5iyeTJG4cb7yMmfj9JxmL
ZnYJWFczbPktpfJxcYPOQHpSbEQqejTtRy1RBVPa7fBTEk3tjw+6aUG2yLpqKSZBZmBFEBvgSUyJ
l9ZOuynhPmlkEiY6TQkKxM7l1mTcGKryzE93S3m+UMYybLWTBAOQ0fx5GTz2r2//bugDSjN5SYIX
MFuf6exjy6vlzwMdTo8MP6nkenwWCN3RZ0ic4JNfaP40shdA8bvubQDfMxfsp7GU4abQzEhcfTd2
ENjJWpdRJ/WkfgIaW26IAn1rkG3A+Kqs8b8/Tp6Qnsg9tJ4P1pVXjnYB+ORqZBTkrZn4ANFluyMB
6Kh1jdyPcf2UAJntB6UMbEVbk7SUsIp7uzaLNXNh+HdioynF7qfokGb6YauO7zVmh75n1H5U5hYh
k0PbcR+20IRnM5hkdcr9cQ0cJYxaSwelYjEw8t7CfVZ/PhbqGGxFWrMGiBVCPrYzKKmknx+n0nb7
R/bOIBHn3dwBsGI00nnrQTXUfJRMfyv+2jU3SRNdJisyzq1cOr0/O6uYvyOPfmlhAze9I6YesYIq
1P9f2Qt4Pnxo/HYuDkp0UDiD5OSZqSuPlKnS95U/kJXpZspSp1Iv1RRDgqoe+WUmtNZYuMqCwBmU
MVDRkneTqv4E7e4CIeuOnoLO0Cg8PhoaFGUo0GhEA0m/9dd0VEtnpMnIMmwzuQxEoWkIaAFwbf5O
7SsAFR6k7s1n6U+vgVF/EZN3ndWzDyS+tmfjOdwIlX7OLxYBtCmcf0EpSVpgFouFjpogW0O0Ux3J
n762FfYRFQUi+DG9AJA7Y6VehnsU/fJuBEMUjqeIsyGBCS2rOFhflEwEWcTdiag5jalj19koaXLm
xzHp8GMEWNkfHbl56vGVb/OD+ZAdUoKwcmeihQgzDBwzoP0X3LJ+gI1kEh0tKK3N9OOxI++Iadfi
wr6oQvn45B/Dnsw+o0W/MfAt+CArQcm91ILN9W0ARI2wkRuh9xE+ONq4ARzKI9WgpgxwO/ssWjQT
+HElRVUM81k117Zt7LICrIfXwqj99V7I4Wwdn6i+f4fKK0D20E7gcT20NYvcBCHL4yMTZzjuy4OX
LyfK0TQWivSr/+59sRhjOVrAiLQwTgeamWwQ5P0mpufuFopxAr+Sk7vAOc1JoSQx9blD6llsPk1D
idIq/0qFs2wSKb+QB2nJ7IaE74OKy/Utk4VtM9ulcefNLXgHhn3g6uIE/EyNLFKS1zUsIbAmXDSK
1et2KPzDITDb7GO2SUQ8Wgf6Nl+cOB/rogs5y+Oj4jv1Hj+GorzpPNceF0ilGReUpd2uZCS30aiG
uESSNv6l8o7FZJJFaL9zGga/dUVQK1MEAf1bkTGXqpVn3GYCjAr/Q244Ardm7sf/PjeRSgx4DGYB
70jZ3bzsQo1t8GG5FQuHh3nd2451nYPgBrl3o2aQOUc97Ya+CLuvzeh092k6NBErLTD5vhEVFngG
KISISVxpgSEIoU9vA1v5rqP75U8RCpuZr+m0efXVTcx0jl9vZULwXs9RZBwSw6pV8+WATC3ikYRw
UeNZwaKggRlG2aKNPWEpli+ZkKzcIXJiTQKH0YSJZxBKTb3vspgyRuXaB8vthWTpAzsikkfK3eZX
y6683eLSSFz8taSIeYQ/adjVJa4R9ZowNUAesoQOM1KVziPoVyitpNNWMVC/fEm1Ddbq+n6T6fuy
6piMac5lEZS2ZUoaiRcavl0PrBeWBVbRU0seiejw2nskDZv+lLvPt6QbVLCSwb8T9M3QAia1uFV1
RX5rZqxdAr7skmCSUCAyqZVNR5ewDj9wSt+KWEMBSWjFFlcGFgq3HoOPCoETcfysUUVDNe7y4Ocq
Om9zvV0Dobi0IJIpeeZ8E1ymKN19JWXzicanmKlxi2GNyLiqFL/oFD5FDKKM+UtCl04mqcNmdhva
oaElO4bwFKFIjmtYGvkdGTwT64p5hDcqbmGHwAJAZVUvNlX4oKMkoro3gay0WBwZN/F7PF0qKKyD
/22GrL9TG1TqXEcn1wVi+8pt8vvMxZZ1I1HvWCzu+FyU9ClgrWq1qhgDrHYPwXujvehtZhvx0PAQ
ijygnkn2nMg9dr6xL9GzZ9LNHgNiHIzt85atRqQirAbZgccJWP0wrGmIUzPul6Gjg4XXPvxsPbSi
ndYkCrHFPPvula6beF0fse3poZZI/Wmj4xMPHwOlrQXbtNlVdf5RBHIZ6ummZ2dyJFcrbilk4A9R
D0JDUafCevDjKZ74mps9S4HnBYirFPPcDyWHAswXl405j3E9v6VE5dQEjXvjpjnz3TEYgzMgPyR6
yTH2pqdi87vtg/FdcttWWHkGlZv5AT+jgj37rD4+FLCt6k9XG8n4r2o5PpGwJQn0KeNIkH4IScBp
EtdJKixDOQFKgnxnYWry6/iZCn26XyFmtICRcCr2oKdtOyeiEgki6HrRq5m9PMff1ztgg9JAOKWW
WNHt3ZbPOvM2cPR3kErQsfE8qrB+PV197xgUAmWAdLJdAuEiLpQMAsk6T8vhJ71T2Lw8HDhA+F5h
dJwkR3DeO8JyarfqDLMXzBh3jvBkoV3/Lksk9tUXUujZ5gplHfRaIdcEwWz0tW/YSHYTSqiewbjz
t61OYxrWzYqbAIwt4NPmOdJiDNhFakaeery/12zye9jJV8qWB8rJ7bkwqMnz7ltY9fuBeTS+DdNM
u0JqmbpMF1a8F+DYcYS8TQmgrvPW2Tpn/4pGnTwGzRq9YAWGgFgly+cdmwK5dfuBO+3WytvUMcxP
FxGsDfiwk9nczWsTuFH8rqWYJJyP/m7nqST1SwA1dYRPgvBLPjLd2ICCZE3herL3JPyQ/5XODyDo
Fgf87m9mdHmCRcs4AawaJiZ5aKm4Hl/bXgCCWDEx9rhQrf0pJNzPori7aqgb38xtF/pOMcbiy4BB
4QQjX1qqtVVZJpnZeeBGYS+xjHipo2DcYZx/2WIYUfxraplGZUjoUiIeuGEhrrTBneIjxK8gLdJr
vOXUBnzWcexSl7+F6SPLHKd+oBwOwpaatpHyiVjeeWzr9bLSfD2Eu7BsTaENyUirBZIWrF3yLd0L
5g0icV15dH+iynNaoMmv54sMUR/lwQjwOQ4/gr5bhgYuECxSsSz8WisfFKpX3ZvdJkaxnYMhgweY
BkbAsbrWsyjPXabtryP9E88MwLY6fbwFpniN7iCOGLbIVhtD66WG9SKzp+NzMtakqCac12qA0WD6
8L/MpCy0G1bPSRefcMohetPjK+BUJO6zuccR7uPaNb+Vzk0Snib4BWtZ9lD/u1VMbC9Na1tkWL6k
4/6bm02ok1uNWsdHTiM4hu+379WxJ7vsC6feC9Cfc+Noa42h781LyBqWi1kyPI6dr1hZwg+Lb2dU
5CgthHnY42xsg2A02pzI2Qhvk7EJigj9/vN/kAtVVuxBlFehpzdN6GaNpE5yoJx31nWLpsm+V75s
U3boTaMLZTXA6MPNzxTM1lkQVPBWIf+0rNBfAGQSPBywenKzODpBwe8JQyCmnZ39sGQtMZu19xsC
EWAWelQk24QgKCN8yXG1t3UMmSLHZLIv7T3wcTem/6Br1GY6mmq8xfESW5GfQxMIYr9CueUzxTwK
KsWfPJ1eLS6YPdyfIWCSlBc50lfQJbv343F5CLkaQA+j6Ta6sCflX/EbBVlPkhpqU6DjLb8wM1nm
KlofLFm6o6Ft7ZtbvUgFJ6s6mF84vsCgCFd2NVxydlB9j9N+tGXnPL90DGchTycazf8zesupTpSP
bs+rAHZ8cykSqdwyIpc3g77xoMeva+LH3OmN9ZcnH7+BX5Q7L1OdfilYXU/CYqAxSBK9USURmIb7
l1/S0x0RROUAdD/O9QrZoMVg11W720+TvREWuO0Nn/Zdy9ko3devD6SgL0fwHm5+BuCklWwJT4r6
FRh8JeompMQGLpnn24UBoXOHpHw2sSwgyWcLvoaqhrFyvvSt6fSWMG8tcSZhGOvm8GJE9tVUjGZw
Kih5tWjxHBb0uXvxPqBURMz+/92nYar42GKpM5cSa03qilOaI8+x2WeBks5bbPjtyzRswNNuqhjR
9nm/5KrJpWyZLPhBsVCvzQA6ivbTbO22LraH1e4qAxQJcM2ivrGbrxEBC1BqYeKqIcpUFuYckgCG
eugWE//BhKVooifR9cEV4nRs5hNjFZIeYpFvLxTcj8G3VBgrhoVL94zyW4lX0fUiEeqCjj9zPYV0
lgpzCVbjTL6926bglvoa7FyJ4U0lrzkuU3JTfCs3+chWo7Mv+fy8RdyYro8UUmO9Vo7tqj4hQMqq
AaxV/ra10zMtZGfnBXa0qcK3Z0cqpd9tC6zr1t+X1MolrND7HxGLp9h4us0WY4t/3zzgBsafJIJ0
ySQ4VfMcdiqDvXg/yJkCp4x9actaqWeWKBYYByP5dZ5cjpN6TyrFIrgO/dwo7GH5Ntacig5fMN/F
oCM2y/U1InEpucsJBhLnSsqWNB5D7scGbnyWi4lpapGqX4ZEUtOhEPx9CmCkO4qIO9LuPyyCjeno
lB/YXND7MTneJkKI30F1ZGF9sz76gIFk2vD3bwb/eEmgtTwrjYlW5kIdBrJNDjAoo6d4nHsK5A0b
iNcnc//cY/IfagHC8YSi+rNYlqDQgDH9Jgm+NC+CF+6EloTnwuON5x6hV1Ca5HuRJUdCjJL6KfZG
ciJ/AEAUOM9583h5jSFXJKpbqqb3olgbbijg2VbNTY/h+zxwtTO9+c8aAAiGkNxFI20/Pnup0t/6
0HJgo/IpTCFnjHssfV8ArsalFt04lC1Ly/WWDjUy7V/vcMmbcW4ffZTsGbw7Df/ik1eyQKsUX/TM
uTXkzOMA/fDoZzwQ/dc/SODkADobWHTMahw46c2jKX1r+emU8boy68yn9HBsDMdky2+MxxR+hErJ
d+kGJJM7n2LvwdcNVJS6GFRuFMUU/2XK+nOuxt9mx2GwXNitZdmCQtf+uTwSEq3zvXaYJp0A4qmw
2byKCYfhQtnMLvzT4pDXDnYL00GVWCu+xCnuksT/we7CjRusOl04S7TOauZhy7orIkdSWQj3DyUe
zs6SGUrtThaGdta2mq+BPlqFAgjqupRp38q4Ks9VKKNDo6u+ttwPeLUDFiUxMUuGEIcdTUB+AfKp
6Cf/0ptE1U7hClGqBlMjPwtvMS87y3vh6CG31OrYgo+S3tBdhCGenprjo1H9O8Mz2c8UxRcHk+8l
5edK741xCvzLL8x7x5MZYw27qxR/8LnCQFKZzdhMsWHYAVELlURzqvkI8vqdeVtJj/ink6CL95lT
goam/OcdfZHhDfS6ktnVHS1D3d5//vOgBta14VR1O73vORYx1tjY73r1UbsP+0EgavRlWF4cJpx0
+/zZhRl/J7xdCO2Dc/1h8IiqsxkLIvGFODPRto0bUIFA28qaNaMm4F/JYlEKftvEQ0FyM1QqO94z
3LuewJDvQFKkv7y46fZoKHEw+uV9HVaOTwqiV2fj544RUplBl/IJ6GryhkuWa7ADhxXLy1p0bFUm
Gj5BizS9DA56XkCTOdbpM/3fuw6DbXk5w1sK6l+k76nykfdnoIT0QFvwhpDtZeaG/AT7rrZeK6my
L+yG9KrGEs+BsJSItUeDkPVMZexJj2ueMCW2I79U75Y5yrxG2DGqBBHCCRXw7oEi97WeG1r2jfwk
hEEli9dRe0ve/1u27OXobfisxhx81nANJ1odOegfncP1FeLEhJaCbi8kFnE6O7FsrQtaQM00eXNu
2SjKRfXUPqpPwSyBKC+v07UvhW9HiklfphyhLbuAnwFUN7ms1qENYlfGCCphb8k6j2l/KL7SrELC
dzlQfdPaJZdwcRAvYQPdVZhR5BAhIVWoc37LLMgKbgX6TI8tFiBLTI9J//PBub/DhsLToqcHZAhq
ggEVRsqcBSxwiHFruh6UL4VE8QD3TUAg7JGPJiPJ5ETGTBvyfIAfItl4QvPeLSqX80WRnyrkEI85
8pnFpRrVjq4M0XONOszBXuNdPbXpHSJO0HIqfS9qn2MNb5WEYYyTf+6K4SQ6QUXjiJB/zamIhGR9
Xkw5xzlRQ3BN8U49pL70M0UGPAQv6LPbszsN9KxE+ULm6pP8Q+CjX41qDERWgCPHvEv3iU740a32
2Pl0c3v8Yi6ZEs7UeCaYUWRGx8cfwQZ3UE9DgqnLW+iGKCoeACqAkVIz1d0raqeYz+XYPJf3XVMW
wedOhHLOMu4JtxZEcbnN6jviQTwTwtNtmulMv0oxKdg/wmGgQPBlIfjqOb8I96CSwXEU15csXlkQ
o32KfpPtgfK2f30UNYu3h2jDz9o4BnhMkpHPLC4rtbX7G7EjnLavOg0VxjMDAFt5jNqTMOqXFHfq
uB+EKhL7at/Z1D02CROTIWrUq9q5twO4AMT/9f5bbwTqdfvLk0pXzbKnHBNO7BSHAwa09hFr6Tmm
Eg907F7WOwlZn9YImwNUd/XpuY5YvNV0m0rb8qxHYhl4jNdxClYdTrHJ/212OJxC5Gb/q2SlhrSj
qPYJV7pjADLIKbvwl+Qew7xcFs2Me06wjIMNhPMxLrJSGZDLvoNi8YyvFk/vc2tGNduTS6A/ihEm
/QdXtR+CC8DkI1jd4jdZaQGtn6qTGuLdWdPpfLrVHOlXnzmV4pT4cL7Vhqnan/zLXxn2dD7iX+Q3
QxtMTZEGrFK3UPS7QjF47soy/ZvPdRrd1G4Fa7JrVuJisXQUhAq1HoNwKFI/gURW9bLI0oqyb+3l
lNJgDhO7Ad47XeWBRof5n+lv8+PEhuYLr6c7dXeWNiNTU0tjLhiXzgliEo7+sGHlRKQzVaO5dzsc
dl9y2KSFolUx7teu0vQUwbqeCzKRYY38l1xPNcgITdqqBjy3XRpx6Sy48r/ngmxef9jYb5uPbiHn
Wk2BTkNJ6Dn6hwQzTeV7zPlM1iexxv405bUQdt54K/TydiXMqX/sujXxpodUPCAjp3FYikluHKmq
DtkV1Y0tZG1KH/n7U9qO6LkqptPDup3t6rFLTV870pi+WJcp7Lbs6m74G2pXr955bSFhcgrMe/P1
OcBxFZLMBJDp4wG76hq1gitaXjnUWW0d+uR5PxoWlbf11IswfynfQ/4z1ccl5Qv01PIv0BTMgO97
KK4fooSurwxl9jL50Fp8xJ5rpqUczjdvVwivtHJ4bLPnn78RSPZEGuoMekpVqziokuGg2Pi16t5P
8Y8Of/hZa12EXgKtpCvdiaTv11SMOPE2ufoiIGX0HIb5RGAMKmPVd3vkvTxSoqOsPBiBROUFOV0y
Mx/yeCxAu1QmPAQakTrrKpsIFoaD5nWXwHEhpAodL3z+lV/B1s0KQI+ywik2EJ56Q/Ln7pfh3/3b
PrlZJan2MPzxBN2s+7M8eR2aCVN0XpwQEHpnATpO2DlZvX3XrvoQ2IOYgg0lt4yZMTUqN0/WYTKg
mymcWgIQuoPZV5gTMI2Y9ghBXf5IbaHdqMAsuTfwFz1bhRimtn4lwcPYFc05X2KX6iG7w9tMYXqs
WlVZMdD6/uZOvf4yNiAg3AdXr+DjntUzp4m+8wmAtlo6HvvlfeOyKb4/sM4zkbCG9CnLaEJiHpfK
mSLkUab8ewGg5nUyfowVwN6reRYEvUs6WuRBM+K1C/7zhhrQQN1L9dT4F6nupIMPJhUW++4eSuKk
4gnk4knC5dzT54KsmQQi/5iTwcXcvwfNRgb2lCR9RdkNFI7D8PGVOv/xDpjIfXYkX9jiDlcwDJxJ
3Zt/qUOeSKrh6Y5OSaCjoCIGzZK3OFbTrZzq2Bt1wyCBW1l2Yd+HoWGkeUSLDEOCs03v0hjz2cnI
9r5WlgyaV9lpD4+fYDsU3+oK0ckDmL+04oRJN9hPaCZiQeBO1Fa9CzXLPTRwXylycJ++bnkTBtbA
p69sFfOVzHgEryN0dmFn0QCu+IDVnZeNhx77A6+11zQ/5CLGQl6PDzJ4WzQaogmWr+Kuwi5sMJlm
sXV1tYSS/5UCRN/pDsxhS/87GWI3FrlmaBh144aG1psbDvxzzkmx3vAmc5xNYZ+DwzcTNNN/czxL
50VSX8kwXbCc8r01AD8OxNxZeodxHv2xL46rDI77nK1w2Fb6LmDrJOhUP4yIaoy+w++UBGHCFQhK
mOYoS3kCRXwtAxA/AOc82e88SlRevrx4KMG/0GPLYwVQfFFGf2g04dJsBD0azmznmADrytC/iOO2
BAwf+RciC5EXrZ1DkJUsgj0Yl948fcznZd1LztEKgLWY2PyzShGNmYVGfPPpMtOn06zkeRtwqyYk
14rtMtZPnJTON12Oe9SvvWR5JkDpgjM1ROQAnne/CV0yZ7vFmGAjRBIU9tZuyS68r2DXlB3/yiaP
17W4SNLbbzuTWoGO908bHOHRzWfVJiYHSqm/AKkTYbD01Vhgert2CxJ70NNgarNEcokrB/8T5+29
rLqERPRBtO/KW6vV7h9hp34/fOoj58UJL6+VlWtWv6I26/uWhmYBygdhD/Exq0nuG2rcMtUU1hTt
ZbzmsYK/dGMYGicJFXU4ggluyJkzavfM3iUJ4U0LyUR4lYF32u9J5nkk9HkoYD7k3m7HyogCq5Qr
hrm/ymWosHDv43Poe44pncNMvyYysq+xQPQ9ajOMC8wWIhZdjlD9E4lRQ+a8wB/hf41GK3rbAfIx
/4noA8z2Suf2fFJmpfHAv3INhc0H6v3I8PdtRRidRlXT/3wOfDYwj3oUlgx2f4RZ6IrDzlrZJNHS
AMJx3TONuyThMYKJIoyBBdkVEXqHDMbzgoh3EH14wxNX3Lc9v0VuXspUcLwJV/1oZIvo+UoKriQm
0JtnOhgMnvzED75KlvER116Q63wfDzmHuyirTtHweF3HEVYU06dHBEZxs3fkfdLBvIJzoGfFpYVW
AsE/Iu8ASHOK4/OeObzdf5ADjXZxy1PiVDPSoauLmYWJ3a7H9r1fXDEiSCeGzrPHyelJ4RfSpjxo
HoeX5D/2Uo11SJHYuoYmSaaQVNxU4i7S2al0eOlcu4jFpAy5wRSWvy3DAZZ0VDLdai3fwIK2xw1Z
X17rKRhL+2V2lbPsNuICxXQl/1jHR3cjYECYO0lUoEaB+bHdTE/uhdQbhv+1tDjQO1uYCQCe25f7
e9h558C3Wi+TkuWeMJOZX8uX/5aI0jIuz+YUB1LsgiZzu2XengyA+bTPpAxujTSIR0rqsuzMevAT
j7SWwFPSWCRwtNicpBCr521mxuo2w/vd2JeCeXPIjUICUiJHM9YA/Y4zEdk55SqUai/RBw82HfZF
euH53J0h6oMYQAYOBgoahBuN/Hnvpy/fwh9uOijNB6avxUirCkn7zgZnvdkJY8Uj6+RXYPOT4GY2
BsI/No0mysmdPQQJ94QIluEN1pAp9AKZzv0l2U7zJ0vRKKLWI0cwu7S77FTZklynwgbMoAHfFcAk
RHUHLDpYU6cNJLnSkvGF8wWBKqGgeNJR32DhTVSUYLc13kvVV7u1XFSCMC+ogSNb01Y+v/35Fgch
cC6wjzZXItUmnXvHF2sp3SBvJrK/4VCEN1he4qjcl+g+zl0Cjce9HUBaJ8Zs1HdlyZWpnrrfUcp1
XPLeg9TYjtHAQj1z2jTnotMTDNO5sojjLg6t1EjnoByXPV85J5//XVeyUmamTdTApwwbm43+W+au
LSlgvD5HmjakkDhhFm9HZZwIflgxnY2rZmHlKEcXQHNMIiyiUwadvEe6c9Fm9E3+GYpWM28Zxumy
m+CZV7xoM/Y5mnFEjjPK3Luzf4HiXANmHUs3+W40EsN0jhTmE3h/XOCM4ZvzPpk1UDe5XFt07MMi
QFWzIk8+3nT+TZ0ssE9RA1Pdl53P5O+oLxTWoQsUerMoD3Li9z8d/N5P01X38OXjjjZMkmTYxQQL
eq/6rv9b3DPMPBQjdixjGuT7Bz4o4fTIPt/hF15k7WsUnPARnYKaibQse22+fUPN8Lgl1oZaCAVK
KlTkGInyu3ad/3T6+k6PsNnkuleKK47RgkgB6iFGsfA4shHNhE11z82dWgnBYr+HoLF/Eum8fpfo
B0wWHUvnAQnxmg9CDgeEwd5dRjdfGKF1rw6UvNIx2ZAlB26jYonVCYcK9kmidp00S2VNZEMZNy+n
5KfG6WSbO5PTLx+OeXYIZ4NRl7PgLchsvrNKuXB6v+Sif1PeXrwnTWMBRGJ62LWs4Timjhf62NZ9
v9D7aoNlGYewloWc+A2PZrJqOclKnWFLR5CBU8MVptqYPO5CCzHA7+JjOmS5M1z95xAUVpqpo5bx
PNS70ayYDnHijj+XAXQCOgxqJ4IaaSqgvafdXY4hj4kRlfiqTCuuDS/yz5SdMbKbNGhixDy8rBIg
5GxoL4WitjzMGCA4Xd68Kj6L8C10pCpCb2WSY6IPqbbAieHAwA6JkB6nXpY0vfdgMqQQCHvDoSu1
0VdS/2TmasfK4LOfa1dNTZ5kbALT2E+T0mzITL9hxeK9xauxeeJ1TixRJJnMZqfRKUvol4IZA6hb
aamPmP28l7k3atzBhiMPkjhRVxeOdVL33ZVEGk53m0ofNPcN20MdIrTm2Nklt7SEm+Uvdf/WqWrV
MLO4W/CKBPQ6uC7atdbQejR10mBxMSIpP4vIcoRZP9F/0WsbGkYDaD+csXQ18JQmTeiXk1g+Wlq2
ENH9fV3w5GJRfIqZYUhQLGELWS02Vg3NLSnKebch+vyuTHkm78dPCf3RE/ucZng0dXzN4fgeCn/k
4Gb4bVpMnGXJs/9eB0X2TgSxOMKCsqkZC8Nm7vjjubbScWE+1a+ltYsKLsPMAkneanR10l12qpd6
6V9wgrME3gSs2EkmOJh3Wh3GO+lpGikWcP0J245WNQkdnkJRHOvQreJ2YFTXb9+7U0CNGgEY5s23
1gmbnbvd2ItoyJyJ39gfs32nxxC3TefIVd1gwQiYDXvXdcRSSwdnK3rq2mL6NAPI2RHnLHXn46Xd
Xo/NWkJAyire/e3qRyaHEfKT8yBLT8zUcDgeWpV4p8zt8QeEaDRi/FQQnlf8GVooOF2YuW1c9NNT
wzk1NwfERyXFWrkmQP347LABpcYlDAXjdYUL5chass8yNfzttWytZoINZQjr0BCHtWYss7RYAc3O
KyLIRyhfOHklHPzFXLvexlSnFVFjWlj6F42kTAec8uOFjqsdpfq9EY8aHuZ1+SdEWbubH4KTKcPS
u/uIBh1qTmsEGRl1IC1mghQKYrMAgFHTcutbtIRiBuBJ86C55MwiDNKHSGK9enCBDTgbQhc8gISj
+CM2FbY0Cu4Pj4Cq9FQNNC6tPhootshBYpC2dzd0w6hWj7OjnoRs+Vf2/mfxAzMOzKAKROjP8LkV
cA0ZDubwKH5Ko0zvFl9ogHTsBiNCoM4nzwAcM0I/oKJ7KamVcBsXSS9Z0Jp6SmXGVmsfD7ZSeRfA
34qaaXl1fl2xsbjH1y4QhgzZO2DqjuVSEQCUaQJUTBW+nPhgrG5DrFetGxU7h/mdFKbNvj8WZnyA
fM3QcICdu6ZcfqzcUGVaoK0+wh7hAXCaFRHWK5TMKt/xIyVu4pzIkNGMH2ZPycvoy/4fj67Oy78j
YJjdD1F2LNrh1l5opJWXE+Emh7PFH/LSTEcIJfr2pmsRntOd/P7ICsv6FL8T+Po7esyPp9Lwu7Mm
z3w2xWcpTLb8irrtTGN/QBH9Im77yixOuVHhSpotf5UqkiKRXHCOEeSCwU56XeRV32pu5bv+buEa
TIX5QM0G8q8mXPbnG9ZRrxtIljJ48NWPcqI/ngTcXuCbthsn63as4J6LTmsLu4iOkiXulniTumQj
Fo2bRMsDYUPHPmOP3rU8GSfMYhkSHtY6mZmKnP02N+9h3Wlu9CHRjcoJVK4aLe8KHv76btLZjQiK
WXiYmD5V7jsX3aPZ6BQ+UiDwicSCC5PH75Qv3YlGSSjlH3hNqL0VgOAU+sLKw9muSJLV+IyizQq1
1DT4e+KTPYTQWDRB+hoDaiy7PpOU+jwtuFDNnWtpCkdlMAkwLlqhdsnaQxJmU/aUU4NyQM64nEQ8
bLcD4jt82BbrnYzh/nVxXVc2ZR8jqt6PkMKp3qOzg59pphHIbAZAO4Z9QBEW7j6asXhqElK/5tu9
CgGdk+p/BVFVupxH82wKXU4/3ekVGZCqZV737qkMOO/mKNp5Q0Q9aPglP5KLj8qC74HFbaI2R5fE
xq/0oTULphzYGPT1xwWBwSQ1J+lLm497P2sBta+NisW4tZuBFuQ1VB4MeP+YPwVZc6tQU3YzY3ni
gIIJ0cEchbX5BtRUwA1DtIdia4DHMbq7VoRSoFskOd1mPDOHvB5GkMinduJyl0cSJODxSd3bcnsw
NcE9NuJQD9dPoO3RcU4VEonVqBrKbUy/eWbp3hDGkiiPTVVSzp+CZR8hA9MC6xphIfXzhbMXDYr0
56QEzmAvHsuUWtlnbZbs+FUQMH0wIAu5Drz2/SbtTqnoXvfmxRDV2MDrlDKLXh9KSc32SLdX537J
fCAjYI4TsxWJZ+GGeFhzX8cb/IzrZC55atwac6JpyLiwm68cCtm+SGEUK/Id8FU8Wucg6P3nWJze
l0NePVYjTJU8XNXk9n00jS+1sPN6jZ7v3kiTUekIsB4ENwdGytcEL9xiyo3ctalQ5BCG80Gmgh+g
CqSH8s3nw3+vtdaAICN3X3d+0kFp+SBhwEjAb07vw0rsdq8uQseAHzEL6pM1sZVx2xucjbBiDizO
l0+C2QOXqjVM/KYkggv/R54rZN6geS06q4JeW+9WiaJwAEnh2CTrc5eM5Yla3v3YfLF7YdKmWLRL
VGw431bqhBlUtQwFP6B7lwZKGDpAbOC56WQIJAS2cncWn3LEqrLFpGP4df0jeu/YPOwIBrRZk/0d
0zMUQwL091zd0yYDpXM2lQ4N7Grtcx6iPawPOJeqBStxQas5ThfQsor5ReCxX+V+pTyPMEc2dK34
H985l6EzkbbF1li5oz1kIFUlGyxYx4wzffignanXEEn51L+bZK7mcWd93+kHaPeOE2+mmvX9NFGX
ZR7Xw+T8Gv+nd/vluS37K/vRSthQlOXIZwYxi1Os9Q64NvGow7dNBsFE6TLqg5vuQoiGP9pNPCWX
dqW7Ao8wu3yFcgBnuBzoNN2xWDwn74bQXK+fjdPRZxNo8f41dKu1H/89IAAfC+IOCoX2chjfEJRJ
1qmzCRQAs42NNo9ts9KTnWtkvii59HWYoMTnJvR+bLx7IIuzvhcFqrQaX0+eO1XwqrbJq0/EC4sD
8KdbuLB9zVLnMppYhaXHjDef4G/YaVpAJqLjLawnyqiTgIQdfZjrh7fY5TMwJpRZw2IerMb+kN5e
/f5gx9mHwSavmNmF1+rI1A4amZEFpuYD4INYOtUkLE5N+lvXkFEwMHKOXwZ120AfCvQz6VvxdjP/
7ZWW3SzFWXEUrwnSwddQCIrX9QycmNi/LgIJ9A95DyxX41yc9Ys0nHyZkdVLJ4b21mRPUFJsbyMG
Pdme9d2tgJcnNft0dtfPIriMk4DMzCtHFWCNi9DMOFsqZbktvPdksJ/Xjji9deO9YmN4f7r08tuf
xjxKyoYahRkZgGTZIdkAQf5qAVaWGiggM9zqni9CmvDwsD4cx+IcgA0aYRc6E9gPZV3MrJhFAROg
BsR5BcpDHi6PwQsNCTP0pBtrwCcwpSZXwi46Vi259ZrgH+zyTtUqK2NZGAGOXCmXlmh1zCC0nXCi
beeFQTsuccQMA+W6oUxIcbPXB81bl4ebDT+kjKL28ikT8f45UrQ5eNq8qv0JhSZBlWbpKE10Vcby
4c3qoMiDJPmh20z0HsiAO+RM3UgmpReE/kYKm0ASaEx6rAn7zy3gBapRPSBHcgPvIKLIUG/4DjmI
GJZk7OWCJXNaX5/+7osqsOtQwT2BDGn7eJj8me5CQur28MnYKaK/qECl4Sjp0nGQgiypButxaZY3
27KrLMymlG1iLaa0p69FxqWEdaUXkA3qgLXXt5bcHa+IUmTxtbHjz2ubXG8Wbzw1FtmZ8WMozlES
cRUaFPWzZMqbXXzcXe+PQ8KL0RdpTqSVo+v4RMis2AlJEj0cZsrN217eQk5Z3KWUR8iuvVi0+Nkd
OMjN1M0i57/W+/kXoFDywUYX/Vn6y7fc2O6uHlWX64ZFM1ItZ78uC7NBZGEDeiPOOqM5gYJmJdBP
h0hwsofYmNT2/44QEWBM0ufTwQ2aTbsNR450siZ2l1Kb+jo8AT7nFlrlrFA01cbSWDORCeGZc0jC
gHzqiqPby5AkEMByyuIsgSP+7fv1n6AGwpmQyj5Rn/slXm1qlOSEK9oKdBLXB68QdQx5GffOilyX
jbkcm/bZBlct99ySmHoGNTxNKa50ByOWQku8Rns+W9CDvY/9faJWWL3Zai1YNGYF1kQ9as1k1SeO
tLkoqqrxlgDuGu6sXQ4uN7UmU+vNQbEvwLm1B7Hn3cnuN1yIV7JwtuvbW40tRFIwO3zNV1UirgH0
L2v/yfmH9Zeh3CfvtNyHpp+JDcMhO0+kxC2TRGdMUqd9QtktNDVV87uiQvXqKx1dVrHkzVpG5FF5
RhHkH2MaRdrlc1RJQNrymakG4+3Xjlx/hyr0RKr/yz+VUVgrronNrL/fHek51aTsR8OizMIc83th
sRk4MZAy8fLjPWULMaYnhN+YL3+p9aXWMSHBGGKdm+a2jq6TqJ9APrZHbGIdNKHchRevZwCHZqh1
Jsor4ijX0Alj1r2EvdOOxF2JNsuzgl1sN7p+N5VE/i1Ba4arcZwMvnvvZiXZtYD3sFVp6nvyV4Wn
neOVKKOVyzHrInHooAoKIRE9JvEcxay5HkOVmX7iQ5tJUX/yexKP4p6d8x+UP/hGud/AZCJnwSkT
dncRBEwe85y2/3fd8DKQ1+HX7yrQAYXABJ/sUNYJTpmeiiaUYvZHC39oC1bWnB6q/TWlNY99Igh5
1j8Enn6WAhcDAYSiLr+JfG6z03NMLr9fFlQOGVP+7VMyhSU8BDFGWuxqpcQZQ9yrJjzzPqGF5RsN
cfYjDM5bhHmHQeMkF3SpKwyCX1cdKth8FYu0p41wV+kxXMOJ+7P8JXczcsFZBFPcFEGFdqAqCjp2
eCYCZvxvDwWOQuKmsfOqdm9POSzzrNbOpFGcerVsYr1UxPBK2IjvqyKOSj4swKUe8uA6VTJMiBbF
X5c0eYzXP+CT7DV5AJ8Oejdo/4GPCXnvr3SwW6NMkBDNa3YsxKkeSxj5/Q6EclbCBoeIgrFcg1DW
FV7RcO13czLIsHPrKzGXW+SRqII4RauakPYi5R6V+yvOZWSHQXiJ41c1zt9EFyQV0aPTZVIys60j
gEPe7xX51g9/QHjaHH2teUpXIxxRUjM2pcePH9RP03bvvfUchrJQwWCCYqswob0/R07hLWJUGtmG
4sXD903zhj/jgNXF1A5y1zrN8oZu8yiVCe53+q6l3CN70ncZX2AXnC7BurUlB6oMyaWQtjyTG0ds
6Rfk6R66IlNNwbV+X7gBmJc2spXtsXrc8pILLlVGAjqy5HSmfCW1bzJ2QARqAPzlMV5gxk21l/SE
UkTKYIa013TaSHht41e/rLh/FPhayqd36KNexzZ7fAz4eoPGtq/UQalpbYC1flPNpIcttmigy94N
fjwWW1c+EnHA/Xx2MmM9C9+uCJBbRr2gj5+Y+cJC2gd06Btb/qTMb8D8ZrKb/Tjel515I0ZmJ/EU
A0M2mt6wog0fO/Nca7htY9B1HRyWVsXyXh/NXWHPGBAl2KsRxSWdq7YayAtOooim7A8o1a/+jA6b
vkTYRLAJWwLI9J9qVSOmIZN5iQ9Kd0Em3yTjMS4asar02sB7ob35vw+lvDlyKhh1x9c+o6vIeyYa
N9B0zL3AutZL35ujzsApQ+9/j40TpFIOQcYvk+rbVD6rYgW6ul+9fpnqtLOnH8waEHqNAdAA0578
lWhMsx6PcTrs4Jq2x43TnDIBPPFT5wMirP5dRLb/fvpKI94YKusBSTeE9MZPrcRMo3vrDplUFUV6
931jaChB2XUh/hByiNufxVhAoVVWDSy/kylqXGC/HGasZjcgFD+K9cmudLpEHujkvlGqX6Lejj7f
BKrnh3IqONd5MUkpTWIwK2BfMx6zVaVyEC1MMPmFfUfCQ2PYDUdVDInGnQQrnE/rUNNFGu2CuXGG
mehQw9FMbIb3VfKY9BZDGQzqQhBF0MFj39Mamv7U2iTJbJQd3qHvZNUK14nDAUBEHl6JGskQq4C+
+nZLzEbwb0PfP6cW3EtPUZWKzK/D2qJYuAxAZUcqvivHnAKaxeDh4ltZeuvNkKfx4/d5T0CCjvHW
tFGxKQCiA6xpCA1bwYyOaArKtROgM6XutbSQIgDXE01XI867XPtaMNhv+lauzDbeEcKcjeR0eWn+
LouDzNY5h4qk7eKnDdWcEZgitbMpV82au+uiv7oCEw8lwMIgwTn3syYhogytvA5dtsGX/dN25aAC
YuB9ep2jGml4sLWnVXzp5jgmfZAi37/BTP1PjYy7UYEi1NXIW7Rd85exVC3Nts6cPhrrtG09bTeX
Kcd7vzGP628oi+gHOyRxup9vGHywAYN/cAtyt7wLKMusZFVFMGTUIpKWREqttbVXd7vPPyQh1tGT
ZBE+0FPWZaWknLFlI0XpWosnWERNyMdVAMswGaDm0cctkfJm3Z1/P0JI7AwbbLqVEHlywX415lOX
le/2vpkTB3+NPzhT+PmYCkRvwhXq2YzgTQFFb/aTNp5SSCEpSIUGu4KH5QCl69XA2tXrBlFX+BDJ
XbLapjzIrZXIu14RyWUqPEIeSZT/LuOG3aivn6C/+XmLUB/mavY2CJuFOzYVQkee6EQTwcg3sGlu
KrjBHNezDpilV3k9n9O8e0Y4Dd2ahxk+eLgf+YQRwLLeBbXNH2klaLphQhxrHSqRu5BmvxuzAj6b
U7PqhCBCnPXIUmik+UkpdnRJtsxCnaEV6/DIqL4LUuTA6+XG1yRMiw+aRHgA91pd2aIRz0rGXjXi
5i80q+H6tPuZy3aF4oKLHK202xU2Ec0EHBcBDUjcEYCblbOJqrUWWCWsKiackFrCiFR0l0UxnubQ
tNNeKs0XpiTr2maIT1wo74P5GZKvcIzPnW12fDcWeWMc1O9sw/claSR+9rdtOhZSHzDC0fXK1mZl
sSq5jZq5dYOuV7afXhrqI41ZxdcvlvNtSV9WuIuz+o56f+n7wmSJqQJ+NiKF7bvDjDkgVh8xck2f
wbE35S1qkbITkzo3UDfFGqjzuf7KcQFdIEOX9OhpP4frfX2YqLAhXsdnm58EI/5PhB23wSjnE7wq
/N8zx6Urk0wWdMCOnxoIk85BAp2FqOgoVfZH+9twKJQ9KvbqZ/yUbjZ6cGiCrXBYVX8OxaooTHvv
ws4ZThPIdlYrSj8N4mVe01rSC1vEIw4vPvdeRkDvScpIuFyl9IU4aCAcWRAchVo+F8sdUjHwDsdA
EU2Lr2a+60p40tG2/4g08473yVn0CBfqBFkAE8bcl8EVAfUYZu4T6sl0v0h8BSdtMB6UALkxefvE
8DzWvSejqJ+OwRQ8//9VaNMKDQ+NYBGSK6L2eHPskthPlZNtTiC6lmarIEsYCq8xkZ2XNCDt2nPS
tcLesPqEhIZep/GnaHWmSqx9/ENpwFp+wIHalbisCFscIw+hY+5N9OyKW1ArJWNLXdvJhGYhAUKP
wv6dWr8VXTnDM2qLGcywxdluIz2pSxOkqlQGMqeDIkpoJ6Lq/cd8U0k6rWKDz8SyuUMMBk9C//Xr
gI1nLN0JOb3MYKrJvpEnkNff6yKgDv0gtmYJRjxT+bGkcoaQVq0K9aoJPRNw344biOOcx2HBlFIs
BA4k/LgHfjoZ2/p1ozQDV2TFGjyBxX377TvQN8NHtgPkYpcV3Jn/GjW8hy0OHQPnlFdrrX5zbjct
oLFZX2+39VHWd28M4v709oLG/OdjMLJmaXsonc3d5PYvABFC6efLn1HvPjV/b+7x3zTy7VbL9Md3
+GOeTyQHiJ0xlkFR2i1K5jDx588nOhU5YFmoHEi62nPSFayVewsVbS0uhM0Mc6nsOoo/EiLSB8MK
tvfh52WKQUVjf1+p0RSixLWBYZMUt8C3rs4i8VrUZN9rgCcUceD6Gi+qpoDCrSAOsVjTGTL06Og7
M2oIdyumDONU/gid3OZSbvpMMXVUJKQC7LvWjYYvh8kJJVdWQUGtim7dv6oAHIypaaMAyLmzlfSi
pS73Ta5e9r1rZ8rl2l8APrmVNC+xB96u48dWkCZgpmnWz8pemYbM2WLWqpjGGFtQnXeSTaIGRNWF
nhpIUwVNTQpTCaSLZj9zEaMC3kr41iXknfpUIzTxqG5NaamawQC7U1KXhmSx47v2Z7nktdeEk8I9
VQ8icMo7HboBX5f58txICGPUdbIgvpFeUo58QnEvjxfCbk8xXNw/w6v0R4VR06LhsZy5N8cqT8v2
RCIvHg9uA1puhm8lZHQVflyIK5zkhF2xFVVxqcybkQ11eWcUDydNw42ZmiJTRPbCmU1C9eHmMT/M
6bt2/2LsBYZ7YyflmJbUX/d/B1VexNKEb0NyBYBRRFFEzmTV+WuLSWFvFmiYjymceERWeuFY8j/F
mr89xVFQ1clulcO0QlDdmgEJiMJ3i2MdQhiu/0AYzR5569ubs8BuDb2xLFETDShvdk5/Odgiu0KM
l1pYlebTxyClcg7LdqSwxvsCcvcW6XFrKLL2xrZAdoYj99NIzoRx/rfcKf25p5h/NLNbSOj/brPb
p0Mu0eKsEL+C2B7PvGYWre8Cs6yQGciIr2f3KOTvmmmHVrChbV8Jz/x0iwQSyqkoCbeoFrX4J4d0
SX/H3P8mT5RqAlQeSST38ZhRACjxJt7NxPHcHt3IhRYQf0w4cfSXtllUJKIqINd6W2gKuhF2QFy0
SJIS0zcJGjJTcuhtv+BZBk6pkCTShjmSNs1CNIo4DmJl8pBfIVMm9qVL69tOUxv/lJ/9vo2F6UNB
TkkQoQGNbKRgdxip5BTazsdhI3PI39o1kigkZgfBVQllQIMaFcvascj7ssVVjh69WWEeBg479kIk
XUhPWoIHe0Zlai8Es6KxImprJteU7bi0X1NrXuGjlo/pdCwIqfCL6iTHdzHSGxwwZ4t5tj+ReHXj
Q5rNr6sQTuWqYLrSxdcDwSCT8Ekjcdbywgx9P+BgCSgs4Iz//Q3oavs8kXcV4vkKqchUjdNIjILz
4aH/Dz9ay8BJ8khwtSf7xwG2SSAcJpEO4e4e6JZ76LaWUkc+tnQclXmXerCBxmyCjvg7YI7u8UsP
Q2OpKvEfk0EuMntISCKB8+9HHxH7yijdsXAw28N0JJYakQt6qTFyLRGTUpDv0STdqlhT2RQB5K0E
AkulVs8dwjxcFFDOAvUWkQZqsoD+8Hvp1Qn6pel1TL4F9lONnAxqRmzUlnRWGdHFcsezwPy6VFkp
xVhWRHRyrs8WFUHIGy3fA/AHK+WZOAJ63VYXA33PKQm2GpKekWCPpvWOtWIIIxeZHIqF4rdCn54l
XlsEtgev1Uq7156vhqhg+revR9ci3p+tQ892bWOowAInnnGdcN6PRbcmKxaNHfs1XHRS8kBgAqr6
rjCh9yRfz8B/jsEp7JhtU5ureGBwrYBZQtw0YwYXFb7iGktaALs3nPpxMycHMd1tW6KqUahb9Lsl
XTfpa/En7HuOk5Gsso05hPn0i61dMmJ6UJ4C6YyWnPDCngHUjAaMxInuU7v7aIpw5uXwGNzED250
0a4qpVYkhT3Do+UiY9r4QC1kS8NV2vA2W8d1Rwd+4Y4P+d2XffDeuy5ZoNWIjCSDgSO8OCYKlE/B
6z6HgoZXj7NzOOP9qJK0DtOh5sBV8FfBUCZlsydmuTO7C3wpQNFa4Niu7tj3frI6m6tQ6GA2YoJI
ijo+thFqYPkmrGBZFFtQSqvVzZMTc6WZLj9Kv68v6erK1fpIUvGCYhVoNQ3HBbMCpUAg1MLvvOUu
j7HGmi9fB/vChLyK1MvmHKwMiMVFpLtlW7zjcmxsj7f0L6uJ3TshUH/2rqWQNma6wWc2Kz2ShXf6
R88BW1kMrJZN+w2rOb3T0xDXPgO533kkvzcH/10FH6tf5drzI2OEicE61n1H6g1k9OixjlmAGMQa
+7GCE2QhgLXCGQFvZucRcNWxSyRn5RhLZ95JQZcf727Df1yNfbaaqU1tg4zYoY9gpuYbpJ3gs/KF
P9QwMuXzDRiCwPERwR9T55qqoQkMUOCY2gxpdPdr/4BgL+umQIICA5iGNMdByCW11hXlw0ZutE0b
kk2n+7Ax52NE118Kl5fbBocGpGG9Rl9/ravyRItysb51wb8Di0SvUFWNiBjR2vxZYRo4rqvpNqR0
kL7GKL/SeUcNxtZgTSaR6l2ctCy51wvnBR09C2hxD0Gkrx9Aea3i28WBhlF0gkl4pF/mh3QU3vym
gGv9voiMzZCJsc+F9uzd63fYGAMShVdPaq0+vuX997MDa0jWZKj2RL6u17kMGsh/Kol0mqAj/8+M
vUq/QzB3IShvMfGvV+PFBXJXlMdPT2havb3UTp1cbyr+nECxNmGahLhIMq86JlYCV/S9iCLQ7duR
K27tmqGgdj5QTVYbI+ZjKqd/LTJav9xuJMz9RgMF8sGCR8V6UEpGVpW8qZMX+7Uge1XOEHXx9IuS
bTS8Kak+Z/p2OyBBLcQ86GihbK62oj9NDrk4f7AmU0FawuKhqeBPpG3SnOa49ai3ybkbHmBJCYwB
xKDGA9OmCMk01AY4t4sA08gEQyAiaqPS1KVKW9g1SAS2rnmABcHU/fhVpaZh6iHrl22J615Ytoad
qLxeGIJE8uphMdHyMs5gjkr/hlnW0DXmS4AI7WeSlvWdu5xLeiir5/LW0ZNwQtW2KHBUc3DNTjEx
CPVX5X8aMLYb9zcGU/HVLL/wUhLq9QxSVwSca9Oz8eUHge2WsUYaomrqLaJyooShlv1xa1JS8j3k
mNrWJKMq1B4xhcNft9whBfsK7LlExJAAYz6uC0gInMEnFxwsOdVHopY8iASNT8DyQr3i4PuKoo5O
g3VZfzDbd3X8dSkwfYSJN1uNz8mxpbCiA/UA13hScu13/KbSXP6k/3Cxjjn81h0HH/+fiBrverMU
5rs4vJE628LYpddKK0hyiUrWwAEwy2W8nGHO/xIiU0fJ0fPCE+z0RCo5QEa2Prtbz0UzIVoE5bpR
GZgxXETcax1MHUUYz4o15032vdtPUJoDCovJg4/abTD+MqLQnLp0BU4j8+adJlsV194Vca12X+XW
WlzkmgsCJQHIKHcxyewxqv6bh+KsHpjajd08nKaOzIp1kYB+ocktmjP3zmkugBFg9CiSEd+RERWS
TYiCTu6hfYbJ0fbX/bC9WmS1+bP7FNEB+/ZJdDtyJ0WjrMqqE2MRgczurQxDwQmXGJRJYkenT1Iv
FN9Z9vgHDaElpRLjTUWtqESnof1vCO377m2wnvIN1iG+Jx+zAne0ecVgNGWnp7/MMxQy3StAQdS8
ashoH5A5UppMjpWzkjPTqAdDvbr93BCU8xuSzYrDl26QlZK9sZeqvEBenADSncmly5OtOxmkSGtN
h+o3rI4MDfQQMkNoffvWb5qmUjoyqoB6hI1SghgX+/Drai8JCFhRd8O4nv0l91Pl1PZN/+Dw/Cqp
pR8Kla8UPSqMPe52Fs1lmR9XctfPteQMQNxG6T+Gl8ApIKG4DPkHhyaYgMa9HTXE5/5tF7Z6GjQ4
UgkZxVvvSTYS7xvJD8K8zuQe4DPLodTrgMgjoLPKshLRb+7HCtpNUpnpUv2tj4GMqX/EBwYJKpn2
F2iTG/ZfudcoTZ7cck4sJvCTZR7Q3fAiBDiiatD6Leix41394VviZySD7OEA8p4Mb1J5iDQQeScA
3M9qpcRoH2VwxfZUhOD3p0QNCyn5/HfJ1Ps+/JnygirjygdKAtfh35zt/tgaGcoe+c1K9bwWmJ8S
GOaPlt3gs4gHcbFXXf/ADjz0JI+EVxGuwgbdC57DMq7W6GzILfibpXJNSZLVyj6j4MS0w+UrNBQG
z1Z9k7zuyNNewWfoxBpx6GgY75iRaQmihTHTr6zcKtmneul3brGaKcnFz7yYnzNulJ607X7/G1dQ
NLAzTYTXHxmWGTpxVdhp79+lz4SOLbMzl2FBx//+CG4aOFXAC5FtbmIWFtBvmvzYG0C0/frwfwKk
8o1Yz+S2C2c5tkBCcJuIKl14dQCfPwiilTMGyoIqebNWIE8GW18Z1/nCRTWlYT3BN/KQlM37MbYI
RmQ2DqbsY1BnExMX1fMpkXlPh2tzP70Phby3Ep947UNpIyDoYB3dZlXkREL6gFcbXEzZOTg8aQT8
3tF2LvXLhVfzx1JR6B7+mp+W7VbeXhmhIpc1kzVpxVd41iv3Gp/aR+NoV/b6RbvEEpiE8CDDqZdl
11ED7DVmm7ejmgQrdrLeClIydpykfUU7nMpIcVSY8FgpNWMs7f24wBAH/3ElTRdHFOJ6DN2bQfGI
nIbHvrv5KPN98DSyTkL2LrRtD/jM90XC+AdYz4bgq0SgK1boyTtzasc1wYrs0qxsA4fux261bUch
5BPYi/DYY5dKWVklczFXMKrZW3ztrJI+SfWW2/sq1I4Cj4NUkfGCsrN+UM5UZ2xiq43Z0VqJOANf
geWoaTaDtDiivsDeCKbx64tpPKNgGooRQxYKqUIVQYgz/FB9RhVop7Fc0TVSBRMX0EL68UDZT8Mp
qu7QrEy5UP4H0zw1qURDwPG7Dlqy5upeMeKQWZL/oMZThWKQy266DjoTuN4Db7vQDj5lY7BS7vz/
rBTiu3r5DfY96z9RJIUgYGeOw8F/8bftGMSmw3n07KERp0hyC3yYOvJ0DZ+6zy7qn/1qZcAbgmez
l1i90z2Bb7eySTm2zsIdXPn8jBt0L0sUm8wbBJgnYCFyVbMBNuPVtE4AETTGXWYlzt2dobbjoI2O
Rr63eCLaT3hZgwhSeFc38qywaf1JqIYY7977n8lVSsE1iYQ2xcJ+7nvGOa06ENr7dszX1pNdZa+t
345g5QpVjDoF9NnoQ1iZXJrf8JndZsS4HyX9YxzH0WZCqoXZFM4Noyv0i0sDOuys3dxrnqaDRiQP
MpJ0hT27baHb08iunshAkQyZMGK9yZobO5wIlNFJeXTUpjceR00Q9CJTs283cSt5HSyoyUJwPgyj
Mb50YG8YYHBUyd9aPzZSA8lIzY855iQn3LjEf2pzD6GA5jofZC3Ai+ZP58dlv+itXuF/joYz25S9
8ud7ThaCgr4shTKWLEldWyxZjUID92lZMNSyrbAi4CwmRG9z/22sVGd9BLiMy1z4ShJ/faPYtII8
Z+JUphKsVMFb4hH0N0kwsr7Pz7J7DJ9pxnVggRXk29pjSEwh/B+aiGyJGkiueX9IoJ7Mk9U/9sc5
4aX9X6uSc180QGGOlDFrL6kp02MZjAO0S+NBo3ArVOiJqeCBQd43bFXyFxu0eyIlslXkDBTFLtGY
4xpCBfZkMIMrrvRnaGKvLzYhlL5RHqtsWOfIXGdQBN3cVTYhmD2zBSXNysofON5qjAmXnPCmYm+g
ejgCUReX6wyzYFBCE2DrCjqsB0v9DONAi/ukiGz6p/qGwXzqCGndqSLKOnflTf93OCtNvvgyHe8a
RlSdSsc6pss9wxmpRXJY3Gk+aAk64Hyb9nq6HuPoL5+jRKaBczGGwBy352eVyNuUe21e1+AnG0WW
vMTIwI5WhRJbXrcjFgSf9AwAcZyyQ/Hoeej7Mz+zk2bYUt2TH1N1GsP8+pWlAW1hi8scWIIcPOWz
kMmLYGvdN4EzSHTA6GfasIbuWfRhclgJpKIGp+n7VkF0YFMP9SqrFzTQek9CzjXfnP6Q6LkbS5wR
ZKKWCEV+TctpXhXKaF3WmMAHecqKCMbXZ1mESO8/9zVfgS2ulKWz/KWh4HntKEtfieC6HRM20/ek
W4FS/PI4qogzDMPp9hzIzVDZgxEItfJmTFziJYzV8+26w/1FmQ4ojHkf8HviNSuEv+oL+FGKLl5i
G+uRkrge93fpFj44IaXwwslIsU0rKQuBWeEf3EYcKvUOG6IRYcpqMgCcSZcfY2G1BgZjSi0IvCf2
zC+2EmHBCHGqaGksDGSc3ZFLIx2JSZ7fyQeSru7yuHF/aGJ411y/juNDBYQxO2MOncEiz+vMzUuO
g7cbkS8KwN7lm7aWaejGf7IrT41skl5N4kf3QT7mJqvAvvquOCSB+JXmFKTE+vj9xpKuOaP5A0Wx
HfTwzjEmff7CFoZb3cpZnR/wbHVqmDPdWunHCPjq36DH//ENHQ0P3iOYoA7Iy2y5R5Phv37omsZo
5dcDR6Cm5CThmMNR88zom4RQz94dtIRjBAMVDB+d00TvNYRB06hK2IQBMpdUGCXgRWNwBtaeCMPa
NaDoWVLALCgpRsKZpgSmQO0dGA1u0Oi7q94pjNW6WxKbxlvG6FD5nw1DdEIdF59U4X58FUD8OczR
f2DDZfgKgQ7UH53CMThiVgZyGen82cOn0zhqWA/VqdUtzoJcf2HHIHqKm54weJd+ZuYgTVP/asY5
t78KAd9r6/L2sSI7YHFz40xpu/eiH2fDQN09nBjp7XG4t28HfiRCyQPC5pJAnqxD3B/8nmUbZh2L
DlJvcbt8p3n8Tno3xWq2kT6YT6p1GX4LcRqJnM16ztTlwuOERyNb0XuCkAtUJMRhm5CIjlFJIsRr
vQ4EDr813d4QAy8EJ0ygKdfQ46Eld1Iiw2LjsgAEMjx7Kgn+IkMxtMNPRtO4T7MuhUDzr19kE/Lp
nDRsY6BPnFKFyGTXWxOPLJ1FjcXa1UIKxI2Cx00hdTlVfhsCzpL/hTBoOHYWG6cLBijI8ml/A4UK
rC60k+aXkuKQuVlhanfMA83j8D/kVHwztaQsRacGPrG2+IBLBwG7zIUcl2SXEs7OLymglqmN/H+G
iDArSKD4fooqzTHcugI8i+vc4923Cn3WQk1flLV4ncSzRdnAMlBoZ2j6KG2O3AwwKQWz0NTC+akk
HuwXZHkpyQ/8lFa9cIqu6sjH/pP27Bj8azyBKSOJRT7Czob4yDhMLglwDmJyGOza4UnR7blo4MvK
NCxFhHVH0U4OnaHXNXZ96HRcV790H2GIOWCe4dlAF8Rzi0QGTOsvj+S71RBYZMdJJueaQNZsWXXj
mpU51Lr+6/OHmuuzIQhgw+itq37Vvxg02od4kHNpQKHQSBxQhV5Gjkl3uec488mM4oCcBc9ZdpXz
QuvXwlBi/3labHFLAddn4qse1nuM7wJwKRTdTLk1rofmgec1N6hZukcmoG+BYpLtiIjx9O4nHSBK
J1Dk47v8hV2Gh7gXNpxFsyXqNYA3B2kzXgjjK+hoWXQg/7ayzg3VUsb5nUNXJUL4NaLLJupLyIX7
7shjHIX2E0Cu0n+BVacD20jOilb7rtVWqAtgqKsonTcx4GC0IM3/nWjp7gBY/3cCq1k7sHBW2olr
vZ3Ol/JJWs8JxSw0PHIuJOlqoEsMpoJH8Wzk+iCcOdNI1WGRbTUnjm/aOhES0jG+43ypKDutO6Fz
XwZlg1v+eDw3SKMyOjIZMklO/xwEFDgaHgHjNOtQ0rPqXgb6edTjAW8sHhfkJn9ut1hmq88i6Zyv
uCTAwyUow2PaW03F895DtsPwXVc8z7POM/zSq6+RwWV6ra+PJVtmhAXl1vBhXFOtciy/5Pb8T/V1
8HBYi5AeMwjCLXDC5FQ1xp/N3LN1hvQVmn01ukJRJf7RK5+S8zhGHjGyGhbd0gnWjv1KegoOoRd4
aR/YH35SxcXtYi925gTfiinBS6HCe5regyEsagPDSLbBII2QO64qC6BuMKSNl1N/OfUC/v+yiO5X
t/npaUObvzOuuxXhXrM26PRyxm0i4JgHzNJAKgXkjKQVGp0bw9PrP8cWoiBGF6/p8GbZvSGAKO6h
iYzo59nOrnWQLsRqLgUpnZUPoHmmq2cjlN2pC4dLwawMoBcCxiCiBVFRhbhTmnG5GrOojEE2ulu+
yArg/nK+Dso4mzGafU2IKdmFAH3ZEqAKzgTw51WmVk9kwvkHmD4DCaQa0l5yuneJAHP5EXfRGEht
H0Iagbm9MdBDg2Bsyi//zAxoIluvebPEmmaNcvu8302xaKW6ZjOTu3vWhpuyyFzQJYf08200tC+u
wxUTItM9Ik4HA69K+pcK1RbVTVca57VqkkSrphmyvoAv4FZwnh3bLhE1+dGWuw/BGjGGUK3LSnjp
36BFt8y/X6Cqn7V0yoDEniaBoiNInyQAjzFl26/tOtKqxSdRSURok8gJ/YOrVagn0D0ZXsEYa420
oVPtYEPSXzRReNEeVg0cW3pb6YCFDrQOhQD7Wy3p80MyxcIz2ZtG7g8fLZ8GDr4F8K7ni9iDb2DY
wK7BzQJG32Joj1Tb6HD2Rtv0fhRClGgDoN3FF5zJbvJDcfGRvkxomQp4Bz0ThHSd7gh21Rn6YGUP
3KG8jnSgg6Stwsa/wamCx3o2lZQac3qQ6OZJb8nTaUjhYKGumbubQPyUytVheWp0F/Cjg0IRhZ38
5f6EfRq0ltSxlSoNyVauvkWn4UMSbY6JqjMtVw9shYQBFtJ9eS3j7V0qNXCu4Z3olImMwrs/GsTF
KGwZNUA5eT0US9GmR+xNXzOa4UosQS8F3TN7E6J0zQ28FYTa1vVs0D0kLYbohvXx3UHgCpzCo6j9
BudoDefasHfIvSizVCkU8QE4Pr8NMxp0Lo+Utui+UQgnibAmsdfqzuDw5dKy/btEf9mUbxwU9/8p
fr/cbBsaBZseZdbI+YKzop8aeS5pLkVFh9z5PbvvREv5LuOW83oCmM0wbH00yWeqIp9OJy+8fxgU
znaJuTJhZCG3R5WjsNBwuF+E78tE2pfBT+qsz7Hg3CBVDiJ8EpPNW8UYvJHT1mec9HpW8e1e1jzW
Qyu5A718kNtPZirYaPA/1Iyva9zLXf3sxaQOGnbGKj2jgjQtrVgWVrBe7PjC7Np7Nlano683tm2z
bmUxtBevy8OUCY72HWa1fgrvIjgFz5Nx2L+GhnRLCvPSscAT+ZHQw6Hlz2SzuaSnJu7e0NTibR4J
GRWOtP+cC2DkXaZRnUrxcu4AkgBZEjLKDKtIUVB7ckNU+vS+8B20i2EAE8WVTCaBGlwxstZHRCFB
MoLTM5Qj8Hme9vk8CyoiPKHfHhx6/pvkH7ROe1/Kt0gITvTk6XMbmPKlLN8+GzsJQOBOVYZcJOwN
AuqzZgJVdrggDPM+QjVx2vQIlkGIWvoIeWBg0ISBuQ3EEiio8VcAAAAUfisjKtJjkufJCgoHntsc
InulYhqWiF64+Anp8w/vrIA3Mz07rx3G8UMMSqMGxUN8uOQTDenOJYQjWkd6VtNVeaZHnIDBAZoL
e/xDt861kxKPfCYDfbFNEOh6z3gSOwYGDm40t/Yh5YBYijDOaNJ0Qr+q0Twe+uhmae57kitibNFI
jQcfS6yZjDf7U+fAtX2JXd1BTFLll13dXKgIVqC393JMmWEQZ9GA6+sBJtYFAw69k5QkuhB36drC
BoiULCk3ZppOhsVXIETuAHlOj78Ua8YclGOfoy6aQFIwAEIJp+2RdRhp/4sKd9J+iLHJCBwmfpk+
daZp6FRUrQsjddkhrRgJSoVA8G29AUu67tTlFkmJOa3T4plfhpXiA0G38NDYfd79InvYoyLkRDtb
tIdtuKSTU1H103eocFkJhCjBpLJogWa5mCPWJOF4bOkDa5b6LHoPSoQQFJJc/khP1Yfd73imG2hL
esp8ZsvrEAMNJIbKPyBDbhZNzf/o8DcM7paWYWqjCM06NrTKPc/BOyxwWMsoV7Ey5rH52AwTzlaH
UZe7vKdb4jXlEi9x9Z03Qhh2vbu313KcslUvKMzDOBaf3y84CvBwCbbjBTASTQFeCJN97Vw4Mqd9
ieKVJgJV/5k5B7MNIu7HtoND3FZQAEEQnkY3oY/oRsgsJOr4krTfzFJrRHvBwGLpy+twGoH1Im21
IRjQQvrcstVHmbub1Zq+DdAHnipJ1E1wwR6lojgPaDJ7vUvBRB+lIRaryX4pJQgvOl7prDHEisuQ
ETFO/dR2NY/yDLej8G8JodhshiMryTQtD8tYDBVbt6wpsXIf0XbZkTtHyk9qOtuwdtCSSz2Oirag
EFkkU2/VBS9PBevjaUJASGtuxXy3ZpsifSKyNKe366VseAH2ektbx9fG90zRxSvTSSquXqGMHDPU
QuBBH37j/TNl5xbVkRBaEbz+KmlKpXJ9M3RpniAdgF1lp3I8idDX/DvlbBOTvG4JKaIAndHmf3On
7c9w2udBD8Ge3kUBTkBso8IQCE1B2pggzX72yS6AkJpYdFY0HaK6EDVc9T6/Q5mDAj2f8caSrVJr
HSgGgraNFhnbsM9M48+OJYiV8tWH4zF84k4Rd5US0xy1Oo0l9bYXAkk/tgvjaalIB0Y/sD4Ah6SS
0ABuaFIvrJ+d2lvwZoXYa8Mq2UQIRdbK65lZlDdd5F/F3oh9lCMYLIFrjK4EOP7u/xwYUupqYKCF
fZGUmPyfdDiHLxc8gdJRkcAgfPEYKlzkkkV3JH7b0jb3SakusZyFN0p2jkzzkqv1yOhEGQBwwn0l
P3cSY0kBPjcqosXwsRdnf+CzyWjmK5rAzxALFkT/cVliCQ4B8/hfkSm3ew9Kd7kkfsVxAZn4tvSi
KfnoyvsOPbkWxPJqQGvHYYUMTGK71hmlbvteOi1fTWZg6XnAaQ6oKJzbhsNixsDa0JLyzYuEA2SN
i1Bityn69yPzYYKMdbnvmFtoSOcXHjK6wW2yNfrmnNkPEEF9h+PPKKeiUXdWp5ZcXF5e9rgmLgL/
qC/AFu3ZV2B23CiM/ia4LolHohrXLDxHSnSycdqoN36xpkODXK5CBcwdVNt2yk5LgQ/HH1iEg/+7
PsqVCdkFaCcM9WJsfo6nxyaMCEIzYxLXlGTJegcMB79yXQJA2g2w7IQL3dPMMKzcymWtkilnhKrA
bOoasDUrwvIddenfr9Z/GOBPLkyznqk4QYEuQfUxe3WKUgpuaZzX5BLosyrQjxnily4m5kc6spUO
C1APXD3o7yjp4QUCzozfSrq03DEasyFBSsxa7kYya0cuW9CCaOzDa4F0Nd/+UzdTgfeLeNJEb/is
8QFWeMcnba+RE3BCSerj0/izTFciw9xoNYLzBp3SoNZRvYc0rOjdf1FmRMp1pIFK9Yyvc2sg9Ps7
wU/GQJRzfEeOGW6rmD4+DjO67+ou307fv7U4nB0gyh6Z1LwRf5+5+OPMdvBB6konvGNbaOis5aeO
7Qui+Guzjn2xEWEYzRCfdoz902WjCO/Vv2i9Ckmu3v2jxmPrYRITSE+55O15+GQsUqDNtWBCPrlo
K4TDdlUMqc73Uii0b9GfkHLtZXI1/KrGmZMUkh/jqt7kW27if9J7/8/xw7+87g6jemSUIyI6bXaH
wEi5Bt7/t0MF/FaysfNMOD35e1VdwZnKxLVNEPK7rkIqY2iqb4i8//7yFcdh+nWy1btaQk1HO/Z1
8Bv5/pFDfGv2ebrAEH7NU8pnchiwg5Em6Iy0JYFrJkO5oQ6rnqvAvgt/Lux5NtSLt8ovFpWoxb79
bknXhdtalXcvpIRio2Oa7NP58iCxSBINyetAzRXU3PM9azQe9QiE1PPyyjM200QcjGt4RpQAcJ1n
6d22VV0GNvhRBIkN2LLAFgRmdiRkn5uU974/aaTDaFOQBLySisEItfPBe70KqtuCJWk+XEsjxdEJ
cnKBKKfrKHBHXwLSfB9RyFbzChe5luagYNOFoSHKp2mkFBfGy2jcm3TsOsRi9RNlqPE0/sEIr7cu
e2zFZEH1UPDdiXCI1BFHKqt6kDTJDtrn/XYX833NupNvEVRRbBFyoxzMHHXiDYd2ZaTTHkKk2gKC
W5s5OFTZg7fcFo369nHg4iRI/G8l0QTiyGMbk1Z6/B7Bszr3vGvRwQUhyXhrxiklOhOzhav3nJ3+
HDT5OsOiTYlmZ8fAOl3szzOssHZZjmulXgtiqScU/PNlmBiI8uc61cO/8fd7vhoq6OxKS2UyOTO2
rytWU3QebcUxrM6qfmXdv47SgKYsyXNXkHk1KtiyAEKFsjRylOveV93BAqUoCekZ8u+DD0IsXMU0
ASmWuMqvs3E9IOko/E1jYb1k8zgZ5zZf0Rr/MtcsWAbp+/PM2Zb86qm0efiP3a0gOgpfgYbPw8Wu
XdurxEE2Z/tBt22Vjc26T1fhF3IaZP7HzGWNmOrGwRTn0Va0gJdTrqYEqZu3q6HS/USJUyCXDs5h
B7pNdrwE0IxEVgsA+qAGFptq4Q+Dii3drnzk6kwBdbjdus/VHwM4en3b6pgAoM6p20OzhwyJDflL
b/hS8w2ApGVcN5VKcn10gSlxgMoUy8KM3Se8+weKArBXkuvaSUI+puopsI8d1SrzxL82S5qZHHX2
MzrhiJ/Kb8LcAwQrjHM6/EsUJkV1aqIb2LaszF6622vycGQ2RDMucjlxASz0qJ4v68XQ/Ue23zBR
t72KKR58u66K3+UQg72XheCgmkszdattOz8e9VmpweKFTYSCeDR1pJl4TTs20A0e+nTuWSxVGxAf
K3OAPkamSMF6Fz3eoO/dwx8DmPHhW3EysTn+pKtLv+92KMwiOYhEspyQgPzY+FFST4sYtZTO3wRj
h/STIcPOb/fstJxMkE8XRh6bIh4/sVIZ1VsRbeIA2DTxZUccrM6EUiG2xYX/GY7whOYz/s3gNPY3
rCtBqHohbPZHiFodU9Qltg97TlNpJ/BC3cr84Q+QQHBwX4vp8PUjrZuE8tOydbLO/uCjcdepTnZF
3BI7ZMfEljPH6uJm9s52kFIhu7xtAYshf+i3CF35+nkyElUQEl2ht9gJ4e3rL9hixn9Ix0Z5GzWT
UFSQXZD7hrvty1s55NprUh0pdPNfYiISmcNJqqjZnhq+CfdGxRbwithKlc6Fvq6TQH1CPCYXjbma
kL8ZQfgUS0ev3UZp4wAip6XPM6Q117R3LANvvCNNwU9NATBpWc1pSww3BHurdE46CRpPMAStTu8x
GWjMrAncRr6CUNegneUqSxJutT73Kx8Ibv3UfStBSGbLRbdlSz7VEQKmEqVJQKw0tR2tnK2X/vEN
ws+55RItZ26y9Gz8gd2XADqxTIM5i6ST3ruJyzWhuMz4Blrrl57Q87T6RPvHhvIHGeCQfnYMqCZN
vz/TlHOurjq0tF5MSOEQpeLKIzVqBg7QVNOwrExVz7mZw44kndoGM8gvaLibShn5RdxFzamyqfw4
6TUqpH+NFA/0Ya/zrz+0/JIv66gjjqiXSrfL3c2hWAlgbMnb7i4mqN/xNJ1CZVjllx4zHlciopcE
zb2EUXez4l+smaJSfg24/r0hCucjxi88QFvo+i80N6Q4/5vlX7LDBERwEoU8/C8KSFdFW0bIdmjX
skTIbRYQGw63LE64gNP+EmISMDVneUDDgAGCCva8xUFGq+IZcNOEU7FpHou/ceTLPADZxSL5qmcE
qbL097ypTfhkISLqa+QQbhaVuYkbW/G/KzzPuoRP8GwJ1/76QY4BHznSCUkaDzVYCaKVUINaYHH4
u/AXVyWA67wBWGzP2HOM92pnGI1B6arrNm6lFm6OhReH89zIy/BvWJYAvJscEQmWtpNqKwKEoMqI
7WeJsYV4mDSkRWvKn0odwCBTZ6Q+VLhGP8j/MuB4+0PUzuNvdEEKa8b3qmeGiLVoYtH6UERbI1bk
dzjQTvuUNvW1/kbZFad3uYCKYu9Cm5tcyiLbasvIvpXwtrx3sq/rluHNbBZlG44VypExtP8a+ird
E7twdX/y/sszd/OrY+5qB0jWMvnGO20VfyrKFP7rkTUDJaiTrUm1pK2Rz8F1mMabfNWlrqRnG8NP
YIMZqAl08h1eOgPbEdI2DQ9O7/mP0uwbJF/X9HbRLSnqg0Rsn/mK3EENO7XqK7kyQQt4iT5Xzbyy
l8KJqppz1Wsklqa9x3F0ISJhFWPzY6C/R9ITU+aItpvQJi0G8bbU3K0BEaOU0kGU5ZLP5e+sIn2K
Lzo+NlTSjG/amtdbN/+vx9vbfdM071y1TM816FQ2tVlGhKeiA5KwIKewfJN4DXDT0qvMpem/VnHR
ljR7mjgr20F3kzBgqGhgJDdvLc8hsJF7vAUbYEefWO6GjIQFC8zM/jRjG6pOpEdxoHZj8txw8TMx
Cz06mAO0v2WwSjeSUz9KReJX3u1Mirmb4wFqS0sSZsmrnpThEGGVoKnLMigFj229OwTg1WIip1fL
QWtSKTn13soWX1r/ST0bikW7fEQEl0bO+NrShePuyKlZqUIn5zX2anWTqFmJnemcEkVHwxglewvW
hY9CaeV9p+dkeMgrvQ156Ppu3m3pwUUpYGW7SzegQ32dGJpdn6WA16oObEAqKECFq3hItvTCY90v
L6i7B6YntTo3560wdvoepOrgg+6RklQXBo9JPpjIGmsJAQimwhB6L6HBSB+gufYh154Fhq1W0m7g
46jkCY1IvqGRCAvTRwqdFV7/P+AdUUtjdbmHkOEYGdx/lS79R4Gtj0oPp0+ShyfD+X5COE6Wm6aj
4YT30p+kAvguhZpkCVP9HUG6tghNqTdObYboRhscM1anIQa0yHgJLjH7u5HnBth9D+nn/RZqJ87Q
0NC3T9y0Hac+PeXDh1x3U+qm1YDBzLAPCK3v/b/0urnMXLaEj309i63yPzTKrKG9G4H+QMulKjFA
9El9v0YR9+duDxZeqUDm1bqyopq8hD4dLJN5ZqAH1WdcrFFeqEVjbA4qIqtvhEnKpfSC5Zbpxdr4
cbN4WdPHmTMJJy7CqtfNwK6AZDz/LZiRx3j2htAjcsRdAuLT9pZO2ubNs5r/XMoDOocAFvyZktJF
3WZC4fMuZarDEJs24uLZz5Pr0/f88iruHW4bb8AoqBVyESKf91aTAWxkWEjS5UKGd+iP8aG1asNv
6PKnm2R1oH8Fj3A6iBxSI2/ekfHkKsTYYm+za0VganmOFOpq7kD72LuOvGDuU4XRGAgbZ1LvkIxj
2J62GFCTuRhZbOZq+qcsbqg/9OlCniuQD5RmgI/UZgrvwln1DXNfIJ0YGSLwHOGqA0hCGWkjtwBO
fI/ISRPBjDmdKat1cawZ7eCt2GMJhFbBaB6EDqIraQ9qQ8TmIO7UmBaQXvYDLKXY5/Gi/UCKp77e
DVtFGS+jA3GX62DZfuwXlXkeazWyT6DINMuZcchBBR35yo4yYyDgz843ixJ49vKexTPTqBYLzLGG
Jcbt+EIPpLEyNd/AC+qwhJ6zjyjlmWRT6oS3/TeBEfOWy1RAex5RJOzQUkfDmhcyWYcjn3xfwtLR
IlqnZzoQEFWJ3aNXoCmM3G1HQSQdAumXXYq4F7QljYdW/FGm9JH+5pJ0ULhcWM9GSq4/kwAHcv2q
HMIh8/2Qstlj8g9fDOFvjiqyagCpQN+nxyL1x8j9RzD+jw6Lm9jKVOa7+yMv9DGpTtMwWHxEBqXk
PavBttYNzgXT0W18pm5GtIPYbVtB50cOkm2dae1c72hmR/sfbiuUsaBV9Q9s6aXJ1zD4zbuUKIYZ
j2PU1mW6oeDC/PCf5xtGz0CarU8Kw6XbDuBVBPxbiUG6+mquV10zpa4rUgzu88crFcRCg+i3E22b
hy1gsZ1rQ2VAn42ii4mE77P6RJ3zOg5g+O6XlSgiokp2Flisfo2/8a7EoOBUFJx1GwJ8AfSanyTg
hYOW8/5SUoTOuR0wLn0wUITXZNiHQ/opPCzPXpHLTsBytbXLmBFuSdzBmcFUQZI5aN3uVFOcOYOp
b1NvGuq8qDJlNSUqiTQGmy+5Hxmf/5+AGrGSJxCftqKmd7xlZ8wqF97QDU2+OzoM8JygEgHW7FTm
JxUHmtPO1P8JItzb619OOLBOlxg6Yr2BrQkO8htJUl+dmV3Ko3JkjQnt4HWLELjf5boCjCF2/E3z
SvNwkOgOqrurL+BCfR4W7wkZy7i9ymbaaUTk6yTNRqqBKyOyLs4KEmmcdYr/gR6KJuvjqJqxipk7
BffxjqT3V4GmNq4GcLZV0s8FNcML2MPVFPhE1Zk9dsrGjXqOlH3r+/4i56uuiJBbAzOwQm3Rh6Aa
c49rw1b2dk7HW0WkH4kgzx6ShL4thzhavI2ZbTms2Iw5erUxNBKs7TcgOSDPguGVvSlsNkgrCUi5
3mIV0IJ8NMytzx7q40zrDCXWVENivMaHJ/OANWpzruDAY4UtT29bKXz+9rcT8crPVx/srwO+SMpe
4JEmJBMF1XOVifWa2MxyBI9md85Q9h76h3TZOAw7jukt1hqJ98QCbi8dKHXR/GNWImWPRRUcmiEz
jGCP2b6FWI9/lAJwMhkozbRhDZT9zHSYXIkiUgGuNm5PK1FltGKXnLOje55VBYaqU7cQ5JlrjEQx
0ITDJA25Yn4+lOPyZVKtIKSzFhxXmvFjkwz2+W4rOANXyvyZzzmvr6wMHqT8RBWrbHjihIo6mYF2
FKo3NuHIJ9xdNxljgcxEDFyTCfWD6+xm84awEPfGT6U/YgdwmEkwAhyAXy1OUIHRgSNaTqoKY2PQ
7bRce0YLaO5LWgT8403UjdaQ+Kx4//4X80bVIHY4Yu9KA1r5aqszPLN1BNBLMYEBAEonW3HGQr5u
glRi9bwyCy1/asvykDxsQix0QUrRAC5kUTUq7QjdwzPSrEMmTW+XDT0Hie2HaUumLqNwHv98PAPy
jdHeHJwBcEzF+RMn7sBEN73a9+eaYVYI6pO8mjkqVB2ckhOY3Tr7CaKpOIqCzrgq/YOi4z97V5me
T80MWUU6jjOhubUwmyCm8Rk/vuMGbvH/Sn8fEd+3EikzgjjaZkuktKEEFeDCbPE/5XovX4q7njgn
7Aq1ooGQXdSD7sajR1YewQSEGexZScHADTkDhOK8Scx2aQ359OxBJbet3UmXTJ9A5lshG0wVTpcy
np1m1UiOc/MMAr4cIYaquGC48h3ypXkA6Bv3KXvmzqvlJxECKnn7zOwH2N1JV3av7+ypRmj6EvHw
dY43YJynW1wOFrTO5xgl4aj75UTC2m74mxesiCoeudAV1J3olEsZFJ54oqP0//u6fNOU9LvYD4mn
eWAGMonuw0od3HmcvuHbhuXMmCTO4+iHQAhaE6e+k5iS24rcnQax8XwhZfhNqgUzV7cu0xZr7lNB
TRU0HNydu9WCq629/RyF7Q3KEpVW5esdZU17QvpoUOrzEWNAKlopBgBfJb7UE55y561jSL2OKPG4
PbLr1gbzpmTNoMSKrXNwuBlLrrgh9+dK6XoIkueV7SdYISDaB4uC55Rsi8g9WW/m3W1h71/wnQi2
qiaZrBtmGE3HwB7Ny9+1+jHkjWr6XZPnEghsVoHKfmCoinVeZzW8MIg55tFcAuVcC1qqqIPhsiJ5
t3bSTZQSIWVdekGDRhUMKacpd0knAeXChZrWKRM5LjdadWa/q6pZE6pnlxscSBW7HOO31jqicLH2
TnhSQgV/+8EwzX4+mXwNX3Ve6JmEGo0IWdhFoBPeEtxv2S7110O/8CwGBTXuJw4hzZ2HtGJncTiF
vap+EVQa0l/rOaAH8W/6LnvB+Np6yhEIxZ8YyMzUMrGNZcNT8DhuajSvT8PkeJXXnRHFQXiUm1Ob
DBiWNe/oLPfBdZXRx6On+JT/2fIU8b6prPf7OJWD5tIWkT53+y24CkmEipTigwBVLO6+rqAPbcaE
oikx8ogOLF8FktclIcEe4f24LxfgnwCWB0YdjLlGdhklBdTjwVMH+FOEtvs2YTaDT1SRWfAZT8I7
Vr7eFqjEXfj8TQtlX2cKuYZOPA6MhVBXQjz7H+I/n8v5niCPvtoS80TnaCliHonzWGBL7JscMthN
Ds5AzQpnVLK+pb9IZA3lPh6Hzd1hFOIX2Sw9+dX2YkEurpKHGCETmwKB47sv8VYA4AQMYbPmcpwj
pnblcvdZ4QOz3DT9lTCfKtAeryuoqfRKjORMZNdR198X8YH+KsN8o0WtcZ1PavrC7Bw+Lpc7B2qy
aJPzET/DZOmCt0HXlm30ZbgReBgmiReIl3NyB/kQYGam9Pub6OCQVmvIM/rFEmRQZpt4LsMLMclI
96iCmyuB86hNboY8dGFyIpUfzywPZZWgBazTkuoxqXmk9c83QjISHFle8HDJDZKrmid+EjMYfANT
lEZjm6AqpZ3Ckf0XNOyeF9Z9TOlo3t5wD05UZMRlH84qIqeCErcCbccrieIIMAES0knvoNB4NDXM
rC8809lGfEJkKwyjqmfBywiHp9vwOkZc2LN/vdUUMuGrBDVVA+ShFRij5eXY91S0wrQuA/N72ClN
qD2zHAUniIG6uzSkkLMMa2Bz9yEqcuMf6fimPGmR4pu3/R1vwbS40NI1AyNBFaAE/RmeiQ4+9h/q
rz2uHboCJT+IXAPk5RlO8SqyL0XIb+9FE0QDzqv/kLZc2hNHkhMG25g8bs3MYFVJox6mP5nkCYM5
/OztZHTEEYLp4B7o0cnBezDl33Dj/fUBd+5CYRRSj1bjcXAwyFuzFtYyEARTl9ZzGtYDq/VOQb8k
H0Fl+jgUkggWTKwb/Bk3DQ7NIzjZG3WULG3GYxD1Td9W7FXaSwAbmBnEG1pHH8xCxDYHEr/TyEZw
VkW0/MNg/d0da/KKRwLabtnpm6UqxZdCIFcZDQP6mMrEUppc2SthGdI2UUqJJ8bXgeZSDjww+PNb
8oIpjCdI227ajNTRU2WRBgR9DmEL3n2+TPEtf4/wz1utzi7vZz/4gpE69hHblD8IZp7da1FS/Q3V
IHVDm4PRXbNXDALaoasjwp9cEupEaAniabxrOUmjgaoCswNPPa1rdZQdraixBNdZHZWequVYN/Jj
YENAXNMxAgJZnQnclNRNrr7b5ipwac8MPIJ/1U0RQ6EOm+Z6WmMPgWnznmQGVlUWC9XKkWt/tvvQ
xW3AZoF4VmwEd5aoUeVRR+JE4grZw38BLUa/6XrbPyN77ugxqYge2IKyrbBXTUCMSgv8Y/zoGqWZ
LifK+KJhC77DXTicn0JMjKwuhb81Ve3zIWKyMj0XVoAgZphuMbcQyOTeTM3DbdaxcMyYmFtgle+/
gPD98MnqVQOEtLyIWEYQ8JtLrrC6vr0kKBEgZG4XNMDMq/GNK0GNnRt3TEEcBWjOBgeHn++1l8Wp
G/PUwN+9UYI/9Q/5FmyUMKlR+mM0ttsI5r6L8Uf2u02I2knss6GJLa7aW3fprW95F0vy0iU0o9Gc
7WZKemnaypxK+ttXNax7sQPdNU3OF+kOjkafIxGMSgBnU5+ktrXKQGxr6Qbgkr3HIrmyhupGUfAy
1dD5ZhTZmaDS4ZYdfHyHUto34lcCaq6k5mG/wVut7yN8yuOFBkkW2/SVKptip+rJfKVHqb94DkGs
TUPWf97Joosj/Li5JeN8YTm9oNUWpA7i7crabQLZoiVX4gt5al18E00CzmvQgS7BY48unjU7SHCO
XoXXrSYFT4nwPkkAyQ7maX6+Bya7q5Uq9faV3T4RoQtXp4/uWNsDpbACEqTLa6HbUPJhqCEHrTJ6
V4SmGiWl/1UADBU3lUxTAFk+JL1JZgAniNmkwpKS8L4u0Z4LsG2Wd7UvD77Yz22Y51bldf24S8pN
2eHr8MM/RUbJrSJVXpl+A2BHuw+9Pc2DHdZe8IgB4my6RNwdaKUBqhlBgzEDWaSid1c5PrDAP24D
C56fppIfOsHX/SkM/DHj0RZ4xtaQBOooym4GrH/Q6BoU7iKUdMH/C0runG+9V8S92wEbMNp7xwtc
pKp2no7r+g2B6FQ5USbcMJBNX+QGBwWYgIOPL7Y+mCogQHCgjmY+gpKnY9VCizPXG633Nath4PYm
5uIa+StARqXOfUkCLfDNWm0l6L9YqaNAnrA5RsX+yxexet5wWLYBoAj9lDMDhvjCDeij8oU6VQGw
TQ/qA+vANsuNSbFvF9o5uxBQimA8vHIKZEVvt7JErRGzmVKANhX4C/sSHbmCq5KtzlFAs7PUWNR/
prYtcVyITEYHa7Ie9qHi/ux4xnbSWm5CiVXyZp42UkmDkF57wIWKrNcJlg7r/jE8SsBzfAptQpw7
Dg11Didp2e8L99anTkC/BzAx4pUxrWuK0TT7exaQv7Y54sSP6NTKeGPHixL4MhKIOMWfFVNjiXmZ
468jTdQBtmg9W7NOhHv77XTycQTPYI/FzM7j16iu3hoMMqhhuQg0tYRPWgjXRi3xv8/jtGWurrMQ
tkAccvvyaDxbaCMXTd5OuRpZ+Z6/4jZtX98hwOecCWWzI+Qg2oPzIaN61wOQ+TFwrjcodJz3owtu
SdUiTfEzkmvG5OUzuYf6gEsATUCYj0IE3/ueAgKOR87iq7pynzat4477j/lakX3gsZjchXPQMxLY
auyQMlyFR5Hiq/Imo1efXbrRI4QurWM95QRLjoYNjXVVBPFyraaZ5v1+vnBBjBYft3/QoFWjs8Qs
TFuWV31fAJnXYmY01jx1k38xVOV6ZHukWIw0HhK7BLCOvoZCIf8APYoYq+Xk9NTLvl7mGpP6ukpJ
k85QqKCou8eB8+wfzN5qt9+MNOKv5G/umkHQ4TOjG6bvs3pndW9AVQ5yVwwAOtUdBD/qMuB52jmZ
eGcwoQzU9Lwq8N9XkX2XVhgicsFXQq0GP+suPAwHxsH2OaHRBcbEYuuQ62bRD4mfhG4iLuc2FIE5
evzzsQSNbKzjWpmRAkynH1V1ggE36ZC4k+9Td4BuqqenjiHK7qbWvblnI54icJVlhAHCIm0MaXlT
w+k9Od8hmnpfFbMjvq6/Wjk+B201pjvk8osQ0OCR2+HdqLlyfy4DVUnHB09mzriFLWgm8cjK8K9w
XerIPINmMoJeKL8bwk0yurQSwaFXwPNkvGM4zUwxWVANWO4qprQ1HyKufKtu9N3639Hnym0RxEiH
w/r3ktNrA84Io4riGSziiDdjv/tfnU4HVQOgJt3CdQQP5fmp9GXSgfJTRzr/TPJ+try5aFy+BQNB
+Cri64TyAs1mNe4ETyXiTMgv+CM9HS8heLS+UdYtxByY9B8c214uK51UBJrWPtrYLyf2qkNw1rJO
Gg6TF0Gyy8ijDQudHqFx9VyuNNpnfi+ECoFutlLQnfFZGSQSv4pDWIjKF3skOBLpFr4XZkrPjsaO
JAg4U8H4snGtPW78wjHN9+i96d6gjGzQDg8fr1VvC2qAeeOW2g4jgSy2zylJnNhnfmujTcHWum1B
ufU2Pnq3bub5jQycDZMVhvGcv11pZUa0ObaMiUQP14dMLKqIwV2UZdjpKjzlhlcdoIpj09tPPvDq
0MFm0Dyml9MoFXCduC0+ycbEhsnwvaHRcIILg6gKNNUQEFNSN0I+q1USp4dFg0pbOhP45J7HZyDd
44jDi7dNamZhgYWTYteSYg9fZatn0R8J5eYyDOFaj+HbTsDBuUTbn1jrHlKOl8MOIn+O1Gtra7MN
mB3YEEseKzykyUjTJuWtK0N/RhH9IaFyoew+fIb8RtSsqu9kH5qrzlPrQT5Fge2gENzqdFm3hUrG
xPezv5kd6fySXb2RC19wEJLSj/DUP6O378PcRXeg2GnugdJEmWkI35NcN96NOeXyzFvdEXX5ps7w
uv0ZLhho6UFrXhhqI/I8jkFKfjt/4gi8m+jtPqZjIJYVtNhY3vPK9ICw6qoxcX7vNuWm4NKLhDtv
Zi3Cj1kspdU7rAoLSqMkqHpUyU4e2Lj33r2bBAKIMIzVi/uiLeQuAxpC4agMsQhEvv6amrCiDjVT
HgpZ+fyhAxh9ipaIV/dW822HSQdCooh2Bjuvzyvz/Y2s51BuFDw1YWKISEyVYRGzIzmGSYz7T0WF
nL9J0DiIc5d9ndZzdiVkGEDd90qAzxENg1dse/oGMgZuD4Dq6wbhV5iqHjjczUOWXn79zPi17LEC
RUkRurd/H9PdlirjnKY31w93V2rySRctggL7lGPUoxQdpkQfwRIpS+FMXhkLhhF5ThYlRvMIbLg+
1RMoqC1p3tyWFJ1sifRKFrR3gXQVwWKMz7QsnR1kiHc/lgvzk6iwNZ5y3EWxIuzBQKdFNsxid1Nj
TJ0DBEBhGZPQQnbzxItw07rOx3StoM2Dy3aVfF6/ajuXpi1BSSbp63EzqPEAICYvEnpi47jImuhu
BpjHqLY+coNINFZaMr9bK44afiuXn/YCgiHLjbeHA1QGur98MvBItN2h/eKOORl9qlR99fx0mh29
x7vXSbod/w8bD4VaRouVU4Buyi9Joob4LO3aDWo7PxxDVTID2wJ65I3FQRuzba7wWhdh2lJRBncy
JyQY+joMCNJgOAmbiDeN6CrRWO1HqmRHFXvIH7WQMk8F89aLZM1ZXZKEYXk8VlX+6Z6qlGM6j7u1
n+FnUWmir/BECWmhCUyqdTDe1IoFegd95HzNXt6zRDmD5eE+41mURw9H3l/UhCv/G4MS73Rw2WZy
DppPz6eIE0Uxk/l39HGnotgQ3s9Ni6HpoCUZuPjV9EBLJP3fBZ965qVkhXMolqPV7pwPZNH1G1i4
N2KCJfFQAdj5fLMGnZEP8SUzEjilr0cpAdraPgm+CS6y9VX9xp2+1tWmIWbxxZLX2fPBaetWL9A/
12Ijl9EayHVzL0izLMtNwHxl48kXI7+CEfzpnd3wZKWfeGGfkevi+jhtLzLxlxhRZ5rtlyHBy7If
W7SvtSWX+NI476iWNCC2nZRCPm3yYk2GTw0fOcI8o3C/nZoUjPMTUy+sOUYd89vzLuSsdZwKp6tX
tpjT08Y+CGrdG2GkptemYfcKUa+SvoG0UHXdR3C+QsS+seS70QbhAvTcrF/uPIkvZ6cMOab5QTLF
lOWoj55LN0xqFvtR9H10ixoqoiyW9m7O33+I4/0I6Zmkuy27VTlfGi9AkmbbgdkC7FNasqPieH3N
/7Lw967ejRJr2dWE1fIDz8dJjQyFhs/jhBChpCYTrWjb9DyswYN+Hb8ZroBztHZqag9qWYC7QH4j
JX/uWiuWW87P/wgrvmkvnLt7r4VHqz/QAzSW+ucOG9QvhzQFo79MUz4/vXpUQTABsOsKt1jP5d9B
vNkFsCx5JbypDaPpOLPSlC4wzi7lXlrr2T2jcV9zouFJcX4wyZD7ch6I9QjRAT/ENg9ymLn0SUfi
mUYyK2ms0DLfMqgyC852rLPiI5/ny/yMRnnL7bb8mlsbb99cYrAUGi/FI2D3wDfI2+qdBdF1XDh8
FSs2WX07v4FlOCmJ8w6syDREowXAGLvrU91u7kcm52iU3MHLNgWzSxi5udk7QUkSVvKhN+CJoKqT
TLHbnwZhK4a67HQ4WiKm0/0vvnOhOR0/snqXR4vRMGo7x3FsL7id5jfuqQDCxPAeKLHUjv20jkqq
q23QmrcdNSWaLeX5aa/4F5gGpCQPM2Kjch1CoiQoFb1OaFHV7IbysZbK2sAG50gqhmQzNX6ylA9/
mE6gIYbRuDYjhPJmzziKPaft0FBfTQe+0gSPyfZTtfsrRPs52R2la4vKbGOFdjy06pUEFgJJjoZT
Pgc3tFIZGUWNXyqCuabi1eUv7cKlCU/evesvyFgiy7ZCBAtgU94IO/j000G1upb3ayWYaPulK5VY
P//b4/soCwhk6t0pWXvzeGbZeIDKeq+L/FxnfMxEXj6HC+bvIa+4qOKAVD5j2LcvMFJUyciDrIZk
25ZE1aFhLGVs2T35bNApnH/Ov4JybMWHet6qcYCC75gOpRYZanPxeoNbhAl70IShl1gy1QFhi8pM
J9930yaG/X8vNGa4iEs7Jgd6ZHV2p8LK3pdguvRMtcsqXXydzvZlP8NaKdgzUgr2QK8gnMMr5ASU
iUBaskOS/CtbgvoOKQ/XwC90bCVYX4J3dwd4t/RLLIHutOWWFk1UJA1Kb6mBdZ6DtwXe9E7aXU90
/Q2CSTFQVum7HvtTI5Dj0RUwFUh2Lz5RZDEOxkAeLe1pzYu7FxFjrl76wU487TMQl7Zm50+1hfQu
sduCbJzQLWa+0y+FdDMl5yyJaaAibOJjwH5xdJVxjIC9vpxIDDEmSq9h4Ox5A5r2TYqrdDgFuEKv
cSYnLXkYrcroC3uWu0R5kW7Q4Xd3L8W4ttYeqwzsRmmKiBu2v/VfP16JdeTHh0vNa7S50jEuA1qH
7Pd5gAKvR4e4kmRu3g2o4NQwIpfX/lxIAnZQ261Y0AtKPMnv5N7i6H1PUjms83Ucmk5ojzJDKPI6
66UBnNWGWIluvZVkDu923VhHBSKm5iW96jSXglLHcOdM0/QelNiIp7c/1vrRyPOQfdua8wz5Zsre
cyzXd++Ll5pcVRgCgCE28DKhcCzTeRFd2F0YOvCR/DRYza57pWrtkTgExVdxHLiBoyGQhJoQWxzR
0Ks9+hENhToPd44aNl8Rb2V0vaewrj0ld9YEgZuW8Ijf80MciUQof4QQnkcC3JkqCch5NXNmzqNM
uNO7pSNZRTIbWO/PJzHffbKiEB5I79ztzOxmW+l9PIMXpQHFM1pWLKtGSm3lKl4CDIVoqlK0PNXa
fQWb+lvZEEWngF83mCTUZcb5qhmG3OY2djU3KUeUQDDP6fU8xiiMzb7d0L5sOHfAF7AfQ6HifDEd
QQXMgfjw09z5TPf9PxFgw68/98nKWDdUDPkdBmDbJZCgy18qHQgenltfe71q7aMzXS0xDQ/cfh6W
60I73oyYHLyevqcTOs6uVu9nNHdKrK+hkVreOIn2W0krRQaverwwksHpT6zbpDF2zbshyrYruKIh
f1tbqvF16K2c78jsUi5j7nJNetAH2d2d5UHTk1/Pjb0ps2l0NyycMmZS433DdulDRouYzeHuJADw
+GZ50mVDO6DXaUtbnI3SQNk0/v9ybvoM93XfE+eztoEBT3zvJkuSZmBg2+/tYlo9aEGVOGWQVwkB
XAsfX5P+EmZe/CEIMNxJEaIevoXUvHspmm1mYJXRmoPiijQIqOr7FmFLVKcT2srTebLUA/G/Kg04
ezNl6k4iGOUF7DVg1oASHq1kZQtA8XtrHuIo4ad2Kmq9VZ5bWOGcIpr5Loyr1MM/8qU/5JD8Xl7f
FSlBLJ1UCYLxLRqeAllvPzM94em4DQfyowra/0fJltSyzm+w8ST5NAoFSzkmHP3kRaxysM5uYYWW
Vmlx9lPm0GT0mB1rXVQH/bOaKQL2ausWL01mieK3euCkk3HQayo4D9QgjpZUvd5WEoJfSsJz4uDh
B6cP94tvTTOorekVuPjKF0UR0n1fRAgbVS9UWYh2SjWtxjWj0qdIBqDGKjbmNXCJfzG7/F44rngf
UdQK7KPchFVxf/nkbKYj4b3jvY1y/LESvsuWsyhYy1kmyFkejIiISmosueaHjmyQKsFiAUmDqVJH
IHpFQYmL3z6dEepVkuKQ1urTQBE/mG4V8n5TJ4DV9DTu9eRc0+3aOvFYdgnR0+5rMsSGk4Mn6F1I
1rQwVPL3TNt0A+A831UQUdfd670JHW9yN98C/wZ3m/V3L+zSXPtI5njvhdxcEO/Rz5qKTeVfBhNT
wH7Z9RrA9yvsTyGYTA4957zmu0WmWaQ8TStxSr7NYzLBQjhTLyO9p9BbNpGS3tCFPIhojt1U4K6X
wvVF4BgJkyw8MgrnzhRlnpwGHXWUwWSB95vO64+U3oDN9x/AN4P42IK2NyNvi5V8XErREcNSBQ1Q
SDXJGjEI5H+32qgH/33j/jkfNL7x6In++kyTwsm/OWR0IS3hJVDb1ieV5S+wHXiBAkRKIc/xakWY
Cfm4dyehCEVDvGBlhGDOAQgFwHuXZMkM7LnNxbCVWtIzTbaeYejo2u1yRRaONb525ih7UHHiO2HN
WRGBYbdGnUDQQWtiNv60FbvxplWrnwyS6SMS+cPZgF6hLCENbr2Os/JvAobbTwzJy2nZFw1zRWYb
pOqb6VJ5+XC5fvmcXBl+nSilpnhMCHqD6PyRAltWccLKgscT5VAgJH/o77k+MIQVNn7BybURqnYp
HmIwH1nwMoZjRHkmJzpMkuM2ha6PyEhwGdwTAorTPrF30aBU2M62lYPTJIO/NqF6MVYAjoGOayBj
cZo6hoVB/+itulRIXBEItRQ5YtJ0qjP6zbtwrW8K5dc6A1mrys1uer5jMHf4APXm/ZNSWA4q7YQg
Su43o4CbIdLMkQYmvI/WqBEUJKRYBF5BDuRRSPZ8YryEr8U8dtcsdJmdP7rt4sshYvx5u9Q7If6y
j/oCcjFBF8HoiQ4D5eLUO5bQhqtoCJmH0D96KvwqKRVCGQ+DKBKsuzIwWXm21Jrg6Jp0EOYStt1P
lwmS9fi5hkdbpi0JjJjYN2SVwZcYLVvuFEvgQdXbK0FZq8RREGjQc2+hpcgNvYikxeyfxWETlK6U
VIOY2n0tDUMXnfvysWT41tkUxghojgFBxlZWCrraUcGZNIzOR72aJinBKuLjYE0Qi5p+QNqgBZNg
XjeM2du7Iia75BOoT+mBGXQNENX173tYYbPce19ykw5zXH+bJlfsbhzjItDvY9DNxrEXBrSoBuxM
YTs8zDxkfVShaKxVkHFuVFijb0FpIlmlVbNx74A1h1g6ey+o8R3UYQcdZsM4Jn6b1jpSxElH0p69
3vYXYyP3tsHC7kYoEwKIiCOpRhTfhe7ItAELDU8hFo8V6NqyX/Fdvms1CEiZ+VimxMm9rbPAIlJ7
zc4au1aDY4OWhzKi6XJ7alKLoymM9RcRZYMiTu44rdtbaCpf4tnMOPti1ERAmJ8z5tiYGhl0wb7E
vKjqth8R60f0QthQ5uQOpe20H0o2EpOYAEjiZ87zlxwewjg7QxgbVT6bYvD2F5kwAGCPvQyRiN5l
MD2lRc9546D037ArY9NnTReukkrv09VkUda2T5N3cRyeiwEyBPw6QFXtq2RdcGsSpC+R16JwLb3H
li6Bsh41bbVagOXxvAiZFDYswzHHNqzUjZ08ElRcT5eCIeI8d59s7ZdnoBBjNb8zMf35VADKVRbs
4L/wjH7EQz2bAVtGmnndiq9RtBpGSHD+uKso7lZ4FAqEwxyeGY6WmulRPQGrnm7nF7roqMWVVZR7
uiRBgBWCQw34Ia1Uo8Ubq0wuZECzdtTSPXwAlp+vjmKw50f0AAjb+CAlvH52niroWptgk9rIXBbm
8fNqPGZkhW6Tqh7rEK9v4HG96UdKWtcjcc6hJvi9Xsw243Kl6yfGadBbFUw566oCGNqcWLZoPaj9
+iS0DwjFZ2nkke0tUpvDrrZcHNXysdPPvll1+2ysqnRqL0vUPThCnELlq8NV91z/ErMaV/DGQiAe
jS1RnXVAVULAAv5vLX09PtVEYo1Y4iCxk9e29EkCG7TTu6WO7YTUfpln91kEdcxepzB7S0Jcgzaq
yiQNQaCF9+UZaIwjNNpjGNclq38JvMT10d0/sfFlUwsnibdHrhqPQgXA61HGy0eyx01F1O3ncbcT
2ayM+6nzuQig8XOCuOe/EMQjWv0y/DX6lXif5pIKxC5jWPORiqXxP4UFGYc0LhZVezbiwAbr92Lk
PmGkwpNyJ7bm+ifVw0kcUR6YOv4q8eiIM3GxKgD7bjkRzDd+SlhmvKw6FmznLcHtbgJNb9MU2ka7
fK0OJMQhCARMPOpFHtwWmnjQQwtt/c1DlW9RidthKBkNPPcUG+XfVxstOPMW7f0gQW+nX2ULwa/t
yEZfPDzxc8XY3/l2e8RUZ/i4aQ6wwIdaHurOq1yyS9ZLX7iaumAd65YfMwUravq4D1W6kZE6qTr7
VEMONk+ALbtq1lfrhRanHDnoJAmJeEMie6oe+3sexSGree9hyvp5ArGSphhssKOGOyTRRn7bFQy9
4nWSZ9PstuOHWvT2xDekZtmUEepKO2VFces7dyPG/lEMYAIrcOVddeoGKvIj/vy7XvR1Jmj14UWb
cU4UrXawBhH64Y9HCJiwzev03jxbNHtglfTSB20ZFmgBHYwXFDzDYDz0CESz/CAukE8m5Hmx8ujl
NkqXmWAnmFSzkKPN3F42ps3y0XSP8L/oT2YJ3ib1ophOu5g+N/h+1fz9OCT+GFOSJEBW/5iC48v0
uk+jWHS3/6x85iWc9qi94HK+QicjAvFsQ293Q5w5TskBRX2Qn5Z40u5iIvUJFyHBcklhex1J38lj
Pu+GDL/2OV+e11aLRYNnOqVlrUWO//FxtFIVTnqmWIqoPxGFXSvngTS0qtrvi40CKWUiRnPqW1eL
aZfCOmNdEHDs7Z7QrKRGDoA6Oj18hlxC5OcIZZYAoIbDrnTc5ga9RVhHiIGGS3Zfp7YEWtio84h1
REHzAnpGze0MlZGy9XTxBkYgYOa+fWdR3NKUjaiGyw+9UTbx8g3t2SO9mc5YGc6+rAw1RrHlC4CU
5Xd8MbTC/7EBiXeSKCbaXzkrNEnLFfbl/3wal+MrypNwcXdZmBTlFfrB7dmD6spCgwMR1KAvX7pV
1PruzToQSyOrimpjhzl3sKcTlI3hLlN0XWZY82Zl7+w8+IStvPPLFcYVednR5Jc2scwK21KwWFYP
3BEFDt0o1LwFr7gtLpk3XPkVIfxcHHvK6EK5hL28Jq6K3O3AUBDFrXZ5V7nqZnoADwFVk+QyyQHh
+WOIeF/BCLWGC0C3eAaKhlLfjRsjE7ggWozuiYKJWJODEB7cLVPak3UcelkMJYeGHtUsbcH/aHcB
5H9tpwazEcwKgRK2bz2/+DmlLutxcLCLUL67I/R3WAGdaZJzZ3pG0M48vVCnhrh7jd8YfClLnO1L
RfP16gJtoiF7BDCI3sMix16YfU+ON0avEIryTQosXbJ+D0NogZK752bHWhCwroIPA7BTkIatjgGo
W1715sKhxjrvGkhQ/TZI9MyYnja4LOHwgd4imh57eW6lsfVAcDDrGRZNMmUlYGjAwGgUbdLyYgao
NZ3uYv3lvO7DTMZkWEUj1U1NbePUk9xkCp8cIz9mNy12iaVmPguzDGFSXC2eA8VuVRIBG8wb8xXK
/BOiqQ5d66D/Dewla3wq0LYrE4vIUXkqIgiotOkaHSIdiQc+x00cFHdb7KlhDjm2Q8E6AKZlYHyz
23VuyYRXhc1kf1pqaRBXFSUXXsYDFVZX9Ir9MCAAiSzljppoeAGBTonRJP3k5IN4O59RcNvNXA8O
+z7t2/KYmaV4uuzVUvN1gpxHP23N0Ftif2dfvNPTQGTAjU9bj53srUViZE3Es8r1IZSgFJbRK8JX
C1CmT46fEiocQZxmyWyCm1f3FkghSBIAu+7HQxkPOVrQoElWDOKNjal8pDwA5fb2K8WLIoKBuWWS
EfJFTV/nZBKVZS3KbuRN13IMHQw73rZeCJwsPsvKWn0ZiPljGgGRoNyaCia89Jp2YKWaZnCqIw4L
Wl8UUYkBjyuOvJftLR60uBHviro11ORfIJGfxHDtjpN++owNUDo8nDdnDu4qhyBwRqk7Xf9QJHRJ
j9sc92cXr35UUZUignLwme9YXY2mX64NmS4Vzk0pJV6dt7BpoTWOYn6RwUOGZ6uESyMtsLT75Tib
vNBZAJSLwssiul8LKq7sVaHP3tINaSfWsUClDmpcsR3RBVWxeM5uhx6nST3NANfk51wpM7eiYfXp
SPAYwonW8nkCmCGyfOlPoCgQ4CUiLpcsRdX9ZA0AGI1VMptw4hMDka7Z3JmOtNrD4kHlpjoQS5aR
P3580ScFhnGseUN43aqp2QhgBcWmIKkG372CJJ9kkJLNwaiFgYEv7rQQvQHikcP00qRNWjCHzaa9
8samFULOwaQRzALLggO0/lUY2CXa0KegWoiJMTdHwHvDihqml6UGHOcUpMKNPNYjuUjianPDe9Vd
iUeddBc9Gl2YhaO32LfZazXLQHybKNQXD2jRDsb7S0gpDerqFfhINM9ux9x+ZO9n38VjjAJqZC5B
yUwosfXJ1YT8+YECrZ+O2E4RIBgTG6PwC+SfFROQ56Ll5R5GGMBUJ2QX680M7g6toBYJ7HMhFL4L
lSyp76jKiniHukjkdSUkXKHgI8sQCrfUgCF1H2KY9sevIQvbmZpDbd8+V5nE1tLnlseheFdJYZsp
Avjesku6I8yW0BNVOLGmZOMgeS66JlmugkM6SWACL2yGIcChpGQ4oAMZoz9cjDpEH8hVPYR1TTxF
rtHwbuZj+1HGTI1AuWIshG4bYIVe457PtN23uLxBn/AEUPbaPoVFbLfMmEqqFGtY/xTXAw/gETRb
dS/f5YbLMkppDhk0ysdJ2NYCzrGrYfkDrICfdk/lBXItt9Oslg3gML5o5aWhtjnNrmmgtmxBcJ8H
4J6CK5p47x1jdR6OVKB8ufNMzrpRsPr/FyeIr4nYHaJark/JBLglOqwQ4tA6PvRtdjNYMDzJICOT
8FztnCkBiTukjVKwo1lXyTR50pnskdwlFG2WDZpFYmuojvlLRtZTI4bpCrUkmEGqZgIwg7TQgOd8
eLgBxyxtegJzgC7pIT6+rdYsbwC7OW5sEJywPcz4y60Eh4NxpH+3UXIT+54sq66KCvKwI9t3UK/5
G8IYP+7NjgrKA7vK2LLYweVc3HRwfWkoBweqGlTdgBGmtJ3kEJrf20074txHRq1Q+REQpdwArxFX
dilhnPvgzIfIGzyM1px/1O0tqqCCo2YPdSt75TLTqBJG9XwAWOCTMVa9WjwquaDcwH5C36Z0PLH2
rFvpkfVbcxMEaYkYECugTRNSPbyH5PL+Q2CCh/hfAaeUbSkqhiCS6RWzMFObgbv9xnbXq8eI0QDX
C2KLUvHhVFs5iStq7w3LLcIZBeKtLFcVIMmNZA8SS3zlGkHqxbvJmaQbbo+8LtQkEhQHjD98S42e
Lk4zefRC13H6hijdzY7Z4uJgQ0BG87i2nhp2yrHqFC8+mBOnzFgzBwKjkkcZ2DpLv4sCz5mw3t7E
bOtnGEAQttLWu67/6vUUuGzjPeyTf3N2g8t3617sIi8AIPOhI/JbC+JcXCaoD+nLkeLn4LqRgYah
D4LvaPoUHA5LhtEKHzZEsTA5cbM1Xape/EBldlTFf65xzkMCy8K2SRrOQ7HyQkNg3gvEa06+R9xV
W5/5qMVa34K5DHiRWRMBx8xQYT9mJeocKpr1vzpUXfQZeGkxd9tciMGQnvc6Z+QDTp44HF1+nxuM
fpn1/YjPJw3yDMgMvUERQlpyg0VXz5mZywgH0l6d4HnEJG2Kw3p3a69YoSeL7VVDEq/SsqE03Hiu
og+Ak8vCSQlOE03pNvVBZQuXZXJ0r7fFM88xxULbvYbzNaA4aLRI+IOmgf6UsJfZHBI7g3IkUbYA
7C8px4UQDA1cjVEFYAUy8q9OPnzc6PW60P/Ix+9V3ztKhIfey4DZt5doAUkadO8xcXJY18PFSTdg
UtgRSA9hfL2RE7DKvpVxXyRvRJlnGZdoFVmo9hbz0eQrK38ShUrhDW4HztDx4ix80f6k03csfdc3
siqdxwVE6XqT9vvKmGMP1t0RS5o8azFKiavqsRWfos/6LB8Wbsnz4Iw+YXpxVMZKAFKx/I4jWr+p
eFeYV4daZHaOoOCXOe7cdPYtE/slQ2yymmACk9MhQClLxaT7lbRjfhV7CjhqqW0aMeTQwR6jp6K5
vYKJA0grmj3DddYu3sdfi6Vf8YZd+itYWQX1BX5oJV2/3gwbASZ1c1gglWuzhApOywSPjIVW5ghT
TfeF6LCUZ+cybiLrVoJkxIbOs/qoC8eUL0ajsSZ+X8p8Ay6lxEcbG/RprodDd+6q9rz222wcpjz0
lq/wSW7c61qWf3u5Y9AaNCckE6isQmqMmuANwXrCia9kQgavqs23Af8m/gdpSKk2/qd/J7iu3gz8
zn2iSIyIzAlf72t0mY4PDEUISizU2VY5Aq/BgEc53D0GLaX+671pQRK76I3HXOPxQ+oAYPBE2VRU
QkrriIv43sQcUBF3+xOQrDHEeQwtp5ze81VqVWfeI1M6fizlGd1TzwrvvEZnOHmPs9SZx1DcKT0J
O6fj93VARcSHencLRQliR45Y9gswEChum6GM7eP68/umGJ2QCllnyAbz/4p4BMbOr+VcIl07++gC
I3JWgl9lChdmKPbec5ybIqL77iPxZlcMiTdNpLROnSri/S3j/lI96qox8atvKipOJOOSw4Lv2jyR
RuzZ2eJv0bkKQ15F69KqHGbOkCLb9Sf2JEi7Ny/H2MtW1YemK0cQeViF06C1dnBcq4O4VoVO5Z7Y
fyATgxcdxeWck8ERhZCWm7JKJLjUOmDOKxgS9+kpRMmXWBof1+vfsL86TmcKuKifEiOpo6w3hEPC
jyKMsVkswJjYtrlTXnG/prGFn3qGKO8Ho8duzeCaO2hg3oI7kEikie2J4mkY/RiNsrkise5DUUWH
6rxJ1lNK/O/2s5n0JNs9o5ZQLtcztBRwO/qgLMBirSc1E9P4+ZXVy+ONd2JsIqXhF5uYs7smx0hz
PnWCx2p/PhfivZea56zZ+qL/MonZeEAfCNLJBFLZNC+Y1PwWQy1pvnI5P6ZWJqnz8qPYqtQIIR7R
HsTIOdfRTBxh8mES3mNoX64lXCOAIj6OivnTCUx/lKE0LTNPdjZar//YYLvKrUCgFSSPvcswD8Gs
FU80PQrryC9wnWe+X+V7eeQMzrLG1gQ44lk9r8yu6Z/zFPYeJ0KPZ7fxKTIL7EQKvhp2/Zcqe3Gi
2R8xMnHb8WYu7L+SJejn58xLEMaaRTlCux+I7qM1YW5hadiRT2DBe7FfNlfUxL40Md4K9ZtO31Mo
ePIC3lSXNtqdCULXZuLG7EIOkdnJLl+G4bU+XDl9Vs/9SvnEm9OG9UpFONcEX/eHiA+BuyoDM54Y
05zpGTkjaIRgmNAY8YZFs1PZwpwgRXbTSHPj4YNX2lxegoZboGSAVaxtN/ybIcWC/x9FS5ILqvC5
+fhqXzPT9En2ntDjj2d1/mIW52C6ClyergQANgrJx4GzGP7prOVrX2rI1MisKxTN58L919dY0jkR
gzH7v7B8KYoyQYnAAdxWdcPqFhfn4pOGJCMEd5JLMZ8zirRA/oKrO6aeRIpHcqnpSmXcz6mqDXtG
xkrVB+aCeu4uA6lz13XvepD52HPAPdXR22o9hcStQ85vqvHMkzWpimY9ouDgwk7JqjTU0jppziLX
+n91kFS1xPMck9AXAHfAq/8f3Q+IYxVSLIkUx92lrnFa99ec+R0z1bm6ivygGQZk47sWp/aYxVjG
ZqZLSqbp12uRmJIUngCQuNcV7BYbpa7Vz0UMciJbs+SMeFgx3qoxxe6hKtguyzx2ItqI8LjQUqaB
a2+PBZ9Jq6JpWnJNbppO0Xu9KnP9zxJFVatax3bYoCgJo48RQSPt7WG7uBERoyt/NWY3L9V9N0NN
u4NhWG1YmIzmnihQH7PiP/Z0Yubqst3oecMIWJelHJtFCRlOk8pZkFq1Sqkrmb3I4AbQb6E4a3z4
wPkiXRlN1jpFL9Tc2PPharayg7RfHVI17DGryb2xhNFOHScckiawAFG3XTAGuKXGPc9j66g4cPBZ
vE8ZPo6SWVEOwIZZWUycJnXx6QquuTRi7bdlAocBR9p43jAtGDGOMiyzs6wEG6qj+R0NQAX7rn2R
VjJu0C2c4kNTbO5eFeInrBLtVgQ2vtf+L/7PfRH4xIpac/56vdRbGWa2gP5ODRfg2opafYyomWXZ
DphniaWWrS145sWOh8rPILURrtp9diPB/G6/KX19gRoqii3K0Ft5R7hPTzDej7EQeOFs0tL27Vja
SE5bFajHZ0k8b/n/516HNm+fU9lJzRnnm2MyWMo0dBq4inZnHC1tCcOe7HFVeovUM7+cJhIXJfNF
90jUthO/hqBo/2LDOtbSf5LX81KTuDqgfyhKKp1dMr5BYw8es9keovz0TIXquL80YslZHs1aJtsf
pmMhpkEmcbS3r7/D1uPLZNi0VxQVJ3em2FnY/guPFbQtZBLnI1J3YH/99I2e6go/jC3wzduh2uGA
6rDgjUWDQncabrfhxm0039xvIxvIStImGfNb0GKXAZ0gbvxCKlm/Cng5X1m8igS3zznaCdG5iTUJ
P6W5J78dGrUtN91PeVTuURvhbVllCuKchIrRvU3RnQmO/h4IjygDbVrnGMhJFUPSshuP+5SbHkFN
lZyKBlk2NcMR3kTT/d91E335hZRAWVBAYa5CsVQgZorAEZll7mwrQnYFC4s+rslN70Gd+U+hNu80
oNVnPMjZ3C5POeZXHN47chiN52C6l7MLgcPPYJTeBFAax1dyFGCOB4JjJVtanaHzdKXpwpebG6r+
3jsyu5iLmbi94K8qZ1xUJwupOOR/MTOI3ry6ICtfbNlm1b7t4PyShiBpeZ+uAEnqrdgfc/05z4rP
KY6mcmH+xX4PiAOoWyBuRwIGZxndTy8kTynM6iwZEawCeEK0TSfeJC4QQSX5H2GBYjA0QSVXze6j
TxF/geFJ7ajokDElF7mGT9hSRiW2ddmkZYlC4+OkpS765Wn2eMh6DYe5/DsceR7BqGcmskvULhjE
5CK2jh6TjYqlFVOlY7pbQ4Ca3/r5I8uJDwQw3k+diahCNxGsMEWUW5Fl2BDx76g11mPSwT41oMuD
w9k66pbtyc6oPdQVkHA8jDRLnv4hW1i2e+YisDHGmj6xbn5osO+ZN5q5AVn4gx/KuI2/rCFhI9pw
yK0brlA470Ys2uZvSB1e5pSb4ZwmE6GvUrQiQk8xOCjvWw/5whAovVdx6ATdeXvR1LzEu2+bB4G3
T5N2athxsJqw1jJMY9vFrRD82cazir9g7WAWKkIDrdhhtke1ereCAEe4alHRhNA2Uc2G53ViYL2M
UuRTu+lQN43oXVDl9jVVULvUIvAPw9FXEjmzZaG4BXJvM+MCSr2TVaRJUzvn/ZYX9iFMIwkUpXIY
Mw98KroMvk7RFjLOQhPWGgD/4H0q/NwKJKRce7a0rirykk9IBn2plf+ZSiMPMW7UzS/rb/j8G4w9
MSsBP6n8EvI2306zG2nhKIY1vAmySj0BEewT61ppTLraR2c2k3xLhHRMsKgzfS91E4wVGiIBs+ie
3XjtHr7xvwcLvJ+L6WGg/zjcNn7rA+w3UcbRqxOHHiwZ2IYSJZ56GJ77/SagWO/tnk5aqwDpbVZN
kFcy3jcZaeBKHk/ECC8hXETKYjz5v+JEdPRb0ILl+PPNM2I/AztEQHGEpC8ICoAdHb6XoUMyBVNQ
o4GVC7T7JgNEr32g81of0mCMLm3oRa5Sj92xudXRM0kB1bhzAxzzPvRJti4WeL86/IrwwbxZtrb4
3NLxou9nXsIbBu7TjKr0M9Us7Xbup6dNkWma3OAWznA8uAxhfZBH2geW8+vpxFmom3fwqw+nJPRp
phTMYCwAtf42Zm/TUtL4DbH7lduHhFfe9p9BAKqfvSfKfKu17BNf6sX2PY1Yr4rxykXtCk01sTYY
FHTCd/qLehmTE7phNrJ+H7AzpVao/1kSQBCvPRlQaYFhDUgiJ2776bDzPVTPA9SjuLCFXI0TMtX4
LszNh5WM7AKybjHmbw6kTqQSVmp1q2wTNJGp61u8gYgBoJUlSF2ATMDdKJ1/geP1dGLVWfrK+mNy
Ea5Ym/rAgl7OIFWqRZWWRJVCbiPk1t/h3iWer0i2f9Yf7lJHoYOoXmEfjgRB8iMdWK7ZkpOXwNap
2kRicmKDqe/jsuxvV54st/7usaz7xqDsJ9sJ29EobF89GJWI07zSX+XM4gWuBFcEq9KSm8gw1Kpu
hFfDdvia5/D5TV+5jXNIGLodhWHh7obP3LlshQxAUrX/lhNgGsrZz3LkhVuHmF9p7Nb+L8sk2D1W
c/NOcTsvnPsnJDzAbNLsanBlJzKSBMK+MOmMQAdSTov28RitOBds3R+eorlXlsrvJIUo/vzc9R3a
VKliWK0YhnlPy4Uq8rrucfmkW7J/qPq+pL56IDAEi/bV/q97hC3HNVODAaQN7CUnnxMpArtJ5dxl
S+euCD1owRwsPVsl/dBggcQRN+lM7chETEXKILSdWBZP3auu7I+5ng8NYDFT5YWc7ywU9iD91CTn
ruE63CfZYCccJe5cm4xmIC10AwUWk88o2g7qwzZIL8/RcQaRfQp4Z1xCbBaBqTct/KLbeZwhsPv8
jG+p/B6OTN2EiZTxiyzy45KkZ4oyUMABj8tj0eWfFGIIPOfLBfJu4K/PDVZZrQN5w5JRLJgP1yoW
3wjkYwALHObwlXR4wk5rRjaxQL4pnelDZvBXesOM4ak73AsMbI389kcfgLESiDriAWSzNqqZOL76
aKGEt/DXxYXzKDznKdM5OzdEqYJu15YGloq3YXNEeLDKhf1oxaLBS+GCyN3rpbgj8QEiUzMKxLBb
XdkYJCCCTZ5B61pANPrnOG+TKRzxbQFab+X0B7YjAr3zVfUezK3AjEGR9fnjZ+a013oIRdDLHR5g
MNySARo7YpQA2DmuT5wgSVCns7JGE7oonIfhbefyU5I5HUTaSiRmpwYs8Y8OMuDx2cd5IyDX8mKS
mXHo2xwvP+iHNuZkALgDxbA6nQ/6CkMsPPe02d1mk1e8K95h2kRDDn3OGQdS3f7OyzvugWv0EREO
1zSOpjSWkSilbpCmtQTS09vI7/0Auan9jWV49B1aE7aavgtoXA/B1IE3DsvrX3n4BvqCQxYU4Thj
Xqlt7jU6LMlr/1/M/w8NLfjMvTtdJP38KIYEfzqWR0fMlvwCH6V4xtvwE8vcXFdoyPS7j22k/p1B
lT0fH/DYw5b6Yn3RTswIbP7MryCp+yuzryE0HBPnlDlAaS48jtGB2XGz+qBwvPX4Ax/ZejkzE8nM
BeUGtg+P8JYNL/dnoO5+TJ6atq/jOEN+QkXe1AdAvdUcGS/BWxl5QfIPQ7jrcI0dDZULU6LbOIJx
+blUnHZIT9vWNDfxz/ABx/ktgCsVq1216v/XORzc0G51YMc1iAQ9kLbFEUDRMOdXfT2PULiyXfzh
4vBzxse54qsL986zczZWdmeo6BFwNPg/AbYUKjY5e0FHhXTrmoPeDgzNtC3zYShbSkCDB38f3GyW
uyWHa9FUt/NnjnRmB7IHW9JKjgz4rerkFI9Obytb5Hmwg5zkBG5/MiVNnm1UGY6pXr9idRPFYen5
tuMHCFi5UJIe0Ov4Ve8BEdtsJFScgrCiV7yPXGG1F7CDJoM6wLbssPBM0Joai4E4u3XZsLPlVbu9
szDsanEqfz9P0jvbe5+nUEoV3gELhp1DEHPX+OKKNzi/lgyh9clHmQ6X0ulGXwbZReXabHRLz4Ma
hSwcKrDfWYsj920Nn0rBB3wmMw2xKCr39rP51H38Vcj3S0BF/SP16E3mSr62S0SiHrKXPw5LzFVK
6lzGag1hLJE/gp/YArDf29+jBkGRmL8BiXfgQoRUhFWJ7lR67bauXLMCPberRCNbKWP4um+idV79
dlx2QNmQ2Yx8fGnMW5yv6qGu+nDOGTa6H3WXBGLeccRRWU8mvBFuqVmfz/ljMKHCP4+bTJFG5NPo
6ppgj1XMf4TRnQkEWI87TkC89AO40iPMKScfNZ2UXP6Ku3/LQpoU8/xsdymZlu7oPaz7KM23OFqJ
Xaixs4+SW2+kguFUGNx+LxjBjnBgxss99u9eN/J0elGtA3rCgv6s8b6ZXTtnRz5rIOvxKuw8iBhf
g6O7vaS71fgnvPQtzXvyMjOdPVLtb65QrmTRcr/jWTNmpap5WdB14EWLeksDozXtmNJMxY8C6QdS
YXp7gaICcbsWLItK/VLlavOEiAyaaX/UogHST33JY1mTLeyiakaSCkz7wOuXbiMTDjD9u1Nk7ZdP
J7HOQ5Ttig9rcCT7XxfWPXt9o7KUxUJyy8fAcHc49LK1vlvYUPa/LbyV3XUZMUCzOWoWzA/ULies
1N/kImQoAZfG6sVch9eAxQ1eEpLGADbXgVOUC3Mj9WaprGbatysKosBseTqZG6w4jb2LmFu87Ydk
L69yB+LtPxxbgbDeGp9+X6DdZxULLer4M6B61qtBAfipVTNc4sjInwoRh9HbpnHT3AA5ask6nMXP
MV9EHkx9SoMebp+DlDnpoGC4KzT+aJYd1OmoxakOmXC5ybfP5goVVF69M4zp0p6PUxJdZDOAcsPN
DtUftz1Aj5fCjLtLoXkdVK0QRz6iauczROlpDjF/yzT4LnezEY8lsfGKUtE5QEK+M166T++7yEBU
Snydp/flD4YtoXFNhNHi/F7fthDPH/JbnV0M11C9C7tyGE21JGPdhU4wyVfDYgwWY2XnQgICjlhH
Zzo/C6HzucyKbVrJajV4xm3SbLcSqzDXSeza16XbUXIukoybO9Na0+LXvPN+hV+/F5GeDMEJbh2a
9NbkP6RYGndV89zpEBeLaUJN+f/WRmgvMjjp4wfhkKqI9ma9S0YBXP0ftudkSbuguAHU65WTSIbW
/j1ywT3UjD164q3zfkoERnHoD3OlqQvDCw/nKMHWjLhOo/5/xawG9/QlvI0NaduJzMNGYUhPDIvK
if/uddYSL7VXNUDKmywTqda3LhmvkTx8tZniY2dNayp2Em9cPEfWxfa5Kf73JsOOkL7pKQNwRX6Q
J4002aGvBPRsvsX+mssd6MZDClGzLau3sUpFjySVgrfYpQjSPRV8XUbxRurh/6OXfnMyoocA+dPL
n1yzI888bUQiv7H60EBqBlwuVjJQV9SAfc55JCe2G3JIS5PSORB10RM6wPyPK4h+07E64gGbxCRe
r3dG1VDueYf2E0FanSA1GC65/KWqtp+Jfm6GW9yN4iUMm1mbBN+dwWPaBPSox9NrHQE9AAzXqv69
hox+5ZwuMpRs4uGJ8UACBRaIKweK7lMhTL3NOul7AbK1h/Qa/076pLKgNDr0YgeDfzA+2DWuJtPp
kR2tuEgiT2ChDE3wmKEi1g14ThtSvX87CY4KlXhnMgI8yOTWYzXE3X5WFnqPDypJNp6vE0iPg2+g
LEJxBG1GiHCJ9HG5S7uQBHUhpltEZJ8Net/Qamhh/xk+kYbVmGygN/29soo4Hi/lVH929Pye8BBq
V+hn6eV3lcXe0JsKyPCiwL7f72xqfCTBqBb5o9mkLjmu1CgO7JgV5Q3A5CdSLIcAfnlBClX3MjBz
iOuDHO2GU7Zv2aoBGMldhBIBUPqazUwGYLlgi+36RCM5wQOrXCTXVKhQbfzUSSF7tDkYYhK53IGn
FDNGJPmXXzT5B406zQUjwqg01SGStG6ho0I5x/37esJQcQgLe5NzA1FW6jRnkHZFO2B3WJKHvZ4G
gpjL+T3VVTXmS5xaz5Pnu4MaWKCvCwI660NvbBvBZGF9ARC141c36NuMhbIcV0MSxVdh7CzoBLgp
QrnZJHII8Mzyhu7cSQUft55wHqQqYbgkaIBGct/+kvvQCk8Pppw9GdTNtZAphvZcbGpUfKiJsSDg
iTB6RHQ3fk5yHakZ9NbMbP38AZo1ypcZwo+HhqBcHa3XEX26jjOC9Oj+/YzmEui8yaV+5z8vY+JJ
a3CNH2hyC/27einqZNqgrpazu+R2NJ0Zex4674ooTTyY/shWvM7TemCBXilHbU2IzTnWHVM9unGG
5zNrgDF0Ky3h/c1Il7d2SRNsNhitdtqA4Z71wx8UKMZmj7y36fF8nz0YQm3UtedGB78PMZt0/opV
9O6UbM5YdpENjj8MISpzZ6KGq7YEHDPBEiKJmEckCKD0Ro/5ri9rYCxWFI7x5+9PC347IOSI3Ar9
2xCuvV1BJn3dtlHL/CbQgFXkzEJh8Vtb0c7TDZd1xSzvFaDDrLiRwOUOZhdKDyUgq/piHbYny2sN
kr7sa82p8nqiRbKVSppSidRjJfmbKpUet9vcJouJTXe+HgObNghCbIgWmlj2y8JpcPC487tTPs7G
Ze0oZPbsT1Aa+aG78fAXZxSIdPZMw22kzBwaiHEU+wBI9AZ3aiwp6kQ0e85m9APMO0sYOCSr+WRO
tJ6aVKZJM/ttmdx1YScPcudt8AfzWUIAJe+TlnmoK21EuBzt8iAK9almpgy6V2+35onBkGaDXt/0
M0z5OFEO9u4FK/bZtlFPdETbxGvkBbzmzABqhHzGn2k4t9HU4t3JlnhxKOnu4ozLnxa6v30WOcHU
lYfWtlHBc32lHdyCduaxdG+7ct7nfxBC+Va7YzpJb8Wh4513gdeNkPWPoPDvdgemRvIgcUiWgG7U
+hLffzkYZPCXnsfr+Rdd5bOT0nwECJGMDuOrx1PrlHoLa3yEy6yGRUGTzb3q+SQe0k8BKxizCCd7
U7pjE1esOydXeW0mFnEzrJe16gUfdfDYLFAtIlt3NXo0vxeiD9WMSW1sIgX/PKMW6qn3ZAy++v0w
1woTluNDheHJNRCZjNy6bcRvmxGm+UdQ50+rWphVfMAYPj5cRt9U6f8OzKrgqhRNdUlxemyh0oBu
l08txhOXq/CW0tRvxSoh4jHZiFSG+BFefrTtZzhQCNyCV4r9aP1ReKBv2f3IYq367LJbVDw9YsKw
D6EcLGv/XXDYptZzIRotAtnxfhbwsnXz85YsX7+Odo2ek0MeiBGUa2LHG+uMsoaEh2HoanzNjW0N
WLTjh4RthFrpP5fo6dAcue03dXAprkrFP86vXIvlESG7vZ+2UqlYUFqd5pUo0V/Gh4EkwUcBX1p3
5QKpl3BwmY69UjTJl1Q9wyR4Ij6+UAw6a6mQwCr0uY5ue6sF3+ZC85b77navFsalmcv8QTefU8HI
QE8Gb644OfZuT1y9+PokXiefHShS+broQbuBZItw/s7hIDrhtUWbnSpXgweTa0REE9ecSXyLrjL+
VMBePPjYRJ6uYHiX3zyBHmYkBqYuyxvqZzH31mn4zLBouRNkIA+4unrYejE5GVw0GEb+72dhIN0y
8s/fQ8XPLtwdjLI5cVs5xB4AFgb/xMzQzMP0p6/iMi2hebBxAsRxXg79ct/WIv4OEWo9UWle2oCL
4AfghFoVR8kSkdrRE3kofDPvtLV2kROPScNAzQgNI/wnEB0kZ85JFAbe4xTQplc/fswQn8GPuuCQ
jqziINRcP1TBnnBFoWPRiXsg/lhKwVvC65r2n7bxLYU6e8oSFFGq09wGFiTKrTW/Rdh2UK/dkaWi
aWG/trLtj/YITKNPiI7PNnem1IKFrrBmyod9WWY6sjI3x4/VTPsSPJaeejE4RiUTXDcdd/KRKw/U
k3H5+JVfkpmLVY9IlUZZOBem0S3h+OfjiATP1S8lX8ENeSX4zPAt/AVeKLKe0SG2zFLayzpS+Vor
v7QHDpKecukSXC89tzyP1IYe//nsGwGdG/2mDiEoCFSvnJTwbt7Kz0wc8DxdaaV2rwKWzfr6+QC1
5RGpUoQ2xXRjRtQ9ZNqTCyzMXv7Sv/cGqGQxZe579/SbirEKIDIXmgeOtOA5zi/nlMSlHtOv0PUQ
GhILuECG/6gsq6CBDDI3GqbWgkAfD+BbUyCJ0qjIVg6jloVM+hRByjCOO28Q3/feOzF13etXSG7t
Wr0gtYhmiy/2VKe5UTncHMSPTRivIFst7Hx5St+26FCKWWj2O3Y59enYV+iVPhZbMmlNzWc3uI9j
yU3wLMnJqs47GGqV4Xrn3E9s4EfAUbYZHBeb/a+6NM2U3ZHNxqY18GpS7sNVa8E9LqklJ0Fx3Cro
wpzw6lqexPUyY60gllgLELd4qxrsVq/CyR7u//sFJZIQor+TFrhg0IOHkrx/hBIMv/nzaLYTJwaJ
TvMxiBOSvY89ba5QK3xlmiXd5SHBUzTnHVY7e+PMgAtuzujFsSRznkE3KMrWkTkqdJkXmnMFyUf4
S088jNpZcUEHNKoO+By9PNiOJYyoMGKEQQpiNfznYhHBbsov+QF0h7ViOQKhmWuH9g3ZKXhBTEO6
/jFJtWeigQN8DaI7VHcIgCbPxjAijcvpLpTITtAf0u/wyGaRVN451Se1JJANTVez2aIVcglf3qT+
wTMBYojMBbWk8pG5QMPyqTK6qoMXqg+IkOp40sHRo+9/USwwsWdJ9gpd/FXNAqfFOYlGXEfq9hPn
xQBCST8bHub3VA8xrSJE1b0gLZGrVPEdqTDSJ6hKKZWQYx6X1XOxcZD4rb62An253P+e6MN9W9qF
Em8NqujIIRaWvpLaA7Ks7hsUNZD3puC02KrbF/Yh0oG/TAfuZSwsp2lPA3ZLLJJPHMyM7k7BnxG3
az2o5s49/rbbuSi/ItHuw/RjpDLwnIhwCcg3dnGzwNMDeFc/oucBwEZvWu5Y2TZ6fL8fDb1IwLoI
KWELLRszzUXsPJbNMpeKeIGqkREXN1AzVPc/ygrfm7yc7oLK6+H/Qq39Rac60lw5w4jvheyOWbEO
v3u84KSt6KdwHDwkwCbitBMxEVZHeDA+hxFsmrJVUw8cpICWdoxi51dhG5Az0msbRAyHhkL9XPDI
9qpsxJJIQkuvroxDcPNMYx/BTc31DkX1IzzxSFiZwTypaxCgbWseoeGHnaTx29WKHpZQFjgqYCGX
UIFh8v/YQuGletvi4qf/qbKqf3NR41+yPNT3RCuWq4p69U6ZJeBQLoMCxWMZgLGmfH92EoiUMDNF
L0/PD10/fMt7XJaPB/48g9VbmJREkNcUvzybWEGABBv8KbZQnk4DA38ag5VvrCAm9BV8DZGcUhnF
olHQtt8w66ZBvWMrsd6tmzTeS8wx9l7YlHYdXPSLoPRkyfO4ABAI/dDCagC8ZlJn+iQeYL2Q/nK2
sfXKCvTs6L7m9ggTwOSuTJVLiviF4QKAc/W/Z1GzaPwSyyT0imKOqVGX2cOQIbZ/OjF12wiuOQgW
DifS95x9TuvrFw5MyQGQhykRnh7YR6kJ0EUlnn1oveAH1r3btuN91GdGQXH885W/EhQYXdcVtXs+
Yuxd9NYbkb2iAOSPqjTDNPipeGOCjTZPxR5nOJZQWhwh1BwaK+1Ji/1xzQh7tbOfFIJstPxAeA2q
IZhFr9pTPGIRAF6RNPNbA8LvXyLk8tm7/RtsGprecDTERvzEPfTCzjpxz2ExvTUNuZKrdEHNZR6n
ou8bpvye0jw0Jf3LnYLgWpCYy299t2wKp9GiajzO8kndblIj6GbHK+TslwyVAvnU/dps8sG8WwBv
tkTykHZS4CbwalBd50OxEomvZqRU89iJB8VifSFNtTAoqH9G3Sd4Ge/HJU+D9YgkvDNLO58ZTBlv
sCWuGZiAK8LVdGbzvdYTYPQ4mUtnpRtEWKie0fTW12cG+W0uZ46+UqPYl2kBm3pCRECUZctELFKT
dPNVuY/MSm8gXNVa95BcR+1j0/GPPMDNgTQsW3GOKimrU6HR4ecZOqxCtQF2VFShhxytkRH23Gf8
LZVU8Hs9+jsx67fcs8Srh+/WRrG6DSUGoPashhYYRJ2PQyGKLoZfb5gjDq8USj3RYdoHv+qR2LEY
b972d6WlLdeJ6Bf2PTlC9evfpHVvHJAA/upd7Cy7gsnrI82Cg6GKEkwkbwKA2t4OVCkY4zCcm7yV
1JiHuFGsmX5F7QDG0w8xSvguAnYY05bE02ILCN+GlU1lKVd1ZKPZu5a1v91asNp5+/1Q3fUZuNbT
pTzQQpKM+IavwXRJTQXFRjNuyfru4hbuaJcUHBGgSxLaHkYnGcXy/bh+quligsesQhxvRSXIFC3q
gkbjRbSUJBKbGaYkwdxB0flzGQUaEMP4Q54HN27QpBpQIuTHCsJGt7H8eevBtI0Scaj1o4dV+7za
RLUnMXdg1aHI90XmdAAmh4IWCLpmg8IRgseJTxJLRcQa7OjpfxeQdQZy5+zlQ5m6qAima8fteyzD
GRpKfhFagMxMaOuwjlNVZhGpllnYTLjKeLzNiFFtOEkh9/mtlbjSrkUc3q/sUDm6H8BN/95wpm/3
ubsetfOM6ML1KhqwXhMDjIwUw+GRxRtF0FMG5e1Cs6h6uTuSO1Wr9HU66E7ipR+EZR7CVyRnSscf
D11RVvEtUsjrYepa+OzZFHruG9rfjjvzXvmWeXxPe9Jkq1LQeDfRe2e8f6Yduynx+sGGNMUWzE9v
cXG72M3apRZvJ3RwftCA1wWU1VKJmhuHc56ks6Do/DYbx9ZWYr481rBGvwFAQUP/HcEaIxHMCynD
ThHe1rGgdi3kdL9f6PBA5cV12eYtpk/ZDjxpsOvoJQaxgfFayLZGkkr6/t6Ablz57onjQ77T7/J/
pqA9ExfQ6+Mtk4gtybyuBGs+B3AmVwYEMCSk4x4gYGcTKd0pkZ64QXQV7bDhyuH+PXEi45C6ihGW
dwdNmropwxWQnN0LQmaeku6roei6ShJFjalAp/l+NPoQI150Mea5dhLTl9JF8fHd78a02YXlsciS
24qIms0HvoOG+55+WHOLP94LQbWNtmnEt7xbmiK1Sr7cRabMxinf1iWXVljVPReSBHa9Q/lsIMQN
YK4trmF2JbA/tHq3KiTZiMD91epHv11NexD8C19EkewmICfWwCdBdt7W+ouCF2tMz9ebf5Q9BbHV
LsqgsMOqhaTGqIUf8OQEmoUnu3V8eVz4ragsbopd3twW5IuVakHNeL11WhXBw+EOYdRuCDdNhWFn
RrIcJbynX9bcMSjPufAojZ5OP06eP3l+4tz66v4+MJrzvsw6frSvUvbdD8/ekLxN818JzUDxU4Aj
M4VgyZL9LosJe0T5d1jhZMP4FBWiHtOmPHFiSPMSvF/8TRE4f3dexTHrcrNAck8pExLbeJ4OdcxW
/uzIL60w16iqbWIIFl/1o7YsrRPhNpehelnK8x38asjPFquHAB9UuuULJxYxWXwgGmFVabRGm92/
CoKVhNyihgr72YxrRLpLibaAaFN5EpzqFnRlhtnC764M1rcc7Pl9nzJ/Q85yIlB6bCe2gT7h2sWs
xGZLjCCWpJLkxtjbAL3CJAbOULf5kRMWebHIveCFPG2DDt8wsVLKUgCEnqwEWQ5jtm+SV67XdD2J
dmasV9rF7SSGonYTydMADyD6StVfItKUKQxnlapWb36FJ5xxr89hnUjTe3+I3QuPPYGXD12bllsp
KM7WdeFPCqEzxawkIzWjeC3245TPCEkd2hhifbVCDmEowyUgpLxyTozyk2HwrUrb/c8ufx8FPnNu
z2H46s8iSW8MWTRDfiKdZZdiw0YmAkdcFvBlenvlZ335Tv6NBbpObOfeDxfHQr31TKpB2nPtm1gh
a91t1uzC3ts+/jHaj6bXUg2d5ROAMvJIg3KwoAhWGxCkcQf8mPzqxlN1F7r+s4Op+aw0iQIEoqir
JxjskClG8/RzWxY2ZqafVxQC1W8Z0zBIF2aYrOvOVBHMYS6hPDOenXaLyOzqpv7tvvQDypOJlLfe
JJjSrYG4XENpb4gC6farA0ChEwF/m99NsyWOAr/zSHwFfbDD69HHACysUuGhyWDQpQvhKxLj20Xb
4X7xWgl67xesn+OEs4rByOOE5hvLCpBAKfXSGO41HRkNpnIAGaqZKtzT4JCYrXWsXrk91MGokP+7
eZ9ND9oOrzmdBuJuJ7f8mtFRTy1JQU0XwBWrqj8X2vj8lCA3mWqPhvqAift2scfaN3J1VZ09tCPy
qSx39/Ct5vSpqtPT1vVoqUNOXlhJcUVYoQNmwDv3uGAVznbikCL21ixli4mlJo1Qm+5JLviG6qYb
PDe4LrmHfDsPitLo3d6qvcHJGYszkJSFep+e5hRPR6mTNKFbqfX0hSfNkerYo8iv7FHL5/sihcLQ
OnU1GH4fHy/PtI3Gu5LIDKKf57HM+LlV6YnQwo7fOnHcARYYYdRfyfrFu/BA6azUU4+BSQLmr52o
JfEVZaGEh1hoRs7+1Ss8OsJqfihK/tLoGoI+6Wb5Ohm5xJQqxmIrWVOC6kT/pVv8xnBT+BuhvUEH
/ggjatpOTjFLIa1twxZF9LYYi8mgP1Oc45WYhDrXayheSndz5OI6TBL5+WxoRpf7a1JX4jfBG+QM
DpJwcLsXOhj/EKDL7McacY85ZdYqT3X9BwHFK9tjn6JoFO9k0nrzt8VILsM8tcr9gThJTc0CAAWp
Y9c3EodUhcVlImT8AsfvqthvwbYlWGwKEpWjCf2dvcxu9PVSMoVXDSjQllR9e4mb3h9+0LrftZaO
6yNfn9NVJC5xe3mFdbNQy24bE5ZRzeu6g8l7I668uK5Zs47/ppRgXfKveyLgi/s6RTkZcMPwDXLC
H3yYVpN/EqiQHz+W6p3+Chn3wJYl/t0+NwKe6+NvCwjcU9DG5wnBYo2vm5NTniTBpuxQOQIsJ0ao
52diWnZuYd60B5r7VWUknh36AabAzZin+/xfpTnALVrihnGwiTNrUTExVvH85fMr7dwrEw/+NNT9
DpTNRKpuwlMJGWCLvU++ouPPBpPWFQm/O8i6BrceDP/evOc5BmG0Yu1w5tCLgQPxo4Mt24xhKWK8
luSTCY3pvLdiFtxbdpEULwAi8INpUTOVAfI3qwEMbvHY39XcnBwsNpt83CcWQ3rA94pqZ8XWWIpH
ezpcNYutYImcLeclfNoUbh/zrdDjcbTmUkKw0DH7qHmXW2Ri9iOplB3k2VfK9G3+SU4YixyJXfkp
3UpAzfyVswhFETaRJv9rXuVJ/NonTXSHLe8FhwP3K+lMw5TgWmqL8Rkc7YnsSfxc4GV6Rov4Irqd
57MZ7bDDBScYd8fwxMXjaL4Wur9SvLtiH9Cn3M6VrwoogLNKa8ZeQgR3svR2xGO9AiqT/6/duOsk
r8EbzfAqbJQeTBL9X61PfMFT8ne5DdaPjBxgs1nlD8ekfTAwD/A3pv9GGp9HExJJkYPw2xnL+jRG
ZivcrYyDDqmOBxIN2y/VfeT86nQxvm5cyC1YbIx78z5m1caO5dGefMKhIx/hCTD0J1upanVKRJYl
0JsQJ/oS40WQXQeidsbq0KIgprJ7db8EWsYTa/BHnx5gvseCmmQQRn4SW+G48oY8CYbpLpbu/g6Y
IztYVilyY3pBnW2+1qVWL24O0Wl3pCy4XkYoMwfFLkgmq5YY/sr+YW1IOw0BR7gw6ElRASuyLURV
hOGK/n1JITaXyH2vR9a1KGNb3j1yxnuxrz5JJ0wKotMM2inWh3X0Km20QHUJUv7UtRSHhHiTPIub
VA8E1G8T/Dis8ga/nJmrOGMrudbD5C7lwnF8WS/1qOo/p6WaoYLLC0YwozVRkRSy1rJU02229VYr
HzjGNFiCY4G4M7piQ72h+iwJiqr0ZvSIVyyOQo3aqRuUW6FXEZ5ehvxn3wu7K6mQ5ABIyM5r+VMY
y54zHQsMRFEcFGTrE5dAuOXtnhvY89c6Yztv+ZW1Yp1LG1HJjx/fkr+uzY62r7d9633cDxDk5IwJ
EyXJD3hCG1AuQF9DO8RIvAB3LPteCpX3av6KtZ97JfeK8osa0OfHXLpFAZFZcgGhpAYetRwaaqDp
xTw6/TFt8hYjzFvxDFhZEKe59z++ysQmiS48NiH8S5Q6YTBconipP7lqBSVEMHmsgyhcLEL0MyFy
hYNCm+78+ZjzTBhqo4WnjQ00dO2Z6MOlAHUP/bAoX5TNLoRvfDoreDlyLSjFkwUhFjnoApnl52Xb
NREVporYRhT2TNeCQ66UerEUzsnkGMUUHmQo/f48ecH4h4HTDXMYid84tV9FCnatjuJ7W9fAr5mq
B+d1Zl+NnStfBFYqOTv73L2ij71GItT8RLPR2tXXtvF9mtcZhJ2J9Z/mB6QNGCmddMdYgNijp5bF
L/8vwXTgvHtTCxnnsAy/8AyA7YnMIa0GWEnx9DHqPe/kiOiofO2gaKnRUxupGL4hTPG9VmOEXaQZ
xaskIwu5iJUtbNdFUAvpGDipyabB2A9UltEZcXJ4KMLn1YTluO+l7KsU0PXHw47dYYzKCf8rCYI9
qqruXX+JKCQuGeLtmfPOdi/vyYSkMjV9O5wbUY3m8TxSdwRn4L9LhQvzQ+/XjUk5FoAyQvuUtrl8
kE/SGUxHt64Ja4dKtiZ5ua7PRtSQmVKR5DYDooNocrFQApR0TCH4TGuz5ShLQkLCH/rUmIhWMfxH
U3KOHcggkSUhByCTC55uOpSqGpQfExOG5fTqyYrz6jmM7eO5DFn7Ix6ZmFrzLV9hvpcbK0oJBtNs
bkDwPoqMDDXifRh8EiR+aEZLwIHteWSpbmPcmCKDj+5OOWKQYrr5Dg1Qzv5EK9mnljZvDLO0oGES
u1x5eLWCcCFvaeNhfsqm/0dkmlf2UUBdl3Pz+XvVenTFkExvFCrTFFoGt3RgFTsXrNJ9C285fZ00
t77j02Lu5WWaOyFqQNfCcrLtTEAWKqzG1b+0LIF0f8HUrYG4eOB/C+rnQkQ0APB21At6/bqx+rTf
grkvqoIkMywSx6Gm61DigUeI7ilVUy26YYbmaXU7ljvlo72/lBJpl5NBLbHBqwrmIBXcJYP6isfn
/k8Bpc5omA7RCxogJmfyoQHlcS5vno9D7tCh/13sLATwP+b+EletozTgs3Wn2y855ixWeTEZcI3w
FFEZ5PJ/GlaCeJmQpcB3VVGnZfnMh/Rn+y3pwp3E6SOZZUrpE6zx2C+gyUJwFx1jyPNptZEe6Ai7
loMA0dC2LhzcD/DTjl60h4nsrrixgE866LPvtj8E8YR8enEI9TCcF49sFvvTWLXFn1r1/n5oSQ9P
YYuTayd84JA7+O23EtLaeU2WQIytz7EqOAfB3RJFai0+M1ySlp8o09ZbbsBA6vKsHM1ygFscj52W
FZSnzM/bChRD4UWbU/sxujEbqxr+BL5jGybwYJyAZjt0hDRtWem0I05V8l9JkBHOstSm+PESE2y4
7qVYtbUdD+glEwYleQgqZD/jgwqGQDtOpbzZfICZj0mEPGmRCoKCWkoTV8LnNppRwIG52097LpMc
LKf+029omM1YcZjhoXH6EHvgpW0KFJfQSRhMADjhLnOl8vYOTbSo/GrSyRTvMBqTJrmKA4tAZlsc
QDBIhwVLEkS6t0Asv6/6lvt9Zqg2Se1Zibz6Y4YcFBdLIvDX9KwZNn+g7Mm1FNlyzDLu/2EU0jej
JcJK1u0cf5Sv5JqHWe/NeLT1bQcqRCK9H4WAFv0s95/MFklvEJtvM3SUOsI4K9hxW/cLhbcCKg7q
NERS+pEBPQzCHdFTxmFtJvOqq+8BHR7prY/rGRklB9NEVbePwPgDmCdRNL0sfMBRJPnmVa67WN7L
AjJyDef1nHlNNAvO5L18hHnKBiVMMd24yA63UBqdkG4Gd7kvLWDYg4YPgXnkn/dv4lWUIdYunEjs
rZdSKjiUMBFjyarQqazl2OT3XkfjMVX0L0WW02ncflPBvgjeybtPCyQ4y3J43zlWSRgOwTX6w/M4
8IJ6IPJhrF24BG1JG52BlgcWV3wez0NeEj3AyMYFbn1ecFv1ZFMC2votZ9IL1kQn4lJcEqrfoBQC
ALQBg4UZauv7cHOZ6pM1h5t2TOFQsUV+kmBf0ihyavcVZaqrG4p+J9ZAYP0W+cnFM83w1dRgmgxz
rVB3YeXqGomsq3otdbT4+G9eOKpBHEIjnizJBzum2YEIFdNZQtBvctPa04bQ+0tO7T7y8X2vym/Y
HM49+UBRyZFE1y6mTDvi4WOm/baN/Jf/LmYkDN4umXDVhVFD7rtZFOi4fbl0c4f9l5oFOPRqVJqA
jFQ9RJJ64uJey95g3XhARJ6aiMWXHzXFqtZgAVsqVeBKNX8hlHdTb6ffhps6RKUwjF1e6Gy/KfpJ
Iy2yDzDRNnykFc4xMvflGJdduV6Rdlgey5cdaZkhrWjUNYo1Fn/XwZXbs0eqOg/tLgKgFaslIn7T
sgLPgZmV/KxdZhKlsiUJxdqX8CDuMGW1U9Dl+vBakXoVmx3k+BX00/M8K8TVndZtuPWNdS5O0Wf7
ohDdm5PjIczEMgLSd+w5DQHS8p43ZDi+eT4qxAS+oSDoQvDIrwS+8TT+MMhKrxo4k+79QD1JcIgr
mUvg2R6l7XfR6xiEuA6UmWrlFDq8meYVbSFcilBGSoiSu/UR25h2k0iOfIp7ECmFk4Ppwjf7YRNg
P1LkOyF1xgqJNd6GCGdLui3z3lsmLdK/9iU/zqPF7/Sl9jzGSJ8lXQwwNtrlLElzdr9Lrvy7s2Vc
p+0AlPP4ehC5HkjIUV1vnmtuwYkfoevQifrJA9iKYpna6+OgPnfcSY6fRyc8LFHl1N5OSwMnOWTH
IDXK8z8cAPneI1IQz7FIeRDfjG7J7MhbXn4mSNeDQ4jsjXXI6613Bvb6TBkwEZHNwiGPMfhMfM+t
2D1W9hQ9h8V1Ki1/Rj8E8mx+f0C5hb56fcrYH+z6cCPNCIqI0Pk7ClU65HrDINg0nHDyoFdRHjfj
6WaALURhZefFyOmwGCtjPgtv0hHMZYRQ1B1X+6OfavwD0ufPFUzqdHSN2s25bDl87WsfiwjmVU7t
31he9tsHMiblB/KX8M7DW+Rp59WYxFrGlCs8DCRl5TCAVp7BXhrZ3P6opGqwawEfbGmITCSQjyuF
WRXd8BEV1UEx9ERpwK0VhNFf7ZE82HX/oj/lRlN5D/ehw7ter6JMlzMSUYko2N3jC2M2LAxyI2yN
CQnipzT//YTLS20cjZZ1iH+MVirXZThcIxeXAECiNoXThisqu9qaXS6bHDdYvkHcR/VHc+kB5smt
9YDNP1rxkpTS9EW/M4j4PomDbyLkv8QEb/c+y1DY/4UGJ/r0RWo4zo4qn5Ut43Wh40nQw2yB8dqt
PjbDT3m6TOoSU6kJp+fUmqoCg21NA/bAUqOEUEjI+pF1ls7y4EQh2BwH6sCKUXTfSoKJ7nWDnOqZ
vre/QcEwqMkeNkpt//mXaQR5/AdtTlLGn0VkLNaZScpxEkDUYsXHq6aihfLfJ6QxtxnMT4rnimuG
LDdoFG/42IHm4KudxrjP2j/ug/R3vehl8lu7Ku7IyC44KpCUEZnoU2tttXtcUISWBp4ItGigoMYN
8kCmhBQwkhb1f6jP26UnvYkFedgJlEfGwR0UnRai6kvSkaYS11tQS6vEJlzNX+YWXqRJ+hXiX/3S
vRO6CA56jOFoou3EzeDHySjvDrdBLMMUgplitfxz4Eo613TS/otGcxdaaz84c6bmkY2S6cRjZJw/
0BXdTLsL/BXjxcrn2yYq8HBoWALJoyvSvTZ6fVmeEED5WRuNqjNMgPLJkDRW42I3zjPCcElyLyss
5GoRWVAPL8y57enVAWwNNjKW/c3YDLs4iBntK5v7vneh0IqhpXaCHz9dEgNraXFT85D0KM4fNdWH
wkKLwPatzFEoUuqFZLd5b/FJiDdUM+X2TF8TdhrQtPfKXQ/XlYA1r+qkcxbThCmK4deniyAJuAda
hdc2YZeXhnVhWzxUjJJOibxkSBtkJiVzCm8rSnq8mCyLkuW7ft+eixEAGxGiw7hV3UMukpSXFWZW
RsyNBpi2/uIVONMt6EpLCTQbtaYdvQJ7telPCvgf6u7Ay7RdUceeFxjTnCSnwl/5oG0wuoiopfbA
GN2AbPX++c12+cOxr9X6iOgshphUn5f8N63dPG84v/+paRUloI6Ly1jReVVPAUVx+3DSr1v+DwFg
hUvgj1gCeOQITX7v9U6z4Bs7FgH2kOyr4+XIM8ldW1Kf095lltQWZgG4Pb/vggyTuS014s9/Sa7Z
gU5/jLtz0idoDWiClju49gSyf48kuNeiN1/041kml0ZYcs8f9OipGvSH47ADQ3TdqO3ZHoBInjDE
6flJUetVYN0n7sUtMjagFPwD7z5douDyZs2N8UiqtZBAth5gFC38j3PgTeOXoBKdgLKTyLDMgjqR
blgyeYI9VzG9oPyDQxdAi9RhvPeeQf9P+aV6KANJLClFqd56Sq9KR0cN6LwxIb+rjWjbV6PGXlvC
SUWjCWG8dLMVl4wXFZHxNt8uIPSD77qPodrDtW/aIAhZ7Boa76DfpOxpaxwQXlNpBah0kyEnrLbF
1nm0Q1WIDV7r3xEihVAwRQASUU8Dm+8tL8JFd30ij700KHISjZP5NF3zAjLFgP/hEsBZq37DWi0Q
i42jbO6o78awD2cm9xQMEBLfzUB+dE0hwiKyXJPGeGg006d0zViBopbrGIw11S5FBsg8J86GCU5s
8oF1tWv2EdSjBeandSlRQFPMB5OXID3aRf+v0MIEwJiJpRg86QIHx3tNquZ8y5vCrq5JU5tHafW9
QPak+zJcqH0WKz0+nyNnoLDljIJLzXhpFiAjLysrV4hJmSe1eaE5eH3KfQCFdOR90Eg3iGsmUH7j
KwAUutmcmcfBeW2NRr9Zddm+A4Onllw9f2iziIa28exeRCNao+4VOLE9aZpqyi/uhj5plgs/3VrF
a4jkcOEZVKyBUw6YeSJNu2y1DzKfU26nbk8nqQ2u1vLzlbq4knvO0In8hFgiE4fMKzu3hGq3ww9w
c5PYzLKbkUW50OAwXat87+PtTTK30KAIxw6kycPlGq+EbE09J0N4r9TBl8KD5Frifzn3rdHXqJCk
3ACmnkIVdqkyXWFSqsZwqP9ZijBx7/lEkmQ+joFMKYMAFxx35NLnznfh77S3kXSbMD3wZAj3FPzg
rl/0MKXF3wG04e5Em4ZbD7d97Hf5pj3+j+xkR7Vup64pfa+DIEAIN4QJmLymEeLXHAaBpY6hDYNT
v5uVwJI3O2gniOQZzd1kOUcNqL0/mATj/HglelBH1NNx6tpYUOiI1xYR88s36Nckn23FiQKmKnY3
lls6zPE2d0h9mYEbJkDr8fmFTK+SVmaakqxTHASEYlJqKNsIuj1fE3Pab6ldRQ+cB12zeTWFiSu4
DVOZUO0F7T52BB2ifkAuYm7aJKCtWlngEqsSKdySuKaw7c4lSUI8VM3B8aGuxucHbqvvTMS0Td0y
ABpTCUOACyRTVYAYYB/42hNJxIyuR/Ze6UGHW0Lnx0fcLwMInGdv2e6YzKV1pYL11i/CEjpLvor6
x0+ymMCKIiZGWCD0TXsKE9ZGWzsmZbsegjpxg67kGveEF4CSAQNutsJtha9XSuK/rwhe6kEFlkbE
UzCk49g8Q/dOczkcwK2TQZTwisv1wDG3OQVXAH9jDZanf7RbW2/feY8VWtDYg2Ti09oJQYI/32Zr
HB7XaLhvl1B0svEi1F/y/WIU9gyx1LHnQKMMP/1OLHY/9h6UbJI9tMs6T2pAQACtd8uXXnFEgToc
ajS34S522uKY8knn3b7YP5pdj08moKZEFLjqqsk9Z/tjgLEHbkGxO5xEPmo6CiaaWGi3qpjYLhAg
Uqy6iKACHeGsp6DHIlzvLGlYITt8aRZxDxF3jQYytAeubO4nxiCkBWw0LFNoSVFsghrLxTaYR2Lo
kt2aZCWv3KehgKuQByTnQRHBXoOJ6aHDSK9fN/+/wiuVRUCZvveETQ51ptYdfcDdvd08a5iLnI6q
9WafYg9gT11AEIKs3//26kJC+/UEXCL8PBZoRKR8wab6KaqI6ndsKF/n8sa11xpMQchpRSMH5TXH
BJ+n5NMsmzA7kcHEaY1TgishRleRjsVdw+KloQCNroZ89qlc5DCuFugoIsnzxKAC9rHIktNQN2Rc
P8W1aFqaxVbhW3XgDEhbLWDpAzRp5gmH/1S7T1gytO0MvLMoVyNVRkomZxE2RLQRbqNWyRBW0dao
kiiEyYhkXbcOtlwj/w2EeFGnDSPT02bkg0DtPflm+2WBvI8IfoyWv+KqxalIKi0f9WdQfORWfrjf
E52+1q0DBcdZmADQ6s974euNkSwnycQzTraq5a8QqaTh4DNoGos/It2BIBXi6rUibCW7HBIJse9y
gPgHYlEBmAqI0ueA4iMPp6ZZE4JWzR/q4zBVk0uMPiLbt24SMLWB6GJIXsaABLnD5otAQFuPhIDF
i5/+2LONJO+kxjDKCAITNjsb82len4eCK8fnFkmzFgbgO8QvAe7YX2w2nG5QL4shF2GyJAH62gPN
xgtoc+s70t+9KR2wShIzpvww9PFKLflW8Io7JenIDNf2GLr2XnI3U3yNRQojKe4BvWarg1wRovLx
UqSkahA+nsrkDqUW7Ig8KcU6ETFt4KUemN/SyrkleA3bzVgwzoi3EPZHzWkaZ9VYn8NVurEnj3ll
2lOfd5RPXhEiQB6g3G6IAfUSOsoG8rSdpHSf5QYjDMsNlifffCJ/t0zLQQxVcfUUhJv4UGEJ3f79
I01UGmjMIQSYUe7gDZJJpj+1YjXNYhCeE/LjTRKGdaloWZMKp8Yj+mxidFMHTLw/HZfFj6biF2NT
0999Ej5LWjiOaSulWbKzJVArcc7SDCQasXaDZ+/A2hIx4lJUOsiNmaAhirTj8CxBXF87isdp+oQm
HKLL1/h5pq8P+pHcPY0jAKdeFT+9oleRScKZN1qHkXTqVYbiAoyvmR+W0MCVkvLxHkRRJw+OdgEj
89MqcXxGMZOIrbtiHlxetkUWa5Yg/2dg1JEIRU8ipKMa2yRoYyXchutWOGLDlUPCF1VLGGLijaQs
SzhS+IjFPY6FRh7F+zoJmMi4+VWifmFtqDQxBDSjnBm0FgB2qYbeJsGL6y3mVjkoGKLr4PU33dPU
Lu7teGwCoqwM9g8J+uHjcJfpalWxjpbd0Eme6cLA3sMTmf1m+YuHSEoYAwxKsiVhMt5N3qHBl8ku
7+e4LA0GIobTzuw1UmT+akYArTtUt1g2+BTJL66HOOZ+WTAtnV1JtkgpAQhUc72bx0tl20eaydVM
NlZHUKfqm/4spR2gNDKjLZrVAyDgNbcdqsSew6wZjHcRj2GSWdVCv138f156NeXyOmdPDKvGrlqs
1/qQq6SvZrVi5hjm1TgmTZgPX+SkhUt1cnOPuTDG9KH4Yp5mu4gKp6peU/E0DS/Hm90o/E/QTblm
kTl9Voe8wQiSBCBnMDM19vwAg2EiQTjkJVa4lVcDqg7AHqScdyuMCx71fnPpu3Fdmn/KoaSaSTYV
i8ANglE9QfwxusXFvRi86XUgq3+6x5FeziAfvQZByg3CJxtaWZSXWVK7W9jODZul/Y5bXSCVCexI
c73Vt9q1D3Pi19YBYgRpA4YH1UJYA1o7T4y9wXgF5nCe2EwDNVHGEFq/j4pFdI4INOO4dm4irdAw
ovVTF8zOa2BdiPNs64P3GY9Ae0hWW+a+uychfv3mnzKmF8d5L1cksfyudKovcMqmUa1cNBjxDGZr
1k/hRqjndzW/VYaJeZ6FhadpjZfI6GW33N3xtclYzVkbcNdC+rqElZo01mBnb3EJOkaU+peTCJhq
wDB4KMrRgZot3H0XKF2TORBEyMM+QSzapYW6UclSr9bwUk3mtcv1+FyWJhZPO6+A4gTE+Y/xYLrE
ciXx7HddR5l1n2O//atu3UrHEixl2vYvwFqGs3lqZo5aBRfiVPQ0cBssAl1MQsM88KpzitMj0Rhy
Z4SBX9e76sjl5nV41HM6jsaLwgzcLwDWwghIF8onQ72EEFFaQ/II5JbzVQO62AezNUA7lOF4ig6k
SwDTMxGqrDDaN32uV2YEqBC08DoprcUBmDz7uedPWiy7EQv8QdwF9ncd6cWaOiPPV6xQeXJ2B6Za
aK1GkWKg8etFdsJW+B3j+lm3vyYR61hxJatx7VhrJKtlDwNsGZd3wJ7op/XYJWwp42nH721ySJDg
o4P2zaPTQCPsf4PmHVHP9hjhdiEJzKUi3MfAlDtMFYQTQhLje+s+1IitGq5WoZ5VC847kRWkXdsO
UOK+RxeHyBDIBsTsPw+rn4XS4O/4JBN6IeeUSsDbsqiWpdSahkfH/FnWmx5trJVIrG4KqDyLjndW
Vu5pb9Q09UQUUIg40hffZSefdaJ0zzeIjt3Xyatk2hXBkT925G0Pklbu6ukWoMPBd7No9j7baDaE
1vJJ0bvxRPkFkKeNXwcfN5/BSxS6Gx3/VG4gGOoC+N7DvjLU/QvGPjMyTKFnidA/DKQQVy+4M7Xx
moisAw0FPlDKH5NIgybPP5fF1RDBwRUOlmx0AgqKz6Av5zAeiuYMzrWbaLtqncE0nGAI+hinsfnR
BC0iKPHFhde9aNBZoqeHJN6o463mCNTdSzhh4vDOu97nxqVt4bjjeIKC1dKO6We6ymgq+6c7KekK
x444fSrIhrUVty1d4ToUC2mXD9+KDEYHnhPoI7S3+/gp7ColjtzOT5XT34XKEefZiOuC0RraZ9qr
aFHXEw0mGLcxzBuBGiiYRI+V2mDaaeAcbYznXAJAg/vI728xDpbfSZI7JRx9jeDXncbmqM9WN/3A
ITZWVR2tiAm6qv4+yFW/BUaQGKFrdfypZq1nTkFvriFucd+svD91nOiL/vlf/R/6DdUyVq3FP33D
hnrn2PucfyHSPI/6RizgAQubSigj/19vUmRFfsXHtmWJHHnsNIB1XiolL0LCYrSRSjBvrUvLqoY7
Z4fx/cE2jCgS8pWD2OekrFbf2WkzYQ+WeXOuGQBe5c9zK82yb/xPmQvBCKs1BVdjAOEMboolYnaS
G6YaGo5JvYu4iGmLVFP+BoU5fYiUaq3/Va3H6FLRa9QzuOzar4RkuGl6V4ZZb7VHtZf0So/WL7Dh
P5nyFn1RBVZQNM/Z2BVfTjioQ6BjfNB5FRjIAqU2Q99/9TmTVi+fffB3d38Cvem1MSq+FWLxPgag
sJq051gxPCq+mXJF7lCs8voYZZOzDBY9h4KZSn9nM9QGgeS3k+NuTvZihztKhSbqUJwCU3j8e63Y
kShAk8CV7SFGM7fUCq9Sdmu14mhIlYNw+i/v/2gdhNTyNN8aai+H3nqTUlI/BM16fcBGxdaTXk/W
Mu6vYsK82IfOT4KuPileEVw1vXrql1K52WvHTHPQbQh3tmwMQVUKzYfdpJUVI/lgnDjAJsKfK87p
fLBOl6mskWnbG3RqMsVYkzZkfLmS6j9wzqZNLMatLfVpl/tgQOQdskI1HhMlTcCkZ5HiRhQpxUHy
RVDyD7RN9s1H0hIkSPyQIEvogUABb2LO/PsRZNH+eBJN9JZMogwtiOz9iS8AhYHyxjW0v5hf1LuH
toehqWJ/R6ZgDzSrOPc8dMBfBRC7+lfGy9QSuEgE4vsBfXolYaV+vlJx00UIXDiuQgqtaqOiYLle
X93rQ0nke7pGMfuYKVihibaY786u8pkctpFxRcui1VjXD7uukAP4kviX0E1O5oy5Pcq9ZKEc6Y9b
WuO351ohj3qWuG6xdP+mFAYy1tshV6+y6F620A/MM185TyObdT2MHe6GouAJNG8VG3ki3DwguLtj
mu1Qnm3PIxYMpb7thnkeHHXwIQoTaqjI+kZunS7qh9YvwZggMK74UMIccOBTUTlMfI+Pmgzi4WjM
6Ix+yWhqRdCQWLWJeo7d+lvqnoVb7aLTkmyc0eT71y1Lxl2cvxu+TfWYs0OK7BnVpR+gtQmkz9mx
GY7RNDifOQht5yo7JM7AKgDl9cyKh7uMwpMgEQno45k6HWuQ9zRlLFPj4K0wDk/QeLEIFHZfrqJy
+TtMLvncqEYDLcjGdNI+rE+FwWnJJjGUNcdbQZkiwoE94a6dvIhY8dLCvE5Nqtm7Jyf3wHJdyYjN
I/pWl64nJ2W+l7O7kOqr2iiomeECjpXpdTWaUCOccnpsMd8XFdWAb2DnxkFOOdA5qReIT9/fgzg9
IHyscfAybHNTbEZuOIVlULWKn+mEqO1v77kgm2ebsNwsMDpZJehkodlEr8iyLB1xoEANRw9SqOWC
ZXz4PF4ZBdnjI/epvjIpZWc8ehIuHobJTaQaof6cHb7s1bz/oBsGI9FqNtlhXv5VPMPX7bfjARtM
T5AA2ZXbamCTx+ubyWSvDrO1b6Yq3ptP8/4cPpZXVOqW4Us7YDkE5MSsBmhtBw2sawkuk5TuGc0Z
mngJWBvm2ZGe7OIsl9h7yDzmMBzlewFn/CeFZryrs7Jv1AbDfJB1O29H/nDTLkPKk2QZlthQOtmE
MtLsoep8Zpc6FTaiFLsSXbXgaOFcZByICUH7zSeuxWtSJm9+6fBB94M1Ln6KyPiCpw/oipqAB4mY
UPSwkdC08kqQ6B24PW+eAVGcdiTjg339+OllzfQBWuqm9HweVOUj7+8gr29e9zy6sp0U+7FYIKP9
YTbDHBZG1QaRIZOKDxjTCcXiy2yhxuJhMWeU7e/Kd32i9W3hwaxkg8upY3bOGG0nsMz7gL6fjBZq
fqj3XOepaQj7twrpL36iwI/1DUZK//ErZlcOojE/89IeAdm8AhFG4gxCM0zqe6I1w0BLVVNMKio/
/M+HhfQoVphtIZrah1KUf/HbJimJXAd1dGVbLjmA1ocwXY3WNz/noLDKsNxpwX2vQGWVjDipAxhJ
oxRQlNE1JtXZE1kqToUDZZOXx3MGwqjwHqCzFV3z8wgWywUOzuYvXMm/OIBWaYpOMTkLXJWe9teH
IILYVHd7OfLbQDg9bLtSiOP+NVsXqXZN/nBver0YDpF6QMvzTiAGGHtoIXyALQr9CfjHMhndU1T6
fil7qy77XOU5Q6uKHBtsy+eOGA6EdxomADoYz0xWKj5MgINQAfHEWdzuv04SCkUumlJaXYV9C1p0
czC+yAVv5PGO3NSfufJiEkEG3tp6L/Og7JhcVtyZjfqiOO86Pe02oVa5/LH1w2RJ4FKZb/t45utx
g1wtPVhRqs0PDshfvRv16iddfh2fjpKDhDYG9Z/L6cJ7mRqqkGephEIRNRQKqeqlFZ+a5uDPDmwE
OFhtbUmkqqtPkHhQIlTK/0NvUsRjCQVmud9mUmscPAdy27ySkW7RV0SJ9byhvQkkPpriijuogE2c
D5xqkyE+AWgicdhYF1desgyzpUIfmFSY1q5ngiFhGdfWSiHtwjNM3QMRl21NysmsK/CfUfe+4tTb
fhdeiRSAX2Nemw2lqK6fK+nX7aq1EL5Iqy3Q4o23Fq4F5bR6leQ0ThUbw969X30sNe7Ng7uCVhZx
vB/cUHpQzod983YTxpPsSrRFb8LqN67naJzJ6G81Pi6Xr5pD2PHX4z0627vkjBaIfqcytpAFgdWl
kui3pKnyEh6RleqTM+riZqTQwQ5wmnF2JzbptxaDaZk/8G4C93QDnpDbupYRX5L4GbIRNfjuG6NW
/xINBwzT5zrbHvov/2+pWLa5yvzzl5wArWkTERvyGPoJPaIbecwIvKZCvFtVMRcvqHGZ6CS6RMVK
PaF8misN9eaP/G4wRU3xMhBETBOmaFhiXa6IRYnDd+nfpXBs9JoHqNBUKzkAyZCZCEnQT3i/tEr4
AgoYkFy5LhpYu1CBFBiOdWGs5oh/I3SNuF406vICPg+A14nfYxLmdB7rnCTd5Mk7bAqNxVKaO5Yq
UlLMLArN251x3ePxXkAuR07wNBueMuU3bIRS6pXUbNzp4jHiWHVVFIMFx6j4uHfSJRfu/7wCbaUU
gURYAM2U5D64Rs0zQv9uxjU0iJod75jwy1BeCs3EVEIIYHPz4UjjcFjGJPCpv5RE7eMUVtUwIYHN
TXiOr5CezmJ29yLwWNKvfeN3ARQN5DUesS6H0lqdkGkv/OYTlgQ+aYJR0zT00atZ9ZXRgl0i8/Rj
FahvzZaUM/TLaqqkmELpJzOU8BG4Yn03/dS5YEUuaajKvJBtPIirRnJqD7//qcUYbjssDFirWKHp
nsdkwQ225Ba/HhRvi+BjMGtplyhAZyFk9tVvh8fVDL0nbT73l4wwg9y6tNEYQeiI55KTwFFwldYn
KdiTKnZ4MDjdOy+G9Wv9w26zUJARSKNWgeSy8nA9Gs2zBxslH13q2Y0KhjpGYl0n25gwhAt46lNa
hGLLD0sOmbInn3JAbGB1uZ0kdj7vMSPcYkBRsyMt75JBt+3ZnEPYONaW0PNjER9hWWdjxw6gKYAT
c+/RaDDNViwfxrEH2YtL5f4BrqaviMDuM/+tpmDeDPqkLERS7IUCwDncIRI6OgIQ/yutJrqeAm8k
LJKxU02JrrwR4JQ4DHDYncQqHffXAIdO2D/DAQWcQv1Zkx04/JhSK/4ajBQOooPYj731h3dfNKjz
/9sZOevwHXFm5sXTL+p0HDmIT9YvqIDpIpmZZY3vLjVeVGdxyeYsGdrlP075lM3BZ6pJwtSSGR4h
ladckl6uzX1fT7E97pZE3IXattjtYNNPB0e9Lg/fa3hMZzB7R2X2jbHfUysXjpNJdVapuir4PMmP
zsrgPWoUP/Hjbbadhd9PvbmdiOh6npFZH34+jJbg2Rfowetjg2zcoVPSZkJOlVis67vydd9N3UCB
KiiebvgcEprb3eRrkVWivq3hMk06+Q3q5nOw7aA0C3UuQrlPFngViyxxl2kKvt9G/u4JnOfjsK/5
lhFHA+Mdo+w38le7E3NEcMUGNmRz8PTgfogD2jsjFF2POBRszxexpBj56IE8rJU4SAOT8Kgqo3NM
gM9ZIkGtO2/gG3Ayo8nuyTSL/2J3Ltl/2e5EZg4Hb1pVnDgBdZ+AmcAZj+V9bxf6c4FVuXqK+o/e
CtAwiRJOIid4U9PL7dRqO5RjpxzzZ7lWJas79hnuuY7x2E254uVOFxVMrf/9JdXNy73zPSm7zjwH
uwx+2QY20oFHvjUXr6OBTBvxo0goo6dkuq9nFVZ39FrqogAirc++u9m1E9jdtECwXlmKB02XeLpu
qabz06Wxy1PIF5RSPjypiyeUVe3aVflNTSB9iCS3GZkv/LoKXVoxbsTOn2Ry6TgWCmzlSXd4HeM3
qy5ouIrpODCBvjq3ByemRy0Qylujfch8orefYLSNClDW8vVrd2q2wSZ/mPxDgOO0z6CdzHJv2U4i
AiZaMPi0T3GECDsGOYbvD/vgQLHLX5FiEyry/zvrK34/kSadN0fI733gY0dfUGA69ppdTHbyjhCX
j4SwYRaslWOJvb3AdFshJ5gRO+Lhq72Ofg8kIY4q6tBH7jndFS/ab2TfQDNQs3nDInlgg6rVHViA
2DcHkERaDuVfuU7HXYqK/+QqO3VQ5MpA8aFmGpQl5oBrAH0X0eXqTuwxBHSSwU10o14RLwZTcE4U
bBkOD9ndqJGzgOxF4OLQyG7pvXatmocu/nSVH6rHYpxvTaH9+3DLISbgQLDF+8x5r8+oq9F0PBGw
koYYziikN1fL25S4rRqayglSXf7cv7Y6bwlobQMHiKcQg2rIAxDotr6cf2TZdji2fsN9DfdWzB7H
fSu61gDQkJnlhQhIXq2eLuf6eEd0WUndC0Y2GUvlAbqDZW/IgD2WVPU5Hoqb5kxKPZubx35m2PRY
N7+nZq6y1llxX/wL6GSeebyu41Hi4g3oGc9nku9i89H8gMKUYKpDJWv3JpNg05evRQylatx9u3/p
uJMa7KftqKgBGeqTAlHHUQZiMZxqNi7OgThcjcFZ0/2p+rS6RVDfo5bcIXpajHyDOutVMdFRamL1
a7MPAy49LUWO7GH5wKnWvQLWtAxSpqsyMOXaX6RVG0DPoxRTYjqCRZYWoFoN20PjnWO1sB/EsFOK
6fhB/62qyf18beu+mbYLRqLveyvYTfl3TKGqwYVkH+9MDgkOOmnp99UIPUIZMsOqPcpNLpwc1o1L
S87SlneEGXNA3mQpYeyFojULCmLvaPB6NF3rsCxN1cqzDzD/11dhiR/mBpVTtX4Y/hu5ZGLDvYO3
dK1SDIftATwr7KmOAP0SjGgqR113k3CB1hK6OUYoKv4MVY6I37rVVer6keKBZ0M0l12k+KyBH4pF
PTpJlJWyWzVD+Hh1ZdU6+pmu9kST2iri/yspLxdeApsL18+/1cZ3BgkLXy+nghV8TATU8/7DLIcX
ujnRopnrcPLfMNUU+2naTO0qh/IC8cU5vWP7SLdHfA8sBCAjYu/Xuv8LBk3NXv+pVJS88D+pDcPu
vYpSw1jnhr8mROn3HxQvSKBdDh2rP66Cw+I3IUrkbjoIlLSKxRrwPQ9r0CPFWf6yarzdwB0rN20h
HCXf0Gmi8fLsuLDMLcnr//CbAKGJQ7CojuEYHQMdvaBzwESy2FyXRCtJi7HztOrbhdLr6yApocO2
xiiTG5tJNTsRF6/8dCcAy2tWcbufsD4KDFcQRaCETnAEfFqdWqoTLCXFe+9HHzAf++idEB5JH2kq
pc2ZD37MeD720565jtp7xT+fQkVNkSdwcNhKP07IdpFqu5vRAg1HTBVvxl1HcQbVTlr+j4bnuTDf
FBGrReO/lhbKQiJWuPwaCLAZh2B+smcmv/op5pVzSEOwKp6W4i5vybobSdJiPPHvJSV35SD4eWKq
wtyC0Z9Mgyb1gQEDnplONgfoEwK7G/n13AEsqpVTlxVGSDjc6+4N3T9FBLrF9qiC/eWY0y/UGsNy
4ghLsROKAqRk7lJkiSkrCLC3qeU8FWrVf+pYUMULTI28DXkhN1cDfQgHYIgiQTmXZtzndNy3DApl
1bf6WDL5xU6SGYGPl1nDDKcOc5rGSlgWdbPs0z8AtOqsHKSyGWH+wqVxEBsOvUYRBxt/gLZqiczB
wLw0LbK6QWljmVCJlyHHDrCl50jrZLFQCJ9skalFNH/2p6kJybc5v0oT8bKHFVm1fLxHKk/HSWJk
V2r8CtUhLwVfEz/B8xqdzVMjS0iN0leh2kSzScSk6DtX66bbkhJ5gjHobGAQEIIKGzA6XJyhIJjE
bLGozU8klKC/Z3+HC3P2zqPSlPr9qAUpF1A+vgWbgOqpXLmk7dbGxy5sk4EBR4XpC7WCRa+oY5SX
O4bfzZtKmDPueMa6ZDbp7DZUlEUhW2urVqpZ88oxUS8S5rVbNFwQS/hVlV2VQrVSHrOV2GU2CCT9
G9+7cu0cX5Ibz5tb8mDCVpEUe9bE0BHIZYhfS9UCzA/INg9+jjlXBaSpafJQLrOOW5HSa64UxN8K
AJnB+0T5AI/kVgwbyU40lUXkuS9xf3cAeUIwP/ntBt3xckvl+QgpBU5hwO8nrZdFw9hp7VLTqk5T
Xv9dOWjwo/p2eK69SRSLonqIGoxX9o9Iwy2ksf42vZtrKfOSk5CNqjMvrdS/m9v81TohL+bn9QoB
4J1uuhBhGISaJTTSB42ftXP2aghNs0Gci2Rc7ez+Xh+WSe6LlSyakF2adl9J0rU70xiumL+fJFYr
HlxgRrtWLrU0BLv9glVa+KJqhfoR7zNjC/LVCP5hKeGV/c4nPaa8pYXdQiWfmVv1Pss/Qwf9IM82
dMB0eSXmtn5plLNVVJaUGscmhJIRZa47lR4XR3Tez4yWZIZvds+jGNVRfxYFFbMTiwwG+2k8CAQo
SOkjxA70qZR6M7IPApuawugzyBm3M0x3XB1wlwOkuxXhTAhDkOZjq+Es5nlClN3hepq0XRRk8nKO
gJU6hiEdWI80DgLOg46/jwXs5BplJ7RabuuYjAF9jpaYJEw7MvzCV3fZStUacf3G6exRp6Q6JuV4
Aurz1rZoN7kMqaWVz4YJ79IlZUs22UOwn6e2b+dWyv9cUBWUt7+fSy/JzATEGli+jxE9bQUlLk+F
OM619Z9G1lqh4SpsDNaLSWmRIuYWLdt/aqQwkW8BdCgFcVZLUOx+xH3ywbHVjdvXtuYlQPal3V4D
w0WpazNwfHTGGAU22Ho8ho+8oMgZlGxzO5ORrBcKbjIp77kxkcYnHivNhjKWvlbrpu86RW+11awt
uwKNaVbZ38qhhIljjae8iFiR5nHZSMGAeYrQgS39cuXcnht3YLFg/KNiDj8E0M8o036b0o6mLAWR
LELHsjSugarNHpNBxIdZ/Q0agKMcJIWor+SVgSE2uBGwv0ZebNRva/S7HnzKT3bkasiG7BdnQMHd
ACSHqnZZ4294aC8+DfNjRL7JDB09e4BtePpzYaD0Zr1P7YTqvfD+xxwvYdj1xdba430+/nZliBxq
G7XytEt6mypnlcI4HTJ0maw/ZgaOEIZYL+64YfF72rtYSqthG6HuhyK5y9UXvsWApwV8k2Gc8wvs
XA+z4xNIIjXcOkoiQXZyHnZU9PTkY0xlrolXtW57OFAqr6Ua4WZHR8bioUaFHoTWSiurIgzh925X
gNBMssft+kiMM3s9BShuzpk1UmrpgBA10SnSzOVaCMTeTEAql6DEs1LVIg/DQjM4wgJpnfES2KX4
+NLoYcT2BvkTY3E4eyVvJscgqMDDbAlYKctIMHTv5RrfU0A91lG08ycOS0yPqIRwPq6GfBK+ObOl
+Agv/T4vFPvysWiV2vBKuHkSSnAb/7N4I/VtlojzHWxeZ1tGencH3DzVOIrF+JA5lnNygZhibpnp
VSshOFwmpCZk5CB9YbJS6fruCVKn0ex7Yx0hFdqimPaya6CbFGjw7TTYNZOkNXEma45/AMNXkEjS
dLEhvgheJDnyZzWa6gynXMcMkNukkZ1xEBqQ0CRuOzwxD3qJXY2Rk7em+NTXpjZBOPtmqmbkUT10
MEpzn7x+meQWc07rXaAQI/UxnlhatGLen+8oFo4KTPA+mPEssiywTdOzUTymeTZH9FaylBnaBwzJ
IJJKa0Ii/KK5xNC6NmMHcIh/XRPu1SlaJs8prx1zCmkwQbZPbiFU+tjkjbQCf9NY3UUCUrbBm1PG
/tUNZbmzlhNkTRoESW9XAeE6X/6zoI+s07P445HsQ4cXfi/o6kkI5mue+CAWJP2kr3TKmLb3YPnK
Iu2L5XExaLxVwgdfSG2Xkbrs0rznjoBmeMk5gbcdypCWIauNvAx7+qI4+rpCyo3A15q08QYHjrl/
UfpcUxaCjsqKypmZrvApqyGgV8dmm4EKNCI4jR90Gw6I5tAGGmnzDMD/HPQ6ImPte7Lgj515Qn7M
08EjxcPZhppjfMIz7iyjMHaVjGY4f0aQcjW/61C77g2VOnd5AM3FtgLfgqJjMU9MIJt1PpE+Vsb6
PZvnaAG4xdfZxR2EzY77vUvbiV++ao7xSdc5kbKA+re+nnXDpG0YfGRIr0zZdCBdnSWPKw6Skfbp
FbAIHkWUUZZFbVtI6Gsygez2Js48YkRpBr2bO04ccF3EphrP8ihyniuQHDIfe9yK67lQiCrMdjbQ
wqf/IslqCv1o4xmvOcQPpZ44Z55hXZ0+ZQnkqvFQB3w1TQdJ2Gqcf9KL+ptB09qA3LnIcN0s/iBE
3m+hTq2D41/s7w8GYlv9p3Ws7/YFz9A3Mgvf23cbo3127SipQbRmmzmjQ7p+Zl2BEu1AhCKpjJwm
nx+qZb3V0QKaYRxSCmpZJcBCQPr5dN9/Ed75RvwFNJ7FgLODYXzcmHu97vij11PoCELAnhpDsuGY
vQQcl5/rj5gsffjfn8QjGKurYGArzOLtl41VsWD4yTkygmT4SdH48waA7KyPhrnRZn69YSVZiAoL
scv0K0pU0UUjrGX7zLOFbgvd8YdUSxCiQ5xXDDcH7XbAUHzZwJ9FZJoEHfJRhcO7Hqm30iM3Akd1
hPWJiDnw4X9e6bSRAVdetLJXkJRYAp8QvWSjFkDbgWGR+HsoHovzChF7VW2L38tiKcjtZocXTwTR
wJxKxnDncleh+9iqwjb3FDB6EmnUtpfrPoyOrn4QFDA5+qWD7IatZ9+CjLxLgPXq+JdzeXbNEcYE
iZ9vKyS4px28g/gmqMpiG2Sww8aCXLcRkaGJLP3YpDWxTyz9SSvLclzpRh1KCNWFOyJojZ4yk4k1
Y8hkqqrgIjlkHyC1h+U7W2UMsgImie6qOyAWuLLA5iuyvUUzQIxazMiQAVAwQIONgok18ZEiMVw3
iU+6y0VoD7xGfF+pYSKURHNx4TR5wQb425wPitcvhZ5MSBFkJihd1GGhuzHW09p/SBWBcguNm2q+
uJgP+g/rhOQdv5jmOaVUBUacvmXFRmW0GNgxUlfd6joNosR1pAcNrv7RpNjq6plNgxDrgTE4Qsj3
qBPPSghCd3H5kLQE5bLXizUCXQUob/NjN0EzN2C4QGCvR3J66D1DVPI3yoBjKs5fAAdxdMk3TGxh
Z2cC2QnwOS7mfqLuhva2NLfMokM0L1zp5nzCUpDhN4oSnUb4aYcvdLdIHqNlJW54O6ycZtVq92BU
Hxxqli6yE0ZqdgOcYSwtwAugKsFjws4O0x/wQiWDN17/FOl7fEIJYkrWOJ1cGYlBybf7e7syYvq+
GdVVCTwd0MfsWv/F5FpOZs8aUhDZAfN1/sT4cURcq1XtjL1cIoWPziEp/05xo01o2lVCrLrVljEz
XszwuiH1QdzgBUzSVwD2qmcOx6uLLOfCnhaMVoFjTnOxOSLkewdF/xqc66vBb/n++5yAEslIJ0x4
OfDgkObPfRTPx8udvRs/kCC1PwZokSUu2Q2aC4IA43d6j0xLv+Hnps/XOFjCfPzV7YbvRR+HGCR0
WNZQ59ihPbMeljyrQE7o3UUkHijHkVBjx1uxrPF9SUKcDZuFxx6i0WKfSa0TmNOWWkvtkHbN6YIW
joErk4PQkmkoKYndxAhQsulLyfGIyzIMOLB5RSo1rACGT2eX49PVBhRLXRhbmIMxQYVmDelBhYTr
rLSjbomajzmnl+pG2QPhMVRjwJQMp61q3AVWRIsbO3BLlRkB1gS1aRS4ZIfb7sLGRZvepPciJQVl
o3xEHcE/WHGEelKG+4S0NHEPlcALw/95oOncAasZytnQD2ZdnvaYknGC09jChIRiCjCE6zGrFQtI
kPqIntaEoiGh2jYsNspDbQU23UrT80lq2Xvc4r9lNzT5oBCM3EcePVdxxl7r+5wjHALH1ZKOTOp9
A0z8iRQVon6l+LMF0uC0xRyU+JPOWS2iFpJqKJx9d2EzoFyWvHcx04cnMxWlJo19+W8dQhvs7Bqu
nRT77kCgI5H+75iioL7GsQX6bHPyqm6XLjCIoFJ802yVtwY0WC1/cUbxNUzTgV5X9Mjokk/+tWLU
VJVYt116D0fOtsPWXmgi5KbOwOKw95lEU7BRgRz9PrDs6ioNJGajr35G0AU7n8aQQVy5nUkzrEsX
pavJ8lR7kWtY1zTYMs1ScpZnwN+w5syKY75Ninw/Wq+NKywVB8GgOga2KP7ZI7jFWJpvM784gvmO
o9Y0rHdy60trzVdOohAQTTF1DfluCOcb5opA+CYY4FO4bCT++6fpF8bnKlhyQ8c+oSpi1Ic9my1N
tzTI254S1LRP4zoT/PoPlOTANjju90jfjqFWFAKtXDXmif9PHx3GdaFyQYXMGtUHjh5sEVlOyyEC
jJxDXe/VntBcnYrJI6eYfEy8SnKwpwYXeeULIVuGBUxzyAe56BTCC53s6k7WqcVYgWMeIe5G6L6t
9Wxcjfsd3THroGxRrYt0GM9O4/zRc02zLYLjgFSw5fkTkvxph1R2FBDt3ELtBYR5yj4B3qTEGiIU
3GAKeuSAyboZyRU3mdRIxBC4dCPzCJ5nV8R+0rz+tlJI//WdjEZLlOPp0qGvKI/R2CpOrYKwDCp1
85bluXGuktWG7Jgb9emXP5nsbW6+k5QClQXfhxMquzECYIesS1PH0XJ1fab2Rm0NOHi8In/mW+0Z
I1WmIDw+J0+eKlYZRxazohUEwBBFmqxPwhQiejn84aiF+5KSKpBR1yHtIo4RI5PWETKvAe0ark5g
tGeDfHJiTyEERZl7DJsohA4wZDYQGPfnesfPliIPO0p+JB2PBgj5JRc1Qms4gH2+B24eQjFetgHy
1dNGmmKBbHSH17GC1ZJfU4iIF1jNo1M70NQ5N3gQoibi4Z8AwMEGMawIbOg1recdcHu69uglGiNz
swfpsTbQjbF0wcKpGbjSuKSLfxwURKnHpykK3olcJUQSaTzcpy/peRI+HHpyVU0nP6pnFUoc5kAB
kJndYfWqqO/ZHDm+5Hz/nGIy9r+fbongI3ohZD+U1xnByJAF590iyh3ZjQVyKyPM8m1y7VCDalpi
zfcq3gFHwfNpQifhVoLSVHEigY8OoruB8hl1IkLaI5fj4eTgTNe0uMRj+0wwx7kF30LS4o4tJK5P
j96177WQi3l2JqjW23vkMYAIfrRfan9bicol2EPOlurf9qTT0BDw+em/nOonTf0YSzzUawP1JXns
dCIyA/Pxa2v61+xG641rhvCw+pVnQHG6mg4TQqu7aLEzxIH5QUIK1gubcurqdHiTpPz9X79l8LYr
eYq9wvipuX3sUp5SySBjNsN7iIZ9ArBSNSmD7jMy2KCeWBr+LWTBRrd8QxiHutrgZGUn/YR4s/0f
5N4iabL7Sg75sJO8TbHssAhLW2mVTlc3rbkNb8gKnub4VeYO58Qe4CDOZKEmm8Q64mfZuUvMJnrz
rNI1g/2yu73ZTNRJngMYrDtL3WEWwGbw+4LQ5uZfV0g18gkGZNNfvHg7o81tnEWf0e9S2tK/LFaP
8UaAFuJdxh+4kKcb3Mqv8nrSQEZvzEpUgtNd+kkaODeatH0p7aBNdDUh00TDiHUQcoxznRzjxn9Q
WZg8bml9ZKjNFlAm4exwixuElW2vnfeL4o3r6kYc75WcZxfr49WfBjVZh6c9MBF+xGGKx21MLIEJ
UuUfyQwp8a1xLEIuXxel3wOvVZbdnejKAopsh4HUzeoIivyghINdnqN2beEoORbEKBBRoAWoKXJZ
vKrl/31S3G8znYmufjYiIw/YHRzvFY7R3BeUXiePIxPplqoReXQxnBMQJcRMnnYDCKLt+XbaoQ4b
BeIXeeEcqN4jpl5gFnbZG3dCsgCtuM4KDjCq2GxFPWyj8/IG9xuGB6hAdLXlJfptNAnAbiM3ghC5
p+5jjR4MgOraSdPF5G0j+6UAKdyIfduxeL6lt33B1z3WQHBFSidLp0dsjuimk+RtLoD6VhZJtFNf
AY8m3q17792w0hupfRFRgNbKHdIE3Ty4TEpmygvpcv3r05gRwcUuGxwLGXOGgEmvnllV7T7bLdXf
hRVVB2BlifivUA5Ogk7a8FOH8x91mXTNF3bjmSQsEN5gJguIcg48IS2wDnvJco9hpRpBYTOqdtBG
IbgKHjs09aZdfCGgbLzXRmVFepf+zAWUJaQaWcwCUT3x+Ux/YSmKTaHc9mPOHU1FsvIFi+RpW6xj
ptOx95/vw4ZAU8UUHsjZkQJmvohq0XgLeDNe8+2OgRxM34/ek6eBV/42s95dApNY9THhi2Ng//Ef
EZ6tE28RrlGntAslHCZTEZmzsC9Wmyy0jEdIj0umsA2OIMImlHoVg3pzSp8Z6dHHy6NSv8oKUPgp
++sQef4d97WybGzyeDg8PhpreL/CiFLsG5H69ytstUH1y302F2ft0HFsGtgesax5mhXwpfX3sw71
brGCAHheBgXK7+IT4bS5l+tQxVHyDBW41nv7uqo9K5i/Ky/WsMR9oIsycknkoS4uw0CQDDV1XfSx
3KgJ0YPh9ogHC5jyj0ECjwklKGG+3Vo2Jf/yI8YOtKkEyDtYYQt/urb7idw63oXpXrrs7nIOvivM
9a8o9qB0jvEk/yIyq3MFs6HhFO4vghRbSLSZK5kV/2WqADdESF6jfWSENB8MtX49jL7TT/o35HpT
dJrY73ktIFypQy6fkdL1cQzVRY+Zs6zrI0NbgSZ5fIBm/aMMvmjQ+vBQ6lKzcu9jhyMV2C+oTvZs
Hox6zlg5tLwITYpeRUltPhfYTozYdhmRVLZLzSaY9PXQXtWG2nlSQqJXQni5YFWmkWgmLZy1Yi9K
g+R/YZaXcvjbWY9gGWETlJtOy9hqmmFyFlq9xdp5qXF/cA+j3U72BrShnwR3eLkIs31Rkqawqw6U
XHGrSZ303SssK7+NDgpUYj/HKI+L+C8aW4YemAK4KNQ+/BhLMcMuwPmdR9MyEuZOEJ9Mi+kuhMZ8
WtxfCb5dvr6XCN3/Nqd+fLTEpkLqaZIhf7/iEkmoyXhAF7WTZ4VNE/GR86c9cY02O0WgEYv1kuNh
sx6EXR7ggTphvYznZdv3Vn6nc5LE2aYvMXB8oaXIlpP0pzVLWfWEw3jrcbMva7ovDB84vqFSUGjO
KeWtjlPQ2JG4SLm0IcFaYXqkDle3azZBueqSmCaNh+mekOoVCXk1/SnwCWSf+I70Iew6grg3YSI7
hY++booJb6HQCaBMrZx5ZNJRLn80Tydh5ZNIsHH7UEjtenXhc/Y3w1UJeP2+YlD+8OCMCDoZwBnj
XJuROC1CG23s1fqFQjhDR/N0mJJFXckQdg8dxve83f5v+lVtDTTEC+sZaETCd84+rn/U4qbN93zj
HnNupRZihQWe93yBC045JsL3jH67qdhj9fXJMKLlq9IDxte0gI2emSxwOuoyCvGHVykm/Fmkbafp
cwK7bX9Yd8w9SFJ84q59rpxL+KaxgzXA+Z0Q+FV1seVGe8QBM7/4vyqJv0JBmdaXHPsaqjb06Rug
GHjTHsWhq956EcwKUA/jxekyn9i1siLC/EZTEOR4nUbx4hwab8OctC4HWXLbbhnU73gsi8duSIf7
f8jCnUd4Ab5EjbRIA/uzAOIpojcn0DlyFVE6zX/4uR/sgc4uwZ+O3ryiHovn7fHvwOp1foLBChP8
kWwNTqQ4q8+R88AMrl/vdYXsv6mJxFxkYmbAyDN+rW6h7QrumqbH8qfYQIMkVyni84L/hSb5fdFq
9uFi8P/8C+pqHyQJzKYkCdp7OF6LHHj/6eswl4NCs+OXu0LGSs75d2A+goYtlzMGJtdg+6Z3mbKR
sPlJ9piDq4tV1H1rIHuMEDzl87HFBxTFsMibpmWBlKEhQ0EJkSqMjsKO1c/3UTLvcAPEtQCOkwqq
jzuPBnOlxweOWfcDMmOTQ6IvhyPE/Uva58zR6BhrXi4IAZBDrOObwJPbAFQjEYdh6LyYaCY7okgk
YE3p4iY3jyVY/jO2wZmtwu4gRf5Ti3/eVd9LCb23suyucoModzZ6XWfmhIQ1zTgm0lYit8JLG1DN
GTsDbqNKoZLe8VGmslEKeRfp8H7aDVFEmd8H9FPM18S10XUSsKeM0KMOPUUNZAKD4WvUmpzX+kht
m4eIGYZ7GRj4+w0Smpcd+vHpsSXAyYre0wQYFSIyRy1sT77P3ihc9BvP4LVt47nZaOHkzCSvHbEw
iI/Ga1UscgXqdurR+BRMtl0oJ8OjsLX4Seg+brx1r8Fjkx18hCEkvKB8XfAXosV1qhuKaetwXGV4
51/0Onk+MzSKbYbwDtOyaRX6WvxO+i2PBy8HDnSvLh9Uk8WPnx48vmOSVbH1tcbDwZ/aLmri0QE8
aRP/a9hTRgt/7Whr7CmpsbPS0lARnyCUeadv5+a7v6W+bCJGZddwmKUV2nYvIe6gexPYkfq9v2gs
s9HoUgiNTyS4KX0INsdHBNMojFjkPlmESEULrgAmQu3+ut8bUJeIITGLG0wNrnAwuZWgCd86C07y
UfSfYUzSGqlgRGuRokLFlJ7CWfov8pYrRRPM6112Ko+zfrj8Z8U+VFlvzqfZz+J+cs9JuTd79khi
1akUz/eCSByOQFSwsC6AhPIOphpMREWixbgVrGjINQHXxCX/vD/UhzXPW/oUfzaipLAAdT17liWL
/Og+2BFpJdO1euERGWSSsnLGFkcRnQsw1XynEgt/vlDpg7KQpcXzx1dRVSkgr9N1Tz+Ha2kyGIpe
IjesMmB1/VOa2qRV5dj/CzplOJq3JU8sjWdGGFa+nubbohsEpJAVT7kRiImtirIkuGcqXuG+B7jw
Ijq8Ik+CKzAIABuo/9JNwEpxzgGtjjLvGIxLx9T8oEuW929IkKfQqyl686VQDRfhc4l6ATeC8rqd
XvskQUP9KqSYO3rTb6CPT+TCG+4raqPzeoaxTRi7XiwHFHhBxWbmEL7jZZUsVXiE7YivE6j4F6Qw
H6PLQhg+cuc3QzxBqWHxDJjI5D8M1Pqtf/kJ2xI/FBhHroVKmdcM5yK315vzNQNw7j5yGllB6cyi
9CeRtrd2X5NVIy+zW7u8kU7xsKa2hsT86M3T8Vavl7NMTNAbAb/IBuxaixxe7/xkAEh6NWLxMehB
aTyDmg++TkTEWFIxTJO/RUF3Dz3l/CGwAB+bT3FTsc3DG8DQBSTwDKWEr92aV7wShAAL/vw0bNzs
e3K77spbtSZPe7Q1vfUObZFOWs62OmV9RIhnwdPzfTZprOKGj1qc4Bl4c9VDANYOzioXRDmPYimU
+tXNWRETQyeSaFRKveNlDrlEMFjOZv5ru4rGkF2uiORb3V88da+xhY1/cPzfMKN8mypDPGLiL9qe
bxLSxLSwI5J2zNbWkVlKlquxDKkcQz2telo8TRLC6J4Kg5rZANGGQvj4W8U5BVIWgnFK34yK2k+S
xyqBH3hat7Cq9yhJll9BPA5eF1MlE6ReuvZEGNWdRiKwGMafVHnPz2ViwfoxeOevmW+nN5jOtzv9
qZ3nNFwDAvnhQrzSWYEQMikGBqj2iDHjOwKjbAweGYN3y+JO07TM/tLInnVvUmKvJgpTzeJFM0qs
y62+t4OHeYsBC7pyJZLUaTK17U0ndUk23T/K86jtyG0I6o40lLt93aqnolYep47knqlWxEiDqvna
DeIh+X6BDGzN337IXD0J7DjRQMiwVIiduG5zfyjzBKC+ANh46kCIIzVwspuGgSES7llsvjM4mNdE
csHlTLo787a9j6wYwoinD4AmvdM5zIMA+HfW+U6L53y7aIv6qg9DXLc+NFwD9rIr1OE209MQh7TX
n4ggiFmfujKquLRewSiqtgNSqKmAU1fecTKQEkj9659cjfS3gH9Gvt79SclhuD5nV5+spKx5eo/a
vemGeHq4Krwaj9U076uoNEahA9PSAKu5kSwKDRQ/NBjDG5j1yrMJSfvBHpfwl3eUmUHopaCH4joA
1FguEKyriCbUkD323wtceN3EEKl424kJL+FGcfgLlrsGYxgnpN/arPjDxZwmcSjzY/ZSIFvnspuq
TlPo1vv4j1YJeWrtF8MQa7wnKU9G7srmqdOkmkLijif3C5wbT+oVyHBEjHhNFcGRPVr3eEVuc5jF
dlpfd4lrMySG+6CJ5yVoKl5ITdjauATuI4qMGuNqfnlux2ctiSYr25a0N3QxLSqOVejW4gRJfUdK
+E84sL8Y5XTX5uKzy+d8ETXj4yXB4XlwJgltdlLANkPz6yatEunhS/e1KBCW7lNiJxo+ONjIuaR3
7IPFxJdsyEo1x47EeaXLC1ZfYRp7Hw5OuwWoIawuv05QgfjqUu9UhOeypoZ0HbuMVp3JsxwR8wXt
ife1luU4aEgBmAlIhjXuWDlS1f7QWlrORuqUoLnJR43wFECnvlG/TT8BQg+p289QLs96REtYbsh3
88L3NGzAoL2jJsV1Zmx6aMnjP/E8H/5FD+ZaEIJ3a2DfmUnJb2qvkBTg9rpqEnEyp0dnq5turECa
xt9heCv7G1gFbjeqKu48NBmvXV25Ltv37xt89YcwxEqqGLU9ONWo5XXuVRCMw++JnoA4ctVtSRSK
E3Xs+Ti2RhSoqnAFribTo+I3TB9QqScFeGnpgCAnzNp6jURdpHW3G/xrtPrMSTghYjQaIcafdvD3
wMSE6hDvvlqY0BwJWzIPl4reNw1jnfsoY2Eo2T6HHntmn3uwHoz/jZgbddm/dVLOnFpsV6rsPXMl
eHJh5rW4CkQPrj9/8QUlkDSheifk/w5pgH8GRx2Nn4IfZ5wBodclQhwsUOpI+EYQPJ+7Zv5HXbCO
oUMfMGh125UgNpeJeroODR+yIn4V5r8kceYFFTQzti2bXeKr6tcvcd6ar0J9wMS0F6Y9crxB6WNt
ra0meHA4m+wAhvf/2HkjBQKKvU4ciwzu1tph9ZhBFtw3qJphYHzlooVVLDon1B1RP+MdjKq8/J97
MY4hHvRxj3/F/5SaGZbDgyLjWXq7nuA5MZE16ppoqdhG9tUnv4pLS26s2CQSzPgsWl0bmCevQgQ9
g8aRCmE0p5VopVoVlXqe0tkyArUIWWoxdOmxmiDYrJ144Ob0hWCf1nVJk5fG7hcygecS2tDscLXn
bxXTvtdz9MkHFXDCyfz+MLS83ZuRoW1oxvkaefUJibKkoTGifaLU4QjzFM8cVn2sf7+n+1dIdbYy
XwNB4K8PcvGHo/ykEGfPjGtasGHOCUEz5MLkv0DuE28WAOVN1EEa7j+MMglKzylvapN5RkOxMCC9
pLkVZrIatY5dfwNoesHfFAHStlgS1MibdyZI9Jis3DFl5pWPJ7n9U66E8qinhG8jdhZPLosRnoVO
v7BS8pEFHgPv36fbsZULrkD6TGjShA1j6FgAM4O/kbaYbrj0V+3FSC1+YhgH+pxsDxmOuJoE+TME
VbFsrl7Cz7LTGSZRbMTwUzpn7o6vPx/knuqt5fCHcJit4SE+J0uhPxq0qiglpiyitB3gTNyTrtAQ
nkpcimu0t0FTDQQ+MGieI6cVz8t2UnNaztfRxoaTPvdpGvGSzSXSYmx4ToM3d0husS86Qm6pifnc
l602bR40pBAZOHyX6vKp6rpnW6LskgN0Wx5h4qIidfMhVT1QodgyMLwTqTbiX+UEB3oyPu+xsD7v
PiS5dCBBpIY64MUAoMnvx2W/mEum5ouuwXm0Sxh31LCQgywLp4veE4z555NNttxlKN4Mi0GbasGa
/OSg8/Z1niFP9F7kcnUtHYp1N34jmxLI5mhrzgl27paPQA9sgXwG1EyXcNmY1KW8w3wH4rfAB1lV
f8IxlZV8l6C+hX9JEy5SECQDeiZmUCq5eaB18gX/SuFA459IDNOT005llxJl74GO+y9g/WWKWLg3
tzh2SdtOyTt+QY6v3r8VXvUiavPAcHBhWpVMMKdJyE00kNhStHlaKC0T7I/hd+1asCyPAQXMes4c
qkym+Il/+NA6qGYsI078MEA/pK3q3Bw/vVPzwV2qXNwmq/+r/gz5Y6L7vvpYN1oec1l8v08P26Ap
yTVzq0eYhwe6pXD80DhUiCBG/KZ6HCzUO14pvutkgtftobQ0PJPI6r5kgxKaTRg21s00u6dXGUcB
Yytswu1Tw+b9QHgkHdPD/lFtkhccmLxRAHDQYE9lOB/g+YGwIujjTiLR+LHEqbqP/QX3e/MLEL/L
0xhUSvpi5i3RsZyqu6bFChF3HjtcbRm9pJEGxi2hUqdUcCjwmu7GLMz9ariHuiKR6rIP1q4pWKBN
4eL1AfV1h9B7FDNqBrR3D8YoK4Knvh03K+bobMg27luN27vlyBzZLI4by7jJ1NKl9MoMoStbt/sl
wQFMX5U52JKg4p4WpYTgsWzWN12o5xz4f2NziGhh6WvE3WaBCf6zjDi8HFGG5yHo43Z1z6uMTl7a
RzoRNadKMWWx+ucKZwoaJwgDN7qbBtWmZzCMNC0nH9vkmK6QzQnNKaqJpgkyj2yX3v2rK0YfwFFS
ugyFJY+Zw3a7O7wfCG615FWoheC5FFd93vswCnKPnX1pHQRvJ2ApSDBqnFabCyIz9Y1OLGxiiVPC
RFoSy95hthTH74op4vdyzq4IR6lNA2ItXw/zYjBT3i9ORyvxz+nEvxMPztfz97vfVCFatrzKRFzB
MqjO1NkDLzvWaqpgWtPGwoKFbv7Z0vQE/n5FAVWlQWbVbX1YwXTwCSpL+fPX1BLQEw1rPQCvMxKv
qVKDVEjyrPaGytafCRM1upeuJNpO8Nx18RbFFyq8FhflLd2rBYYt3d2fAoVfTLf+RLAEPbhLTKla
uWQztUYIGwW9HE+zAXJfh1ZrOlowyIzt9eS7go/Gw6m2EwMlTk2muWnQ3EmzwKUmtZro60FL6bO/
NEvbID4RPRlSvxdkk/8MkIIx/KlFpUu6mlNRLYtAZCoZE+Uu7/2H3u4eyk23MZN/90bzyelGN6yw
GeV5sAss/g6HyJ//Ecd12WOcHP1K6IHapL2c8yYr8LJQGYo0Q7qfUhhkf5r5JnIt0Tx4xcAFycEc
bAtAYpz5rcD2ysUuMR+NdzO7zny+XCD9myw/WU3iMi97ZrcdbDaISRXo0909Rn89otqzmQrMRaSm
bgapznX6IIcIExiXgyuBeVXV2LNP97E4M+RtzglbjLXpYb5kdE+IrnmdhyitZ2mC0LyccjonqX18
sEF5iV5FKyKm9AEnga4tjUwV0BmjImN9Q3x67IbR/NzYrt0ifbKembadyFYQhIYVQzL3b/Q4EboP
FDvzQ9pSRcN6leSChI3qMe9hJGwqQAKvBFpLb2lHrVo1topM7yVi4so3Uhjr87B++Q/3oHNJtemL
8Gmt3zJir/w2lVE8OT1SQXDGZrdIvAOluABliG0nnIXYBaKpfxQHALRMh7oD9CfUuqV2n/SHtDss
4X8kf7BYglFyJxn4WTD0Go2T4FMZJmfXMBy5kcsMnoEjSfo46MkgOSwnQ1G4htaIkuJyZOcVpS2u
pms/hfzcp4hDD0fFeeWuZWfwtSErDMPRBYwICjQE1WzAoBZADkEWg5KTNV0qLqeqFlfqjyVym52v
I84uOss4x6IDe+PQr6sc8DsTTj3dRtnTP+q2PN53Y/MQ04MHSFQho7ZbCoPv9iGzCzJsnZjMzo5x
pc92mMhQJiIQIY4IQifV5RvqtHJq7HJ55yEV2l5I3/W0Cu0eNxvNYw6TFQcOkT9g9FoQ8itnH/rz
gGQ30VuLPKVaidSBjp5z+GST2UE8MT+eVjEwVzPzUznguXQOwPedZqiywYrLAvBGI9VTSAKCDmB9
aI6h0EyYa9kppv4+ZEnDwlAuG4hLck40nA1wUvuBQ7BMUIPnnx3uluJlv9+sUQsrSvszI8S1hseP
50f5SzNmurE5aAX/2knC7j+K7sTbG4xGH1z64bFFsoNGC+huhr4SsYdzSJZFVnb6UYCakJI8VNGx
Z70wUWikINel3qIX/20vO4y5RxgunOY0IB+XwYzJIc6jydgPp3GYspB1a/jqXqe7MZhcnWfNK9PY
OSuCTyMu7EyrcMXkO8YhyZjJFFCpeu3+SR4zDysxSZbQINsQ1B1Wiyrt8xGLjMXKKaWVyS7RjpGl
ZrVy1TW6Fbgdw9P2ru+aHAixFh1CORHo9aYGe2YaDTVbkA+nPhjUMgy64vgDfU7Z3U9qs+IQYoGb
JmnMFxgFwu0sO/MpR5iVdzLTyK+josrOmMcOhnDU1nUcw5R7NwWJeSA/b0yXqzU44fGoGreTvvQM
iY/bfzfJhldbm5hWrnlTX5mGIFPanH52qu89ziNWgf2zEUlUMvWlVCnzvvQRJHZNF7NmXY8xOeyc
ZBVyxt7pEEQ4pI8SgYfAEPlYxYOBmHfUqz40G43HRbcDs1kYd9f/8UVQa6Ie9Yj+TBSAhMLjZ23V
mjI8CzhoD1OttSvDtkDHTlRWdmbnj7bVU927PECTpRAjFq3N8aSY1nHKE9hbs/R2EsxBT6ogPo2n
lsfujgcFyKAPPXse/tLVHwMXSaJKz+A0Dqc1V2ygoqbUT5zKTLaaEkxoD1bJKknCf6ja7VDDNfpj
b5Mrs7CfDLxjreZlb4ysHjUf1FrNttRHCKnsVQiv//rpRV8M82CdpHH6KLKFvLUz+qRzK4J+hEra
ov4iQn3fiS8qUWTcr9A1Jp8xdB1lARgLTVN3ooQe4B6TNSzTduD8ibhCRq5pKKilA+Bu5YxHtP7v
XOAXft+JQ76T9icLf25AvJx+R1GyGaGRjudbJxX4CT2+AJ1E7ItPnphXNGZDd2/tP57Zuvcmxu25
zXnh6JtoekTe5XgHtap+BEaXnvklZaOgpbE2ottaH1nkmw5pPINdSdaQsun9dvw1nHBhk8tn0kXQ
zd3ZmNxqLMX+ie/P4u4ySkPJ0dzKUoOnhB3b94gdDI4I8ywW5oCAAbXf53L7ML8vYbepUeSly02h
FFIeW3pTMXJuetQwaBTnsPywUYePKGyy7e52YRCD38NMBBrbRCH/22gxVqjSXU79qt18mM9aM7AW
DIpkxAbASrSuDU1cTEmYenvvYt6ZmHFkcwqEkl/Bxa6/cI2e1NGNOPd3NmuBCT3jpNRLIx3RMrcu
gar9CmxkZPuMC9mqJPTbhMW+wqJq7QgpD5GUFyy0Ckz2iJab/vd2LLB3bB+o3rXIAhnFXYqiaNdd
XM/m/gOIuMx/1ZZxLGYHHorx4Jjj3B325GV2FBvPB0CS/HL+1QHEoGfX4GcLfyNFzOlVrcQlCXJI
ibtIyS0JUMWmsG05LcagZs1GIcJYz7r+exj1PD7bQSDogFJK8yd8Eam9LeQeuLAjJJy8tgNW0HXD
axoKuVY5i5NyPPC0A2fWYekPVnWtElWjdB5kHPQWHhprbiTq0JbDuHsbLoXD26HY+6GbafIPevtE
DsMdCImF+uTniXKWmHdM2koM3sjUIBtauDAhlTL7d6crsjxD3J/u9hslfWlGRFRokRbSWhpOGyWv
EN8WtNrNxI7amGAU3pbdSf3AurPhfe+A/Rra9QahbqFXWzfWjh3qhQM+tTMNN9SeCbdCcZZ7uevc
VyXU3+4LkHrV+eua57QnTAjF6Bl7MWms9gNOd10C4C0ZGImZDgoH33hKgvdBlDjy/yOub5vKiiKk
5cae3kgeO7Wkke7RVBaIdi1tbtzsXxiRup/RnMmV8XzROfdBgUhjYhpAtqVObnDE7BFwANoQujPC
trZDcBA4xAtYF0gI2SK45u1ACj4BWSofZBgxguhfj/nw3App8QkpQ3lz+wxmgvA9o1ufEuaBDgRu
u1vnpu5H44z7d8+l3EZfcTb15IrsdAmnWW2A2e3LNfO2PAYzhKkHvKNsNZXg2KGhl1De6lq1Rm66
mxkHlR2tNDvJBY9jdCdEp6wJRIyN8M1ZV0VttibUtg24QdVhZfuc/ioQ/o2cGBdcnqv3Loqvmy13
uElnFyIFAxKQF2f/0rD/2xFDqgRO47YxJV9lz+Kg4OLju7SuuQizhdbE/GIar5PrrngYz7c8LzGA
tiWsyx1YAAh8uOzM6eC/Qs9EYTAahNWy5Zd8exPKSxvJ1U+wGavh+rMI28fL+jT7RJ67nxSrlG0G
/LhjZgircsJE2Hy5xz++QNs4q1KoW6/Sjbj6GO0dhffzN3XHx/NfUm/ROKbOGHXLbxfIlLU1aKjv
JCtW5VcvhF/9qBSl4Ux5mxLwBDlU/ka2GIBV4gmy1Y6tEWA4BjENhoxfuTGocCzstMnZuoRH/rVo
AOh4JQPmYY4yOVdvqOaRBWeY4scVYWfnS1H6QDCc8qu5y7+3wGwHOv3/DFvaef9cuCBSOzYFfeud
bBB0qQz8LOQwSXhLXL0lBiCEPW1tzLUxviweLDpXCYYm6fdOe6iKAWPIurg7NwY9mDBjALp0m1sS
Ds8ROni5wPnR/Us9HikL8QtLsXYRXr05P4NA+puSp1FiDIXLLnLmgEynPSe7iw5y59vd7125GhM0
eITo4W0KPx2UGXJFjTR9055Gc3NuZoXxsSqLRWf8V1bv+W7bb0axVcaXKXPK3F4FhTAfqxdMueHc
MF+NrpOgXEy3ZQS0cxWQpkQ6iH0YUkiMoq2zn7RsDdhbYa/anRyQgxnCYsR0Vf4h98JAfpLpO2vI
ZbUgjzebPb481hlxlM6RLsp9tIMbB7oNQsvr/j7c+9k5xo1FuYG4zLHZTyfBtbbvKWhzAUxfXzCW
Rg/WUyTiJSNrUxalu7Lw6Xuw7VIfyrucrmUGFz4ZUdmhUJML4AxLQvDH3QyRkepmELiqTzG507/B
xsnPCJ2Td6V8kURtpWSj8JkGCAWFuMNMcyt+Jvh8drPK5pQal4C9BT4IEYRILGTdgehg9BBdmUOz
exlIDNpAVq0tBudZUyuMUqhRjgy9vrug7KOn4ZsQZql+uk50ndde4dOEFsfIUwV6+tTXrYt9a3PO
4k87mkkW94O5hkaZEwOpB7O4mK76SO1byjGFUv5Bdd19SqfGW+xdeRGlXsyl/g/k6deXMSs6J+fh
zmr6DafnpM0oFd8023sngVkeZgoC75j0LVbxXFMSCXxXzvW07dbdk1z0csLEFdoo1jXDqKKLZzAl
m+Y/MOTC1G7FMNpsfqxjRl/Y8a8P633WkXZmoC4/QePphM+ew4JuuKLOPqe1ib722e5vBOMYtqjL
j8E6ViKz8ICD/pqhvj/cMLBNX63ws1ay6bRTInCHQ8t720pAGA2YnP9/7lxSFyJtyn6PaQRnw86X
7C5QLOJmXmgsV9r5S/ZebrHtWhoBGXrI791u2Sa2vXKeKiNSfg2sXX7F+AeV4ZdBGutdtDPgst28
va/dE4mWnK68UJMrWH0EAnJwBICITeLW+ow4ny+7+RW422axpkEyYzCPhjBxCUQAK81Zp5+jE15u
QmhW1aLOVU4CVlhEg885/g5vmOw01LbCyyjqVWSsHXB/GpHR6s6wSk3wYSimKrwWoWKjjFrl0uTO
3g6eqVkMkP6hfgUdLTQeZGBt42DkVnjLDYzO8GzwR/06yp1k7Eu7A4xzeNlS9xDSdKKOlL02svRH
W5ZGm8hMiMAoVCcOCyLvcHqv6K9/GtlhF2R6DCSfFmO+SgQvt13VqNVSWDdJpT6wSjO3L9n6f2nx
nvSKMLu/iGP6VBfGLxjW+1hUNWikncSzql6g/EWGjiKmXhllFC044cOhOgX6bgfe6WgaedM1BPHO
PyDaVZ9pbfsISJYLqoZCKOQvbdtgzEwZyBxEuT/qiB4wOoRs9wkBNTfpv4aQZCIMRXNDdXrXwUYS
lFTgls/waRKanMZ4N4eDsRoUxXXczhSU3PxdT1Xfbz3O570nOAFR1yiWERNXQEB+esLeA35FExCK
2hX0U3Qu9DmPC17lmb2HnD5R41dw79KlKzN/AJSAWtYPQc6/Fe46Ee/P4xzydaYCBdpma1HL75QU
tXQjBQcBLiTRM/LLN0SX128Z0hVPAxYtLGsoJWD08xU6t8ZdjiCN+8sOAiB+Zn+wtYsNXxK/1sBy
52Ja9LWmordcILkjYiwl2LmoHlPQzUYnstMTi/IUU8VFt58G9Xy9Qxzx+NXOzvSZKZ2tKNjxqchS
D4+yVAcaWmBx286gfxAWozL0f8Hkr70hQRvqEXdiZdF2pXf0mJHfp7HsKZCROa8EEvEcIItYymeZ
sCpH9tkSHU2YhOzjI6qy6e1n3dwP+2yKHwCc5SYZjCJ/Oz25mapI10UD+xDLUez5wH/r7Ge4w3vR
kAXejpvtybsKvbxiHycjSVq736IcU1ALPD6/6M8KDANnb3dTGF6mwkZvXF9987JRQsk31/uM9adh
nALkfViSR0JpBuggPx9lkyU5cx80eQfupcAXRPn1q5qUUHSawswKeRk+SzWM4Giv2wALWhyQ9O6S
WwjGICEyUVAUeh6o/yFP7pKtX7jh8wPgJpduFi9KJPO2TymbpQ4q4LFRj1XXp8eZhQJU9EvxovFO
Iu/GapSiuwWlGM+o0wkXeF+ESJYJ693TVVq79Ymy4V+Y7AMQPQFCneT2RO/a2t3CDo4aoSW+pq0o
g/zaIAL/TqQSWx+MMRCSyXORs44UerLSok7lmS1Qm/mgezNZlyuHHrrNodSa797JZSpM/IAw2glT
WTNVR2tm4KhfDP85C/z6KJ2TnTBK4N8knYc8T5t4vPnvbnDBnpqLvRDuWQ+/HpbBMoKqnzzkyYjX
4V9pZJTBbfb2S7pEqnc3nthiJdkieVMG0bAw9oy8ivCHY9NZN709zmAqymAz2CEwLwIscyzhFNGX
gcyMQUQDkAQKvT7HdgOL5PgK18bm9q0lfBiaz2WAPmWNPnUmGkz+UXKgyRqGmMPMzVig/5/V9iTt
6kIzJFuXLxVADRLDmA7WNbDjxeQ9d3ROVcMDbdKupb2NSJU5prhMgje9Uwa/2m4MGYAw169znJ8F
usoPYPhtSWHuKa0/msUnHzR0XDvX22PMTue6PSLwAsGmlnqjQop6iKCh6B+AB60NmKAtoclb+CEY
bBC7Lo14RNXG2o1Zv9166BeJ0NHzSSGsr/UGTU6ov2oTccTZgwh7GEu8Do4HBuWgWLgHMdsJUoeh
GLM9mpMFSauWjbPETd0c4Cx5OaLU5qy5wmsod50Yk2qFrFf2J6X/lgO3HB+a2TT7WQOLWqn2lR7i
q04S6wgGiHpMrW0nlFII2wC+MVKDfL/VMYYdqpgoxd7lJ9sDB8ydYQXPWRJifd0/J8exdzin1vFd
jG4yKQdOU4Y8AKCA0Zq59+uleYqUdFgo4c7uWMSfiMrjCGGPY0DQlHCGrFZog6peTHk3T35wLpb4
dSOpMk/XpdzHA2lAQyNeg1fXz3yIRnbMhFiufkW3AjOguEHHp4AasgiJzSC6Ki7TyBSgsfuS2ojn
P7BzTDaiLXT+O9qzfHP7ZutVcbZ2DWNyn4D2DjR5CIPNBQRqCbwU1WroIzO6lubX/flbPqemFU/v
PuhLdxGEXTa/3A2Yx3ZAXtiCWxUrBsI4+qN/8d8EdCHOLByJdUTbzvBdMm3z7QexBp9YdErQ902D
g7qusvLCPvKyMZkq5LC6bAPfgvDxQCVEqr0d8y0PYyqBC9oMfk4lVLurDLjjwzoHM2cz+GUp8O6h
ptQxXznzj+4bFDKsRlEIad29YuG111U4Oik1GVnsB1vV9XVpr1P8YDf7ZtI4LNlWX9EcsWKjWW8z
T/FiDHVtf3Wd8NaiktP8LBk0BqB2o6laByD7M4VaqYGZ509+MlEtDSITgbGraQrWcK5rPIUAxYVv
zBLs1cME0DiRsb4aMXphlfGZBI0KQ6p6WM4uNXrw8rB1NsxS0mZyL3eYlYae4NmjxvG1o9pAT25t
NSh3uCm1Vukfyfo5/B8DxXjhRfsfxXEtw4JuLFmLCD/6lbay8q7ddl4u/ijjTrAm3dQLsFb4Apq9
rUIo1TBtXKLBSrpnqlynmENuWSqvS7tcTra9cG0dP+R9DJM+xwVgQTAz3j2PiVq9xcM1KqEQDCq4
5dvtB7O5ZD2U42lq4wMNjaCogo/LxlCkC3yl4aR4dzvsYIncZbnWiOOR1sW7hylOa8kXSVezkC7P
g4ZRqBa5na4kT9D4qY3IGZXUJWnGQeQlvuQanpzI3A0Nd9YkfooVn6QYaXn5m2VVyUbXu9kcZrtX
7RGZemsMiiqQu6NkFd0Km7iixdPZ0gjQbE0t1VvVd0lbLESRrNLKOIgmqrgg3V1+3l7KpJtrobIx
/H0vwrcBtYSw75Yx//kriRFRE+kfR0Jv3r/dQor3p1HKaz5nwcfq8qDIesCitxBc6LuYbvB8cyuY
+g8qCic4UYYpK8GHtggTrys+kbwf7DuKS7f6l3fCokRth9Pc8BIARIpN30ry6HjFUinGBhX1T2cz
WI9G3GMWNZAclQCphcQ0CsaPzmLrAq2KpQVNjbxgEqgwO03EIswF7Rlw97hJMAtyzesB/Np9kGys
6CuoknIGuIMwOafhyZWUIQgF7vzWrEO+INdAT31pHydu/EiR5rImUr10nnAs61LOc9rQm+5+cCx7
C4txU8Xhj1U23FSyYL6H+h/VLX6GWhJ74I6UOLxi8GNoJhrnE6tHe3T8LzJs8sM5Ny8uX5HDkxHR
QJfefd3TeV02Ywi/cNRcClMahuCnLSbfwd6LwENqnM4dfz9jj2zBCmakY+qg/DwExzTY+B9Yyk/Y
Xxh92JnwNrrxTNYd+1zLKhgXeq/H02iTGn1L47tFI8Ugl0WS0OfwIOCQrBwpqUHrpcIn5v3fdTJk
Qi1dfsSHdKBvsHn1Ckck78lkuD9BwPYRhfGaxz+C0pYC4FAAeHYbceE/USDcOaHpzfuBpcYfmRfp
+6gYp3rscvfvS3bUGOemUki3Vora/zvRaoEzbvhWFQfj8II48r0NTxk8ISs03SyNv0rsRLiHoUqa
5QLcMSsWPkOhX5mlvnjZjKSa85lXVUgoe5wkcpnFgqQU8movM57B9KypGtm9fFijzyek5oWhwoxA
wk8MUp43725F6tjWgD7h3QN2rgmXqAxxPh9RisVVP3wrFZQd2r4H5ltYUExwFI5n5xa6GdhJUAiY
cs+OlFtvVVEk0dB4c5uMkuDjwimsZfwIjkhzUh+SveUAFO/nFvqnBxLb4TYQJLYpNf6EyxRsDhRi
hazPfNtltsnoAbXFzZ6umcwSjjfdHEGE4BGR7gvXZM/LG2shFvlm7by5ygHWIhYw99hx5zOW6i0P
hAtVZR8Oc9VCq1VEZYo6/D4PkEYAZcQ/GJf05C9qL70dd6BmSjb76MZ9UGeS0FVNE6m7q8MtbDTY
aR/ULOn9wqTplklpkKwtlw7t3BKAnz3N7QsI9n0NUlSID8lpN+jUl9LApSqbN8UBcYLcehtvSZ9Z
EfwnIzHnsFMkqOAulDJUn1sqF8MqGiMpnSn2q0waB+LY2ULqHTntOs6AFE6c+k968X53CKwx7CTn
ZcPoRV/+YUeTC2Di2uHG4h+fXOwlGgeNq7zWnAfoTR0dXQCb28tqVb1GQAfbYhOBMkix5WEGD3zq
wMvJdiDQNI8uOOpwQb0sIZAPj6dDm2WQt4erjjXLWovMblrABimWFdlYB48dvDOGWmp6VE6eJKfs
4Kj6AFmni/I4zbMTmBS8x45DKLpNOHzPGL575YWRq2luYbfAJuWiAiaTiA1HgcTDw7wehfxvuCaY
l5kJKvUBj0cv7OKcxLg2Fa3vWwZQWyKx069UmZxVKrtWITrpbaD8APUY1kp8n+XQ5zKKxBwnmqRK
X2ENFFv+/sU6hdrxHyceuWl7cpW4vYAVEqLvtIMNQk5a/vc9C4CMbcHYoNa8oQX8Hh0eVcPvfWcX
4rZazXiE9SQbGuZCXoUgRFAmkKwPTuTxP/jno0oSl107G0N2CH7MVwOe5JFGf+JrxtL9dRqNS7YL
8UO2gIGznvPDgRlBvwftOToUNY//KxZrP4Y24YgKKrTO2GNzZ25KWQR6s38F/NBd9+lrwtunnklF
ojWDmaQp6t95ELjAJhb2+ATSw2hrQ530/x+cJXEZAIn5ysVsMR0CATzax/I36/QV4uRPvv7y5Wdy
RZy6bbIkYgY5vve1HfRU/SfISfA2kx+FRfZ4ukcStz0jlJAM2BenAPOBNhJXkKLZumkB5o60xw7h
5qvw/Zi5JULkGdN3uFP9PpzW4O6Oz18+yx5U/An6ELhuek1kpbS5QJEY+SiuF/1KZlm5T2eGnI6x
2wMlLwbniUNomExC66sWboWcvmX94aUNRASZMwEpTb86eBk+wFSBjAmdf9jfNWfWpYxWtWzgZ+9y
xg9ir3s1blfDe/fWqMeb+VQR44XMqKv10QQUJm8ljv459MG+HIyhB9IO8P+FEMK/b1Q2LvaJ+ZAn
qFHSUnDnCG2iNzUosyF2QNPhsYjgYeWSZD8IRS+gO4swpyxrvBfEpBXR6G4sfOJlaDQIE/U/+Fyv
0xpIlRGCMMm5f9uhoh0AREhohhvRt5VwUn+hIfFh1zPiD1+cQ5umLTQGPPxD2hWgh+cCUgnkn8aK
Lim61VdomMhj7CuFxsRczpIU/f26bh+t4iGA3qWsOGiS28JJx4Szo9rYTrC/+u/vXG8q1fu4S7qP
HMObBhyYRjKQ1SlYJhly3mSuCCd3zro7/thp8pgSgr4JNfY0b5v/MV0rFaWg+Uvwq1thRcoTg8en
q4f4QbX9UF+SzpZQHO4A10vPJCZc1CMoRvkuzCP8DLTBxz3DOCGaMSCVXHZBrSqenLtApVz3Y81o
HjB63/QagyBKknHFEMxpWUPJIsxpKBo0DzJzh7gXhoV7qCCJa4t7JYytMCghaOmz196Qsrq/3dlH
T70ViWFUexQo04uCZJ2ylg5u8ahqaocH1Xth5MMBh688Y/6WJZzjwkybDcr9PzBc9J4VrRSgOKO5
Db9mbCRYMY9cojOYQQ5Gt0sb/l9CSNW1X4O8mswVQ8NyXICxMswTPSYgeml2rbI59dTxopK5rOwQ
pCq1ESSucufep8kWD2yxIbhKYXeTfVXCJ5F6uUr1NIsN3jRYfJGjR8CTumnNzK2sGlRFZaFoY912
3NpauCp1rlK01/90bfffFJXduk1YrtC+iysqYgp3jq8ZCks3FGi0io/42RND1R18fXY43Jk5Ovbk
sgA+yEOc+INIISdg0MvOR1Eo4ahbgjoh83uRjbCp/ZSfMJdPNMvQC951w2UX+uaAraN4gOSoj9vK
Wh82LuEfhywD7PHW3JGiuK4nz4G19AvaUMtH5m7XDIGCeNEiLGHFquMBxQX7Nba+/c1ZLOmf7pSV
SnP3FZXnaYlR3TTn96H9/hUwEwuEy4/+6ZUSDKjCklL62QqblvlkU758MqShAytladL9mQFVzuoY
iqmQZVDOjJM+JCxHMm6SgLcQcyhSVvOwdYaPTG+NC3mFfN5fA0c2wpNuMvqjCnbGXzF8//FfiiB4
42YYh+Ri0nNSZpkA9qYRKwHQjVCqKtQXaQezM/CJfPUECX3nXK5mdq+1UaUp6CGux9ateqO9Yuoa
Xe909xcdy3G7qsWxfgF+6I0QerxTeNr/nT1WSeyxxP1rw0CJBqzan/tr0p09UgsKotKfWV5M5tJc
5UhtFRdAwsHCiYJLajRe0MfCY91S4dRwvmNjfOXWXJN8TnetRuzb39SwTyJjMIcBHMZTTjPzhPjD
4fscqP0wXtN7lScxQfmrRaTdoQP0HApDsPG9BCnxIBBCZAYbSl2zemUB6DrkQogC4RXYqWuJ/9Je
liDzlKxUCacGmQ2LXNgNDIw1nCuZACUxR05GXf2UASPmNlMgmBbFPvrW2GHMQbC7cjEiENyOvnd5
FUTOfRR+JEgkOVDYSM8kIhLzekMcC2ZPvU2KwSeXniMC1HGYBIU4giNTMAoesDjdqlTnj98I+W5q
gSuoE8gyyb21xxMKaeBbeCRYYSjORJcNW+HW9O73qPmgyO5gRfqGMXZh7fUkjzjvGOMz6kKwaTmL
/6YgX88bvzx2eImfPc4P8vHaKfU+cP2gm6GTptnilX8ByO+feRz0C0cXv7mMdwJAifSw/CRhgaXd
sb9kLT4kEiKeWLlaYQxr/9d43j5e1p3vWzC3rjx6Qna7RfiwK0stYbmpCP+QRw04clHV8VUnN9La
ElprYEl7q+bNkJjQF1upnL3+DW38ZDuTwqpDWhEXzcj4Qyp+80bW/zf/enMqE6KiPnwuyN+XRQjc
hGhcs+Mr+jaW6gi/98azM4Zhme6jlo3MryShj6F1yu039bHNn5GFDZSP+supU1bXA1XAPaOTba+0
nEi7oUTBKKCIbMLvTJtu03Ozfg/h/JlFaBJFBsq2/tVUWcjyWYfCtHI0ye3od/81wE663nRxIbcP
K8jOyHT0ieF0LnYhaWqYIi8CZfWiUzuAU75g3Udw4ODmTnIjvJKp/ZMPcgAh7XsbsUo0jfUzxZ7A
C+VGjkOej8429ullAmDZQJfxJZke9povx/gbCbD29OpAXNj8vxUH+od2K4XXxGUKNKEiJx9TucgM
Nd4MATS89MjjBc1nQTt/rXAoAPq8M0b2ZPxDf6uX4yF1y8mzkgWCH8qECBe7yt3m048S+P020JdS
40enaEHzrExjsd7WnhXOBQoxB4T2Kjn2sQ4YD/1NKGuJ8UVvUJyxoetTS3x7/dPahqULR2WJpMbS
foFHCoRK/X3KdfHmtlAK5Gd+/MRInS5SuCweTyFIC3LFL2Lqb3qjJ0Y4jFU+fXlQ/oukPwk6tVIw
KepIB3saIRL3m6tPvvS2kDyj34CDGBSHNzNDR0O/G89o0aCSe+H5weP3kLtsbXTmj6hHStH22k/e
QSMfO5q7om205Df1lFRd289zvFMWcKemryMWgyZ8JJjWn6fynwWh4CR5rvpRWr2tdLF98/UWEKU+
++OXc4lF7W/pTlRTfAmfMr0E/U/mGCqU3SqtygTI/M2jRaOTh81yw+ch2+pemucJaNN4qDXDC1bh
uIknmPUjEkLTN/aQ/Zed4huI1OzRG/rRdfy8cSfh4B6fwdl1qxz/tw09anem/gLcLYY0sz3WMlGC
uTppBcE2KotPhUPmPnnT42OzOZUZg+QpkOcHg55veCvU2qDkC4tyeYdufDSbvYBZh9hyI+1uonPz
d+Mjq1F0Ho2DBpz3CrWnZc7l/+YTmijTeyUIxwDmkosxr1QtYuX305yQ2N+3F9VOkzWDDZXZOJnN
4hOf+QW34se6h5nNjYODm3OhrLdnmiO51bjiWZ2jm81yO0KRb/MeWUIeIimEhMKRPmRPFTqWlrxM
zWYAzsSwtMFzAFUoeumu8VklhquThhg+kWleZJU7SGnDd1fZnZAqx+NbIZ/UofAI9V8vjYdZqq1E
IDMPdaRWlDJIPRqPKJi9QZ16Uh7BDrXhsUyAfQzlXk6VaNPtGfCuiqk8LilVOKLVtHn7fUzeUhdI
iJ9VCh6Uul2XZYNNFHrn0Kf/W6pKFSH/M5jGlMddsl1MBqo3+M4rCECcX1fOStkZ/lc/HjdyFv7r
odIQYhmmH8zQDReAP2LVW+VSfTtIAL0gEMrdjGz2I2UZMrAy1J7cozzlIOZUQRysLfYYbV45EYS8
Qgei0r1Ul/+Sgb1UnhZ7nI9LRmielA4dBG1JoyLc9oNsayCCU2KPyOjaqTGFUPp0ctTMoRzBS/TS
wqy8O6FenjvgU1XIldimvqzhA380BApE2EUlsEx1F4tDXDBWE+ph8tEp/03zcLbkpC9PuSNsovIk
iriEVgEsxcnx696lkONMNWS0sBpqQdVzSUwnf3ymnwBRtAbydTrUMMmYy+9shgI2VFNF4cB+dGqB
hggqNTqN3carXOKkb1sxI5Ot2+kJgDrYTB2wrrtbJ8bAkMvIEImE8vRN397kawXSvG3cwaLszWCj
t7+38I7A1aJYBRhIt2LwnI0dMKMz6g5npSyXqll3DecqSv5qJTl8qI66y5FNKrOQoGklTNW/X7cT
+JdnQTZi91tci0BOnb5SwmzvooJXjNz+4gPpLEEa7VTTtRZTtkr9DP94VZBW2S04IPqWxnZpVkaD
XJSI03fO3fmCoGp3wS2LIvH23s2gOVy5/d87cEnmLOjv+HqzpDr3bkc9sEty4EU4GDcG0Q75zvuK
won+zWCy2abXAGBpSswWH/m5K2WPzRUWlPwBHHND4X0Y5FVf1HEXMCTugAbSl//Bf6vaxWWrJZqA
t/7zoGn6qQowbXAg/CW5SBKguzv9GyjrRkwNuhL328Pwrb6CZ8l5Lx05T5YNeBzwnWiLXuNMDTjz
4vv0nHycEPooZ1LtIYI9ZiX/cjH81TweF/N++MAb+7uJQX1tHDOApKQnLS6gR6u+hbfXe9+LYOFP
0M/MeNkFOLb8S0VT6RUGd2xq/KfxwQ6h9IVECZoiXDg/maIsp+6e9RDOlbjWH7cNk8audhZqrrM6
mD2FvRdsYekkOrKvFurLfFGTK8Ikbn1//RYPSlgnoryO1TkfIXqFtvWNy9BwCBsGnqTwkPL2KI5N
yiejCKq/kjTg7HnDlY66kq059yvS0cmk4swKUVX1+hIJy01X3b/WJzRSgGmpFoumDKe5o/tDZCs6
xnc1IMJfgakYvYNJ+HuQn6BaLsFx9O+U6UV7JdGpVpBGWDntk5ibACgQUczSh0FzptGotjqtIjQJ
zZ4jH4uuZmDMYp4Bp+lZQWSYtmcMhW//KHb9cYGMJZexggJn9cyBKZa/Ri2MmhfnZngrl14P5hdA
j2V0f3SnCvXvVLg/RQClMZDXPUSS6ff+dH4SCz3htZupvMYkHjyvtOLe2RpPPJ7eqxj492y3ACVd
nlsPHLaF22W6b6exqwnXo19ljzz2ZNdjtm2J38+7KvkaAs6qU9QuP5Zi1XP8aE36zEL4aCTPGD5e
J2oSS5VXKj9BZ6JJbar0N8o3FiyvpITnct+h1/D2knSyTfP8nvcfBl0kiPUBUTwa3WK3fYHzd0eS
+2es5UgQQRXneSIGVPIbK0huEFCJkkCpZALfEQTaEG22ztQ2fgT3TAMcOQJspOpo0prEvI5+UgEC
evq8esHx/Z0xhCSPJea1IZ/JYBf/hQ/za+6dWFEtQgPFMs+pcdtEZ/74/or2GzjrRQbLYxRiFL37
1nPeAjCXz83nOZaOpnP9NQZNhXTAm7WsWIrEiu+gX0MnPQ1/49MzCaQ3RhG/rWyh/JMrqsAso1Ry
H33NxADGYYaXi3yMbgGAtyuiOS4eDm42U3cWfkRmt2AW1RcJ41yjs2FdpviGwdhZTYEafc4+YSII
klMOPBkl10J8mjhL5ffpd/62iBFE7xdrAF73CBCCuUmK3RTXpmLqDP5R/uxr+OqvWGQZbiJV0cqe
ejD2TBTD/jbyIaUhDVH8J4WVAby6ZCTO3n+XoY1AO7riNXa5hDePLoWumz7tZQ34nhnB6OScDp66
N0nLeuvR2KXk3deRFdFiZ5vTSbgvwY0wlJJ/xPZ3syJki2ScMTJWNgJFacJC4dcJuU6FB8Vo690I
+d+KHsuTJFHWDoznh9+HErPuqZXtQMQ1UezPrD+9sDcXFaOiUBAtETj1q9K/wUZ/5GPn0cR4oUE1
e1CitnQOsY+6hFsis0WCW2Ytqk3Y6mUz7p9ZP7inyqrNptn46O69pk8+DRiYtSj9MndugCazKP5h
HaeMkntvJ2q/u5UfSJnTOroHifzkaHQdKVtzdk7LorCtjsyqHLqOrFnfUDY9STt6pnZbJFrFey+a
VgBzY3bH2QxnaPqRnTPziJew4TQJqtdYd5UTsQEBB7z/qi1ZuqIcRVb8CYqZ15g3dUwfGEj6qjA4
Ct85ipZnWvzBSzQuM+5eE413Z7qKOzkXMD7fqPNvHBD/VjTtLIK+SGyZEXc8qFW6UxoKyRRByRTT
CGJEOYjrKwh2H4wP6TX/6ukxz7r5c+X1cSJvNjgjK3+wr3d9MJd37t5LYuDL+NbVgmBS+P5wkbAw
yDkelEx9z/FEl5ytnNcssPKlYXH3iCvFezL85TXa9tkuJTicE8tdDpKrN3Cl0GRLBd6xRsQkEdJD
uv92gU9MMKZWpstyP+4Pv4YzNOQBb+t2IXatdvSZHWD2tbQpxql8o08j9gd7lH3oTg7wBVS4YTF5
gDD4MAC7OPAkcZaSrZXng+GEiJAJjuzPoNaUCZbPg9lohQxmR0Tk5SjR6snM2LPMExStFWFw/y3i
3c2TmGx1CX5p2XtVtVubm5iVGEXar8OvaGjtNgznvoifUZFuxS7WTGjt3rKTVaENZ9M4XCNpQCbd
wlcbfhqs2OzwODcp+tOadB3ueredyvx/1H6LbdXcOflJVdgVj5dBTzAwAD0EmzUOwU3pt007i+9q
rL5TpQsweCMXlxve0f0BXl2GSBQAb+q5RVXYmdn5jiUGeDUtQiG8cA8lh6RJtxbK9cGW0pi2161I
a79VZZ81/6diT5seQjyoT/F5Ci8tBptp+zMizL+ebO89v0uDy3wbuHbeudapE41v4MnaPAf7H45I
0NLpbVJEVGJM6bHvijmIt9g+7aoXo9W69jFiN7vjrk0hggPg9XDcEHxaAwTKFq5gCjuAwjyKaIaO
vwAG684zY4jh2dDQOLMltJHF0cloGtTGTVoV9/6wFoVKayc6b9iS21ldCAJsvuhw/X9nI/wH47/g
4gRq0JgREYw7TyHVWUOXSo/b4wrsxypKY18li2ldBnBRDQIBIIvlsem3X/cCjHPo7rudM3sqQBz0
fAjgP2H5baW3O1mXDMhr/T4ambrjchzWiBcxtFCopz0tupzExDH4kkjU4P16jP8r28AoBATETKCy
w9sA8+zANEsbSR2HCKIwhSrAmfUU0JiChg3yVUWRldnlIU+lsqXvVG/kJ+nmN7l/eJJxSvyyF7Ov
xcfxJSSvJuVg9LroBE9mJisgTY9qHd63ULP4h35z5StychBZKdfXXx4h2QF9MXe1/Oi7BfBPaNnE
PJmQHjE8lT4qcGBZa/49icUdISoYLI4+Qmy36H2YyRZca51YEDrz7bmS0fgqYjZnS6Kl+ON/cVHU
RaucaVSUg3UCEJbAXErzAxRen4/0mffCxaECMAX4tLp63xp/QThlJl8OCkhPnI9c5w/9b0sTiHrE
JAOJ+MpXuB4ZRcpK4bl4K9lcDEZUkzoU9sSAWQmhfXu0KAlbw95iQgWd6Wv57KUICcuUNRTwnDyW
LnU0/NORr6rzULDfXnakjN+La8p9VJUScaUtj3WJEUUiwl1qXZEk+J/aowaZ5miULTVZ6WZjqIoH
a+FWblDqsHfznTC7HuncsuZ/9UVG8kqdUzGTyLi8gDe8SbhdSNX0HDYNfcsbOq9G/lawjT0g5Xfh
uSIn+M7DAjSRc6j78VrW/T15roSFHm7U0wRaRtEmNC9tSzlNxIqw2MEwxOLT9pL5IyHvPDuHFpV6
Z5CNy2ZUBMF5YYdVWMN3Qp1Br82dl1hLPckXKqAFPKEnlOXR7BgfjuXSEdZJ10IX+mtGg1edhBvQ
h3HZlMAcRbZLQzDFMVTmqFXJkrv7XI3/eVZyoVMEOf4Qq5svfYhZ+21PJdAvnQkEme2THcAdBrCL
yTZdnGmnI7lz+sWe0VGNtctCTFZgM4dBMrCoFZDzR8iptX0KZAY+nJ70+wilxI7LsX6yP2R26+OG
HR52jOFw+dlNx9KHI9jRDG3quHMrIdm4UQqVtiINKV2Fa3WC92a5y4m87nE+iC+2bc8tZBpLd9d1
veoQFUXMCSma4s+zQLk/FpFEWDliYYvBVJH+Oa+C8QbDRvGaQ4nXwXR11s42bG+3VvfWeTAFr/cZ
ZmAVLBIdez45nDW/DE6LeFtNbFrwP1cAhKr6lKylCtkdu6ND/YjOcIFGAp8Ke3a2o0s2rPq4Julr
3hVXPttB6ktMSdhDIJSGeI1cLU1dWBmDxrlmbIma1s0IkrSnvk43L8ONyxfz6EvRIaw5bHK5n2jK
TNOQVi50VUGGx1uMSSHmE1R1Y7ZTbkvaWCrC2rnmTnbcbWjiexvBPhwDDwLYDH2SWLDWVO+u0ltQ
wlRfhZUxGpmRQkgMaol2PieUXPqEXbuWU2ZsTeQUNaqD8NpxrCR5vv99xwgtc/cOIOY+IoNycHNJ
vu4UMaxTIqWYDPGd4hL7a41O3iBbUiGhr7TqkdiYEUjloXojMm+IxLu1EXZItWLSNgQjMC2xzXUd
1oA4U8DqNnD2TjuuVBCTwg9lbKxuVWS/Um+dZ9eE3GAFDjOI0QWOCS06x24CAifhkAv6RnZ6/ZZJ
JWz5HNBXQTg5KZsZObdUMipsUfNCZpztZQ8UrxcPAnNHiJ/dnaCRfTyJ7osqEnyQ7Cr44sVWG9YA
Rip3e0/sAY+97lxPzmqrNLWWTzkTft0r53JpLX1Bj0k2iBWvyxSN1Pk/bJfIuANsIwBnBaP2ihkJ
KzFT3x98nYEnEdKma0RVzRcnf+bQ22L1l8hlTmgAI9lioYUk5Ktpj2QZ6qw6qAallYidNaB9Ho7R
aH948+9WjK5B4LHVl5uatB7qdGDWtJjhGjLUJW6WwDdVwj4PiNFey1LIpeFwE4h94UiuVl0uvTZ3
/Vx0UKbIG1H/DzuD2UryRBh368amXxB55JQii4V3L1sPaYCxqt29X6/S2LUskAOgXYJ2x8+DGNg3
KPJlfcxRQQcSTxbJWpksK6K2eUhP8hXWfjY2jr0Eel0D/h8fdJ81wYnkuNHdLClLWoyS4+BToizU
pDGeStFsozW805Ny6hRuDKw/w6GsUoj/foCqZSOfjuZPzIZsHeqV2b7OFrAgqqbD7dgKZyJIScHF
vU6JZmzskKroy/XqgAObsjMpb1/wO55K6chrrTo8ijMLs3CjYvFpZsAibHFU89Y22Y6r0E39FmH4
yOh7fnOLQsniUd7wV8CBSB1TYnHEqinNw2U1P0dzWM5wzVZYitGAmv9LybfGhbUeZ2W/BPjxTrTZ
eZB324AQAPfdN2+NsmLGRMlK8oovaEC04AW15j2kMW2arFEvHTxVjruvhwXJCrCuC1PsVv2/ceh+
fuybjplm9AjVmozS1JHiCj5lqHHx4WhmSFv/xoVZr2fP+LSLetTJ4tyfh1y6NMywDCOtOh4ejLjJ
b6eQs3pmgGgqL6HBJWIvAx9acbmizcP3Oz1dWznOJlE7Ms79Q42lgHKZPl/o+1g2OHQlWjHq7VDh
BXLgqYjdFDqKwFe/PCuDj571X2HJAV7aLTwm48GOvEJ2cs1O9R31aH5hytFwOD2n6YcaHOhADYxK
pqkutUnORfaA0zxI8Qrx+7rzBDHqXO7oSxFHpCkDAKnPT6PSF5rJ2p5cB8mm/f970f3xM0p8uPwH
8yUBCVLPJ73fDZlV5ijW2bti68ZOal8uAoRmVZ5q0l8cBsfuWvA+T74TEG/7bATJKKU0uAEeYCUw
sZc5Pcy9CogZw81wEiFm5G+Km1E3d1E5wmJ9d6SvRY8vyH9loF7hGLtyH2OUoNsPMGWUc5Rt/2RZ
3uHx1jTePsRTx6dntv6MOMiHSsn+px9xdlDN5k0afUxcYkMtBG6ZrPNiIMLcqxuj2ZEsvtqyxr8i
VjHjSoCEwh53hxJpwf+IDwmpww1ixCvyofD7FDBylUEyPciVUI5oYDiG89v4ggx6MAzEx/LrL27x
uVK7qS76zFJ9oHE8mflxhP/Ag+IalYGhfs/Vrk795tUkA7792UY/m2P5SQsayYSTnHTg2ETHJvaC
L/dN/I//DolxAdMF2v+/edB5RgZAIzY8KOC7dhOEVa1T5U4L28JSnn50hZNSotTpmta7wlPgPqaH
GIL2/ck1Lh4tNl/vTFlijVEGia7l+SHfm1DdtM2pOT5e05j/kr1NpGdZxlYI+qqoQLGB+5kjT+m+
BgmLFT1dKaz9rTMa0IA5HMQaIjjaxSpOLFX6vUzPi++r+tabD1TuAKY5gbTIXxGIVGrHKKlhk38a
Go0TCDRMygKFk5sD3vNusTNnkwTkP46focfiZEmMNUooAwJZOaf2B2CKTdDdlaEkK4FJ1H+oGjlD
e7teHWV/n/Ahq8SzQGgJQoWQtx3u7KM7fLUWduqGaa+CAedlDsME0YKJ/tG/d0N/qejvEYA4KzDg
+Vxa0+S/MWubmDZktdOYu8bhYUPwqv6MiR0Qs/pUZUpgPxjetBtdZceSzPjX1pfFRCNgAnu87rL8
rgUM9PVl7igk10gph9YyURA1IvcYoegaYMVWOhYVA0m++GW42ek+his0mS9b2zTMBx3SHYzIQ8DQ
Egpg4QbB4yuBQxcoKZhM/eANGlIQB0GY8qBytGD1TlVrkOMFycx4PdQsdZHxDpsB4BqNZt8iuU26
Mj9+sKxtS/wZ8Ta83Df4/Kc0MIb006jjdy6Ezz4dbl44jQOZ9QnWqgWkc6ISsltDOti16npSAtog
jCgVCmuHQ/lPmENQuE60r4hARt/szHe0+kHdgdnJ5qVN+3XK5e6pMWKJBVyG0y64p0XbKQM4WTZV
8x8GafepPU+zx/x8Uc9EP/Xrqbes6JgALd8xFJC2/j2aJCZd6Iq4f2uwLSYnPIU//NdT3oDVApCK
piQcJqAOmGTC/UQP/zrLnoRu9hVON0DyqeCOveiKnfD3Cfj4I3Nk1rb72wR91dPZn/O0/covo3rF
ggFg9MzNXuxWP28v+dVkFkZWHi2t+xRIEol0PU7OBKksH5PIvuxDu9Im3r6sLAnZag1G/OjHGemh
kTyjFguiOdOl8q9mX27BLgSTMyNPxt84vXZZXcinp7AWdstSRm1cVUfGAtycf0BucHGFlyvpL5u0
b644pH7cX/PDTeaqXqquXw/3uWGDoAomiJ5Omf5ltPJiy4e6OEcEwSidXvGVN17FJ3kHCdSkUcPR
WbA4slXtCbFD9kmXzILNglzjKTPHzlKnbuJJMU5twQOIxkoJCiZi30XZocLz9MGgycK8H20sCunj
dhxTxwt4cVSSetN4W+uHwIXALMCwc10cUh0bPKC6C4PdO1OEWPu0HNN54xSHBNww19yc17z4f8sW
PPsqsXol7Ei2pvJ4yW+Ftw1kMCwYqUM9OHbWa7+FItv0wHbCtaJB4prHX+n13q1zAoC/22tcdZjT
tno+xR+c6Xs/Hnk72rla3e+OVew0vDegxqTJkgvEDalNwZQQNGM0ROI5D1kN8jgo8MddWNX71SmT
Mba5J3NoQSZ8uTgkAmC+PwuTSgdqt781PZxcoPFFx8zLZsA1bmNGbGO6U+/Z2QB1YeOM6SwB7FAR
g0HeY/PJCLnSY9iJ8Jgbu5izrwZJCTyOrEo6elyTEn7/3EZ0MHiF0peCupLHLJImlK3ZO3YTy9f+
UcsyXcBgir0E3AtHpw3+ApTiQ3ZZ7hvmQ+mPTRck1nK+PEreDAEiW/xJhR3k0zkoi16ivrqyXlUI
egQ5KNsABeuzEKgjhHK6z+YnQPwRzgFefVokHzj5RIdnNFPVfe8J6XNnnV1CaNvMWDxrXHGpWPE1
uCQ9JWk2agWleHRCEnAbDCARn5WBTjVBoWa+5/WuhHmE+c+YAhTIaHeAhkYeLdW/HAm+ViRe+K+B
IyPUhpxo0Z8DBPFtBd2NJtzvq8XMoKEoJuGFOlTpd5kw/HFX9bGjHjAaAevETDq2rkL0Rxw1CN7Q
eoGlQt9xB3GAYFi//rXe+/MfFy9HPQshykdQq0eGfm0x0JmyJfrKtxr3/XdMCu+WVQPCXS1jkABr
N6Ss4HHUoQDOTBrwnxfLXzSuBeoyx8cAGLcDBv7rar+ykxHKw85qj0G3c3QkLD7wzN4SLrngCiiv
VbKMRKF9crGUfVPsA8s6DO2w0UNkRdRcjHRTcqv2QqCD6MjW1s2um8/haFp3/Mg+MkaM4A0DcC2T
hsR0nzA6G+RV7C0sAQD/Set3+iN7JMB2CXZenIxK/ce+9HDcjjosVX2/6w/CWZ3uHJ2hAye/NzFm
jCPIPbq7z6I7EjKQ7yBRoOY1dXs3cbW/XD4DujW8FNqj3RKTD07NpoW/x20PxojlsZF4PtS0/mpU
Oy2v5v1T5RDBNUt0NTlJFCJ1++CO48sxKOjQnetAXAURTbTOsVjWbyLzgBBZ3UNXtYUT6TGTQXf9
EgR/ZErg1YhOTjg8RF6FohOuXGVpJVGtTJhZii+FiQxS9DtHAAOqK+GdAsbxjv3YNFe5cF3ITl59
ZO8XXdG16Rexz7LqfVudTRmaKIGcrEf5JAcT9yVM7FnzLYu9SX7PN6mM2S+FGzK6IPqaa6pZIuq5
jsGiuDP0MLZWpx+sjY2AhQeGUtb7MUz2dl+TnSvueaTMFhC/5hrDpQkMluhYhNAhIlN3CfNI5zML
mnC5hlIJa/tdW6DPA8nUXZ4Z0YcMu9Acr84v4srrzDacmpMWkXIaRMZF1aKylARYOIsbdpc4u+FF
VFY65GoyWo8FP8Vx/D/8FSA1gJZtynum7W1q5N90Ysi7gLOBRpZw8M3QaxHcaLoA9Ymt3gufO9dT
00ZZCHp3Je2bD6tH01+ql1duGLzKzy0QQxTA80gExfoCNZSE6JZSbwlcJDUg+gvuseyBopFlt02S
SFdYNdQ/W68GWFbdqoj28BgP6gSYXYwhmzuYKUCWIZQqaXPZjuNQgGLiF/xZxzNPTYBxYlfXIu6d
bZxBOt/fFDDM18YLotzsUnXqStkMGkL9m8Qw0/aniC7E4bOPua+3Lm376B+MYB97e1v6q8QgDRMb
/5tg1AbXjEkUPUcLkMAvH3Daf+Dj/V2xcavdC9L8BRFNUEMa5w2utkwCvMc8LALD38VykR/5x/lS
Hg9uarfC6NZHO8eTwF7tIOVtkiq74+p3Aqh8waPDHa4/QAytGSaNkFAS/rzpDekniciyE3yMyIw4
1uTePkYbvyODPs8YMuDpblGuwNg/I1WK/vGvs+RhlMA7tzzCUFsl6LlX9v0zM2HmSmE1j7m8QSfh
gA39Z8R5acXR8RGCaJD4UoXYHd+D9tWpMDFdu20Jv2ki1h+GtMYQamGLGGBt5aKg659BcCDnDJtj
R05B6lXywijrmm8n55JIQBjFbpcHizx6nIRh+ZdiO2atDDSXMtZNRPNS1GIzzgnXBxGX0JFQuLdm
uXc8llRINsNNsKtEl7meFNGPXAb6cQOEP//fB+iUSmdQ0VmVCfPPz46X+B6cZX1dCG80OyCO8Ien
ScuuIgJvJyBKX3eXEc1tnyRpNUxcrLYU9FKluvGPDvwPp+Gg/1mNTy9btVaIvdHHJjwkm3WMUb1s
Qu8e2LkO1dzRB8X4t8ohZ9thD6nNmfMC8wLn2/CfjzU/ExUbZeXJM29tOI+uXXBPhWjmZJ3lZ7lM
i6Y4y8K5AXvpOaoMfYq820Rw79MY6IOcCrEDPYpSxX/js5YHe3SOCpzRVn1An0GNMStOzcdH9VB3
P8cdFWQVyk7ocrDZ1zarBuKmqdlo3eivGHYsUjIH6Cqixa19U1TpcHZGRmUqu7VIv8xqsOyW2xDL
mgJqKB4s2C3ZlKI5iyzGMrIAmt06wZY+yifHqCosOXAj4MyVT6vJ/wq2iUUO1y4s9w2hv73qMYYx
j/X29i2rkYH5Q79Geu6g0LF2sqs0JKdOogKa0/G6YiaaoNSTe7TFUdrW4aLzD13nqWQFWTWqwFat
IEQrP5obkfumBQJG4P4/P+EL7AYH4rvm01yjgV38Y9FkFsWSumR+SuUrtWli9L6ifzPLgKBiRWOi
9JmbdRotTF4zUOp+j1Hr1G6E+WQq2CwUUphmCMJoWTcjq+TFYNJvX8bkcjtjXVRJtQMfrvKz+2dI
KZ/6dkRxQRLqJWv9vfDR2OYVgM7qYGxohKMzGJRLNsvQoOVyoL/7OZgXOI+REYcYmpquB58iEN/V
OtodRpQv3ZeK5mQcYLhNei7O8SORtelAUM6WWRX7bz5WPwetTHV4hwCXiX451Lpv/RS87JRGpZLd
oR4e3XYIFnwemL/SDMjZKpASxVdutxhY/n3s+WbrhM5Z/i5VX9hpXtb0l2RF0MOiUaDDCiTz40A8
uzKgIWok3iB8n7nUjPTxramwh/wnbEg9nriLqCYPc6yi+8/UiOYjgYeRmAYCIKdXRAUDLYJxGIe+
qILNVdsnH3qU9MpZKlRmfugSMS4Tnbm77bGdZyJhj3rhaCGBjpiJ5RwbAFvAbT74rurl5TOgFxeu
DeiTznqeMS0gA/UzwOanUR/hPsWvU26MrmwZlTrmtE0TqYRZUbngAEfKnuOeQOGbRmeQK1vH5W1m
H+tFR+bahmVUXHly3KE/deJcjJ/flIaCzduCRkWCFBnc+NQuB6vh/Q56Yz+gUoqQLybjc5wn8FHt
iD7CQtVQlY14NWpU24/l2AzAEf47WLlZOlLXikH8vQchqRZmMpYic5BP1xqPVnga+fU8IczRIFH1
a9g3hNIVuXSrySbw1VYY3PmbH8D2lPTolLfsSikErCHW4ast9+dL6p4xFEbMc71jzN8Y74FVzmTS
IbH0Y2h8SQNFLcDEoHEom8dxeKmI3sB7Rv/881z7IrUY0VyAxwjUpTzdGj+2TwW7LxHc1A6CSXeJ
XFm8uxKB+vRH+jifkhvoyuef7glls/5E1cdDfIhDouNXVXYzeAL3JFlRg27YWiC+yNt19JwPOFTt
302PlSCPAtOx3nwPiNeWdfJyBPbSxRxrairV4j0m+Q9pCtAMRhJreHqn54TD8lFzAoUX+tCv0dd7
C1k3AON2mMsr2u6OTJB1hfQuPuD2l2wT1V5U5A8W1CXBWuV7eSIe72FdzJ1zN/qkrrGRNLSMx8UY
wAqDBtmP2NM4xQaUNZc8yUDlWueQfa59ma4gpVJAlk1MWcdwftnkjH2wxs9FpqX8owz39pSgB0s+
JxGTBltfYz6oosfjGQ9g47zfflhbYw4WRX0g+I5GL9SLxqJNkN1wtQjPlv4IxACozojC6DcGrs02
xMUsBxTDhq8MdApnnCfjXp9YSw1KsZWnpsPreXC54B2/V6NPbUkuv5ha1KaK7MLb8yD6zDe6FRIY
HYNj0Y23gNg+siJGW5S/dSM/qTtyVzEpFJt/yiCF3yFuQwzzT2u4NovyDgK6kg+0X5Tx0dxd9Kkm
8oPEHAY17RdVzSNM3hBInMjfSSFsh+J/sL3Sjhkyz/EI8p2V37wJMJT3TPHLhvxt0MaK8I8L6vMm
a+qZEQOA3vTClSrH+NQ+sYhGHg3uC/0Jh7rr1a7WbPaAN2Ccz6krPIIAg32ipyt4FckdM/LVDFb/
fiZnv8hNwLO8i6AXO+Puns5Tc+KXH1fWi1os/JzN+PqWOdPRd6gyNsvDgDNratUf3Z7J3dhD9PYI
D26OEFkCMKgtYLx8SOMpBldmR9yJHUZzLDhzjfRUzRF/nMe+t2X6nNKrnrMZ1G/ySCNBES4Iibz9
osncnbqk7kKco9vphz36Lksxo/VXrqQ1me2KgODN0g5AzNhGBujSfGzsiWdFReqtdRfM9dozU40F
XCnYccpnOKL12J49pIbThd53HQKHNbLdTk5/Jws3agHPfWSvHN4yGg+84Oyu6SfTE1pcztkiFjhR
Fhz6ehljl3liUvNPwHNHa3X0/84jMQQAOSaUfPZuF2JdMXBDFzSYSh2MUAzbnfs6wuCetlgpmLGg
LFIZblosBBR+phL96dNQo9uAy2oQnu8aXj33KPhXUzPQg/AFUMAb0CeMcnUkZvvegDjV2lxm+eML
A2gPPFkL+gh6dfU+WdV+B+1RqgvnjaSD2bkpi8wEkTWKV54hd8MsaHYSw6KDpMieYBOV0mWy31We
dynabP13mHm8eWZeliRluVQItTMxT/SQaJu8lAiwdPis4dO+aDW6ddoRyoII91JZhqYM9RDfuFxA
C1nSDQt/rdyrBs1iQitb6WSsbU/MQmW9flv8SOcQfv/7b/wwHLCwLBMsXSRRf6FAIDU8oM5d/UnJ
pVSttxms4t2QcmU6/MjiLcVBoRPQVrujaB8DXG38611S+Y9AlgB/4U0Th4TBpvdXG8POE5+oz9M7
WTRLDQxcfsUZrZuq7XiZJAr/zeJrY80zY6sXtq22QI32WWloHVkMGC3ohqMXnL74hOy4LwmmShMK
GiG5fjgW90oDv94o6RoLbfhZ75eOvLduOvjGrQnZsBUErPUJRhrQYTkSxXnr6g/mv3yXD07h8wRM
XE3qB3123WzHPNr/wWZUjRMM/7Q3kt3SU0qdW1CQ+N+0aGeaDwyhY0Px9i9FyG8psI4fIPqyEbm2
M2vQ2cHPkLKH232icnnaF/Ild67PyMcu2fa9rt0Olh+zEclWGmfrs/t70gSDTa9g6mN1Olv8Pmw1
sRwO4pezHrphZaWMlQjpvNXYF9ckCdDLR8/BvBxCpnRH21jusd2Ke9q6928ZykwDUgQEBSL6VRDj
warggyxUD1a9iJQFzRSHfAQ537fFquZ7+vMOFW00rhy05SmJLUWXqyrtxX5uCod//vIhs41blfCY
mCA1SxSNxbq6DyxC7no7G9JowgBblWZJKRRCiz5fg4xyqiUHfURtvIp8OZsEO9GBxXBgw619I10f
or4Amu8XYdoXGDssGbx/+7w+1pMUjqnORiV+0Z8qC2fLf5Q7FBxyW0axMYJIFp7aZzm64sgmGhwv
I8FIRBk8E1Si53BU8H9PY1qgtEX21YSg5SWSgHYAqm4vMWGTEQBke/B5npHQw569PQK5rQd8iDnk
2NkXh+ZkP1u9LP5uM9C92JVvEFknZxsDNBEF85rkctVf36hVF9Ejkz2i9obllMSwL+o1jgVsnR46
pOkSof4yv0OIO4Xb0zLVhmP8vCEZvaLMw/mm4JqXcsaXZeeSpmKhPl0OCv0l8OwR/RJ1QkSxliu4
4NAUmpUE0gDfZD+QqpiG7JTqpXhaZ6p9YA42/RrvMOwhyNFhMQiA6vn2qcg+Stk1oTeWV8RB3U7u
b68WYJWWwKWUz4eHd3XzFvfItog39VQ/LtdsMovsWii6PfP2tGdPt6kn1VL6N5Czb1PUbGdmGUY1
bMnEQSPuTNmC7I2RMJ7sVU6+2yXm2EKzXWAkwhkmrWUy9EWnU9HUjePkXiEimM77JqWPwvZIcpJU
Fv1f2fdKlK3ynwzJCETVeA8yZY1t5rCmYQNg7f5jahdrcl4RvvUZjkV+3lg5g0RRSIkDhV1UdLi/
uitBVDn9hbX78EVf0YNopUB20IisPYFA+55aqKVNA9aO28d80+pT8qjp15lbBCYXwGvJvSD896v4
QSLzU6td+VOE1lh2cxpfl+heOZmoKaIL1opj48TTrAgmVygOxbgDYeeI2wq4m5fc793lcR+OUqfT
rv0EU8MehQuSFfS0xnfJFDGJbu7OGlHhqPTuos8Px/p/jNL/4e+l1hTGabEevcu76MBHcXPPzRXV
Kbc0qh64A98AzWNipTTDsirtRz0vjqTofuYy0D5I5nsHhgkb4nZnym32uxveqiSXxTxd0DmDSTsI
hlfDxCQ9yRcEnFMfv/TwBBB/+mpGNdkG606GfbhimxkaJMIDLwZPPaRLIQPKO45eLBSM/C37pane
r7RxAit+iamUBbsdGbSP2MU+V3KhpRl1b0kW1KlAOTkTGDYysDVnDmjUqcxjPfelbL+W4KN33q6+
ykQlrL2tM5mJMNIgLiMcCoEQ9hX0WOt1DWBaOzKAANAEedEfqJJw5WVmwOqHtUXuNs0tA+SekpIQ
BYm8nAOZNCiC6g1ERJMkUuv2hm9s7BlFKPJ8a36BxdVqKY6gXj+Opd712TCjeexjzBe1Unn+tYJk
S4KLLT61yFNOQmeaC50rf+NAoUQcwT2oeob2iRIAt/4DRc3bO+sfZ/FJdZiCpSUTdBinFURwQ2tv
OoP3Ed1jJxADO4SeV0ir4HK4N2tqdNZR6vsBaynfDqq/km0YieDIxftuOMRta42YI9i/TSP+hndL
SB/46CAO5A6XKJpCqNVwGoId97oH1jrlR+Mi4FTxMov5Scet+0MsqW3ADwVuU/gka0ykhB0DK8yn
pqgnHjrjmLXHl0KWoG66KP7ElmSNQFw/NSdntULdQoXCvQmfeNztCryKAYDcazpQ3WKRUfNiT3In
XxY0vtl0ueq6KVrB4rfI1w1gKyX02Wzi8OR/VBNPt6/Xoa1r7OpNeyrcWXPT8iClmAqt+wCOjwfu
qfBPXh6wC88nS5NSLbAwNQ+tyYT6QUCXQEwPTxc6ocmo2rY3DVrF/y8Mho7WE0Pfbpplud1vgTeL
FgLQhAoC0dyjlGJs2nE31GKPcYP9754mt2zka/wy+ahoGlV5ZcpNkYICMFBjd2dXNiFsL5HyOf16
12u6c/RaHCyHDiW96qNqbUqdVH7TrX5TitX2dSQjD0s7wVu1XtlrFEU+ya230JPkJQwPSgGFpEvm
GcoLTyDSfyPy7ElquMr0/y2f5Nl1jxvnd1V1pgN75MUoKIihk5YcG3KE//SyBVwlUKHzjoD4BlU9
hqSLRyS7FpqkA4wNZ3axmiHvl8spF31927iLEr/6lA8VNz6T6Q4f/i7gaASAVzNoN+G8C9lnfeo5
IYKZ0mNIaTCNuqqmC4VzPZ+LeQKEc+6bJDytNo9DTu643+tgi/+dRsEtZgT4fmAqEGQ2qTqIXFep
i95E9U4xYKL+xbn1NPpEmWyllpVqZq+yz6zEnYpOeQMAPMNZUf7PPxPl0MAPEJ/T4Elz0/JzOYyi
7x/aG5adlU1kLkfLMAGlaSX7aNs14gnemQWXIMAf2e3dbyrC749kCtl3ofCvukahkQi/r8Ky8lE8
7NbPMwvahzVpxahWKuHwIrAV6fJunH9VMFapHnhdHC1FtlmURQ13tgyNREomHK6YNVzbLxOqlXWO
kxCOkMeF5QQZVcUAcxsPwndbelz3y/4DPfuUUfPPtKe6JnrEz9RQG/Yy1S4I4DBIlM4e89EJ3B2K
r+DciO3YTXm+dWBxUUdVzQzqSED2U6Qj5uI8guHXTjfV5lAdDcMj832QZBoe7ke1xv5oiRK79Dcj
uyCcthtbrRd5UVCwCtDFgfnmeI3OFi+nt33OffcTM7emUG3zzN7WmxpVgCyy0OWjY2wfEh1w4dj8
UiJP8rOfD4bg0sSERUMlmlmX6AhEgPcmkESMCUaMFX+zJrePY2INCzRZ/KhkoPi9Th4f6qp5mGuW
vM4nJKVXQ1ORGwGnOa82tc+Ki+lemZ3L0pgJ5n0MAJ2YNYtG8qb5nqBwkXbxsE/NIvdVQy7/bga+
ug0hsH5/7QCdChX6ro04Usn8Bxf4E6r+mR7rpFCT2XW2wsJipmbCqnkv8WU1lWvMxsAEzSboXWSY
n0iu9huQgN52t46VIvx/puSn+09LGb6MQJhoOSwshwePti0Z2RILRY02oWxOao6bUG7o7gIrl0Kl
Jsdkr3immkk2U3jLfHx7kWqKhDKuJhDXO0OZDZNfHVZMxiO5T8oDarpSeBMHHcRWcR9S0qJekNUe
VI5gsqYQdSOYtVqj43Bd3tguQ1fnIGuq0yVURnat2z5PX/6wkJbPNwH8ySGy4s5zYAdt5WDj8Xyc
UYELJ38XVuwlydl6vJ0ZR7OWSf6Y7Lx3mu6SLvnacJAlE/iCTlCcwwp9P8nI6GqtBOaWccx4Za23
06Ipw7zo64ShxnNkkNfHmgqiKFkDCi/+aCD2zN9FVkzgTxfEUhqARh6bSsKvB9q9d8qNYBdu6ecI
derkuRjyjMlEyUGprhPux2dKWY8xgBLwHN/OBcD12VbTTGn9oP6xGf9qHELb2pB+zsEZJc6cUjrU
ndGHumJ4PdwfPAiXkpCrVInedPis0ZgiO4YrzD0x499kllP9KSvm27a4YmOzD6whLhYC/0oep4/y
rELz8re2QUOm018G34INSurKkp+8gUkG5Zry4hgDvCGuwnyBDEXQhhFIcZK9P4IEyH+a7SDkZxMp
iQSimrZUZkEgBx7LnXvFPCm8lo6FivEzEuzvPop/I4FzpVE6o3IiBkaoIkYw7kOflVDIub7Gpef+
RfCPK7jK8MTsK3Z3d+XXnO8PwTdwfoYNJKrzhTiVmUzUwotDxz2otXyu7mBctcxuKyQ9TTz92NkN
jEV06GGyQmPZugKGvX19Jpwm+mFb6fXg8ObxzVxd9SKedYwEeEQ4jDadktyB7tWWTxT1xB9HBVBs
epQzjgnuz7Rw2YKzEhZrCddCFN9NZgiSecMcyMONgN8BJGp7NdWx0QvsMv43vlCkV7Xfkc9NDaBn
fXASFfRBG3vSvNSftCiNrAl57gP0sx6ps/7y+5C+Vs97gxKAv6J3H4rW9hsS4mXidJ4iqeTfFsQ4
eMaEsafK11eH3SLyQAl6SZxef6afyE+rJCsMcIBsf+RB4IUfhFE86bX+Cbd/m2VYfajgeNmoY/OK
UsKWYLXHW0lYulFyNsQ3C6IFCMYWJXSzzXoVujnqbG5a/3ca9fnQApj9Z0BGL2rJ6iM3JefwhftZ
F70+IxnLTagnPoHilCAscjZ3KeVZAq9+U/msv6B+MGTp0yT4uzmX5ASdDmpFMbC2fkd2J0+txQtP
2gMSu2aeyYZsXVvpqtpYOY8dXx5geeu6wpaZlvRQIjIZQRG5q6nasmr8BrunQxoTDypUE/CUYi0C
suxM/gdD/jSvOEVjvzKpGoUa+wjTrB+lI94rfPhy7km+n2jwvCc7kBcnP8iZqZDaHe4P4eL2s9HU
AmSR653n9kpU+ivWaEBWTEQD4Zp5YrYma8kV7qykQhL2FGWGpODswexrkjoOtalRnJh+449d4bIz
73qGeIFt4H9W8WSfkm+d8XYmdnrhZ6SUhZWTrVzf98kZKLJeejBigrErDbN+BVAeQro7MJfJMiuI
ScIW49+d20CFI47y5iQv+rXPcVxB+kwywhdKtUwd1D1Rkrqr7DI6wABZgQt4iBaI+6KM7pmRWbQc
GuupDCcFgXbji+0szMXFU44gm9aNOQ3TcTPFLe9A5Sm39aiQWLrsfp+jsFVS5ttnAdF52bf6Bcpz
lsk3HvLepfghS2Gh4g0VJugRbNMr3CXw/i5o6ViMGuhO/mU8NflwgaqrLckqNg9t5YKWkaPZhYB2
ACroAoK6d7/lbQWLean2mg8iLnxr1xtV+UflsKqPSEoJ4OogsryXwp3m9s5f+TYyD6dmJUoBONar
1AWdGGI+7dPDXOy2LuLOJc5WWOyUvMSEZsk3PSkJJfpSH9jL23ZMUTr7P6I9DCupWAEqbjDReYXa
Tp37/OjsMSbxa5qVRLqXOmVIiQ8E6Xq/A/QaDzzYaKaxqLHspIFtO+fqZUHsGAsezSbIttNSM09b
JqHTUkGJU5ZDwaZ9sa1iik3s79kRQHpuvxYGhvWmCTpUPu8d1KdRJlLAmvXIFCrmQT/BYvA1O825
gmFasc0TfZcg1TD5hlc6NDjKonC/ji5jn+jPxzexdW2nBG9qkJ7TP5zGFyzFaZc/drsRr16PmQAl
lv3pj5ie4b248w8iXcn0ixTBcL8eew2RSxWh7brHtCEy71tZAjcj/YsT87oPkiazjN1Pu4mRrwl/
+K+oSbSwvwo4SHtRVl/qSloHU211Xy4i6QiM6Ayc0qafVt+owvrVEboGP1bJQzE8whcOv01w+5H+
0Qb5XjSICXq+PJxFuY4mgxew6rMD1RK39HbHbwDvlRC+GTJHrVN/u1NvLRMhVAqG1ftifLrL0xKL
nhK0oH/uxV29MrV0p82mcdwgbfP+eLpcnCqYO1khVbQWVMFVfjIstN/zjNt2igNXLmvdIDD0RUXE
3Dt5aJVrSI3k7UERD60K4QicVItc1WK7xqaGoJTtR+loRb8OXT1cG+eZqXxa3bwUIoYJ2buIC+Ld
j0nW65AzdbES4TeKYE/kuNW6XXOTSLWxa3JgRO4ei3IR0J19xlaPwl9cqyphtA8QDSe0BiolvXqV
oacmUC56GgkyrLn8S/H66qcE5+uK5gnqrc5alQ0unRRQiay1Id1XweonpSe/ikjPx4EBi8m0K1wE
0GmxiozSWgVSbtnpMHubNLNbBzM32noFtLRHXA+xmWCzrjTs3R0OYdqNBSHMulie59ZRoG593qQ4
A2Mcf6ZzywhHBjB0PtCjjDK0JREnlxq8U2el7yJ/dNCFLqbXGDfiRncgvigbsysJO90ROJ7XO9X8
aAM8xmtSiVWAogzzPW197Yi3kzBSTw9gxvup9SyOlNL73+lXQYvMLwNXWoUYy9OXeKL/o0JWaiPU
FhaLcfPcT2Ifb7LT669v4wfw6gLjqsg5aZFgTgNc+SIhZTbVVNowaPh97fe2O0p6jl2OkvEY2IRk
7a4UScaYRrmOFFXrsH3D+cJjMGShRJEaKYOpwbf/M22XaCeVq5Oo6/i26Jv47ohOxDYV4yzYe8br
TlV0aVk0xtYiEQEiYvpZ7fSSTaBTkHAQjQaD5PnLUNEJZ4PA6pXg4+hjwz4y6ltLj2hTqcpMpcm1
JlXbJKKSuYGY8mD+dhT+o5Oeo7Lsm+uoavG8zK8OMj7Co6YKACg4Tu746FrjHH8Aw6e3lExy7bNg
N7xO8/RsU5lWhQK5AWt7h3YjVOjIjtTJ5vSBpYWAyp4SZl0eL4i6aEzLYdxtkBBA1YWz51oCWgF+
9jvUzEJmxfCZH5n2njzTgedJctU7HUfbclVmhKDhTgIAY3owVQpImjHwsmv8I8LCYEIkEj4cImYi
ouFtryP/eu2jai+G+8aaY8uLRhfScAVSEnxM6LEJQ0PTN24rjfQWCm3nWlbjGMthqzFZ2C7ytDfQ
XYc+0drRvesAKM9G44erxbYcxNe53iLEYO0cl0r8dO6LO5uFMyzbILS2xWsyJ5tn0UEtlu4OVvoR
4OOLUdvjeWWKFFFLH2irQMmknQHOASEqPaSZa1+yBbPbL7kOhuTVj0tNwOBNs8iAzH+qlq0FWRuI
vNfj4IJzSg9Jri0E6BpxFUhdo90K0VOujbyvaaw338+HgTREPLl8Udx8b38e4utd+dlHobvBMzee
UIQJsth+dOhD+c2nR9IkCiQ84VLMajiPxi6Gk1fFpP17Vhhq2Oe15kyRQiHoIQI1afT97RYMMWiV
5ZGPVbubQussNHfdUklQy492q0qnAG65wlgugFy6iG2VAFskHzlQ4fgmb61Ywr3aZqp1tki5YdOb
D1wRNYCkltanYZjaEKYx1aVFDm0PUtEroM1c9e+hLT1cHDQex9R1UUzAT0PTGZAuIULPOfO5CZp8
vm9MyKz2RbUyMZaFvxeI8/Ir7wEspUuPWhvbxvPaP0SzmUeGkcevsyAf0M2lVgWkcURyJ3cUkQ/A
tRZOvQqJl6uCfLVshUiIvWYx76vpjZRWxGtQIRkOcPBQ4I0TUkILhyMAuBAQJoDEXrORPv36Pyb0
/qe2u4vtwBscGTkMBujZcO/EtMyKLK52b6dRgdZVXgQ2eE/a0MkS5/wrohqTjDtKhb7/mWYwvXCy
1dBo3k1LJZG+rdgMERQIUCdBqIpA5iigOYo8wz6cP6vr6or8T3oSdYT3G9II03GaHA+fPflBzNgW
NEv8DDUoOQ83Chl3j7HRSRVg8bVEWkqRiDCUgGW4hyGIBqRe/cZT1plUP09bwDSNaYP8FyPT+7Q1
dfUktauJ0kexyWy0A6fM86C+cFdOk+rzwy3lpdoASUruBLF2bQk8l4s6MKKnLr7JHmYJbfq+ylsv
9C4j9oYn7DWnIv3QvWXJw+Y+3L72LE3KSlLTFxqTxTCotB7TaLhkPcuLeqv3Zwr8Tq1mSEySCtGu
alfnl9IIsxk1gdUkmdjNtiQ8QyDHP225kHPwiVlimVg6OYhp1GxSBPeiq7GnApdFFQPmcHuAfcvW
1ZWL7GfQAX+MXyMVQnNe2A2agWdVg9mSfIHFfk3+xiZoRifxA+tfeadIXDPD413uZ421VUZZRc77
MPC8XOINmoakna0quJGEaidcTBmWQ0JTlz/9oL6h9yKHSWBPEwdm2BOLEvmbu7uoLoWt6D8Sighg
j1egGZYcSnet+uaAWgc8BNYXj2nljOfk+d9zOHeIMlcQeA4Kqz1mDbGRaVVr2xlZCn2qg5C6jH0B
uSvi92FHeKlEI0qzMvVUFi+uCceAO+TGbqInqfoD0s1a6u6KVcVOQ0BeE9+3TCBPRlNajDKVnSZ0
H7YyPWD8qA8YvjnE3m+/dTpQpnb8WrFcZNVb3ZP0+ztJTFZ41QewK5oglQVv5R6h19vFoAzbTSl6
FgJW7Hwrh4eUyS4UrWolTIxq+CW+lnv8xKRr1VFPjkJdxSwtOfpy3OqRX5eLhOx3JM8qqLd/WrjI
mUCxSIOSQZHJd6wVokPJFCXNHGdQOC/6BVusApNtC2qmDqvDxLT26GX27w0XgVShuWPsuWGDMPkU
3qmSqlpPDjuWcAGRK6yIsksNTEenpF5BMiqWZybv7psyRnyJ+WOqIoMVEKTvwI6M/cWxvDEktnKr
StNlEJgYQAeyFek6IRc4hGioX3ABf8TUTFKMPgGO1Ld8BlR+R3L9fJb4Pd9T86U5bl9IrFB5vEh8
gmBk3jnTWAHZWvDbnque53x1QAPUS5C1r95aG4uJVdIETytK6eh7QjrnG7ZSFxNhVaSMUCqwrRXV
Oy75JBuwCx1II/Ny7KMnF6uW7ZBPENVj9/xBMVCq9oTQupQDILVtY3ca/3LxolRgjIuLhVhHMpML
M5LPgV2vo6CoJ2o4tamHoT/PysPqhyTjwWNKitSr9UZKmSf2iXZFBPfi28DueClWhGQxjck6aqLk
Ex15Ek4e7IqcpTzDuv+WTXhfZTmJOdTaBOXC/P+TOV/lxA+HdvWYBY7MClDar8FXk+IW+1W0vswP
x0iUf8dQwEYG+GMtPinSHKixNwE590aOnKMGbS7H3hcXHiRaIwuHLIdqrzIFDIa0Wb+vtkmunpBV
GUzhnqXUnyhphTXhJgXqSMM4Sq4vUXTGF/t5oueqpPKiH6IfOo0TmaB7D0Vm5ML8ogjbfr33XceS
n5QNReE0Dc8DWdH2vVPUtUhrb29u2sldbWQtMn4Rm28EFLBA0Lw1ykFL1X4tuuTMUj01zEaWGcOi
zWVQQ50GS0MSkrvvVP7DiUjIO7g8Snm3DoOGPAAUL8RR0vVIle73G+O/v74ouuc7uo5hb6nMVKQf
8W0zt2QYKrQR858FIxi2mTjZFmzp9hWZ4TA0XhsSb79so9WiOkM2G1yt5eqe+TIndza0imMFUVag
uyqSeKdXT0vgWjNzw/SZBBqtjrdUg/QoJmR9qEVBrANVtrNCRXQl44DBQ7FbV94Y6YtRK3L3b6vD
YRXfLU00pwxeLwJwNEjmIZJO6lbIX2RajdracxtURKnUIOCj0jxjuMBp7U1tEIAUdcEl61YPJLRZ
t8N+91CT8HMXm0pMW6YCLnXt0/HzHetHhYvU+q6MU8UOgx/ltmEWPm4hVeKNOcxYUEhrhiaZ2JGf
41T7AO8wPd+kqdMhatd8rkAvbVhf3DCO8wPGacF/ttj5bH4j7S8Vkj09WSBNAVszzESxCx0mz/Eh
+ccYZ0sLT1t9lN8kNpshIPppZMToJ79JoCd1EXcAO16XoNUv72jqK/kcsrgCP5UtfPZgwwnx+IfH
Ihux+kso88V9pw0J6QlBqv9fZsI4O4pStYZGPQUi8oP8cjhwK+B0TBqo7BRPkK2svm19sC6mKgI+
//VdrnUT1pUxcmRKT5XrNI429IyjCsSVT32EkaZTeXLXn4VQN76hVuz94P/3nPLBOg8AIc+3HQA4
mdPP3fAOEl8kp00GWT2/kTMGSl3SEDuv/rEmfMTc90ODJSNclngowu3iImo3CAj8jKNvzqVYlTir
/nWAPM3eEV+0uQ7vsGmJqKCe7ZjM+OUearmw50Z51WOjM4R+tEww9ggMl+3ZIovc4Hhb/mYH3Wdl
cG9W/tGzs6YkfuRV4ByfDoCCh1vTmm4gZ+s6JTuutR/PgY9QRCVoV5uWpadz5gLPDLiQ5hYsVTRF
X7+ZurxKmQJs2rViU0c4KnQpTze8uBXIFp/fguSc+Otl3RZ9n0ZURiFEBRoj+eB1CekEqBIjyCvF
yUmms887zo8YeD/mf22Fzq1tOMd8BqYUrkW+z1lKXjKVMSUS5yDfcukxW/gRytmJwaAtvTruSHcv
n1gkSwL7xBfBCCPBpHFbnJrG1fkYdYUX9QKOsFCOIN9d5uyd03cNShus3rkscYHS7RKSLyCinIDR
6vxx6RUQsCnj+85x+nTI1IH82Za/0x73fCj6AA3NXA4POpjiLMbhPIc21EWUXtH1meG8B+lAr5sp
iAUFKkbva4jKwXQ9o3VjPQTJFki1oduMOzgXpA4zaJCZBj67csztB8pjPUYtldS7chWQ3FIRTali
mkFrPg9EfmzzXvcwvSHlLy7IEXRecPjCMj0lyB/yFUdCIV5ttvsInMSie5MhJ/O5rtCpy4KJMLbT
wMIVGr1drk4Z2HkXTK8wxEQ977OPw5OnyuIbZL6uv7pcmZkUEVmNVhPNve+StC/+69Wrx2yKtz5L
LUg1/NM2q8JkkBaOvFMT7mv/pLIhl1F/DaCBcslIUym09DKD2x+hWZfCMvOO5TAWku/Ppf2z8rg/
1QoYzhjbo7XR0DQGgFIdmYAnBuRkJux7naKgi9x/oYW0K97njdDHon5mXOh2fB/WJoTYKQ56xQcD
dWHA9N+x7RA8FjSY+EOUTkL9M/1UrMQZQfohtsdHMdMRRvpVCcmtWZQb4QrsVyQ9JuBgZ6dVT4ey
rLIkw9m6qwLkQuTYERJoE86a0uxOlBU3IRH3z/4Az6mH4GRwKA1vz+H0/Mh11eJGLMMzwwUBaQa8
wAT8Tqwiw12xWZUxYTjBDfpI/3Z8riWvlTM5gUABveOD1yU5fCvMU0sNldtWXdQHpo6k9qgrS+aN
KEYajWBFGzdI9Y5zK5cIdmjz7Z5m3n9E2ksEZuU5GFehlmG8QPeA73kjANSgie6f0NG7KdZbEoeF
aHmiwcWhrEuW3ge23l1V7k1LBG7NbJ3AHR3SLu2BuwLEL8iTmcxC2yUhoxCFoTrj6Xi1O7eVCCK1
GHTIKPHDGtTDhWB7NuJ0psg7LFG/KXsBOS4+yL40a4g4yAroTEVFL2WmNdJTYmBZOdl48idaBK7Q
753nqh6GkWvQryJJkPjUKt4fxACELf4iJ3HyWGFiledxx1ZfjKgXcnOKV+qT1qbjkD+076S907cU
4KwR44TljaogxH/Oc77bti2NA/dYa3SxhU3eBMMGoHndCIqoq0bkvY+9o+r+LpanyDXw4ko4xMDt
D4wxEVJ1p47X2vkHpA0dzfrKUN1SvPEzIy1TGB8xQkdcyhXGiJFdjg5Ve2hEKKJhJoyIeATyRWoF
rs7ynjpg30CATFL7zuX06Rpx9pyAs6BNvHmMv5nZ0PNee8QRndYDIJn9LF7eeFjXGYQGPJzhmL5X
JntpWaGBjywSkZko85EreX0F36Qh78kb04WZUx5AK4wmwEAzZPrJbvj/gWNPRmXiPBE6ewCChPyX
JlkbtBMfXhaWjwfoUBSxMqtYAXc21d9utxdyfN2yT9iDk0cgTpu0mDVEommRzlGRojtMxsbNOloU
L4O7LsfZGlfHxO+6K1e1YdWRZVVjsjM1LikEHKcOOJcBxe6ugRAjEwFd92hTqYu4kLpil1dTezVP
7TCVL2jURqvyHBe62CawR9cVAxooFzeiW+VtqVm3Syo/lTQIwzD61g7PPH0IZHiOHkvmfznH7SPg
K334DFpphnlE9unlRkrLAqdzsHitLg/nFUD5FTucNu39y8113gqpr3t9KPQGG6BeCKOyob9mS9a+
xx4iEGmdnf070z9fkchRX34LL/ir+0vsNBhr2i6gPCrVX88ATXHDIvDssm8Mx0TtKwUAMtumljCz
9YNCKr96c3/L7zax/AwEvJpYdY/MLq799Nc8CldaWn2Cu3bEh9Wxsq/gvutXTDI0bE8WA2oKkh4p
UV+Ef4xQTBpMavrcQIpMldQ5JepJuFlkWhdPmGGhbfCze6809++Eypxrn7lLZLkd1X5wLmTXXxYk
+kyFNTDMpYd3Pqzt25DYz/ETUZbQpJCilvZvz/nCnjiVluz29k/nm6CMDZL/hnIBJDCxN1zThk+t
U865ud9YXMw6gsaJzr4I1M5CheiRcvSMosR1PPeoFZIhK/R2KmK3iGc32sawY5k1EqonmodPKKkO
g+GOae9vpzbtpVzevjDXXUp4cCiJTcbOEfuuASJPWbwK/tSdCtOtrS79yUcP4oX7qqhc6Hg6AO8P
6fI3vKVL8LLWNj4NqdcRUxzdrGiCVFX7xRynR1V4MC1lAPQ4W52QmiPJGploxbapm/Oezfdpo8Yd
VppM8qcgRt5R+cxB83N0BrYDLH97cXgNx7TkgP5zQmBsZZv+On9Px1jODBVYeXmhLJcnhvebqYOA
ri+pp/whMeTTLLIUlIQhZCVlYxhnxeQqL3PFVuBTmDidnctVdhFuVvRnrdGCQZonBe8ttX0Wi8pG
Oo/aIEzhaT2uM36UI87s2WbsNX2ChWIQpN0l5yB2bV9Mj+gkkpO3wrRVjCtOmQemywvuxaGnGx94
ta3mh/qBycjVZXBkQwvtsQxddH4zu87pVVM3SAP9a5FXTZO/Zr7aJrWS1p99CKFYIEJpDFeNMPc+
oKBba1pGw+9jHzUncNt/51Jt6y9NicQhiyq8HVXwNTArmOH/R5N8qX/nTtCW5aHp08P6WBXcn3ll
iLmnH6N0pggQswwGkN7ZuTEqExCGtOpm9Dv5AYjAelomK28mTzfpsTr3GG4MJwX1XGYPzDRDSEiY
TaAtiLFK4zvLhIHz2D1WSruXhamDGhUBMjY9YiyiHJbSF50FT+or4ow4Wg/bCjRASafiVHbk5VRU
+YrlXkvnvp0bRWI1WwAtBFSxCDO5Yw585u1i6HlOwYbq9NT+1lFmV2yW2bdcyDZZ0Jbf3nY3evYA
RcQpyWE0u5el+5WNIYhmd9OBwHyoMnB+of00r4k7F2I9fdCb8Y7SYvCc70mqkW3a/xP9NRt9RKU8
PrgI4RlOBdqmTgCZWxhXtndvStleVzzHp+zLq9VXRCYiTnC04YxrPOsQBFnKYo9gYg32or9+W1Xk
EI9BI/wdYY35ug7PWQW2TBmTPo3xubLXAmOywmfxZiEIrA0u16tWIkb2IhR6PgGEswbriSuzPQSi
Eajkbn7SDxZMWulZwr/Zja4wq7+SDznSqdSzn171d+GtcNOJbBMf9A75qAV3mcEX+LCu+7Q7pzAQ
epHUm/9iRlbyNpDVl3bN/TlMTCV0wLNtGOzdZ5bigAIuLzCWX0tE1XFvJ32bdaX5V6AtosKqgHao
jQX7A1jKF5pgmh7nt8gHDpg7fZXFiDDWVpg26RXO6xg8qrnh6aI6y2AInsUDQVx4b0xM9DBJu1/3
UnbLaHHEc2Be8ygqmH4tcY/u/JOnrzlOZ8D2Goa/DZubrUnkDbhDyFn2bi0dG1WoB2DC63pmIChl
u3DM0Ku6DMbZcpd3/jzQCv5o533AbmxXuHdoqwIC9s0AyhhcPgbMvTcK8P3MDjbfLH1T6qKORBYE
vWh9NI1DLjzdVkgVuXgbag4dTlPEH6cPHCx3sQq+aZUBBkB3u+SsLiRX52Fc5BEzIXv57YFftxr2
VrDHMw3M9cNn+WXHxb3aOxfxBKA4UvelHiNik4Ycdd0abscW8vDe3vyM0NNIAbZM900VEzIyGn2v
+d8G3yAu5hCZM0s5s+72rEEFCc0NouVlgKxfFaJd2gAHDUs7TuPPLi9B41FdhR9a9I0uYJWPUIaO
hbl2NBOqlae4ur5ZaPs7P7hVbjjMDzapcANa3FwSr3v3jwbQD9HjFDaKEBcdzslf9pdeVdi6WBvN
S3GlQH9dietXcnM+QJ/t0QEqK8pGXHvy2ClVIPrv1yVjSUpSkf/duf2H471z57svtYOO8B2c5YH8
Da0ymTesB/nJxsp4hga36yH6E2GcbBwHMEaHW58vjEo1hfkhnoPA3r6VFHBiWERm/yewcN1P+rdU
iMxDiXXdopwURTAiKn9UUjZh8A8Go+8OJHBDTz9yhLZkd6T33O99xibPBEy8Z5LgXiNKssJ+C3Ve
FzV9gN/uD8A5h9LBFeEqzy5OkBqEjOqairFTuvkji2Rm9HODtav0Ltintgo1atnA72kmEPF19fff
IFT7b9CEyrrSyOr2btDGt5Z9hID9YyjojrWVa2TmXVVmZAinZxcTuANaCD2uIQQNYHVYbXO6FndC
CRhqN8WbplRreI5mA5gr5XgTCovqr/lsu77X6lQOH3IoQiR8ZM4BKtUfACCA/LIGbBwa/8WZ9mV8
jkKDj7iB6Kn9cdyDkEj+sypva+IeFOKKXYDMbUm+XdVbK+cUZnxNjSvmRG589Xz2bUEFGnNKkqG2
NinmjhS7EGSnONiOe4aSKbJB25jCBkvnSXpyAuOASaZJImSIBj/wk+4PWQsfdl1e33r7B6MP3sDe
a3SUJdLZBMXKnPOGtT6IZ09q8Xemp/McoKjA5kPVhUBzfh0Li5DnHNi0sPd/isd4q7DUcATowDDK
fGJX2kx14Yom53Y6f11r22XRImOvxPdu1uLCMLoP2kx56MlRZE15X+SeRBtAZoUXBJCQs2PNfISX
zHtm0ccVxovVe03lNKPmnW/chOerwehcLV3UpbcSFXLLfgNPWDzYjOm65+zSwrtVFtKteXwI1tn5
rrfPXo+furUGBgP0OdBPeElsmDgsHF67CeMZ9Mhxu8znKRvcBcKuT1aWFdvsiiSB1j3GPq505Vpu
3DuvhPI+naNssD6FMUzIqd5a/DKLtq7lhwYS8fm+IMRJIq0PwH9oLu3I6tAKzP8gpFLl4FfTVCZN
YtAsie715WJeHA+UWoYNGgUpOtBXR/Y7gjD7hQ8gcB5XRQ8RRl/5VNbki7k3EtdWwFWOprKAujKv
p7LnpIwkFdqG7jFeir1ykEoPTysXPLZO9i4Zvd+vRyXZh4H7h++4jEnEOX0VSq0cdg7LBWhRebfj
Y0gFnyQxu3p3K+bvyTP7YvgxwQrTAGZ93sQ3dyd5QFTn6KPpfYsBGvrxLwQ+W9l+CXC36SaVfsDS
zShlT6+vPPneh+1vhjxUF+FaOWqbn+naEMzAVMKsoPx4a0/krwy5RZZKfhK06+QnxfULd7KtpsBR
XABke1Yjse7zA0SYkUKQEiuXHIEmvGckey9BpDcMf9Z6s1mRhYyjVnRhB/bg8PzyCQKHnOKZvjgC
izXhlO8dGi/SZMGfhrXGQvuFmKNKHZ82TCwbIJsQc19AjCTkXzDogEop7+qLT4qA9QEmbhlRK+U+
52XkSjUtQDaoewkqyY1tCcSFo4m9z8ubX34nsdv2WyadIx2yAOmfFoZV2Bmyy5HwOuZBOK+quYkQ
/AP3JDJ6JaNatiTzmhlbIsUFfL3MkuvBLfUmP0cGjcA41PEB4j6kiC3eNCb82SAT10MkZIQqTcGY
gnQDgv0RCgbf7N1VPZw6YjQUewsv3ThesEn+zbvNibKcCDVtUXmVbVeYxlG+vgwvH1lew/rpTHQw
NxmlRHnWEjk9N+Qo7+VRcXLVhrae7zzMlOFA/p+uT9PAl7xFbj4KCOCMrySVK9zgejILHyB6PVUk
RLY0fkbnLpBsFsbbTkDyKadb1smVpDAuPzCxc3p9b0jOqU0/nO6nJGr8nKpl2rUyQBnfZD644+Uw
b1Iw+zYLxmWcMERxnIrsu9aLRDZnBCNJ58BcaI76GFIp80l2Ny0mIin6nsxbCpSjYbHDvonkFRD+
CtovCzIYQtlqRtKC6qmKkC6YjNj0uANTPukH4HXDUCzfNGASZEuKiUAODKxOLNsgBSKSUM4a6RGj
9EyUakaXVop5cyzXI/ySkEDCZh3rsx/hj7dNjjG2dS0RLMZsIQ8YyLDpA/3y7SLPsOXlJYpc917h
lji8Dzt3lZCPv3sDTAB9M7ii/gGtOgfibPCgl+PyksqItOThh+EazzSpLn22lUpcpEN3p/HsiTP/
XEyDtJo1jCOQE+ORz/HC2gKKuHpiUfU+As2HRvKAejPVVPDm+3ks0ANcW2sEGQRqM2oYknxd9mR/
Yqwqc/YwetgIkxr/7ysF/1GxZuvpDH0S6NOmjcmsuMdjQS50aeTj6nCo8l30mMU1f6AL4+b41Jf2
3ExvAfUFQguzJXbUy0dhQcF05NL8uG1657942QRF4BklaXDwEPpc6O0AgnmzUXvu9eAKRDUK7gbg
eBCl9v7rFYehSi6/hHM4GlSt9xVt1zMyhTibCy4IylsLmdxlcskO75/HodWqGTWqgRkNs6uD8AYf
X9F52YbhkDLqzWxK2FcwZGXuWwWAwOJ9R6PAJ9OmjPSQsrShuH8mrqo1JXMm9JC/MXGGmUkK88rf
nO/OBmec4oxM6WTaBKDEs/DykFUOe4/X3Ledp3CYsSkP7Ya4fLSP+rDl6A/oLoXL3eR3krVRNYF2
Yrj04rzGPVm61L94Y5V1I3KBxXSS+jrbKTONc2CAZyj1eUajnmpKC7nox2LLtieMnzI6UJ9J/ikP
YCNTpV+l8zWVs7Nf+EEtIlLfaVPSDVplyHs0mCnEe3jsRemLyxIPsY9BraPg/MZOF/LozMIO/SiG
mWilbn+Y4QO+zNXwirGpzXs8PRsM95Z+v7s2Wzc0J6Z5ZDefrvKFaZS2JHyqdm4aYCt9bsdSvhBK
J+C32xNueUy0Z8GqFASVXl6Y3y54FtnkHajFbCuZ15zNEoaXCY8LNUR07WzkTipdJLYlzw1uZ/Rf
wjRC83mAUT3RdJGuWZ+LnYnlzVxDCaVhQR/9Nxjr3wJx7gj3ZooypLrI9mexLRUdMVLL4ilSj20/
H3afONReBpqJYkInAQvmjGWPGh8cAe4TS9DILrBeIVdd1pNtrR0LRExjCfxvpbPXHgmEdfZqV77G
ZZhx6TOKGpGHAJt/VWWLu1IXIE/TxM5f/Ah5DOf9YJHEaBZRvSXMvy61VaFegQ4xTZ3xq/ggNgvJ
X8NpOcKWtt1wTRB+UkMsQigbJlRN561PMDAVATIbwkDuYy6IoYMFRp1CQMtTbcq9akkNJQ0Lnp8m
XPEksV2Agj80vl1dxhRrPwHxsHDYd9lV3UJ3kBHzmCfgmO6xAr0yWfWY7A9AQnWBdDQl/NtUCfHm
Rv8901lyovGsbQDFmTPeuBuH4JcbJtScKZV4c85aIqsx5/EsULLqA8rmxd9Cx5jWf4QGjgdMnD0G
G0U4vx/APiEk8UxKBqT2JYbIYATQEeDxH17ShfYd8SjtScXThzdXp3s38srvGw14UAfWIxmmpBfK
eVbQKva+toDRfwgu+WezXwHHAargBw4sl/AkXDayPlUGG7zcpmnGnSRAunUcYfEJgHZatkXXnMOI
CoY3ufZVOjv7KidjBcQz7jjHdl079Utw70Vrqp4UMXY8X5mL8nR9k4aC+wkWCIilkXnJzTxyphLa
Llx5JkNxPD8alTWEDjEMkUwdRdn1UWnWIv0CJb6bEId+ROcvfrbmBsBNpB8otEqBUn0sFvMDGmyG
uhv2Yi9BlND1ShSI0gOAeaWpdq6kc5xorKXgr04zTF3rzFcBtux4CaylCLmtWzjKeueG387JLfuD
jiXH/IOtezwBfCRK+XKvxttOpWDNdKzW0Vntxbh3ilQ57Cy3k0SRTHd+Xx+3L/gHZhWZCONUOmhm
r3QFf+Pf99lyyRFKoEHRbt4Mwj0zffXA2GkCbdYrHKexGhNp61Ww9Gv9te39cSON6Cb9o4RNRdX1
l0zf3iR35TQVa9hhJ6lfFRSjDh03buGbb/0+BXZpnVR2HJRjhfp/Op8URlDDy+IihjPM6cyAgMnz
nIK5cduBcpFDsridpA4g0BHpibA0sX2DiLqQP37gXZ2UIOmL4VapIRsSd+T7NfsJg4MsumjMhl+r
/UbZ2qNXghh9Cfls5OxXP0KhDbqYw8gICl+WYmi4sBxTDaTK2iSGQeNn45w8ukDBqZvDx0WLlrtj
zSb2RCFM5hzsviNi+hOyfGRvJYe0+oNpBI6wMZ1eu3Kwld/F+CDd1060XiBd1fl2ms3uJhJZKsVh
vVDTcYKM8gxv6AhjjQXB8gH0By1USKS6UHgZTiskykOsaFN3feztMn4rxSdZEFDOyDFbazyNBbmN
ARCUEpqJRuF1/pUNRXXCWfTCDYHeFRDlO6pXmc2m2/WnnNIuxn5M2uriZRZulosTIj2+q1NVsJ9z
j5MrdoP0usHm4Zhktoij5FAqdBFJUJuW7FFaMAJU18HDB2djojTLc1umPVWFYNcu466zoSn6qKQ2
7yWoT2eeFxd4pGbXJNcMn0+BLJGeaM8+h1cWgyP7ZqGC0HP8FjAFskprs/G25cG6aRrFqAyiI5Ov
vMGZ9yIH4PA8VO6zKniWcbIxB4Dy3YwdWULozjbEBihhoKa52cmS44FaDc21rOk7tmnK6qks65+x
JtREt2y/7kc9ChNUd8k1JqVJcjGHsMVpzrnYPVB9+azPAPlzqgvPo44LJrrunCaSJMQzTtmYH9Yd
hnUMbsPK94n2fOoAbe+n88xd2IUqStKN3mu53J9r9XwO0XbegcrwH/Po/fba9cDJAhSzchs5fT1X
qApGwz13SD0UdNBw951c+1hwVZvf04I1EttI+truiMm/zZoN828VQA2U8zzzbRNB5LTAmPUBO6Ko
O2FRrZXODySazBUaVDxmqABk3bBQEdipXhGVhLCARHIhKXZ/djn+VYvMviFzquM9HH6bA6/gyTBc
vAHnoaSH+S/dIkHp74Eo83jwVd82KtiAw2ToGc6q2Jm0+VAuDhXNvRbK7JiiFFUW/x/PAtkVZWra
5Y2ipjsVk2YIMvWu6c/atbnp3wBfCcNVByM1ONtxllqKciqjXTN9/Q3dBbi7zldqK1LAot7iWuCd
eUj1Cjfm8aF920Q7+LtpkCkTRRmJBgW8N/6CvW0cHOBeDys5uqYUZwNzk18ccVLbFc+dVRs3JlEM
u5C1N4yHMXBPMha+w101mmtKXqbQ4U3Fae9XpBMnsouEznAetQ1zDRrVGUJhvgJ7apjb81nbJ+M7
+T5va5nXw4yHckcPwuq+o36JbHLPkfGWYx/aMxQ9/f8Q5JMaQbYVqeckpUiwBDJX8IwQrnZO7N2U
OikFuy7oIyT0e+baPbcDyUwkTHybOp7a+rPJcBRZjvsxfzV71YRBo7SC16hWa2PcGIC9Y1+sblYR
JBnw7uVC3u4nRGM6fJH031VfZem0fnXCSRVZGQi7GrMJgX26qf5Ih/wi+3V34Hgarn2OJF60AqMz
gzFLXTf9CuzNgooa5fqZD/Bm++YZhEmxpZ9L8uf5C53OQyW6hgXR4dX+3n3/8PQzfEkC2kMA2jLr
fN8gtdjdCmssRdfTMlVSMiluc7Sf72/pLk5YzYRxNCH65rDescFcWCaNhs2mmGI4LLDdBBbRtdPk
ojONom39rGf0/4LgLG7fnOGcJSNHfFZqwQVoQVbuIVPaw/f2wmN15ck4WwV0iSAcriyBMuxjucMZ
irR+b9WFJvo6cvNQtZK5483cAsZacmH0SNPmDVIFjMa+QEctseoYWQJ0E9KA1VmODvv6u/j6ssHX
FPhDTHAn2gN74QA7Cmv4ChBIh9EO5R8B7Nr9O8173cgYsUB0SoboZI20dr9+hQ8K59aLtRSrkRvl
bTvoAGl8tRmgtf6+wxdlleDrHpkmCxHIZhtYxvYlPOp/WgECIOoP00T9NlzMmf+MuEnpMO+o/wPv
Xl8J2v3bTiK53S0lJqPwCm1PsQ1cR2pVasVmDrAMCAT8d04KSaMQs8JlJGzcqAsnABwST6XmRquy
8gcTupzFzK/TSawMoZ03nQSeko8ijTTgairl7nwtxjylhgzq5t/RgZSfkiPvBPt6hxP3jzcvxZio
Qc6xYnyI0DG+UXW+x/EXOs4JQ6dZPQuJEEuHr5/qsUButaS9JytkPFHUtCKAemigb0Dg/AJsObrs
b1bRhy7RQP2h/SbumhWMwv8gDtkQ9ehIIPH/2PuiS/Cj58K89pNaUXlFs8DsMUJh0bJXkwwcAeDb
yd2P8V82EvIBuRnUH1ViEl9dXmGz5ppkUe/+JoK+u/g4miHSiPr214psRdbmY9ETWDeab+aIhfjw
uoGecniq187eSlrR/8tygMfBD7PxYx+f8uk8sGhmHU4QFLYxHIiyW4LVBImm5JzDOcf6a+Xc4cpY
PGGd7r0q7E7zYH8bU997spULkfhcQ4ejQOzS65XsvmMT5KjHmQ++vJmJIL0tTuwSP5IKx3tLPnFT
mqHkIl3TzEetl+JiLM/0q0gVy2z9ZPtLHtCRZu0cH98UDwb/gICd/qpr4zrTJijs8gm6+yi2nHiw
yNrdGrur2IvemKBc/BaJcw/RbBTIgooTAEtmWkHLUD8SVPdwLl6QVZpLV2AANWwf8z9Mcfzv3Zek
Yo13ZSUjz9C4KUotkT7PCTDuNbFP52w/l75SO3WI5mqKm5VudYeLZ1PliGrOAzgQ5LhI6Sjp4aED
VU3pMXBsi/C/HZ8W2ORAareEFCa1lrTFyVuvYuWwi3fVlLz0TJfcSaP6pVi1uxmj56GLivR8+6oX
qMRk4RDgwPULArkuzG6sPMQw6pzHzEOYOhrlEhERn8BoUpXdMB3EcZlU7cw6TMQXPveZGnaTIatY
AawhFJplotyznqtwleDwanYJ+b69jLtTfWrUQXMuGj4Uct2gmdqRKtmAjbN/FuwB7MzCeukJzh6X
YzAgUxs14b3GlDbDIOgEIyVTev+mhHjbgWl4cmSSFAv53l+KMmKUAG+eumzWzZckTJQnJYyfjrTH
vetfbrDJHjTdp4QlPvEqKueZzL/MNeS1A7Sg26X+ofmBprkpvof1l5DaktHTON7m+KtRKluX1y2U
c8MLSOmp55ynqzPoWfM+1oZgzRrnBX/ifxTPeJ17807JDDOjM4m57zx6UyeJCga/RKFRu/eGuui5
KzyAl72aU9OWwpUvWhhQgCPy72wDGimjD5VXilTOBV3nrXXN6Yp1VfW/skuXdgPqBQytVwnu2nqj
f4w4YT/3SEO+KbkadMxJtrOew4j3QKGnt/DhOOapRyJEoWSCvGzEyuOMj8MknLBFKagKiJ+oAGqY
lViJcOVEpU8zDWArv5hOdElABsQpvkIpNRiKUX9eWMlM47ew5JaXqDVssWnVsO+W4AJDpJ2rMeD7
AVSJvm5h1crczh7WeFhiL8Kqp8pQvV4VPLcQWj3SS35NDbNg5yDOXAUoDQyzg4StkmPfEGu5c6IV
atolXqAZwZ9q1ZPzR/QZLXn4Xfn4o2cBq3u1zCcswdBakq0oo8o+Oy/WFvaWUEtDKKg62ReXsvi1
oDqpcj9QUgMcwMQCYx0DtiP+pTfqsxMbLlGnbiHci71UZ+AVNgxa8iWW7/D3yN1Qql/+wCe6Y94B
O/q4WW0Og12PDMnOt7ykGOtJHXxumD86o0jEZPPjTzxpQ9AmK0nt1RQKOv2j5Sxavb0OaWbCTqMQ
3hUvuOa1sgUDVGlwOb75NSNTHlVLCcUPZRd738/tWU3rj1biHySzXS78xuiPSxRduPbVtbLiLFyc
RN1FEndPAlrKk4gudejpCTH7RNGTCtra0gpaL4a2Y/MHmMcN0aduI8GAdNQ5ubd49BzC3XTc9cXW
bRY7jr0lR3oYZs1QtBoDHLIsbT/odRMNHWZeMFAmzLBiLffT+PMzy7rNkAsGZoVjDJb6beLvYIzO
avgzs8JyLy1TIiV9k3nKqud+30An6rcO+w/aDDXTjX/ebjeyE4DdLHr2uXMbc1mehLCvlu5lCKH9
+80BzcPksAeYVtIYU1w9wcoOZiyzQspXXJTIQ/lw+pCIwk1jUpuNa0W9NyfpiNLlScC3J7igp7r6
8SDeUE16ID7cIKYsiss0g+5IVdsqGyyXGzZDnJNHll9sACq6+Eps/Y2OqUCFmF1SgXIDuxsb+nIP
Drn8qO24YY/sDPd2jv9s2PqR1J5gU2Nu2efCmogeGRohN4M0upoBcXhyAdVD3TvPwtP/uMpbTHix
90vHDqpGU+yQn+un1lzjiFdgZhIRjhZoryc6WtkqXZfhdO+P3TYA0hKUzgffZEApwLqeMnIIDrg7
+bxOTmJT8PQ+yX2a/q2/rS+KrROHYfysstnl5gPgSblzR3/cs2/0UaPM8IdVqejVSWJ2DidoDNS0
sACkLY+HjOWiOimrChAtYqgRFJSzFhzFfuihDKxYbjx8IRhgp7f5ZMSnJAhoqjKSAKdgooVBQlop
RwITJW1vEDLarIaA6lJnX3gtoOzzvv4K6lCVg+0HMpv/vk1uUAI7hELH6odc5y6GwpOMex9ioHRj
Z/e2X9IOdhwTo/kZlKJVllzWV3KC9LnJAy7HQd632gjslPDctU1iaY5DrsCkeMZO15bsEYRsG6cQ
eGRZZid3aOt5b4x2nNX+sOqY09rK+MCb6X9SP0C4PWxCNeqcJ9ppo5fu781qld15JUTwROK9Tmph
kMefoNjc3BdNK1QYEHaY0EMMoB6SPKUi7AmL2G3kk/jtudNl48F4djacQHNwWwH5LfSyt01PV962
oo0OZQW70a/3Ko+pSOPIDhggjik8q+BQORnXgFpMhrnF4Y/nkE3vWpy4CA1TLKbYjOIaoXoSAn7h
Yum3X6HZoo3YrEIvuSpbgjlAcD+gAfnfgwP75KRcsQP6v1Es/lrwyOg396Xlu51+HrQF1Gvb/wlF
sLrTjI1pWdE+Qk6kQGwkNe1FqvczZ0jO3Mmnd2Yf+xSsltMm6RKgpdr79gpsgoKE7qP8M//WtCP+
MUo1QihteWyNLsdp7D8ybPqG3VO1vDKyOqY9pNYW5TWLpl4oG2BL9g3X6fu4V82XKA5qMFNxAhj+
2Efw0TBGV0DDJsGLr16alTptSjTClxX0GNrUfXMhrHcFOOEGCoPG8iXI/E6OLbm4t2tVg88go9/l
raNvcmeikTvdIMOKtRAdaJW3b5x1a4wdGtW8AtlluoHhTEKQWS2lZXtNuEtwd0X/CkPF+Mg0JP4u
OgRKcS4hd145HMkjkqRQZwe4GFwbZZeQ7Bz7Pa5Zlxwr+XB0SdmNja/EoLN4+mYlUfo9yEbdXULk
AGot1zzBCaF99zpW1vfCvoVp7M0u4zZs7PvYwD6oLrRA+zkJ5U2pCT23VuuWmAldllG5gdbU4tTk
vSvQg7dV+r9zrjzqoIHnnpxQDEocyuxfa+muNsw9LcBUpZkshvXOm7H5r2zIikOlg0a6dBsFOvUq
Wy9AOlV2s52xHE2xjkW5Wcwe6FnyBtrIbZrqiZ63lW01L0TwG3hNGa9aaNT/scqJvUvsZOxg0RU/
ZS8p1Ckqn9AK2OSMv13LtRPZ17aNskJFNzpmWTXDjX6Pxb6GWEIYD9ekDB0qVZJtXU8u5TUKWr17
Q+Yfhnt/CQyFAApShPdaf/h4kDeT050lO3dpvgvqqrpJHGbEb3WPI61Kjti/Gx3BEoc8rKofxH6n
6kumGhK3FVLNbwR+5yl5V2TufTtM5zaIDzkmVsndJvFhGTG/ngTZgD7TFZ12oSxe2idVfm7qyDow
EU2OsmSB2t86YBbaLiQ4zg4q3cf+zWGl8YHkRcAs2zDZLAF7Zc+1QUoloGLnL2RpGreR9SDs6Oo1
QG1PV4G/Jj6UsS6Waen3MHQ7YiwXgkWAs3m1eKGRK4rsoQubi71U/gstCHGA8r5IU1nJsFslgfxJ
BgwIxb0Oz8JxKI4FceuT4UN6DyLz//ffVHXa+erRkBP/GjP1aHesm7ozdPVmfb/+zEDMMx/WdF6g
DSwFS+kd4LRFsN5kEBBmKw4iTXh+8Pb+1//NZ9ml83vXC0BlnxVMosOOl2n2tZdenuvd0tq0j2tq
PhxT8g/pvA+kv/rEldFFKv/2YOBB1Cd8W2y5yWq7amDhmz4PpF3VPemQc9vbw9sKCgzSf8kU/Skm
5KFA1SB4qxsf2JqnCK93ABb13KtqyUM0B2H0nbzdH04oPPhjz5d/NoDafQ/HoKXecuCaayUhQfrA
7iJrMTj/l7KmIi/I6Dtmtx1xO27imX3ZpwhlS/wWWA0UKGKDHn1kv3Yp8onPXwa+GVAOdSttoIkt
GlLAuE1M5HRCJDixhrlVKN0YzXGHmxMuKwhlIo3dFu5pskKJjEsVwR9rnQoQhkjSwbqSFb+n0NfM
w6y6RpMuUGMGM1RZwM4g5AoGZD5LWpXZm4OEkX+VAuvatx2ecUgQKgf4fKpuh5fKClAoWOTjzc6W
+9hh004fL8NkHC0pvVTbdgVhtDErRsQLahyva1af0NUyXjLuSdfPrt6c7poUKfKGbBhAgT4o9gpi
xa4UObDytA5n07u6HJX/blnoavAsFSbeAt428TdDQ06w5TuOJNJ6fe3qF26+Mvlck3ploqTAMm12
oPpzyuh5dtFbTCWn+WVaN4P/+fcYQEsxeNPGNl37auOY+0S/dmOR4j2Fuztq4w9L93OALQWLp/NY
JwYue//YdQY1vUfskC//TO+8CBYUsGRS0nAmzggrveh4o6FsH3b9Lc7TC3t5xGr/fsi4qvb8RHs6
9G4rRXovT4pkoi0hB7J0xahcGuUrZnvry+CydoSYwvWlWHQHPqeUA6efRKnPiK5EtsSRsEFR9mOe
ARUAbT2HIebA80cdy1FdHcG0pKs775UBMyXSTTvE5jXx8SrbuSRxCiQScHB9EBzxKXjDltKce41J
A62Lc9ZCrrUFGh8g3F0Cw69qGvAfsbPQwtfZa1B/8dyoiOn8ORbyPKfbFZHQeP61vR09fSEmxSrW
RJje1qMP+hmGY3bwzfCDUGD08UuNN10BLsnqAFde5RwQp3yQJxOZco5Ud3ZhhTSyReW6+bRXmaC4
dADBwI6VTPNo37tM5yJvrL9kS3EG80LMkCMw7hFyDoX5+LjfMAfUX8EtmejbYBH08olJWWQOYun2
Dn0+DpTx2iHGLzZcpQcCjPHc+EP3dfvv4ZG5vrI9m4Iy/0D1mRKvil06GqBAYvdvUEcYTqNIcPRF
l8Z4iqZrRjqbagO1m3tBYOcs/PG3fyCbOxsssFbWdtTQ+ImY7lGP1wxAOlGeTNJt2IJI7PdZ/a1b
/rUVQRM2Sxk4ZrwogiB5Ffsu0D7Wrw8pDKc6ZpzZmxhejsbW9DQIByLZCJbXHU79nWTEvOyTM3cD
C+A6kZsnCezBLlBYzyLRnXAgbZSU4x55+P9P55fccD5WuwU8BDhynO4sPOgzgKQp/U5+E0wnj2hf
ZgHTOZoGSqlmLxENdDv1K6NXW8BQIQQ0zL8yWGjU6LoXkuXdvm6MnYXhrhJGsoc57385zNCN8jgI
X5saTDJ9n5xnMMWH2djxASk4x3hyn/WIhtjBYAS6Vy3GT2wQBZ45JFS7wWLCFTxZBKAhKO0xz35c
Q/8/Gn6IS69vSVwG7fyrVxLPKRjJBQT2RpuPKNcaW3TFzrvGfztwDUEPKB7QjZpkitjJ+qr7lQsx
HY1EBvqZDh7AdyDzdKvw64YsR99KI1pcPUxYzTzUTgOkZWbTFWnMonfGRWYJpa3PxHQsCUIUSAOy
W1ZKQBB96jrr2f811lITEcXQNEv4vZdELOZtN+vZXaA8zHlLghoZxk8j95XUy6TEDiStHS4zaa1d
0ksrJewZV4RZ0xZ/uswR0D/D5SS6XYxDoVDOKKlTLOt70V6vlXIVn2vhdadDdyt+H6Qr+B24HplD
gKkcaqmGjyF7kLSL59VfnoS6LLp3xxuZe7TAMkvCK26YKaQVDevt+cV4hN6Lv9wVtT+2boBl0naH
pGjzqwILLkOorJNs+XPxHr86BHiyhXRfadnAyykfAObhWNzxxmYwavsFN0IlYBq3Hi6oKvGy4OPK
SGImZVMmEcvTblh0YLLWjvHzn65ngV2MFNLPUZrFfjUQRzzdUUiRybfVB7t+O/SQILg3vGDDMQue
5LzQpe4R6fl6Q39qhfBhdfGDdiiFoH8puJimMpYJ/nwetD2eOlaQFCRuDfy34qsvx56ujx92nNtt
GZczuNKJpqgF4QCe7nWUL+buEkCKe1Qbwo1o1UuRc9KmruP/wH6rZblJFAZWW6GBGF9kvnNuVYTq
GN7VXslBp42mB12IMgTe7MPf7xrejs06ppJo4x3RB4SYJ0ZiGu9CnMwc5cBDkAFaQTebSQBJNaxV
pl/A47dDyBV7HSZo8cruNBaO6vDsqYJxzHdGXLNX/zJGRRzNA5L7gIMJG0ZDrpodSd6RZ124ce+j
n6fVfzUs7wCyXBTl6sY+eEd6X1RsR1/o6ICsCZOuChtckwE3FBPZQz4HRKDBk7QcLVQ8TC8lz5Vy
MEfWceF+4OYOjE3QDbaYSpKXlzDgqBt02FSmIQN1QHqx1m4/u0d2Hd2yxIWMGUE4jKYqYagUih3w
pGFxVp1DQ+CvSmuxJIRQTmzDOGkOL2p7bGdzQ6yakAlmzGW48TNnPEe5p1Ifbmk+q+hziDJ5ZX9u
Upg4+d6SWTtgG5rfllnhiqYV5xQWun9ZbzQFcToP6MEsWeNUPSiM5CBd5bpwqzOwxPyF/Bp4QLnK
S70nX8dKzZlNUtnu8qu7Zvgk2wuz0eAWr8+kl5soj8vFLwWrD5Ki4rG/hBP+Zn0QRJxMIjwz6cGV
F14IsvpB2uFKx3jLKGZAE8EoRAYEWO8KVQGs3DG9UHKAlBVs0ekD0LiA3tN7w7GpJhpTwBW5oJ05
hr6GbYrHAL8m9qTt7MwpN20tvPv6ZAAcKFkKq8wESV51KYt+sBTEQxIXEGKFRXLWID4beUb6VWSp
fqBnyzJOSrx3hA/AOgbkDJasS9LxKVyXrsEbeobIJ3jz+JS5JchkkV85NnEYkxoE2TJKCdnHVLql
duWnkCIA1K4l5ezVei/9Nx45d+JyPwXQ55EKQ2Yvf7uNFFawiqNFkWyvNNWcZHsauzMV00/ee5zE
HzIutC2EkW+UAqjSAF8QhPqad8lcmjQsxUd7q+03RYCVKJqgHtZctA1VLNkJvcKAe0ISmzpImAYv
76VWBaNeHegIPf4ep17YFZ1Sp18vVdkmh0ClqSMxnwSF9zyd8co/zmi4d8ns2kXKjTx/jU7FNEss
tbtWTwMSigGl2ZPjkRa9Oo36/Ota39YVoG0r79cix0hpus30ClO5ZNPiZOupWTdz8I9rDEx7jLGv
KeBjT9hY4nv7274A9IVcudGvjfzdt93YH8+rUBwUIPQb7yzpg1xXguiLWZSF3lbzoCmnOaUUno35
O/Z/29cK7zRPQ0oNjxcKFfLBQ7zkegAGEjYp+sM4OMVstBZl090YiTvawG5j8pFgSR+EiO3UjKEi
hw9rZef01YQDRne161CVwL2hXefersKxTWZQit+eK+6YhvRT6WDZtA/M2+MXc+cEkxdSHtInSoKs
dQbm5LtFbTu1SGZyLa7DHgo5LZJwFnMdN0eCWPNVQtx846NdbrmBCn67a0Q8W4tHNg+0cAmGODa0
ZNIAfqftZf3FP1IdP37a0SLYHDqSgldjTRfK9AZJ0gDy8mS2/qm9VgvKcpzsn+SZIF78rzwDC8UB
3y9BsWFmwHlaRZHMqQb0DmXgpLu165wNVQ+VZ1lepNXcl5LiaUHA1PD9LIbvqMEzcxd/sl19IpY6
QnGM1DMdaXj/VbBpJaPK5clGKtaA7g3psO8bvhGXpRZn7x5jDzAlvh8qh9dSXsK7O72XDEMOyI9N
aM6u6hc7UHmnONk0yNk1/GpbUZc/mRu2SDK8WSU8lIY2M+de9OO5PNoXDTgPiTtpvYSp5lw0Y270
sgwV0elT+TWeg1kMzflwxjVYwMZBj+MB5YnRwY8DCwbRq/oDlwUXohLjqa3ktsKRGVAV7gMfudJX
3H/iJwLFBQsc+5AclBQYZigHFM1/Zo4ivu4QUYrF9rFdxdOj24qeVIkgIt8kGaBN3Ub/l/uADQCs
Y6mA7KgLWGB2V6oh8eZVb0t1pLJKhyGKZr5X9G7yglzoRIJh2GyxGadXqNa+vDtwZYv+wQkJnj5E
MKmU4nShnFcnLskQweSBFfMnFVS5GwMpo29Iy4hehNL5Uyrj5Meeuc01fwuOT4TgR9CBYUPgqQ4J
K9D9p09B1vjFjud762AhN4P2MXEuKtki/7Tb1LhNA5P7pWtmHFMX+cLn0g2mp0FwLv1/pOf3w+LX
gk5Ux9eEmQrf+o6er051yslAoV0oSXFt3BvowjCcGWjopFL8tlxpaV98OgxqYNpLpqC2/t7IduNx
NQGAT9XTPSncsVS643sbzu2zYUVGch6Z9yMAsyBCxaOpCiAjV7M8hv5yUJFefGTDLe1JPeYALaAX
330QxT8GjnjO3b4KhE17vKJC2Xy6DdBZ8gx0xIqiE4wTRO7c5RHUREp7+/4Nyb2FKpo1bwv0afTD
wMj/ZWIm05CVOk/Mc2e7/LmLxn2tk5voL0d/O9dwYo82KnjWEo4dlxx2ozfTsCRskr5gsIBPn83E
+s048H3Rrkf+i9PmuQTcO/JcMUGPa5nXvhA5WP59pInq0aM27X9S7GEa2izJ70wwF7165SQbmQKR
RkuiG3NqREZHcZU0OJ+8gH09v6o+4VbJW7AgSMFDOSMHCDpzTny/4th4vYP+/TLpGWJEp5drHT6C
KgQWMLzZjZdFAh5pO6EM/OzFT1ea/iaSlyHM0Nh5qFyqfvNFSooAXtwdAVlzkgMIRgOyFL3ssqzm
D+L0YDYjYfvbK56PptgqliCncR7fcUPrtYLcBPZ09TgCavC96UMbUFur0j0lXGiGCgYDXQbJ6DGN
ZKktAB5HCgCDzSIAsc4xRnCrIMv1QWSQUnG8xlF3KYO52l61ZF+rW2vgRFk+anRqWPnQT7vtqGke
I8pZBuQ/nrwoP81BmCl2pX0fqjeVA79e5Tjsa4YLrCl/ieUDU+UyyURVB0SQ9xO5owS7TxYLLW8c
4NHrhLTAkSuzDzj98V66kQcMmJ/hJ0BirsYBHscsV03OtEnY6kriw3mUi0y5+cjLLFVOvrmQ8a9i
6dykhJn6KmF0Zz5ZLbV2iq8MkS8jfqW+DwwNIvNmvnydoDC3hCKXkM9B8/FJo7AW6OWuzCpc/LWt
njn1oJQusRqj1AqzntXye8p1uJQDgzK8B6+vk+i5k5ucQQ/wAu5uanRBk8pucFdKZaIoGb4HniI9
rkQhkRKBqQtm8PFWo1MA3l3RwhrvkRTzfhxbA/RrtkQYnPI+HFhDIeJENNE7KOBuZoVxz0Sn8SUD
Ns42k6OVItYjpHqnQ7mH2zbpp2AyfNubqfjLONf7L6kTzFzt0/X5G5IYS7Lu0ilNE9CEDbuz73Ql
yH4njZ2UauAvfNbZKPOusnDn3lqWQz69NvoNoo2pL6AO7K2nk6DC+cu/f27N16eyE6zde1AGagGW
rT1EnNg6TR+3fCiXhPyUe3NCPWv/BpuTTlTBYuySEddFZXRN0U58UU4ForCQT5zq823WBRozPr3W
bWcAkOta8ZbJbYK9d2X3oDuBlHV6Ec2ERoXofclbR+OPuvqTOxlejW+/DNQFpuSNGb609xdx4cOc
hF/ScUEwFXHyLA3xZ2yh487mbFv/bojTA0Fucuf4ZR9XvU/ggu12Z/HIEcfcGjHDEjMRQddQg7d0
Zb97VVcA42NmABQIj5mAfU7uNqT835hCd7H/i/LrEhrZVGQNoT4cv2JhnUrDzkk+pci4W3RMXIdM
UdLWS4t14LdVf0pfjtAJzpmQfMFfcb01sIC8yfmHnKRWTO2dnAdi4aT68J5Z2oUW4dW/5rljjG6+
15D6SEYa6VZTo8k46A8fbzMABa+cUekhYAiAOc6sqTHNa5/vrytP/WMiN1pNiZdERlZib4BuGnUX
9lBPsZPGQNYmlNP6lEb62lNs/JoUC5JiNV5+OWEFrWzUGzCnybJAGaTrcdUIkNLNvn7wN6PprwbH
dFfWr/1aMfEtyrG5cSknEvL7bvXn/2k+LvlDkN19nyhXCaiG50TIAW4k0HopNIAx53NLR+/KCQ2E
WRR2AMQQQO5QEi82weDAiDMUjj43GG+l2wDzJEGgni1/7gdIqAkAvpQo/qT+iqYY+02hqJcnaC8O
/J9YPrSJWUXwcwNZpWGye17igruPCn+fgj2Hj8EwnFLDnEXNiNZ+zQFH1oel6SPLtFmaiL0qOBwD
cy0hU/7J385dIjJuzLZgDKu7rKwPV8hvR2emKg4SULW3RN1tXwfbpaQbHeZ11xyOpfE7YjrNPISw
eRfR/lAs3XRE9GlBmP7ppntF/9ngBMr/ji1HXjLS/dTySarIzHpPJT0z06SDvwx6DfOenmClK8gi
ua6UWIU19C3QrGTkNe5kUD3Mt/74eTbqEKXMIGFY0jKyvrPqdgiG5EqeYbgKEW4dgDJunMgkxslI
IOtVnKWh+qNm0/crVMidyFra0I9NYGjeno0N4LbZGrrTj3h43PCs6I4lznt+aLfyeBaFTsOHl+dI
QOE8dL2jRSTIAse8Q9n4thPjMRdend/RSi9kh4jtIfxfZ5Rs2JrvOUz7mG/qfPAufa1ccf4ndvsU
yBbP1Kfoulh7cmV/PRZU/J6ANr7Z2sYgrAaLOMEQSauWoDWIAvnghbMeIh/a/napktNcEqqBDa1u
sHGLdgtCPUyc5g9toDD2iyNnMwoNYGQoE9Z26RRoBw8hlbTbPJwxSz6T5PuF4gYpHESOZKlBQmZf
qjlBTGj364IpRXVrF/Vvq5WpuZJddDcbgOrB5INFsp7a4bWeWekiplcOmq/gEUdIlEjPtqnWOwke
svbI123YM0UtQm7ok5MPo1J+jDW7Ghp3eRaArPMtyF9Vk1n2JufBrA3HiBxoThS59SVwWTFPAqkz
oZoPPSJeZLbXKqV+wMgBVG/Mt2Uq+By2RoWcWaRaNxQYY3n57eo0Z5TRqJjjms1+Cv4zrU2GW1fH
SbaAbsrTpTbdQ7SGIaXNd1kJkEkfpSzvIeIRbPEcvQlQlpmt1cNiLqeF+/NnNlURa+y0VVwxCsNx
MBzd7aGw3IahVmhxh52Ym70fkTShdw6+ghM1IGScsYMeRydLtUrIX3DYhCkoP76gKV38IE6FYpFa
ZtpBQ/CabaHNApSCOZLomaCLJmw0w5s99FLYsidghA/x4lHfjxY/8lilWq4WBkb5hbZSEGUB11+r
KVxYB3FE9SfVe4JdLsL1yxJ8omYaZHD3yNC0w4fj3DqiPGqljuGGVZo19VksSGW+/9OTbunbn6Fb
vbEmycN8b0ZmjCI0Psz6gNpXx+Pj3pQqffFm+WnBgt1vsi+f7Ivz49QObxb+1zNVVkAvxMbuxX7y
B77KAQmleTLl7FCsoth/7SRewHf0sdYwXK93TTklXfBGSFKYlap2VUs8+12uxgEl6GOpnift50WJ
ETyyXVPAZ3R7ukKkQ1tV27U/85wfh31XLxhTn9Z2ZRLWz4HxPHWH4M79PdqqhIEnNYMqE4+9T0pY
sskq1FDSCv0QGmozof4aEDslslpzqC0rohWHh+o2wVvWfOdpKayzbIOACXxbho2fQOnx+BRIj8cQ
64yCGY1X744fDYCmTFFb7CESdeWdnr/LyEpSrJNhVeJv5of+XDwd73kfVGEDnpkKe+Nx0BTOMs9E
9APQbp5LRXKpFY7/Km7EjsNeKw8NCwvwEsAVJvmEgoiY5A2TifSSkoBKZBCQvIiB7uKK6txEQ8sL
BNfw8YQHtpp7drwRTAURfX36nJS+SgOBA+VKY8vcGPrl92l6LsTbK2kqSPHSV/3eYqiSzotj/cIT
DFRJ/FZly1fzhTwgX1TGkfRCyeSpLyx9HW0w3+EVJlyFx+YiKXE1KqeUNG8VEN/TrZMvQAbmnl/g
bj1ZxfrvWUCYLTNp4GZLXbE0jLMrMEyBB0bDXmD7HC46TXzeaHljxu/yu1lMcbfLTLBgwqWE3K4g
6oJkrPVIjWrFro7rBiFh/kj6pY5fFi2gPLnNBSVFkm+9Pia8b8yrhINLdPbU3Dn0zbLib02uavqQ
MVcChIoxCZ/kBYyyi+pABnPk3o35z8/HdMLcNF+1bO/W2r35rZaNvQL3+WLmVg9nX07z5xxA8hdj
dIIOWsyZFuCz0jfdsSupXo5iFPe1wWkq5aSDkTBBgWCzmdk70Ik+YccV6XGcvmu+IYWhq40E8JHy
gOZbhHJTs2tsK0WUEfWTQjMZkDj8sszfesNoir/oBfr+VY00oRlWCOr8pmaPIDuKP/WVS+ZS+sS4
4b45L18fkDIGBjZ24ddHhEAZwPU5czFNL6BZCZvqgZ52QMxdElWqWf7l1iNc5N1huhjKMbXwvRNV
RH06zMpaxs7r6lJfD6L7sfkGwnoE9X4+bSSprQ/UQhKpvKiT20kwNe9G7StaNQp6XQhWuMWySK7T
1U+j+dAhnMLDDHC62cRury+FUAQnGFQpnxS+I7nsTCFil+TKVAv30QaZHssqtUqwotrYjGglsY+v
LqjzhwDuCaP2TSNXGlwHDks+G5sURmc7YYTAVytFNEJt9FymaLc5sB8E3kYkW43OW/tFueHfd3fe
sIw19eEQJkMjmtHL7ltS+phiIqlmdZyDRfz45q84jDGVB/34+lJjtI1l+/THz8EcZ6kjO+H4fZ+t
BsN0SK4xMAyDXgztTs39wWo16IlP4cwmTsv9R5KBrSvZiA9tuIL8BP2RgVmATKvwgvoLZAL+JI/T
HygQNUolO+w3QJ9N/Zsm+odKcxVuIwhKhzwXY6EO99KF+3AI7nXU29VO9RxvsLKVCTRzi+vwlZ1F
8LWGvDHZXttOSUGejpOJvjDl5Ik9VhLeL36duzp0bK6Lx+WFZpMOVVEJ0aRsU+S24AZCeGo2qMGy
MpC4bxdFSY//3PZcbbk6m3pE8lSMuVXz4mdGUZYWE9DJmgMbT5J5okoFoMpYLZg/60wT3WcRTF8Y
aKM8S4TTrF+lOf+p7Lg3wlAE5c+U+L/8fp4sDg3Lz7BVGe26Prcy0D7IUog7WuqR4n7bNaAK1259
LCa9Pm6Z7o5Gw7xdvD2eZZbjBCjAvTJcLqeae3n9xJuF/ULCTh4ED+Q1io4Ex6Ecoly+ntObNMjS
j+ghP0oZk3O2EvRkCsTy54L6Sh8To4B12V6s+pFiHvmsF93lpk+va/rkx5TZhBZ/u3+ukrGk9jft
4tyx/AKwTUlBBujTg1ecn4dOXKBKFJdOdo1hgy05zRN2959hSMXP2swy9wgEjV9MN1k5Fdd5ZIW9
ngJkRbVaQpx1d83m5YQsnGgPTg2N5DIifeQgpyLtvbT2fOd8lKl8hWn3ZNJiCxXYaMEvAI1i4Zeo
Zhn8kkzX5ClVw/WYP9i6fDiVXNfiuPE9d4M/Kbnaf5QbCAzoCh41kFSZwlS6FzEyMVM0Ugd4Q+OS
XmjBSpYN9BMWUDn0R6dlVCdftEE02+XOgon+mOGa26u3iSHuzjOZsTlTwNiuWas+MHPxZkf1PIrT
vnGzfMJncfultu7FI28J6YpHCK04dJjTPCHWTQp2lPhSa/UwR3zJroxWEK6+KjKFem2oQHzKKe7G
PtgnIAesLBYGor7Hy/bZ9T1w9RJjL6hdoDa5OjR/MzwgvVmwIhUzR15tbtQqAy+FTZ8B9bud9LsE
DmHIJWkapT88yE+VNf2r3qfhPOw9IhY9zXrxJqa7si3qfLSx18khMm26EkvG93O9iuYcfjF8pskr
n44AQWMs7xAYV3tV6UzvlUFc3avnh7/XVIZmbJ2f2gbfj2ev9acLZKiW1MV9MLRA0ld2AxsEFBfw
B5SSlKXRna6Xmq+41x9Ocz/P/wJ7LqwMNguP0KMlE4+MXzuaJ7wxWea+zLVp21eW36AhjrJW8xpG
RMRF9JkbkBpOX+kkmXQ4S41mk5cDOLhYiyF7ASElYeAtrLjjOEgKDOGkC44lAyB8RZDMMutqIWu8
q7vqNVroGt9D34hCV8CC0RLE1P5DPOwiegZRBqH+J9JawNT1cWHQ+5iLfnay6se8gWWhFEupf3Fm
qSM0o9iWlEUPVnURySmthhZOiZiK1LJMfp/gT0DnHoQJQkDMboMxnD/sgx5RLxUYDXxuZTPlqzQd
47NBkY8QnUDDQlA/FjtoVNA4cehdCcKYvWX+ms4pSswjTFN6jBROpdzX3dtO6tEKZGLX1qznDloD
EZqeKRBn279MEBiJchmapYRN1TpZJevsLHZLCvvu9dvRo9XuFwkGrafeSKR4dDlCuPP5Or1Fg+v6
GgbJ+U7G4T5173mj369HjII0eXfW3uoAd+rYhpp5xYXd+fwPakSxfeW9KjdeXEHEB/mHCUUBylZP
X0WVqT1/4Su85HeOndoj4aADdD13HJZsDxOt15mq688XmirIKQnKAz2TmwcCeU09al1xUf5Cob2K
LoCDSZIY/GXup0e4nH9WB4TbJ4RmML2PmlWIBio7lo4TxKL8hPshCBcAY1RiLdgVk9RUh6UAM64R
3aw6cl9ZW6sLXkZ5pMqEMlP3XTcRc7a9RzlG6hTAQBtuD4K3yq9MPpbY+TEvwWvIB94khZ9mpq4A
8soUT3lPyYi/bMMpPRv9BKXfGrbd3rqWb6eqsIdsYGImSAOPfrvaU+kLCDhvp65kAXiA8cEKeZ01
qPtj7lX9rWmDNuhAfsp9311UDBKWUJFiCN8SJPDiyxxiDXpeEQrVEnWjkjw0GHmQVmMJymxtM3fK
ho8u/vOifmOPSCytbJdwcR2mRgPOKmzbmk0wG5o/tOYJdtSExW2AdZsRN/DoPYbQQh6SxrH7LN/c
Lp0iItnWAB1ZdgiTFMz3fJUIWySRukuy8bgzJmWQBDHiFY1XAfxsD+jKMIvLpzSjh4+OOQeLIINd
xDD+dX58CuTtKG3nlAiy6AnaC8frQRrNJM6psnOCj204cjBJcFgz4cU/Hka4ch1BzmOU5kEE7vgh
jQPQifn4jShg6ySQv4sS1tqhRu5Voylt8azdLxOOpVFu4HvX8PRr6w+/lKRtto63ZqDzltykewlT
/1+TYKbr5uzji++y/SzDUbMKk+Xl8YJHJLoYsE8OVLX43U5SZhXhKU2eGXFBlXMOpyK3ygCTfFuo
2PLRJbKg1E12hNKR2q9BhM9FiSVkkERYhmqQjQyb7NL5+vEsOAvk8ThULAZ+0u/6VBKZ/r/Zi5lz
RzpdKcmz8INfqDrMZrMAjoXcUrCh4RExf1ToIwoUots43R+Bk9vONlPBvYkUDC2UyZNXA/wsMdiw
SbPQGCE1MGomen9DXg8G4PLU7ycRkjNWdNuqEH6HFs6QRHioETmhJrHQXxA0uKl7WiCrtgR7NyJ6
YhhUZL2OD5Q/SjnRovHUlABhborAlXBhvGvLRwXI4Ze5TZXuRWUMmnu9EuQ6hrW50JkDq5yDz/C3
jpYlHrpYgYWDI3bOp/dynJ+AF2o5oBQC8enNYr1SXHYNMNFa08phJccE9Qaw6n7kjAdYFL3ItOqU
LWpEnfkkkpHQ7kOnQR/s7muw9KSyxilNI1HZGEDRlzhN7Bsl90/+ap7Gx8VvFowW5DyoPcmUqMvO
5KjWmXI2sr8aXg+5WQ1tbfMG/QvKE1HNEL/JnjMUHBTVGf/2K9EBmg0rXG8hnsPTXixM1GLEWG4O
slHYCBmLCbu9qQL/p24pE7Jtgu3g37XatRtM4/eyHqLp/6ZxyG9VIL4v+Qj8aFS9eyOZD9buMpH3
5kgzTFY3Yz6o0whTBHQkBPiVaKSTTeCtSSnzquQwUmp+dsGA4rH2FsiKlUPJrZNm2C+6IuSimHPR
Jt7SMcpJ6JoPmsqPxB01AFjjuAt5/GiGG0xyN28PPG5GULh8Dk/pKFbs+C8mmwbqJglvvAmYvNV+
lJ63cTi4o0PIPLwERdBnE+AB7jMOJFRgZCEPm4iZH3nqf6JlQsFXSiQTVZ4ts1pS1Ij3F+wqmUFJ
lCRi/PpQQ3OH8LcLkizfUfRGNzGklgMcX4gnQzbF2RevEzU5W8d731RjfNoUC9EfcoCbytPp/DZD
Wr3LVuqDwjsnoo9v6/sHh285RlCpeABkcB/8i5XQgi/7lIL8dx6MtdPq4EvA4e/Ra8aY5g0G4sAi
70D0bDUlD44jsZSR08OBsCs9uU2wAtDN0vsRga2Ow3LdXPBokmeU1I0pDs+CuBiInS92c3x7M5C8
sZsoVzdYih85OsYkxLKLjpyTBTOoKHyvpMC9KMoBJ8+DU/L2IIBx7KFQDDEcLfhs0n9iXAvGyvZ2
85JWtB/LNgNcQL2sc0BozknZFSrNM1d9bX2R3hw2APAlg8w0Ys0jGrXGyWDZUK+xGMXO5X2Vczss
sDT/oP6tDqcKMopEFuiCALZ/cVYzZsUD4lBKpQ2zpnT5Hvbc1iDXPPm4I4vO3ndhXMQOpKHrQPmW
jcKuj9dGnALlKORTTBuZoH+7s+5nlcDvMKMJlSd4MecPLW03iaGs1Z80tZa1FwvZ5/YeFAnIbiSr
b/r5LYlxWyJFrUps2U1rpH/HNvb8Ibn1j4VzEgDlF5a0ypfuNBklf9txqKcIFzDJLWq8RC5XioRm
kPVCE/CKcAArxhTTKVxuZkt2PXzqy99RZPynDShkXN0AYtTDaqPRw2VLzVAbsJUUezSQglgaGsYf
OzakAyJwIfrTJe54wPg7Avbdk/PzPwS4haTECs7UfRQWgmnrtlo61t9jig06ghPNp8NLdvgu511a
jtnis6kMKPxsMzz9Q463Gdj8MHjTfNa+qNmnfDSI/5dv8/0aZ6woEF88Yw+D3GXzBYQwjTggff1N
Yt9s04+upWQV5ji9yAvbfNIslzQ9c4J4lSPDZRcERPrbIIzdEvX+6Oky9npEbZndmLpE28Ao1NUH
S3ZEpIVssaLFs0TrvugR4AQfvYMgv/TbL3ckybhyaeNBwa5JbVtNmFRWR6hGfU8gGCaMjrIpdWs0
EwghqLg1k5/Oytt3kp9S5Exq/51wvtXcxwLPYu17ZzpRriNd1pJfRlQGtfI/Q0sNYInXCaEOqqT5
yUhPn4bOFtLAuxhRjBXCyKO8z31iQlwGb/7BUsHyeWhEcXegjC/4ILWT2ZWB6DjgykRAFrEBAVKE
woqZ4UVxeqHOV+9zQr17Bk+tQ/FSMp9iUol2swfSv6aTyFrRmbSvBLgpsk/Hp2D1+br/BDLGL78c
noHbLB0cxlo+lTeQKWp1sjWfLxESCwq9EMVKdywglQ3HyBfi6B3ECtk0cwpL80Hp3lNWkyEqXGQ+
qk171yWfEZbGgRylJsbQzm4MuQqPMOyYp7udnWvz5QAT6IN/uuXLjJKZvHFlWMSp5n+CtAKrKhVT
LqH75ru+3hqhiOMp0cMcr7DJm4/DP9l1K7FfS4UlcXk+84465Favomm1xEEFaFUeLOxv3vOTEA0S
rgb2XDzwlYuH/sEgdMPetVvboN0G9WwVjJ2aA2of0+BPJ3FLm7scIxk1B6PhpaCAKpHUAHQrRNF5
YLieCMSAeofmueEkgIXzrTN740SQ++hm8LiBsi78D+RlV+m5SUPl/eTEs4D/cVq6z3+ol1YvhiIH
oZtMq6vEDv8NDY0DdwkikSH5yrQGB1CMx9za9XNJEaGEemSIhfowhI7jHhBabRP04JzNyofldmEU
bbAg/HLrjHXHxYcqHXZPn5qdzsDjybOeNbQZKL1D7aH/CY9eKSo06Zep7I9rJoodNxZEmF4rbn2w
3r/4hpt8bcoZSO8sk9Zv242DW+PEccC5DLhaK6JKXCIjLaUXa00G5B3cLVk8nhcIg01bZ7fCkbwF
8pOgzoAZIwecY1G7jgry8aNEh4ReXQX8urNduPzgFZK8OsNrO6BdMl/+k8akFj1NiGQtyGIL329W
kxSas/ddbpDxDE8jUCjBpD1drrYd4OTL2fBXnf/zR1uFOr4hLxoDKe+F7ivati7T2M0S36/vuiMj
xgudNVxhTYjKYYTPNiiiqv78aSQOMYsVwOp/z+wdFwYGvfarPk7b6uZCtG4RDTzZSbbfkW2gmUAU
CZRPVA+c9AZcNoPEnpfaZiQ4drpjc8SkyFsaBzxpnwS4buRJNZ/ElZGi6ucvIk7C0mjBGGsh6vP2
1la7V9+TaQEPZqJEnF5JLZnt4Zzl45uhvgs53iEo+ymt5W8mMJ+lh9s6Iqxx4Tq3yxxKPyJEoTpa
14yqIK7wapgsA7JchUSQl3fJLgwAz8ATQLXy1VxceZRvFYVNJkTOh7Zhjhv+RowP6b/SbKBlYPzc
zSJuq/FScXyd+Q8NerOYGggI6qB0Sg8dUrH/hqIEUCElZip0smpsPtUeLVO6NVWyzdmrhvAl/B5P
oz+zmzyAMWwejagSEg0hPsRywn1ikl9GKZguUrWPM4f4MOLXgUX7/5WKrY/i0TRDonVmIf6SzjND
a4gvWl1GtLtPeKZU+dTWiksVWjaeQlikvGTIgyDdcxTTuB7aWVRBGnlJeCvy+x6qhPImlZltj1O+
nRY619QMbfn3UQxg0oSovfDSQ9Eigytn9qjHht8GcDoqkF1TnE8MyDBAyzW6TSpDEzw+yjN1WoKT
dpaJWzYs8Q95R/Yfdch6Rln3/qcz2bpsUMAbRTdZ8I4Ax8LDaA1CcE8kQBhI8zX5WutpLkAMgoFv
RA/HPdGIOWFFra5TBCDHII1ziGPH0aO1J24wsoyEZXXBEhGVLrNZSyUMdyy+nEyFuMLMHJ7WYyec
6wMBnoTlZ1zI4zh1yFBXIE/PeMKB8BnQMlXk9iM2h/41YDDQjC5iqTtqBVK8ivAHXARPw2Nifcpv
RtL257CD1e56pHM6IoO8GroXEXM3e+rqAdNsqlbc9m9N1wFOWdxaGAGXPC1RwcNIMC5XuofcP3WV
E/SWaz70jhpbGP3zDmqJJcmsBzbvsFcMtQVuICgoYTvkVKTQ7nJp05JUMfNeAk44WQM1iqqS6Qw0
wRt5e6KvhmMqifnm4201vVjvPiUMTHeoZqxmnDP5XVgwOnzWNZjA6RfUWKz5scyXVTtLWpcPvIvU
grt91y1rb8HSM4MfBBOeoS8pLJCe4TYDCJxMEA2ckFsAYvYyUj2QUCsT4WWYpEmmIWP9zMjqolNz
rYz4cV0+9DZfOVrBRclzQ5D26jZ6T4Mmyi4NuqAnw2OEiIeuqxGAliOn4XTNp/aAfG0pQf+ACt3q
rYeZRkpRrntjcz2Gl36DWBPfn6KWzwzS0KtX66dBrLdb1Qrhm21jG8+CDjm5IkLlNb5skjmnD6Am
N0xOULX7V312gIu3i2nzrxPusqvojE5q1gBTFdSOxyzqIwtgTkHr0/WPN9lEbKwhRE2tkC9VyUg6
NDgkwiAJzZzZA6ZuM2oVmSKCBwo7Z+5SfsAl03WKzN0oVulM78k6PmU1pfaT89xw3HfJdTP+rVms
EqIXv7Vq8BtVJ6QWqqg9hnm2THJ0nnLi0Ost+iMFbFjPLXm7lmWEt1VAAPdNqvWI9Dt0jAU+1E4w
Rhp+eXDdxBpInbd461vPFNEIFvvSSVpHMdwYeZthlpPAssc7JZj4gUfv+rch59yq+21uVmChoHch
zif6CHa9YVBZxQXKHRYs/osxagb37c2/kQvaGxbo7fnPmOkgzJXu07oFSL6cmqQbF2BioqiYGI/0
z/1dBSeQSzdMZVmyu+ZCj7nBCZPXOadNFe1Jg59cYCw938ug+O0ECa1iea/xssa3tKBG8FJyofeL
TG5iw3oKvIOyspBlOQvg8DXlyng2mMS03J2EEGxuOua3qT5d2vxAZ6r8j3CkpnB32lxHndg+rsa7
TswOlHbA9YdaLf1tIdP5UkeqmwucG5CEfFWB4mrQUrl2hHGT9v8w9FWoMXKzqj7oRTTXyUqiSkoN
DxKCJ9Yu3Y0UR7EQZcSNRRxP+fQ7QSqWfrQK1hBDtwTMwKqhPMbXFInZhsrx8wvVOmO0lEx/2WpU
FfN3Ux1xlenSYbZ7iZew71DpDHHsUqXwaTFDLbhYybm1/7uFs+7IxuFyOcmOmoSX2YlIAva4u53G
Uecnk9uIFTQceqKlb5mEcu30zl1lQFAiem3oTZ/H07cpBmTB9L86RoPg34fYw+W+ooPvVEnptobV
y/QPBiI2GmBwYfsxN7pk86eyEB9lDYol8//MGMeeh7AJWhRBIzRAgmyHBzK5DTbfo1NyVuxaM1jS
JdyLxZlOaPJeGdwtHaz87SCvE83uaclvTO7jcw8EqVGAQqm0Pp2Cc3DYu4urx27YhRzsOTwikq7h
7DYlpKadk4dPoerfGzre2fcGKc+A2lruCgnnHMpg8a9XCyKCalaufP85IHXGuUOoc3wuLb7rrm8m
6XpiSVA6BGvrB+O+i5kfss6c6ZEQ+idFpRY+E/Zc6AoY97VMPhUoIB8nOHyGy/2g6mVnDBHnVqou
OOfRiX5rUbSdi02jomnwWTGCEj6qV+EC5MqkyFqzHJ4V+7Tuxceeb+FPqHEYQ10RdmIv+v3r8Z1B
Ipdek0gCTclNaFpA8Jli/w+ziHSz3U8Fi3LuYnGdMLEWfMTpGooSOGZ3OPk2e3oZcHrrExmP7elB
tggjF7EJVF5VDzS/5vG7NxhEG+nh1vx2kbRgG6WmokUQZj4K2+3jQaK2WMbaOymtjwstQ9H1vLDT
0lin49sXfnm4q6IXbzxwVikg007RYBHSjlmqvL6OYCGelrsIlFbolMlKjFwWI5eLXMqL/hQje53I
bjzMJqNpj43oqTFejhad3gQY9lFgepM/uFx0IZNxbmi+pk3AxNp2gBuIDEjhaC+YS6IskU6vGZEV
QYigNFllRFsWhac44D/cC88tLwZUxe7z5xOrtNEizJ6K6mrO7530BiR0tLjqWbtN1kVOkz9V3P/F
9omFvJCuodHKICrQ5RZR6ZMAyBzp5rsyeboNWfHDySM8d72JRpVt+rXfw6ZYVTLDG6/JkEkln+e7
dDkKYs2gheVaqcTfa9gQTSL+gDBBxeWPfiwj7pRMBKAWeAw7RKWIMnbp7dnFrubb6LWlKLQx02oO
YKAZISUDZ3SGJ7Rz+q2Qc2kCRJAAVasq/dCIqwiQdHs6Nr2XANiN7AgK375jWlDdefCXIstfxixL
Bu1+D0eWDo/dFtqzzO2s7F1ukvgmLMNRrgCbfZeBD8p5TuCKjdAwxhuHfgHlrGB3/wNgej+2vr76
pODbIuEOUsGoynyyEukhGtcY8JnMjJmmTHKJP2Mc7MG6V0egvvfWFUYQT5nfZHQmwxkOhjkcUD+A
6wgGrBqnJ/erw/iW6wK5X6P6RlNsi/dMLO0yU5U9p4IrfkVlGrc4mbi0p8tDm+NWLSrsge+9lh3/
4wO0JnheIZRDe13Yq+c2j4+iURp5Oju7+VS0zYUiqNZmucRUAaySAx0D5lQZ9+PgbBFiP827yDVX
q4eKjngQfBYu9przXjqat5x4xFZ2RzUFcvGr2PJqy8679yDkIRecy5Xv19rkpibrlwiKyH3ZZMW6
1k82wZTu8FA7sGVMNaDSGe3SCOwRYBN7L93OLrHwDGeB1MSZWBMyoVBZ5IkwwgLdZuCmBkKE6RMp
QJmgCo2QyMVfZyxsdvYS4/cTR9Mihz/VLkt8uQNu3D0AdaOTuOaTHd9doSmj5ujM+BP7NyvrWAhT
vCxNl4xljZi9jWMBAxU/ejEGfqkCRF8wHkWLwwXdwbPuRi+tRLQsXQAZEDh+GVx9Z5MwD6w1wz6O
lVQU+B+wgKgSGVbabnPnQ27HcvWYv36TLXph7fmhFkCX0nYIIP9HrjjKAmMAcJW5KDZrCFaoT6DI
C6nygCRVRKZpYqBHj667gkovY8br1xG9b5iICswUPjDkTIWDwPvt4eJ8Owl6pwf0Wca966J0/CB/
Ul5guJAfsSpxi84mfWr0QXGY37I7j6q/sMNowKnZHyUH7CyWBtB9nxV8JrnCfURZI9IXEEQgCoNr
44SoS/qEbi9I59Bj/D5Rwu9vIbgVa2bFTbxKMMLqP15vMtNohwM1f36jDyPQA8qLc9OrnvoE2K0P
7/R5ZnX76PkH+GglzzGsZFQm7AyA0iT5nXg1X5lI5B+KL5vlwCPN9vxkb7HoNm4nXfQPyHcTH+Io
L8YswofobbKq/dQc+pmKnjpCgCKR15av888LnP4PfmxPrOvzaERzAV93D1wdPhvgMbls8N+p6fny
ANhiJtsOiOipDyqhIA1ecrG3YN45Buv9Y/gfArNNONwfoh7rLw2O2ySglrKT7Ii4awgcRMgV00F5
XeU59u3rN+bqq5qX9hVTPrWhpX5eqk7e2KXK5xAoGaTgRwigaqRROD9aFe4GdSSdfpwD+oS1IS6Z
zXEDd6vxDexMHzxdqvRJpSFMct8FPJKky1T6ll2BOpOtm278lZEo+Jeh/1Ex6MWCg6q+6s+j20z2
hJUYVG8bIuwsl6PW6/4cgbZhjO7jODC/8sgJqhMZmvasm4CJFLLN8B2bsnB78mCnnpaaH/NzuEim
XHHkZyTIth1xS4Z6SbvRIKpHg87wxfYL/rzu8xtGQOoWQwiWHjncX+GeaK9aO0yxjGzE7jCJlbTF
+Dy6ijXGhu3MLTFvH0HDl25fFQsaKKJEUmraJyg2YOtmMmzrwH9M68ugOILwlqPoweQnT4tPJRbU
r8fGyh1C5MJmrXoGRGN+op9be7c/opO0O/vzNCnBQkuyiKxFdIx/aPCrYankj1O+ELg2RniRDYXI
1Zpg6ga++G8HSQ/op6sypw22Kck5uI8B7CbWmtn2Ib+3v2SY3SlBXfKCpOrJ5eiQRSV0smDR9Mtw
4Xi8K7Swxlws0Z4C2UIp18FNq5J2e6RDWiXVE8IpK1MkKNWr5VM+rU7qZ2S6KcdKpgmcZGsKpS7k
WAUkJr3/pNy3IrwFsmN1JTDcv2CCZZypJxIM/tFJ44xdtxs6iPee1X7TnxNNayLpBhiYy7J6w/uX
oTVAxD1MoNA0ghU5Ihfk6k2uxV8txNWOpOgj+uxXAAmcSeSL5jbLs3QwaEJOEVkt+r6IXH+hskA4
UmMMSXZd/XwnYbd8TTxDVyS7J1wYW31F3EnKQrxJCC2Ke2Shlcz5luvHvitsezqkiSWElQn31I8L
x/gvA9zxsZpjudGG9aBxkWTLZ71osQD/q7twwi18tvf6spLOAKFQwi+5uEkrFLy60lAbcwx2mpOs
u7GQ5g1gyghML3NgjMUb7YaFg/8xsTzUvyHozuEQYnmGd9jf4FaqAr5DJY+wTlh79cYUCE6wTEur
towBaufIrCSxvJzax2XYgd521RbAsqayq2gSFyUc0nuQMB3P+kgmT9dxfNTH8UM51hTs9vg3GM35
AekgzqlL8uBLk+PHlRBp/3PEAiymfGQBMJT/69ENoTI8RdSubTHaFLHwlSqeMMjzqjUwAlN/BalS
HwitK76zEmKqdKyui9dg1rDm1ZW4cqiRGR5fHhznIFbXucrBd2YqBS1TmbTMXKMJciSRzn7tBtuJ
8m/HHWXTlaheJ4o+s0ZmB0FxHpP+Gf5emWdp0X+C6FRb4xiyx7HuIOGuzWzFL5EPK2fIlSwx3qJ7
xWAPq73y/79XoMYxGA28zF/6e5oqBytowsdNunAnsRZkRtYcpCdnXAJLqmG7s8fw4TtXlfAcBW6H
RWCeP/W8gQOiN2OQQYHix31pPJg0So1/XxARoeHONS9rBIz1T+H4U5QVA01W1jIl6RV73ntEjliG
Roy8DZRSkEkOTvWpqo2f0XWU3eSKvRDOHtjnQD4ZudlAtw3y4StbXyc+qIWBXWY/HJ2M6u3PXg/+
+mTCbmyqU4C4th2E8Zde35bi4J7FYCoU22clNweUBKlv3RH03EFn9Hc+12V14S80LVMv6z1m8C8J
TFeAP+jsjBx7XlZ8X6X4seRVedCxwGvarxgEZ+tLeWaAXWEThUyrB6gkbQbzwUQGBagYFM06CXr4
dx0r08vJYbymN3v/vWZxTosflJAJxLpIg4sej+Dux3LTI+g6TC5BwXXqFN4br7ohW4PocVZo7/Pb
XSZeqnvnOoTOeegyKl5cjTg2LW/hooP7O3LMH4StP8RCeFNk/RWqHDP2p25mb3abtvb6nUdAUqeY
6J+1czMZ1TtDJtbCQ2U8wNeiLOka588fJDD57Z24aBsAsZAcy4Gyg9VhxbDBmud/PwZSFuX0UGXj
xAopZyA8NAAqRUUw8UVTLimDxNUYMKs/rKCVYWkITAkhN68CaCJXmWMV3HedF0oWEL2ddDHmojG5
HKb3prAEQhL4y+LKdrfvwarSCtLTOFtGRON3K2BoIYHUAkgH59BsGG8JxeHK377oQKNzFbwOOU6P
WAIpoTimY2nge1f44kSKRn4jUsTl4lCGWFcYzCrq6TP4A3ZYVm5tS+qn8x+iaLHDNT0PSdeouwqT
t51AMv9rwFjImzRdBQJTssurLEa4p2XeI844kf4QMZvoytevFoROaU2yDPynAWDDy2nQqb9GUU71
n9fmaqEo+0+OTx7O1Z3x+c9nMBPiv+b1mHJ1NSOZQPz2+E+Wd63Yh1DBhejU5wWbr9fAfVMInF2H
bFAKoPYmT1sbFAMwDrVuAWAwXWydBuzptpWF0FXHHiBJcc5eI/ZTz1zj0wQkYDBFgrBFec6ewq2s
BHVONhKDa5TecMEO/r9d7gKhLygiVbsdyVpmYr9V3GWjd2lnpY1cQVIfoT9UNs7aKtuyIPeRC3bh
Hl1MnzPupBBGQhAgtRhrWywy1aw1miY0xm0mY+Ssw2ZR1/pVSj2AaC1ZXo4pDF7YTCadeBZiYNcG
JLm2CR3/hZVlsYEXhyw6hAGMGGSSIXp3+nJMJi+Zyn/Y+I099zL+O9OV/oTw7xx9JGJCfdUFY4UJ
7okwOA3Zk3nHwpvJ/8kWeAT6u792t9XOcd7jIvWAhixgNIgMRdPAZRInNFcD656+lOv+tAsr4IdR
FW2XaNfMsaZ1CJ8GYHzEnsP6IJlu+nLI1kI9ydgFpGuPqnbVJP940eb1ZlEQ6M3nAhnkReC6Tngn
9e7j1Z5LHT8nnNLhFNFtBFEQeEwmz7XvjEXsi0YOcsIg282L2phfMmgqRqGV495ODG9a47hCKiHA
ZoAOadVAJHK+BzVPmeyFsFQkVLUAx3CvtSiD8ibQvVPNWpE8gAZfxteaOZARBGRFvpRUSXxLWzgg
DSRkYHalsa6aJVMmkrA0S9tB+tl0VaudZYy0OhbM1NBWc3alaTKf/nPxF2WWvHeUv4G6YSnGkL3C
2k+msHcUyzPFQmDx8f63xN3DBOeKFZsi0SxJKYtC1ZSFXZ02qHXS2XHxpHUi1ZF0djVFvFDgROSR
9DGtbtPZMIvqeHclI8uj/aL7lK3Vty2dazwBmQxpSQ1pgWhWT09XmtCyd1IrOLawZtbskiH/eRDU
wTspWZtobZif0ITklt+QiNsUo4op7WBS/ES0bTeQUrK8kdI+fT8BbeA0Kqs/hfuWOpS5BC8aeBcY
LbFbc3mIIBe8lIv7YIBUPMsTc4vi+msLyv4PkGCz4u8yi+ZbDBgMrKXkSXq7OM6O5AvmWMA0g/J/
F8KAoiLDFlRVqyRgdCFPfprHbH58CVr+RXIWzigw/VteJ/oXKzD+Us1310y4C8GTQ84YRUy2Eu5V
3CoMU5pWdipyygUD58YspfPOcIlony+a8YMwBLVxyPU1AKFHIlnp510i9SvGXQnzyfr+Yj4Sz48w
nVBx9u63UBesPljUPc7VPEP4FUwQdUzM/maKAjGIMamkM5QU2oW1g7cAWxLvCsCFNLLH4DuDnK1e
8elKjmnQZ/GGDdkJ6aicnLHQ6Aut+Ay3iNOsL26NTRBEf+xuEz/Ky6a2X02+h5MFBprjzgAo4GgJ
pDyI7qon1UAjjui96ui9CU9u1a4wrJCRg5pedEAgLOHt6r3PNdgB1diPuv0Vl9KY1nRkJdfGuc/7
Lm5Ll++U/Q7gXzjWCNn2Sr9nOHVPQVD8Ea9xkQ7coGZOctn1yr0FP1jrdSGTtpNJgCR1OUQFZxYx
qOisQ1Y30o6+6gw0L797QqaHV5v5s/hmG29hys8CdhBbwSaaX2qqXaXd7mRHUT+6DQsVVxncOn9u
wWA3NHOIcZ+jzc+0TYMznLzlrRIn6pZ0oG8gXVU+axLtAe/k8CNcYmgCSgPWpjaMfc0AjlGVB3O/
b4TttQexPEzyOobCmE4DUT8/ppw2++lmtIi9reUy4AASNRBBTpGFbRaY2NEVXzCVhEX04Vn7OCYG
Zgrxd8irQjMykLecy8i/JOAmBzKGXG0jjJXjM0MT2k1VEpkgbnSLweOEF5DbVXAD/KGpJ9W5gzoo
sLEQqTq8v4tBhwYQk1fEAUSKXwwVpZYn/g7o/SFh92lVSRywiNvRKMpCm2okaiSdwiBOSICN/nF9
uh6I8fkaJS7yuqEC9nTBDQNpbHvC6EBv2BuFWeojQj3IUcgDAOXyOnJ79Kr262wPYU6JXGL8JLFN
px1m6SCT/956OsLemystqAv6iGEwpDNQIdl4bfOJOIzlNyNVNE5B81CNpQY+LgjJwh4wbBq5+jev
qbOS3XWAJ8L3EBBFpwy+O/uWDBqAp4wdwXDjajqcRtozwGgdJhTmq9jotbVpLXU6JYIKKPJXrt+8
mQDZczqA2myGQuT+hbKDifC+nsEBqWnIAJRvLWBfxapb5eDqqWZcHCTzPGnV/b87duGg2MDqUX7u
WzalAUB/DQd8OJJ7G15QtlqcWUalO3Wcwmpn9c9k4m2Nryu/asvuGUSXzoXpivmnyrl7vjCBMSeu
WgKyGi/a0e5FGYEJWSlsMH3qSg1yTA9kiMqUJDo9ac7YRQYPWGIPgq94R8mOpJpeK+45Cc4g2xUH
rD86ssomv3MmZ3z+5qFx6UH/EyL7l0xHTHY7crumWO9CYjbSOfie4kxcg7cEpC04w0owguwYFNlh
H5PED/nWzGVmCeKY/+1e7EfPS1j7Ny8hYmHhWKEHm32ex6xVyVZrfcK0KVxQjUUlBgmfbR06jyDI
0BvThAWq/Gi/RexLwsoPG8JklQ2rtrBnl1nFVnV/A7n4RqF8X5Phz85QPCJwm4cQc6Pv/ABBdys9
Vyh7A5TRlB+zjAAOC99lpRlsBNNgDhL2x4VcrijguNjgEJPR39z6cLM/KH5jI1D5Gp6ZqVgi7Bbg
H5bXXs7ujKGCevbsO9M+B+DmozJkCDQvghy6NVDSpgbnTYcNb5MXXtyGsFJLbwsaXMc4SRlQ4sGM
o30kvHoM5nxL3CFvwO/q6KogVsHhvT0+tS0fk1UNkxJT7xNyQSmroyG4J+D1cYs3NPak1tSspZiS
aNA+71Azq4qlms5LixEIYzTJyp5n2DtzYyc2CCt4TNko2JaF12rSj37HguNWeluzYgC6fNFuMkMb
qjO/g2YzUlPUKPeiJ16g7U88osFKzzArfAoqssbXQ2IQwpniLnI/M4jMgg/2FpOviD05mWZe5LfL
u9Hwe3GozoOy2bgX4ONPjMfmS4D/nA/XcS2Ydi3gqSCnSPbgCB9zl5uRHnnoONRzr6kU2DPxtxO3
vDAOBzqlvi1bnqrrcrx+z62mKvJ32PTEuYRX7lLWWRm7jDjwyfIg3xWegMas7Ro5APsCaTqy8+VO
E3fTFftcDM6EHjfjG22eh0Z+H3Wi+vgziUL87D7srZaWpRnqxhtaq+cb/dbXpZqOC3ZXqf9YMGL/
kUqyGMYU9nUreLCZpABKBTySNDmSIBjIV31enxKW9xlNT7tOzyAVeh4UmSJVVRDmXtrWfSvCvkiF
4UY4kq+LuL1FonH3uuXzNa/Pl+0K6/1Hz+5zRJIW10TOdTYdZv+aIcLwyocpKwh9Q4iZWj0T9CbF
a0IxhfXkCsc+mCffi4dGDZR1Inh92mPYnJcyvi5Mfhkhf6fkkb61I+nN++hNNP2zyZH3C301JD3e
/+Z80Wu9T2MbXFKUXuyA/YnbsjdKYarrivEFgRTv/I1JiVEyVIzZXnGuwWpW4e9UAT/6d8a4biMY
/IzxIvkw51V3bKnAQTW7dRxmo++gl++6nPTztq6LEYtyaJWsRzkNgTajlUNSqo7qMKnzBpP0rcN2
8j9ye9reP0eS9FWfhkpMXQ4lm39zQ1xq6k3Ajx75sYcbqWvp/zFP9bXTwMJZ+eAgorB3HNP5CbBh
p1XOdUuT+5Mq+kg7gNUW6+vGk+VZ47ImEN5ih2Wxg+QMPT2ZrSa645K0/vjfQrXDvj5UiEZU9fiF
TSsPn0Pux/TraaKyCRWQyYAd/pidnLEFR9ewhS1M+hGH5EHXZXOoMs592GS6BvRbZa+gFkwGQM4+
F48pBAPNT2WKsJdrCoJjKdmh08XXrdGOuhT+zXFComlyDNHXupOVwnz/LybuY635pm1vgkMB0GiG
mxefEwPT/YB/h/P1EHaeWz4uBxcfUdvW75QuoB+FSmHfBcWVZdIMb2YDZ1HGLZ+egFYxW85sSBqk
MOBmZzaW0TRZNDiiXakQeRY3IzoGHe1TyW9CMOcGnC0WzrSmswMi7W4AImPCErTw2p9ry032ASbj
SzSaud3Uauj4GLq1BPJn5EbMFEBIcr4onTB109YPAbQf33AKqLaTFuNK5eZVp8WV+NdIVwITsIIO
NSwlnSeqcI7097hl4M9VkabkAmlrB4wZfKw73poS1g/KpdisW2qFkPd8NExamklIiE2H3+moBG2C
NvGsZsIrBxm6TwJ74j+Q3xrbjmtYQ8JysqF5M87NXV8qnO6+i0GdC0mip8zATNTcpzvhnqHD2B1A
a7s7PUN21t00Pfvd50iBc/P3rZhZc8o9KjkTZRAnPKroNo21uuZpbYIalCp6tnnaMwBs5TaHrVzZ
SlBoDpxP4PJdjHwHES/epQRZZTVBhaj9Jbukjtsv1VDGRru4bGBTdUXR/API7xRnb7iRK6j7PMaM
z42UcdBO8E3Dp6uBMgN4Qn5YARtrWGuPK0vAL7goKs9oGQZoQMXFunqUuQc2Gjbv8XB/m/rt3STV
B1lPeg2YiS0hMLhCHizhXgpADHBqWUk00toLq5JH82r+LxqS7YUwCHeBPZYtfFT0wNGiyReaI2nr
+x5RQzfx6DlKYNGY4Q17p/nPd0Df85v3uqMjb/kwkLWcCsV2rJaSH8l2vhekTo2XxvPjZsKRyYL2
4rg90HC4rxG/d9QA3J9Z7X01slhla5l4bmKc4/Yw0aj/LLFQ0YEXdx3s9jvJwq/DRsXtRkDEZWA/
40lF13JzmgEV10hJQ6JOhMj2iDuNswdKZR8p7Jcwb3gzEFAJTnUWHMbTUjztvtmbmf6ow9AMAbCE
gaao7v8lZeSxsHl1i33wa8UKDR1+KjAiziGcnLBuec2PxORe8c0EZrqxylSMnb0/V4Tt2TpwIxWB
W8Rxv1gDetsI/4KU+boJzkd0BtFFxZ9dXqRWcU26Hl6J7spLFKOfPSOJrJJjERLASB0msIB7gBQg
uRcYeHT50md8SDl826pFMLSCLch5rwgEP7RTqZWNyQXF7sntOEWoo+vqChroN70G7yXZmbXEVqAH
0t3QvVKMbgT3gCdGJLj7oKaP28RGwhNl7ufVfSeee+73XazfKZ1YMxrN4+qzSQxE/IXV/UU0L9sg
ktKo3H6tHHlT7o8uQTDC+Y35hkmALHZ3WrjTVQpv7Zo+No6/tM06hwO9PZbkSsfpKezKoLtFhIvg
OC6qTwySXjp/4WE0oD/vK+3D5JUMZKsh11pGZTnWv4FIvUez6KyYl6Db94/L9BORZ+lJpxbgMG/R
+CNgsTok9o74cRBvsTMgP4oDB6o5G/X3YZlVsA+ueeHA8j/IICx+MY+86SUpLeRNdhxXpvK6kvEx
MQS9SAo6wHAySDCUCvwN3M86WdsXk78Y7gQ1o8RqFq80PEWgQB3ihrDpxO5Q8LbRmR0QQX5N2uKu
r3l16ApWEEaiPE494366bK9GJmoZJW98jDPCGBcXUpeJSQP8x73bg+stC1WgI1J3RlvMzs2vguDa
1Ke2HbQVI+ycB/nNseK4RCSoQ2sOympT4QfxfVcicxkVpMRfOX/4cJ6tbd0IMhzyKY9HBFlE6P+q
g+n8Da9FA46VjFunNxOp9eoE+mKkcYHdNP6tf1sffbalNJTbujDB8USnzkH58DMSZf1IsHq2pDfs
eRNZ4uWnvFCXI3jcdVr4GaY8DpSByjAm4Zfi3kwvEJbdNO2dBijKeQwDW9RtdkhufkwbXkgolBxW
KyutN6dpLyOUN/FSfHjRgrg1JMR2F0YVMtoFLqRnH+6EC21rsT8k9OO9rXsTysNVlVA/ifpodUL2
2mJ7AjGxEacHywrE2fhDD5GLUcu/A+4amhBa6FUf3QgpYCgvJPF1yoq6hP4WFyUEpXlXkJwZHRby
1YDFLNVRXYF2y+nwaOdQKTy3nCqH1AejirCUisPMTpn9SNCw9iLBVKSy6esQZIkjgRhhWuPMFSZm
MMOuy2y8zHHscG1/1PFxSfnaSjv+7dq7hkp+WQnqRmVimZGyODs16sIzgo9EA/EX+g7hvs0wVpFz
5MrKhuIfUDj+NxaH/3e3gyXyvRSqQyIV/QV9Hm3mr9No4Xn7/KqDFGIB9jSg+odLBj0vzWlJwd6h
UDHjAw2Rg0crKZMnsGMe99yz3WDUU9p0so7Q9iTycmQXp/WjhQhDuplozLhJ9lPwM1klrNbj9ZCm
rRBww+TRV2C0Y2KJry3J/mPoIO8Er/WuwLySrtr+AF/HhsnSfP2H6lmHca46lxfQhvY8mIx7q+FK
FVfh4xbe2hCuW/B0YM0ojSZmkMLTT0WSlZ4wCoHAzz7wFtwXIuyxZ7lXEYkJg59qUb48oLTZdAeh
+/1ap6WN3wtjur283v2h9cBlqybPH0HKu7SQqthLWC99q0oHwePMYL9uX7qhT2oakznakRRMCz5C
eQ7ZC3Wk9djl9eMJZzRdXm95g9DQJqucBBDO9FTr5aghW+G/sUnREcIINXOs2vLDNG48raReFzl3
NHdQuYd7nbbwdpmSf5MLyBgoOdc0ZSGncVIbck41FkwMz2nYxXMZA60RZNsUswVi/8fko7NUu6IQ
TWvEzvxXYJdmXBdhFr/Ba0wLHArCjtBRItymqMY39xuchi7zHOhwwix+mBMVa0qdI7o75BwWqK+l
c6VfyhFnN10g5JuJf0lJRPwz2m26kgEqrnPyLI3QtfJVJpHfl3G+seAB9eD+3rYi2zwS0hr1zPwV
F6JHzQoLVpzqqAhU3azuR9LnoTi5rfPekwTVPsGkl5DyItm/041qZ+Zr/xjDK9JNksbFqjeWeUlx
ndkGKZykS6zTsfhXIPTW9PqoshqK6GSVcADihbVwZJwuejgAlDo0JgQ++YuLvcHRMM6Ndl9Broxz
k84gaRg3ooqCrn0FviOEQylsZbn6IBkx5vcHepfE6N0BfLrBWM26Irto6LySXkpenDexGNUyf/b8
Tvux2s8pDDQDmxk476Ym2dDOLbOD9PvYniiploIhCM0S2LN9cZd2HpOMaCIIzRUGBWtZ+UCiKMZI
5cis7sAqpAKkqxHV19iNAIfBvKdVAcFTXFQ5O5GRd4CNBbYulLoxU570gHuuLOcO3gvSCWjxdawY
kUgQuiilF2Sta46tBEnTT2SC51w1iDupRIJw/D/PiRx3o/CdJAl65xfRqRagrdQoVy7U3Y7ckb//
6w5OWMURo+wstDhWiLTT8HYgTA8eOOhBkP3side/uYck+6K7s7HSSja8pygtPAl3k7C0PIs9VYeF
Ot9gGDfAD2ld505aNr7Y7Wyu0FdjIkdkCTwYgTPDYZ9IqB1S7BVcJ04+2zBLkJxAG3fV8oz3tdWp
rCUMs1EcMUKrOF3THpbOLjzYN18KDt295yXv4ws+XoKZHkmfxsOFF7fgmZr27R3U6clTEbL4GYUi
5oMDs87Xih8Fdtf0+7PC/cCG70e5FoY23QhD+UXqkXwKe9xPnCgGDh9QdQqNAsposghcLkzz5wSA
Y1VmrrByumQGJfFtYCT7+6PF14D9TLZeYREDYq7ejnd++5bWz4hiF644U3JF/bh/yMwgvQzUiNmk
HNyx879+egyPECv/DehYmNiPPo6bDefQ3xTZGmF2cdsi7h5KJZW4beKf1JucFMIpMzwxn1iAAzSk
yhx6ktfbJduuldGo3uh4Tu1S+Tgcp335lyOcE4yfGlgK1jNYUcSC9Z83haDQdqgU24/gYkUr/nhq
fRDaSaPenoZGEEh4xBBU98jYuWf5XnvMdLnfeSo9y2lBR5//5TaqhkbASBcBCn3jkQ64V3Omhk7d
Ym19N60busXETojfvC6Omp9WtM3h3emIX2w610MRGha1fn1lQjAeqXmDGckGGWVbYpTkljmOFwyX
qVKlsJiwT1SgKqlt7uYReJwPyNYAiw2sYGC93N174DWzDtFWG3bwM86WhjLJbzNYVcWTh2Qv1Gb0
gUmqinuZrU2glFEqg5owQHzZ+0/PqfWR0MHA03lz8MMNNsS2cNMgazJXdkINrcjlcak7cgM82J8C
M6c5w7dqCFquiTHrf3jAlzYH8TEKbbYs89j+A1YUBzanzylJqoeOwQQmk4rcGVqdAcVo9gyGv7Xb
Q7MQO1IhDMUPZxQowQ2VxipWNlwYVTdzA4WWpoFP13X1Y8/Uqx8M8y9UFW6+iHd/VslBVvF1KqS2
1drYK4oK7BEYfYXQ45iJ8oxgV4fqVfOGFZcEug6CBGAZ6KFsssxg+Y9D9RuietW6nOCqIQVZqN7f
cBt8TLV2jcIOspT4G7fqq9g/5Z5C5zMvLe6MYh3h8wzQO06A6g77Dd6N1ouf+OflBke6Pe3PEzPJ
UXsNZ8YVJ13c6AfFXeIoegLQjSUJac8+cjV7XpiJpb7NDaWOEWsi1MTmwoeP0Do9v65zdFkA5wu+
RyUqafKpn3KQTHInRT7mSJYTu9aqt8ikMYffcr2on8bWI4OH4z/AxC1lVnQoSkQOul5EP9VoLFDI
Yassnp5ZxtBcf4eGWuH2N55qWOpUPmJfJQ2zZiQg1VpEROKkQK/73moEw77fRRgUyO9NZWJ75T44
d3Pes3RqnQnZFzrwmWQ8HPQNU+c2+mqfsl2r5zKSQDOVHFDbAAMsXgsa0JKilNJz4obVNkD9d+IP
d5o1n3SN5mODuCo+YFHoB/Y12dJwiVvBV4WkAFwrxr93CMUbN8iA8VWuisoMK6Coh32QlAcpFB/s
sHYSRW+VdW70XxDXiF02IIQLGs84KT3/PhzHBBGXSZf694p3b/qGVP+njRK7FD+yLtGRQ6KBfOlC
50BLBt+FVN44xmeWqTYQuqjr1hwspmssv0ND8V2QbZcZ2rRJR8ChPk6RUatYVQJoDeSD5TV7b9Kq
TmHFVtrNw5WB8ycBmYlUtUssCwAi6zQsqnky+/rmM0TOrQXMsNYEaBldvvla0OJIxDSdZ43tJUba
An2ao14ss0jZ0qRHMrM5aHy9I0bv8R9Fb+743IqtWW+K+R+rGQtVFU2wDaUZgY5TFs5ZaGzoId+1
atcj4C58RcmRHkHot0Oic6dys/BMBgpjmBd9dFRVIxTmFuhMD0C06lkg3CMarXL6jp48Wc5pNRFd
YgiSs3FFQLJ3lAaHLAGtP6dzJtWAaSanqOYdZi/9K4PMXzI69u5D4IyP655VVwsg5AVMJoKLfFlC
XD/kINtue2Da4JCl8gXsJNy66k97zvn+WCVT926PPDOtm3bLjlE3WJmXG6iKYDNQPS2rcTsi3y48
irXDOw/8eBacJPnzc8GipGKfMlNeZ0KZGPFDwnrJ8U/c+6PttJ7tsGZfD/hhAVXapoZECeYgt6GK
UEN/srqEIDyVvPP52+UJeF8r+hmcZqez+vc5RTaPDWvXTLen1Vk/IekH/GdfZP3S7kWJ7dnfGt9e
sUNWQIANVicNZEClmewxBLrX6/7694+U6zU/rP6IYM7GWz3ceMH93y6rizjc5gSgQl7DGPOOhORG
OiduU1PzHCegZpCga+O5QGWToYYJp+GhaXSpqjWTq6HNgpZUVXR98I7h5owMepGpcoTBo2Rfj4cY
9OAI/ft8WipC7fmmsBpK6kIyoOHJlwv2CeanJhhTRsL3Ofp1K7JKv/cjmZXHGhAurIJfNcawuab+
hC0acUAZwSxH8aptv8JU+yAWhjTTNTxA7xIh2AEYSCLOe4ACGWEGTk/iAPM7fhmk21tfxhAzm+eI
tTDnrSyjnsneARptcbiBvKHMjg+ekFA2mLlqc2vcZzEp1M7TS0TLtFwBtRt8k8Jhud4B9ev1in3Y
GN3ZC/T9HOT/JClIoEErurVnxVq4GI9jumD2C/bgTIzsNTVOI9j/Wy9jN6GuQl9ZZKFjAdvo7GZV
yl/v5GHwNMnbEDl+MdxV0BXFGeGjpjo9rF0vnfh0bswb85P0K+Ps4QjuWAjr4ZPb3nIg1oqx2gz1
c4YeGAKE9qSfyrcn4iXw7ZYsTNu/a8zV1CjFHGUbER3FOBOBBa1hIappcavu53QLm/MLr0naMpll
EC/6XSvnVcABzdqDrxcTmZwNefDoiYbUNCd+4I5HklD5DO0lNFkBLp6M4SIN4oOpru8eZavrvwKe
pspm67i2MZoKB/G7ZmkQhywRfb138rD6QNX/AsVYyqQQ+wZdRZP0uxWLt469u0yhXDz0w3CEWSei
6T9gHSAGurzYaRo06LvEYhFGiSL+aLKD6zpHHZK4i2NpI15I+oc4sYBuQxCnbvmgMulpJoJttkBZ
AyCWtwDh+qo2yZNwI/6wq2TnDukHU5w5tlpVPIZmP+DzehDjapNRzmvKS1nD0lPDf1N2vBAfKyAE
/6LgcojVwmPG1Daen6Qe0atb0HAZBP2dvlT01HCj+1WJZdd1kSpb5m7CiuCNcZG404Tmj/XRO1zg
nIXJgJTtQ3KT0QH7iP5ohAKeQajx9IW4NFm6O+3KndPZr3VNcX33rvhxWUGhBsxK2K5fX+Bjbr29
2+HqSCsTAXs5Ahekn+w0OGnXdL0/piN0pB0wNlRTEU6/HC04JiU50Rt6RoY60HoPzG6YMqJFuQFH
QtBSME3WlkR+Q08gpP988QT9GNo1PT91pIIX03EUgjEhwcYe9MxYc0mVMwWQOLj69TyuWQwIBzRS
vX7dpW2QewuheOpAOx2QsVsR4aUlQdgeu43Nz/lJKuT8WBrT+7/c/5bqrJ0oTMK7odHLEV9DmcS4
HIp69HQrbWsOIJdnQCCW3A+iNWZfhoeMUIknyXB0imKj2RJUUU7BVH8O3XaLOU/bXnQ4q2I/+44k
HGnFET/AaKW2i9lXJrzH9FHsHYHORFqqnNiHyUHuF4aYsTlV+vDAITz0fvWskMAkHnsASRr5uCjG
iasl1fY4oo1FmceqgMeLKgTGR8YtUnwoYeCW8+j/ZS5bda32lip7Cc0+ShLfU42Hu4zNw5mj/lJF
xWSBVl9hYyoYucbr6Sg5/3gfs1EgfoRtg5vACJBp+CDRm+nmTDqK91dUKypHsT6wOxCNb2gez3yd
kmrpzr3hpa68IABZfg6xVQbTRHy5jnNxl0Qxq6vn5cevo/PP5kTw+QzWnU6RAEnZMXuVpkYJQOVm
5hvwLbDPC5sUcr6hjTUMgL0UHFiNFCoYgO12Rv0s/mw7TL9qGS8tjMdkb6p+PZzkbPFVV/ejiWg0
0U3O2lcx8ZOuGxWlSraKI/Em1ga1nKvlmF+vQAde0ndlNOM7eJ7F43XsECOpPtdUR26BMkx+dPk6
Bi37gvADzUB9O6Fi3yUvnZJv0mrpjSPRHsJGyeSXGe6SydREk07OXMWup0N3NRjLjShvl08ECfTz
9shzkpXXoc5sIWZrwiZpsY8yKVwxJOBe7eFUPGuzf7rS4c1ZEjYFlVjA6IPwarG9UEyqQHZ/v04B
Eq3xG2P4CRLWahxM0Xb+ozTPYUgxMIzVG8GjZBazrUZ6agnHGWxute8+l7xZuL8+g4aL77WzlS8c
BBqohxogusR724yZoO6IsKW7+FkEiEScYMPMQaP8xdduNR5nOOtWkNEGuZe0m7CQ6gv/G0XILNfD
HLH0RFXUZbMvu8Pq1X4X8MbqyOI1LctVTVdxlCxF+8cq+LEUFzmVes+bgFcUzGqvghtjT5BbO0Fo
HbWqgO5GLFHfwTbr6hcAQUIgpx5MKZqKSYdp1Pf5sO3hcv4nt4XxZa3MUB9/spbuBlzYOq+ePPBB
cwOWO9KtLv3EWkMRxAbD8qVTRxPtEImRLxNqi5p5OVxT7tjSlYXmF5h66C5Ot6Jt3TFqEUkMd8kp
Y6/r3Y6s401swHZVKcydIsS41iSAUBPK/YEpDYJ4Bu5/AuR7/KpJ8D9QsPcuYOlRgGJSKyga4qzU
RzmWfsUZF1htWn0U76BAF0CiN25wBBgSzjBAR4pIEy8ydDGTwKHyaZfczUEDSZShwY33TlOBjk0A
XsHrNfP2GVpzEIJUp8dra4DbHTolPsMJwIgrMRD2cZB5m5+mHX9Bo23TtHynvvAtWcX3NNs3KyX3
K6drfgc21OqNUjj7MDRozqpMehDujrsjDZ7xP/Z1Bx5DKLEPaa2hwmVoSrRgqvndEogkmuUJf2Dj
39kKYr+tTt0lvVWy4wEllOUZKtytaQ6/JM38u44MpViPrZI/10/5z4DmARMP5gZy2EuQTu99nhSt
Th8wBGX7dfA9vcy2mWiXBMQPS4TGxYWhG8BFoLZK6z7zBcXs6XZvaYlE1ZHRs5Shblf3jxEQ2VeG
UtbpeBPvyIcDy0XFZaz5qJXDz5612y/j90XJIAF3tIdFGUpcP2YVCT3E4bzp/E2zN1Z90+zZe7/b
3svIlS13o9JeQrpMaOWwsiw2CMqIIZH7iMqhR29ZrzZ89tI6SGg/szJ+b7z9x+meJdH/jmU+guue
bRDPGeZ/JIt/UgCO4ST/wL4sJqo+0mCsgzvT9mW2Y3ILDOi645eGSXRY9pNEare0KcLXkRIDjzJV
SYOaS6SAr5m6fm8rTnc8YPHPeUlxb8mJgC5Mk9EvIed82zvo7Sepd2eJT9PfU5S1u1C3okFGXeua
/oiTq1pjwaGXHZH61/T28c/0AWTXHiiDWExZeV24XDKL/1RYFW4ogclm9qJed24a0TT//lTEANTO
byIiFrSSaSMx9qO0PBtxcIWddXaTHRsldSP8oX1ohbV1HxyRyRtHiaq7ak1GCPwKvFoSqQhvk04U
tZjGysqpVw+R5Ww9avzIvbj9Xic5vQcC/bU57hGYZ6YFiHSvrwPGycxjVey4+hDo3usoDAq4lGP7
SEq8Nqi1A9pmPpQxbmV1XpFKDMoqzSxL+qWdd4q57wCMFbpgq2cwQwG4R4P8Ty/a2t2cdsB/DG5Z
jA0V7e1pbQwdLLBRgUGWX3TRxTvNW3b/zavaFdWZnQrFr3EnoZOLuRxQYPBza66VjEDTa5dmn04r
aNNwB3Z4vi3wqyXHrcbIAQv3cb1UwnnWIWfaezWpYTRqEhVjioBVYv5v/tTCbARuBsCP5LGU9mO2
QBca0sQCUVsxSn+h+0P4vXwDn2OUgJR8hQ93x8AZYdPAvK+trbjtKf/VpN7rkc7BvQoRBzXHMtVw
gk6sQvtxJj4GbDiHvCRH5oZQ971pZvuHOiFzM6CZIAGBd1yPP9t0/qhVT/G02NUF1vRB0VdgL5dl
3exIWn6BMtLl9Fao15/Ybpocfvznp7424fh+8A1g6yL7ycefFqRjDUrelFGdrWnuxqUAhZsnpEVL
ECDVYuzctSmCtZI+BKi3UkBFvA3j/5L4MBSOdxMEdnWtcgkdxmNjrOtncrCmqjGCaRql9fAsUVKg
0ReJFdrlPpgrikF6O+EwwxkrEN43zgqXwDdWyV08Ain5kpF9+7Feb9pqRbognqgHRcT0Gds4hPnH
hjCLTcdY1fvXmYyiiGsBRqIHZy3z4LTD97DpdCK9yR9RjyDc50T4s6COInASZMBxb+f10WCCtO88
wwCD7SuuqPrSx5bQOKMrHFQ3KNYp7vPbaVw5ds197Ahz77GwKpHg57c3DyIXdDzxbhifT9CI1Wg3
Ip3GyoFpAAuz7u0X+Q7WpH300/p09eEpUYO7+BeBV0JL7KFOmAh9FnBtkcbrcCXAnVCIOO2lG5QQ
V6tdtV73nCxHIdfikf7UNa3LwcQtqcyJz+TLQ44VAGwuHU1xY7jDcm87IMqt8mXL9ANl75ZChTEz
uaxGuLS6nNu09BfhQYiuXTGS0eVLkSyQUq3VuiQ2uWqKHX1Xso1MRhctSZlCbgUqqykEENhe5DCj
0WHWnpaTO7dEJL74YizUH6HW5wMagusUN7LiVLEbTy1Y41JbTAZMCfak59IStoR030/z735inoXx
MWvfa9MgWyJAzvsQSBPDBgZvP4cEgTzd+A5XRYOcQMEbhvJGJwtLnSJqFiYSvTrrg8YGAsocm+x8
ANnB5RO2l/wrI8OjtnSwqkPGKKDVZtwa26Jj9XYd0XKRHScDt2PoGmNHSwnEIoa0f7VPAPx0OHdr
Agu6xDSBzOnL/1hLlIc17MtDncEjva131AfJJX3RP8L6rK2H+7toIAFy7eGlkHVnbtJ+WJ6U+pjg
dXbvtV+OXlke4RciyiIJ9N3mAYDEhXoA2XcJ2UVPrbcUmDOWEU/H/o09JJtJ81Mn43GzwBgGqGGz
KRVs6deCo0nzqDJfx1muLnSOGMAgZQ7LwaC6pHVjSg917p2/GNzfa/TTNPhbV1oDtYgyP6HTxjLj
4vDHzqyrBgzM8fio1fXjRuMDPqJ8acsZJedXVv+yYjkob9ljTZ2O8oVl+ITDzDpUYPpRoASuc/kT
KmGKt2MwPxeS4JYvxfQwggxnNo0QBtpc9is5oZZW2JVjTk6gDMYL8ZANN6VRqbAFdFpSP823Zbb2
Akx38RMQF6g1WGKsjU8Dw8dq0DU8G70zsuuxKNKp4NTsmJQ3oHz5UO7CtXV3Vlod/dPATkLP8ST+
b7345R3U9+t/eaoLscXUt3KPyWkG+e7FHJ0R6G+PSLh4MQZNk+VCit4GRl1ZLgW5hY6VQxJp9g79
95m+hU/tUySxJZGoPQ8LrkqqSH+EcgyXps4u8jjGEirKBkHk6EZ95fgJY6qONXjts+e7pDYj1pju
2nOwXSoCx7FD1loPE0ZXkjJn4GIzUnqXc+MsZ1FEqqG3yngJpOgzTwUam/Vyn9JzYGPn89JTMp+O
qY9ZEEW5tGPFlIwYuDASsqh4BXFkso0XfKeSmDhP7kzL1XbbALIg/RsB8r1OYiD7sM4S9mVKA/BE
LiCdbvTI7Rebg82iSwQ8grcJ+2YL6GYlU1ZfToLhOm1GAHs3LUB6Dr+Tw5nIMfMKliLaZzOm9F49
Mz3OIFS6hgUilAbL17VQD7OziWdyAbHqBbwZnQm1KTdWC6L0/Kr3Hg+3moJTo4OzY+DNw318kcnj
+vTqiOokHsFuJq6TNE2FWvR+D3pKC5ue4dgP8tPUeCvxmsNxzz6w5uuE0IkLR81wfVMsDJEgt1/i
5BQrUxeCjapTVhftFtRszZH2ABgSA67+gaqX0w8W2BpK32u+76MHClBUojVDgwKATdqZBSY86MOB
dHn1PCLtfs+M6AWXVOjYAMxtL1r+B+oEH6ytwm0vt5+ANlWMx6SPrRvRZ8w7FOkbbeq0X+1DPN44
VzqmnIsrcaI8I8d2/Pp1aZHcV00jYJZ7fRYw9dghYhn+k7vS0j37LPZHGOkEnuXGrH6PkDLwtYLf
JzunuydY5bSSN6KTAX1qxyNm3QWE8xVJmu87+JBJzFb/JcKakEymL7eGXorHZo1L6PwR5jk/o5Qr
qgNoy66o9BvxDouqA7bzC5KDRyCPsABX7yFtSvojbkCatdRn6E64Pp14xRNLD7B1wkRvPxDFZR//
gUANve3jKIjbEV/6bwzX0U1+9jphRdx7UrOfC1v8oN3xtJtwK79zMUnx+MkQo2RsTgLgpLahGnBf
MciwKKGjJ/IzuGGJ8KBx57AbVMUNMagY58RnwTPmV9lXSCMhe9zTr3ywjwZ2hJHGqxhX+1WY/9HS
B+5hkEvNmFDjt9qhgUgAtVWzTf3rveP+us3QVsqnzhfl1Q2/hAakAlQaobxm0eHGryfngDXt8hlH
2tkodqqOwcjV7flTCC+aNGdAstL/JKbiDlr5ATxD0048iRY0Isf3s4kuJ7n8RCpC7JVfCgYmRW1Q
D73taNcsRhg5p3N9n8/yOvvpkeLW199dpyqo+TfMejUATSporvuHKUjfbFDfZy7U6IdIMF1L0GOD
N4tCjyAab9a//2ZbolIQwdVOLMzjoW/m6vhqmbU2nOUmYjbyNz77hgyZK8NGIPuicSRaMP5EYIOa
GK7Dj94A/yTIqckgsAz+oZFroPZmC/cB8FdKBpKrvfkmJ4CIPnnKJOq5JA+L97vO7942vCNouOKQ
+tJhdSF4qLbonLkYE3CSlpYFtBw1rfVraie1lmUKmemfw8IEDOpfXz2EiL+M0Rol3UIrVTpVMCKt
b3M1b7sRyvA9vf7/Ou6Qgy+WfMTP0ACXeFukCVAnrR6SycVQvTDDFCW73J+tsSq6GFfK/IMQh+ai
/3BBctmzScjTHYfJmv0NxLgGV7+OdnPzpSQcWZTM8G0+FkSFIRUFXYnVIB6Mq5vVMHY4Zde8EkH6
Y2pra1PJ5OC1c4zukB4CFH+EOcoOFJ8kE1TF0Z3WdjPvcOUA9eGenhX3F/msuIBXwn9IMfg+Dei8
2JI+vcojUU9d/XhRLGsCdh6k/c0lVv7paw1njX9C5XgO0L52Dt/wjJh0mC1Omw14sBhh4ybA041c
Rw9aslwb8s+pxg6kuvh27DNPGMucnfTweNFS2pdxNA30HttIBcpwAx7A9k3hibYlF4MS60jqJSHR
8241wvUe8GfsUmMyAcYbl3ccATdQ0cu1VFEFTFNfPlg3Nmz7NMnVkhGIzKO9ukUmeOLB4E5G8Sqh
MvVa7FacEJh8vl0aKVM74j2EKZMQkngFJtNGFyr4xEaehdSIHJtJA2yJglNvbUOsD5UceKKxVBeU
GW9Fb8wuL5UV4wKKir01k8c+8dT5XR/3Wig+i2BFFcmcN1aSeuGD3i6cY2gwMowx0cpyTutlAzpi
sGghUY2J0phAisFo/uGU8FwqV7n1iMEnfXBJNONvyEiC+tS+DVMWgVjeXALigsSlk+w764YaLxP5
O58dSvupexaC6Ok9OLZ05EfcfFIoYtykyqcBxcdNbxj3iheHCX/yR2B2M8Yd2cClXZaXsprLbN6E
P4RzoLxf8JeyrLIb80WBk3fF1CbbZRJb7wENjRNnb6pvX/P94oPUYi2ZG1mlfmSDEC7Z6fBjzb4T
/81mWnB9jm4XqDc+d1XvGSMnBfPIrcUmi3Bg5l2Q9vz83HdsFnFHLFU2TtCiclizf1SZ4/XLpVco
4+IDthH0udDrttti6c8C/TEenlXz4B1wXhPlNwXqMf15+/J7gFOBVCTYsYDtElrydJfnvgYy3Zzs
3f9dwsIE8aeOg4FPFBC9djkKHdvziOaG+a8yeOwCQrTfKa6+2/FvA6RVLn/v3CVI5Kjmr6NSiv1/
+5gSkBHDonpvWlRpulFuwEsSP+IYUN1TB7kFstutAnQn1H2Wm+FZnHK2YeM7RjGuogvKX0Q+wFin
tHl4tvEoxUMJViESzLnOzM58xJqamn5YcjhbwwQ8Z6IoT5W8wVBrGkipY/sp8wuLeptcVEjg+G01
k6ozBh6gk/Qk/rBiZ8xoZilrVeiTW639Atgelz7rCHla9xsE158YT+l+aeSr6HuQk+LYKyEb5ka4
9Liw4iUqqzAlAqrVxqPU+B/jqwvvoVJd2CaXPBgOYa9fW1CC836J+FxZwZZlbhLXl+lcb1Yy9JD9
58kYhikYbWTIF4cvhd8yoC/c4gzCScnc6oJlQr7qZ0Qc0LxAyVlqp2JfgkCReoZmE64+wXSZ6+BF
7WgeuTS7BZOOCKw5oXbScGYFhi7ZiZ8X0w2D4PxAvb1ytrUsbGgRzYJeLkxFHNZjBzjV940HHn2K
mrPrBupTh+ovgxt35gw3WIxRtW5rvOO9sU9wXwUs4TCRxIHNNTGBdO1FYwSXZ1WszCRRKjVkJSHI
JbIVy8MnV6JJKecbOJRXK7HfGViWjvaUiIZtbbwkK207/G/FQe16sf0Pd1NOxvst91YqVzoiU3G2
KwmjF0D7lnpFurMgf7ONBbGAEkuy3bwsORvb6MAYO8iWMzB3BhoWme5rdcmifyHp61cX64yXJJ9h
BffdPpQLmCvBeD8zj+t+jncE3Ea5LTlggCeCOkklAbCGdgRPnhMRIaH4a+zlaN8wJsRI2/vAq2w7
x/KfwY0WX8uI6L7rmGIdCwIc2Mu5Gj76v07HntL1NOKEpDCXiqW0Z4RMw6VMenah6qq4Sr/3YWNh
wf+VFsP9t3zJqnp1Y1ZBOdwmJ/GMtb5yUpRLghi0mtNsgVQT06yVsc1utx5NcgS+0ary/VKGnQnQ
Q/TRipd14ntQHWlaQUVMmazfJrc5JdoNpab1nlR4LhdfRCe5FX68QjNKozHBk2awoJmFYw4cd2IP
iEP6czLuGEywkNN7UY/2dsgdYC3rbfXg9j++RBdTtb62Pj0lLqle1NvApS7ag0uBoboDRnvCxHai
e5WrDReMfHVQe72nobHbQNYhnzO1owhG3Jm2l4kE/+XCdkDcMORdCqDNnBcJnRp0Gnwn9oPcFrdb
0AH2h3J/zm2MMGI0R/1ZR6N5YiyPaPujmBMcOfDp3ohcEJDj37raKbuW1uSpUvbIoVAaiFYxmZLw
K2ID24RDB/BmKlBuemjaZ1mE4XCEr6MNAUMjTuEc+D9cAylZbxZ8W33/44sZ+L8SDjRR8lPx8Qb0
GmuTgDs4QVeiqNL8m5VHOEpw7c20DgI14BeNY74Je7ka80GeY6Zzd4Kl2z906C3aMVF8u+muhr37
7sTTwHSoNrkwk/2QEHKnItlWQYTlwgMrLC5sKjbtcbN36zlErjflpz0LDWJwcw22j/Gmy6veIAJ3
hh6Z3+XOZ/Z27lOxJox0JIzouaBEsrj0ho5oKllboQhHsQSYBqfdZfr+z+PJnD0X6evSXP0cnT/O
i6W0VIKwbwk8F3aacoZzm2983mA5jK76mRl/g7ecTSpt+r6V75qFNnziUtZyhtlcAQB4+O9L9CAE
E7ui1+ZK8SL4WXr6gpyTWM6ky/5AyO0TX5ymi6eVFLtm+kIf0ejXnO6YkHA0BUm6xumdZ7bw5rdZ
6u90mP3jBTPTKaN0Vcl/y1Bf0paTwBAZvdySjH6P59VlwVnCr3zBXSLh6C4eI2Lf56rFIBqMs+Sh
YgibZwNhUywaV9BPCr1WoScU/Qahu0TRbze/fO5hGDn6LJqs53XNG6tEd+KHEybt3s0vnywN3ipI
mCZ5cAO1+SBU067Cc5LNQjfDChEUa2MvtvrS7S5lfPELuorOF+ijtygNY3hxi2T/ypxqIxzHeJlR
08ajDVg5y6StENMNLNmIYZ64cxqyaV+PlERV5cSi8NfyzJgdryvtoiX0vvz3I9KJIU5TM02D+S3g
x5RiHasY9QFK10+Bh87yggZF+MvMqwPKbkLKOXa6tOm9CL/vxEk9quePT+Vv8M0rrAlG0ZM47CbX
TY6gffSYXbCL5IBKkR6AFL+bLHx2jRcKUyKJzdIGMm4qAhDD9ToQvlfZk6jM5rU6Pu4g2nBdITxx
pUB6skedoDByt4SbWgmC9t5NFRFDR4OHg7i2W63NxgZIl6zj7C1zuThjEKYTYGtSa3RD3LhePqgu
nCvY9CkUZvUK/bR3rGvwJ0RW56n+QLpudI5PEUYkItuk7fKi84Yg2AIIivBX7MsCqFBS5+G0slrZ
iB/EIQZxWYPLx8HnC7+h1b82/GW9biS045eBhpd/yzV0pj8ayawOWNtLy45bMPYsPxcOxueX0dJo
GNTfTPntALMTcamr8xHTbmykw2+2g8BgljWuY3U0uAOgxHhiaev2CO/jFf5BcFqYNYkeITO04WEM
JxXkn1LHXoDokcXed+gAQeONKrteRurDMTdHHpRUDb5PZQ+6g4KrddetSu6JDb3Mlgr/QriKnVsN
KVDnyIt7Bi5IfCjZShFsUXSDGo9h//eSmQJXUcu6gOycM6IgDWc977Q35mjWAckq8CsSdsHjm1vb
Lr9EkXtDCbffb0eoW8TKHo7IUJJpnvQHloJbCQ09pK3dkge+kJNefAjaJv/EUyznhhTPsrvt5PrR
5gJUB6+DdLfM3hdEfOigbwHds20BcOKN0Mb/BHb1wuXiIkmpIWYftQgEm/UisAXEFs6NCD26ggVC
5VOlN8Er8tmtolTyMjP25ezbbs8O5xXfaTsLfAYyYJEVGpOR0zo7xcD3Jg6hij55Wxm2ynKnFLOs
x6aRBH0TFUrRIC7eiZ/CzjYGPvOSFJs7xmZvweb2XiyY64XWhxu5X7RBqCjnsKT+dEairfr5s97J
3nHt1rTdV8vLOWRVDtgirNZJ3hwUDz0KgIyaNI6Sy8oFBVDlnB56hQoGxPfF439I6nLR2wp6klqc
uuLzs+PxsS13iT/acbbK1p3H6CIAeg3H6sR4o6betRV1n/n0Sc/TlZwFidS937kflhPKrKmBqizN
4sATIQdkANcVBE1heMW2Q3lsNUv8Plfp3Qgj3UqGUlop7r7QPMIEkWBm4KHEJ/xVoys24N7+Cydu
DxpnyJ5rdzPLj+wxzdFZi7QNBNddmLXyvtscZ07e4T8ze1HnZF7pSadOrsVjMR74cnLDVZnxCK5l
pNpWH7736B4d7ggtoDCcndEeGEFKkZUQtnpEwzJDhdGO7TKTGe6fzAnAangD3Q7C11GXrwCs/25H
C/zCV5AC/gzKRtDeV9iCLQSdNynNWVHNPX8TjbRnKpfLMygTLKesNtefx2TSlPm7xNWJ2GtbqEgx
RsjOtr80CBnAtzfVr5GxSCmUhhZ4d24EHQBi+B0H7/fsSIh/luNfnjRz7N8hkyVtNFYzSw9jIHhk
NpgBe6KQ8YVGXkSJP34S1ivsL7z2cN2vduvu2yIrhWCgmMwhquwZ8VcfXPl+TeH3oz4mpFoOHUo5
nxk1zCR0jmw1cs1rRueGBAkXp3tF/ofUVHxoLAu5MdkgcVBvHWRHFBUQ76A+eMdEaIEYTCds0cep
sd3gAmTazsQWHY3sDmXxqLML9vDBz+0hh0pZfiv7kKnXdN5/7G8TL9lLvxKWtMhSapBuXWI9Gaaq
iYAr3cosiT58x/1WauEz43GEKvgqiViQtxqovhk/WcbQ3UxxsTMCvU4U8npNazrP5bbPckXhVmo6
SomOzFNgeK94aApjDooneQDVM8U3Ui3ji+tOgDUBu797C2IqGEhslXXPCdyrJ3aisQH1ESLR1tR1
H5asTlW3yskMwdjoyUyOgMxOzMZdAWSOABSix4HL849apdjSr76WnTnzgXW/EwsqoaqhW2m3cVK8
QpUr+x5IBr5tn57VTyWKmiMuUV4I8xTQPSimwZ6Kyhsqs2RSDFwJies0tzw2CQ2eErJ6qXriB30w
XkuiKwsZhl65XnUJRpJQPSJKHx09aEtvgo7tRB8xf7djDishMLSIEeKX6FhMdph5BPGgmQZJiQ3C
yTH/MamReXrQ5dzJS0UhQfXzJrn51wA+YfCkpJxArxY+CjYVaVJDAWF0Se8P1HcV3f4kt1j88+E3
8glyxxAqZ5myhLlkOFEiDeCUevDR1EdACG0EmqaQBcYw2sWnPzmE4yiB3FKiNDa6KAYNZUmM0ITk
8SOqnVMFVYNLZvG50AfCB1lC7nGVhqU9Lebx5JIOL+Nmxu7kAh0/8wnrJhDh7ZBFkKqWMHrGeC1u
i4fCPkoz9lJjS39GAYRBIS7nRh0iAFKgmnr+spD40RTPHvlyfPSqX5WnBNI4tutU2ba2pq1XCUEL
744ViTWMCDlpHCyzdUOCeXLkWwiJnOSsb/wE7ayX4Gs1kl10dXQVWEPac+LJiZTf62ZAdOINKQcD
YYjPtq1+U33gVyxBQY//sjolHusEDodFQ629lRmGEiuaNGe+4p0idl52vWiLokWDek7vc88lLUqk
azPZjhK/b5Dh99k0KvT6VKo1pI78K981QZUVMkz0s05ov53fY4h4+YP9AUdpnJe+fC/H7vrXWtBj
AwF/azx0gbvyld+U+x8E4bQLPCkbK3SvADUtB4DLq2P4I94+bc10cHYNzFQUe5EGFvedt4SSAa/a
wRGOBlSbH1p/pyU/1LcM0tL0f2UHhcXru7JEgCaV00l0Sg6DdqfxpusTJBwUAx9e67fwMZzfBFms
04dCu2oDctk9jT3P2qDJGfece+G1clsmNvNfUXvi+gR7JlY1gFk0wwa51vcL4nGqvVkmP0sZF458
BDmjO469WkrDVV1f6f51XkcCcXkOLKYbsJt87fsTkrDj83HLBxvngDLPEg9hXY72Vxzj+j8J5JCv
gtlRbeLgp3gb7is0/of9sEboY8invhEVOQPJBDn5t9bRGeXmeMabVIYe0Lz8VllFyoR9Iop+FzvM
kqFIJxgw1grikoBL4Rs211GQHLucYLJLajy6sM2XYG4NpNjcsOniBWggNKsWI+hVRwxRQZqQE65f
3Zy/+Wn4GH23Vc/rxNcytybr/06YeRLaZ2NvmMApUpv0kJul/eSFLdEB0ptNWynwwqZ7u6UU8Ebg
NyfZ6GPHRPISgTOeVC1sd+WB8zr6caSw794P5buGqrEe8JV/wEIeOdt4qbIGPNuT/xmfyqv7Sn+G
b4LsU9ZeWPGPe7cwM8yil35Zbk/H2h/yDeYsBicv04zZbL7eh+zLkYMCaK4Y4dn0vzaX3b5Nm4Iw
7aeJKTDoxs4lnD0NTdgbmnbLyA49rYdpcgcEFdFAaLvt9GlE8f+s40o6xpZ14MkN7NnIJ+Us0hef
JmgwYpd1tM9VqaEvTUi0VyLINDhsMWdEgWWIn7iasULqBKHsuRiJU7k5EVLD1PZLH+DIzB2kKrtI
Vn2VWXEmcvOa6jdEoQ2oYmDYTE/FeC1LBi68R7aTEkcobjVGPbxa6tZhCi1S9gBq45YFdYoovmXQ
YIT3+hQCWqX7bNUV5k+dQHvGIdsYtPG7QxPsYCnG7CeLXw4kvoXR95y8VWwwb9LiwEgD2BnPMN9T
7RhdeSwhOYhuZ9Ua7YmwBSBi2YfsamJnLo2A0heQFOJ7vjrDp3cjV6XazAA7n4XFZFgleS8Y7dAj
62kGBPlqaaqJLxAjIsx8+ZKgaaOhcnrCbjM3lAET5/2UCCqobPZtT7TeGqA/uTOAmrqOP4HuZbAl
7ChtmJOSHeogfSVmmGhrRMxFQHPDSHDNuNEkoHTRRoF+zuMCH8qPADVX3QDk76NPQt8t4T/335Rx
zkYM6HJCuYQQguIztLzXAXdJStnRefW+P5KFJVaX1jZSEIYlAeAMTymZBVPjfGVlPhlkzFAEhbTv
G7laFQRstbdU8Ri3qq+Tx8FCPRs5+rndBUp1eOPXUiOOiwWCYU+o4GNqFuooVa8RnmHd8P019loW
HOX2fQ6H/GK0B611sDdlis8vH0W8Z3+Y9KQZBnmTkVVcEUjxC3BujyYvi5ZjRYGPoprJA960l+92
i4GXtpbqGvkP5arTQtAmUQG69dXrPni/G29pinTaysDAOqX3PK6nsWGVmg/JR/n3Fnjj5horRV3c
f8dTg3Hji6JiejlzZuvyICCKY9Bxa6XdaP65VtozBD0TU2bV2sPZunXboilWBmhslNbTOlFL2sSD
T4u/0+ISUWK/yksuPDOai8yelCcgUwG+p7omUL+/RbDL0UsKN44HafZR7R78Ibu1dnLwuBxKGluU
rmpEqOHRDiUrIqKeWrVkNWPmaFdygOLKCE//ctOS4F8Xhl1K7JHIQKJNDz+l5zIINvcwkUv+ReVY
DWp0mcE8sgaurlCvlCeWU407e02H+FTRnhsRIxndfizanM4gvi7EOFG7C5HOTqU8yRIZ58NYN4zR
q4VufK24hg4844X3kuRVHSY690vEFCVy/8n5S402fWzeVPPjEe/8a55XNMISxgRArisZlH6NX3Uv
QD66IHjmngU57f5uvj/51Kob6Guoc3um3nUe1tUlp1bw9LuaY6xWAGfafvTICJRMc4uq1gpvC9/t
m9YRAdx2drYmBQ1QOkgic5yA+aV9vC97ryEVqrChkl8t/XqzWx4gVtyROLcQBepZyB6pvXvqhtDZ
l2BGjT3dKKFTfPdSu4sQ7GTrC+7gS7vlFg4ZfL3U4emEaoqEhY3ngXLn2jhHiBWbKt9FmTUb9Jiz
5EQKLfxznwAIHza4tQL3s85nnbdPHuxldkgDwMn15aEJttb/CTjOZzU35NJDgRhzUjZZsey8GhnD
n44WUjpFC3k4QH+MPJ2BeF79Y+7fZ0t3oyRpdI/YWSsgj4MC/BOUE21WwFDKo/dXQ0v3jeL36Vbe
h+xiQDpb78HkyGat51oDjEW6v7oerMcerrqflNd+M/REiH/YByldectPKT6pC7VFqxWK9/L7Fjun
79KUiGDtggpG4TzoACgekdWcKRCz4YdZP33uldp4UmGq38Os2ABa7y4zGuKU+5jaJmydpwFY7NmO
UArAa4d1yWd2W0VzGbpZEge3SR9GqEAn9rlZ22ITgTP2Y9HxSRtMh5X0fZ1erSAKPU110+s2t/SS
R8XBs0ux98f8U1BRNkmq97GqOUaT3cJCv7jEy11MjDrWG4lq46mOFmfg6NlpWGeKXuTUW0Z43MZ8
XK/vW127jy8KiXGr+RP9vdpeQeeJsqKhanIYKmS8p3RTcS5knIol7OB5iXUf02nQkZ1yfFMZu8R3
feiZAsosTQ9wRZUuMsY/TvxfcBBY6AaabJC8uX9H7Rl1GQ0MLHWPfvfqXdvPBDbfjBovaSUDxRiF
XinPo0cNmzJntNb0sJU2ox0SoHTSsRxaIdXnjnF6rfwW+iTNeW143xi83SZW+62+1niNmtYZ0wGP
S9vMmvfjh27TZSJSttxuDtTPrAS9H6nP0O12HskBeWa/vVuzsjiythTCI4cTQBpjBdp4BdCAvJVY
Abz12zMlI2ANdpoKZCry2ZoSawwp+th2MKebtFoaDGASZOyDUdBm7sOgH94Yh8ljTjD6wiNr97zZ
d30SCC1yKpf12CHtUQ3r0P0aL2s/yhBSZOpgArURIyMb70OvJTVft8mgG3DAy0sZbFvPT/wwVK4o
QFzJDeB2OrIsx3aeCvC07viwfseK1f1zDJpUKjK0APq/YUATJVEknywviveTvLdjnu0ezQZEkGH6
Yu5E5imBQC1mTindJdjDDLqmzCF3qPC4c5o5hNapiCLD6v0EKNGJFusg8PPLrpw5givnes8WsvLc
eBhDCQsPuB5f6oPy3kQBLQx3qLQD78ub3/qCF6a1f895AVL3/ro6hF77Un4O1TrTRmjl9jnYEay0
lK5RYGJoNzk/3WZJA4/VZMTmc5IFjcvk8m4UGJcIuzfni02SLJSfH9+PQQVCdAemF5dOSnqWub0f
1URV8DXCCiDk2U3JwDhMbUPjzD6JXygQjX1wZU2GGKp0KY2m9TbpXqCJ0vJTuyQPRhperuKV/hVt
8bFlNwZ98DDU8GDy+jQtg6lBt13I2Ny0Y49sw3MlCpaoTOUoRT8RPr++D5P0JUpx2EtuWJA2h7YK
SNI/LjJezROxvjvkQz+xAiLFp+7VqNNXvmJTSgBlwkrYjsg+e4v620rSQ3MYe4xeNzZ+gPcAhAC3
LXXD8mqDHtxw7lqCN61xX13kFwURV8LneUcDufKjxxUKh0XkzBklkjZCPGjzxQLUgSgOBnlpJZpU
uPS/WnhLxyW1axSlp0G8Y//L1TxXkWouvwMRmp8YLaoTbpHJJUrEjPJ8hDjOrxxTL9GAPIAYxstN
lRs0+C9LsvFkjauIr+amss1XwGE5HG9ln1S18powhmtZzP32C4HbAQKxvMbpYEefTknrAEQ15R8A
kDztCADdtfubD9s/BNOesORnye+l1ZxpOjawaeO3pHHzg0bJTD80GbRr75O3T0GJ1kpmoC8vSHuq
I46gfzPWR3Bo+vvz4E++FmMhJlQTMtNOwQPryTn0GYluG2GwYrZil8US0kiBecCdkN1JAGIJC82x
MKwCM6GqyVM11E6K75wwX4qZc3VwVEWtokJNoWUW79SvS8sPGbY0Lqw3d8AcwrextDFdiIz694j+
qc4Ap+eBPUbR9fpgYWuz4HGDcNU+8zmq2TZ87/GfULaZ4T49OsQ6PIFAF6zAckrcevvKgRQR/Ix9
lolGDmYwsTC4T5qGfRvgiQHVuN78l6ppi3BXU/JAbQK9osOpfe/tAZD1AEeFK/jlJUijUTE5+q4v
gCfMnvS8f5E4Oq1kBxcKss6VgoSmc7SG7N+F8h8yX480qVSZncw0KHLMOkE3ChBDprip443Z1GtP
84k6XKFkGU0V3eWqbLKJ1SbkchGevj8OLgMyl5f0Kq/PnfAyayK5f2q5krbmoaOd1+mZ/GKFOD25
9GTMGgqarSvfQsvIlrQx2It9SAAL1MRTCCueaOPFqe3F40IxgvMHNDTfP72v63Yxfi1w0bJ5WWoS
J83fzNT3LWUs0PDxMWwvzso75/QivOr/4BtFJCdZfvOTqPqwEMljAkvG5QFiyJm/rQaAKpmLF7jc
Zj31/vHI8QgCxflrzz24dMs/Mpgp4nT3ldyM3dSBBwULLfoaZgnajP8zgiLHwxM0tsqVbBG0gr+T
Uzu8eWkPt422dQdxO+AKj+2rea11UbBEb8o/Z28V8B2tyxpnvWfGMdqUyXxLLK/yt7Z/zflFNw68
SkzmDXnGADrOJUDULKbZ8OFe9Ot/Ojk8/LVJCmoranmy795ZTPmoCJ9qPFKsIZcpJ1lBNdlozTB3
3IbMKCK6cetwlgSgBZSWGgLZWkzJR87y7TgU/z4gevyCYZmD2Cpo0WdWGiSvxtpFSppgg1kvZ1y7
v9ShRKsPLW0b2B8KqRkszlzww9++g3MtHwz6xq34tE1Uj+72BW0GP7hfkveQPQRfAMQpdbmaPlDB
+cytpYS8I62FWhNAEqO9ZU7Ua4BNn5z4mbsD5I+m0CvVkuWbzDQvIbuuhnCVE0PbcS/3nLdNMAnX
XPBhFrpWKuMdnbiJOHyk+CBjXNVhmjnrd6TlDBhhdKLxHV7IDdyfAHAvsN0S1/zsESIMPtLoDuA1
rgFqUxg+kEVweSEOutVSmiRyy4WCTOhodgkQOf8cYtFZafsOAPITgaQxQL/MyodEEq0eEvka+4QB
7rlWP7A02LUEeVzyrhruT7b+iRcOGzijSoybWpEY7AB1TE6p+fNl/WfCSt9jmKt7wY50zrmm5lt7
p9i238ZGojl7KcLdQAnMPWeXV/WDVLnq6uObuXyPgcQ7M1xwFFfXRBBo11WR7y5u3dCWMmgxeH4i
Ic7L8zpJB7qiCie8dAC07c6M1i52Cx8R8O4n/6nepTub4+VsE5fyDQrGYFgtyy6ADzhP1x4yDFau
RAlfW/GWLYgtGByuwkonM7KrN2u6mpzT1+Huh65cdrQUCzhYNxkw/OYT2Fi6K+EsTHFVj3J3ZYKs
g//tEYL6/MdFDXWulNs8RzbUPEektdzGpZxYJ/S/0kpftYC/saEnlpbHWMOJreAEW7bgbIRIpkrc
NavDcr+6KwUYztnDkoVry7it0bPx4ceiJ5SOmuoTDSsEev2ST2uJfd//mt2t0TnEdmBHf6N5sDE1
48OXFktIUb0WFNRBte77rpMkpVIf/QRiOOucY8xJVV+e2Achursd+Sd8rTZCnURYXPSeev+EDttA
pT0QvaCcTWTHQvBMg3wWj0Njzj4qKaTnvzRru0LcW3jhujSxuPEFYoq2XimYF5pO18ePiDfP4q36
gRXj9wXmA3+7HDQBNPkb2caatfwJxEUrTcS1csg8FIUwYiHe96vsbN3lm3SnCjmmpZ2p/6bUBoq7
jJ6J0G5Q4BtpUhisJt1XxW2IVisOUD0GfGqXF/M8GoAm99V6ZzeuiNFAmBMzGYt0PkD2pFpu6E6f
RTIIvyYloio2USHQXVs8e4cvPGmGUnwpjjs1Vqmppiq36ptxcQZT3i5+9JCZPSNno7e6prLvE+4/
bSQu2bTGBP8lYl+ov61mUux157kgZUCg2hMZXIki7e2Q0DQXYuQ8MD/WljIznCQ9npVzodnhpjhq
hjxppHrQ2JkKaa8RWkZnCsylDofXp9HvL+UWl3LN51+x5qIRfre0pjdgu+s7WqAbOWgZCefoYcC5
Wzyzg4XtTzwQ7169IE6r3gClJ7oPIX7G6qavU1FRRsPErHJbU7UI46d33tqOQ7UF0Pv6jBiX5JoZ
gLvzGXz4mnTZCDDtXZus9ggs8QH54vMaj5/fNDXdMs4V7K+5VygSSrV6T2a4AJXTSDhnM17GtTB8
eSh4uzLbDchVeHm2FNWL639zl+dYMgyhrfCf8EwyUWQnf91mM6KmP4Er/g79gBfKVxbw0OLXrMaA
fOjFYNoyqZYyXKNmPeJe8mSEaT6QVZEn0/ehkNhBuvqGYAmFFKa1T4YExj33D9CQJSOsFbS+JnzL
+k/B0mhDsrYtE051mdRLMu2nNDZjYQthsCM4H4ZT9vIbnjI+rXvksASMdW6p6updVTrzeA2x5AL9
z3bS0BRizvMT+61LpTebSnuuMub576+frllpIXn80Dcn5J4G9ZOwfnsTMMR1YS//q+iFW42iKGTr
DWa1Gb87EPkQj7V3n6T6ZckVUt+hUjpXnz/p5DmRBL7/57vfft3yVZNFnfkG3t0NmvGUK26BMSCZ
7n6pKGShK51y+OR6lEss5OUb94X0PWqCKmwI7puKV+ApaaLm5VoeC4roYXJd6WxN6Nd4FuHdXla1
fqcJ8sEb8m8t32N4XdIUvD5IQexL9tVHa1gBksoL3EG9sWrDc6G+ESPuBc+8Tz5sfYxfxmDGqGBY
lFFefrJCXGSIkPQtjebs0D/VJY1yvEbz0cqqckAqkeLBv4mSaWDSEFxfevkT/ETLof1kC9d27mlB
RnZbJvvP4+gNs8mbjmKQAaTjcT10YmdfQVbbSSTw7BgHva1E5HSahiVC3L0WOYd/nql77j25Ra1G
ZAJ4l7HlPSAD6VIGw0xbsx3ougmE9Zn4xUPN7YpqmYeqMQR7mW5njym0vySVAKXR2mRUBjcc8dsz
gfSQD2PdtlgE8X80G9VkapxTD88jxBPQ4lHBI6prXnvqGV43yjY+Ngc68HmR5V9amu3v1X8aVBcm
0M/wcQbtNjgiUdY6z1WJW2oMX5vMZoyeSVLbQW5egnUFqT+eSlbTGpbzLp9rjGI5IhMSceZkjqhn
m87dS5Vmt3fVwniYulmOfb+EMAwSEa1wgeoHy7a15X98vtAIA/tt1dBk+cCk3+l2h3//f/j2LlNm
FemqUsQBZslThFs8lndfNODrFhl9aiMe9Ie3FMwvLZb4ffPLi8eoWeyJ7uEW3PRodW1bbMmfYVoC
PWjDRWE53YiQJ8lEETiq5ItY5t+dWUm3VGAlfetrXv4ush0Bmn97zRnwm1hgLFqSWEQwad76pacw
y3urGgZAD2UYG08YWFBw+uU3HSgNkAnH7ikJbVgzPSljLU7PQ2NVPEe4jgprCDgLfYVnlb4rljoh
cctmQZIx7ptAsSO5V76ZAPSabf46kNotsa9JFM1WKq+FcKBthpIEWvwpoSqZJtor14/VcczYWA5V
wPhz+HzFfLal+yxhbieW4vr5PuYWPHgP988rpVrhoc9o67/l7WaleNf5PJw4iSwp2OkZEZ2mnrRr
eyLsKJIhJxvxqvtC+sTs98GV22JuDevlvqT3pw7rzFG3CHSjszSz+eYIwWITjeI8SOBZcjmuaXcc
YcUA2LTm0ncQXVYfboD7EG0E7wPr/zTMXi7VGWAB7TuI/lVEK8wYbl711bMvvKYFchtj5sBXJfez
hkb2f7q2hHYNkAixy9TCd8dNrXfr3PpRqRQ5a0andqlBP7QFdKss+tNBuV3G7xEvG1rxfL7gUsJe
L6KECdGU+AGufK6r4BacpB/jA7N+wHP/vG6K7jS7OTDEjpXlffPzu2GTfViR9OX5wC7NvRDvRNY4
mUYUYeL2HHhGyDL6jzVAKmZBWQCUpabaLpe8en9i+CZPppIpgf3jcTfITHhFE0ZDjfe4vB2xgblC
LcL78si3qui/gz3ckmVXzDAjSoexCPoDdq/l/exPh/buVBDBIo87icRfl7XJPBGHzuDrdQbASA7p
qVVOPcBWAwVdjkX7gAFeYGzaajqQ6Y/NY5O5tCwhx04mPBUehcksMCcN26fKABYBf2vYz7RfSiCJ
ILZAi+iuoG7S9zSPiTzURmrly1hSe94ufQs2IpKHAc9Ls9g4fxq6z6Q2KctHHxJUC6fQE1a108Aq
H9smuBlRD5SkvHAqVyZLJdrmltq+0RB4wNLJMZON+6Ro7BGqS7U9L1wqLv2ujxWmOeDtK9cY4aVQ
/+gJLPZ+CWCgQR4Q6MSuM02jH76hKfpBOCjeVXTd5Ljf/hJu1rF2u/T3sOCnltAq9tC6UTlUCcFx
0CZ/dNW+SYz0n3KTs6tMTgDI08fXOXt5VgaDhNFRAofgiVQpSxRrEpn5IflScFYCfeVwt/lbA4By
3Zkx+9dSuT9kKbiFSKWdMCvz6AqhhIClI5aNVh1CTgbY8e+hXyBh8ylay/ziO0eJZfAf/QjWteiI
gSMsHIWD7j3H1XZgrKK/FVfVmsz0LmJMtrmU+ZIVLrdZMx5WxmgZZWTx8xFbSFhwEcUsK7ysGm2T
bsqpvRNGN3KkSSMb3xCCRW1Apr6ORXzLBwiT/aF7biLVkd//OnTjfuvd2YTpqNA9Djz6OZ/fg01T
k4KBMU9oBsc14ZITk8LrygexHvMvvvmI8Htk/Z+5b0FinN5SBdZ6b3SJIFWRgvYsjH7H4oMN9BVR
bhF26z7djoy8tS2E/N6wgQ9TYnGM+i4scagAeijiMWxyzc6Z9i8sgIbKlyAgr52HACplE8PDMUeq
jGyW5F6/dkSyJ0RBEkCXbwxLQfV3bHpovVPJJRC5Gr2QPv0Om4wjohhDOVIf77kjZAXw2t9bt/qi
VU91+FjOYio7Om/se4O90FdxrYnRf5C2vlq8CeibcGloySSSWQ140xuXQZCiYfgCc/Cx/n3/NqFN
MuFMGVytZlYQO6NPlCV6AtNqSpAEa8dwl7dEk/RzHvwbHAt6Gs8a0pKCLFlFN9JBdBt7flrQmzlp
VLFNzkIAEAyx/ky5qI9b+bBMIjAuhCpzCMQXKVSxMLzPSKQGY8zvkvYY3MuSVxk/BvtFw24mRxA+
9xY0lOuOWe/zajGK5fP5bkt1iaaQiS4pPv2hC42r9n0OHDE5bROhlgU/58vwP/o8vgsNHWsjgfLU
8cT+8lnyjPbHqvhDkdeSWvLXIeXM/JT5zyVeUHaLWN23Ixdx+KVWa2N84eDN0pIIBu6AxwI0klFL
7xWl26STzwXsPEpO3K2MGMRpSoPBoTQDAZ4vBVs73paRvz9CuwB+JLQmwz0MC2u8rPFP3Z2MF1E8
GJxcwirbmbH1sp71EIJcwwAhwNkh76vhx8BDA4P1zZDwIEBAEdTwjXXg56JcDe1lP9KssZ+QLqWX
AUYSdxa0qr/0zm9CLts67LF/YNZnrgZaDykCJTixV5Zk86G6FYESwqqZuV7OhFagCeKn0zfcJsVE
tONU0PG2WQu+TfcF/Lbhn6SSqPXpEAkm2zPDhqWfR8jIN4DGA+SvBKOSQmXy5oXe+4G+wUXqfPq1
GUiGzSm7zF6TPVggG0kWdKDplWVlBVZKvT5hfhXBGBcqgQTtxcKqFVsaeyQzyFzTtVg6rRlOTQNM
BPgO/4nRRQj7tbHfDWbVhAfoEGa/7PMWFbXkjP7KYmdnoSuGldapdXsLh+uKyrtlpJObmHZXzho2
WG5OIQLv9ARRyH2S4N6apCLU+K/738IpzC8QJt3DNwwRVy/7ujCZqrz//yj4OKAq3jb5hWqB2NDl
y4mtBQyrPaJyE5mRlMU8wchUcuchILUMNhsgvP1lsdZexcVCBlGEukdv26HT/x1es559yvolt5e/
1jF5HF/mCkSY7i1mHgvjxy2wB4fatr6oAfd/rR2n6c8PLMNkpdztj/qsmzv59FtJK7Zf3E0Jb9HA
4T/hpxcqPVgXqSBUx+eGP5c7QH34qO9n9o/vfoP6IPRvRqY+JWRtViWOAO8goghuyt+XsQTdOxgH
THtK+QEJ6DpKwZVRr46W78ETakk9eoxwz625MiFk1vC3q/tEk9L6ki34DX77rzeqeDacZOmK3yDe
PJTlMzJrrd95ScA4tP7LcSDhjJmiJRfKY2SIPFmCDrRDniOCvAhjD8NjmpeChrWhJrb/l+An50Qh
ia6y7VHtKpFLCPABRuBEsBDSXUionzkDImLx0w8lPlYiuw5jWMJUeAGkfrTnsdz7Et6a4J78FEH/
e2JZm80l2puG05NL85jGlqVid9GH3UBv1ylSLqOh2rATeif/xN5O2FPlgoGlwyf4rDbkipRTUTh6
5knxSldTVDxb2Z1RF+0alUaj4FQoxCQMzuW5fpoJ9Ndl4YpnItVxSM3XuakQilEPyv+yr3gYN8Bl
x8YGh+R09809wZnm6c2/zofqWj0IV9ThKeeAAC+PH+u45wWaQeAVs/U66+x/8Wv8twCdxpmFeu1E
RKopYiS9/lo625KmLAAAdU38eVX2UKVi2Uy70uW1eH0H5rfPNZyYy9Rhg8nYtzRswhLSUNy/oUv5
sSrTo3ASZDoi93SM2n4ZkXwt4JHM7gduUdiOp6xAivNt/mKcSY8GmKqozlBnr62VR8v1R0RdIjf0
3Cey5flFdUOUc0UX69eZGXXOoxYO3DlaVeSfzxIws0F7YPBi2sSdbUS8Shfzx2WLLAvozb3DY5Jl
KPiEKV8Sbc4H5Ro47ZtzZkCSC+FUi8qCvsjzNwTB/dIhXfrcMMSfjFVYdHvuo/ex4NTVBsj07vIL
KnPoSrjc7Tbh1bW8Hp0HRAUCzW68qfN+jTtCuv+iBn4vux6EEmJ58xidUsyFgcvZL2AQw8OAzP7T
X2+AfrM56nwoigUVCkrFoKi0jIOEpr/uHHpAHvxYBelH/lNvpic30Rw+NP4+bIfYAOuX0I91kvtl
uZdCl7ibY1rNGfOrOmi9OeGs445mz2cIqCWyN+FyEWqqjpbZGrUzO13hIjeXm12CIRPd9uVAou69
wO6rnmIMdmzqiXaJu/DS/tZnLnuA36voqNQHSHbpUzE/iOAWOF57clhZQ2W9ZOTXQk1W1Wr+RxIM
rvgfnimF04Aq9kMrsOamYvbxyxWC6Vq66+YiixYikgiOfoezdzqEqdTq3c1d9GmyXd4Mw8sfzYW2
1qZnTK/reaLIRUTgmzxGsrm+VdrBRFJDmH4eVv35UNjyQgpshWNkCy1T7Z7G14edRnE+fZ00Dvh1
DI5WuYyIoZDvQtbB55QCFGf1KLKpVeDI5c2Sf8ox++tdwJd9P0wo6PsfrNW0lOUtSv5mXct67nLg
xkvZ13KcSu69q/2OjjwfQsQ10eMVK+RuxBJsuRjzyHCp2cAk4pPfy40hmC/Ix0a68aCDE/1+Wioi
5CndXIfd49/i3oBC8U+F2tt/+dcf8WXXePz8oGR7MomtL3V7vYGdHKoC5a58zWPXIERsSxNfaObR
1EmNVzmazcCRA2iQ9gtv1z+lc27KR6W0MSb8ik1E/YXvnYRx9vuysmgwio2iZczJqfWQNVEuDR1p
bFzLU9lL1wiuMpze34NYmOXSIPo3ySpP9EztnR7hdpuERmzCjyrnB3ZODgoiH/0nE0KXDmaCQDeL
XNdEodW8epwYKsYIuBEtMxVQQXl7OXKo50ooU/I2nVS6BSccr3WnD1xZKpio/cFxz1e3ifPiATT1
SbCbFoQ5I/FbBuQ8LwIL5U4InmuehZI9QBGUB3AJD7IVi4qxz8PTJcd2n8FPpPR2HjK+bNmJHMpi
eGjRixMc/Zugws9Frrr2xLeof4Az0snufD2w1BVnfuqHWeUylH/XzYTChtJxi1csUXZOowRQLxpa
H8CoYBwf7xSD8D9UhOm3lK+ACH+VH+YOrk8pAN9C3SloVCFJW9MaEuCFr6hc8JedufHdxXXHVVOb
1srdhBtliHNNhragzGqLqGj7IJBUbtJLJLNsdZRon6fmvKgRnjw7xrma7uRZx06R9KVkpOptl2wt
EhwVZYPl7ytzuIsV7EyT1hTVQsDnaBGhTI5Ec+EIvvYNJ9I9iNfVNiLQkTAPPUHSH4GW5zFfGVGI
cOtO322By7o8Scifyv/JXXULT/nFL2D6cVqdr0+WXKVCS7QbDdPbAHEq/821lmezPUp4Er9t88No
kLdyvpSxDDwdUiDKdn0g+Yc/QvLzmU7Sy88sjCjLX5l5olewtE3G/KISJ4TOnwrKO7FV3F/Rx16W
YTLT3jzySJRuvug9A/HtKi+HyvDeRZxb429Op7KxlKS6fErThsHeGQeG6WFKA4ISefgZBMrIq9hJ
smuaKtCThgEsT4ZQhgwT35zceHBvO7vkGzQzt7Pj/aSnKvrWOojcVcUbcsqfDoekg53DiWTogTbP
M/8UfLFkLB6LzdVN0eomDi9NRCZ24LjQZYlrK2FIhdL0ZgUZAbXqA2vEmMgHNrHjqQFmo8bSz0PW
DF/MA1RspZyQtJbar/YFGh3RlmGvXHKVhZD8jJMnnZ6IAJJ8GMqVyoMTdJc29qt0hykHQ4wSsFrz
FdOKJK/RWOxugO9hHA/F+krfCywPlNMdwtYJ/8gdmR8QFjNANWnIzRVE1mc4zAEEjAIT6MkuR8Eo
jGTiIcIjs31j/KM8fdlkkonIkq0EuX8fK8u8hkOq/URYqh5ImQg4Ub97gIh9+YFSd6HpDgYRRKYJ
/CdSG6MKmHE5eRTcfFlKCHxRkyGYKzvj+XP3UE0/iBJsLxKDirb+mpCX5j7GpPeHC/wiOELWCDpc
O4U6h3lP0fQwaFb+pDquLkhO6SBkaYHsEoVrARLJINR6lDLbymlMpnHnNg9fpIOdbK7mFSAkFHU2
ODfIEp3k8ApV5jpY8A3IDlqIPoW78Y7hpjaBHGMI80r2IcuJZQhupDvRgqNg8AjweDykbYFNsO3d
RLxQGyb1At0QQpYuUKpbl3snGzT1nZ2eXMYtI0/EXHB1OaReRwFcwF+KkVz6eYwv/9QZ+8LfwWAk
k/GTlUGHbGNDXMOTYJQgfJvKAYb5UyaIeLBAcke5F5BYwZf+HBtYPcpc+p1H91XeE4/19K7bJ7Ed
DNBsEkKqUAngjzzObHb8VI+IoVCnM0y9pzA34uWe/o1ZwUcvzi+U2WLZ+5ZUpg9juyrzJnExIESy
ijsCIj66HGlrch36VU9hMrbTvhU7J84Pf3XSi1c4aPAHlaHlgxjxrtsnVYLTYUVDnEyYgEfe3hyo
QeM8HCcf/9NLUNef/VlrCKsg299Vl7MSqSHGPtlIc6NntWNiXVo2c4FxGeCUZcaP3q2EhKZb9xq8
YG2S5Wwf2l77L70iRIb3GurdZQQghZTy1eztnEoZNJlvzt2hyOUcYybti1k7LV1tehZ1TBSq9Fv2
Wa+0Lq+JQLbcIK7oEB2PGSkwC4l5w4Eg0rjlHV1VRtiMuOKUdpOSfAIJKSUWcy7XYmrd6W5pBdvR
PkhX9ZmsRv7/bGcgTCKqofilui2MAHcB/jgM6Lq1v+HGttw6Is5plgt+qVy1B9MCia9S8qp5tBww
pwcHm4O1rjpgZHIkGukYTugvKoPcLjveEkAq11SFwxifZVW0tjJc+6rGK405yf5X43bUSWK0BkfZ
s7pvy9DGtGVIGjN4jISjQZJmw5FiyxrOm8P453JZzswgilHNYT4T3wTajq6Ow9gVvc7Cuj85Kgtx
b9lRWG9YsBqj0bhPBfAKmmeoTbU3/aaviDjTCk9kW5vKiM/jLAn28duD7Evo+kVDRK9kZTgjhG9l
d8UgY8vgAmdZ+uuSYJetGcbLftRAhmNsQOHn8D6kpXjM2NRy/JrCJ2WfTSy7Pdg2AdSNT700h9DK
eiXKJItrBWlnmtX3X8ynYuZJckBk/wCAyUriUNuWv97GEso7m2HbOdsi1CUZcSV/egCHJ1ac+SZd
aPYL4OAFnIkQXDfxGyiG+LYPB9C7jOcGSfsD2EMxkckwnBrxts7UENOiCuvfSKucg2ZM1LAtJVlx
wa9U/Y+eUQrX+4N6Sd70Lz2SuwCvkqiTPM6gDh3w+pxAWjGfrwH4gjLvDeJC7sWqzJKKtI3jpPqt
OarSSvLOe3w4HZNy+6kvFIVXCis25Vy7zZXgGdXTzEOql6eZguAGZs9dVZCzFk7nU8thp3ezkrIb
kSsTU2Wf0h0Ca9n58vsPhZ81E3Mdehslh8jKbRHYGCqgN43yIr38pqv8P0Z+2xsNC47CSlqfEMSb
nYBN7k2jxy1sHATxgawdkw5JjfTnHFaUrMmqaBNau9v2NgxwHOPFHR6qouofPXCYzoOnBG5E5Xsd
AnrOf1b2dT4H/itjKvO+gIEHS6aPOF4S6h5JTdacjq3ipKT7yxv5b5o4kEqMBx0U8Vxgf30lbNri
FqQwLemPNDSw05Am1zMph7LUyg2atkM6uXQ68jo5bNgqxUPtditAAdZJ9UvCFrRhaXlqJcG1zPJS
BcGqY61jAlWTAamDVs8A+zagnD5IO5+avNunJ/AoHcinvAMGVkQlguaI6eTUW33YHfIoyiZqg251
uGEiA5cmXYFEheeW515nZnYANeLPMAYLBkmWgU5HY3mDwoVsUt0AqBOarfwp92K8e+GWQ6gtduTN
FzSHSVqHczcz6D6UnCm3o701e1dbij3Vb3s2pjUiGRcS+f8cO27HIsnQ8yzqxV9DVgcdrhY00jVJ
zdWfTVtX6s2FZ9q+6dE8qe/tJFjOECIgqL6u/yk4vsIZbGOgyyJ9G+ShgiHA/oxhPnzlE6bnvaru
JCLZz0U2Q7prH0EQjMHXrC7aSJhXeeiRRFBZ05CnPa5atAj0vC/2v4wosq4OwN8/H2jZSK6dgrxG
OZoOG6SDrQo07MvBpx/6lpx9S7tCWAVp3RkT0XT+g3zQYaebfcSLS6X0MCJ8YRMbwlkUOBSDLmyZ
NSBHLP6fZJZ+Y/58xmI3VD5FyOVt7+yzspKVDsYpCAfkUbLd3dqYNQyAW4NoDC2JDhndFm9Q8t7m
mcz+Mv71ZSVWVTNsZde24gwg7B73WU9blmAArJJi0k+9oxdaOudu8jnyTbsONpn825HYg0B0rTL2
FhgPRy0S99PqWfbczrxwH6r2DhsooUqgkwS+GWBZGarNDV0U9adHXBj3OKiBLEYeVud0yP3g04gH
KyLWSlRdlJBtM+dVJ194wBtIjJPtxg4WpK9/ZIGwzNaqWY2om3s6Xi8HMi/bJdBtxKWTElJx6caB
7Y2/CNiRrlNuaR6tpGPCH3Y69ayN7ddo6jakVUHI+GqZc5N/ZSszbLlo2kQW8UapvsxBmYockKSk
fhGAzdiSjXg4sHp1oT6A8lM+KXtz5nDPoQG/2MVTfRNalVGLwctoNSeWHVwRep/OVZZc8/0eNdlb
isBx9+ODBKIFBJnqMTvOmRxiP7YTn9aEeJPtkSQVTlQSm0MFN3wk4bwRwntiInuKjB1S689LpbWs
GLlflx1fcY7tU0XiRXoHk3HQVd0UVnS3Pb5+oqOpBOHy/tsRdwBxIu76LUd0tpjNCDti24Jy3uE9
8a/z4ebv50He22n/xapVH3CR0r0Ra7lb5G5qOjHeUAcrzHS2uWYHMgd5n2zvczxAxNDQKFAUpOML
0dDjh+bg6IYgkha3EyJT/TML0hwiEaLlKPsX8DQAl7k50S0VzOsQkM5EiCQxcSIc0FMeAqydIjqW
OOvITlTSpfZKueJbPJmxATLjwhdQHAXMfN6oUfq3qUHVIQ40vrDF4WwJB4+bCT6o5PjsOA0Re0ow
tivRxUjpfxyYE22Tr7Sf1WI0nbk5F1C/JVcn7iZe+KEHEZ/NazWOaLIOFkitfesAWdFhbHDgfQ8p
+aC8LqIXFy+l9ZRhg7fTyonyFiA/MvXxpA/X6rAKuliQqV1SVK37BitWxvrCmV2oGJNjbkvcjbK6
k7GTPXtNa1LHQk0l6JvwsJ6ZdocqW6nHJsMRWeWBgcijakYsFxxU//4+o6taT2O3RFRtdf+IBpbi
dlhLWSvcP+zjMQ4FOSPwkwmWhEu3V9aYjfa35RuKvhSiEqniS3Imk6idym1XLmJKbZiUQ2wTZpaU
fGrxfHoyppwsnH5BKTiycrgzoRojwCo1sKn9dsd4uKgDPIJ3tDWQyW2UBSc2OIy9X2KfNjhm4bIL
n808LmL+9gAEeKlM4SXANI5oxyzbm8LDkmd+lz4qPzTHttk+IpCCUiz3QlXG6KQJUK/CzPjryRO+
J8KsiGmxTYByxqZwjnS5epVCGrx1ppNRlISUkYHVMbkFfly2Qy1GdaXXi/W2VPQLGY7KyBv6MQ5b
WytuHLs4z50MWhuIxsnWiCpzni3fWjPh0DSNyXsC+1ENwWrrUdqZlUVrRBnkqtfyroo3YA7YMMah
uaYZERnGAl1TD6FDcsCbfp7pzoo86BFvOcLG0q/mPiXLzsqILVd0RU+aVSJFguFvRwOTuuthUppF
MgA4mV/1+FkUGqpSJpru+jufumnDEG3NMpal5zQ1n/xDBvJLwhh3Hb+fsXIAVxnQ3w9a69xMgAWA
18FlqQNZtrMyuH3Z0g2j89TPIvyqWkygmM5RZN6p1qZpKRFar6MzkEU8znUQCtPixQ2NSeC2u27j
bOK8lRlphy+OPHrotbSkDLfC9TWbj4Fp9KOTfl37myTNRaGhEe6bFcPRP9w2PMvPSXX2pQ6L5DY0
ahPypUuk0+SoInRE79l4zOv/bVw4UfoLi+Im/MQ4URSPKr6hxAWIrZlnimjTWLl00u71ZutDlYkv
1obgMDM5XINzuHlP4iiXojTlPU4L/76Gwn47Sz6+pgM+ipIOFxZztpcjGiUx0MF7hmsLH1s+qmMv
ZokePxTSYb8N0Im9Fyi1LFEN1t5q1Cx6pFGq8KR6Og0/zQRruGfKX0IDBR9dxfQ+sMPMlQD3yeZu
6yWmZHOJq1NTmq1bU9X0qRkefMRwIBtDxNXZ1Oa0k8/TMT1MoHGOei1UHjlZUYat7c+O7Bg6tciD
3LKyciVQq1UwinqiLe/EuEMrY+eTgqrfeeppKQlJcw0MKEREw3eBnoUK0G6tqdqXISfrYHRkenrW
N0pxlzy8F5WRiehfqeDurKAQElkchYRyhNO7PnbE4ZI/Uh9D3eb4JjlIufr+VEV0fceYBGAr8ea7
1tMHap5OYmD7ImZ53i4VLVYulMxVl7wlTUFaplcb+LNyRnpKM51vIbzo7tnBWhc6OrxNFs14/rgK
sa1tVAReteiLGNqzIk96kIStRggcYpPzbVQNymiXx79QtDQlQL16XXXcVbEa0SAVlMZJNJD3QnuM
z5RfjEilM5+n8bItOlNpJT/dIZ46P1K7Rbyz9dQ7uzimEr4/Izy6EJkUvFZMrGVCSmXcpXLayHdb
qAhDTWJ8MGpy32H16enjdeNOMF5h3n5CziC4qPnnMn31cYFgQLBYW1GFawmAYC+ed6AuU4Jrr0yp
G/kPUEfODFpn4fOFBuMnnCrPN4bevp/hlLpgUDWyI3HMJLHOv/9vKfoIInjxziOwwg2eKzTy+/LG
Du91e+GZhuJTzUw1v0dUqonX+cDLuMcId8IQMcyx66c6rpR3X8gwLS6E+0ktdu96ZtIDPALyOc4I
s0l7JF+h6MTN4T9+YmjXSejhsyz70du6NiT7lBjs68XHUODTRvJt+jl1I7BxbBvFxgRof1EXRrvK
cVL9wELz5B7AKjwisSVweQZZYyGQ1oxDclTOqurtUXe7Pajgyt74Dy8CjHc5y+qIvQbdzqKwgcaS
doMygFtJyIc0Bca+wjItwQHAeSJ3mPDMtojfOIDjG/svETTCafZbULrS8GaeR/pagAZsIQJXLLoj
fBgseQ0fnmcOWKlZYD2OYVrA0YtMIVlR6qCsLaIsr6LnnmJXrBMCJxc2YRsXPi5q1q2fL2Q8qjve
q1ZjVBxQSFxAQSmSnpb0Ro5jCew/0nQ3f8f8cFuQDn9CRGbNlQODTPW5g12F13bIKjD37rXOV/6k
sDh1x/8WjOFzn5QTOak/QwVcmCy7R0hJkZVNAmfl14SwGYRPcjsOOcia2XGL70guS3aMpAvNQ2R9
f7JrZDcpMHKR4GFKtxqHAw5tHaAjWEOyJBNNfQbPyrwvCWjvSpjwK9VTQQYs4CtpH0qyf7kpb2gg
8AqDS+NwG7OO0ESQk/XZr3+hv3uJFNIk8gdg8Xq8XUuhchXftB9p8TpA6lvBUEg8qEW7fViTJ53T
W/aca1TspBruQVffsrCnISTnrAD2x4t5XITrLRn6TewjXp12tpVKlRDkGp2+Faxg3IMAPTdGh8hr
4Naj46qLU8MJMNjc3acAK2v70xw8AeJOG+FbCu0aGiboueBhmTi5VBXX76wENrtQu9VwDJnrSYQa
41+QpeNnNeh2J0IbW1zqcKIL0Du/kJq8eq2Pl6YD+YK5FQBD7zm2eu//OFCSXMPDCM7JO+xY5u3O
5aTrpkoY3TMEROzsqM+iS837n8Lc+XTTxVB5QCZ+/04AZqPy+LhJ4lBlg+bjbduOHUo3efohYIuf
lJhwsWIhbEDZs2pQNjOIH6Htm+69ONju1d/CBlSee0zLMSbPQ3g9IRd5nvRoBCUVfxw2Md2+UCUH
cHx7TMgNuCL6XbxUGI82wZltXl9BSm5SYd/m4/onEVMTfI0CjY9n3tTEfI6xVtU69d4TuuRUO95n
NxG86Ttlprg2MfrzyIretgGtiTneSJ/7u77x/V3L70gLepaYR4QH7XpFuog6BhXAm5JeZfWSPr4A
9V2gvsizkvll8x5gw72fyfDiUUJFJcsAhedP0TeqOca8mWL/hLZ2oY+CoKotjLmQ9vlan9cJdCNT
/LsXm12XHpMs67uOpci6fPtPYCbvq072kQSN4NeIuqrRsrHpySIdupFt1BFN0nbFHPSq4zercXOm
Mk4vR3+e9n/ksbg18Sk3Mf2SKa/dnEscxMlgJT0ZILAhR0pH+VV2et6roo5jJ/NS+XiKgyuz9fsE
/xPBlQ5ydJxY4h70tYCUZfcWqf07z8TnN2OSVTEwMw0F7k3sX6agx72or6rWqKxnhcRCqids0KhC
G2dcnS4lJgX+z6IbsVsJeHJcrAZ2YwjGC09lzNSs0nrQqDAe/5Bo14MjHNJWokGN+B1cuAQchEwC
fBL0hnTwbXALIXlnC60MfaDJOR6++fYuqMbGIetGIi+LW6FBWqehtugEOzyt30NQcP3oOy3ke3Dl
MNEjxWnUxl5R0JCc6oBhogWzbWpjiqSDc1+qOTIpAldv8o1GS23QSP8HWl/182DzZ4OAU6nl2MIx
b+q2/VD9sCFWKsFfR47+43dDo92As5kaBRJSM12mY7/Y/tZLiu5i3e79d1M4xZyRF31s2k4GYNUF
XAogM7lDdGYx0tWNnCxb3evDghye1G/10D7ujtnTIW673R2tAmUdrSLcbTZQ/ojoSJdqMJHkaUeI
keEsTSG1xsEP0gsqbtsR6o9LKbpHJ5zXxu6ujnrYstKadpyxSioP6tuRoE44V2JelZIf5B0chuU8
f7L9/NOudjj22/AZMEF9uebbMuYWMGAzSgKggWZw81+anGQ2kbqY4fR6dbMKY1qCyvCovWcU/QYM
+9pHlMM0gdVI2FVjTrSu+Zl5mQGOhqGPWUp/fJHVokqmES4eCv9Ju885nCAwrAd/mGvBzZj3zyXE
vbhhsJTStLTgeDS/Z6jbNkgzl8AIfHbwg3WmjCcoFu9HwZ8MDC585zOzoPYtO3qbUlLBWl2Cz0F3
jC72E3sAzaQIwKJD3HO1eRgc89s3ZTRrNm3aPtq28pf7IfLh9bfMEacVkQUIxheYo1mGIDAkMHuV
6AJnlt/U65nXiCtcAcIuGS2zd6fQg6iB3nBlU+z4un/6Kf0rugkcTExrk2MoQQsJJ2xaj+5xgJLY
ctVp1L+cmKYtqXzefEDW1+k5S2x82QEP4K6hHlMA/bsRJ4MvJo6qhYJD0mqszoN/KjwrTyDBtvda
i6dOsxpab59SdSu2V6Ql3tn+WrjnUKcl2waQu1Oszsq7BMjIUWjrIxxWT8+uVyv7GjB4Rg3IhtFa
C8rpU6Tan+fvTqWmTjn9qOPW9/NBxT1WRS6PIuzWgznEzU47pgGr1+SWpTCgi+U48RLdYw16kGdH
wapfhAMM8QEqjFRZaIUC8Guy3K9PyM/08HNdZl01t8ZRKVcRYtNmtxqBdkoT9+XU+CATyIBlAqa6
WJJIV7HqBGxUtQdDz4Xf2EKopfq0Zwq71izZWdrXreEivawVMyDQQJ5qrfFO8cgu8i8uXjYx8y7V
GU2d+8k8xK52+JgNOmtBtpNpHQ1SQV6LnN9YgVKGSAmg4LyHZad3WGfN+yvKCOKR5IeTqYotzfBU
sjpMFDKGa1uL/Otp8JHF32yyz7vhBu4a+R1jr1R39W52kr+1hWVusKPs8Lh+lgpo9Ga9n4DyTpJi
grhEOqf9tcXePbrWAymQZuLXVm/yiKqR/y8lhQunlN5eA10eHe2h2q/sK0aCq9VgLQLhmOaIt2vz
H9oAtkShEzRQvT264WhYxJTssAcTj6SMmHkIkW+OhNDO28w8yz7vEA8FsrB53jedx0n/t5B4cmOa
MzVHnQSFQuuH06aUfMJ6C5R+/wEDSdL+WaItETzj+ykoc/O5j/ouP1Qp3u9xx0FH7+vcjivPTmW/
i/YGE+3cpWb0taa8kcC94RCJrXhl14wTU4DOH3uFNBhkrqZQOR+KTAHLEtwFuVf+eQHN0hv01mwZ
QIawsFn8ZYX5Nx2MzPPHfphtLU8KZiNja3ttK77BGeTX83bTUHB3DezHl4TWVgyzGTIifHnewHKS
2Tj880HQTp6X0js5DY8bkXyYvUe63SgVyb7RDapOQpYFfL2vv+WR6wY59YLiq+x1XChPOy/1DAR+
HMDOKxzAHD98DFzZwkLsy4esw2s/5RSD9NnGNR6Szh6jOsmzZxglQKJr410EpHHtVzOSNzd59Xiw
fCP6OEej6nxHl+Nu642wkSkGR2zisOfphl+wRYhjY/fmHlgla3lKjWbgOXJUmiIAld9jpbYD0mlu
dANqeJ3CaXMIrF1O2Qtw9AlytlNLp7xapo9gW3m1XewQgIPq4CYvQHP8/jtRjWma3b6X5iDV1VLX
9S/eyjVOAy7Q4IGvh/CIITuzeLd1L6FfDUHsgC1y8NFFcN2NPaHScBYG9SuWfTFU9CM44loFem7v
ZeJxUiPentQJKisU0sv9fUTMOcuGQd8LvPQNoVXBSmd7/3WM2hcOS8fFcuOBhdkeibOMlA5xo4sg
TMk8J0MFlg0L57TOqVY/L22IY4n6gEHyUV97oRIWVsPd9Rciy1vlZxDZeNgfjkknCp60tFo/B6YZ
VGPB7/Cnt1e94p/bejShyvtewpx24fl5i3SGAVPwltt4Yvke33k2SGfTPuuKI1EWmOEUAgOFZmZE
yS0oQgxnHmZApNYac7hiG36RGNjqztx0dXKXFfB/DfFIKJ74wnaWtUMYDZrmpc7OxbNL4nDPbg7q
QdkQ6SM7Z8mmnStbW0zdq3mUELKrCfeS0m/iARVtzxsV7uBdLVS5mmP9Jj9sJhbzqeRRRbf0iuYT
eZ9uVlPbsciwc6tTA9ugIuu8Gl9Tpqwgcb64fIiGdWdRPUkp51cTJKJ9WOQ+P942+Hx+h+f2X3sQ
wylRKnYrsqaZhqHxMc53Oen8IJWg/RusPbHFq5E+gUG/X5rm6Mc1tkY+LRO09uAjTaJeg5w5L9M7
Bit1d2lwtWDa5Aa51G/OVDEb0soTyd8zHgEQjWDwhcpnYjYwmkA7ax8z0MfWdI5iiFagh12j9Eoj
KKQbbFUL4JAQW6mLmjn591Q1n+G6B4JHLfhwXcGP8PF6AZqQ42b6j8zZjLKoKnxdccs9tNK92hk3
ko51f77+MhjLpFLXq0aGOyfInxMHf3SjG2i8uRChUhnRBpEJLRbkF+p/ZmqIwYe2pvmN+OpiVmwu
gS3rSaMa0/goNlRmdJZzLuVPKWkpozA72YvSfCxM4wKyOun0ULVdy5B5WKpQ6YzkeOeWw1HRieTX
zaLpLYgTRwlY5yWHBWgUDFgN+5ASKlInDgyHN83aDTaNOJEyYrIqpDystJygkusjzIvbLOKRAyOK
wvS+QRcfTCdzvX0sd40dhR93KoUTcU/Z8DMIi6zXgcYovnRyYodQZ8t7ugPtTv474KemfE494r4S
+PZyRtMI31RP3aavPxlLAJnb50ID9fRnDuN6+1lv+qiaiKyl110LjjpPvUFfhSSxgAAEkpPbmYFB
pvXcRMouv9VHyElLmJsgmji1H0xXGYiJl6Bkd2rW+xJGb1T0kVKsCubjNTH3+wjFqRn55jZwkBqu
w6ZIiWT/oSP1ugj83GkCeRaV5cSjTH+zV5+h3HpYbkl5JG20dADnlP4UTT0RixVjT6uhHXR7657r
+ukjvtZJopgfmva7uMwF6Duqn4vct7qpf9HDnm+wG8mC08OSrSqgxAygZuJ4fJVMQxmXYqxdQBDH
pvHd5JitHRb4+x6SeumKdhI1GPtMVJk/21DZXMJiFktZqQvqGxrGSHeRih4YpvwG4MYU3Fc1dbbs
ijAwjkX3ju4VP/YJXDkWscMuTnMU1MZh9QtlgXCO+qeNNLPdnISFHrSNJx7ieAh7Z82cOFYztpU0
iiPx2kONeZpdGU3khR1riPQ/GmqXoCHuhwFiP27WAVqxnI+pMXfn8M7oZn+eOJlpLTmtRjOo82Lh
5RlzuWzeGxbcSyvZTgbqWsYRflnQ7kpqFcwjLaRJpt6AwzAnenKqgl8MCRX5cqpv20R6E8Oy+hPi
4rTED+Zkr++pEDEDgW+QVJt7yHPj+tZsiLQtP4eRff6MhU8bmBsosogoKTXHn+m9nwCYVo3sSD5S
N/uK7NyFHx3sULCuXVmoga6YeNoTkSOw3aXemtXf2lkfOTz0ASQ7EkOgaCNuQJ26mXb2Unq1mpRa
GbUiWhSE62ITnEalRhqhTM9+3SMjYriqB1HVATswh0HWqfNQYlCnCeBL1HPWGxN5iZecFMAs0EOq
VNDOtNvLloX1Gb5ppGw9QQx5bJO6MSAaD1vm62Fw51sXma8QMglUaI4fSHlt2YcB740/tOA04AUQ
9/KbMd4j2YgTUySc9mzO3Hl6atAtoieAvwKxVfcA9SmmfSR8fnv4799e75pEH20u2DfzAdgimvRt
YTHzNcHfpzpMTF4fl7MC99m0En7MGcjN0uVUG3YvqKGr53e0OKx8ZrfquBqoUZ1NYwFv5pd42YQp
2EZMYcMpJgDx3AsZm5CxH2KAYGZ9af5J5R+hjiU1uQdB9THYeszO3CSjnNS+a4J7TXe1UJsOj9FM
OIWGimqU4XiIe5TZWSPYDvXhCSNwanafxX+cSOtmL+neKXPNX5IYvMpEFmw595nR4v7OaoOsLbNj
9/bJm1tyEJIAUomuR8uF5rpG86kTNK+vtAdPPWQcjSJ/h//jSlTSOORPk7xP6JDuC9yxP7Mum1+5
UunpTJ3+WCZaVmk6/akXV2uKzuLGVKZ22Kbibcw2ZBfnK/pBCwtRcNpNNKw0/0QDXz8uMFosptRR
1+RPQaAhysvJKHPcFgB4ja+tnEGJCAvO2z8DSOU7SVHel1cIEqQDlRLdi9LLjgkiI7FCcEMHWaw1
ZEfLoOYoKI+m7o9m2UvLw/yjGC43RDoKVMOa8Z3P8+inOBa45gkaBTHiry+jrXjUEoD7udDhOWSG
LFIIPC1PMOUTOFSbIuypExY5jnsjicj97FZOY8zFWQYObMbvIfcbAzM+zI494kCTbVVTgN6SUfTy
WBKRUL9V9TNXs71zrd6SNvMRrw+PmRsnJdpAOU0HymAKi95kfz0S1k7tjbF7OnYHg5YvZRfG9iCN
bvfwsPzyYPfOBFd9GSsfak9nKzipX7674ejBQ7NWvrJi6RhnIAdL7x7zJWj+Ci/xUFZJ9lthRs2X
bgvl/MrZ+veFl9Mqr8jBks4qiSG0d5RdEMY7bubeuNWu8DKxbg+V8w9KmtxL7W+Lt2anv9eHGmJr
BBO9duTEYn86v4QEzlDXaRCK/9cUEEtjYQsteTC349o3WUbR7v9AoeuJry4zz3ug9Ia6v/x6i0or
HumFvg0TgT6uB7BLmOTqhUhQcFYmzNASJ5aZuUA2GgRKx6mxlycO40MKMoDM2sKnrsuqZ4yiS+Gy
KccNDYBtOOIYyCyK+kY38lVRZFDbuea80nuTmQvvNBiuUXQodZLx8hB9TK7UBYJbJDTYdAcT5rKG
kGp4Ra9LKhPFsqMjYKezAlXipaX7CsD5ZamayCEQC5vSM8nsdQVtoMEjeO9DrtG7Ua/BtJGPlpbH
eGk6+mGiK+DRaTicOuRWOKheHg6EOOyHHr0HwUV0BkUc3/nIHzGs42rnob+FekDJ2u9i2opuaRF1
D83h5x+GgoSWmkvDqhUobRsgKMnBaoVXU60CSEMsUOJ0Xj0R/g9CM5yxrMZvmJJm5TiAjkPMk+gB
nwEVVQnc0xzCSFGPLHkokCYxggffS5FJ2ZWz1mMY0ZQumFxUoA1r8cjO5WjN0cGSjUoI0GlIvI2w
5KUEQsvZn6WkVxI5hQNoIQiRA0D/rFi4jVM/ecg8LXExG9c3Q/w73/fNPuAF93p8fFgocMtTpv35
uJ9JRyZWz1tVK3fMSb/nBYATNVBcKEkM8wgdmA2/uZd692kR8TJw7fmbz+ucB1sCJ/hNSFdgNEnb
BeT57KLtPDa8TKvV7UMpClrd/WQQ6LrBmnuaK1cyz8JLsCtGYXIE4Y10tnR0blyONRS1E2KxhNoK
0VJ5/yZP7Ea9dqtKNVrl0UNdc7G1LoGduSpf3nnydZbL8f30pf38fMG+ICwLml8E1wGz1DQLY51t
LAu3BRdHzi7FHzdZjbDrz7nn+HVtZBLQ7mAyyNgSLkMFvIHCnK+ByG8pvqHvZBdtRkKGmWP3EzOz
mh0phh8GpQCrwEs4ADfwthyd6oRrUSNmu/RzTlV2Y0wiRJ/I+l+BQQAO/VLhD/fQ/Lb3nKXNk+4e
3/FHXzY5Ufd8s6/u6WVHjsjojE8mGjj7cc0gsuuuWAJ5GrB1d9rV48gJJCxQYrA+guinPHHKZWKu
ZI/YKpU4AEvi//11q0x1P8Y0c5DTDBrCQTxs8T4WxJOi5QCdCbE9tX8Zpcn+GoQOVElrN0s8ic1W
Ms/6GYOQz4GPxb4CWwDAunJpDExLzgAISfqNWClWRf6/3OKVLPQdpHPpVCH007cumOHiSonsuZ0K
ZfaKw46Edkph4lwD5JTAOzIi56Uy/X7962E3I69e5w9DBK9tH1tDqh+J+b4C4FJBxqlgfEOPchLE
YmYpP834cr6YIIk8NjhBYZwfVGkHPckssfrqkjrNVU6Ron3i46bx5Dtrpl/vDOC5x+MuvAGAvrtR
Idl/BxLRS1Q+8RxkCPd3gZpHjXegNVaAJrOrLpKVvt52E+EYk2cYa/ON8S18iRprPtir4Suaxg5e
RRLIgl8ikwXqev7WkDHYoJXHbESPKmEyXGRT2B69ehuob0zwgCA2jJVx+bIZEL+exoEWEKkLTyes
EzwWlu2L1IkL2NYGCitlSRvxIrCWurYCq2TJicugv8kfxYeBMNaB8mX5qbx0wIXof8xTBKTM4cXR
ZhkF3rycUL4shka53TG+78mk69bsTKaRytj5RMxOV7eV05AKHN0SeKfUoXfF1R2kebBHVJ2hOAqU
PdW7doL+fse0TfZc20+9FYVgcFtCDx1K5UPe7F0uIkghbjolbxzIIQN1CMKimIuHQV8zpuC+8Di3
5d9AOo7Se0GGohYOGJdfExB9pVzIniU9DLZtJatFftZBOvLIV/7D+qbi39oMX9sJfW+3Oa8THrRI
prr/Mv/eY7qzxSUqscN0R/DrMf+4Tp+sbUVItl6sSd0TjzcpcI8tkfIvO9nkUG0qBNWl4swShrdA
FA2B471SLEWyNZ/61He7R75OYgs6xQWKKFtSmuyxw6UC66y3PxBwWa7RyTjWFQ76jIJfKgffcS/Z
4e04MqCjRUQ9kL4QhdthFBWN5bSUsDzKj1kgpxDplvO3y5F1iHHv6BY5RPy1hKPBn3yIyhP9OECL
P60kGsZIx5HoI0q5jHJLrNPQvmz3eQ2V53iAzy0L/vEbr6ckuCH24YFKVTUdldDjIwNbq7T/9Xu3
ohKFXJla3sHUXCjLLQ/78Ixtsp41zR0r734JPIHnuNjMVe0BlOt6359ELv5C1o8+0SXAbYFADwAe
bjQD52lm9QnH/Z9aPYx0uV8VdvV7WSzpmeuZbScoL5Ll4UL2IOEM8VFEXs809TygSbCRQjL41hAS
eNBn5uc9HfJ94EJ9biouXWp1nKoIe/Caqyu6uGfU2Sxst9V0SifOv2Pmpt8DnvAljIc6BroyiSfx
Wc/gfPPaxastelbeSQ2eYYX5vpMI+CFcJiKrEv34LknCX1edlOtIrqQYvKtP6N0/sv8axKDOJMAR
Iv1fDa7/kPlfQoGMUGeearDZH7WhH8NoAAlKyRTJs+/gyTM7PuQC/ike9o6RMy48y7L4IirQFQdQ
x977zxFgLoKQjRY5jKx26S5t+0UWp6r283Fmoux6qlz6qSyof1M/D9DhTi5IaNplNxeUtwg3DaEo
tLoK3QY70U+WP27D2e+cGMN4dfDW9uRGnCAknQ+G4Cp77A6f7wwN5tJISFPVyEXwij+n1NpYBPn5
XqSTivw9FlgQCPd/lwAsozbkdpdqf4lvfldWfHwRVYLLfM2EZKQlPu1ZL5aQPbrBOPoiiahCha/C
zlknxDmzweGWybg5KXSfrRtSxxdw57b6D3lejEIlIfDsrg61IGrZ1/x9BB2Jdzzwv8aCyX8cobgo
f33IHtam0lb45VLa6MYIsCXqqfoRB9MAjrLL5I+hmzvQIDNt1Vgz4+IuqKDU1rIMgr+OaOzhtGNY
kSzauThTyZ/dlgUkIwcAgcV07KX5X1//gM5nhe56juBR1Twwz2QpZw66gh2yYLXxCLq8z/0mRUsg
n0Ksz93Bf+ozVAERPRBjDGGZiMtBN6o49k7GgrgcnLgUcWsDVuLV4MRStbjKU3wn1p4Db1MP4y4R
EvheO+Es4KZhbfKWgZHrHUq8Inl5TEZtPygvqoeLm5CcNNeIcGoUWSU13nlTtogi/xC9yvDy7oy3
BdeJC/vCNfye+uoLZK/5Es7NGC1jfCkW8e/qW9fRnXVbEI9HAJ6u/xUEDQlys0rxSMpniPtG7Gre
52QDGzFT1qGLRYjyJBv95gP0ueBkuPOZ9hQ94R8ERsBo/M22emDpJkuiAFLYuRd3cVeXgKqzr1FR
loJYsCyeogR1kNorYo1r7I3jTDrlTR5BQzkk96w3Q9z8ag3HNzqsBBCx5c9Fym/NCkiadA7UGINH
NjcorFzHYfZcEe7wlx6JIkf6kcb9jVN2QyY5Fvhz1sgM+wYECtRXRSaLr3fGaBkt8m5XXpe4L4H2
PrOvAJ6wAGWDIe+U/p6GsjDOGfRnCva43ofEavwi/PCu65+8JXgNhDo/qW7jHEFh30gMIEy6s0R/
n5gzCI+MgB+MsnIc8HZT8OBIzIgxS0FjHxWRSxRCaHTOixDPQ8zdJBnUxovYDvZql8woXrYqoiiL
hc7Yymbj6rh3WpguUFmkVyv5bUgj+sRV1nH1KlypWO9DV1RRJ7lsOfUf0hMmMdJBrTbxm3JyEH1E
qBTS8RJWd7QPK4fafn5ZvEoN+7q9ttxFaqKUyI+mc+x4CQXZylAwt7f8U+enZrnnN8qkSP6aPDox
0TVfSDbRqkXWrfWyy8cIn1ILxZ03bSqNnjLxhuUe5tjO3deetE4GnEx++0uWPncbGT33zSB2+rtV
UJA+18txY9k1+rwIeWQqD0wQ9tnmq5tvwwBb4PGZ7oaQ1vuh+G8mbeItGtJ9okRwG4jroMt2+4LW
yi0q5fe5KaU7Ijnf/z0JMllEzoQNRo5ZolBXri8TAEiqcpo0EK+/BVRiYeGrMWq4R3petkL5vbiI
jGXlqS7sqHLKkEkjytFenxScuLn5SbENTi6Qoi0tfgtxtfcDji2YT0gpsUipUIH0piZNd303Or/r
YUK69GmlIpNEfd6T67WNeyQydbrEj6Iv7PqTmOEtHSgW7t/JQeb/8kWmruqpV/VcEO77FYGFKrBv
VuGBoITNteCcyTbzwWgWxqd6O5LkysQJQ39PSph36XjglntfALgSSd9xkkAhZds4UogjI702GHYv
jjV0VsblKhSOUSPx80vgzXnT9mTQ3Le6eerNZZJ/XCa/z2CNE5xftKZy0OaPTLkJAxL1XXbIVGgr
tNTCw2CuudiaDv4DbMcwYQA+CLBZ+OfCrGO3a2W96gAiSNiidczVkEKAj7FZCVkNJ5QOQwZ4hj3l
f+2b85znrD1x0P2nH2WhkQ2bXw1TjLO3FFwWVgeS+YVVqoysH5BESYPMKZqwP5w4ohB1OB8aJEUa
CnVQELkTel6rF4r+Ic6Ho9nZ4QJXJhAo9Wdo0HgVpMQMLuyrb+ARIFz1cWXDaouatIidiWeMMcA5
Qf+4TUarclSvdzhC4EEHHfKNu0RYo5My0SmFVNZM3MExvACTgG4cc3LRS7bM88BSLW9kvcROhZQJ
ZqEr0Pn2r8B0svneU2Uw2Rt2zcrJeqHyxD30kijacwiik7Byttd9DPiPG7y3rWgdk2JixBV+OVDy
sgY4AY3AC/SIoELylzSf0RlgAk+4JkDvk9PYwn4dONsR0TkrxMSe2qM2egU4vXcdaI2sAJiOixa0
CzAVI/3e4rKIiKqN5pF44SU8ywMfoL9OyEz6Z/3JAamFUN/XaeoyBThQV+vnhS9OibI3ledFdZSf
Y6v7MCxFsYq2hrFu3MAqwzbqLSaJdPoRLozVik4hoSDlrOJQaFCHgfHjt4q4yaIcw6YO1ATw3np+
m0UZVwslLAZiMal8omGbztgyAR3IJTDSpW/+IloTQS1tUoZDuU1bvyUzD2a3dNG6WNBOpuG9IBnH
MAouINqxGflhJXpnQ+QzuUDjnkGySLXAqpjUCgQJ0axP3gP+lSoC2qu3Q6BJOQHbXvXAJJEvgI4d
r8Nz+9oqGI4uRvdikn5zY6L/r1tRwLWHqsfktXyA0AWZamFLB5HSar1XLFrAWtumKTZIWI2tCEQ+
6r1sFWTI7Gunj/nPNsUPDcc+YUbFY8ukz6X+/XYZi8sFoV3SQP8h/BSacMEMBS2bvJE1Lg1WkijO
qsG0stK1ye4Su0EGzT/UNc/1VZAoeLzuRtHMhdZI1r9B0qAUemIyJ/NJfA6eUKq9moe4fiKl6P7C
vCaLsYj5dghr4IBajO+cLKZMxScKClxtAHZkHzx8dVCNC1tl4YTBkudHYnrGBu6F/WY+HBnBUhcO
AvPg5bsbSUBPHma4eKC+QiZPjvlk6mgU+dfOrnLT/FSXR3H2u9A9dBPNUmXfPH0DIWG2wXr3UKvD
qzyXPrcH+Xu0LrHaOCuPvPCW0eO28G7Nf6WSmxQcRrVZjDC93Vglyw9jUkRyId+ZTF/OVmXamr6P
Lqcvb0opcbUVegCfRDYzoPcGBQu5Xj9d+dpU1e+Ebtce1vTseEF0ZDAm3C70NYp11bdUQQ8X+4wr
V9FrMR2MCcKC3nDxk+k1VrPL7q6WEVZLqnvtd/x1yBe9KEtKQpDfD7fjlH3qGDMFxsKJFSO8q2fS
Jq983FrbKaj1c+CZfmpjGym5uedfV0AZQo2AFoEb2cq7+d9I3MmTe59IOlnhIUtFtI0TbHxN6KuO
G0B5B6W32VfLiH5AockUe6wp1C2xawB5IchqPAGvITa6IqYYWOknJI608Z9phiFRJeu5pwqdUz9A
5mUij3tnDAQytBLi84vEq4Ag2N9yfY/kMuz5MdWpiGC2/ZWmAFox5uCLlWpvR8I8RP5crflaj5kL
Z550viztaL1FcnaoA/jjcwKOsfkUXK95a6ARmZjNjO135Sj/12yqRrT8VIodt0oVzWcYOa4wM87Y
inaJKgEBQQ79pUUjnz0ur26njsKkA5vBVcbEpyzOvXeHLIfCuUFjYYoJ++wVIRHnguEIONM44/a4
E8hiUrv4I0MxE8jfQQ3CbxDeK5MHtjNz6zFMYbdhEHwnMift7Ioxo2QNYsV9p9GxFZTqeiUqSwfk
VvCIFk2mQIGG1uLi4XgpHNTUkL+SSe98SUwlVxZAfq9Or/VbLM42Teet12yvIZb6N2cFYen3u2rI
7DPpuAmgzNEc7lA7cw+ELLsISSDpxPmBDSXaPIderBq6lBYFNq+MrdhSpZE0l2B54qe0cAmwY3J2
aWs001ZTQ8SPTDdU+uwmXpFOc0yh1CUUeoT2Pqj1NntfH+DZLttdVlDFgltUeSUsln7GOc8XEb+Z
hAfJYC5nDSUhSVj6RjwlpVmEenrE886SP959dNaVe4bWyMhT8MAmj/Vnqn243VthOOb+gIfsrSG8
6iuhKhAzKvbL2iwJ24IHyXQ8p8Mz+z6kBEOzzx6uPYUxHMkkM4BjR1foDQWUBI6xvDdZ1U1iQ/91
2hlyjEEwEFrPeRnxXxc3hUIxmGVbs7zax430LBybPCT/Who8Av+cJ2Kf7jcJBHOHvzyyAB+Z0STe
qdTsnXG1V1/nwuhe8WNLSkWirK/U7+UK7S9uMHp00aA5APO2+nLvWYSCv8Urq0sLQtiie1KGq9oT
niLn7fjHnKj6o8Y2Lc4k4066ojd/YUz72uQriR4e/62biE12AxI5TWsnnvagJES0/eahvpR4scUP
DfwJ22T0WiFPp5dUO47Qk1iTPNkC8QGnsTGv3jzLP7FqcHxmxFpK1o2Fjkhlr2H3A7UmsdNS0CE/
vmhCyZTH0nPikjGGZhZLjwmR3e+OvDf47tW1Oo9J2FtA/gF1gI+tB2BVEMEH1yRm71Pg8h0r6bXY
jvbxFz5cIVKVKXQm2F3zOB5Kd2GBaXKcmjIiYPD1ZwDSfGKWLA67i2LXFRi9XTm5BOd5lrx0q/v1
YQElNl5ovshISMHC/mKus2vfTmI0gSsMXPLiKvhhSKuNeLr+LtqBpxHOhwNzhsLXkAgGyXym0RkP
rHf9qjhB4f+1VArLSNlJu7oSnfdhj5Z6TC1YLRtO15nrYI86r1JLTcmLutiwSeRxlxXpGAbQTBhJ
SNjWW0V77V53evAUMarTUdE2GP7epCqkHFTGYtsGZBepgKPVYodnwZkr+pnxMwhWLIKno16i7DIa
iuaC8ARWUi5T2gTWRh6/PQghKqFPxl3ATgjyLYas3B1qMd5oXdOTUwLxYvtpydaKGpfRKN7m2JC5
20xjZHIPWPf03NEguAcCEWiIe0L5vIj38QS7Jl8GmHbc1MX98/lxrf/05uFrvgHKdVFmz5Bjf0H1
O159AkC8UyqOWi16JM9d7mHShWWsuUBI+0Wq37qobUhotzlD4t+92rMtzg83nrMeStwUUUA/tOSF
ZnsbcgBsJIzQJp/a1tTck42VKN1TR8Bov5ukcOtn7V98TDGHbDXCrsKjpijBHnl31qfKuj0HC03F
7xFJogbvCvTlveAX7SyH2YW0pW7dqhcHP6neQVOLAcwbJLD1Gy629WDk8qDLNroNc4i76vQRqRPu
o5b6LngCWnRhfFopeF/TSfvxNBsBlKMgiRkjz+n+oRudgKXfMVL9T/4AOchFQ5u+ic4/DMYSRBT5
AAzujsAWxl+7vA2yxjuCFEAVtRscPf2VYNrJNBq/cD4gHnaqfSsG4loaX6w7OXKrmDt7D6bph8KV
tlyfq6kZziJdiPiomN4vC1tFDJq7T/8wrLAN/pm0ZjiYTooJSsBL2mqrp+7UAfh6Ti8myPWVL7wP
F0p8W3cjpQGCAoXgN/6YEfz5kiLz/j/SOkWUX0K9vqez1f/pOwVYjJg/1iF6Bbs/Hdf+ehgvZwz4
cqESJUdot/dk71bKeiVSumOGnStwZuk/m2xr3K9pJj1Mfe7hNU06X45fis8Rn0XFJ9V2PdYgbkbf
Lu0GezY4Ve3WGdubM4S4dSL8rv1Ult/WvD1/32ZUR6Q2wlnp+o5FL5vJmqA2Q7053mTxIFZZ+qqv
e+ToQHoDpJqyBpUW5CaZoLXW2AqO74Jheq0NqqnxVfDjKnG0OQH9ECEUXbqku0IpIndhoTQqsDEd
48tjFTCApUY4u1D72z+PYSnOjdHzvA11dUMviKWo9mmlue/kycMunjdbgMrURra7X2U3N4HiVPeo
nOTcLGQvDsmoIjrPjcUY3RTORU6bDTtfP2NW5jyd8NhXg8pUi2Of7hssfMRMxdm+AUat9hwuJqG+
xvP8vsMGGO92N2v1M6dJD8Z5+YFrNaPrkTwTiW0s/fshrV9NQ0ipgwf2bdMkFNF9kL5eXFVr0u98
lBlOkvH4q78Ww6ZijxJjv89oYcI01Qqst3VgWgUBcJgceLIUNSr6TT6heh8R6r+qjx1N+fUZLnRA
p8S/rAeaNAg6V2rMLXQfFEUTjlCtbFczguTCltsPHJHX8m8dgDeXmSMoDgc4d4xs7+jnVkY3BcjY
c7KOhkMI4auDLRgwd8Lgs99IKwAK946VOCl3BNZeVal5ZMaxOUmEIudsS8f6VJgr9wY+nn+t8Dqx
X/vQkWkz3C7VkwYWr6rIJY5NPfDkl0iro2AIT8awyB9lXG04pUpfygDT5TlgN+xI6T9lWypLLvJB
As+0AS1W3sD1X7touTm2hbaSsX9efVj6tNnHhTbOUBNZ6cCVYJ6xvhm0M64qfXB15npZngXbfC6o
+kYI5zvYLoQLDkbiN4eI985XRkCDrDVEy/y4F312ZPIcFxGwWH5QAJxcvGT8IUlD+MK0oGXKtY/1
QJFq7floVDJxJKSDdVN0EB77WqVYIJB8k4z7olo5S0NNuJuA2K7Zk2tSJhzAUKiTjehosoUwN8k/
0lXgA6Pe85AAo/G77xnkYil1HuN04DRDdcGQE2jz+SuXRkTQqHLYhJKp6P9Ro9KLG2XMi04DVDZv
Ra3sZcXTLULVacc5B+74vOGa6tic+K8f2rbJlmOONnQkXZak5hEIcGSNI/fZxcf31VJBgO2XJ3Kq
7hjZvNQyPIw9wrh4AhLwqIg4BndULMRGH/MmJBF7I8zneMxm9MNABpqpNzrJdMJOeMp0BbYrmjKz
s6iJXTk080XbNPFgbzbv4eg+aoQTNT12lrLL5DUcrfuYW5rl3NKnV38XPW+B7Yms519/7xDM9ewT
LS8/zV7zFtw9E0YwnBLLRUOVpyg9qbQ4Y9/8sNkmEX1tBiBYg731oCorXaQHoiZ9XiRRBwbjXvDG
quCrt/ZuYbDbgeyzexFrd+sgJvjWNe04BJlfKFbuxvvsXyAjvFblddu4UcugbLQcFd8pRMA4JJGX
mbWBlXroE8W6dxXNplOi/27LSSOqDJwF3NItt/tGjf4NtEk23HFiSF1iB6V5/LWs5szsPbSdDhOt
R/vnUeUHa1CTB4NN6rrb6ibWOaDRWBUzkYdpo0OYqsrrATGYMy9c6Hn2gSB/yWDQVwU+BNgLKhte
5MSh/wwlyzzlsD+5/4abeecYqxpHSx7Koq9d8qTdfwkCmLAX0BnPam3GkmT3up4vR0zF/CeqEMS1
4dU4EhRcHfpWVVPkskaj/XOQ2L65aRAvHBbgrD6hcafW9fgt5ViyPoJxZNIrBxmhD0C6ilLDx4ea
3BQ3I1F/N1OOZQ13cwby6004VjGoXhVNIKApXnGMF2id3HRPjSZs1GUIwG65iI3g1KCkX/9rEnfJ
/5pZ6b8KRsEqdj3sOrYDH0xc7u4grnecUoAm4BFBKQzkcXu6ZSD4nEY3sTR21/HHQNPVzN6CC/Jx
+bGcizbwg6BedjDTgR0CcWskQDSTMx2UCqhDHAYVB3WX6wMd7p2HaB1+V5FmuEEraCp0BvFknawY
QRXf1LO26NDeFwmSAWti4Feoiu6tplyJ9nbSCQ11g+BRA3nDbJI/Hc3z6t29JW/M3B+iIQWR0pTm
jK9JMPOcOccNkNKSSsBDklo9cCxXu2RRaFqizg0TDhLFixGtSN59fBb19bbnQ/dYDXB6OfPp2R3l
tmcO3gCfwyEPVhrsG8i8Y9B/yQOt6l1STBN7/90mWoM+I7Z5G/7RGPr7IFiQ6b4vDvbjQVNJUyYU
uSSBV8hbC+aiATzJVifb3XQK/XNDzJQajq0Z/mJAb0lq8FXTrnUv1dHoJrvIYPueLyCCAoCyTjYW
6CIttTklxGei2TDH1wnE9isVTGvfjlDNi6A90+b19HEokmFE6ZGmIuLyMv5/d94+0s+W4GOVlzX9
ZMJ0zqOhKvFnshIPm1pB0B/3lVqcr53cgYNPim//WQKTBbt+HQsDk/Fdd4hBbYEd4hYtirOyGEWK
OG12jvsyVimRfV1trebsolMQRSPIfREAeNjdERBnbAAVFCoKf+wTJnbnXlQNxVYxVxDT0HHSJxOo
C3vb/Zca8ZTJSdbD1owde1luIDkhG1vi6uXnWXWFvavRBuLlZTGNDAF6EXgK1lS9LasKql2EirYY
feUru4Mi6TDNsYWnQs/iMcdVF1GD5POeaJWv3fjn48ta/Uh7h7o9PYc2fCzQO5p/s/Q74IPRjU+1
OBQ9zZRAlIKSmtKxE4bCemZvJd6Q0IEuFkRODxoOQQxUX60LVZMim3u2JTL1bKkIzZK/v8DrERNV
PzSjr49Vbf9o2LhMz4S8NUBiTeREUXhgDRjShVuid6HEWNeoEGgM+kxOrMZ5qxFgJslCGRCL3e4i
+UaKjBRemRGHDvC6b8YwDxkUV4f+qm1BJZsqgFY0OivgVIzRTfnB4V5f+Dlgk6gl/b74eoDkvMHY
0ifiy8fK09XZNMPkYMivn9ZcXQ3LeuZqhoM69uJKdOrar/zL//iz+atsB4HqZQiHsT8nxSqnhcCR
M0QPti49Fu8cZdMa+Cv6OA1VBb1DZYnVejTkFTZvO0nl46qOvpuD+uLIQN5m13lHu++UHeV5vWRI
gCTEMiCX8rpyDyvqjzkrlwVGLL846OL4FSDZc57Zvs1zCEAHgBYX3GK4zefWwijTwU6+kWOIWqir
B8ohhiZ63MHf8t2Qd7wFtYf3sZBYWJdmM66Z3RDttloJtQS1bFDQNHp9lCHYds+LgC7YP+gn8zrt
Sw7Ow40bN0RriySUQvwQHmX+prSOL5a3/Trs8RZ2c/14fGiPqlYjXk3UUzNIhzZ1XlO81H+CJk7N
iQgB3ebXbdrhCp86iq6QcQbOb0f1wpae1dqzqpHUVWWsZKTpYgh03TgG06qRsXMMU1MKwbXieUXs
RQWsUaAeGbd5BP14/wLy2MaWSk2mSh0IQr0UghKIvPzJaSVcfenqxAsrvwI8hqmg5a639R0Mqncn
6nt+3oKRRlT8kQ40Ys+l8gYPz5dsF7o1GWM+4ZTYUXoRg4ikrzmmWyo9YEYzz+UYMJCef0pRG78X
iElTS37f489FiC7wOOS+h2kD+kds7z3xVgQ3vjXNZafIlCSgFgOk0voeopRCYEsR6qS/Ncvvazk+
CRg4/VRl2LWo56481Z2JKGqzw+LBOqtGv72Z9kYC97/9tIq7t1j//hMqHUIIKGdGBh60DqkOUwkm
ijVZ0WEj6TzC2HE29bl86MTcL36iI4QuvmgVf5T3ZAZeroFM7hStixUpCW+BzvMtpmtiO5B6Qpa4
nvbe+0RPKgDlS8oQlqNh4t55qpGPokgkXjSv7L/rEDFDZ11dhd/gMOjoiFMaqGjZucG5hfGo5FR9
B39o5VnFOm+cvNC3N/eqOu8Bnqmsfj7vqTfTsny5y4wyfnVlg/bPjxh2TgXcreKxn2HRjZ70jMGv
0AUte2YL/QgwHGGztO8LNMWEe7vPCah20yyJeabwtVs8hb7E739hi+2qoB2B791XzCISLscaDZ3i
1KlDD4+YURA8iYb/tGNB9cDWsRjb8QBN60hCnxqDMHGQ7EEexkrNsb7lvkwk2ErtGYDcLnwd19lN
x9VAwC069Pyb7WtSTp/Xd1ZoUEs/KLMSby4brz0doTZpNEgu7GwYigvRh0xsfzN6Y0sEp2R2Z74j
03/I4qOlj1kXeaPJCjwUvKwcuzLsT0sDVlWvNZOOYPdY9TDIHXPUefYzKZ4bbfFEUprkg9bPwDzj
t2npq94/NavL3XeJev5oX/XdCmH0HJ2LfeOd9DrLHbF960hXYwVMFaXHmFTLecUeGgbchNIG3IRo
4X7XeCeeTJWVTvcKlrrsWrOZ22xXpHqQvmuGDdJqy3Q+NTFOE/NJrESKgL1jCSGIByvfs+PGYX2E
rWW1hue60EKBxxOAJawYNkYTg47q756UMcu2Dx6gs3DWgW+3WA24y5uhULuYsSCDaWnjic++ShsI
R5zHWU003SOSBPPPZyvey1/Ch61SBY8WT3MHr/yyKlsZohrrGMbk2sVwdIIimkTU0FTZSFmMGCHd
lim99mOj/KY4jmUW2kzS/x33ZQOqP05TnKbHRXllZ1zH6Nid5o+aDo9zE4dLoVwBufV3vUi6TmVQ
aLuRik8ZPzdX1VOa/chapHi318p24amfQdzD4a+BN8Sjd327djwkcEq/V1wYFTdZjzMgW9FyZrbc
mT3MGXKk8iMJ9FCviTZ3S08JldVxyOR5ZH77xBlb5KKzLljQKJcEDvBOAPLxfREepJ9FB6NFlp+Q
bKZCX/vnvxd1LNC80YM/8tZuvhWvlg/O0/XGqldpg8Mz/FVVE7bh8VtM1kdVQJzslxnFLT0Jsupj
GoBwwQZugoxhaNBfj1BG3Yb5/a2uSk2b7xUEl46lA1vAS5GoJ1U6l4nDWIaarILN8EBN4F9xG9gn
eEIS1bTHcE1NIGQEPGkilVhSCIvzRCXMSNKF7KgNUcLHyHNvQUY3Dqrsn6qmHDuREF88N0/nhZH1
cLJT1Lxi7rl2Fw5H2Hna1a7qsUjXcLc7ur5hbe7FThVdvRGRXPB9PoSdHK7qC9l53SNfJjCueK+D
WCqyvybAEjD10PJkBsZT0MUhQU0XPHSNIhPreabXyjoH5Z9A4eEzA8PXtXzLIsjHR77LCRsoEt8R
r98IQNy/05C4TsY9cBckvRa9gUdzizlSzNOKzx0GWum1ybkI9O+7Eh3yHEcTqHbK42vJRY0Ojti9
h3vqRfFKjWpIo+Ndcwq1rr8uLhHFrjN20LltVsS5vr/jOnuOOJBSIMwtba0IrZJqLfjTVogRWFXj
umJaIsz6XJkUA1QztzWS5vPTbY1/9gm3XUAGqaJf9nnWuc8gddzCEEQFpaYgOQ9TEm9yx4vI6MYl
XpbaoMM1x/SsB/MyBInOBcmI1U6x4dGduY22+74np23cAdlFhq2Pjej+rhc2200+Dpt6jPxfILUq
AuHK/LG0OEclnDEYE0AXkI/IDPX/kOl8NVppr8dwuleQsr3svbhfIi0SGT/PatQqLz9OPaQNCzRa
q3kqobR2BaEryWK1BCiq8FdySUOTKnsAxOg01QIh1Ku/uaWGEUZEqDE1H+X2Qw2uXfwidC69o90w
c9HwnE+vmLToCb7hBecumL07aVZ1GTq0cyrKMhNpGyHHDBb2645lxqri/F/XYQPOHCq0hDbqcBD0
8sH4WYH0AkorkhmbpfrKek3IfcOT54dazEeNtCQMRhm2JwDIc2Jcuk+S4IZtKDVJwsnUWZCYMIS4
FKOPw6cOmUCrcl6iI6c1154qFoJZ6qpQkV0xOfvvKUJzOk1CR7+ut/6dvRi+fAdtwJqmNLezzYdw
jl4UZoQceOKsp+YBRxH0OsmVb4fB2DM5xN57v/HUmahw9VkbYb2/TAqHBekO54wQ9lOMs5NZNxj7
LYYsVdKHf7sW728++Kxlp+Ie0YzKKajlbg8+W6SRoW3nojUqrTi4GsP36ZvpWNJLH7ZDneKgRIxZ
X3jZvl+Wza9S+cdOg3sYEiIkoZMzPgbab9oBZ8pHmoRz4gNr4Zh0J0WcfaeOlpTjlDGZS+XBoJYC
Pcy23DWSADmfg/owku5tU97nxd0XT+75vGxl0OLgMuIOxDhQHXpr48mqAk/JFW1mK1vjpT0w6Cwq
CizP68OCZr3KkstZHQOtN4qn6l2WNhuCDbdgxkIkBIkZHpHFh7Dqp35bfhque5wKH1CWCsoJgGfp
bSe3FLkQ4NkcyPzIHa89RklYuKlGHsZrLyKMuO/89RmOfB/u227XZSjP7qpr5vqF0yzy2HYF5t+b
hYBKMbYLQOOix9ctcM+fb///TQBNe3mgkeXrLnC098B6w5NDnUko6VhKof3pCEObWx4nfh2yorsl
WbblKrBYGFSe7RIg0zguJWXBo/ACfVzL0gF3zr1cj+XqiiLKmJ4EL+ZnIgQm1wOElZl6bV0aavSL
GME2Y+WBoY2V5X4n/CeS5rAGtF8MUgkmuAmz2i4Ass4KFjWGIB7bQdnzYKEdrH+RhSIvp5LKDzP6
Nd1L4QMMoKRL92dbLx/m0alHhHS6dmrf0tCdrUBDmf2o2aT4H+TghYTXmP7wnZCepUbNNrxn7+Tc
EzPdNevskHgkKDrDbI2QhN96bgw862lYpopucR7PmP+2TxwVpZg66SQ3VhbybKpAZXAYdwjU6pyf
svUEN5kgVs8cAgR/+ctftyWWPJYQfmeewwzRrWzZecvpBfKHCRzYYhHQFB0oCouYG144FBmnFKfI
XKA0yUt/iU8w82quXc5hh5r2bFc+oAJYyDlgZtlQOzroNPSXOPeGieeQWj/xzovgmbTuJwrgW9S1
91jTdIVgJGa4DlSWpa/OIsmAMNBYSLalnrzFkzJ3zBr3ncUd1MCiRxufpmltl1IgBni9j89c4gki
pjVTqmHzCEhDUy1NkLXcmmH4AMHFj97Ijcbe51RSeq8ZgLH3DoHHEpmIbudx9xWonsZQuTXO2kdK
A1+/eDJVr0ERjtW5dALjIDqUlqvPEUuT8cq9HmtCkQU02fiflgpUftz6VXwcOzHHrL2n6q/L5kKo
HWuciILIR2RkIyadbhoBNtnoSerTsUvnV6X2J9MzPNz6qXHRfvLNVwNRJa2vsf3/7ZHtsptfIA0L
0tzsNFgqMOSYeYvRXa612LImshijftNrMGP+vkWtOJIY/Rj8ej5SAPwEhrNwy3F3Zpf37XfLUUYr
DRQmOOKJJrQ2qFMlFsXdzfxhY6uBnzBslp50FmQ3KhiFfuBcIOZAdCwbdqL83OYsyTFMNP3mpRqf
Ru5j3LxlZF56AXqfvMW5poBocLJZk1Ojq0lQcF+yENUKpyJ8+E04zTk5HCN6xoY1JScSEhV9E4NC
vva+U4M6VjPlR1fhBP/fEy4ww9avuTS7wqkzJzymNHXq2eOnLAQ0AEj7iKdeGniVxSYJuonOVqsj
qDlb6c+3vvZlH57KTo5blpgBGN9JBhCLtIhXnVgdUc1/f9As4BiwE78Tqb1n2/RBYftjdWYuAIe7
3HViWYMzfPZCruskPXXveGBZZ0VVsb6G+K4Nrr47Md1ifRbWs+hbe7PUfWxco4+frIq9IjJXXdHg
Q9f6bt+omcRGZfIPhonwLYzbVREqYPX93Z9blUryO8sz/T4HlJeC9DkeicpW4zqv2BCqZDDtxY4J
q77nBvh/HIezCyFyUq3r3Kg66H+LiMq3PzHnoeXVYzRgp3og+hF/N0XSr2s1mYYYaCn2q3HtsZ1t
+2IjOn1TrqK54E5j520hoiWqpTu7QtMISKWTaTDd9TSE67XESd2zOYYf2eNUS+PDv1tv5r68u0i2
sDGWI/GIkA6F6PoDC6zkoPM0+uO5wKomPl0PX7X7p4SfSvS4zYejk868BXgMN1+rzAViD//eJNou
OlYJyNvF7SjgE7GQapiBcy0wYB6JehGG3/EoghTiAcvQU6+4q0lQiKCWbEDzg7YP5uyBSULdM+7B
9HnDvuTcakkfkjNOusmKhqlq9UAYUwSi1U234DtpUPbxwv8RVYf3sO3YJMzPTboQmVMCAylbuP49
0LruyyfN2NAfDE/NyQWIYtEQogjEo1EP6ilXkut9IpHUtC0ZTDMd8rl1b92RfjrYkL60DCqWYxL9
Dcfe6wDJ3TW5FHgFTn0LIMPIlkpEyQNOUJ1R3OPoYLwwgs6LLIvJCjbHnlS3yZ6zTN7Jchk9s/rD
CfRciCZRdI91j4xUXxkwsI2vMDgTCFb87zSsuYrciyoB8qLR/4H8UIW1ozbHVqla0cc27B3BiGoW
kHRLIdrcqEB3QSwyCKFxeBbb9aAgvBUE2OrVvdjWQq8pQdJYLauduKiW9VU513Ii7L7ujqgHOm9X
+cRKR3ZKCqEVP6R0ppbuski02FeZF9o1fWnuQ1SzfSvDAyozWCNTHT1p/p+SltSvn7naebogQIok
ZLLpDfa9b+OlliXQcpKpQ2xE5s8S8OEkJt+lqxjIH9OYnFUJieRfFe4ooH1RmCAIX/WGPK112kGJ
b5wrdo6BWCMdEP9B2DS+McMiCDyjJDlF3jcdo+ikl+hjk6DGszPRrl4QxPClv7soRm06tfe/Vhc0
DGjK5kyoqO2Og/yYNFqItQQDmyNhhfx3R3z5tjPdIJK3tVc3zZZmZ5haOrt/bnmrCnxE9iaD+8bs
AReuQoTC5eQrTzD07JisSaJHiTUOm2+2PXxkWc07Xdjcm04Mp7of4nwiJX+CUwsgbeNxxjb3ZR4v
8h4S3VLy0K2lcB3mMWDuIysCc+S0pZFeePnomAlxoKUBUIC1FUDnQocD0G++3GZJs4esI1GxwIaD
JAiTAX211Xbw7G1kBFnsu8WRR3B7at/gJ+jjTz14UHuI3Vcxgo3dShhjAkJ/vHbof10Rax+C0PFp
aOMmd79Ei6K6e43FRa1WdOs9v7b2crokmFw0u7yOi2t9MV+JXyJAaTvWyDcMoSD7LBQRt2meEmvR
twM7XzynNrI8bQvcPIO04GEoP35eqtV2g1LNeicSiVEqQsOALQVYc6/JMQk4/CF6w4FClViz5C98
U4nHq31MO8/bhGwdhsOn/qqewg4MgrmN7brJ0FmzPWe5bXwcKh6SchmYPow4FFgJimbeP2+MQyge
eQp25WGLH3sQH6KEfKrPVUI0CHr9V1t5rrWCMaFAXiAqhd/FwBerHMWSoO0jWk8Cxi5jZnxJ8ZAe
7D6TjsY+P05SVnVW5twafHy5osSCGg+sW/of8ZQ33dm4Kmz9M1LMtZjz0VsKyMWuOnm7m07CPDri
idMziRMu74eaFdsI097lO6FhfjBc/4jx3PpdEPbO1jhhUPL09Owep7DyXELJxCT21PJLWBM38GN6
i8ALZoXMMB48/7cMCiDA6DqV0tAvFMpCI9OvgiSIfzHWgehAdSCHwx75uQhczZ0+WpsqGbxK3M5V
7wlb4muOhd6gsi6tbi4Vxx7KTnGTmqS7yqfYROPeF6wonP3ai1sBfBpERHmY6xKgHaZnEIc4S/85
ykHVUkh149SiHZ8ylasF5ZLJth+WGgN3mULEz4SKotn+2wP/URNllpKlzId0qcUi7CMUKwSnoMlF
hFrIKUFDLvc3B7SVKI2A9MPZoWx/ccYJdPgEJESAnpDnQ4GNcHO9KLjYOaVwoiKMUfUUE2OP7y1t
iC+bkjCf54ww+1oYZy6wOvRRxxZ37Ushx6ZAwQNWS7fe/LiaJ/alzATGFo51DwuMHNR1DYVVionF
6/RTnC3hpvlRGosE2xjR5cDdwexmxH9soTXDrMfFgxoSXCpLxWQn5ZJ11A2mpe8QFteuPJtBUTpu
e8Yms2EOQJWjgDIJVCo+Qy3Fs282Ldh5ZAj8mV6miYVrpnQlLZOVXBJbo5/zhfUzcAabYYKLh/Hr
6xnVP9AETTMM2iK8Gm6SKEBTCNBHyvPbLSfPsu1mgpx9q0c0pbpAdvQ4MaCfrA43PiU6nAjF1r9u
zMgipVlmQx4NFAwiT7XQnbyV6RE1I+aCvLxTj7SF5XqM1wbY0zbFAK9JI+e9t5mjTEvsJDlHCsv1
7blcZ6eEg+UP6P0da8LzcpzY3pU9Y20+ixcuNDB7YQb0CHmIJzVQW7sNKKltRZA8xm8Bawwtb6Pl
nwqYiZgYs62CKw9tL0nFW5X/0WeXQ2q9W9WhZfL+2Jbe75RUzTLNrE6UXjPUvKPveYATLrvgQ8rM
TGaQPQvN9FG2IyAHSEIw/78lrM8C8SEgWqD5wjqjj9VopV/KJ16Gbnavg78Wd+1NrnrlF8EZ9ETh
xT3LdcvPMat1RuSy8U4kTWpy2ZnkAcXBFxQ9sRHBOlJjFCditaMDBL8xO2ms6H+bVHc2/6wShnhQ
W0hPzHXoNGo5BQ22FOcZFIlWUT/TPCToSGK6P9LVRRN1kajb4lZMJZIQbKehVMBpyXf/vqzcgwo3
6v8jAAX1PrH6+zZLfghjZV/ifdjCc09HivEV1FctjYk0Ps11+cMVEOhB9ybCQI+pCICpc3ryGyua
ruITR3CZbfXd2sAQi3J3rZLmVR5aQoFw1PrG+JGDjCX1ZkkkbpR9n4ONwqPf067se9CxiKb4rWNy
kBrOvydwAb+33852r5168ImmvMGtQrs8RA7pG/x2smKYXMIk4+fi3gx9GZz7AUaymutVJTZsUOTw
ESTSMe0Eqd5eMNN083U+QtdawpzyZbxBycidlAwfTrVBBNNl5iT5klhZW/wpyNtk1AP8xaH4eW4g
jJYshOISGWejz9HXF7iIuZ/68dgNB5AFDYFeuw2UviPxeIAhFrLiwlhsXPyyuXvAEmvC2F7JzrzP
/8IgvOgs6F/mPa4lPRlZygCq2y0ABKo2CzJlYWRr2RBhDZlBIU1+Rgv9xcJYK0EHf6nxhtxADkC8
wVGQw1vgOEB0JW5fkERIcezb24tc4o3zZqL5P7ATRjPFOv9ir6XmfCOhpDaFtsALn4J7vxpKgINa
oOKbIZyMhQkVYLKu1eJyBW9Fl1+a37p7SPG/scyiSkQSUqp7n8Bm7WzyJBpFoJuMwNf79Be1UqXB
nn9YFYhWcTDfU/0LiAd8+PkWhZiBISaxYE0gXWAxY3Tt5lP/FTapcznxaoZTh05Rhyg9aMy4bwG2
BFpHwD7xMyg6/0/+C0mHUIJI8leIWwPDcrh5WeQXYMq7yK3/PgnGNgeWGFfP11fgerajUAf/2g6X
KWDoZDBJRnQ418rtlI3Rss1/hBZXL0D8eF9or2iIxheDkjm6ptSu/v3k3cS1FGZlGb/BnG3qKCQW
3XSvu5V6ANTKxKTvrZWXHAUOfHrstcIwiKj4opw6w/hB08vKEj0pEhBDsFQyxXezYUKO3OuBERAC
+1ST7Az65Fdbfg8MkWRpZECA3TwUKrglwP4UmL4semell9tMXdoQdeVR+Et7t1aH6OPpsxUXYOOk
Hf+g4jmzpeii7vh1Hl2W7mwXFgmAUjVu/S0Tp5WqTdxV3PlzJ+4NXRUVChrZc0lbCS3MULn07maX
7M0jRtTqPij/CmRiMg+r+kFRCoD19WwPZfFAzl06d+s1/Mz7bNmOS4g7YBhbI+ZLLSBE5IBqLHlZ
bKIFiO3/hjWDdwsg+YsLu5LUgnaonpcdPfW+Fyl7NDIfr1qWMr3252t8fl1NNtJ5MH9xsOHTPnHy
fWPI1YLbngl9Zbfg6Sme115oHKh+ofBBSmhTmRvFm/OyvR7IZcyGsomuAFFZQ+iqsZFOw+k5a8FZ
vvtUNZtWQ1DViYlhF97KocoHecmh8LiQFmqnnRywlSnC87FhWKRjWc+3JkBZUWSI8ggepPEEI0rU
JmQzB785unC9BnyI48Rlqist1HVEAPNh57y4odfouFjGOkLRcl4B63yGVOWhrj6Qoc6s+GittW20
P5UfpLBOA4rLRH+hYSQ0gn0Tqw2FbyvRTkN1InYakiQneCe3TZCuiP62Hythwd3k5iU9PX5+1F6x
uzln8aCgnBv7EKJCVKGtKzWLbCEzQMhubqiXhuu4/p+63id2EbDVDlJ4c3bWLL+1G6gYNMx6b3yP
OG56wH32OqsvLGoa3QQKIg28ISMLU09BQCqaBuyMpFqzL6RMEhlPOlhg+5JoLL3lpT/5TMHDQEDO
uKoGPhlJDMbFYOQQMJ82J+s9dbqlrlYpF5yaPSxNR9Ej2nlCU4pM49YYkmU0uQmDshab7c987TFp
nfL1d9htelcwuoS5TfhcIONkvbzsDKkTh2vQiPSxqE1Xk4GmAoaKNyPUI4BfjoGQKL0S08IoXYLy
oSuS2VFgG+eOs9JiTvF9c9/+WAGwf7nl1RJcf0H1324oSv5x+3M7w/b0cQpiNPA0UOYKIF5tgpoO
zDBRmQ2E4JK+xrRRTI044FN0n4u2Gy9ofrvKOSR4GlMNs1dBdFpIMpHoHdp2EQIEYEik2OndInJr
TWBFKZjQlQ1ehSWIMe96Vj6YEkgY4gZtWjoRJYmIdDg0qscvXOLr6a/9z6FiB+srTeb6v0YwqWcU
+5yq5i5z0iRJReNIrZOy3whEQ05sIyHskCdEXcdgEYyuW7FcD/FpHKApsr5U6B3JWOIxEIDKSaqi
SW78GKYz/OIE2NpNdQTiy/dbpll3uoTLNYamCkfQT5HxCTQXjWfncPK2oZCatKgbQqj23/6a9znY
T1omW/I6w96pVYzXPTIRXOraL8BdgtvQ+49poDviCA422xuTLkLpyxVNoho/ESQKAmETPPWrIqlp
xInDLbCRhZbq0DQYRPFn1j6kXG5jtYrVZstMQKKRDAeCfDLqDwWiQX4bfMhflVt57AWNdXVzTU7m
kl2JvLS8fYzXHaoH1ehs+sfAgPCbYQoB1g0KomseUXXOYLMozcv0bRMos8bi5grE8VA954u2wZUZ
2Z/xUbOF+5/SyjMsp/s1jmWrlAj+9AYSsy0Mjgr0CxKENzaTTKZP0trWZoXDQOhgUKaIv4dt0y3z
PHecOC1x6AZ21R0++f+LS4M9pwcwLrPryjQv4mVDBu/py+37Djb6YVO34T9opojdFTiA6gk0FUhl
LpXX/m4cVQyBWgSMeDV73Lk/sbzYikY3kb8HJGlpFXQsbLNJrS+OHQlsM04eX6283KPKNZOjmThD
7U2YlZg60FOltgCBBOh04QAxxIWMQ77nINIYaIJWoovtphxUfrhw/ot7eeWE/kc0KqjYie7TJr6W
WgMxYofUU2tjrUQNfrOHSdoRYYQP9mjxS7fD9YcD74YQAt8UghEIc16RcGD0trrJVMaSpqk2SRkj
h1H136QREoA/tsDCgpgrnu5RnkdrpAb3rig34xf4AQt4iFkcyqgK/jbgWRN/qEyKt8JUjF5l3n+7
7G8JhJfQOupLLr6E40Ko7JtIdUbYyxTPfqAEEM9559Gf/wdy28H/B/7Xnjo2InVXQGg50CVVYX7K
3NWCchf5s660L1dlHKjNF38WpReVHXSylmKyRmoRht+9RTRhbfjWhOAsYOrVSDHXwgZb7do9vamY
CTs8nZMR16FCNYI+pMqkB7q63xul0y+wetOJMISrWF5rbfGkMScsxitOSyvHvTNw7TxAIPCgGd4Y
g0Y07Lyt+lBQxLWzFRi0S2jIkUwLT9XoAYgW7AyRfPzQR64gxLcHSZSSPVu1RjMlI84Ub2L0dBXt
SZR4CJftFXWnKqIEkpVnsbVqPUYoxg6avSFc7S44sew8mxhya3SRVhpiJSRb49M6IFZPxAbxcyNC
s1N9rBJhMVdQKDwN26vrX426dDFS8FGrsaUwYVNOt5lXX5Uso2/xqlQbZqYn/uPTzhQTqCNEYnaL
8pfYNiY1K3TwPWGQjk1yC5U6ghr+wTlID/g0qe5BGvBLTseOOJA4jk7Cv52LuXgZdFLETgNfiFz/
HhB+eUlpFQgctQqTa2dmpZmfpm4K1Z7VamsZ8SeYqICnx75V1lVlX7hVAlAS48Y6iokD3BJbscLX
aNzx0lKwoy6PcxWrbIqeWilbWNtM0nlM66skiuXXf6oqcOBBxru/GtkJgyrO6TOPKH7kZD49cjJ5
DUVnYKIxgAiOae/U9xGtvdg4KxKCwJpl2/3F77hBiehBflRkhOhC3Yhd3t5mHZZBaF69nB5VlXht
8s5/VjKAK5LK8GnUlCbwUQMrqwN8md/6Zq4JXZpGRB6g5eq/LjPxUZ5ZLQwVMsynmR77fibfLwnQ
8//TqBhCElWDTqqn8n5GfARvVj3zRh3YbRRM2Quv79YsFT6SihN8k86GMROgEupc3AfZslqMwpJY
VfLcGfFgLw+a+wPus6OKg/m1/6B9z4BtYSNrbBpmlpQts0jJlERC7vZ8YphQjhq/ccMGTkUZyT1c
GtT4UL/NEsaNZGGOgUfjjapDANx9tk8sDgLYufgup1vbX4lPrlqj5xheXnorP4HywF6SjLriFlwL
fWbIVl+9TgHPCxqfbymFajftIM5QCwXAJNLqpPnSBpJ+YTHjCCALmFj4PfKfeQfxq/tzr5KT+Zji
8XaCHedODaCaFO7MHDRSduxskBzVYqnb5zifGr9RsWKGRKx4CYTeAfnFnsFUO2EFZpZNp9upy9vh
466is/ipRN1QfhQcgyQUncvjx3tYgTSmAqHQPJ99huxVNIs/NaR9AVXFEgRpP3jxIm/vOYj8gpG/
MEltnTYs7JoCZI/24kq0XAIdabPjZEuhrf4XIllSuoMlSw+0egv8+0d1sYukSlbY2Wfn954hxGOv
h9IrFUgfxqCRUsMAo3jb96yECfv81hHKxL3Q3iTV8QgSnuIaQtW7ioyWlEOFrzQE3HMxrXLZ21/k
w95G0zq89MR+FlO16jdXkfIkj+SaSse/VUO4bdSfsc/wsHekFkScQJFlgjaYHSbiMcvyiW2xu4UI
LMbetxynQeTI30NxlOFkv2QLCZTohg8mpUyEg+MxObG99xpl7dwCIhlbRI2n/4mUE+0luA+FWPnB
e9vzR7cC5B6SCdzTt6YNrcf/ZiH/pYXe1yHhY34SA1RICdGheUZe34yPAr8oVKs8m11Be4yA/JPh
oqljK+GDwyu5M1pq8aTf6m4i/2wp62STz+eyJsBlsz8/XiM9PaPojLFdd4vJwbA0dPpO+Jvm+q3p
FbxNsbARsQbsvpOdf2dw+Cw+szs75ISNmOBeVAmAs/M0k+PjeWoPz5EbVfMoXUVpXf3j7i59PTWi
qFIculdq/Om3SP/plYISQdgiFxNsouxZTDdyl0cN4KiRKq1Gh+ZZ/Qm32KkOrUMDq8vjoQomtzi1
qTskw15nL7wPJn/jcctC4JPlS6aW/5ZMRh6RAW82IybAED7CMAOFhDkKkkTNudSM/isrevmHo03c
NcKsVSk+ielz7gNiKJj/qjpsKSYKjHlpqpMIZsf99Zi6AoMyOkzr6NH06GOE/ZHTOtcJdc41zmap
TwS+n4iWCfYzNcKTmjzE3F11jausq6dKeCXAUv+fmA3Wdg104uFmpXq7AqpnRfHE3A/ff8dO35LO
eobg247dhb6A0AJzA9IYzSaFF8MzQ8P5BvekVhSr4e7gMAd2m09oq1JFDj0SOBcwe0W3ZSUzxBVr
zx8qIVnw7GnVASSCbIl8S3HoIwacUb4nDFWaCI7nS3/hiuYNZQtfR+inm6KsKbTw+zsmGcXu7Zn9
cUfYd9CBq5lfJ0CHV+yI1E5GkEvhhj6lQY3FTMSuMy3A4J2w/+1jiY2ymp8RBtgIieXokyGG+A5u
1SfSEZODPCo7kJwo8oytTIgBySS2bDjf91wTbKraUcu6To1HwCVSX098xkyYBBZHJo+Fk92I7zdB
pP6I87JQFuQ8xqoOsQEOAwjDOyvKaDi0BAyui8bP5jUFglEas5KVOqdwDzzB/8csqCzyx9SSxSHg
norSS6ccw2uZztIG0Y1PSavfdLeVbB5kcgx5R9f2Sz7iSR5iKTsdD6oAHIg4SDH5JwbqBaySxhT3
bfGpDe3fgERHdwLWqxzf2YlUn6FsfZCcBYJJrujSBRylMvMG3BlQluXVAUKBTPMOa2RQSuVGzJhu
/LMyeJimwGnvY0D3DEynjc/vfO1Uc8muedY/w/uujt4fYnty43w3b/hzIdx4QD0jSTKW+3xebnvu
w/TMw5KrvQc+GMbPoQGGIleoYraROejDya5WEp4djIrmGZe7VT78CbkYKUIyw0fQWVT78wCSfGpa
T55F1pC1CBosxxutT8zp1mDl56vo+F6dp4VnHV82nJq+Ve1vTCtTXUlsH/go0DN4ZUM6/+mT5S5K
P+TRWpeQZ4xs4lXCFXYpD5C3HLSIy1eSiO1EKFBE9r8Ex90f2F1UMjkFaRmGWdb+xGYvYyU+gQ8h
TsoR2eXTtPN9d40M7Rh4VYUFKVi867zrnEMBfA9oVMeEB5uFHwpo+1ZqNyM/LMeMwd5bQY4BdTqB
mURyKjhvRm81Rm7cBwG/qWRJiQI21PCPtTnuYm6daLsIN+fQRd7Zj+Lq1vtGNtH/B7zJluQVwsy4
4EXHEkQQKyB7FklxLYWThqI11oum475CJQm6uJkTKfzpKQzYHSrLkqyaFSCXRLRPlkOr3LI1tEi9
pN7ZUuMTyA0m61ynE4S3DL9NX0Aw1OXpZvOxdFq4I52BDjowqh0ZGjQOr7Km48dwvf4l68D/PPC3
4qbEsa7y0taWRaBVAJDog+B7Qd9c1z7vRielAaJIE7vEa6MJhHhU0ZbEuF87AwQkvw0GcqSUAw/S
W9hOM9A6DlBsBfkW5mgp52OcF7t50zf/SZ74jrBeEy+Aww3FKoPdc4Bdijrz0KtM+HEjtYp2G4Qk
3ADsPK4zAzaixHxQrKQO6v6kCvWeAJzm+fcEXaixG/JuUzbMvyZJsYxKIp6eel6LwP6ys8TFKKCQ
Gb5538LlPbVbE99GYUmqiYLXm0gMTtreqIhhvVyNBrB1DSZmrlxG8QaQTv/aERP0SZMLSkHA3IUJ
KaUlfgKDtuu1r5byoxt5qSobbOOs9iB/3N1XY8s7ZfzD4egC/1ARF3MEuIsJjLEiDcIPFUlPQ44W
iu5q+pWsLkLUTnbej9ZGjT19TCWFTK+oKIMaJ8ZGyloZTrU3UOdUVruRoTlHZlW/zu/1AEiTe6Rb
E9g0UOFs9BoBb/NdC1rLIPfWbdGnx0UWQRXcRrNaiR/LDzAaEASoCmlwMFIQ/FMOnlzt+wBBtWBw
+0xzo9aNQ5U2FQ+h0Q15PJ4DdU1Md83dVyEFW/mac/QH5ZVX2TfxIWIEhZS6b7YdDmVkUC132O7h
cJcae9Auclqij4QT5xofCiKb+mBo7ZXsrhUhY2rvg2tmTYrLhc2g3ELm0tCBrkgzv6mHGN9n3CJD
dth9ee9sL/D2cVJhDVx2E6SF+5uHKUCfJSR7Zx5gtoHR68uZqrm12MIh4I7vre5J7VQVJ4SIr684
RD/vW3eUHkDPBd31wFgYDlAnOrmjQxHbxmSqgpgTFRrk2cFDfwwbnJd3BN0gKD2v7O1Wfq+AmYd0
5WT8XTk/aNoRQBF5aXszKnWysujRjJu7/yr2NIDVVGXL58k4HeZ/VZIlZer9aigKwLs3xFbC79/X
p2DO//o/OytX3ddQX+3Kdx7OyX1O0/XMN5JGMsVveIyF96m3uvyyjhw9tdn4xbpVU09UUqcRbks2
rMW1LUeDv6pd3XXCvukQbWf/bYmgOZAqa2ydu/wGc4DcMRxDVLg6uDE5o5X0CmPJ6ujrFilCUTrs
kp1AwQNmNc32Wskkp705K7KfnqbDcbp+c0WHvAGeMhJlywMZjJEkhMW6OXodVnz5k0VzVHjghOKn
0VF2MuUjy6HudO05f40D5kimU3yiR0g8YOsPnLImibE3ENkTgggGt7SSJNm1mjWUMCs01P0+FPir
Si7m/FlaAzmua+mi20XUXKRFKYxDiGAiO3mvxU6LkBYvCeH/hxICASXJbKDmJm1ASLOZtoeixj3k
9hz2QA/QVW80Jd9SuiMSzpQ8FaP9lbFnbmMN3KcsL3q9EyKXxPjK0CqlCJB3p1lqdflLw22kGhL7
UbejXM4C8cG0udSTYAuCzbiHglPwU8jqyt46ts5+tUql5tO/pfI56LF12cF0r90yURCm3iQ8Ec4C
cGNvhXRdoeUPTu/9yiYZS3wKMgfQNPdQNJbdOEETHFMWPO4jaUvBi2WGZ4aEB5HYend2/NAkqxse
l6XQhByRutEidR0vSXrOPbLwip7Qtfu3/J1qocL6De7ahlvkgOHgnnJ9STWW0r7yAo0rckmL25Dw
QGcrU2PS3zVnd3B3ELV+KGU36vajdggMD7/LVi/OMSbpLDM9z0x53JcHZpSGxCUM6GZGHBfm2xeT
Rv7t2u2lbKitgG57cdaHS36q+aF7nbiPtDEPNFPb9tVmDhZQLP+P27CT9tOk/KGVtr3kALJNgayJ
SRQlURra4e225Qj392DEoG6lF/qcYISn7YVV0yOqvjt+2IBgCVbhPyr0vkmmFpJ0E8eOtwSwgxBW
Uki2WjcaWADgb+PqdnFPBFpOnDLs3G2GVZ0Po2tmYx4V9nEOLPvSndBSx899v8uqyv+cEjcKIEkP
GpUt6/NsQ2OoV5WjXK/AhyLdrpA8IckdEDU1VLR30JnPq1YRFrPz+3rL82bCDKUjzoHVtdo/W22W
NRWUyMm7ZaSMc8TDB7t3q/NLgxoDnLqSTMXnNAzWvqmm01pZdskqIL1OjhbLT1R/VmKVYyn0t1Xo
QIoV0fHVbjOH2JI6MIzSSrZ910ZpymH6m0D+102p73GE3mnLEWaqewpRFUr575NItcBtWvsmaqD2
s7SSef7AxhcQrr+Hiwr3L2B9gj94IwARWazkNIuHcGoC0smEav++eA5a1VAvP2cPJnZKOLLUM5WY
SZ8CxEvBWZXsaaA1vl/3KbEZ+GR1W2o5LCuDCH9U404TRm7aAdu+K3M17QCc3gqmJf3HfUkpIYHi
o46gcvCk2NoNMflmmebDA655uKhDJa0YFkJAOpRGhn/JcpKTfM9HfrqjrMgV5oZb5WSjPT/MU1pK
5Xj+tPvkenISCvNfv1F7gf8l5h9SkrY+Al1uF4C1wiTOlHwyZZ/Xc14QPOy0vT2epafVJvfjVZDD
YN8r3t6s1DkPYeYPRAyx9jOoSC3Ic7ZCsUBKieF0fq7pIbLvdV1juFbihm4s+zMH2BudLIHRLO4C
fYXVCyfC5XkzIt2gYmAPQq4PiXTnKhdf/wH+pBsdjTPkcxwiYfcZ/lTJZcfxE4JExS29DfPCQOa4
+UGfAyucTqztbDIPzqTAECFlHDBPXWEIFWda6F/aiCVK4cUwcsdiuHLSmLI//4AmY5ZVcfxo1fyL
Sua1dX396kk69xWlW/YKiimcn+WWsuSqTTA1d/AyHhfcvA7pgeWiHmxbMSRnXlZnVU2WPfUNYoFU
SBABn6nj7dqZvjA7jOFiOOdBLqOgqnvP4UlOpQ630HDixgrWr21kkANlG1fmXR2aKPHdp9OvCSMz
FcnlAHpo7PH9xw4mrwjbRcWP+SsxlaSWoEXuHXnWUA8g6Au1NjTU7FBjbvANFHnH3BS5cZIquHwS
w78j43fYHIp5kdTSxvz+e5bVxvAVPTzb98Km31tUDBWU9N88fYVfPjVReBZTVy0BC6k9Y1BnSLrf
Ej5weRHHtCBbR7+n0YsNhLn4qWPrlz3n3YULMPi6c30K0XcMFquFgHQrrH4sSofu9QRW6gwKwUWf
Jj7s1L/Q6gxen7hfQWOjFm19G8KLubMMJS7Il2KcWjB5J1jKQzS3/kvbMxSNI3YQc8NJBdJIu4G/
sYA9RoN6OCpmW1sDFKqzJXQbIWTPPYJTgZMtQ0vDpN16yDNpU+aGSx/Wlrno9mb7UvmbEqw9fWuO
0XgWIyLdAwemZJ+FBYnyR3xHKiFS0GrSd2khZKGl+2gSnwERQFpY8Hovszj1kaiJt/49O2Ug16/u
GT27gq63kkqokNCt3S7J08/RtMNns25QMlO217AzO7OsOO1OPxAsQ8tGwQ+1xP1cQ5Oz+Q5+jvT8
b2IOusT8P9glfKI2YdRavzOF6QQWI4oHLjDfEzMK1zNcXw0+mheHHpHge9zqQrdub6Oh1GWaxgSL
KrAoq9jp0aAyczkv/ovfjmNArLi6IdK+8wt1jEJ1q39Iqp8T65ax3zuNMEeEXRUiMfUN7aP+MO8Q
prdTxPtr/fCS3ePjZir3VbJPsabFtvzy2+m1BTxEKpmvfX9bp15f91hLhethhFHUszyfWPmIf8Mv
zkgVcgW/VtQMiPmK+QQMQA6BJdmuBFdS3v5jSP56fJ/iLnND9ZrTIK2eLEf57k7cI+5DWTGDSWNl
7sctnEZAgWED5PeeZ1ubXIyr9dgOkp6IQMXR/v6y3mBPs4+os2N+bvA2H3CPA9rHO9XLqh5mRLiL
RrP/SwBYrVl4XBLsWKQpU4PEgGvc0mGjeeCgULYagvjEmcCjF7Qr1L1GOKeoBqyO8wx9axpWjXA/
ldubXLPpa/YIIVWKjEFIj81Ueqyyjfn+O0MzlbaBGz7pCKQd2oNpp+YrB6grye0pdtTyEl//lrgH
NhoZE8ez9AqK8gqX0G++k9Y48nlD1NLHwdolTWII/exO4RnKgib9taILDxmYBYnCNXWWewrIOc9n
W26PG3WQWd25cE+QEFTn9419qgrTM5UhSGeljvCUDX6NkLb4bi+JH8T4DcjYe6w2NiEP/DqQwSJl
EzfXkn0mbHLdkpw/fGOVqoYvLBuNjTnjdvb7aXkhlkzDkbrZ2w1S2EMxEfQTMPYugumITg5frSZz
v1kTs7onLaVhFo5HaBlkNb3JepbS+/9b7GSiiMLlDtsDnMI77Fbt88Cwajxx3BzMPJ+ZbL3MvHoa
O2yXRQkFJC4hZZ4K61BEQ8Z9NTVjbg9M6NFJIjpjs11OSRZtbGmhDAwAzI1zfCkdajIxtPGqr9n6
rTuS3JqKswOiGSfuQhbL5RiHEKZacJYjYZLklDKYllFegdrrdFnPR7ogIGVJ/MIgtyi/FQ0R06R7
WUmj5OQM/p4yHX9I8FGxygnDFTPWYOjSimyghSzK20Nkuvz6oQuUcAG6fxMwgw1gzUJ2/tVdaJaa
aeN5rXdxdgU3Coa6Hf4yxmmf81V2Ls15jbdh6bJEd5bfeMQ7l0QEA4E9iPJWjgPLcFMJf7CiHf9l
uWOdCmxj/UbsHQgNsW8pxClqVpRyWZxN02yVwrhhIqLAzafSDDZsExDn1PkphuNZ456k8zlQ3vvy
tA+O+dlw2O9lHMVoD3tNiKC6g2kS3KJR3Kp8DUmze8diGdkNIrBS5tXvd4VEq8BlzueHFuQ8C9bM
NxOLcmxhivFKN1MzSmUmUg9x/u2pQM//GEXTQs/qI6OvgYxytH97Agl2WN5Xzoht+WuuCFwWi9H7
/GVuMqgoABSO8zEh8L9Rs42MCnXwG4Dat3wtojSIGrTu2KbbHk+N2DaL1W+sHmXqnb7UZpBbe+Ox
ZH3wbdtLv4aslTMefxsTOpBVt0XKNGNin6d5mvVcq3Bitgsnadt0ijgLjAvzDLbDofK6b670dv2e
6KpvMEOguJmSiAvSKSv2/PwDXijIbQlNg3s3NqgouSKJ3RjHrEpS8iUMVDsZ9qx6XK3yHh0rc/Ug
ASfCeRg56HNMMAlT4JZzWHZxBMTKcinjjp81tojrPSwaWELannCMmEKBGNY2hhbE+Ped3lUzC/nA
Ms2UMLsJi7uoRTG1A8+u1QAWqkiSIgA/ZFzzCIGQGMcFQ8Dwu3ot5Rn1gg1ZwJ5dNuyhpSZLHfAK
B9W23yOk6KJriVx2kE4Cao6cSrAdLfDZN6fHT4VlVMPciGNmmUloJXBg1uSE969EG1zom5NjIHu6
Di8jO3mOHhjyU6qQjvG7ogbB+euYPRwcOWfQb/v6IMLVsYhG9gEPQz+1uSPSFBQUXgF/e+wyR3wh
eLleZKXq4BlFx2IPrGvbcGdUOTamBHLsyI8S5tCRAcx872SaztSZ96h7UlqxpqDHiqmnAERwf8gt
dAU0yvPftXMQsGVhB+iss4nEWycbGchRiH9Zi3vX3JlGqiOIQXpJJ1LoZyXTNa0knoJt4Y8cQ7on
YoHp4Vwo8jSrFxoVo1V8hWg15oGJXs9wvtdGbWj58LHNXjyuvyL1eM/sjLiyQcnUCGYapYWouYM2
e5CopS391gLrAJ6PTHU4rT+AgIVemkM1hGXoE+t4FmFGt33t//U9B7zRwgaS37CT5jzPzWlrbOU/
x/npga7/Z9JgfRDel/gO6IWl0iJ3utuAFXh8UOGm+Y1aedUme5W5rNs9EXOecZExMF2S68PSfqZ8
5flL+NEfPTzuF5YPBzDl7FOeL6EEjk/Np8sQkFKPCelpAVQP67u7uJZ+eStYAjykcUY0G2jdQB7x
Y3OajNe93Ifomfawp17iwwfityf4ZH+G1xdgcQNl2LdAX+aTr0KnLlz+LUI8LiyMcw5K4m6daevz
dF3hz4oZU+vkITxKWmDH2hsTIQ/vJcw4v06zbpFQGoKZRacMaykK7qEW8w089BR2vASgfZ0Tw93y
Z4VzWEMCt/2BReA7mXs9t2uupKh88nafhuj9Vr+ekXD4a27owGWDHozeYKBSO6SVtcdaMgqkiqw8
s216ltK7oXV39E9+d/2oMN4udFBV4T/BtTzjlxgWQgejAq3uMwESoyCaulcUEja5u/PvCW/61cHB
1hZoVgfjr5cYuwS2EexZF1D7eqZVLK5eV8LR/p1h00BFJmcJMLvEJAKSRKFG9yRPPoLSaDxwtAEm
kJXM7m3IgfidqWtml4OCiIgFRweXHs2re7q3mpue3rrmcUksWZuXVJ8vR3s0oPEHWafmh0P/XNeX
s2K+zO8tmU8WICooj3niBoVBFAP+EfRCoDXJWkNahCNW2xiK/xn5X5qyB+GKEkEcDsN9nIkTq7oU
ZPBuk5GHfOxNrpgv03QOMBTseYFnjqcYO0oWCxiY+4an5Cc8w2rUnk7roKr//R2G/6tZohqjeW1Z
XPrB2oEDiUo0XZPv6+hp47IqtRO/9F8qkemK+dR+bU6Ms433wMJJ619Ga6AfBuCW0eh2R4sEX5+a
oGquOnRUE64RU0KN9sW5+gjkLGNUqYzpzn19Jfw1ULN2mrVeM8nRmNdZar/bHxIeRFvQOqTfDbmA
YREz94VN5KA9ugmwCAYEpGQMhCC/zFsIN64GeglfdLA+FZAkeLCGa0muVFCJvLU+orwGBT/qhFsa
uYETHs9/gILy0u4YRu+c0RykhjOda+r0NgQJVpB6GX21LwERMypH6SK/Ko22zpqjA8pyoxjzJCS6
eiBZK8mi/+UaDdPjZlHtJlNILJJUytUXb5VtbLTUYtZIfbmnvqhGy6ctgkgXaCmlOpI66AibdTqc
ZPo9k/tU0iI7McQI5V0G6k6FV62KpGvoY7Lzer97Bx/u7SEmNBb5IOrEyVuLwBFw+oJCFFkva3HU
1upMCYpLFVsRwpYYaQxiyWviqbBhJiREcss6A0Rngu5wnclrHqR7OKCQGEjZVkXDAJrX2BijE5c0
G1clEhNrKrQGeB8ukbo2xtos36hINuXYI02e9tmsAGDM3woOMbTq3tRswMR90fESR5g7P61UxSvZ
eD4mcDtXe/zzsyACoAlyl1qakupfS4KHk8D+gkxL9L3bLR9sivbd0g53ugS+ywO+4a36EpE3blM9
+9oUwZ9SUezS06gQEdh4kvqxGrAo/L7elubat95fFb9GKBeuKqXpeNOw+HhKI+2keNt8nvOCiY8L
Mf9n3eNp8BBukTSYuGwZm1EviwSKH2BwkK2xFJenpTIHpdVVoA9GHftBZMUcqAolc64XRPvyHh2X
ATCVy6rGfmfSm9WVW6Ml7r6hKSSYUXCnoywId2oIHhKqMK3iQlOpefm8JYWibetuUQzAFJ/mSr+5
qquG19+rojipXvcdv2rlPAQbvaYALgEHnpIc1gu0DbA2d+0FYT6zg8dxfA88Qk5CaWtCLMPNGa2i
ZD0uPzn+YsqixBRbVQUEXUphfMLFZ/Z0megxKWQL/Z1ZlratysKWpvgBe3vQMpJOGaooDtQYRReq
rqpaSz0bVG0ieQkiB6p2uWtdzpVtri5rNNljRoRIndH9tleE57/QbBU25QBQ0ekTUvHqNj9jQrj6
yj7wgoEp/3LdVsNhjjsys5q1LKE9YfXXFpI6sREEY27EYoh0YxJl1gfmopvyGV+DDggWx/so8AAA
yX8rBvInsiTZzpIyuWMyRusETvhP5H0/5SYGDMZ6mirmBw2Azg8yw7UW27csUXVjLmAv3vgkpSjP
FH4JjsDwa2t/e0NOgX2KsmSvPtdXOqMB+CGecLFMn1TRzS5m9FTd3BlEVuafpZXsC8TxX32Tia5g
lfK6CCspPMwCNse0dsnKypbqHJ+pDGkcMTjYVLNAThKdTpBJBktZLymli/j6Sz04EwxEt31R9rxp
njmeeDj/X1K+3fyIGlUOexv5jqUkdT084yzk1EE/ExJruSrwdnWb1gwOx+iGOWiHNhztGIYt4LDB
oimX62DvnfypmsbA5DXe7pklCvAW/ivCnze9vLt+jlKKlnkc2TVtq6khK7xTuIG7pbTfuNmNLH2n
s7giocHLe75mcr6l9gd4hsZMKYVFQ8YGJlWiv0JPX0M/az620JwEYCIRPIW4PoTj4QH5PsMGgePx
nekneC3DJCrUhwxVifsjSNb+M4eiL+tann7lxNTHHZq7NglH065Ev0itcIxpYuRm/J45L5488vq4
rdz8yUMtKpxK19IzkvLk/K7CkVsrNOZq5jeYblK2jxJmDZ4S3BjNk30ZTUHzcoi8Bt8mBZ5c2l7D
fc6XWVkbDVVe/uS6gzBdN6huL3pwpcE3XFGOLC8A7igmZEzhJDRaPyshIL01mr8fb9vn5GZ+Rpxh
88zF0EmpUypnKJdXuWEWbfYXq0T7Uj+7MJDXxedfzwxQa3rcAwIP8T9q4W5BwRWeZRvWI/u7kAxE
X3fY0Ip3PJsLG89W7K7Xh+WsBQYAj4a3ORMbMwjajQqJ6o0wjfxeX6ZI0cg80jo2j1pG0BlzkBhv
pUGLEZqRHypfnRSpWl3XxQNtkTw3c7vNpbQcrqLbjbnb7l/AAEvitEs21cuqMJTJtFcbqc/y1zeI
n9Qq84YiibKvvn6lLk3UQvZBJ+BaICO0Wq0gIIbFuuDTPd72L5v3/JHvjebe3u27FNKG8omrcHaS
ZpgZDvkkX7xcWxwWydab8RkFTWJXWrO00btA8jYzEmO/xrwvzmrr2ccgAALyU39i0IOfuWQqbfEo
3ccfBGSghhaX9T9igvMHstchQGbpfUf9EsApWnmmlHgodHAmHW4hZq6sc2pWLgLFPU4GRspBbL41
zPa5W7dkapgn1tmWfPfNp3uqZZSKvFBJ7PIbUSAjlnEmQcYjbjD9V0QQwvwdCAo8zp/jLUvAMc1m
yL1sitlnBRRInvB6x5B5gCvqJ6G1lEMW5bJq08L2L8UIeWJOGNMJHfKbW7luu2GPJtKu/qlAVPzi
QmGcEQ252bUAipINgyF4rP+vh1F0dxlYjzFag6CipE9IIviRDlTOeDxQf2dM8fLVqTlzHYV1kl8f
PMpZpwbZXl/QoR00nXWVCnsiFi9Wxl+T4zxqNz0wnUIxOQSJ9y0u1+++dBCF45S1q7tixILoutGD
PxWygpv64cBxUMUFfXx58+bYAjAfTStEP1V+zC/Y+bTE2nAP+ob8yg7fzBjVkzGuwxJaFU3qmUPF
kKSbAtf1pGuCU+6M4kobUCeRcKrszbCNb0FtGrs6GLoNuCUCU0xS9DTlL1KKm/zUg5gUmE9+0gNz
8m63IhFOjnT8KzMze5MDYYe8FChuQcntM3bESxDBm8rIRpwZLK8w0GJ6mnedpkeIhbEBWff7EPoT
7UUIOUPkW4uFfhcdjUqcyIbz/EQhbL/pqQ7wh6GNHVxqii0YTZkVjhjQqqKMjn33KjdynEeoRTMV
x+NLmU1Pvst9Yxfv8M65zXp9C5pEDsHZzZbnNGzWGZEyZClVRWf4JGiP0mS/VNzbKyR7Yajmg2ku
gBjEnOgoV27tY9oiN2Fiqf6lvUOzZGQKdj6pXPeDjH/cQaJNILPee6pzVDhlw/UmGetKDqRVPxiz
44eVaqZ/ZqjBWFpvlIbDormJfe5X/z+56/nOIVO0LCrGXZYaPCwV9ZFbbfqoWGgj+SOSgKDV2I/e
vQ7CMEPzmu54s5Elq5lvDxT5fu2i+tUmKV4WKNDl/fw9WmXByIHVUFTK5KEj0lavAQ+gQVyYCFvQ
ZvTfaS26Z/PzFpcmVAXEC50J7l+YKwtBGsYkXt1JyVd3LkJpKoT8PSbFUkunZcvfEBV8gDPFUfdY
5eJAjLBo2JFdgwGyt5LLsCS8Hw2pYaaCwlP8ckT1tfq1y1dgktUmafr8rurJ+7BBI2mlsz7wTa7d
Y7LHclNzMq228X8xARj8WdHEdB26CowDN27U/vT9as6bJo90oSvsWB2Vsz+hbZOWMA789247ddiX
A0S4lUza4UWGt+kWwwSWVozi4vMlFTeUvGZsvYGMosmJ+GSJ8mApa8UnG7u5vIYhj6EMjbCEfSo+
ECZF+Lsk+oUsvzST41YbRRpY3Z3+vcdUBovXFcVGhS78uwnyvpylv41sxyzthgLBXPEWzE9YPSgc
UGLskDR9w60wYMHseO9d7Qkr9YY52L8fJpN0vqGOCFEYFlLrU8dY7HkbI7SKDGkBNapcG+16hnyj
3Xclg7xEW1tIbH7xzBqcLrMvS2xD8JAKQS3YQUFGEUh10VX2FE1Q7Ds5rayRnEGiR9qMlU8wOd6P
NIVT4kYiCU6y+2UeTNyKY06tdepv6xgIyQuIqZFHHrLaEXYWt6/hzaWazQ2y4x4E1x1sH9UKFXKr
7Gu4tE8eS9AsrenWJmlZeFkWOIMOa0Iq+tlNHcNcyV2p3asKDIp2zqfph/XV4p4ma0Ti7FRBKf6n
9ZM0Ql3s1VGBaFLEaOKd/bewNXMmokl2Tt6GZR1jIsO+s+0eWThrd6hSoIb7VJIBbV85N1y5YEoX
vWNm+BPtq+jWLa0A3MjqCuKDGb7S+Dvj9NlbxS2705ellzKCNhygZqoRbnm5VuqyiRTgn5C72HWk
h6K2mi+9DydYu0MjKaV8ygmHEfoQHBoEdhN3iCtCEiISztGNxnW2uiQ3sr03/IgzigOu5DLyQre8
/j+ZhrH0y4rCp8NHvYgLyiAe/uW1YbGqkPHFOC11wBuFgO16Ka1t1lH+OWn6KM8VmIsoubiUoZGg
XUImYCq6yPEGMPKgg4wBraZ8Myso+qiB/JWm+fqTINJ68qM4mozBe3cLtD1uQORX3C8n1WIKmWKs
GZ3v9isUALoqpC4twuG6Q83MoWfMZOpqLJ++Fd+K/hVUiyI9usuqaewRUmOab6nZMH2iQiUbHDlj
ZoGcreDVNJS0cC0njWVDERkddXDsq+Iqdr2tMXmypQmoYNfW2vzZoqqn6oC/TToqQUbxFnszmxbE
46k2vWV4ZYd9fMJ7MupazaI5XXHvVmtED4QPsqUFT6hI6laMC6mBU8B/0I2fqN6XDmh8hhS/qj7Z
+yEH6V0+A/A5yNZP143Fcs5AyVmRiyXudIzsQ6dJsDQOGnkm/0BWCEaDPIwZNi2u06pdOF+QHcUz
hzFv3HdkoH8A2VLwcnUGRggBGono3G7jI/QPhu2L9qUMyl/3ahQn06k0/pn+ApTss+47jKXi6R21
H19BtIR1cM1GIefGVpSP6P8Fmfl7NwJGqlUckysbbTVjGyjPRAz/kyqHjDnTOhKl4SJbLeOffMYM
cVQsbovFTXmc8sNLzR0tuagD0nd8AtKX3d78FEA/l1SLJntt57JSaMqqol4mhNeZkUv4SQxmrsZ6
N4PpmBRM3FkRW8HhAm3tZiKkUQBeqahh+EV6UnRCKKYnLUjG5LHogWFgVC0+c0JpGyhoYYDeH/Wk
3WaxG/fr60lAo1bNhFpmlALV8zBqooRRqL2TG/srqPIknlQBgm4Q1xAGQ4w33/jpXxC6eCv0rHT1
bqeH3jVnqYDSoDjGPf4AGw9sqFhLkmpVyJDOWcyxt5GftlibGIvubZk+cnb1sc0dVJerPcKHwh+B
lPM7Ot0Y1He9pCF/7TGpbNcKSO0kxp2lStMwZJiEEbid+be2QAoM3W2lU9zRf2mUNSBEd2VNWkdm
lKxX3z7fZdgXoaulVQa4V5H9XDCscCZNEjS0Y823FYbwsb8+bOtXBT3jeEuWRTHp4i4nLc+ta+IZ
bRh5hGQszWLytG1bsEAWZiXzuE87Ho43A3oM9zKYhgM7vQQtHxwNDd9pTl6A+a9bd8k2l4Vl1s7K
/cENfMiv/FQoAP2zI5IrRl5O/0LciumB0UKqQcd4t/OR8mzCGRyrWmuIIHn1enEcHm+e3KA2mUmt
7EgapiIytOaJxlHVHq1iyp6wpoqWtmRHoWp3xQFk5Y1aEoLRLm8+P+kZB4S2H4bNEZqRmoAK87wu
Ely8i3Wg/ORVLx357ZqYA+DzpnZilN3377smPv4UXbqoNeJBp+rdzKEi/Pwf5s8eJ4Oz40W65yuH
JJPug1XCThp7ipc0onSMIpqV+mT1RyzIO9BH+4tyF1fjaJH7zx+Cu70TpeHjNkXKpsniiPPUWnxo
8bE4wTj75tr0pgGkJvZrwGLZ3ILXrRC+ufnl+QDh++RnKSCrFzpMwGqNfiE351oN1xjjKUGL6UEb
UGq1wmna0VBnY+QvIHynSu1rFyJNwUAb8y6kmaqSk/6FY98YSRrkCwvOf0FpsvulV/FpxlTEPFt3
Sn3ZxasqlzZ3zgww7Jr5wvrzCjCTcGP732DqIaHrU5k0Ea1W5vqzca9BwWGpATKRrqC+sTdBnx+7
ymUnsBpqjzMIN3EPVU9Lr0hTVk3jic4THRDXsmkjzuBYCJGgz+aR9BhbG2Hn0NWis47oC3raZnpd
8zAOQN6lHzW2tV3fd34y6lEB/EhqIdPzmTxW9X+YgANn5bny6Q3m9qr8kvv1HxAaw7A1sHhqUZri
vMbgk8QtpmYscus12o4McFbHBOpnJkgc0m3XCr44gzUOHp1ONlXdNGD9RY0kP8kzlcLojZwxy21W
Atk+za8gvyYMfAbcpeKl3BXot3rlDK/kUtM4xTZwTKP+EOaEJcEXiwpkumLXxeh78MS5uNxyeksF
BfIsGPDEFLHDkT/7IrRQx1BxFBlov0v7zdnS4huYwJioZgnobkQUdsTvjKfIPDi6sUAgItxG5BZE
E+5LG9VeN5dgIHGm0dPXQilk1nfPV9dDbe0mtbLQwewcnmNk3JYXBQ/2zQck+8PTdN3U1ZWi56+E
erdJI62P7rJMMrD9IATmfdtviKJBP8ZETgAxGw6F8xUCUdijflaGigMVL4kGxZuErkOzfEqvt7Im
17BSw/sK4oHHQGOOg8vCf7COgXI8yQCqvPSNpWx6sVWUY5L2xFTkK+1K+YXWOrmJinIr+gGrU32O
TE7UTYGuS5NJyU6ubZu24ROsu4Jw4VOXbsfRlleQf1zAKPkptZ9+Q7pAtttzI6e9FE3iQxYlMPUW
OsTJlbzgZSqxSHe29emX19oHZ8fx8wvHEygfCgLAdZo7nX3UdSlybQ2b7heqC3M+TmU12GJDGAUq
9bHPwgLpNPJLHkaBxsqk4FJ2+/XHmWnzcvXa68nhLPVtAcU6Nr/rsJ7Bwt/Xq6Ejw4ua/ifHxW1z
TJ7PxhGXNfG5CTPFfX1uhaQuRkAuQit/8OwNs9boB+QEBwsnfruTwDId5aQeYaFyLtu21ZiyZNXg
I9qLafigQ87b0hcKJkToAyw5ZUwdl7E2Wrjlh5FdB/VzDppaGkU9Ejx3xAEdNOX2qsloxwCngwPc
cP8/kCrpvHCiDH6IcuMlUPVQmxiOfLk6KekS53WTC/FOIEDEz4J4WY0Z6JGbOE9PV29N0WEXd+qh
xhT27F/s93QV9RLia00NhvXATqYCvVkOrEJGHwekALc6htoaPmI/3uAzF1s3pRYIVhMaqOsQWyTT
EPLQwuxBJKKHi8XwSSAobn59+JuTMbyEBglTeWZA2KO39Y2Prm+44aLal5LXtsgMdj4ObHHzUZsN
zXSNb4b7k5OyOMqiF3deqSeO831bmn5xbMpT8ralj8FUcJKqfpCyD72KCy8RCfgEcAL/tFUNY0I/
d56K/qk5ku6Ul0Pn8IfFtqry6Glx3ayYjIagR0mFOaPS2oq4lJ9fe7PzG0QQnbt+cbLbgTqWY6WT
PrZkLjDSo1iPieD95YjpDn0ZNWTj3assUEVx4hR2GBAVmW4f/ypgw2+Y4PsxA0/TM+T0tOxtiazz
/hNj90+aW2dTrGj1xUphSclfWeQZDcv9JHTRvETZaXmtrQapnGSgGVQ+ygDHUuxhbU+oNGMyE4Ou
G3pwAZsRDffBlzLYsqt63iNFR/nuomBY4w1DdySgkTlUy7PGqwAG3MM2UDIXLg5O+ZZzUkwj+oGP
5BkEScfIf7saGGMy9CbZtEFdpiIHtw6Eu4mmrkh6l8Q6BX5+9Mj9TZMQTumFnu42Qizp6gnBI6iF
EtnslgITbZ88/x+2zqpoYgO2NM3VP3zT5ZFPfEbDAHRTIFTC6ZpncXfC4Qg7ktw7ddBFDXY5ch4n
1W/yoemHFNyAoz4mnRhizQ7NhaJZKVO3buOd6V5lLUc7mrRq5rD2nkDnuB7AzVMPDwHAn3/gLJz8
7xCQWh9FR5n4wgTO4AldNUxVsiuo8OVMZOVcpEm2gZJL2SG2PQCPOjMqZqmLR2mbj7/dmDyxN9mU
NJWqjaL+z7HldSKNvDrDZxz9rNkkAkSYFghlbslvnk9S9rxweUywMr1O9nEebFVHLdyp1GzdzOlc
iBRWI0X4SfBiSB6XtsD8p6h1/whU9JJ1iP1LdhXcBbOn5X4rNqHEedWah9qjYRm5ob+qQDQBVVg6
9XYEj0A4Hxgkm9zyl4TTs9X/T/6raKOj61SJW53Pb1XMmyMm3iT6aRyOW9an9WlyR8A01ht4XyqG
bSaqTR2E4nUg3cVjArovA1MUUwCdH1C/qWfQZu2QwTqU3z4/RMvzLQgTSaFEKOYpR7+K5V2u1EUY
iuJp7fjf4JS08lENR0w9H2avS1+89zEAh0vzX+9+TQvotLN3dG7QWVnDOkXfnQ1G/4tTLcTlKTW8
rXrzgnVTiwJmQ2p0kLSvnzuqFMfOLKBqhOT0bXcw7MNT95BmILPkMn/1KQLc3sC9Dlc3Eu5EM85M
/I14OVlmu/n++ChB3JO5sNVmUfx6OJCQgiUAEu6RrMBfwfkeKf2lru+tLC2JtvQAa/YsdaZ5JfO7
HqU8wgmWRGQtgpzmyycqy7/9eC3miHaQe7v5TLXvd+KgQmcjpf1oWPFdjCXyKEFwL4jeBpSPFXfy
fzKT2x+EgMvx4UXBzOCA6xNor6muYNpXWcxl5aIcMIL1ukm8WfVQzN5VbRaPCV+4pAEpWt9h7moh
m+DmpaO2fTkVM5csIYx85glnmPQAE6tynASqhrVBgN+fbSSePKKR5MAGUFXgsHBs6YJT8wEyuVA2
DgU0cdaQdZQostiWlu7x2SuOz3BcjlRq0Ll7QqogxmRzZq5hgDhDBAGzMih8/NeshHMLf7Czys1B
wljBhMQl0ksGN1/7JDFZmnvTcYNy1mRbgSXaKnfuchfYeSs1o8jLRPrVJTy8A37lKAM/Pm0LLImg
1E2oZTe/ssrvDSQFiYQRY+zg/ScITsO7Xh17JsQFeOlZVYj5GEIhfO39UHvyDzBm4p5hIPn8GJa9
mPMuXELn+/jr1tgo8tFTnySUp0hq1vvCn+j8e6ISc2aYr8HiUEEXmYkW9nJE0Az4ZCA8VNrOossU
I+Li5u5KvDHJ3dFgxTFKQ9t/DrDlNi5+TftUizJ57VJi7YttY+Do8kPJs032cvRHduweYAVbWqfg
eU1SiczqtDK4Ni+ndPrJeGpLEmaHlaewXxl3Mae0nTCXP593fhmDBUmL8/+3nmyN5r6rzSoLjYxQ
Hb600R1Yfkq3HOoclRGcmQKTxJOg+T5tZ1W4nqOOEkB/FIBq7SBwEcvYOB0gIXPc3L/VgaHm+MNS
lR60xLzsDp3xPwUnGAFw7g0GT3+hnto41CMUcWs0GKTxQysaejP9rRJDRzQIPcG0M+NHz6s3tQBx
/Ix6J9HRWHXBPMX10VgMbIXgDDeTEXgQ4ZkHNSWrdlm/cbDW3E5k/G99FtXhw4z0tB/zpmAYlB3J
qaSSla3/o+SZ3kFcniFSLQp3oCXR08gtf18nUNuR++p8xTHPCHxlOhvbgjVjqL4pKMpgHPMkfbrK
rCZWupueL8qBAxaEN++c8EOVEqF3KuB1H/2v4RLVO0lVZczd/rTRo1XHJovLCXHzvzu+dPuxuPwW
kRU64hi3zrAiL11T3p6wNgJzFTWPm/xiE0zR66c/IzZu2mOTEXtWnuEzxA45NkihzzR1yajtG8+N
6QQYH23InC9gFseonv+N7Z/2p+OG1mK/SHBBLbyDy+dyyLX6DmVoOkdQ74BcQLP+cu/772Z0GXDv
sWJk5Kdl/sQ/0FOzY1e9oU67HTyK/DDJ9znviuVFNLP5WHwfKXmDSjZPshZp9qDDRtgkoTiCWesw
cRouZKGiZDDdsKE4wKZLPDuNifwGIl95Ap5VTEaV5k+iAgLeyYgHJbsch/JT4agT7d9/0f3SUvWP
VdrEmJeUbSymAgx5T/Xu5V/Lo7nxE/bfSfPU8yMPYEypBK8p2Q385N2m4CFdkizUX500D1RmNZ0L
y1YRtRU8MvVNbK5ICnbxYPTD6eeFSRLyk9j8vchvMh/C/Thwr7SzmpToc0YIaK6ix09jR6mphcTD
y6/Xl6RBGuu+VbzLRK1JTXj3Y1yRobvsXLw7jYLsTL8MAa/RaTFc21mgyPjSTy5vJqj1ySe7lPGK
t2+Dv9THM2U9LsJPvSPq0GsoOsAk3N07WZppyh9f6E1YHEl9ApsQRCDehty0lMzwTBno/HCaAlSq
+B/0rCKGvX6T3qVgQb0wj4laZujdSlymVQL5fjikxKzK1/QFUCTNU2SwfldGb/O/rSBjWavt6X5V
OGYkGo7r06AK2Yy3rfw6Uu5e3zOBLbMCII1rVWf+ELv7X2yCO7Zq4WV84j/WZIBR70UZFHBz0LE9
3Z11hHUEgfEnw0LW18BL3cA4fDtPh6QdkWFtHiyk6p2LSmGnhhzcVQn8Bhupxtp9A7dCDA549OKy
CPqAImIt7NQxEPrtG/nSFBtNPGhQtlcwGnr4ERkX56wuTLc/VmTrwoZhsHEFHrnkzu9iZmlIeRne
bul8fjrJ4Z+o9ojS+L9KVaMGnPBQMviqaeZrKixW+OAcmqNoWddmbXRLGUSaakML1V+iDv6z4I2Z
4F2R8poF1Aj1InH2quZXYT/Gb4jcJKrobgmFBVQ3uyP72JuLNT2BO5+7WIOtIWS8pJWn8d1d0e4q
DPRoCOefmPwdREwNmBbwdURBi5yzqAgV1Kl5xAXiVJfllcGLtBXu3sFziDmxKIIdnbcN8V5vAFX9
3l7AFKT1RI0CCAsfm8gg8UL9BJQmV9gHPlNmtHQwosHiBILUZ9yrETkMWSB3WSfkr0nrAlQFGk7L
RRK8fJ3paUiXr+frLVZIpwONfgr3mrKa6bTkWjva1QnexqhkXeiv+W5CKi/WH0mWzoKciAVoEn23
Mf/hikpcnePNG/KK6bPwkZxgd+dtWf/nT+uTzXw3gbVzEVs8gQI4/n0yI2EugL5Yz7xSwIrR16U0
4uOf9jlMIWeHj3BqtN4fSWl94QqiHiDy/GnGqnOaqBEf+u8POpxJbRNVcFCKhMPNJ+8areXp0BFD
AQk9bwWAxovn7AcepSoSmfpr+atCrcOEfPipPy3PHfZ91COISWu/QsgdRGAFnWfPL0RsST7/y8Iv
vQmXK8qcGpVG8C8QQJHx+XY7DwVt/BaG0f+OmHzElH+H8AWyt5g9RlcarRvDDTrXsUPWWc33XiYF
1z5q3Tcmshx1Z0M7zNSE1fxOZGOYINKLjjXPH7qhUaxUXnzoVrWk9cQnDngmIljZjcy3065fPt76
4sxPFWfNdRKUm4drsytK7dVn3wlWmaLgN6JK0j7BSHOnd+3Q9bFTwF8QDNbJUDCt9/1fX6FB0Au1
7Mj6USNRSwJuZeIuTvC4f8IA0ciI5kTi1xR+QniPb/qWOpEgX4NH9/DxhvJf20vP7lAP+J0YABHY
b5c2fBHfOejGfAKXdjHS/Mw/zWEV0SmlCmhieFm6kTA0GOcGZ6eQ4ev7L085igx5zooJnhqTJ0Be
JAmBAzT0ON5BJKjEGL7z+5JILj8FF+jYhriNnB5lP3Aa4cnrI6oDVWvmqCNO7eUXBWAr0BX0Mem8
o20oMVKlGt+6bYkghYplERfgEld1Zti9dxjcpoDcRK9engdscHTxT0djPzDFW58WpydSnbgPWsYx
zUmOwkLOnyt2M1SLOQ5K8hSp8sRvPUkugdCZ7J4Kxw31UhsXoNyzXjgWNws1blOOJcMw/WfeXbqr
sFPjXaD4xPu50VZ9wmtL79gfS0/lNs6dzLbFr0QOreLSkXh0RFcszOK0BjO2GIumN5vyHuh2UMaj
OCw2rXlqXy5wVROqORVoC0554dIcD6PF613R4cj5TcsZGxUtgLRZt5whdimRoJroVgionH5Fo03t
ELUviK+haJ7unsQlWVPqJTPwghRh0c4Fx/vTdczh5JVREsq59FBlNciBD44AY6QKbUGuMXcMPN0j
yMrTw1PIuLl39JJ8sG+72DS3ha7W80fnb4Nl12m+frx6qwF+8Vw63d1CIdqzCqD0YGI8OYL0foyC
X+VVQ7XyNAcDt9BQUpR13nBnhy5cfRpo91k/trxZIaYMnDCrq/pEVJKpbujqP2kbx+MSspxt2Faa
TRPkMKWQTYtkHJhn4AJshp7Nufh0HoEUTej+8X8QVgQionESRqdCS5hcpX2v/AIyy425DTKVhCbT
KkOD4YfCDlSVuA8HIV1bzX/L3I5qjtHDnqYhBK3VU9yrULVs5ConKXN8DeuyyivSQoaaBjUparNg
f768nnxXMXWuprYXj3CX6CoOKmF+d5vXuCpMG1+8l6cHnopVb27FkJOv7gbAHohVVX0BcEmVDcij
Vpd9E5DaqI1BabUFUFwBhvrBQxk0CB9y1hdhbN7XnZ3WSW6M3rnYhabbW8sQQ+6UkImYUp8PGIPa
fzvGM2XV/aS7nlbalJAjH8FdJ93ja67WU0tJDYakV8ZafU4qibSiDCPDvLlRM0354bJEtzwsubHN
LqsCHnGHc2CkGhnNLkgXrRpCzocDMghhigZFM3fgPir+7tLzXIcxmHE6HRCnv7zKSLr61FkgZgjW
TS1GAgo0jFDpdpIYlx6MTO7C/eKw478DzPTNpo+r7m9gzhuuGRcbclQdTznGuoMOnYyyAyaeXNZw
Xm8W5iJWwv5Cy7dzCEM03BEdnoqkM4UJ9XTdWNnx6dDyV5tVldkw5reqcUr7h9AY2hyIABMudmjq
meNdTSCVetuiroGeStan7I4f9LlP8DNQArgbMDtCIldtzykbT+zvzA36dbfR0vH/rlQxLJqz3GtH
idxgNnh07phsZWYrpGsA8li2x2UM1tMGt7HomwxRxbd63GpiHESGs4Sr9lu5Wfg57kGgdfBj5aJ+
gZ2ctLy2G5r//s8gbUttZsGXqsJN/RagqXVIXI7BhA6woHxpl+XJah+TxCycQd25huQ2AqF3/LXw
ius8alYTTOZtvbnTo/uuP/44uv/X+3tIQBkfbXbmsdl2796fe1+fZvfVvJUVmbMqKP+jb5+ubksV
AmR6IWKgIDI7rE7gR0D6uzkuOkYpe0kFFfz4wVTinYGvhWSTzt3Ol+2wsAXjk04TEgXQSEA5VbXI
02X4mcPyTMV02P102+UVGXU8WrUaaf5Ykn05sXwkmrXU2sOyXe/XOFCNtaA+ptmnY6Z2G+OkS4CZ
nNfQ6ANxSO3k9/+jamCIjIa6lKX+5Ylz6bFyk+6ndaeSeMIW95hu6gcZYryIuZwV5XxvaQz7c4yJ
JxhLExAxszoRWrES+06EuWVOORebZ3OIx9hUiwfGMx4OC+FYGsLeIJwo9JUUPnJaRsqRT1Y5XAsF
z2P4E7ZdLwcOSJFY5PRrsUD5/GGjbTmDJWITzhmMZkIYFLHa83WEZUkg4xxzSbM4LnXVRb1Vcjjq
GhOrkcTTvIVIEuf6GL3wHHw39SeLdUAuXX06zwFaP1Y8gQ9XFOrnCy392Ckfv9M7o2iQ6GgaUccC
2ZQKbrF0cXdsAdRXYUK+1pUfsS62yuO2axNQ85k6QI5TPw2qcz3QEtpcs0e6PO/a1LJFbi2rh2S6
KLqjaXF3ilo/VF15Tq0XXINybMbaDx4GYNDPR/oZDL3GAqPl66uaSKGDkDz5yWT+e/aPEOZ3YBXs
x+caxTxSMGZZj2u7uheK7nLc0r3oAFSV5KD2LCdFYrI1YC9fLa5pc06d8UYQGAVt/Uf/odFyp28r
g4sGEhslu7eY+zNYWNqOHIj2fEA1QkaeVvhnK1Tqq3kdUsEG12bP+8Xz+qgNNWwsK//c5jrvamSp
+EKHROu9nyaG82IkwVBaIfjlw5a7oZ9fWuXAcIL38xNda68qjZhaYn+KyKYoM3hGJhyfdj/CVu25
AnvgSQ4yFklww8ivewgrsx1dETCGTWuOz51mAyf12RwTHO9ABNX1VfEmdIm6LxVCPkeqDMzAgvnu
dZoc7LbrKDgG0x3bflFbnn/ep52rS3hpkjpBl+mdXhpNNPvGrtugC920enLGgucWnC5eii6BcKD9
YOstXB/FN5nrUK0Tn+xGcW9o/ddCRM0sp1wHCBW9A562akv+08KRe+y5DTw4BJIUgPvvTO0I/Mgk
PPwrNuGbcZH8jIzfcQCdTWfBMWkv2Q5pvYQKl4cQLGL23WtP51UKVCczHvVIBDeYnVUcWT+rcvbQ
SO6ItWMTFVbr/NgJaEU0qPEwz069v9gLV7psiK0ewtKOfLHW4d0aYolEKmztGz2g/47jCpfDuk/H
Qow3hc3I6DB0IArCFobO2eCXyFsQ7LebpYKTM3xBQ9PHXIewI+QuEbG4UMazGzHT2okGYJNHs4nk
21ewDZpL7TEQCpcIgXHflFgA1YV6QBSimAofy1uO30VgiVRQXxw2mnAha6+km8Cqi7sCZ12ubPsH
eUAMX92ozQNk1JvG8CPtSeZmQ+gnmfKKdcLV6iB88Vm3I/6llXkGFZz1cGbGMoBjwR38ciUrisVu
sgh17mEH0WqVubBFAHzUMDd7nSEt9Cqo2uxJObEOwix2cn6GN8URkiP+SldZ4i6gvX4dWknhe23b
TGpTspRUEV0Dp9PJEXUibwOAfXwKxJE0exUwQeUbEptn7Gn1nbSGcDuM4hCzZxPoJj7xGjBuMTcp
utWCTsm54I2c9m96OeSJdqPWfbPnr4m7Sa1YqDVT6vmNll71VQSMF7jCPloTKVsgyATP50ex8Dcy
fxZ3/sMD5J540ZC4vHLHdYR02UX4KRYP0dvVSHS7R7txvEXm1gmdXIEW/WYDzn5SzVaB0P14u1la
TdzSXassGGbS1m94eB2WEoh2RwU+FxXcw+vClHVJgGC50WD+A/EjtCqqm6M3MDvfR5Ey36gJKJKh
KLLT/s9+2aK6sbRkVsK1+h7dI98re/5bd3HqWA3hHuCWrnwLLoFB2eUL1VWYiqQ58UCShXzaVt3N
tovgYiF0BlRcqEWLfd+A1A7JcYrKhduiGruPBnOv0wXOcJz5I88exBWB/o3EvMq++rW78C3FthOQ
1VbyyuM9zSFFbdtwx0Z7ced8a3Tir7dxU0kzt9E7BeWRFVMhQaat4dYlpmVRjrvqRWKVlomKzvLM
tIwAN3K+VxpsE3N9YR4oLLBk0d425SY9KwbWsrrTV/TRVwJvKIa2BiNe37Bo1celtpmgrpiYXNx/
pIbC1BjZGgRKVr9aL8edNbUL9cPEWoF5h7ZJMcFT3m3qZk/hvDmPKxFx24t+U0nzJJYAyHyy5Abu
x3jpa8dk6WqGb0TXNfL2qiKR69PsmjjXfg+oq5IFApKK1yBsS0dVszk/m9OgreJ1EqVL7JUWaZG9
5lcsiLAdbVbBzC4oBdrHyVtLU4I6JZavOwWFXpuROEUuOJ2Qu4cjlFh1pST7TWkRk8gJIsuuSdmS
cEgyNKrO/BV72pO/NAcQblWJimP4NInXAt9EWBS9n2jKKgdgvLlbcrgXSMHEoDtmFFz0QtR8uVHH
5A/gx8oNgNub4mQKkWf1zfuP9LBr/7F/z88yXJek4Q/oUAtyoXvD7obm6kBoTGS7RSDNuhdFR4aJ
ReHIvN+ADHZJW/NNBwzPaWOki+XyzNQSz0kgjKbq77U2uYOpDLO4n/YrvkGk1fqaksB/iCrv+eZS
WF4VGHyJomilSOmkBjbM/6yx0aOZjzC9MJGtbBKegyQnilWAXt9+3C74JTvb65++sZjIZDWydOmg
ZvCMOOOL9475LnBbDUZKOAwRWm+tpPcw6mU0TUI8BP/FKEqW+CJC48Zrt5mcUDO14RV9ozcYF4kg
CCt5e21iD2wW96Dusp6SN/YXjh6dW/7O2kV+GxqgppyfLF6faXIG8QIVVkZ6cow8iPSXUxQDwQ/V
kSfV41UeDXt/ygXn6ATUaXNV3JMhoTc/ZgWg3MIKpGEhP9zXrklkFeaFVZrwpptchZ01CqFcOYV9
C1/cEHkGDQ9vngrXIQX0IIvv6arr4z4lTimGFmE2EdbTHZvoGJVaUSWc9B8LHt1ol2YVzt8vExfa
LdpCyyT43Qy/MTmyY2/nIbXZt/eBDRz8K20HRhD2cY9eEN3/AVq1HVAAyTLh4ot7bPZMk/8wlUOx
kvt+iC8Z2Fw9WqEKIsyUr+b0qoMXVsC9AZUv741sTvLUEvXEAIRoF1L/C/hLAo/ifoTaHkkI4sRL
qTlhHeGtcXbNPXpddK38AwHLr+fgzBI+gQP7gQkSb1N/j1NXBxX3LHgYcVK2/ip6Ec3G2aDzLsWv
7hQkQq66vHq9p2cmKfVto7u9ZLWF8KVFKweTsXUazwDcXPqGeoTwDG11aTXM9pQwr7vh1J6ow7V4
j8lrKfN+vCEJrvSFoOstXLcXMxTQNQpT3M7LmUZ86rlbtM6cRSz+CNYuWHMkCophLWPhyKChL9Hr
vyhF6RySF9vFOuDQZEKrMpBeFQ8MZeq2vzQUp/6943tppQbvGkCZ4m3koZHLndwBSOhy/yhVOUde
cIazSWCcuZia+fLJOkRjGZafroTLPI80frzgFm4/zayHlCiTLqOvEXgYdKGGWC5LL24ZMpk6Xlsr
qOL+1USdA/2LhcPaLyFN0LzlRyldXg5HzARsA9I+8txEsMZKFkPu2LhPPHBh8g6vtLTKVgbKFT5f
Ummd9DGvDqC1g+iNpeaOjJw4t+dbNnTqIYhGGZ2DOeyrC+GFMtN8SjVVPJoCJqhfPCal6Cp4SX31
65+vADN8Q6ccFmVLmBOugdVjRx2eiRkWyDNyUZ5hlICey5BsSd9oRPp4OpDZLfEiL2oZUHlmRJiQ
U3Geu3ULYwkwZKzMWl1NST9BcPBVxyx1Vi4aVDzjNEqvNOx9HM+ugBosuoToAZtdh16d0ivpi8FS
DPIk7g2zCkB768d3tF6a+K/2RH/Dk7zQUX9DOzI35TNaImT0MFAK6z6JmdgXYTevAFGeH6fWKeKV
8kutql7ACzJSZ5IkG3DmwLC+hF7Cu5FvFjweT77bqQAnnDcosYIa/S3JdqOBh7jPuFaS9XklYiyz
Lc598vFI1p06exgQrvRCuvX1qoV+tAphTlkzDE8LUMiFcSwJLnf6N9bB5iCh41BfJyvgyB2RNsQa
cvRsJdYAaGqwunFhGGRRNiEbLf2vlGa9NjGNp5kbrrMqAvQLXscmVM4iLKkSGlj3MI/QkpaTutJN
uybZeLrkRWu2Clbyfzqph27jhi4zfYNPGAuekPXOuTf+Kli6Mxg7c5ndJXICH8c8TLyAsxzdMpjv
BYq8ztpydxnUGf5ErTCNzpuevf2J+rOQKYh3yy7oxGAMJmSQkuSCx9gSyxvldO73YEaSSVIM0JIY
SCsUVJ+BGZwpcxkE+fMthdET+ahxv2J5V59cjQ01aeNVuDCm+4YBP9HCabT4GEQd2uuypDQRW7gw
P7Z5ZRQB9z53d3c+ZjUMDsqGillemDDeYEDBtg/zMoT530EPXjK3cRgBKyI2Pk/TZI5ICs9yhCWv
e+7adiFXK3jFSXKK1dbV6CDwxNpNh4FIOdXiNfF6ABlnax45AD2gaVDqaD6GffekyAhqBsvpr5CH
N02BAYvkUCXvG+v8mUjbCjNHJ9fPsT0EdRD5Ov9N6KHfiEVN3kUAEsAyymmz7dRffzXx6auFfFWh
z41MwAPM4OCxIq8J22rhhWag78drMutHuFZWycZBANNywtg+QXKkRXBZwy6viAxxIUpXIKuAANud
yr7Z10nM1MFXCdCYpo5ANxb9Hywn5laZyBm9Bk4leVcGABT9nmnxHo41QFqRJcuXzKBWvkULMIqa
xeQ05gBvSgwV3SAaD5Tqk8JO0gzgSvuPVt9g6+JPWnkk0VpNxP7Upap1BDdp2dI/jyQxrCuei39T
TqJBUZDNOG8Tpf6ATBADkLZbton41pUsRvRnpAA84o1RJ1Yhr4a9lNMnN65pzBYSRrKOuv6RhRi/
pPHME4iPqJNPprM/laPoDJU/PDYkCO92ZjxSF2lnsl1OdDcP1GvTbmEYDoOzcqiKg6Xeejr4xn+I
DaCtezvJKgs3BXAE+oNt1tBMBQ882qwaZKqkxLcHZpg8rwtO1gN/sckyLVL+sFZkv3Zg11NFtzbT
lbbKYEgOCixzkPqRiEb0HJDg9fxPlmjr0QewEWo/9CsOb01HGokWfRpu8j79xxqstTMXsnjjkbtN
LMZgfebjwrbjPOeH0GYfu/o+7V8wXDTFyWHxt3CC3IA6fKnVNBajH2amWmQD1K7JG4dpV9ZZwT+3
EmHMuITazH4J5oU1J0eYdqSwTf6BcvEd/06XVqaaBl5plmErboFZEVaLx6G06CTzSZJaa2NsUp4X
dV1t3+w0C3HzQVGUyfc96xTgcXFcj+QFq/RIpR5vaP/9/7c1WuPJ1tLy4IbZpKk+D7/uEa5IsDiG
LAClcfgh7vi/VKyo2UDceFEDV5DxFt4pr+RadFN+7hPaDUmQDtJFiRDU9aGDGrmVCRHxoYtAy4Oh
+te02ZLfbSthQbCLRh63pH+KKGc3uer1hVdho06z6pCfltbw85o5n1bYLIpc74hZ+PnrFVW1zr14
aMeYSSC3+FLWcGhTYSEQNoQq4ql024V1/rYNDw9rVmckce3ZNyP4ITa6yxjm66CwPp9o83X7gOdq
sWTsVjayTiplepkOKpqhYOETIgwuDjBqn97UbRZ9JnhCcGCt8fJY2v254iWUkbfrYD3n63lJpgRY
qhYXGuxCJpHujPsFNvDBO98fSqjif9gha2sIbwBKxoNa8MB4orYVRfwshIHLFyfCb3haZ/gx3RZn
FSXdCec6J3gd6FuJdozxTSzR/dK0HC5hVVeTKhkDI8TdDkVMmVrfx0fKSGq9kXlA86JnD44FVYaR
XEebxgY/iksvKBYSkHAaDDugNTRQom1cb6P01DaJs+YfuNNcK7LHaY5CL22uka3Y3eb/bVV4E9/N
vSTAS6SNCAQTtej0FkVYDH6fXkYsNxvrfanyeH00jFp2j7PsaOHWN56/xMEqduOBA+TI8d4noa0u
WaZPfnqFl5SG0oDxBs5aJADTiRA6RJZPqVmYSDRXDlJ9dKZ6CNEOWNAvZaXm/YNP0AI/010S2iXr
XmqYKtG+wdSt4kXMcSVwcR1pASNYiozmsYxExv9Vp6CfO+fMALbFbW/R0DNwVBC1zo3cVV7mAte/
eXWzTre6UJbsSjwcCt1jW4zZQt1CRDVgtA/Xwnu/f1XxBt4hvSswMCkG/2rvHq6/ACSilgRrwFmX
pAwZTIjxNiusvPG7BUeKRgynoygWua29Tkgz5vZMfj4NW7C0X44hbzajbqb9ewKhfoNY1K/Y1jg4
ZTTwipVVy9G+32sVgrvAURFjlrZ0ywbvAor3RTLh6CZ67trWVtz5bqD+AE7zMllCf0JuyyaZB95z
sfEnV/bVexLvdoANt4UvfmJC55LZciIxNiQR9ziBQnz0wv6oJObzf5pk1oVLrrn1YHT6kz07LzdX
8YNq1wgwOg8Bv2PoBZLRA56X3vRlHQRPIse2erwp87XodBf1jY0RsHOvagCDnp6e4CozmkeVUHq0
wUKUN6zcvZMdnkWCJIDe95mtUfJ91Ey57gLnVWfrNVSExO0IoOlxtM7JenafXQ5Ci+RIdJ/JSx9A
vg13md9vH363nvn1NKV9HD45EmnP1rNg2G/x0Tg28phW8WdKeuSR5aoSMsS4mt7nNKjYMBvoukGh
kaxCPCLWNyI223Jsd7Dd5jlE7PHnqkiWZ+DZWk3wg/d/fuJ60nagVIwdYKUpKMCujhPIp1zaz87L
f/8Bo9dI2Tyx8C2zfGX6ZfBSXbtF8d69IQTMNXNdKweuFpqFjmsNwJcNInqawGvrsu3itVfCxLQ0
QhdP1ptcBRtzfIwQHqLxu4B5cyVrm87kN3Xa0HTOVCc1qiANCbwVR9mOfe9mrdITBXmwZ2LJh0ZK
hYN2RFKsv3Wt7SOEJxP4oRbuLrkO33xDkod7dCVsfYEWrcgEGzaSo4OaBqEFMtJAa2A9mpMUlewf
QK6onD0Nbpfvzh5EQdMj5Asus4lVABv0KGfUPX8kNkRgikI2Ddbj2ECMQq2+ErNei3TW/Bji/S7k
KmYsONQRjWgOPOgCeVE4DEKJchE9pTJXRfoen4qwm3L8WkM6Q9q9quAQYeLZmyAHrOVUdy0OPuh/
wh9tA1AT3LoBXmKX4nMB/ulVOBOzDf1ZCWsAVrkULMkrDwpoop3PUkB1wkpY2aTZg+E68rGCbop0
s0v2ely50ng+TgTSx3lb9/k/y86H2y/GLtZ9yuBl6Ned/Z5inoSIdiNCd19y1hqbpHiVXc2mpH75
kgPSX4+/SLn5y9SWmGAGD6rAz6il6sgzeVt8PXh3nofAiU/Mbzc1iPPOwk6TxHI6lCm6ZbJF5Yy3
vYNtHmcPKb71JdL9UIgUKsg6S9Xjz4/32Q9m+O7pNO/EjqWSon0JmfkOkh6It+eRwGZDSSQXZBPl
/MDELlYJAWlVgQ/2d4J/zaowpOE6vAGVniFBDaTMRRDi4SvwK9LeFl5FxdoFhqrFPPiDlSc8gXLY
9jtbNmSvaT9Y+qZuuLUS5Vi+naVnqmP5vA2IjE/4S1otCdqwPz9ZL7cHVHiCS/Lw7Fp1xHrCn7x7
a1l3o6tyhm5+cS0NLJMyoD0CcEIuIXCByW1WE4/GjcVUVlZp6sLJapGhGSUn/fRKeFzCYGGz3RLe
jS8uQPk4BTbAqaPlhqWXOKO3TPfcY1KJLCwqDKMpCn699yrGEM0ab0DQYGDrGGWZGF2a7aULas/y
UZ3cuVQOlAHg278P7e4eR0LNBl6cYflL3+tYR9qY75HIEmLAwhLBDnMWaosp4XAzQs/3sG3Oz2Sp
NiMsMzA6fUZsqiqr7eZL2U+7eUDi6WwNbxNP4ysix4xSr5agOvqzLQBb/zcwyBjkg72whA0VElX2
MemPDjHy5j6u2z0U8hnGVqwaoFiCXC9eizAP0pLfvfOLcmM0T1F7ZtQMmrVh6DfnALaNkOtRibtX
B3nSrSxm1VVHMmD8HyuTMPbxHdKqbiCz7pvAFqcsO/vzK7ZuloNXrdOYfkmW+wwxkjijw1W0Q3wl
AXcjqsn0YuuVzdi44eMHtrgxhZbqQrnx7vr+gpVkxzBDiFdaiueIs7gnqE3jDLyHvDoAzauAUj5G
tLV/IxRB8aKXfy1Q++myAaJwtFg310iR6QPNiu3/MLiDWD5aQ1IP0V2AGMIzFlV/jRQyJ7yL2mV1
yDQIffOw0a60RPjkTBlGjm1x3s9ux9xjU70d8kDkAGuKsFgJCSDJyp373TUP+ANwbAbfIzW27EWA
KvWWDx861WMck31cl+cpjBFzr5pCi29FtqySTXBjGg5mCxqTE1tRo7o6xZ+mkwpcFBiAEejc/3c0
fdgkXn7g/fSer1papzRzevafZ/Xo3VavFnUEEZI+KMj7OThP+lThrHtU+2X6RRmEgBuxKUkJ6f1/
Oa9xJOCVB9niYwh608HvWH6xQXM7WzskPhg84YZ1ZHEgL/gzzQtetpZh/pHXVlmzH0QLP2gTfpN1
suNuhtE5lEis43QJL/1yvx9i7XKUV2mIKEjflxC5s/nhtJ4Z9Dux/9wJLtnhTYSfcGyzvjpy5h4K
Kl9vVLegwjFAA6Ivt8qkYoAAZo/xQRN/fOaYbm05BwbH28AMm/OYbbJvUhdBcEdC65AoNALule+O
KD2UduQdyxDAIqHaSRsI3aR2LB4oJtc5ClhPemJV2IMODL/QwHuD0dwgn0I3ryXdHxCu5Rx5d4nQ
9dY83lclOjcBrA06j3sgEbq6D+33RlPQgOGKTwo9mnIZE94adZ1pbp1wk4jd4OIstMv3PnYrsywl
tZU1qaarzAhxkAIMIc4epGlnCgxwmz5MF1rgDLNDAJiG5V0nXzshBU4BdDi48DLnXoKRqXSXOElA
BLQ29W3PF5XxTgYUe56AlfaM8vJrPsX9S5hboWcDbPpBrTeUrWDV9lVhLWDKveOIY6C7PbMDGsa7
ZJsUBCkvAuf1GaFj8uhAB2R0eXI9zDeA0U0Q6KATl/+2EqCu3tDc6lMeBhX+tTjqP8BEAkh71WIK
MxPjHPZVMZzCuHvK/SqvSDNhJaEacmXF7w0HjDmmxEBG9qr720ADJoO4Iqi8uC7kLascyzNDbymi
1cgM+FRAqfWk49hCmIgTXUDWoP5UABZzXPFBA6NDSrIHcgt6fEc57xQT2jCB3EE8VhioEMQat83b
zGk8FFpDzfz9a2BzgDbCdYRbxinP/jMCSMgRuXrliSjMVPFkTcQH13YTO9rnoBTIjJnDbxblQ8vF
LgYi/6vpxfH4XUVp1olbWwR+z2e8JAHL63VjD0gX0oANjUEBm7jWcWAedcbE+YZeltsVLK+88Z2D
tyscfoZUS83AhHVYsKX3oeqkJDCywcU12vuwyIydyNizD80KtJWkhmcN2IrYTUYU1plKihKON2qg
oU8D43wJVyz11LeNuaYXkP4RNOMxvDeCbRkDvjUv7iXS7cbzELHTOwG7oMX+jmrXyF9FTKrLZ+MW
RtweNi/fALWa86CQoEExhr0LmNLXdNYcCuv5JD62apcS5knktAEcHdIMpGcqJnH8bEw1JAoUpvv5
GSvQ1SH3ASezHie1gAT6XI+chHJc3t2Zb/eoBzafBAW0ZY+DA3slO959BP1lgX71+JHxWll4lHSU
Iad7zFvNln/kaYnjGfdixWML6PTMZLrdQcUmeN/WIZDQ+Uj7WedmgxtBHjc44iZUSv3HBd1UFWEP
G2RFVmdm4/5HSMuEnGxstO9j0Am92eNxGvPaqTHs0aGAqvUinJcUPTTPmpugooHc3z+/lXf4HCD7
ozvLKZouv+Rjet50p84q24mND+RCzpxPrNMhGyX/efSfW6kIC4XsWSljwPHaIC4/3pScSRGUoaVA
D/BTDs/GlwXPAbHT63yUBtZM+byn93qEp2lbWojFVRDgHMhDdHkECyUiUGSKKiTBQyNEtMz9I4VH
VvAjAlzPLTCY3lP7cGUR+CVE4zSg+R2GWwSdM3MaVlv1WHFGBi7EoA/llotjane3t3t4kAnM4gA+
tnAdOswbmkLQSowJvcqoD1rWJ2cpDREaT1IElTUV4flFdMowfYJIu5Ng+gGi9S0iNYFG//KlPVF9
IIttHHzseshmLR9rsYpcgxKom61T7mZsE3iJicuX5g1V8FdWPJxTApjUc5ZTty9A1Ojn/gE9B74+
VxAEXkpQxn0KYKQ8gy7AsqVtGUg2YKopQ/9laRJ1qm/ZLJ26CsbKJJGr+EvMtsYDIgjMHYtgFieD
xmlVSABanXrKiLJl16FfMaWnJQD0Z8IYnJbTaKlNx1pYdqwpHO1l3OrarAhqrWKYYRP8TIKyNMIB
uwbJhl0jN/AMjdPLFCBw68m7xaG5nESfkgA1SLc4gP1mvPlv0JZwtQWW6qpE5MDVpWqX9Q5ABBcp
pnpHW3IstYYmTkNZfl5qGC2nSmQuWBKwxGv6xBKS+bE/IiMtfWLtNRM+YNqI3UPQ9ASrqK0r2q0C
UiFqcPfc0qWdRo4/zunxgHCE1EXMYjxIdrfa25HalQ16NXcU0xPGjcWA2G34OQEjYGLTmxkOkPEw
zLcRpJEqJn0LorjZYzyqEWTNBo1JXcBUkS1GClhfY1vkd1EBJr1oYWqxJVYCKKPoDlEpVMxRPUwl
TXq2tvmhWmTPTIrjxAGVYUjeuOfmg49nuNs7Q4heletNgxKG/vgnJAWBCPebsCSF88Y4xb0NbJOF
vvdQkKwmjLN7CRusvCBPxOaQd/FSaHhXPEvnd80xMHfXaDDN7NVMFibPE5ROq/gt0yzSX3CVdJRs
/Gni97kj31sFrLZc7a4AWAJHgsAaoKJ2uu5SWUWrbxeKn0Yn3mAQtmBplK5uyex6rA9jO+53g1wj
iVlFWuHEIp6FF7Zui4c9Vb70SMwrYwFASE2QdoiwacHhgqRh4Svt4/2Qw3Tq3MJ+dGAJ/OdHGcwY
CQpjDl9p2etoe6HLyAkJrIdRfj7sSL3eg4yUnIq/ztS10X8LyvaRlfJu9ctLu8cCbxe2rtPg1JGS
A09fzKIdmBXB10YlIoGBOCVpIMx1ul6BBp1IN0soR6nx+yzhKh0udTWnFY8uVSEXlvqJC+usX5zW
K91diwx0KkYUwmsyPzSR5lpQ1AKuRFz5BRkO+Jfl2Tax2zuMjSuUsVwT4fZHmzYec/WF9YB3stMH
/Eo/1agWPgydzfyscmTP89HQfonfDzvoVCcBZyVug7UYlglVdKJJnLX0iTGuhCJJZwDupcZAjZ2t
D5iDIvHCnjEnmLwbGvOdjR6f5Hbp8iZOGtCyNuiZTuTzbxey+mZZSQPuRYjP+aNr6M6Iby7AwedQ
X2mZsije9tKdc5ZD3nViFTaeXqvMZK2xbrgNAnLBQ6VOPjHwEM2JV2MuS38ih5uYRvY+ruemzk97
I00A0mh7FpvFiUdwtRrGra92DWVddnCYT9t3NURz+7tsQYS7/X+2sJOOIKhZRJyoplday2HK4Usk
ihZnLv/d5CeF2aF8vZEPPNe26lf7fbKk6PVUtX2azPH1eo9ZWJs1H0sm4uQCmRhj6FRzm9nJ1TTI
e0eIB8w27RaFnM4sy6qJSqvtfjL9h2ZpoVPCxt3lf21OWaRVAK+oZcuzAu8WrjwpYvSXlWwMNP2c
3uCXb3ZGDtB79wybBJeDbqfYf4domooJsyEn/AgIa3kvpKR0l+MQo/Kytxl0eS+Q6gJAOKXHujm1
bXw6nRTnG28grG6lHnca8KwI6rsM45OP3AHb5gDxKVKmHJmvKQKX27SlgtSckcYXpSLMJcORv3MO
qkbMHw/kjzyHzFI8DxeVdW2E8gUfTvHTUZ91eO6JxBjzz41NBghzoU95b1HvTJjV2919yyyeMP1w
4FGxE+yvMRCNLFSyxM5wEpvnmrVVfEtRuiRNaYZ9upj3izTnO5F5WawaUeYPuY0zF1cU78iEBVSq
4/SGuJnFGCtzImD/i2esxlzmsn5PxMDhdTB7xF973yuPm6JVbhQmqLkdMdp7Vq848nLqMqxc8NDV
6rA7S2kwbbY5JLhiQ5sHq8MJH4aapvBnWtS5QpIVblNfuzwISN+Z6jvClj1xAgLR22VOOqmzIWvL
RNpKFmEOM8c5du5riSur985eUnwVo5xYpabhnjNWU50+vS35kwb7QdWeZRdMx+UHggS9a8qRn5yR
IwZvgv2n29b0Tshk5MZbYXNTs0Bj+4auTjPeEk6dpOU7pPzEo1DtKO99XRrigMISJRIRfUZ8ld/O
TUetA5prLZJESxcoYabJdafJI/Mx/uFuzID6USrqDHGf5OhWAz9BW/titAnWSEpqQFIprFl2w90l
1nyE1WNrROX/tze9pHX1iuzbrjlUoNGNqRkEYCC1Osoih188vCIm9D53+/gOCvN5TWE0BwEB5xYt
5me2Wcu5Tq/zVFRLnmXRssQfGg0yRv1cLspq2L4GUV43NnjAM8vPL1WVo3WIQdwD+a1P0uW2rJXP
5l5pPQLbhEXOFa0E4xU8FPC1SI94zBF3SCbGYJ6YBQhiIpSC36Nxg6RX+krpIBLSTNBhMBFl3KfV
gyILQX/FWyGrJnm8ujb0lAsKX9EyFVhZcrEyGJJ5ICAhswJ2n37beLsYwRfUkxJV7JltbUjCKNXT
iY3+YmVMD67p6bwkaiNckDu+D01wwAmwompBpQdr4aaUUcwXKXvRZDbOTF3D+sY3++1NiadkVasD
tHFOOBkZGdZD4XoTJosIX5fsSlGxq00rvom+v7O3sWdx4WhJlT7RP1wMQJ2sAF40ZyvAa8ekQ6Y5
E1ddkIADbmvJri99hhvsrOzOrGMOC6REIpCJZwfCt3cDxFOTbfE6+9IHRxGDCYUSGxTjTtKkA75U
IW1SX3hLPBujEyJgw+Od94pzK/VAG4ZMKIU0WZcX1fiOzIBpKYXKpNezrAeaTOvva+f8/IMgEtPk
OqCgZcg2GeONWL/P9t9sIceM3/qL5gudK7P+3QVJnLipFuuKOWXyYMJb1AZpyluo0GlLv13llJ0Q
+GWVIZl5mLDdDCVXkPNmtU24kmzbgv8fTPpxdTj9XOoWp+ph5DNy4VeJHMFs6TdZ4vIoBd7NlTvk
OwiOCeZ43pGkjpPTQ7GI8okkhdoj6rOaV5flAEJXGR0TLO7Ijwe/RwnQVJxAQDCdhirujoXNFkVl
vnUawDTKZaEQ3vZRs3EMXKvPdJpqXVNRdKK8VGuaZtOf3apNIW99/yNnEW3dUjLHQykmo30Ej2sp
3JRBIEyclXj9Gg+Y2/Cnth/ebvhVsJbB856sqRs1Ps/UzkiIYSS/sXZ3Cq7KoY3hP/W1lpeLOZ0S
q2moKVDCBzd0ecot593s5NINVk9iQcH7CMXfrneThxJwFJRKNVcCs+Y2kBLnHtAHOf9fIQ8H0nTP
+aGdPmWqzHzQ6WXEOqXoV3NDM9erz+rYNyagoPAvgUyfA1tGjjQrsyvsHIw75oehC+6Z6BS9aVzA
1C2r+9TPveehbGU8XXM5ujgBHkn5RuLv4xFyJky2WhdLpiMuAH1DTfz/zd+a7kBHhzwICp4ooy8C
IJj6ys6PYgYX7jOliY0cF3o6Zt6T5QlJlklqg+OMi8RRNObWdjbWk4YkVW5Yksc4n4aiWX4qnJAX
m+FRq98lJGKSyAln98zp5WjIfgCh5GoxqT+1kfSG+hrj5E2R03oW30BOEvlrQExl1yAraXqecM91
pVyP81TqeBpuknN4AHKJQ8Y+yF/5zlFWUn6fqBqlklKMEG+2mn3XmkMXy6afqtXfto5GKWb4ZuiV
weVp9Z8CNpRRIfbyLNRqmzIEInIqkqCtyMlcp+dMzjv5hr3u5I4l/qLsVF/BeRN6ePSD5Pjp62Gl
CkHQYASQyGC2fMp6Rq2DXEsRNA8Y+rH9q2eZIzIp/1lDcV3o8++5VBXU99gSwEKtnZSgJDtPKFpG
swStoSu/FHfTIRJMuvZcOiwXvX+WRJ4JL8KhfsDEjo5OmTK4MC3kmG0nsbZopKR6/qdSubzVUEUN
DkTnJeU8X7NR5aYBgudjzvj1pDUkXAl3Ea2NMNoxqj7xqEHAMzXBGQvTAMb5Vi+0HY0chQE9/zLS
mlXsSRPy55mU2IeqxB8D4vx93znnGbD4lhKEYVjZjsUoDB8I9UJtPRKAT6qkgpUliA7bptvIGXw1
bemSooNDO8b5C0YPu9FxbM2d/jQ0f0olpMDd5YE5Jyo9vMnHLCN0KG9Z2QAKW7tukYqWnoe6NHhK
6NW8Hx7t/Pu4JLberPhjMsXWsi8oHvpma/kDtlQiQcHmZNw+VycfrzPBB26Wi9l92qduJZvCcNWb
REsbb+iWH8EQwIPIrFymDI8s7pokZEMX+CzKPxZGWbEddAsM4VPVJzB2IG03gMyonO9rZGPMvhMe
1QcQ9us6fJyCZOR3/3c4yUWcXIWzoKTkGboXfyUCyrirqltN0ef5JXMBqhLltgBwy1LQXl8EMP0G
4AVO0oHvugzt1vU8J7BuiG9CVuIxgyEvcWCrO7wZJlHDO3dtEAdsL/sgBrY5q+FH0Cs+D4l5O+l+
Izvhso3z3L6SjCqejKyuyrkynGz4BGTq7vjnBnFU6p9HvaqcbjFCYN7ej5dopEtLvUSP0Rv567lH
aNGxoC4e9rISJK6WdPqzO4S0C0fVpt2CG2FUtQhK04z4GjxMewWj61JozhmZUr0+aOWsA5ajKbqy
zEC/7/3S86LAFwrzkq9tcKC5UcY3uG4O0iVi0UKP+nUI+UPWUYBBZGJ+EKjNUljw4YIJ3qKQywM3
pjtQhyF5tlAHX17RKSpusvy6ZOv9WNQUoASmoqYKRm1xlJoCu1lTUPsIvsY1GIcpcKr4ZCnUsTsi
l/5F7j4oAVXh+caaUPGrXun/9teaicKMLnSmwEFOwbmMObehS97jEQs1I6MBykIEVxQQUDQfNwfq
DUXCAQSzmhaC7FnBEoB8skGAUwW5DZy6Kqn7WiBL2WtGzxL7yCZXfzwPkkcOB+dwpr0wjEWktcf8
RlsvemHe1+1YKwTOFYCp/Tq2jwKxkukbRUeahAOw05iICuDIxUWd4Vjjlfx9t9LrvuG1bqjS2WKZ
607kGk+OIYfEh0xGyrF11LcgCxQBcC4uzophlD4trLAHVsQobkAj7dAIMdoPOwIJirp5WJKzlMka
5nms63YUsle8JFPSBFzzoYDCI+bh1r3eRg4fGhZq+p7v2c5CjGkEjE8wKIi5RVOSsOzE5Yo2sBKq
tciVNZWP3PRNDB2CpcjP3cU3Y6K6/uQRkVaThaKlgPtz3HL1xYpVfXejonN6PpZgOl0f1lvOE57k
KKmyQQAtQydu+V6Z/4IndpAtvxSLMzbqOmlYMEnWq+pVZKn+cwOIxH2c6yNxTRKQAd6o9kWgWPjc
oI4pZj797YqxfuzVkBGk91Gyqpx5lgLh4M7vyW81p7ZK41IAfQ3KKfiJcXCfHMK7eBfTQxxubKdp
4MZdtQnRpPyUGVZwtFPwLATBbMl24m3rbwa55h4MtEiSzHg5ajzzqOVz0/QBoI6R+LJ0S44rExwV
Rg4Pvce8G/QttxqjwALx1ffMJl/rhV+1peNM/Nj+nFqdl4UQqFW33DdVSfL0ENCdDluaKHReK2af
f84qfAg4RE67L3jHxphcKoTtB9Lv6jykHpy1uToqrOnNPZiGa1Cmyyh+v5vnucooz8TYIAaNALrh
7tm5SkxbWkeizy4H/gPtKb8CZ/rAtQJOf8AkIlK+/U3pkWsYy/q/VdVhgKriBvAdequFa9uoyrwf
VZWhM2FoWF9fqSy31Ny805fvDiAfYiF82H0mOTYTwhtC2Ee2ENCV+XL7uN6Eia3FtbMay2k8CdXZ
E1XhFwLsV+SKnMOMtF0JqU2TaQRyy78SlljvBgxfF2M6CuRMCtWEuq7/ey/OgnaDTS0A7dWV139R
uLQHtaiompXqUDelvph3fooHILKJfTzs37QFXhnp2nwJ5nSolSZhZkzOkdPy/M/DzfASgkeF/z5R
7UwdPrl9aVUDpmTRiQCVstc2CNpVlc3DMIGlPLytcP8DXcvlAlK6+6I+CGM2/umnA3PawrrFaMlB
+9auzjpHj36iEsKeyWNLmaR7OnFEXxQYLZY/dUmxLeyo4TQkSVTobRtTF1QV7RXdrIsxn0V69eFl
cd0598L7MOnVsZRiQPKJh7SzHkzA8qcqJZpkET6FDnNXfN4PmqN3qYQnAR8dGAjyfSMU+RDurwqm
nVlfRuE9mdJkBSIo74OXXwk+ZmZTaL1wJSVad6R0/FY5u/uBSNxTGf58G1qOW+3V2kc5BggJ5Y0b
o2P4YdMizr+49RKyypMzzL/wyHl2kgm6nhZpff6QH2PYq3hXjrOe7xwJq14dubVbg05fCi4u6BDG
Kusui4Vx5j3o2XGa9Rc8ShRR/8N89CfEYdTSRwC+gfdFLPugU3Q3Bmpz0ehNO0jBt2xbs5GgASfu
2DVZc3eAjzthBFYd0RYe2HG63fI7KZJqdwlgohoH8sQEC9IABQsuRwrCYVKq+jh+E3cvwox+3tf7
EZ6k67vYoxLtAj5bJrGrq1UFSKLI8hGdKQBeP/OZzJhxqgr/H+NSH5ogmqZs5DP2U9d5euM+rebo
uXnOwQ2EsWVNcBFvqoRiBkb30PyzDCbFMRCRo+aMf6H9T4lbeXnP1gHGNzNXvetKzGLGdovg4z+r
u2HKwBUDCbqQuIG+oLaiq0yfGhHImkSjGY7yIWOhag3On7jWE8l50NSD1uClCQgDybKVOk4rj5zO
3m49NfzKKimTmE6e2Eci/A6jYSQEnS8N4YXAFmVABoi71XoTXIdBWYblxAKPnMlCorNHqkSNrbEn
j4CetYTfGRpbbRxOMoi4KbLr8Ffz44xSjfENuIwSdvEXVrkAjNMGLEzbOEUku0ANYdxekfC9eN/u
XhzdYTdEHqKmE+ckRDr0MrnDrlw6AvAFxFniMeG+/jtenu1VgpD+WoVlzBquhNV3JwYaohz+At7b
U4axc6x9gowsxMlgmoxMzDEAsVYbyPCeCuNXckBf0Ic+wBUzbhWqETwMhhpTEYcu0OiduKFfIgL/
fo7OMRnSHtHVbrfDoK5K0MRC69Yg4ArNZFcvnocxRwJBWeJYivvSPNl80dNIut8zLYliak3ef3pY
FTwlI8PpMy4rQXhl1cGUvmUz/DqJizhHiP7es/75gL48GI40juStD4cMugtkzysLtpmCxDi84WjI
UZlYxYCN5I0Zr5xmXICb3rHk4t10raBSZykTBiiV9zFE3czfAKHw6zaSYvSUna1rF2D0RlLCjk8L
ta6PGuxTz3y9WV1gTWgK9B9ImZY08lqSETywRJyNeZGxPU0g321N7UI1KtN+wOcwHxN4G46WGyM5
XCK3xNXE927VZNkPkaTYjuDO+g8gFpRFwFWDxD1tabyP8ap9cekhNxoZtTlqXKpw2X1LyPCJoXtA
+6D5J3wjBNOjKdNqqjTbhRgpuzE7xuAtJNQ/uDS73LNj9X8Hacf9zOV3C+oky9uZCFQ4lEOy5zaq
9xjyH9S1qaz+mBq6Pf7uGDD6jx3ri04Mk81AMpSX+XbyG+L4UpPIM4vQhFxtTEUaAOYp39CzldoH
0XVTywvsru/Uz0rYvnvWwJ/Ck6n3ZSLVMDWRN7Py3y6AdSvBbL+8SXItN2IWJACWWU9Ppg3UiDFi
Sh3SfdZJYtFnhBIpgh6SBGG51D3S4qY+cqiktEgI7O71ZfyHjCVYMjLv8F5bIy97dg4Vajt1Nr+9
/AoFHHdXLcfq6krL++138YwhTGe9y4+keg8NXyc3mu4EcxoBo6k2CLQ6Phvzv8246vCqgY5xYLe9
77efGFnPst/G2+jqnzizS4+VsVfMDRp1O7Ijsejykcar/cELWsFYQl+sgqr59QDYPmF1wiGTDPP7
/3absSlYTyGSPWvtwlP213eq47mJFWvqYnjHq4s/HKJXgr/c3sX5MkNJSXyoEWZAFWGhnCrYTpu7
iW4C6fzBuN9xhG8nA/smh2G00o0yoa6PSWokhlZw/66hQ/P2l6JCEdUIcQe1UVYlSwaqzMo+5xnN
3EaJYnwnqkMXNVcADYJTMoTdhwzl0H8ErgFyTODg3EaZ9+uRfvRPhMEb8zr0K7UqvUfu3c1MvwNx
zUvafMAk0vCBK9s5sq6Hey5Sa++vMExz8o9c40EcwssZ5IBrferkCfemtE0ORZ3MzJFdhCYWQq0n
cn60OgawSdFvCjlLd47aLgv8nsnzxqsyzd/NBqK+D4DG60Z/8ZXDgkdQZer3dArXQEjINmfZhi9L
tZgsnv3QmQcX83OWafWtOrWoYH2zcChtX3/IpbHUFJBfG12pnZMfm+hzSpCsSnpSoR2OLT32fnY4
eK4VdHpk1cdg7v9g0pWvwVdGg3NZcdgw+3cSWXr2YUyIrDD4AjW5SOfHgYcQGRJ5Q8QLh5LFOmsX
TNQBDHkgsFbVQUARvCXSPmKp1brCXe1LuB0ENmkdn28l1yaKMkqs4/cSpbMgKymSEnYYFUPwp19E
HniE4d79Fj6R37/7x5xvOQmXJ+aN8GPZaJppjttkmytvxcSW0/VM1EQRBacehyVCZMnoypRBDBn6
SnWM8ZM+0WKGFDxZMdfemb+qpcPa9tlU7bXIclkj4IvhNNDUdSJa2mIWA7wd2aLOb8kTrbEXboVs
RE3s7RwqpziORE1lpx/Yv0kqlHNejZmjAtD0lOJMWB9ZahvxF/Uts48QRUvPlMmVU0nR0gQbmsdR
Xw3+j7LqydCnnOuXLeBIaS/JIgZsoNHkMHBinL4pfcMzUY70YWZ7xYLCXWUEg15HwaTOAmpwXvAQ
9sTrTVqAgKRuQIW1s3BDyQ7Gl13SutoR2CsHlC67lYAKS6KehOFaGVnahsPq2QtMy20Pdfrsj6UI
bfgjVylMe744ODZiAb3UlhnWiSZG3TOwymD2vu3GpEitshPxSKNWkElfben3TR7ABI9makdZYli2
f/A5f1EKFCqaaW6Hx05CpjMlq82KXTf3YYGWVLBHkQHnKffakfQB4VwZmdrCYsZoJ1t2ahk5t+Of
f3jyPyn2J7hsPfTC6Hg9sn1mZ4zkVvz3uNHJYPsfMOQ3lzJa2SEuJLf1F7BD8v8ozxtiQYD5GbFU
jjoNG6Sr/UEtTQyEIedf4l3yXZx+dbUmTTMWWAWzSCC7ADr1mWnoBJQ9dKfxnV/m1lU4BZhILgnC
fp4UGGfxvlGdF+RNmT8oNMffnLyi+NdJbnh8RqyMkRNgwlIu08GDI7RWFzaDHjQker/xpgQHpSqg
GQmGDYkvM76hR0u73ra/QQcgT1+9eaAn5ruj48RPPfpsiC7FA+kW89FOq6bKn5fG4wTRAM/RCG46
0A3L51sA8Xs4dtWWT8zUfcu4U+eDA6dVMk+YuMqUidmVIJG2yNMavfmPvxBL4trUeBacnNG1haQT
Ez8oZAQVynIOUKji1OedlffA432dnDl+Hn5h+6CeZd0bvc87vqm0Y0nOac9vAkRHMaE7AKNq/mOA
nL/b9IKNrWcwz4chW+Dzr9768bdAgeZrM7IqBw2cgDDYE8gk4idEk6xNW0YuXkgYllimVDPa6aOO
fEsu0hEaDQ8VrBf8sGcapQDdOVrOaHbJemwMkubVOIRXrko1ZKw1l42AMJDhcPuwtpccBGIYVwaE
phf/2cRSObQvMPYAGVW3Iaf4o59Y5adx0wksiTN5l1iMVsoeejHG6kRU4c6Fa+hXKo0Y2+duzUoi
Z6H/a+E1IzF/WT5pmqHBw+Jc9ImMZU9haB61ALhtbTUnM8HeyriSNyLC930yUsG8YgD05hfhPhx2
ldFBkOcNvAyWb8go11DK0zrCNwzYpjy2MwULMw/f0dTDQfBO5UxD5bEQ+C6ARz7709TDMf/kLJx5
iUquEnsCuFt8J7QXwiHVLVuIGf5jPVKxDVf1hpxjsIZbdd9WSW8QEDY1kxlFYCCQ7889bM2kmx6b
pBC83c+DTXJXoRPy35qzdR+pw4UO+V6Vu/02yu/ENt01Boi9EyCagWT/S4jiVxO4w4uvsUNaXBlG
WX5OJ9fis9RDNhsjrft8sodaK3RU0xJmMv1PkTrJZjxFr29oGpz/0n7pXCgf2EK3DQ20His6mz+c
DKzbZVm9OI6nRpN1k3pP624v9nVsl9YQ2AYuBaSwcfIyzPii80knSM49potPpO/3nQ1wt6LdFu1F
FsrQYD/np6d5IACr3J183+DF3Gz0xOOUZ0Zn82iVOBVOXd3kg0+HdxuXsQNWnxroVJMimmhbKiqg
ikFEviwvrX+LxyZ4UDeKsi+tam9wO3ilB3d0fHMbaX51pnIrd+n76oO1szkUeysh1nAmCbk+MC7x
0YX0sZAFiME9s4yQX3q7ReIyi47YHSep4QBkxKbVI2vUm+wX1hmGkq8WlE2VpEvyW5Li4JTSVYUV
JHaFf9V3Bl+s4U80n6SHkYUDQ9HYxtQOcGNVIHtvbiec0BY/kPdqjDdkUGKpPYny6hXJX5Dp1OtJ
ZtG4NMcMLvz6vaLz3sSSyKlAxOWmBJMUS7g6Q3f4t5MWO5jq3I346/rzJ6/lBbtvdydypKelNidS
tEFvTJhqI8b5qXy1SAKjaPobHzxPbaqZFrAcdWEotM9IZXEI+pmNa8L0Jz9VId1gRTQriW81c8jc
LCqUmqh6CEITanumH4a6kkTAHahhM9FxuA36IqnoiS6jdRm1n5Ufse5ODdJWpb36r898/H3CQTMi
KG0dBNmGijKmS7+OX25zZ97kbStDPTqaqhm9+2AOBB/U0jiqDybfQDopA2zUL2laUIz43QAQ4POa
uJAKjihbROGgasSfsKAcYC3dYdAITZYRozeowImTXjBnjkS9KVF9BbxWs3r7wOPO3nBYp/JW0Fcz
Y+e6O+72bnpzL3afQQ/1gIdYISIt0cfPDEj2qwzxetNrnRhAKnxvjPAPOYFzlLqGWa+CQ3Tdze+t
TqDlVlzSk9vhCDoId9RvVMwTK+npfUpPu7rW4WiUp+zzrgqe2RGmF415Mqsy0e0UA2aViZxf5t9y
kx5RxVB3xGn/rgf6cK3sPzxfSD20Nj/6jLCgn92kB06BF7EZF6HIiikptWC2T/aXis2miLKDyLJ2
GN94K2YxPWNANjK66WmaATKxJ6FOjjLoWWfasrCFChEl/Fn9inpoy7C+z46aqEqvwC6ck/hRFRxJ
Du/53yH22fG3hecLVelCZrPX7IsdB6Eq1dqQiuHHZil5aWa3NMqNBN79ypci9uL/G2+J8VDlZsgL
qIgZHy2CJjE9APlFzBILpxfoUIeWVWdV74fCnMCMCDoo/joxYZizsRTqu7OqzBbE4IU2wZC0hzzA
xdQBjzCqt6AwplkxlRAHwqRlFhhVEkmd1wbetG42O2418UgEmL7XRq7OwUHrpFu2YczEshFcvpPR
Gw+VrqgcrpspjGQry5OZDhOEJVa/ElHqucIudNZik/zwKWGCAmIcg9R8lZSc/w0irv2Y/nPa6NB9
7gB0h28eRLws8DcRCWD2oFDxUqINkmJxRtgDnfKM3peL12oBbyRYxrk42mPhJs9JXwxF+CL5HKML
MJuN5y2KBmPNbF3Pj3k6DmYxPOa7q73HtEVl1ur5N3kd3aCUR4jhaFNsrxRDL2sa46qS0ZAh2L6Y
X3hZdfshbGnttHPSHAzqE1zjMJy4rxEVYdqpHLYvU0t/rEEOrfI6gynUCPqvgwWi2TfeUesBkEXE
Mm9u4eZ8XirLNtq/eLU2WkiZK9x/xG7pMvMBGFtcMnF+ERoje52/UD7kJ5qBxKs+6Co3sVrZTZSc
v3cAZkOOLKkLNB+8UrMwppelqJ4EorJA5kbrnn2TtDCQfntvC3g3vWPLuttVAB3walzLyylYnFRI
irvTlICZ5M+EfYkkOSPcazdAOU5Q+9/3cejeoTCfM2XQamoHOlOcIDjwvSqIfFz+ZmKsnGve85R9
e/DI0I0Bw8Pu8YkEjSIQ/th0JOqMkdzr7NWpjbbyYzyE+/GP9OUtc75WvTPY2tlA0KfxXlRfWog6
KselETJXn1WWAyAhyP8wq/MVm/5rM1zHr5IBgx95vyomIZU0ADhN/OJrkiSIca92gC7xnSxV+mTf
Oe3Qh2vHsHe1iuhkbkFelEy4sPhHCBU7PPF1HBZduo0CEAFtPyu15/2zuqShHMJ3+nxsg4WKjrj8
jSihoHzAU7At7utBqIhsnxPwMgFmv7DmAbvMGTnk1QEE8+wJ1gls+GsIC4+ETGpQ3L/VwW1Ofs/h
oWZuGUJ3SlPXP5U/lD6DiD9JWtyo+2r7cq8AissjOx1cld3agIrksp2IQ35Y7OhePhUuhoRgtTgS
8eWMpMtHwg4TJdhn4pTWkKg5kVP/IWA3gXEadxRcx31/8SHQ1EMkq+5wUzlK8kDQ7svDFhv6P4rC
JQJ8NPx9QRc/649b7V72Zg9txcvuuGB8oPdeocPSKmFbow66MzrbDVWyIFkZ7V7v+dBftt7Jj8ai
hTq3pitX276qP149JBv3NiP4uxavMtGhfYbspku91m7K9uFBd9gM03iNsc3R83bCEtt4ucdFIcOg
KcPaER/AseYKxudjFKSMXS9/98KGhEhaP+YA1yWNoj8rdcptmFQ7UvZdyhHxTRtfUIUyWZHLlxBF
6/zSGtk9rU1qGSZw0BWQVWy14udmOHmCrnhpTOMl5M8+jp2sRXxJaZ6PUkVOJOvwgVWZj0mvJp/9
SvovzIErLLJEHKF/OnX8Re/0RNbmh5uZ8qNZexqNOlph1qVHz1ELaYHA2gOEz/6eC4SM0lT/+DxB
o30ZO/TpZmSlCSVlahLeb9PIZh6sMqHVdjhnQI3igK9fLAjMrUjQcueL/ZSA3tT2quFGL9oCWdmc
T4wqFJ1jfe4r2D/IMRKqeS2ScgLPTR3LWK9d30brHHm2KIAtNEd9DR+FBkTCtizWuLBBjIhdSful
ZRkY4HPVrf1vJjWl1ONmYCmwUNzAhoReMzdZI8cnc/4HkfdJ5BSwHvFjBom1dqBgRggBKJkDsP/n
+FPJ6oGJGHOLiHF/JnjNw7k+CRFJxrKWC2BayhhO5mlUSyUXTYNViDz29F+w7PjDuIXd1nPc9wlA
JPFff+swBAeV2+KeVCK8S2I3myp+zpfDnC48yvLrD/lw5Em1WaZc5EPV4Xyfo6BdXiDlxlco8Mjf
ir4MY2vU0ynxl4QxiLiC1UWevPh4J1dTWqOxR+Lyy27fQ7XmvvJVuVEQGmAPhRr0n2yWnUphlPTX
Ek6HvM8OTXBtDxewR9yDeU3yBseHVZxCWIJFpNgKfzgK9zdgw233U2y8UlVjxfZASUcjgrTMUxJr
Fi7/chJNDujvUgKFEkIFXWU7S+UbI2WYL0JOqU7CvwlzRcsjzA9GipDYf5C+wr4SRZHKMy1b8ozh
br4zeachumM1DLfgFX7xLG/1COYrUkfvHLvHzD1BgLVyDXfiZuG/e6+dF6rQB6y0Ml9DzfscMlim
bbK+b7pnOg5JGoDv7doyEWVNIlOk9pHDE7T4GomGAgqcqBPPC5zTiOUIogRh2Q2+5ScXz2LS7S3W
s7DiuWf7Kt95x5UWVZC8HRVRK+Bvbt41J50atCbL2rxaSmKq7dPw2864nKiYzvdXHsqX1fs3/9lQ
zJd/9KGDFJKS1MYFoiMjoCL2TjUuAzyxwPZlRibFNjxDpq7G9Sv+IZtpaHLi0tiqOqs9VkfXGOde
amy/BKBPIv+TDDrJNYQWgDt+aFVH5ZxO1P5hHTJK9OpSopol/YZn/807TL50g/J230Koz55fXQQy
s0xSanzL41y27HLbA301yMTYGQY1YnOPRZwlLLjoSTYnFN4RfKMmyn1CbnkIFhDdh0mjNLGjh20J
cfQl9R407TsDtgQPLhO7D4wf18Ao2YouGA66gD8Wtb7vUht0CkX4HggiYs7CjRAbN0Z9KcYi2e1r
QLEoWHvRbukJNgkkIJav70lVtbDCNaxxQh1VEu2fcw2sTJPwCW9cMRWAaEd6+6sNSheayD0AyNTe
20CJPm/WaRyh1ZewyzRWQCxPVwZTBRSvXum8gFpSXz7U/vvZNyAj7HeeVxDftFjTZJdNqq9C2kR/
pFUJtKTqtMybnpelzR6gWGnjQysvWCHEX0IcNFcOYI44TEFGpBWnLwrqWumPMJiqSUzwlCYM5x7L
v9H99RsPJX5ZNMoDnAR/mnl4AGB3TdOl0lk3yRrPkvWu6p9ZowdyQf8QtzyaCVmfa9U6PliBniUp
u4LgZvHWmf1ITsIt4weiWWTeisMJNURv0jOTpa1M0Wq1QxRxtL4LVg24rQ6MDUWPH44qvP2Bmv4r
JVg9wZakElraqFVRxQytwwzHIdo3KagxTms0bs4cVlA3sqR3P+GjcVXSL4sBBpidmtiSkvajXG3l
Jj3rgZ0ZpNmxEOyqJW4k67LXdAtifE5dHxcKVzvp/taIb/9tgrwlRSEYCJu1SLSR2eSYUNHA4jmz
c9PTIPeCGgIPxlD+r76Tx7IhqNyH4LMoToRWkKgGYU8I4ExA5TOavZ375vC1uklhI97OHf0CTtW0
S+Buv62SatYvUo37kNsaHcwgPbyOvHEPJfgP1eReUudfxvjhGoPDDVUA66mlDXxw1X4FZmzR21U9
6J5A1geIoKMcLcqNNrSxt/QwC/15kIeHO1KV+tM6XVeprtjSz9UXJ8811EOu9RZdNKFNJsnrGpCw
lUtH8aDZdv8JvnVpK67RrWNLt8nBcAcGUBSX8PpzeQGpK6Nhivz8CmV1AbB7CQFl0N3V8Howl4Xi
2DeY7RlRRr8IPr+XICHfBvGCxpjXdChy9PfBmtfTU2OB9kaDHpf+dxUzALTW729EPKRjgGD3oGcU
prhfAYRnnumHrJOckZW+FFkCoLhkNQI3mNUwpnSZoW27pLsVceTMSnw1nEnJwHU+LBuOGgwZMsQ+
tgddwSCGTbjhbR3AnPV6KsxXZfVczD7OvL4qFNel+ZyS2PGCpjlLAknUnjs3qm/Z9ZUBexxfzT5x
32acWs9dFpe14IjWM7djzQwkTTCQF9XqtlLFTNDQq+J6iYgvRkZyVVugfVkzOqd5ovDKscGtqNn7
Ryi95Yth/JfDmsFKq3HuIVJfgdZdrqbFkWYLymbJhDM+mhWMJA5S8nGa1J94OJO+2+HhGJkEaOLV
l2L3CqxvQwpUCMRWhgeNYqONniZOZSO6W6AJ9teZKY/lRXipuLXMsrQk8Aqvj0qZuQahFgpbQIv2
slb2YjPI0VMgBIevut6AvD72OIjRwUp2zwsfEFoQ+YcuriDyS7dTLEUt9RD83ClP53j2R5LRdIOz
cL0i3il0Tx/kBH1R+XMn6OFU2NpLvyA3Q8een/JBtrFNvqTxXq71VXnsqypRuh0+ddFC5gRAcFcN
gGcJ185TYMYL14G4jtqU4HjW0LUzKvKUvPnfUJozuCssrMlzAaNcCRUILWwI54pknIuwXRUp0Ds8
/DHDdTlKuVt+NTkI1g+JxGkJ/UkLEKIK72MbWvuutP7ZZ1D2PnePnJ10JgO3zcKFgMd/aPNd1cYs
85vBcoKkrn7e2ycGPusfPnCAExDYloYJXr9aoBZ6HL4Bb32VTJwouktHYd+pbBng3oiC+PTljeXf
ZQsARExS4EE1ju8thQj9ylpCEyngrMnMDKbagleT1u770Ui7M/xjNNCtqIT48i56U4pRYRAd/9h5
11pWImWzMC2UtU6KraXdSt1OHjBNDYB6IoZJhPPFzQP6myweqm/ZgDyCwvnJAF45CzRe0OZ+9K45
E07pjegAtqkLpVVCUZr7u7H3Ssk4H7o5DeAFtcO1OiogrSLir9hQ34BWX+74NmnbAISwVayp97my
NXcE1rjPcEaRgYgHdAzpTDtQsoqpePzHKtweOXJdL3q+txyupkpJFndM7x1rCL6jG8OurUCAjD+Z
GH0g2J0ZaTHfLK+E9Ap4Vx4ZHhKaxprSh5cHvfoP3AEFjaO2WzGNAey8+onCeQdnVyntMZdOhh5U
cSnw9JRJ8KKghF6BldACBEJK3GA44SoVnLY3fJ/302+hM5TVAFbSKIRXlfkLAGe+8MyPnrq/L0m2
Pl13L2g7DPf7YgXPf8O648OkO5I5k20MCTM8QIjIOeb6tgjtY8CnOVjm+aUGxmOEWpCHKt6qboyf
ix0GFOwT5pUrkWxjI1MSfDHpRIqUnaQEmi4rjMk2f47tE1bGi+v9mjHV+29QVwL7y3q2ySeq7UxR
EQiQ00RyyjLcgFgM8hrVfQIGO1dmOOuLSRxCuP4SRpKyQOoS5oKJO5R8xjKFwozv9kxUt3DqpFP8
K2FSfTByuBwdEXDekMo+F7MkinkODkNhvbjFg8tTGYsHPVmeAc6bzTmatwNeTm3wTcVga9zhkiM0
Jrg2lq4Dho7vpkgn7jsY30Qy9TtegzRbwwsy7UJok5d2fJwc4zs/0k7wPgFQnThGop2V3+BBY0x6
XrP6orpY27/tx1sm7TDpTVw0h92Yz9m4sdx+p69ug9v/ifJwSELdkQ6MfdymgVOY4p3+ZcD6hAic
Gy6dvfJS9eBXZaTHsvGFnYLldMlDvpgt7isHGHwoBTL7RLW8grasVbFXFLLcVU+g3vQr7BAIuHaw
haupY/j8v9OLdL9whuoEKZAk3HhMby9VPrvHVL4oRzPeQE2coKn0m2/E1rib43sPX1RBtdpEZZdR
PMt9BSD3n02yK2Kn/Iyrd4M8mP7i42tHvL723j/tmOYLu15aif3jhUkDdwD6Rc6Dzmg52I0qXLkP
Ftqtgwq/c6S+m558HhqDkQyOgRnyU+T2tkhVpoMiF+8mla2WvXanmO4bC8Jv23ePoR5IHu4i3V/E
w8IJIBLPklTZD0kX6EOq5MsDN4624S8XcPEQfAPTWE+kDsXZRd8uUu+Tk6Ea7P1aTjy2883hzuBv
/MnvIR+koe56MCTmLubLLsya6MwdMU3wmPk2s+Ss1H3RTFVtKv+Kc74rlPhcBKQv+cc6oZLidlC8
OBHuvJTEcbB22oB//w/1p3M27uFH4BvieufG8BQDgmBEQnaRSuO/dp7jGiXcSL9Tegf/pgutu3+x
HRMqzuUuLhHYvmr+idMfgLpKNEHB6m2hxg9wXKCiImc+E3kWmf+AeYI/SPQCBoU6AT/oqJlPz/Vc
3wboegoukKjxsPE6I1BqVkC3s4sVAxQcNdqBAtev9gP7m81cwA+8UPfrW6lTBCdHFvmN9zguHAJS
dIttp2ntr89M4QPyZzAptQGRBqTXQEXgRacGHPMLs8tYh+49m0QEil2szYFiAiiHRTTBF1TkWrLi
uJA43QSoaHKinj3dbVgRcXRqY3LTCvQEe6EEbCLLCC2x9l9BqBpPwsIHXVNNhzx3if0U80j3a9cA
Es1WHf6BfJBWjPzDwAI3b7g6oafThxFU74Wz5SsYtw+ZJl2JbonTW/fkfuYNZVZiRjf7l039RN9p
MtWLVkUM5Ou7iTjPwFEySlwJDP1NPleWc5/17oFQf4IWnVVp7ODrKvOoEcG1OQY200DXtr4C2FwT
1J0QQkR2JZfIsu1T859lFvRIIN/KhVyI/MRtT5oVYAC2GhT8+rP+keoHUycnCMYBzPvHV81kHrCS
KEXCkLFiqHZ4n/jqPQrhY8+KmQzCvx67deCx3CRINFetD+Q33pRkpkwy8XPJJ+mtHfVUgF0Uzs/B
aBMTDMbNiEwL4oYc/HUuv7wNBWMCJmyuor41Bp2KFWNfF3taptfeoFfimy2TDfmEJNFGwwpzRTdH
d9e47i/IQI/xI4YYr9xhpQMkhHBXFF46RjuKtiRqhP/3XIeNmnUe4bzR/ji+ehQSGMS75twSWK32
0upZVnkkZ1cTZP826NNiZMxdmy7BME3WU71yKZq0s0biQqo9W9eZq5KiKIGlqe9CNqFMLWYgG2S1
y6zuGKC0ahAIr8Zx8gJt3iC2hB02vcwD0adMes2qsdXqTP6ocsDTURhv0dnLnWoLtuTLi7OZa+Pc
D0KE021HvuIfRP8YIv7jJ0//eEbKHNLK3mGRhXhl7PLNAeITTQYBjH/VPdrvLidrrT+pHDRCd+3y
SwqlsdybqJBva9///je4PNkOj8Jee8XTyLjz9D+jE7i/W9gjCjbARtBWrOooA2+7FjhgiWg5jH7Z
8Xj2YrUQQpoYtBFXok+kbURWCiz2mQNTMbud+JhkQ8Q4g1W/IflMqbMVWBRpIEA9PDUpNJ5fusU3
3FD7BG2Ve/pzECf//zdhtQZP2IOW71794B7fatnm001xbR0zdSaLoBlPAZeP+dbCUwiTJBRC+OOy
xpSw1e9W55mw/MUDwHUolnpRWfFfAbQlnUqKmqMwH8a0+/TU6nygdg6By86E8K+HMCUrkUz8URyA
3hCMEbcWGF+KLGoKKSZu9mxGePX3CW3kw+ge3M9FjGT+Wu7FoELTuzp8w/LonlNH+xpkmLeBqrhy
IJrHJBLvR/AfBpMURFqzjx9iYoJR7hvI0OMLPMmY1BlSToss7RLwPbyjppbEMlY09tv/VnoPXX32
610vofSPazYNb6jS5t64kqvRJqP5lPHLdVd1PHpkS0cdE0OYwlpBlAV72Xqd+BC2zUmxDqwsUr+q
Fr/vSVLySz20rC/3vNpb0zV4mi/dbnY/KNyLsfyMJ8y/O7Zui9fUM4igUWES/59bOxwdRz7acYmX
O/MGmO7AKeSYPjlTXFp7nlTQ+IXJZBnrTaRdDv10ZesDrqaeAPX+fsWnqPrNeKqk86IyOnzLxFJT
cyAh01xDyluiy6AbWSgi3GPMAhixQkxVPAuMc9BjEtE14jCOtuhhRiy/HFd3B3FsNsn8pgJa8s/+
ETrvpzpJXUP92tDWZ2X70bdF73heTkS7a8TUd9cTr8P6BPqsA1N2plT2FNfOtv0gakBb7hZf6zGd
LXlDrBoKGEu/aBdpNV4FFErfmnFdyijaMIJB8J7Z3YJliBHOz7YhkDIcnJmawiDAIjzs2KRUVAxq
kT7sww8Kg47bLmDQYuJCcFRc/Mn3Ix+bhISBQjJITq7XEZc5kDUMpj20Ng0Ng+mFyGrE2Wdu0IqM
DlsTbklXUKUROHBX882uyQmPSornFSxsUGl0scV1OLyfpNrFdfSssnkd1u5QhLAPm6A1yCEu9mBL
/EKkLCqVhcOfjWNG70pDSk/6BFmVendN8U7rRpnF8JsLWNG9FU/D9i+guANY+ojn8XrEFxNsiOXc
lNvbgnp2ojOe6T1cLbl2Mao9WV0sUmBU8q2LRfATOL4pJuK4Wfh199uOhC0FvUPL3OXwOL4GMKPW
6T7ZXjwpbGAHuqlJgLvV9Ynu8loFgYA7CMBV0VRQpKv5G38ayjzcDGbXYxEyzT6S2AdawJ2ABmf+
vM9vTIEeRAILQ+KeoEZPcv/0n9rQL93OMP5zfndP1fZ+WBZ42050vcQsA4SqziqWkj7cqVQktSb7
xGd9n18SB5l84eM56DHpS1+lEY1opmiclYFNcTfkA9sOnIWF9PyjCIs32+FiStNMEoiYQHCycSdT
VxMaF0s9INY7qRMx8AzzxpD097DA8+zKcemcF3/8nM+izVKd0Hkj1FsPmcjzxMMIReIdti9Qfkii
M0EApfvLuUYxapvo539caCkE4hmvFMvE+RJ7TDNWl5/R5HPMPALrFxMgVDDI2mbxekZ7Wm9oxtv5
L631mqf6t3ThfvUi+XzbY30RsyQw7LDsq4gkklOXLDiJh9VUSU5bUsVYCAmrNyte8OvQjxbgcTNh
Kv47Al0IeQAwtTPNXTnmVe+KYliH92qf5+STAbbdYespiG6AGJxBZup90tFzstaBmA8u9HfpbNd9
8XaQPtjpRDKfGeUGmYrjl44il3cQOf8qIMWySsLN6ghJlsciNFyCWnNTJzxehcRz87htUuLac5V7
f4gzFXt06tZYofIWDgqF9Xk8ghuywboMCla/nD83WXJVLPBeMFUYDunDsOvnNWRJGPgC6yaTyDOa
BhnznCMLtrB7Di5AQfdhhwUOOmKeyLIoNrxvGljV+p9Vj9ERQHRNE2GJWTLdJNcKPTXkxb7Iz0Ge
Ainr04IgLdmJwzNrbCMe0j4uw3VKkFLOOtFPqjpiib7IBW5lURLN19buJiokr14/moazdwx1NdoS
OXiokLedePOwH5BNz/cOYCNfpxcPFzH4WC3E2o2+A/ce50hm6ScHK4VFGHOp5ZAhPcUjA/I3aoiK
kv8RJDGwF5Xr9owntsr7qRbMxfmt5/Wg7r+hz1oRTiGgizdiCsQquUy4Z6AKpBjtBTkCKeI2qJ1o
hkDNuBdWs5lQhvo7O4rhQvLWAKec4uliyHmoXsKv2Q2O70vNHql2ythiizqmxzxUVFGIqozfS2Mh
5GL+Gd2YY1iODhHxPn7GB5+SAJ6f7T01GgdgkfpGNP0jhD2Ku5rOCSAgz8zYy4QAbsgQQdRB0IFv
0Rx0aA3OrFCkQ5kDGQRQeM0Bfw+KCgmgeCW6H1QeuvOfhhbvL4JXOIReI5HZwxnoiP7NiRksgy61
LiWQfkWZyjS1OsNN62nJtIE1PifSEI1Y3o0r9fRVlFQTxQ2gJSVXBN7HUHyueQ3FzWQiMnVFd7bJ
S6Yg/Bir4SCKgj75DSuzLP5fQ77D3FnAQUr134GxC0uJoY4mPHQMrWjqpHetktp+62ANWMM9eVsA
OSR9/IOfFTJ07fiiwmaBevAw0yyTyMgFSADUnyvZctEnNvqPlKy6wSUVKU+NaMJQJ7jb0XTMhsBu
yLHIPNwTqAno+8ukhQVqMnkfGl9ulsVgts/O/wTP0t29pW+runGqqpgjosT0nbXZA98O6zzoITyy
If/w2BtNK08J+hmLj/VnsUtHCCJ3PGl1yhSt9fF2zwoj/SHhFHym/hYyrxkCBowD/TJ9r6E3EzU0
r+OnHKtgLk3A5CHki6fYOJyMtgjUYiX4o227Ghoc0E77k4z/87Z/2ywc8mlGXaC6CXTiIiH2gFaC
jW+otX2BhcK9PB4GZfW6nEH8nUEeK7Tfd9h9Nq3yheqjjxdDUq7xe9wd7Zx5JctB+MqQBfssrs5+
D/cVrBy/fcX8mdlr87eWQ4RvYwSDmHnkbqwfIGEx1tN7oF5lPhOLhPt+GUjeUOnyOcpm6iEhdcPJ
qWhACQeFGnbcgGWA+i/6/NF7A4XdUo02BgFqVdZLU35bT14OWXD7netkOBLKfYw8EhhbNdEc0kpn
ajtC+baId5hSz5u6R3gebmi9YPE3dDPFv6pKAPtiaz1qj7/toO/qHkD9/qnV2q2R+COZ8JfD8arj
eGQT0ZURWpK2XV5SxXumwiZjXJ0uEiuTAlNj++z+X1J4HdyrsYdj73unv9t5VS2+ge+84wdTqdjQ
YQwwbPZAdIK5dJRby7C2ZNbUEbyIsgvXb7Wc+PUHdFr4YCY4lmzdCgsC5krCU8BtwAP7djbS/Tfu
tR2uJA1O7F5YwsLR+Frj0M+i7IhbT0wAxtq+aLBUcJI5R5GbOSh92smU9cEPFG48N7CcwEHCHExx
ACeMGM/3C58LueWotBLDCcSKtT+W2b6PzpmNwxKXTKxlWudBIwguzIbXjN3vtqDkXE5Ie+3MISBG
Ay8LIC/E/cMm6l7GwlJ1cBWqj+B3yH0lN41Sn4ANpzYMPQJu5YxgMhnOiy0VTGHwUIOT66pabCms
FLwnDybfcuPZuiVL5EQ6wmSLpQuKo4UMrfcEmHc+cWeAw1F9mtVgahll3N4Sb2URzsW2ZdGfBX3C
iSaz1sg9q2lbDY/+7cYqMyOVI12+BBxPVv75RoF0vHzbAoNwsbbhQqLsWC8811eFbAdsEI7PUNN/
6buBih2GbxKl9zEqO8TBQ/8xRd6Y7DzoYyx1/kslsVg8Zmror5hefmxe19pxbYEt3WU44Ea8krls
1vJK098UQin4Cu06GNMnvq0xluLrA8iab1Gx058jC77yQcfXm641o8QNlEysKDpYKIflva6jCNiu
PRAKUsNbyusPt9P8M8sd14GcmHk4XRHLRazlQ6eZrdNV4y7pI809iyTnVq3hdaZzrqhr047vkpru
qVCEJKi9PxARsg2t4x6zuvjFqNwbM8GQbZaO3yG4JKY6Qzm5QUJhglCM2Ji0p6ZrXPLFcdLjQXu/
LzKz/404BS6Kc87Rbp0kPQLjJEUgsI03bef3WwIO8Arh3a8xGdT3edRCb6yGtoZRRDWbiV3GL+Hm
hAs/iL/vIG1x/Lm0EzjO2P3QE5vUMwTiJBY14cDh8WK2DUfgt2bL6sx7IrDJTX7r8ug/KdrSYznp
4rUYHlRnDiqHMKDdd1JeCrHYG74NPdGoAFy+sBSevUO9W/GqU2l8t7DDg+0ilqPy0ghSFjLRS8Ig
qrWowM1TsgYbde27rOBMaUpFGd6WrZhihng6VKzEU3LoG+hRAfI+MkDVoczXw27950tjfLDvSFL2
VBmTTbbdxRW5jLmGoBUncfFdPOdt/NHY3ceJE8huZEQjsqEWQrDu+WsdQqwdIA/fWDbwYPzRcYQr
f5NNTDk/DigK2u0RlXPm7F2pY3l4WhW5KaOwD+UFAeRQuHHRrMURUvqLcqZvC/P2i1bvCW0ZVRvM
AAnsV6IplLOhpd6BE2ITdSZ/nEePee3F3DuyTXl4eNviE2YMNb88rRgl2AUFlVFb2dvrBLZ/XBvI
iaMFjtsThHQPG7+9jfP3bnm1NCUSY5kztljiDl9B7mtHrBk2YdY2anwtogznbJFwBpvQF1k2Ryg7
Ec0hoNv2+Ctr08VOJEKLUk2Pu7apUEsniPWsEpUIx4sSpkMLddd63LZQiJIjNjkQMm4mpkJSH4+O
eK3lk2KDSd+odBgtxEE2IIGq5zdmJ7mQgouyVEpWUy8z1ogti3btGLH8lqUR96GAKCEGkuj0uuhI
BMsQi11swKZEa8YCZ6nFDZ6mR6cZlu2uk73BXf6w21kcmLbpSj/UI1OoGMCwopodubDA5NFtzSNj
sPdzRlMagosw01OkzwOhKV/uOPpU7KMJmsV1amad+CHBEgunPYOxXNI/18L1vpbYLW9zJBlOemN0
M9GooXaftCOmker8Nh7aVALNX6xhrfVgrWylYx5CUNBIaUfWiCpRsN+AYTOVepwi5KSKcP+DOrKB
VDt+iYB/n1ecYsssFgCc8xojvaNMhsDnr50SINW3oI2hteqKYfoFwTx0yzC5nGBBKBeQ2t60iZa1
wTSNIvV0VqZ5P0APeyMp7uu9Izt7T0yw20pzQ3qOLpMGJx2Hwd+5wMTWFhrUkdlQ5gtLhhfjwIY/
/Z8V0CknW6uz0t52aQxX49YZcANMvuhOHwLqJEKCg7XbXWrjNIPEQxvx2gzVEB7TKhYIYCQdaFk2
bgw/QtgxeJebPZMSQsaSEjK0qcP4K7R5Z6pFiDKba/AwEW+jn7U1o6D/JLfVtSIPmtP3As0DSf0r
YeaHz2WwuQlbdPNpYtGpd4s+OrCN30dHgDZnkAbjS7Yu5EJb7B2vz+kvlacOnq4mxjDLyhgqgQiG
3IFmfuh6Ql5BQNst2/HKwwLaXljIhplz1iVWQUSnUMsNGJQ9tpu4XgodaGtX8+QMrNByLm2RwKK4
TwE0d6GPbi7BtR75hJJ7rftgJK59AeEY6KA0HSQ7xHiUPUJt0wZJmLtjvDFaKWL2aXOPxW0LJok/
t8zfhjSU4jVbhZyZlGilutVcvidffmDRS9FZuTbhdgfeOpequQtzn9qx6EpuERFsLjX2+QEzfc1I
wDgx5GC44SoVoCCWZXSdZQ0gfAViELQoqPbvLugHDJNV6QjNGdZvMnahu1m3V3hJEoiPkvzQTs8W
mdidR1qzP0Dr8sHFrviJ5uCdfhb3wNsELhX71LUhdIQoOKH/mURnEebZxxUHgcZr6v7ShnmSdWLZ
Yz52DyLfKwgDq+tue9T4z/3vi3CerGtVsXhRmcECiDPJn6izD5LK7GfGMYCHXXhogQOK8iBGbklu
86k7dP2ACHjeDo4YT6QijykQchFg00qpxe0PmqvJaTWUbdivTWhMG0pF8R5evM3yOiR/E2bBUcxd
TS9jX75+YXaEAyjQw51T91Bkn1ToXsInyc8i1dfcWMkQQpAwG95kb6Z/09aO34Tf772tvz+e8kGr
ekcBSbpq0LdqmIXTnSwN4zf/IF65zRMqVjLsvOTUhnb8ETf/9P/4EItuyn/HOXGE5rrPidqmjeLI
AMy99c/iejbCTycYhYDlknmP/ZhAGpHckQjEfOph0UreSIR8PcGL6E2LmAjIPKvlAIYkz2Cerrkr
dnWHzpAUSq/bIUF2pm2xiuFFYMjOthh4vdzAwmR/eT/nqgXdM5Ff/QuN4fnXH9LswilRmMMNpw39
+UtRi7+NSYITgHuLniPGnIgYxfEYpdf34OYi4U9ctePnBNUA7t9ZoKCtNJPYAL/ahavUi18CZMVA
UtOE4yqM99jbaNZl21N3kHggmBiErxdwZuK/CCkyMJPKbQmOuPWrCZGY7y7rYMhiDHtzaR9yTdq5
L1V+HEMM4I8OTLmhpsqsgfS5EXc1zb6yUtEUWMCTaoQYHueBQYIaj/lcDFn1vr9hiYvz8Wa6fUaU
zXQspZp7Tu5RbMtihwmmuzUu4FzablOAytd9Bs7fr1L9QZdroAgvmYYE71XBoGUZ3u4W3ylrTDw3
855kxmb4NxKJ6R3+rN9Btbx6xZzm+MuRErcxpd6DKpeovIUUNRgYbjhrJvu3ZnVyEOWNyXm1K3vH
cQ8y969gOoAYVNQrnwDUy8AWDTNe38VjWXnMrX9+hYBtULHwYDoChbJfxEeCLN9aqDouMaB+ET15
jILV983+Y0G5bfn9sDH7SK4Gji80z9tG0MctM4O7/0q9Je1PynYhpTgjY9p6gECJFKRy4904RNqr
y8A6+01bLA/Q/fKO6ikHWF/DhF7WHiuXfq6otZUGNJrxA/xWU9nanni7QKn1qZzxWwVSnHXMiOat
HIF2AsLUwZigcoFZDxbFvsuAsoGcRqlOUSLZxXdWwAlTskxKIi5yIDIumvCF/zThDvseOsTkit6e
GmCBI+yIvsRIK2KVUxNx3KD5IvMZ+gBMlnM2QpDGJNOBmziFgBu29GnnnNbAQ9MBwUBOzsR4BWx8
VbWaqXwp21rFO8+m8by33d03FxK2bU36eURcsMeL7fBjTMeT0UzQV1E8Bi6hK/JN/LrqwydWFOVB
HT/u5B1hxub55k8qOUnMptyqPrLF7HNnEEtjACdavJXgfjrwgmc3+MVOVP8pNMN9z3hH9g5tmLsk
dlK7L+V8yvlQndjlCvAr7vJwITXI3KFUOP/L9hghd15jVyNmgEL1m4Is8hn7yDpavj+jzgJGk+bM
/cHW0jm745yBHvAfSn8SD72Q2c1tJesyM6qsBsXwN70XyFtX7Uwu2HWriHOjClAqH/ncoLUGOuEq
tnpGr3gjdKgbIddeJAQXq1mSm2Kk0ZbuGJexV2zruvbIK+0cknUW61NS+Fham+tJTiiNO1CsRbY7
eSAGhgg0Kc3ETb1+JcMfbnpbl7Snau8MjtXByTBZYNpbmolrS8PRrVPMCQPEg0r8aWLQuxyYyHMY
dKimTNPs1+DxlcBlBMP8F+k3pGLIac+J2aCcRl+rZl19FBDZoIUPkpu3Dg8/8s7Rg1Q7ReU5Hpqz
PIEaSnV7Wo1XNjHnuuc3vC/6zFF5RDpcVp6RDjTJu5epvYIYeCsFnlzZIgNB3/h0bPQgBFXnQL2m
LUVVR6iZgn250cKt5oL0m8X4LhQlpVnc58cPrx8iwGk0R6K9eMA4GkxdnlBLxASkvDPFUSiQalUs
g2FdgFR2VkghMzz/ie/JdyCCnh/a3gOkX4dI5rJnHd6br20WCtjx/woklrHYcHE6kdRdXOrfANVf
qVOOCvbmnyrERTUPdthTaENJ6LuVgN6ECwinPFfj1s4V9bjx3L4XKJ9P4iBOqNiUx+rL36bg+SMU
40zQ9qmnLifQSHjGlo8OFhxgmsbqsl9ly69py6ZWQOGw9mCh/ktseNQ14KYHD5j/yO+PbSaNHBb/
VOCVBC0hJCAqSscTOI81UsgxgazqaBuxOPgiCN5nZmQbl65XaKfWSLCPcGgE762913hTHiCDr5vo
Yo5KIjP9ZmrkVoEgDzIoa79udvkLgEaOUwtisyktC5xVA1SSdnhfklG/CourncYNtjFnfX/5tC1g
azbRCpkBHNOTvLIeJOFMw+JV2fAJuncNU0RBR3I52gXAtc2YVAP5+ClatdkRzywGH052zWBUjjEz
dzAkmAjlnMXPFa1Q/fq81+eiO7Do4xB+BihzCLC19G3dNSqF51Tnd8PRcjxlRk0LpWQiBMOnHs/e
ku3JDgeevtevvmt/bAsUrbUHVteshkNm0hcLFtKI8ju0Sp7tLWamxjskdcarKlbDVCm1WarMzYPj
w27VvnEIA1NUt7j1Yrtwn3WdkDYVY4XeOrX+W5qsRz7wZXWoyzINPzv7b3zXfwKM+lk+CZweXcBV
4PHY5SV/IojiXoUcPRU1Sue8UmLBiHmVcMCxx4eOqZKVG0K1L3HidjkJ0+Q++3PRhbgug2LQKKjF
VCfRLHYanUWTrSmrGb3d/Q7hAmo83pufpCXd7twyOV4bg6heGRAFs8uxC0hK+s8HXp8DeLC5s9lk
GedA6Ojx1DCcqyT5oh6QNpBjRlOe2qogHYTVn81v5dp9GQ3rgnmwWhGd5EBWrWvVVRv5fTMV+M5b
0QaHoPoe3DOJ71jqveNm4m0LUSRE4Rr6ozeUh0AQJLE7GCvlj1bM6KFTDEDf1UZ4WWJrbK/kGstq
R9m91SP9YVqWoI0oZP3H1g3RWnn1a5bTBSBGIxVFE/TK/KBg6crc89BsuKNhNhyMjdDyBWHIVcLb
roIwEJVMjn0CyCuEol0F0JD3zaLgC/fz6NnJBwN+OSWn3qo3Nmr7KGD7QbDva3xeyBAAjmbPSYTL
2yjnFjJCNm7dfccB5aynJCk5+tYLhZ6ZgvRPZZidBjC2y8/MQ3ZGHzhsH9iIlUnY74w2CUzxPsIe
YbkVHcmVdgcSYZotx+UpghwqngMq/SMeJdXFFqrbGUBmqVNEYhZSOrvDygIYnP1efFHW/sfWIPLk
4qUvGQ/XlEj/Y+j+6pbgGCTEvhL8wjd8x9XRnJ3epwPYoeV8m4poe5FndeQ5wL5fgsejRD9bxPhY
N6xLzGZ3rGpK5LwVdaKiHf9/DZwsDx8cgDCg6a6nWoN9IhmF+bhOqWuVzum96jyUmd8wKda3UGw5
8jygaPEfMPJ9bO8OZhEtx6S2H4ZTKt4Csi9qVijmoa4dRO7rDBH0URLFjI4zc9TWR7MM5DfSdTE/
JcKM8Sl8tORZG0CJKwC+pJZjwDdeehmhVWaAmOuY0Fb9d0GGwKx/9qQAIexOnZxmaber0EsX/+g1
ej0CWuJcnBOy6s24PCe7A66INXVJgOHUWm0V7pqpYMLr19DU57/wLM9MF6Ev9TXdiGeUuymd4uh0
x4VE38owd4IOkFzzVyxYBBCaDLVArD4RZA4RHNdSjF0IYGNwM6Ox5Of45GjI3b7XVzw4E4LNfjXN
YMJoeEbMiPnVGiuyma/9YUliA35GRUWe1T7OxRu34qzlR6YQmI3+PalZ/fRQYd7WofV24QyDy92j
tOr1TTIlcVsgWYnH1i9wWLuzsv/Uq/nxZDjieUjDtX55+jiB+jcoVyh90AW7KdR7VDNWoAA3/V3b
3mwRMeFDEPEv27YUiNIrnrOKBMf3UOC2oyTmlhpEy+dwnq7IGEVkLRoWYm+XPIUI/xECDh9FTEte
SSECqqFVILVzhQ4tkenDTFWJUg6vVKO1ZaUhHyAWDVn3AzF4X9AxPZarQi9Z0JhOxaLVRHwW/Xo/
m1nMZL9urafAqEDXKYlRPegO3xM92ImZtvr6f7aAbZfjRXQIkDuD/+20WPR3p56m37V0Pl1Eih41
qz64jqv7SvDRwipWoHrcZfeRvD0GM3TfoOHlrcoKklD88g7csfFKftJ0MKh5XqH3IghogOU1PXVH
1pHKrRq58JaRm4rAYcmRmEsBS9UQlZOLcqPoUym6RgffERdMXG/25whgQ+B5uRnxriLBkR4PgjyX
/AQkKYpydtCF6DZYbi+DsCGsRv4NI14MS98Lxd/QUB081pouCni6o32X8o8ulVTFDI28HAvlqEQN
lRJZhHQLlomoCB6AHPp/Q6qDRyFntWCtJ3j6KCrTiYTmN1fBxiC9NidQFnp8T/46lywzfdiT4TQy
+XVsWI349BaaPKjLshhkaoPB83gYDgb6BX2BNslUhfdQQPeVZZJgPGHFTqiBePDbRRN8CI0jbXSD
BB4sKjXu207yrOSVUFbCep4rmCI/Nzkk1yLuj6UA2mMpe5HlrGxyze2G4UMMUKFNyZ5FHLLZOcEb
XsE1M9YX+GjTYiPDt8v4UWoZCFg66RtCkWkwJ72XBSM3WtibonxzS6dArttN2Poc/sJO96s8kBV0
MyhmZa5wTkbN4x8LytV0cI0Ewe/A2FasqInGMfIhzB2vKOj5B0f1JqNAekWiH38uusQXtB4xs/h5
egjwT+f2veDVLfZX/3PByRsa2kPdhBhHS7oayKAMLsH8qCFCpT284IWQMxy80KKyJAkGvSJYpfti
N31sXU9nBL1Ttt2g9jhMjvYaU3dIQ3/OOFTEr5vyEyt4OqFnhqJyPDuT5AqQMVqkwegTLYPkkkKY
c5nbDLPlpUde6C5bMFEmFRcE4krdSHUkZibeTWO+4s8LCTZRL8lnC2KEGl0dZj/XFzo7aKejysUE
VY9/BP+tzYgVF2uzDCeO1M45fwsWhLINdPzIiuTIYcoRnYv7nQpJs0AmlMziBoWNbXxyCpzth3Re
iUJNsWuGplcPA3JKhZQMrDKdv8RPzcyIjtY/gFsepVslsnmTP3ET7y/ghWM8kz8hbp09ORbGFUMl
eqcwnVFUWrPtnnQ3xV1VD6ojaVc9neGXWqBaMj/8UfVqQ8hGY6ms7C83XykrNWinEVEiG/kWTI7s
cV3ZXvf6AkOXyl6JsF48cxZPaFlyy8JzqP5mi+OexnpM1r1xqmeM9hqLSwmTqIGU9NtwNZhpsSaa
Pxv3B2uM+aUBkdBelRmk9f377k/q93Yo/HfYPHMFzecGVgT/W75LZRUaGky6boMY2ba36skAg6en
rzH6w9CmjMMPvR8grMyKFo7ly8GdWqAFA6rd/hS1VRnNPbIy5ohgPHS5/qaweibNoY+lLek+Ekhu
cbg1K+9W/MegLYEQ+EFW8aXTMHKzDATy8mUXCxcsZkUEKL9daMfX03oGOkeM+Bwvub6/KSO+DH62
sEkXc3tb+q2AQk9Z4NF5BWicLpyUcJxu46XRO/PUkgRSSdqAamw6rB+0NnZPqYJln8RP8wd7ZE4N
L3OddbuWWYJq7MgFt0JnXIrrvQZ9RYidxpPG3JpjGHA0iua50183oCDYYHeV4m0AB9sUdbP2qZ1j
bAX8m0PHtTPBr4zIqdmLFEincuBjww+yT6wFZI2PfX5TR86OF5sa6G3jDLWuiKeLq4HLQuV5XCzh
A9AfYdq5hD6xzOgqarPG0yRgwJ74UqATZuA39MINyrEFygaU6Y88zKLWyO6wz+8V2fGStTwpbcqo
7vFM/qNOEJTEGuuvavXQua3U4JFomnRpEx6l6LAGkMxvumgLfCjjZrjDSuUivGz2y1FZyRoAsNr9
G6jpzB+W6jk+bFN13OmAO3tNoVHXqEdX1eumKfOmXWfi8j6Za6IT42SKdB7HA6/GvS/Lqa1UasPK
LSmQKkLTr1PHD69b9LVeLjmc0ke4sZPnB02e/QCE1VhfwGYesnlYJSiWDfAp84Xpyi7nC+u4hzQu
+jO96T9IxokHGiWa9JRdfNtFMsstiWHEeAzRdNjjSxoTtDBIHV19opN+/bUksjammMgvHR7Yt7Cp
BoLAhR8h6I1nOMFbEtK92m/uj+P6Pw7e/76Ng75d0JQlQ1v7i2mV3HfV4RxqWotNCry/eqqUYv+F
Q9J1hPYonOtsm7tnl0vSy0DLucBoLdDam9RVXk4ve7sn3jej+I99LFNCtWGwqDg28uEsHGnJoyVQ
b775vJYiIXOWgW2IcoTL0UBOOjqX227pDVeILGHtAFrGcOcngCa/X5ML92+gXKjZiaAbULUbYCeh
mKP2jcv2SJHwlJ6k9teYgFjvnJtZB3MMNn/U6MJMa2AXZMClI5vvpHHy88z+LpnwWWLxTtTY92T2
ZP34yGxHUyGiXlH8kgRloz9jb89JCukC420v+ZoM4V2nH/T3SND7bv6X6k5V6TA6kvhQSWslD8he
DOMFzFzCwKMtMWQZLAv79wX4x32rLSLq53MsIKSVcMxOBbyC1Fk5fNGO1v7lImEdD0a6hbhuM8uY
cX90nBYyseBXnflcrIeiYnqm6BNMlXTmLkR1U1CBll6jzQmtYr8sh3FIS2HLm5xLj/kJ75HNahZY
6FD/9WOcrs2Py0a3UirKV0XAJIuoJUv6X2AASyfeX9BMyoTaMAQHDoqIICRbBmxE4gTnZY0vIVK4
8dgB5WKvQMd1BDfW68+wl+ljV5zJhUv7+Yg+gCCODojnToil4Cxv+TPPUL0DJDHySGOUnHLaz0CI
W4T3uZfKro23NvirxDw3Ofdd0E8m/m+Ufc+SJ4km1AnYlXEtB6m7P8tbbmWY+Hqh553OdxG0ScTZ
AVTk9KI8etW+QkqbPbG/h7DvCf1f6kxTWbZeMdVpkY564JYmdNfTC0enEiNsfVwqpuSE1sqaB+vm
G1vFvsjZie9mej1SsqCAZHs60eXtUViEnLyb4cTHxo331dxvoVze4pwotndkvgqNCbHWY++A+QXZ
CHXM6DgTSPMEz9R0WZ3PTxac3V7bRDnnYxOM1E1AZrWLyRAKivY66sKA1rIu5pZr9Nw2GOOVGM4V
FfxW48dDkCQnLwIfbXBUoEIQMK7qESr4KPV9b8llIteYB/bdZZppwaWIjaR8hPnzrPp50734+1Nq
/W3zoJm2L5Gf81wyG4ayC9+yfBb47klcXGo7fZcMi7zlb9WpztOTc+pH0iwfb0n4x/q93y/cuMq8
QrnP3Qy9W4QJ5ae2xr9QPxUYur1fSE3UsC9h3aUbxe7mSwRExjSMQTeneveTNCpsnkODqzCnbQJN
L7R4Ui7qcFLSpz1SGIkpAhzQlddr3XfqWli7zE4/g6IxzUGR+tTM3s4IeYHBmiatevD8kKsDJbtx
PEjE3rgYDWveky/P2pXjPJ19udvpIx4E/qM7h39Qc5kphr63p123AyzcohK2b2YNwBI6QhvJ1scz
lxoRhY7O/tdlomaZq+1vWYHln0TAcbJvCSIghupeTrOXeo90H8Xfz2MPi2VW3OmdGo+Bhz26bSQ/
znKhCylRILA3ES3znDdu2Js877VYthLUHML/bvNDS7U/84/YSZW9eFujLoryKaIuqJv9DP0fvKKe
Sx+nv5N1lEVb6JwuwfxiSANldc10MGsfBDFIb+BvnMM/vmQ1GNHAT6Y8cpvZkU7Ou3P8i286LZKr
xQgfpJ+o9uPzu4YBKb50lmUmhxFXAhQ5/9afW9+aRSpc8w27CGnYjNM0lcmOI8Sx6HfMkR/cgpqi
7+g49+n5jjDbzLITaFUzBlOi8SjLwUmo+oQoWcOvw6K8ECcU9VmDLbxN+rONovb1bBw7P0tKwqf5
hVt9/QfM55Huc9yK3MF8sUE04+m5G1/in8FoDX3mH1wiUByBnD/ZdxZl9wdqfEA6ARAZ2zMOkQ6b
pl92aK3yfO/OysuP8OWtM0JE3f/DCbFXAbRRylZKg5CHnWfNAVRJU932fknwcfd+a/wIRSAmc4zT
KQrdLMGbqy48twvBwqxi1NkxWbk0zpWlXO8hcSeBfZsuRDQgk/5Wzg3JYelJE2nqCpeHk8UdHP31
70CsA47yAlv5tupL9PVbP26csinR53iux+EqKSwBd8z5rYyev41hiRjkJrZPrS9YcE8ArvXYq46K
bMsPObEvRjtzKzzZe+ljpcN/IciTmXWRc0TlstFKw72m9F50gCe3mATAYjrygkrfdFMBWNHLj+k3
jDTq+ObmrA/ys30ADHT2PdRCKaSeOa48/jZz7cdq63QEkPmtYCdRyQPlZq1/TsREhgc5cGnqFCTO
6s1f/wJQYgkfGy/NS4VnFbIPYBYZier4EOYlqLk0JEgOJzWH2Lbo78ptmIbLjZktI220XeM82FYC
uexRUx0RO1m/qX6jIrTv/JnfxbJy0QdoodZOjc+0YloY5Qd3VPbnIw+L7M9eg4X43G3ovFNmc7Q2
4lC0jmR3tPto2jlKcpxYTdBSDGeiBSZBklwWOexhFpU9GSopVdQZfDqnZVL6UUkEEpB81eEfP0u6
X5xfL/72yJtiA5qcP7fDo9H7U3xQ9FP/EIDYVkFgN63B+t+TYqGcEZa8OtXMzmOHLMNy3cn2mEa3
2mnDezavPmK1Iu5Xy6Y+NuEDmsGLQ2SxdU/KvGVwZmrxY7seTHS+xptMMhc8qfKXa7yiqYkTX6xX
HBcvhNeTTePj1OCLvbzswWOSqnQShN57oaq1zvuD+weZb9lHhh8RmrH4cicFJbGK9ZVDWDydNISo
NGa6MlICiDdYJEQqWNqRZ2UQL/0Nc3L1ejM4bmp4IZTuHymRV4h2cSRr1TCJkP78+BKk9SGopeWP
NAdu1k7lbXwJgzo64Da/wNLf+NzPlAXPw79TB7gJoeLpUJ+9YOlT9mZ5/MoTcynLQnpa/R3ppRt8
2ez+Z2jXRlCtaXtp0WFto8cWyhmJLrBxxfsvCK938MChinT/jaPU6tnK0qGxb2YM0tabxipuop5e
ScpzGx9TVXs4VhwqiuN3IdyNq0kpIE8dBf281+f9e4aQcqiJtKjuc8JWsopcYqf6fsKE6X7AISZx
w+wHML7arYb+tMmW+t4rTynoO0aD+6t0rFalQCcRRr1Ldig+fpvmjF07zNoTgJRa/kpC2twep7ix
5lXi/bfXt862TE0SDboUnrtN9QU4a94hU86KYZqvXseFaDyQAp2votTdRgcU4IYgWzXnMRwy6fQk
VR4lgd2PgKw5SzPwkYriOyE/jgriq/nVeLcEznJfqRh/g+wtaReRpJ15asS/qe1FnqiWfVsaBl64
eTcy9jWVu00HHerX/bhO3N0sFFFDK23sZJg7/tnsJnOAqx3GxmQAdBNYScEmEvkzpSuJjwH4YMon
icZYBwn7r8l6KGsWBXoYiheLXcFDuePAUoxGXhxa9Z4xloenxlGZbxJZ+0gMNiGSnUhuw6cqPIzT
Zp1iz42c8URNU1dEUopssYjMqNAnUxWS9+V6Lefn9+mE3E1rU/8uKXl8Si5cUvRLVzU3deawSWYy
523+jQJq1u8tpjVNu5kPbZUPt7VFt9KWYJvw/+bxt9G0/7+o6N0eMfLEX/hN7lDzh5pBWqVvAx93
g4AjhUQaNzOlozwnqBZqFkqADTHZi2tg2IXGHWpvcjzC+LIbLG421LVagjTzF/iLul6Vg4pKSKJz
OHwwRUbo+K8sx9xRPGzpch0n1ipwMZHzr2t0yuyGseI3TlqXk9MryMQUaagxpxyTvFy6PbpB5hJO
JMxY6dbqNnoQDyqWZ8HO/gKOdH+8bt7yFogYf4PkzcTWOraJdebqfdzPitBIl/wCz5y4TZUNsd0C
HU7Ags2kU+O9aDFB7H6FKMbR5SxaOezvEtU4k4tZdhIddTnOnldcPZhC7cStXr6nGmJhKtSmp88s
zq7Mso3Lcamd85u2NcLY4KJu5hkVjb8hvGeK/Ta3VQfpRfDPKJrKiGsDbLvAN8JPqiWzL4lGplIj
2WiQf3eqB15LtMTeRQogfhxHxvM7Z/qDqPlhcrCm4+DYaXcIo1dqQRxGbMpYao/6HI43D+18aUui
BwX3+i2oae7JVepsfcJkssu8VjwKL6qi43ttWx2MHl2/o9pk3ur2jGlA0tAmpK7nMWQFkyflcHDF
8hvR4rVG/yT7P712uyc2C2f7CjhbHGRYffEZwc9H26hrJnXcPjoC7oTgdAwsYEzu0S/Ge6h0z0GE
zMhHMSW9B+6ihnIU2Vp0CFdvxQv5clwQwab/zEZJ1xFNf9iLAq5Gna6SjbkJL6149fgBhb7BEo6Z
73+0EMRG3rmGTB1Pma2tkh/PoWLgGGd0bDxL09QLfMNkH7Wap7vIYyVLHpbr/BHwkSxXHhYFFwuG
DDc5pjLDP7PfaAdksmkwCEzyf3ovp7g5l8j3TIqpK3O0ZnsOEBkJXkR/5dOV5pSnNEi9LZGEveQ0
6kKrgc+MaBuuSJuRV8YnYx6CHgdxeOdJ2xqkrmbcCFsEmqCyX2F4RRMGVv7LIiZoxINhwhB4GvWn
gWoUphEjK4Xgsf1TQuL7dNGYMqBKP2D3Iq21CGx/upAJ5oXgs0K/SnlmvjTZABvGhi9u6dnDnLet
jz1w8BClUtGbUF5lqfgoD4N+fJ1uXEr9OFq+23cEucDFkaVb4klTkj+bbFl/vlKfkvxtBsd8Ws4U
Rw3YJrLWkowM0VGHI4VnOnPvtzxBy9h14hHJUsppZhLqKoYLuYJs3uiIPQWa2xQ/P6oIrWi7CElR
3CmCGbZG7ppRUbuvxJn6iYtW+PaPI2Xif290g4p9JKzZKUtLHM2ONTLt/XK9y9zngFIi5EsaZ7Ps
LYxI8IC0asfdjAuLhC8Esj3hcSenikZBI6zVt6hqjvbEfW4Q6D3TMjxDFW3zX1jpZog2rWBwDo/t
QvVCOlU2s1i6ndOsEQYWJLGuQJQj1vcIbyrgxID9QG8vZwkn8J7ZNvjfCOmea7ge8/kZVv/E1+Qn
vFAOGhgOO7gq0B1TQBeyGs68Elu7R/9+ypEl+ckL6jMEnL4gghZILV6YuN78A+tNfEqijKMxpnGJ
WFKkND/5dTcF+CidSPGrvG+KCGO5Yht7PY1pf1DFJrVymvivbA35DiZNwwZjicQV0vUTijx18jzy
CcgsYITOLVrS4Vjc5oHs5x4vhkQ1nFXJx9jMG9lYtTfiinMMGYV7gzeFxQvn8sfFqC1E3YbuOpkg
E2/NALUkRMlDnT5vJ7DdO5O5szU47Cz0jALQUKMzV0BYspKXiSY4Rr+enKqb40sfH69x/T362kID
ObyXddl4hka63YtYzB5rtNj6ITCTTQ8+QL4eQK7UQfR4TFQ27Nf82C63c+AmKOqJbcdlWziDDS7P
qzdHpbeQblQXm788Jma4D4Xd4tN7Z8syCpmunBrELRp94vcfaCAoLV1z+MFMmv/J/ZDaBY2fg/Ak
2iYHP9BbH9vpNurRe7bBhlG+mLhS2HhyVIc79C+UEv4rMfqu1OLZuzvfIOWJ4lSQetwzbWpZxA6l
Q7p5BVJDXh2ha9MPVCRUvAYT7gqm+NLx2vi6YtQYmb10nSex6tL/VK802Ogx8G/DE7M8lmHLnNEN
GOQFtcugzt2V6lgn31GcKr5r2Ib6Khsocu4+TJRC1n+GgJ8kT9bZx9g1mOYYRkoCezGum8dZs3XG
g5YxbDn8fkQmbvXdHDCgkBv/z1YGnx3BIoyQ2WntW7zypE+oAQHWEE5f9dIqDocbjYB1RrmlXS4q
zYURLIwJUp9K3Aosc3JKBHiQSDcxGd1nlN0Eu9ZOSEmjEj/rIr4R2i21w5ax838sHpvk49ibC4/U
vHpK3ZudGE9oNrjNoyDEzvMpC4TlUaH/fdljIlE2KcoWYLAxG+S0Xo+bH7rlIGN01ag6GxO42StN
x2VF43Gw0bhOn9roZCU2fmTXjsK9lCygEdCyh5lX3QQfOx6VzTDO6Z7lR+ZYV3A4sMDUX5LBgVcZ
GMdC3MvytmsfAR5br8fGZT4aFIBOERhotMTpZTgHzZ+BDe5eka/TMUKIGvH6Sh0XIhGgSS7TPa1c
bdeiYqVmmpF7ojMZDQFKsoisNBsytQ4XEaq/C89lmjHyWBDUfpt/6QIdnmjU8zp/J/nnP1K5KB2R
7p0W0pv4/QgIrvq1Xx/PLLGY1N9AGgbvyYz8f/Ai57eF57Ku0K1dJHygvC4b1eBW9/qTeuv2Cnp9
b6OQU0UBABmm347RZqhcLxxFAZw15240r9eLoiAbewps9ecvxLLWiV5jiQ+DvMvUS6QiWIkAAp1n
5JBZBo87n1Psx3RFtpXNSQ62rPBb8pHRlu2G8Mj4VYslu63Lxfk0IsUIfYrudbiBXbtJE/vnaKJu
pZUseyNmCMb+EtorBba4dH0IkTJo6+/GsqbT+E+mv1uLyiXDZwkA0LVWn4CH9k9HoCUJQOccGMGl
2sYPH93c5RGDEPkhtjQV8JpG5u7aYTxpVehvqK2eol5klsivx1+5uurpZCru5PjfrP7+/4f4Kcog
DiyDKJ/4xYEFTKG+qPelNOCK9B5Nr4xHY+3V8RSjBMBzK6eP4T2usIEjrLRfe3jY9b92yWGsO8QO
qODlDV+NxGBJURsCHVvA8+O8Q7vVgn5UlBfl+Po4jeht1fV1Qu28JFJREs33ZGjRQKpX1sMBAEiQ
iiMS50B1auM0p74CxD2unrLjrWKPAwNVP7kENO3Y5giep2osB5Jo4LyDJBsfot5rkHtJ1whG8sLS
0yPfP8u9IvvNtOf8vkINfUF3/1FHGJ4r98891Hh3+tl808Xl03CbCkzUXQRQDW4PVqVqNh+tw/Cw
0q4e/qOJAuLvCjYrR+tEZ9D+0WfgSzNBRRHJ1/x07w25nWd7eQpsy+g92bnPL3S3neBialemRI+e
/7r/1UyVXNB6FkbNARp4Fv2V5hT3pWfEB43z9j2H2nYlu44by7Dxp8/CCn5gUMOd38bsAV+iX0Ws
YFi/CNDCv52SgXfv8lZp+LWlty88PBgXlTs3FC7t+A9eLpXY8BVvp1JrLsxPwOxuVaRTglzNVFb6
sbV4Jv1nR18q9D8RQyYWU/Y5un2HHeYJOtU/obKYXG4ybCzk7TNU4uGXVkVq+z7WmtMJ8TOljEl2
LFYr2XuSSleI7d33oK48g0oZ+mjnC6P43VvrDmhHtfF9FkMALN5wRT8KJlfhSgfiRpDdeSvwBmsh
IKI5Ea8a59nrs+L/8kOSo3y07B2g+ymOTrSZh1Mwh3iatyI8lIEcsGJ2z5zN8r7/qhlMfoi3OzyP
XAXxFiqj4d5+ymZZus+VlHUlt9rlhSI1JBkCnmF11z2W5YIja50npxYUMXEOVDYyb/w7qHJG+bE5
LrvN1u1HaDgJT5dXC2Nq2nAPZUpEsSulR+5D4Xp7/nho2n/RM+75eHmTjOKjVoy85vp913TAqEeo
tp9ehrGA8bbwMg6jPYKQq7mG05RBUfo2qW9i4ZMt66BFf6vEm1QEVAnVBHB/j7+q7pc9RriapOuw
eKZGqzhp2KzYxc2Kcy32wTlquTtDuWe94Wvkte2vSxbfZAodvGZP19RDWajQI3yX4ggtcmYa4Xd0
lhbB03zmKn5v7dnXWSM27YA7OLcfVr6qDeMdHYDgGATTryiKPjxzVwU+5Wu9zsMnlJWD4UVRNg4o
IvhQNLjFzBrPdta6LejsMNtzTxXHVi1YNWoMdcIZegmz0VWYVwLAym97Neu65g6L8KOEoXNSJ64f
hFS49T5q3dd07DfDZ5PX9nuQU61WuX+mmD0zMdd2z6vKWav5UaBJr60tJhTYv7br7cAtSHNFRk1h
WfmPUddVMpBBtlbDGEKuqCPzazfvjK9YWWazG6w39PV5dJpjX34+sSDFIWGEyKqoDuxgSv2cHsaK
uBXCSAAvs57vilLVHJ6/efM1dw2eMMD3AVAq/1DRYeq7F57ZOOmq5w0oqkdQbEAedCT57qy2FUDn
isl+26e4R6M1NXFAAdgLQ+PuvPhpUrE1A+jMWpnI1N/N0++g94gjCPUkiu5tTq3cQ5CF/E45svAo
4+qGfE8CMSUjcEFom3mlV9/ilWUb9gM0VgDQGN/5jwXuLeW3TYXD5N0S4OEZ+quj4SNrok0J+heZ
0Dr95nWjapcT2nrMy+ZHcSTNbP0H/H7CtQbSZquQE9T8N2IBPHe05iPpjWepMfIChHC4W9roYgZ3
I+bT02EYvqZadVD03RoRvthIzJkMCf7TKclkrFiZXnCoW10wxZ9msTP9Rw9waYWXDOTRanC8NDIb
5qdfMKmxG801taCLrhHab/fd7GlhZq7sL5TUXVQL+UAJS4XZmx6qSDvM7NeAep1FwExIfMDgfLjL
uZyJrVX9ikAIZFKCBKuciFr7WQkx8/bkRuVJvqiXMkglEk++44Evt54eCmTdxU4ZrjDvCTkVmTyW
zqfXtb2qQvnze9jpNFXf7U5kcrpZ8AxBIYENrVqVNaSxRKOVdLl9z+alHuiGApP+Ufo3b8Yny4ys
x8XAw16/6bwo3HzxP2DQ0oKd1Sqo/L0xnc6NSPKFISx7e6vMBkeZ9PC+XfBOTANy/z8RQUHDoy3y
XTzZ9BdrelW690/AqH+4EfSb3d73mT1Jh8WKuWwcYIvqdzUF2q6pLKSuQufMwtm1c8qtAd3XeONi
zfFcAe2M7A7RcymWtaR4RGwBeXFpliXr8XluohcHhvcMzzts9YQfkSedj4X79W3gA0RZaBNoIca/
adM6rzcexv5E76HOPV4ZPzygM8VNXsPJqLH5/k/CYqWUufdah/KJe+I7XEmQ/Tv+6Vk2n8BuQLVc
tZFMF+4/8KflZuTgsPKtMtziIC5YMyQDGcagWRbK42+ZpwwmDXurktruf2BJyYPdUU6Vimzpz426
UanLbe/zM+ZgqsStH61xn7f0rjvXhQeYa4WR7qNooPtrvrbyf1mWWp7JqesVz37SAWMSKxqsa2yk
J8ozeFQM17UmwQ7UfMqdnMk5VQLH+Dg553tJ2lzFVbzazcIlVQMZv0s5kEdodDjLSkwiOz1bsmW5
Ava5tFbYRHtjhL+1hPommkiClGffKfJ9+9YK8rUpED7dsOa9WvRx1wwtlXy1yWhsS02N72AgrFN+
2EI2s/oM3oWdx3BjVrDCeJ2ZN3gxM19I1lS/+A91PQB9C+AiL9AdAOqUGuvHPUHuWqq7VnBJgxb9
sp4KUzBAEfzjf7QuXZg7Uq7xYUZLyJn3jtDvrnIpdlyseZ0hUyScYl9FOfQhq2g/9saRMAzgWa8Z
/6+r5LsQCkUp8A1MTodWDg8OQ1kIhSuRsLxKdzhYFVginX+9HjxRwKqf8/0+uM5VRfUzXG+udS/O
fBDVAUadVid/En0NdU60B0Av2bJ0qvMPh6T5S1+Se+B+zxH3zDrJPcTx2p7ogbXF3z84QkCE8/PE
YoIR5trBiUpw6bK0C0QC33OYHlB9HdjR6FpvxNQ9trztuYpx3iokrDMV7rXqhcKByiNviB0zbBe0
8VZlgQq5wjw6sPclKHYY92ehadE4mc1xu4iI3TeRtQZpUMEzOG1hy/HD1UVms2CZD5z6cK5Bamm4
5CSmAdlrV3IcE4VGzAsHFY67czsueBUKxR6XZg0XO4RbAdJtTH/5NNERICE908bc8uKBllNRb6bx
D2gUfVst0y2sI0fnCPJjyE5fomC8X59bktHnV5pjHdDkQV5/sw00xM0k9ICLpmUOPHpmLXQTuut8
9WUO0yXzzYnKeZ857NaEho/ShRSJpOEGqMWluvRPDUcy4R40cYQdaBmSbuZ8hVE2n3gGn9EnKhjV
tt4/dQTAI3y9e4aGyRUt7lEXIkxWvOiHoXlkgxfWXT0wbv+YyUdMDh/z9AsZilY9ZPSakGrYrQAZ
IAjhwAdHMSWVYOYlFKtT3BPuN8/NKS1IfP6KtD2YSsruGm6IbFzPbm32lhc6ihboGw2KGdU4Jr+U
KSOz23/NDG4xlwA79iq5Zh78pHKiRh4cCfftVBX3V1x7NtbOQ5z4SpRosd65SBLONdHiukESP6Ju
ljYi77xvjfQFkKH7DPb3puI0w9ju4LffJ0MAAGXr7Y1G+MqIQYwT1x1EdGnOIwkjIdhjvzFmG1Mj
leq7qm4No8cHs+SlmOPf9DSY90+37Rfg3cOHwGLMi9JjDmwonTTaqlot50kgeAaa+LxwZD/ObrdL
8xuiMj6IHaHDhAYYGgkgKHKrS7DSnepAPVfmRmlqomHyzh1hqQBipqiaO2AO347qaNU8RO/Q11EM
aczc+2LJU0hzwyqSTkXxDpxESUz12FpFVTaTFGhuPPN63th4N07pCgQDFM8Jd78QK5bsj+ISo/fG
kKGm8KZ5M4wl7loqDb793YDAwsLR/rRBjnqQxp6ALXaUr4mRmIMTB0mmtGHCX5KcLOuYom0kwfI+
iAROAAN6+V5gnNAtqM72Izwx3VmFwhcGhm4Ij4J+owtEk/J8ClHTVZLe4VZSvesz8MoOEexv5Gvs
5KPUS66UXY2RXI2TCo52W9gpvZz2tQnuJ2Yekxc4N18fivv3SWMkR4G+/d3EFG0kv7a0WCijFeZm
8fXb8RK5H/e9Ss1qS9vYxlLq7dzFxI/MvlE3Jf9FLW9oBBD8PaznfCJ7zByinuZCW+xYSaljGLT6
kzanUa3/kvu05ksQVNLK+2Cr2EZy44waNZApjMPbCvdYU86xIaCrAUKFUI9V7Js5tDaDXHv4xjMM
DDhtJS+WDeB1dTpOUjh90FAr+I/Tgox2a8TAgQYDnxPglckx0o52p0u6kP4dLOScSedcKwhN6JFt
ZIHKyX27IGTLDfOgdsJ3yBQbHe3xqDMkT6fwUWFuZRMA4WROEoLITYfllhiF+X+hu7zXZqTMOYbb
koxusL4yQBVLNH/7zCIlOX9v8CYMend/RTCHQsuEUPE32vEuXaR5AeLV+VQINRbwaxzwf1uMzmrM
hhV4Ykyj36lvffka89i9iUNGNBGynPKdC0+0Wj/L3RX+j4bkjZJGAGLhMyCKY661KzAYLXZqU2ZP
Wwb7iV9deQwp6daefk7kLOgzI4c3CoE6nTv4VsJHmd9XiatWPq4+l83wefLOl4y1b9VblnPK/UfQ
Dgq60iMFMrw7rQuuHLDVrAV6TJK3DCLCLgsIFhQgxGUoqKTtOFW9zQnTd5EHx+mX1+OfUahiDzA4
wnVzvUJTdENgrzR+Bt66iO25Gq4QMskTubQoAaFo7g70BsFvDf+5RpVObS15/5VeLy+bJdJqXibq
HGb7Wy6Jvr8k7vWZw2ws71oIx8MuYA07Jmz0inn8LBs+an7SEP1HdWEtcmD67NZjD8Qv8YAVka7v
vJ6SPiJo0cu9Cw4tsqgHXRmID2nMY1beL5+LyJgY6BLDyHm9kIyuo1v5XIP7Q9MNyGLz26yRZUMK
MRjiHKVm4cvO0+7nXj/sfP4tgHZ9gLN+hd49GKg7byXQoz5G3gbx6Gtv7gDOutQOAEg1PqL7q8SS
MFB8CIr/W6rhFSvc9SdH2I53+jdfCOXVyKrk3AFngFe3d7bw1EkjWtceFnQRImQIVZCbyTE6LpWk
L0XPuhQn6YB1oU3/X0oA2VP1lJs/VSkQdMU0XwEJdOlP37wW1Ja+BT7R9gzh99qbwH/yavoARZsB
uG9f7WNuqSFeAxVzv8JcJebwh8myW89Iu69sm1J9d1tBRBdDvw5o6njhiEdGzafeEHJ8gpPkEogP
2SmheYgZ0CpXxX96KjB8GCokM6HPiDsnovqzweDPRALagk8MZ+8usBQon5CujMv0b9+veDMWb1HD
3EIxUjoBO0CE9GSMeqI6SzJaETA7RYC4MQZPEBAuoSEkWB9no12azGwl1wr38OGT2CVMIN+dLM/q
7HE9lk3pZztwQOVlAxpyBLNp83NuwTEpD355d2vyuofkwAmJ6/C1Z8skWKf1GpmrmUKjhIeF6Fma
8Lk5H4PD7dDLmBaaBfiv5Xr6I1ikAI0I+C3NjtzDGBvXgppaCxfVqnLe7KdkNXwjZzwDoFvJQeDs
owoFrrIvA5FiA3vBVv+2TM3MPOh0rRWKjp7zBerTjNLY2WzOKaGZxswiM6uH24dEJPRKdMEVnQuV
iriZbQqt8FsOb/PV83lHgGglrn1Jj+BuS8JZ7CRHdIY8rrrhY0QLOOzd+yqb3I5FAji/fKCBmEJ5
FtiMydpyAg+5oyPZQw7X5J5B2Wulz4WttRh1jLQNFesb0azjpU4GjOCBHm5Qk6uwr6bsgtJAesih
4zV8GCMpxUj0n/X7CBdaEbFWrRY/qVodL8fTg5edKGCpA+3ivYuLz2yNlkg8VaeL399UjiNyV2lD
6OS8cl0vOus6jyuIgwetjLmcIeevrxOslJrqWR7x1+OUA72U2j6Kwful3jBeNq4Q5KzNZ2jsJg6X
QM2SL2wktxyMGXls+yURrHTBZtxUbmCwWVycFokZ4pIYnzU6QuOIUaafLtMj0/PBrGY8qI++EowP
3v92uKCv4kv5DkdWiq7VdWbuvw8u9aWf6GAuXG+IoIHhRnipo/M6aX6OP0JUGefN9aEbLZFwvBO1
HrAe3d6R7G71UwfDq4n1pbZ5tq6PATkQMrZHvRX0YWDs/xX87uoeR/a4J7IBD4qiGN37oy1OjPhq
KkMt2IQJb8KZ0RwG5b4prBHrbxiZOp25j7iEFQ9Yy1NCuvJS2o5m5jombU47ODSzFYd7+J9HhC2B
gj5uedsDmTUKgYCoHLkYifkPQUh7s3AL/QpKyaoRqyCxgK1zF67jTNWymZGiGi+VOjuGmHLLTjQa
yYsX/jgfyQHl+Ns3UFZ3UoNO0MfwGbLluqUrgl71vU2Zxj0Qj7sCOYzCz/XKqEF067MA7OFutTnY
W+SOk53eooqmWAnlEO2QNEV9rnGYcbLOb/ZWqYMKG9nmaaJgt7K7AO6J3idIyMkQmQmVg1Cdzt/9
fal4meyUFtB2q62NLXa1AIGu+TWoI12VHx7tNlIlpwnvUfBGn+5DsEnmVZZ9RXzaPubD5pyqdz/I
nwlCA4HR5g3X2H4JRj4lX3q4L+PqddT1LFCFsR3527CZbxkTuauoYqnkfWJnfqpvpRl0tcl2YMOE
TMqFCaQTOwlCjq0S6mjKh0btODOcoZWPJzrBckJAM8TDXQ2nNcwdipDzTSNvz+T8BIpS6DLeKyFN
3L7XOmSgUzGjcJSChxRyRvDlBxFY3l65GzOYECZ3FOeM3mkxQL7pYpb0L/dQjIQnOziM7Xp7dIx7
ZLnWCHHwcDhCpgJSsVd9RzMaFI9yrrXsmxgrokTY7Ism9NL37NOnMBL/mrZYZEfH7EmTc4mplVWN
U/rz4ZsqF+cJfbqflhZ4ltGubauNwPAxuhl+HOWq3P/wLLtuD7iwixFoCFuSKSO43Pss6A8oamtK
jEnSV5JY/yRORZ5UJmJeqxTfBW66Nv22arhq31+89/r9wmBWR299W/OJwcaHCVgehyWSHI8Ye0aA
WrISJL/+dKRlHlVer8/MIYgVzJwLLO7sMQe+nUjjh3wOnTTmHW1dWHx64V00VWuVjJM718mcsdtb
KFJathWMrI1koRLoJk4zvHBdQo+pPniR68t6zMG8AV7Y0dv7O99FOf6Cefb222YwZnb+JHoK3i73
8UhDIgRXGcGn1sUhK+r61+2d3G3NM1Mmp3gZmoNltOt0BCykhBMYx/2lrTSQlRUTtZ3q7jhoRuxh
BSLCSke+/rp+em4DxYSfQNIkt/7v9KxNMOtYZtX1TEUj9mX1ok9Xu46peEXPqbRYyywduVGJuMsh
cUy1R35/a2OkA+k5JVB8gCr+8Vo1KgaqYHicrq/UwL7L4MSD3l6ntIb32kzGwxzOowSSzPFpaAEj
BMKY1ekiaYN9t2OFwD0VrryMKHPmx76goqNHeNK0JRG9JOjllHXWToSk2adQ+isyVOdb43djp1vF
ZcElI8WmlXZ48nkS7zUHg8loGzXpaUtaJ3jzQUFuLrgtLBIBgLoMgH4Q/cAq2CfAu768CDVpC60U
kAsPqso7e3yzbNOf+PEMPJjBOWSypx1+X+dcDj3MQB/sIq72UzhqFdmYGfqxM09wmV0hbohcF5nt
4H+8QlFRE9gji+CXa890xxTfpoWhcOHcSetvXQwHB3twSr7VIz/mNxMbAdzBQcsZAwhzWdK1/xl4
qrWOjFvCSQ2SoDBet1+TZfIdTk5jiz+gagLM4Kdnqkm5j4TFW9i9g80EJX96gKPhPbUbv3Vfz/Kf
XqpT/U+OUcFywwmmjfeObilAqI3q79pp92SY7ScmUYoDsSh9rkpTVCrcidj/yR3a5dpjvGftn2t6
pbKpb3SR2mdGkPze1b2EE+UfZXHupoTJj/uylCoj/nJ5yZ4+tyHKo5EkJdD5ZIRoeMxVu2BI3Yz6
8ym9FKC/cHUifqE2ISsCMI550xXVs1NAX9ZHCCeO+ppkLoneybk0PFkALVp8CvCzrjC1oR6o0KM8
UuRNrUB5wNKCgsqYj34RULV+RBqPhO6MV03ehulH13jb5BOAlvKmzRuBccz9VNHuabZAJPHlZDOI
HuUO1zN3C+jNgNz2arip3Hbsb4XWbqGw7Sg5IkxGHJJTWJZhskXp3S1YD4lg1OYHrgoQevhkratL
aVwFuElGNs7i8lNALmZrzLQ0WP+p1GLdlPDR2/9v6BwBGTFE1dNREQepf9fqfPPVhAaYxWg33Ni9
44Mp5+XSzM6g167fGWpAMkpgeB2LmrWo+KWFWzLfz2TFmsv6ypJeWPrqOWQz7qEhGt/1qcl9zLv2
OXsJ+L5GFgkRnPHwEFcRUtigzsJr91i9sK3Qj+ridh1KjsOpntDVN9Ic0YJhg9ZB8+iqlxOm1juZ
NoLW1+P1r2Tu38Eni00J+iA1H2FwF/sSh00IEzTgcu0KqBgQb62fpqJpsAaTnH64ubRaLw/7ugZ5
lI1GsRr8DNyFIML0bb9P2VSSt1KQx8q8PlffTOYOOeLv8MvyrzbsW3fK9EuiQ4eNEtPbnwaBcYfu
QVfLy9CdOEKZ6Ga6oiLdDC0+h10njBkfF4967Bv/C4u8eLN/AWDO3guCUcPfDoKFjkwQtgxxnV1D
2Yyu9t8RdGoGfwYX4/Ikve87XtFqOLPKrSTLRYA4ku7kbTU1VfllT7RMSqCzOVM4yLZfvoJzlCnO
3jrUzLONGB2ZZsPRqcWzZAzJMd+Vm0bXlspbfs0+VCk8ggqKUXDhNto3ZDE2hFrDW8Jp0gTyVowo
o6y5bPnmLCUH4I1GCvbG2CE63FAbP7OTi3ZxkvJn0s1GLxikr5m30PkSnphKMePisf33kb1v6IdV
ZiFxb9PgxxsXZrgDy6O4RJP2d+XZ4/RO3G2k/HsfMb1KBI5EZAXUFO+/Syf2hOfLJtH6pETmwCI5
uNlfLlXM7ltASWiBqfI94rEbrAzFbUb8ZzZzgfHm8h5TimgL/CG/4gXOAgPhKA9Plu4pgms5xIzI
DnzmwtaXX2jcM6FwqI4My/TeOyWPiFhpcLPSYLEO4i4PZSsc4/CWsv3m2tqCw8D+w7o2j5W7yGsJ
EKgdfKMX3rYV1fArz5HYm+UBnvCXVsutE/f+ZgZ+u8AWm4oPiIqwWpwGiC7a5tWyDcsSr/yCtN+6
LaXvoEP7wmd5WL9KweTF56EUKjZsfsNBggY7kDW83ID4FjCvq5t7mPV4v0unyMykSw22WZ1AG3Fc
yvexvBpUEQHZkd/97/FBsM4+yv7YjR7sqGEieEn0Ov/0tQVr+vRpwvNAGfrLB4Y+iVhtptYgNC65
wpYxNy0mlL7Xt1S3w1DWoAJvcXw/rxdiUQBLPirVg8CBMpePVXI5vTq/zL5NSqa9K1jqOXbITTM8
vvL5yqo54qlCF1qjiK61s6gbaGSPtoKQm+2fcX9TTHokQM70QMJWcz/6SHE+2+Dm1VfCld9h7TQK
2Q9tfce2ZR3RTzryjhgab7g90rc8AoRf1O7RquGMxVpjYq6nhC5Uotr3F1V1ym6Ci2vBh9MXnedg
hP+tzu7D7rTqGN6BbB9HPr1SYAnFamWXNi0Km78n9f07K+WTokRFvlhAY7x1/eZtq3ZP+eksz+nN
qYYWLexY2eKVlqtQ4BuSC/xRZegAM129jXK8xc+o9sBz37XoJPaYsgaPCSHnCjGEos6NNnS1cwfv
x738mDKpI6cgzMEpOmy1vQKl9qXDnnbg93MHkohglG2zusPtFINR/YSF5lVzxs7SrOg2KNTO4XHC
QJcBQi+8mMjYLA7PylmbzTvH+/iys/ySXPcEqLqZTgsT1sVDqRdotFxBodvVdh6Hx8pa149ABWzb
QPdFNhvr8eraOvg+8kcN7Nbl0mfj90jUganIW+1co8N56IogI3c6UP8fOAX068Y7L+NbvNnVBCVC
UtpFDGsMfSh+/gAo3B9T1mS6QqmeQfXp3JeCqMPC4DwHllbRQ3MMdvO2coGz3ucrUrRTZ/M+pA1y
ffkIc5cN7lQguhvcE7oetTjGm2oNod1SQtCQXMZjugA2tdDLSnvitup0K90ZsUsB+am4N5Ejj/DR
OhV9FLVasvrbIK6hh9J82Ov8yTUdA4O7KrQ0+Q16mqxRg4HbktLLSXn4liWtGOgbwwaO3GcfjYne
dqPTtY++nL5frLoQEIcXozrFXdHeQPPXywbD18md1gJrcKUAuF30WJ8rbgrYjQIh9QjpWbZbAUc1
dMfbGvUxOKhqAQtnKX05dIYhs9uBGxesTuPkzv/6O0OEgp+Qk6V24f7ZX3+wmiBzPuIKvlg4AYar
E6yyfrzaNscBLuTRw3/4NBNSF6bl6fEMj7UQrvjRTlnQrbNbz3rrm04eyfrLAMP4JACyhrQiM1vX
VEUk+tVq6LM4Kia6WNDSHJtM9wbn5FgHfSwG8XxQFahEz7wcR114BRo0a69wURo95369/9hHSEMX
wEznCxuMmY1/Z21uuuzocXGA1le0YNZz1gKd9yJjGRo2iIDCkyQPlQ7eHOmdiITnPJbG1wZ4PsdN
w1QvdedQ0EWQLJdulHRXDZrMWDjJoi6rlOkjKzqXNNYCQJ82Yd8RfKSS5XZGUDgki3qgdRNmYxs8
63RPycUOuNOPeku75SEz2LINfs6zzhtCfPLuvi3UEfsr0xKbmR/4MQvHihTLOclhf5apvNsY0gUb
Ft6XFTMKXRnL4V0rXBOSty30RVjE3zxVFQDPNjftpVbtzBVBedGoE/ziuzvTePqXRE/l+wUxkwzv
fGNJ4ov4IvEHegVxDl4/K0HPWSm9lP8LFrvqu0ge8vhM/gMhJhKUvjeKHkOHdiSXM1ANtxh31H0I
WZW5IM0nwe0S+en2uF8Vnf2xJAn/3kgjt1PDCj/j925CCB/FEPla7KFYCsSv4tsMcXU81xfkBcgY
wTgSpR2+6xtX4h1SaGchZGkwxjoYwUsSafyd1EdgMLiHYEEN94rnA3oD6TvRrvLSKrYhXRTSijW4
4P8mOLoKl2rpiER5fZhxO8ujevkfje6qd9BA1gLMlsCOhynL/88EtrS2u6PyeZNnXVuimmHhj6Db
vK7fL8BBDlP9zG/VUP6FxUbHVMNRCocWdig1wVmghUEZkTVAMyvkyseb7UVzjN78eGOwV0W5lgAa
TwS8zV17wFeyDyC6eCLgrnI9LnFt1+LCBDWLp/KDkJa44LOTAw2xl8fSIQE+LJKLq1Mocr2iDfef
KVD8m3lAvgnhi1vybcW21OUm6e2Xj+AcLLdWKOV4apwT9FF/PZmHZJBQMFhwCMIe+osrjuj6+3p1
cqmJXpW3SAzb3Yg+q6ZYRkRU/2gXZaoYXoJif1aJTwu3bJt91R5c3+LKqBUUm0YAJ35RiJsziDlv
ZwgEHMDGA3fImztYZy7G8xvcugFSOA+hZCG8Ipuig/ncBu5ARkuMPpFEbnSjjdwRdO8oBeMShIsq
sNH2xuxl1SulUFgsNNYQKqtKygr1rgHhTJXPpGf0tW6rY6NzsBW5PUnWXfZc3nUw3sqDzORX+h7g
weaxwwkSKqky7M9OskGBnzTOfgpTVWNmrNVN6I8l0gYZMlfEahkY45nq2/wY1c6UHfmjunYjOdIx
W0RTLxuRV+aAHJRfG4ScvBxhFeaNP0VTDQxuG+c9qyoHix9cvC4K5SIQZDtIBqK3MXpyEWlbFJck
gywcy0DsSGCYNj3fYLBq9GEq44QIDlt+8Uxd5Ru12J+9SCN0v0K1QmAsWFox8A7IjNK7da+RBwp0
EdJUfS+12EXTAefDHXoH0GZ5Kahmf7We/98FJf773qTa9RZkEgpcFA0SuUxARLdTTp1SPnrTBWzp
L7QeRYSmWsrjJfz68WFA7M3dkMgG5et1oafDAwGd//v/M7wpccCrrExCdQ5zl3TsD6BS5Qh+BX7u
Mltoxh64JGkD9R22kSJ3y8CXPZyevdUefpOyXkTaRBAfFNqAaSzlrlUgkYeYfYPVh9BE20EUHGVS
rOH/nD734TYAzeKvKi/9YkPepJma3m76N9chsmpSqS8qmwNv80AVODQ5dAyYwThv+Q7SCMIOW3R3
+QuE9fU3e8StLJ7Zi0mP+UrcODCcc0YANTirmmXeV1z1h02VywbnRv9Mz9z7+hUGFk2/Ug763aD9
WX6Hohv+xk5Y9ZGVqu4QHZZ/Jv1fw3utfvP4c1AzXMW6hM7o/G29ZamtYOjVHla/vgoOUayGiV9I
4Vd6qTWLpVxPJe/L8DInctpX2+MD+LSUyu1WpJfkbdbFZSXT5bOCX3E+3j49YSvRVPG2ti/P0Ltl
ObhqKQ/n5SvLQcnlYoocF/v2txt+fX2UDo2qdvY9c7YQytNYQGzPyIUQVTKrQSM0FdHIlKQ6rSuG
dZgP1gCJcncWrQPlEImVYRmUw7+Zvk6MNJ3ArdY+zDJUqMNFl+3dJLdHIvt9CkWo5SDtMQ9wujBa
CttJKbRO3IbUndTakNIqiH3Ks6rCrdZT6w9oIxemRUFyz0+ZthFnDi3cbwAqhZsrby+nuXSNNMO2
TRzIDuYkMub3bc/vmdXs8T6zNVqH/PcDwaq/nvOmvzmlu3dLNVVKqtjTzHzbArEpnCBprDtQmM/i
5cD8hauDVgFR1Ho7l4WMaK8/+lwLohFYnJv7/iqNr9GM0BFvFKMeeh7SJLQvi/519jFVtNCSajJD
fHgHnnGzFles9ibcOIU3+Z8CvF+pMQnbqbYpDoh2rbCHVB7/xmZyxAZ9rOFrP1gNYeSsTlExffU7
VO6rTSq7hAJ3j9xCpSjWXc+wEs9GuPLRALPL9bET3MHubwUnK0XQTCRDtan/SFxuaZLhUJM/YL+/
A6GszgoW0lIco3RR/CFG92JOO0tQ36Sj3PaMIoE+i0/zjhDk5IaAvOWDee0ktD4bIjpxyr2LbWNt
sCLWRkCCVPILiKEUEt1npufuVpAaHhfhbgnjp6vTAlsrNoH5TVKPz8Xbr6/5IYZ9ddq5YFvM39Rw
vydG9LDALLkHYMG+ckNuU8LjmGKP3dm/XNDQzzI+RfA1XELMainhSE53cSaFFe0KU0cSGk7RKLtx
pCdgWPAmG9/o6VbFhijm4RwJLSIp1gJGHyS78mXNtDcx6qPXy0N3mU+Fncn0rM1k88ahufcPLsvW
GyvAEJy118rqZZoaY0iEvvtrD8GYUH6DByqVAK+TLxVdxR9z0MZhk3mwGVcnwYFYAKKsFjZU1h1Z
uWp2DLANQEEQdevLVYh29mLl1Oqtc7Z03BJ5Vhb/fDgocjHyBZpMTeZtZQElNFTxn0cHIOybaEfQ
rmLfofB21v20DL/nnR/4oyJ7qULnOAEMb7dY8Sf6Flv77TVwtyf0iWm9RpEoArcjbfXbc0EcNdJE
jDhDVhgNEAxaKg98GZYHfDccpTkSbSRF0Cg8D6Z7y52il19FzSl0XyrDrUBz7T7hBXI7Qw9HpChn
P1V20f669FTVQQTYyDWT2GimLuVrf2mItznxJdNyrlgTcLufNu+UN7I5o9Q4cL52yDNDL+SvrIIr
10WxELmZ0LSZDphqog5x6yPRd+IoFAUeO0phqoTEHpfE3E1vxNA02zCnS30Zqqoys+WJZJsKkhnw
Wni/ZzmAMx4tT5A0S3fzPtdric/cGw3IbNbeVjbcF+CsmSoJhLnNOtmdnyvsCl2QIosqOgEgD/F7
YpVgX7H7JhEkE2WOwk1sG6NIV/3une8PIql8BXpBZPSvqH2RrHUKN9pfAmjFRfAtmpvMCMK4a0eJ
+ggje07/baM9Whb/eYUVkc5VF6kBx2EHrRD52zTR2CX7HOc1Nm6uu3NrYx0T2gzJBrHOB6c3Mkts
Hh4aBusNlapsyaSqu1j/oSPkWdyT/qMnsmuljsLc+kOWQUr3G1SjLajnZ9VGf2ziHf6Ut6BN/kRm
OBS3hcz4XJ51Avy4JnCJ71YvsKT+/8Zd6M1Ss8en2BPiD23DBdaR9OcgSKqhFvOYoSHjzeFiESm+
Pt8iI0BcWAdEhBtLMHv4CBIcQIujCGhcBLA9FX9FmY4IDSoZFBF9zA+9Mol8ldaOlulswOZkhSUx
Yo7BA8dYdbdTBuoZ4WIvNP6jHHopajdmi+tKS1IRZNo3iABH0grq6Axje7TDmF+F5MT/ChQAa6ax
+siwvq99+GBynerMpZluae+z1X1Rci7HqwhP16r7dpYMswB2ekXYF2S16kqQbZhvhtNjc4lfKzWK
P+/GcmjahVqETLuesy+0dmgiZAjHGOYXdbVCbQukJSAMm7JxRcZ7GPNCnpFa4ADrBg8pU4dz4w++
0OvHFUf6emjNs3AY9EB3kQPdrchv4SKCkBQfUwTK/XTATw9QqTS229xFmm2XpJAh4ssxyCFrkpUz
wuPOM8xiyhexMrHNFBfH3m31dPOfpIspbMTEYUp0TnhmFLm2GVjMvL1M3UB68Yojh7t0AdQH1iwe
jSQM2lDfg6MgUM7jPMz3wHn7lK+NgoiIgOoB0AuhWGf6gR+X9Zr6K/h/OBwhsc3sr9M16LPJivwy
X+fPH2FiCOw3dLJIoKXe3JRFg5nVLP3AEusu2C2A2aDK1NKAxkD3VX60m8HUH5DhfhN+7W51cHJC
19qtY8brDVqro5vrKNZypEE8ZGi6AOiKl+3fNmlkK4uiadvpQvRARQADRBVZiHK5Tb9jNjcVE5q7
P5EyYF1Llax21hAqrNybd9drns07YGlw4bCnz7Fnym0f6I026/L4vlZJqA5kp+0SdJeYkxXeGf4p
N7sD7kEkP806mpnUM5NV7XtSDBlG0vG6NCQnkefb2bIJTgbL/Nem7FgZmSnPgLGPI1rmVtE9eNBC
eU9iMqTPzF4nSFUdx0Ff0DfoeRJ69ioagH4eC2RiZYCuCQqePoF0Cx0q9WX902RGURppHGqj65m0
UdThUIXBUboU/2hvkC2WPNPzxaTeW6gbHAbWlJBRFriaqjJtEL2JKJaslj5N0UVVfTsWe+2Y0qcc
5EozxGBNI8JXOeBiAjQGThCHw2CegdbEHD8pteRJFXv8EWmn96RBGPib3gwj7bzrzCUft48WQ5xE
vo97NyLPT47hFd3oLDt9TgAoWLYYevhlV2b0p33GN01xfTLsFeIvFO0UodiEElRZ7UmBbOp3uE7A
CLG5WCOeNpKDiXHibWjRlWw3MJkMF0XpNIdyte0THNH1+QrXUtXT6SLaNE6HXBvT4H5TqZt/D4Kw
G6NzLO1Dl6g6zyT2TrAVjzaF/ZqVjsPvt/fwNaACbHyw71Vrr1MH8PXyyvRUREKq1KKWt92/NuXJ
v/bdT/MIeecXat63kX30/9pv3wd44kNl8Q5AnUtbQYNlhViSzpoi3ZtoesopiNAriiSnPvzfTm60
LzKxD+36lNcf4pwlu+2W/u9lpMo54yUlJc4YuFB9kJi3CKhmYznzukfVTf0Tw3l0mu8ollc+Ej4a
zFI4tDJN54Huc8oBMESlQQpplP61Fn5wLlJiv5Kih/VWMJ7IOF2lMYOXQW2oq3lwst7VPacfVqTM
Y+YsBkGSL5yu0EZ5HzwrT8kX4x6YbIfJJFlDoWjsvsOJQw1dz9aDJeI/5lQfi8fPabu/qeumfY10
ia4K7YOs280NaI/zLsBdlRNdxdGcg8CDNN75EToHIoVd1yTD6OYpm86P4DVLBFbbtxVNI0StSgEu
uaPV8aoLOana5HQ6t2nvNJtnItwFQf42XjVqRIVeZOpvQeZ9G2hLj688M90X2oPPiWXyWYrcReuu
WZkO2MKqdzuLzfXd4KjnK+utlTEEkdj33v0TLadSZvy54yjlmcUwi4JbWIuX5ZkRxC64I8UKYeOI
gnaTNhcCXBB/2R8OLMrGo50cFlzUB32g5hMLhETkrHmvNN0t6ZhviRyGmJqlE1NQjg9UnVIENy0e
3xAicd8/WdMcnQ/AmLZlol4tHEHfNdPEXOHtCnKORJtatSKlgwW2phuUs1ydTyo4Zd2kxamBrNHz
FwoN60o5IgG2R8T5qfSqNGNC97CMym6IJU0nhSShG3Gye9l772m0m5gSTpSq3n+OChal2TQIvg1p
bb+FARGOnheJDhbepMoJbwT7r4IViHTozXCzl1AzuGG19MlRKh/w2MCqHT1C2vO3Iu09KEdDWaZd
3YYT6CZQ2yPP8DNqxcuEeFUMFbVAvCnitLOxbMupvfraa//U15ptvLtmsztT8LNLfEskgEmVe6FX
mugZ5qi+fn5m+sWN4Ycdg8QB6xvUNKP3DJql13/+tK7bHq137taMUCr/yjUjnLH/ogUeqiPhIMuO
WispY3HErz4BJnkAlc214enA3KwwGhlsfcWHJNNAl16dHL2mAIXeqAtbuX/uNQWYtQblOpa40kde
vpoW9P5IF2zVZPTIoFnAISII7a3Ha61vzahimcVd34mUagEPDrIHcwoVt37pAbIX1KUTO2+RufwV
I3RrmcizB1l4LuK/8+KVdsS4YyWEpcpLBo4KqiJiMZFbg0JSrhm/6zJsPzwSM1cMJMEHsssgQOhf
6ogzI4YcgJon02yYfNFLX54W7NB7ZFT0wRlWMyIe1BUIIeAf/FXIjXfxVAKO+6/Qfp6FapBhI3Dj
NJuLesNPwYRPlI/U21S5qOzYa/n7/MaSXCK2ZVDvomJyr4QTomRPN3keyAV74evnk1MhU8jmkJvf
PM6Kzr2k24dyHceGDjNfr9vIOkehQSsWYcyGXBML2G3O8eDIbaJnwzDCHJAvKaWp8wx4ZUCHEQjj
dXTPjosrCe/oSJBscDl2ZLzH+kM1hvfqAyUe5VJHaXaeFEd7gz6kduT59o6P75UU8za2EBcOlzje
yLyMmiHuY9JKjKiSa0rEy7NrNVKCHSpPsP9DQZ6veiM0f3sblXIwStUcJAAMUT2ag1XrxtowapaR
vywswhQqSvQPsQGVzXRPO1Gr+t35py9Gtni39Hz6EfoEtCGmynTcc4rYaR+xG9wUDnHcYoYYKTho
feNQYprcZ8v/edVNZSy/V8rtmkoDhtP5CeoX6LbfDq+vDhzATz9GrIy21sKU/tQF7jNiCd3w0gC1
JTeyM88yj8jOICPEzrUQMmwxMt/LnQDIWmCYonJ+rOWPEDVF26Nxqp515oR2mpTVgZlMDa/eJy84
vcronG5FjO1EUOCtTT42vbk4qrRCCktKMwg5HtotFDeFOo1fV+uN2PqU6Dv2/9QF7CGgxKdaXjlF
tdQzaj3VbSeAdRhQReZVFH8jsdtVFEo9Qgy6AC6yzP6ySQeBqx/+ZrRJhFS2Pms6GZ3ohlf0RKya
WDen7WUzQztJzleNPB4kSI4jl5KbLed3hVSW1BJn4wZxDoW6vngMJQ3XX1hjERT8GMoWwNIwJ5Ue
2pZyn6PTEqxFc1MweWRFOaD3i97IHtu2Pthbu1KWx2raXxlSFv1rHwukeo2+H+TqgeIhdPqz88Ri
7pHHegc46PKkeDin1JZCuDr4/wUpOqChsonD2BD3nCuK2/QHDdo2Q50laliRywGed+hBBwjyBnaW
BbV2Jpsoti5h2yizcAXeANro/dY98ZENA0hZ67ZeehoYxiq+wVdkbMYSSiTRkXu/RP4b81cO6KAo
OWrkjW0gte7sU3eG3ZQD0cF3htfn3j/9WiBkWRZsNXUXdzscwBrssitWF2TzMJXiUxmv4EtxOgqY
crCNe9PLmmONY1G2lf+1id4z8hjDjT/kujz9qdoQTHGs4IvHKNmZXdjp5Mqz5E4SlZFVLoh/a8Of
zmBkD83fnNWayPwkDq4BjSfBwa+9aSV3cG4Xkpbpcf+/dcRyOz5UWFoPKN2RXT69YOlrEYY8HbOv
UNqPZXiLszv3YZyQNgAOoKlyF3MhEJB6kjHNYdL4tBwE3mpdbThhK+noLb2qn2OzMTjZm/agiv9x
ddwcS41+rRuslBR9ToUdQpFxitOS7az/+LR0Z1CTAX62EVHWw2O+dbGxKfCQnU4q3bwbWzzcq7A1
Z9XCAz+R4bAoyVykz0IHqSwrjxa9hSdQ2OPBpWIexcsG39ygGN3jABmUnI8+iWr4gyH3uFceUW3C
4v9pixzgmtjoTGH1y1s6xbSWvoKoHr6uNp+QqhK2RSPS/fx4l88uZ3KTh8LyfT4M1/lsBA/JP2/U
M8nFOZB0wWouyOaqJNjOxhPoZzk42bGZeNrrG9iIuHYwBcGe4bldHBwH3FflIZNwIPtSceh0q9w5
XXsAhDwEsr7TS4XYuNQKmMoSvEYCdfpyrUKjmyFx2VNj1rqbOSc29VVu47tTF+KW0J8VEAw+/BLG
8+CtqP+qYplICeXBSPwou8zZvPy3FQHep+goKf2wAFVohgH2ZtpGoy9BBLWr68RRAneAqW27uKu6
l2oFX9I1tVjAyGqQtgYpyRN5cXuDDlnYK80kuHE6Pt2xHmMxLdb/In109Zg85RZupSzD36g7SMxO
AvpZMfuzO0890+pS7vkC33WFgcQ86wvCJHnbmsIgX/pu4n1Xqx1DYw8mNkEK03cGrrpRb0TYMj6I
gI2F5pR21d/l6ISCQWNXoMWZc3F8pK5RldiYiG4Im12KmWtkJk9VEtoc4PekFZrxLjZ24RH9W5t5
8q4Vmb7XTRYNa1ZRZ51cDLHeG3N0+woIB3bfR7Yd7EpHtCbsxjXrbG6PfVEGZpyzn1lkF/Aeij6o
vvrsRmTBd+jTGhu0E2WdakV8ra9KYWJnZuX8O5Xt5ljJzqKnGBmR4A3LVjEisoeQY1KOO9w9zriz
xzSWU5Fa/BwTbGExc/XpQ/cVxYnMewgHmNyXdFWxfj4grWIC2nJkx0cqNkntgySPFUMSbqFl8ruu
b4VuhMaTdjsevBHYDvRqKfU/mKD5CarGID+uPloNgqtrYGLF71ImaqfQEabjPcSqT+xtWPkRO9xB
xWuSiOjhKUITnGmhQaXd4g3TKZuaxaboqMeqvpulPrOzQ7hDdL0ICGbRFaEvDf1HZRjyGPBS/b/Q
BfPvQEcheeNAcAXB3YZMDBQDACrXwsOtYwbLX8y5XGvNk5pVCCVk8FQJgqezCyY+KyNJ+7eb5EGn
h6yMkRpHWPw6g+C92YJG444KpwOLIW0NV2QWbgZou9DwKo3MSiXUOUhCWWbJj675vgU/gwP4BOLx
7h8t0Bp0+3xaO7DqDYUZ4B7HjylJ4KYhDZoLCJx5XG+2fD0P8fGqiPq9hyfoMkNZ8q15ZSq2JBga
S3JPzXif6fbipgwY31VbDiBTZUDPiaGKGwlE1Xqny8FYZW1oQPSkOFf2eKpEnngMYHwRTf9RAHi3
NH+qLG3OQlsi1xobTil3Sj0fxSBa6n6IOnGyOtpWuhD+g/qdX7DVfTH8MRBJ4PEjB41rO9osglyZ
SmtjaCwi+T147Rgia/ZnXJ5qWvG+nGR0cm7EtxuP3THFc7U93EXimwccoQGTE4BFfI5IpRQUQwF8
nyOr2ssGxgX3i2s1m/wzZB8Yu5GE+inbREK9YL5ZJKhLzwexMwbe68s/zbj8rS20Sg77/z7ZmJwT
EvTUcsInr8cOZKLh3qUbvAW0z8o+08bUWwlNd2D1BUyF1yrquVfV62b5Qo4REbz6nBi+GmystOcd
yvmepCSrRAS35neJa11xqm1cdi3mCDDmxk9x/uQ8lsrk7LjcYPcls6lahXvICXBQoifWEvzdYlVx
CxKpNFxigLmOozHaSnVdGIxt8jEPJpK8MktnOk2ze/U31Q9RwE0W0eKMR/ZIbhKvmceNPKCiQh+R
61tEcPRhnm8vtthi8D1wBQ1ILxrMGfLwoo1hp4KKJZxqZljXbvHh+G3NlPiRjyvUfVVAiXUi1jew
ENgR1w6IGil8IQAmNlOBJxrlMhLJo7s5bU96uhi9/i3DW5PTAgSg/LG4GOKxx39IsigQ5d+ec9Mi
ZTJ9Fmx+Eo6PgRSNDPM47JvFoCPlrup65k8dw6N1dT/t7ECjfQ2DpHmmnlP5XQ62Y4LjaxKdm+Rp
A8jJqA/xEkvxgWTfbXj5Avvs2g9E01liMnqa5Xfu4KrX9UTr18A29oYFROF9me9zkA07/ylLxaCm
kCUqdPR6959tvtsVe8Z/qtHgARXL9ZD8F3Br9TpfI7TBHAyB+Cp0TG7doL+EHMzN8Bg223xukgym
EZTR5M5Nhw1nMTSzQpZ7J5m5DtQyq7Fn7XGnVeednGQp4e6CG7xqRzlzaz9R+MZ1ofUf6gu9zRHc
evOGPs12/E7qidyKa///r7t9HK4tkhV+ffvHzXYHRNoqiPDAMN85Kc/BQnhbAyRjrcEvzvNkjDwG
cPdeeZN5qOFb4/zD4RCHSO1dGLzKu31N5E5QytKOHIFdTTHVdZARrbZQaJI9xWo0nrpeKDBqzLj2
++MxbhHlduR9ovLVxCLol7U1p8r4mwdlHXo91nLONUsnzkpgEFr+ce6RBt98lv1ZI1jGZ2c1NY2q
2plGi8zv3VCaGe2SqpFWNo5W4LwqsySDwAnly/U+rdf19xIHtoa0OHkhwUfqSVIoFnWItHlvqsFh
XR78tR1Fdgxs0BCU7eHTMyvNHJHYd5nq7pq1TtOmySnwZuv1IZiMs303/YWeWjgrLQ/ggunZev3T
PXRL1VXlD5QySH24P3SQXNSRJJQ8esVM2KG4B5YqvpVzD/PeWlMhTidhLLrSmgEasZdEqDj16Vfs
Gtbn9crvlsg18LD7OhdOcvulZa5jpygOurEY7alucyxaVg76o3uPK4gCmOOFC8fBsLEvhZI97ABg
zqkdNl2Vap5LdRxxPl0rMxEpxkrnDTHeUSpWRQ+bmNytgjo4v4YS0mYP4VqQjCG3+2WIOz0A0ZGJ
aYsGBrnH+Vmn6xnOS/HCuLk5KT9k8scaU1uGfyR/0oIAOqj2Yf4BEb3bj5Pp1x1cAb7RK6LIpizw
vOp2zu1tGOcOGjgT/lZaEpCzSCwgl04cAwLAOs+Y5NV5RDj9KtYFtOx/H62rEEKTF5I1l0auo1nX
dln4uvRc9a7R7uupjDQ0L5iYeQSgEo+1EMRGtp9Vha4wjlBXl9rvggj7eGIxbM/sfW8VBjpbXtDQ
mTVwrYK/xyUHBXeDK7AJkBGag7/9KioOKUcjQaGeLNsRqMLr+4LznIGlzK8x/X04YFxwMcHbK+Q/
4CKpkEj/zTIMpp2Zw1WgmQHdflg4jg/823Xo6odn3VQFeecokrK0KZeqcYhvKlZyGIjjl84W8w6L
/ivKeGv1WlWLoJXUyzgUdsiGavI3iKneuwcWqISpSnSiG2eDpe6qTn5LX7dOOe1GU+kmeukpgqe4
hZCknlfkDy03u/zFlRPc2EKRlW312jIuutTlCkqDsF6SXgrclH7hglA3htCIfho2Kgf+O/+oxdXH
5vyh/lF8zlSTW+doWdJ7W6fYmpar84zWSIpKGTOSdqg+c8gInhWWXBpF4MAEG2vMiy2cPnz8j+jx
YR1PkHYjCCtWyCsrSoF5BQuR1qTrbQ7hEOcwtCEx4nbjb5ALGc9Kwj9Jr+YptI6G/B2B7332hs6I
yZiy0dTNagjradFyKYeyEOBZ4gS31GnieUawMlIpeBZLRbPQxAxVL1I8uWJeh/IfUnJfCGF9vY/W
3MPOX9Ro58TEA3BII76W7LQ7LVYnI4q23VEwfXk/C3MJQqJDBS9T7V/J9Euovy9wAinIRWcQEQQ6
SW2UNOxFdFVhJ5HzIWC9MT9SQDRPxxTgz9gJw8vRntKGgEGjULZBGPWWrt1GS3AJNGpUxhJCVcZm
nB8bsnF4VyaY8HgA8oJGDHHPzoNq6zXf025djZ9XNthop8pey1MfqTXcUPT6dnKjIRBZSnyMYwBX
huMmmp3+5Oz9+SWSOP9pGVxvD6sEgY0So5R6c5+h0m5M3/cagp5tANB5glT0aOKNcsZUjcFjZBIe
4hDnbubeROSStVCc/ZTi0uo3adA/SyQZ2XAIabnVYkCbwVnc0dnmx+Y76bGgyeiuwi8AYg7yE+TX
nx9BS7s/Xu70KWlqY9t9LdBLF/WEt33lSfKytb9Nzf+WL+BURFfSNwDcncrxcHLj5Yu0JnFgyf5p
zWe43ybFOPoVIQF7UeNqP5rNwBtK/OqFi5pJj2NbB2FRP0dLMKTxZu6c/5w5yPsbVgAx7BH4bZXE
pDj17KvQlVCbq+IPmi4Ou/Nj/6Oj7YeGTjzbqQ/cPposwl+G3Xv+Nc7pO4cIRVNfbbtdf01o35Rd
YK4LBWYoqnG8j8uPUHwSeYHT6yVIWQM5YCJ1bvGIif9DzYT+oM9rveMGRG/sO4OZTVLlA4G4wDrj
r+Sm87OOwOmUabWBmPaYI4WEXi1fpvEX3c7sa5vzPjWjipJGkrF6v9Bt3xhEGRVrjf7M5eC6h7/h
x1KR7dCjLyCM3JK8vIlJr48U6pVBkFcgGVUmyFMDpllGByClbp+EshQ6/tQinDUgqXEuEsLqeXxX
C1YA62F8gkre7HtmkCLs/fXkKN+h2hkeH0WXZBCOx1krUJEq8Dd2Q5TGI6pmA4Qzs0sr76kbL1MI
rSCM/DA18GhOd0QQm6pAMToAOV7k57i8hH1JFYae5P2Fmp51GpS6kdjxXnL2434tI57+5KDTeF80
nVjaXYEkqX1IkEi0iy0cIWYA6PMuHitXa5hFt5hVhvJ8SCNEN5JGEHcFnDxDiOWzGywxFAu8bqiy
WYGeHw27vqDQZCT5KQ+FBH1GHENxexXkOpRJlOHF4yB94DbpGvolmd4SxUkjb4q90ZGUNpwasXfS
C6Ng8TIS6WP+O5ETK7wk7briFPnpaNTlqdJv3R/nsNtU5l4xBGzAZhUFd+oeWdYdVVwGHE4E57cV
tQ5q8sY+uiVRWLtDD9/r8Ya1wADib8VkgmAHgnuBsr+EA+BR4eBten9pC7GPBAesqnGuSDBIZ+uZ
Seha5t26cuyLLqq6SvAHpAjQ44o5JVo2BXttVQwcPbGkjZrjTuyz7gRXjh8SD9Vb185pgmstZy4n
4IPOuh6stlunnNyBGFDjY2H69GXMhB03OsY6aWJS2Yue+FHtSZpYSoezP85GIuJ4nlnUMJfubcay
ec91+AJGSWMtUAVlQsva4iir1Ac1FAT/OPWdVyU/CtabMqK/QNNpUbVMt8uVjqumvzbRYDO69kuh
OPqJ2ckEZA68vLnxxH6pd6YI9WAcPWAoqTRdfteGTRV1bUaGlcDgoUsGaspYpJdKkhfJHrUATIWC
hSniKPeIeH3tlmoZH5jesgfdcRFq9sBnUERDUtmJXGU8x7YzJZpULmif3+JLHcQAkRpcTz0IPZ64
iO7BXJ4eVPyEMkwqmZFwjhQ7c35Vzy7hoZp6Yjm/5utzTNMwZoTkWGEtKS60NHrtAc2g9p6vTXy3
crshVi/4wuhOAfMkfEBReJ+pTZJF2YKLbbx45SP0HPjuHZ3sIeHc0UX92C01gZ00sUy9b8D56xpv
BNFyzjl3EkL/tmKryRz4jSYN6gHEE1I5EppLt7MH+9bxs/t0WhbK0bOwn8HwTeTnPgcJ8ir3FkSF
3n20ZEmhCMPXwFP4I1B/VRVHJIHFHUnpy0EuDZJSveH/GDtbXp8dinaBU5CEbx+ik8oiXRHMXmSX
8FDsYC0t/pJqn9gyTtMBaEp4uSPyyRhBLSa8OGHUsjkDjrlqoeyP0ZSQs9X9WeOKEPELA61zcDgJ
9DfxYwHDpYA2VC3YM8NObtnNShE03SW9HMCvpS1rcVYlUQmh90QmYHzhvyWMx8csajTK/EW/W++L
zakx/OwJxhqMfo8EFVMAti+PlPJtzcnsKfnxOUvTVW5nfctyemS65kOWms5HeD/OBk18+tgM6x02
KvJ+ylYStBXxadEvg9ZMQbHNPxYdquMP61zylcj1WNPCjfCJTg4l1hmXLwipCsBvYXKLU4MSaBxP
Gg/h6oZnS0UuEaMdxUp8dfrSufAgXvIHx0XHCaX0s+KkPO/qLaRzcTMupN4BQ+gUMp3WEA51hzIO
zSNamhEAB77qF+esn9/rEIZXic0LgPcdTwp8X4X7cq8Cfz6p/VBCDPQet+K0gMEKc1vpG9iuyoEs
lV8C5UOyL507z/GmDjcDMRXte0qrWevrn5Fce7+Qq1023hFah5KZqYHw33GYN1oBa5hzb8SaHDTW
3U1jeLLHG3udTicZoC3YHUgBivF5Q5HxKwPrUP7870CqusuOylGWGt+0RXvYtBb95qII5jVPIiT1
t9cDq4mlINUV5Me8C5g7nEcpXDycT08VZZ5Vlt0U6tN02w9bvoE20xvboC+qnuosZagp/H31vNAT
5fSbUB+C+yN0NQKWOmVJ/+e9eyWWj8bLVQSatsD0WTRUKhME/7c0ZX2eplJiB5KCAyz/TidU6vZG
aZkPDSsTKj6RIT9JMImD97cdcLy+GxVhVHPNc7OoOUf+citH+CZQ90LEAo0qF5pgZ54qZHw8JnRq
Mlv5zSqmkj9CbBjHQD/3R+iLFmrksiHx0lyNss9F0hgC9JvWSVTnCK7D4alfZsn6mNs51r8JICJc
9Azs4CTYWr3glxtf7+rpj+Zggdl1Ai/kADn4kueurW7caPQ5w5/aSlGmUQOIWHvcVmmOwwEnPlom
FzKTh87N/RYeiVUZ7OrODmOnXE1IMUGMVmKHYH1ICA1zdcyLdwfpE/VPn7Elj4hmHk6qpdmnR68b
xV0JbzVulinKyY7apTCWOSm74i/aJI8yBoFulsaY23q3/MsIvTBB97Z/vvGMXZzUtXTzEGsSC02Y
5N/qFaWiLQVbWTFdt+qCu2+0jl6J3MG11r9HXx6gA4w3e/qYj5fYRpPs+1ig2rw1TfFgYAGjDmKz
JryiddoMrWfVcJc9dPoRoYvHalKx0GY4KB/adiUr7z4GpYU5TjdgXen51yjSpWhEWaTKQFC6USYT
gkNDo7oI/R339njHuxhlbheHDPZuA1bjjbp+PgZg0LcjV9mASWsAEYv5GU4YJ6KGOyHI3mgPoc2T
/aA48GDVGQyrH7cU8K/J0/LcGbSyWtfrEkOSZx933OrkqYjw4jKDW1GpWgBz424qzaaeOlGffF+A
xBH9sCFDvG89VMAPVEItZT6JPu0NyCf/cJJAhylLs5Bb9ZOGkSOV3l3OcEOR+crxdmnvWVPP2in1
UUY75aUtxTgp8LWmvtcZ5qUIM+x7ERzP1Q61ZoOmgRO92zjCLQM0FX5usjN4IrrDWj7WJVHCzfqu
WKTnOT1HbGaSXhglCZUgp6HJ8wu6HHuKDFxezT7CSal5CHROM7vbBWYH5y+6cU1Fy+0asWeQXG2p
LLep1DdQc9hWU3ZNU14bxYojEkobTt2/OtLwCUZF8mheNmxmhqQ4nLp3e1EGEpqA/eHSDaG26Gxh
C0T/6i5I9Vc5GjPYWJn9y5LIURvs1dQl3O3GYthvwWeEJeXMrteH+z+PNL0vFBNMZC0dH+c+1v25
Z6orqAl9WvuqfKR5LOOe30IT8sXn99VjcB29FjHh5Zgk+r/OEbz06+cmBK1LK502OqJM3JAUtUgp
9rYYWe+povCCkjC0LXeHKaOGWkfEcvISZldFs3TOwNgyFad45VfYhGUhLWMqvt7zvraIMbs3emDR
T6sPB7yoCxFccsBHJzh5TQmeKVtFGDM7/8ANMPB9FI52eKP3Zhm3DbD1KDfdX31k1pKmy+keuUlF
JVmlHMiu5tMCMbEnx0RPBgPggfheuibN3cQZBbT789k0DTigtrhh+Vx2Ep9k6J0zl/1Uq7C/MLKx
5SUeP/F3I/Aydxv9sY4tsMo1N+96whQhgbmll0ymE1uxZG4PfmxyYgaaYoiig+Di2nvjVBQfoSP4
TbrS8XO1nljVfnFPX4OY0QYyPuLqYNnXp+QyHWkrXCDDDhCcIYFwrA0jdMnd0J3Pid5CBjxVjgMn
6WW25TSDbcMNwt2k+60oI/aBEo34hCMcgpyXgRl9JKI2SDYKtASOS1e/B/nIuNK1MG9YJnFhz3VU
rpKhi0kEkj2jblg3USMpOx05V8mPh2uylMJNNUflzwztueiMdmAEeQdCcO6dBvCiG+hTfqB6sv0R
9MJUPkGT77aHvEMeLjUduBmk2QW14T3TTAPOEUbE+SeMELPfKTz+KUEVd3+wnQPxhS1n8kGJ8PJ3
oXhLEXleDo/Aa3ZSow1gTaUfLky6fM5ZDmKFy/ZF83TainenyHOpm5p1FhEmZfmMIT7Z6hGk22tP
1R/x9WjKIllxlrcfsnZZlEhT7qmAXn728xGjgqQI+yV63E2NfBHpQlnblhGj4kvUqJ20ifb+Mywu
pDqiejVYaYKS5uzx5NPJ1ThcYj3uS9zV67EQKBUbuQje5zZU+qJ1gV1eLSP0klcnRpfz3Ux4s3hl
f+2AmWFKAYKnbxVVNIbjy4JmP3gf4ctW/h63kZTQJk5OsdOndM917MuvSlj1ttDExBMIkVWNgD81
dm2YQXgdKxQgRfEw5vHBe7CiTQ3RipnewOU9oxifet+UzI0kfRrW/tIcoIfxHHcxCYpXrEZlXgfO
EhM0Z+4Wh6aJqXzxKtlCP7oluQLG40GyZVRPJlFd1DljnFiksxxSJy4ObhdIdaeiT/hZ/BQroAEG
SfqaAeVMYqxhgIl2TB3+8QN+xC4eiPdfwstW90SsqtHZf6oXZ2rmQqBEMjz2AZI9ZWXdMUMjENp6
wA3OMGg5E6hX438AxMKAEJNYzzZi2ijXSLR243ALydY9vayPvi2yGhuJeuqtTKthful4FyzLV1wO
c0HpPxojGDvbYgJNocil9vzDl2kmSNO7t0Hqs7s/LteiHWwszAUZzlifDfOguxCH7edX4CT4q4S4
Y8W5rbM95/dWKj4MbaY1SKhAUfjmNyyxAkjKUR80AWDfWQGGw3B4sUoDgefAdAKWacJ5V7CSzzvr
snOP6lwPILA8ndiUfcFpCShL41qd9Ybg9kX4eD5EPlA2qmFEVjdQXAQ6SQfj7x1cvpwysi1XB/Hn
HGtRmTe2/UcaVSE0f3zvTZVm71X61NFe9ed56H7U3ORps6JWQkxVRyj0QbN7cCsRASQZ6vTeX3wh
shnFQ9FJyfpSZh0cEj6HGM5GoQweuBRhL0cdgLimHe4tH3d5Gs0e5a9Hs5WLJkDQYAvT/JJ9SxEq
YzjJpDmw88LSLaqm+dJDJmb7R+p0EMsaqZ4gc6WolJ0kJfXSQQNGlvCX6Sn87n9+E8Wbszo9cSUb
bPMI3yNgmN4GbWm+IWqqPWWVvFMZTjHyV6aFzmSZmIkTq09KW/g8C8kKFtVtbD9sHo03cFhkC13w
kRegKF5BWpjJL6uJ16imOLTRbyMX2FrC2gCanhy7LcJeHT28OkTF5ulSUo0WE5XNu+ywkYVdB6nO
OHLJe+dh7QNliR8hpbvmeVY6cY3Lolwm2Ntelt47n+MJK6sYaW0b7hUxc0gzdPw3sll2dScw8CZt
CRlR9657upXbQdQfMKoFK0bvKvSVzMoyJit2BSJ2cro/yOhqdlacxpgLWVq0WOegj8Xn9DdimjMW
mbSe/8BZKeJGOK7/S1RImcUQYSRgP+Dg1CvJUyOIj6PZHrQTt3dywtlZxXEMQJMEROU/qyv0BcBU
/7zNJtwZOBvS0e36hBbts3T9WgaB4kiyIzS53VvXeHabSynd1J86bTvJ2iYqxoxWxHyADd+d2NKk
NBRMzKoZbAbNeOf/YdhLWcDj+lGH6TZLxEaHiBZaBOgNQGUkL6eyNGvgfuI/sC3xCzGp9k1MFHSw
4AlE92y1Sg4QaQvZ3XqWU4smsfipqnw8x5nkJztWzv45DK0Nrjy9im6GXZREv29HzCQCYYBACz20
1Yi59msnjWBkGnJWWyrq2temcVQsU01RbozpR6rkxROUgJDVIc+R9XQmTmWBLz3sd+bmIhz/HiI3
w3JdGVqTcp3iBDamgR9JA1OgSHgc8MoGB597y0EjtcN3VOBVQQjVzLiGuiZSvSSVkOFmDofW5QUz
IB7Q3XIzQAI9h9SieWAy72haRP7gotmKQzbfMMlQg7Xq5ijzmismto7RLRr6Fp32mxsmAIRhlsTd
ERy/VJVjimjy17Ut5VLBPRbVpxR53AKjJjfGeP9pR/xlDYuwv5Q/7ElneRD6eXjBj55Y/04RxqiP
TYrFdXqdSw4TD3YSFkiS0F7iUGF6Z++NLYPLynfdKEyocr+HVN/b1b+btrgC2nxQirtwHyYW0UTy
AirQpnW5SWvOLXg44DqVCENtPcHrh5QX1hU3geb89JBNa2f39XBJWzA3VmB/i9B803li4vAkChZ7
yY91jnEDA/B8vw27UzxVhqfWT94ttV7W3ZdZQtvKcryyWfml/9lUxtwwEbWOCLzIH3xqV2pbpXFm
wHlXa92y66CTE9HwVbx6H0MRFVawEtEcpFNi9s6lggRxtTO2L5Kti+YPQSbF16x1O6BFk1nJ4SWJ
oka38h1AEybikuQ7s8+7gqvJnN7D0PJh1sBpcUo+E9CQYU84HXgdhehdWo929P6Gbi+F25MT9dvY
fA/Ty2Bx6mRLb/3z7wryunLGWYhAZtbb7K1M9qpBsU8weck0ebTkIvjPlVb5w12P0OLyY/WHZImu
zmr/iGbrWyTYCDYzTQ5eCZFutletO1c68XUqmsbQ5geGacOIg+64u/gF/v4bChFYPwdf2S3lcS9+
zAYtpKVTPDXj+XJUMKxvvFs4veXhJ+Su8d3ZiABEVAdrE1OKVzNDLFw4L5Ce4IsLNOu6c+do+V4V
VGBlF2ihhh460jRMH8e4McGEikaZcQhc03uuJSKEvjBTIrmMVWOqb7TxExh7bhJ9UPHT94l24b/R
wyg7ddMciWFho84XtRfvjBC0neq+1l6JKxk+qgSx5TrMtjXnWtQ6gvRNbi90HJ55ZJj6XEZbhCtS
4XxfymPRZnb9ao8tiZpWCWHFdM+0tEcoVekP/b365OpWR48GpjmBXYnHBjb5P4aRHf9/Ou/Ij0Zz
vDA75R+W3KiTcRkAb4mI6pu161dHpLH8C96VUe9C0tBAuq8cAae9l8ffIC8LO+rZbRWhyEZ0lV60
+tK/vfXCuWmxz1sJYAuA8J1EOJ5bZjc+8pWgi/gAgRlMNo3mzeXedda8qWCjlT8h12hsLiP5wjok
ZcRNxTNmrioJVFflAS7ASKgO6c+qMLEXZOCzBB5mKfC4Dh+qDMeYbMyDJI0+H+iISPftKfm6SgQU
R/O63v0YcztqiTx74fncwQE1AvlHdkNq25A3kIWX2W/iyz3j0yQPMcOR7StBkCMLFINTQhtFFGFX
Vk8jAGkz0lkHmrUyX6DIPLc8BRWlPeDWF/PIFrBW3lcievGCXGjFKyX2ehe0KfDB2rJM7UoGPLZy
j2FFrIBq1wzIFTeim0GR26z/ABEGv2fbXRTgkRLECXAki8tHu/Y7Gi1Clr6k8m2RJkbno3frzny4
oFYks5mXNrgwzze7d4MxkKkrtKieGs1t50/aflFaN1HIi4sBjf9gmZMEE8c2axzzernrNAMb826h
5KYFtKrS416fwDtHvbhNR+EP19mjg2fT7udRytSZqiKHJz0cBzkr0G0i5gj0ZhzLnZiBIQkeLMlx
mET/QPtknRKBcCcFlJ+r0DvscTMvB2lmN+lcPAnWAK61GU7i4r/DIUZN4Q8SRi34rBg9uOZhhNst
oTrlgtK9XKk1BpEmhUwsSeTsLxmGfeatVMDBOafIJwn33QMru9ZiJSg84cuUpcBW6D4hJoEHAlto
q7b3JKJ09eGdjPViTvNdL4RLWxleM/76eQ5WAwFyE9jncPP69EZrGpnunU2WAsfm6dqbZv0Q6lQN
PXM1tATccvBc97GGypBLFIlzNtlSGLBHpkUL1J6/ZxKD3QhfGJST8L1RjhmaVqZK00zvAEJT/m2q
x5SxLLNZaiu0FF6I2kvHiKct3szXLF0Pn0Uo60LZ31nAvMOvSaqtS0no97WsPJ5dK8lIelht4Pmf
tKsQTQjqFXXEhsmq5z3joxR475dNs2Koxg6L5W+TQa6wkWxZLCBpJmYzprG9bORSTg4rwrXAHG2d
tMbtj52pWmB+r0wvzhVAYZF+V85wD75zaMwBGSteXQ5ENKgWz3QpIKnvu7r5rJehy+6HaZ0Z07Ti
9OqTV0HKih7zOOwNcm5Jj20Gvv77+M8YFQ3NZ52zWBw2JVa+3pFfhqUP+/ewtk+kMCPY5dm8Iaxe
8F7yne01oFfO48ygBpRyOIcOW0IGrXuDjb/qrayZXLfH0cWwZ4Lmm/c9koiqlNsqqagCq/bSjqGx
+NN3/fNjT5M8JK3+eQ1INZEXE7+t1SEksJtYcomx5akaxe4glma8575m5cCtekFPBuRjV0V67l9L
gFqEkjEizYigZlpffzimMPx+RB1XRxNdUlA5D47ke2KmovOXf5VAD3sMSqGkCZNcnydnTq2IK4K2
RXpTXm9px2Ako09wcshjlEWsITxvpVHaaP1OOkFoyzMXgdLRv87F3DgDtbnSt9Ic32w33E2XAIQZ
T2Ol2Lg7jbWja50i2hm1Fmgsf7NdYiHl4PcKF5M7aJ3UUaEwIXatusY1MaKMfHMGttssjZ3fQmnt
Mqr2YN12npOcsfRwF2D3D798hFAIPx0EZz9blWljplobEZPskAH2m0IIxjjrV78ZEyit4UGkHBVw
4qPvME3EPJFNgjJss6pNsbwsnFhOIE5aX7SfuFFL7OJ6tjQ28h3Bs25pz6XaH3SziIilw3XPIwAt
7Em/snIiEN9yU/QSrsAoeqpRj39srr1N63TOm6Q6vzCb0KGEvnZX5rsMQzJt+RUxo/Vr5mH6LNb+
pCz/BxFb3vrpRCl3iuAl4h7Xp4uuFxRr+mE4tTuLqDWc8MBhkCzza09szeM77Ltr9k/4BqQ4GPsd
TFOAFZCLwJZEDLm5+56J+FIElmunyluoAjvQFKZveiWl7ioFTY6UaKyGmjx0yBhB4Xg/kfbwGAWW
3JDH0EOgewp9ehZ2ETnqJf1T5vBKlV1N5sfQuupl+kdTfdaQHYmQTcVa/noiPXATEs0iSL/7ntbT
hgDRTwxPU1How9+qJAGcQZcgKCiCHD+oXnllXMh/8yrpWI/pcT3U9nWovSxPCAWCzE37ZW+JSRuv
W/SSY2QC4Eh1EnBpgqzB3SnplO0AhMDxRKZScOfHhB+vapKI3JKy8m28IzgM43iToM9suykArFen
CqZrXenDTF6DpMAdaakrk6HHfF+xSCj5GTWNU1upczDs1QXCRCF/xdtvdgxMhM7Nzmof7YA5T4Gz
JRujey7Ln/fN8Byevp2z1a9H/pVSKmvvhzIkMldqJjQCZ3oGVxnHGLPSUeFlKQ3NyQ4T9+/uAZpe
cEMrDKkTuM2ugLf3vfxF7EuhIUmgaWdt2qf5BmceiJfQzgfrrgF23pZ6PmhO+vvfeyFG065/qz0W
wH7oT3VuwcU9DPw3p4M2UOeEioi0xNPZBJHTdUR1zlN6KRtR00gK6baS4DmGXk1gGTwc8+uATAtH
vtLgRq34m7Q/XDUnuJCEMB6lh40xxfMrIWAHUd+w9TyMeeFQ9pUyIYtKdhvji2pdYPMeg4Y2cx3Y
mOt8FRWKWAOYsfi0ORIVnc+NU8X6bMWqtJV3c7PpModVcnydNgeA7B7HIT/oaB1B0qd2zjk8/x3N
eeQi67Kt/4T9t5kFS63XKHCsl9rF7EnRAWrrMTdQv2DUMdUfySs5A5R0CPRPmB12NNESEav1LOlF
9ynGEOHNFFrho5SbTDnwjqaYzTbNEOzbL6ZWQW0ucCOAroECriefyT5jjA1jz9aBbD1t34VO28Fb
dVDMN5/ZnzptR767Ro+RJhfwhyQK3hZ+2bDNovuLVhGJoQ1sytVeHx03ATobPG/HPiKksUOFiI+m
/+7kKO8XHIRnp8cvO+Gqd6TAKZ4j1m9uAVIhanYyqYA/95tngV/ywK3GzcgRLGiwqAhIhfAAniUN
yugmG1SshvsOFhifl2zIGea9I8d56dRrHvdNG23/ITs+AsOOIC7FStO3L9gB2qL7bDTz2hEEX19I
ViAL0LiSiW+Wdg/JX9b58EWKkANqtCBfCQqhpukbRUMcy4dRjUTH3yy320VP2xNxWb7QqhzzRh8o
Mm7zeLnKp02k3YC8vHR0Z7xg13lfngxNFWqDrsFY8smm3tJ9vX6Ls7a/ubp+rXVDz9lkZXFUnocT
A5uCQ6O7GDtIfYSz4KuK5gGoyCTTPnVHSb9igO5F8StIe6uUII94WZXKRWDcNE3iNxfQyhpXjmeW
RkbYEVXR32JR8LYxJ7JEdv0HyE6eoPoLefLRT6aymx5db+o87BbOVT+JssasjpYh5jOtb5jW26bt
Yf3jE9AUBCciXLYVfTUXVJNyrLH+V2TTefU+naKCV96uhp3q40KZjaO5qEWmO5ONnAehXe0oSzzo
fapAgp3lsU9yOcRdo7ON7gJNR72elq4s+UA7QvYpLzHHujyFZwevftUYKWZYhHjMfEO7RaFZePhL
puhqfYGQWICSFz7vdT7JcrE0OBpriu5xR/FIXzNwhiDgUyq2mt2drq8ILxZILGHWburZoDnaJQmT
TBAv6UC1/59vL27ap0PPFjGRNAGaHaet4qstwk6O8KHNx4EAFbvyQl1AzFEmJh1S/48ddbXuBY1V
1E0us6vClcZ9GpayBDRXqCJhmnGJmVx16q9AnMrZ6XAhRrx1QIhwO6rsq+EtKZESpTjmcQ5IlVRS
WiMsTYmc/CNDGD2fA431AKvRRw/dsI2vVyPYAJt+dVq0ceUe7bbAia2JPE3qQuTeJya0Y2nTc7Fc
kv+k8+t3uM+8PGTSisPEHK3OXuG0/ceHx33dmNRq7gGr2J5l1iAEEERFwrVknOXGRUbO2sAUOS6U
6urqHWIvKc2IhEHDYox4jGjAv8Eh6LFSsds4kJl76+iOpQnhWl3IzKOiSAfa/Y1ky3NRNyIOYZFy
KnsS3X/MAT/XAmbIfCP5xbXDTzxTjYXYQUOTn4KJGyteaPVyPIeABX83vex6q2qdNtQH59BYZm5V
6OLVgRLrh4AgVior6GS5kBK2yZ1m4vLdlUKNsT66Fxl+Rfd20N+YCoATDJ/JTELfW75SD4eBXPac
PJ/50ft7PQt57OrlJva8BnnIGhUivxrbXJkT00V8T9dHqygeqmPdyQj7OMU80c8dlfPwPbaoatcS
9J/RQPfwDCUgZMFsXgvzGgbHToVBz+m7Vg6wkj4Bw8IpQ09esb3RA7FfWdjy9weH4gsRErC3KPzZ
OheKMkpNdKbVRe6fHdh4a0bwHWVia4mnVRN0jQFh/BkbEu/UcEKaJMeOkF4AvoT0KKSQVFyAxRBk
cdwZV5ZnyJENUuSudOGg9P2F4EzzBnxHXAQZw6eI7EW8HHCkcop2rSXFou7oRqhbHzBxs88Kzlvm
+gkKwPRH87mNDrhr614U5XmN3feOtQ2XuervhEZ2mUFCwMH/7c1xM4JUbGzz3GvugKLwED3QGWVW
x/xwXITckUUa5DW96iix8Ukuig1EIN9zU/KoMm8qHebuQ60RnkWj7gMDHczgRZNHxCs7Fl6XjYMu
96btrFYcT31Ooa0tGMKqXYuTe3bU1xasHZA6kLzTlBKcpViLxLC1DGNzTby5Nah7Qwfdzcwfo/YD
unYgulJnXfKxPnTpz4Y+98YpYZK5z9KxLxAX8hXNouCui52pgglKhL5m75v/Samx/Fr0Y/dHZZzl
FRxM6opZMQCFmSEKw1iIm7xvw82AoEeFXj3FotcssCkdVkKcrCzww53RPA4pVklj/uWrvTeu2PA1
dcERVPZq3eOIA5u4fPDBwL3l2QUkr9JdtZDhCCpbQjmmZxxYL/UmoQeGDO6IUyVtY5sKa4gU8Dcy
uzO+jLWHmJMmgu9WIi848f9QznySFY3ox0PkHqlmYKJkwRRH+V6S4MDmszXJjk5mH0x2qYMZGW4L
nQ63S6EsUNVQeWsqsYSTETQQQdAoHcuF6KR7h60iN9U8cWIWw/uFprR+uvy+8F4D+RpQQDSkzd7o
xhzVKvxSpM4UqhSPTUkmAuQ7XEK6WCwLV0qOVL/3tAZp//KnJ2ByNDk4mzTDCaqR8UzL6ZmkWulu
wmlF3+wpfggSU6rl/cGFMuLycusAIjv1mUTtCo+cb1AEtxCowM5DJJGYKpyL7vr+HvIPuFIF+w1Y
SMfobvv/mLyLTLiMQO+REbmL0OniZoTCRiF0PI+aavbJBkgdXn49UeYr3lQYoiG0tsYw9yX0LLOP
R4Edot7Phr4sK7Uh6BxS5txmFS5Bu2GDyP/hszyelyrJ8XHDTnhAEuzG+8gFX6RgSYbBCYja5kVC
jR4u/TaOGQW4vA/m5g20lWFVMfZvc6iIPv7+eCuKcUq+r4OeGf8tvWywfercNqIRYrWmv/Zh/2Fl
wsYzOS9DYqyvdt3iUkEaHLUSAWYOv4yVDo7bN3Hiy1q7oJ1jgn3xSHLWj/FCgh/65PjawL6Ax+Fe
lU0u7rr06uTVPgSaTRec6+XKRr/g+/dJRoU093VDFBp8OWrBS3bJQer+RfI9c8CwitNoSKwQ9sLs
XouYddd9VPqOoq/dgEJNNOte0nXPSXkpy5FSb5MA0X48F66kntRSC12jivTx8dpRJWzbfZRzWYjj
Cg/B6l+Pn/NGGW167SLAEjZGdYeBMhPSyRGRoN0FSuzqWIl1GzCZvg7t3Ts9Onal0AZrQwIg3Vrm
l64sRPk/QlSvtHdYXQP55q3OwtL3Jjl2euaXr/Ko73yh1u3aLENX8JSHT/IT1e8xOoQWqPVKHtii
SOSz8bg+aysKNmnniOXNfs3TtNXpzNeJMYgCxXkPmdJT1aV7eaRy1v0fWmZ72QlmWhAnNa7qkct+
50WzTEUdv/doHK4/llZ4n7syHX2DnRHnT4XyPoC8gQDo6JvCY9oK8iQfYf8jsUIomIpH0oOFTMoO
UCSY6WQqb+1vW15izB7G6kUnKhPFBT1AUvU0kaiiHAvxHu8hpdIDk7QT4qKH3HOTOetbpHLXI6/p
p45l5j1XxKMJ2y2THlGoEB3y+e9p78Ma1uKxnpNZUdvVa7SI2Pc2YcOO5SvM2gZbzJpH+C3wpJ2Z
PJICFAVvjyaEZbiNHrtDX2BCVQhQSrOQ//gQjpgDMMqPmxnNf+yjS4ozjdMz2IcQk+vYeF0rih5z
34er4pBS90N/ef/1Lg9OM+ltZxWeVxqldIihsC0XtDuQnX/I/YHVQqqIeawp8lcuzaZlrnLzFCBi
Qfnwetqek+inJj8kseobvumArugRtUcD/dKqSix7xApprDzg3sGOcWA5mKLzknysbqhVMDcgjNIT
/E1XTLCUGEVh85kkA74GMyXdMUifD5Fqsv2W4GrMOenPniF2WXqWmGSgGKzAxcUktpZVLhlFEQjF
rAr4UrFCnygaBeNm41xO+zzRrMrGS25NtTnFjz47wsS3lrcYeuLcNt7OoXWm3tjppSS6dPD1xYrl
ot0giNulvxCsmxcqLTsRKtU5idHqroUMhQhlHLQWDpWqW+BhSRXLTBmMPNaSntKiRHSB48kPb77H
LXJMluTe6KQLIG1YYFWLbiZZGf3qY+GyAgRM0Ghi/PJLIyq4gT5AFPm5Xjg4477oVbhgJ3KmaVJK
FvRGXsqZRohOY2v9weYviCOahBNvgAtq8ZtzstcqoY0jWGL5USZYdZ3sSDS22mxc4elT6nvnxHiE
wLOYXurcv9xTxGyKPH0GVl+jnxyBkNFeMH2nHlq88RrHWD1nmMq4cuwREi+wA3WCCOPjL3+J2wJ8
RO0JzAFe36Ik7EBTXhqeqDPzqAG7ct+UmkT/0PHkKgqKkWldQdwxHXNBys/I//pULJFWtQtoomrw
LiQ9R7ogkJtwKrBqd+17DHnWPtrcLjP+vrAnOYZoFPKTotfTRfsPEQzxhhrBK515auNyeUZFOuVb
d/U9YmRmV9WJQppkkxbMeLwEES+rL2Ur3UY4VD1YkByfNLklCwI7DNe3a06zgKB1ASeSDKLKR1jW
UBDO6HCEDvVjObBmS4kpZN9JiS0D6mKTyrF3NEKX8l/zwgTn/Z/N0aMB0c1O6bgU52k5BNq81xAx
0nOzfeVJAhnXpDlP9gzeNaF6feIkDnhitpBXss7IUdXWkXVMa39lGvXfcGRPDKzOab9qZg7jndk8
vuCm7m46OpQ9ydLvpa+vg6IXP5S+wGMHWTFBPI5/IDkKwzxUyVFHE7JuT72IaWPDX/UZ5IpGaUlQ
3ODM1B7SJWj/E1iKSiBtaSYjBrwxOblhXSzfAV3DYZwUE96Bm4qbt6VN2Q5IsZMehNPeG6OH5nOB
9hooF1w8H1Zs7bn07btQnHSo9tg6AlQc9z7qv24jWH5aNSSs9KiDhXELRBygkbcDYycoboqa9PFT
Pl/EI0vbJjoVm2YHITh80K2f3Y32B32w4+lzC5g3sIwue4VLi1Ada1p2y5WNVLZPhHPI4P5izjyk
qptB2Al/xJzcuJCsJtK0oyogKAbekShFWlAt5Or0jUmJ9VoqIJVeU4qwFOqiTl4ZWOawhQxdlPYP
nL5XB9v7M06Y2u/TKYVFuoy9c6PU1cKq5wr8EzPH6g20y3ryiF0nyXO/olPije51HcKw30Jc2gn/
z0Iq2MrgCtnaTTWf2LS8ehp6Y7hnjLobFLusJ/quizt9y1BLqqcC6Ey7ovQjmrQKOLzheWmcUBz9
VS9eR+QLHbsCEe4gK7sKUhERbF8cGWKiWLkYLwJZvSdkuUqPBJjWTEp1UBr9wBqAnZEFRE8BiY+E
BU9o5guuH3RQEq8lCCBEI2d2xT+z7cF+LklATS1TuOLVVXuv/tkgAT9QMHbBmJoybF9mnz7mN/MZ
y1kVy5KZXqWQyhv5nfecj5tivzCuUHuoh2RlRdtfrrvSsSlOELYTrgNxiykfuM3qfFJ29oiQ54V/
j63I0R1uX1g5+jb/ddSEFEiPFuYpg7/+rpz35EpPAW/qqzw8Mj6VxrwJYUGd2OP87ra3B5Bq/pts
9WtEnEj8XPJdTBZN1Bxx02OUhKBJ27jctMkV/HAj1rA/aKctUFjh38BFOTrVfoiLKHReJSbnUBlF
1tSreexI+H5cteYGNVUC14lX+s5SAESO3HQyKaO9KjNw1oTydczrmbrlIBWaKB0EfSSWAn3VGcDx
H5oNpsze9x/NB+NSMOnkY4+yYPCgxi/14K3lYR/xRASUGo6XejKLXTewJ5NRjA3Qr0bmYPGBAo2Q
2nh9VM4PGkbLDoSi+Hyl918f5kWm42dJwv3cT+QEu+3N7K7fHIZRpz3N6g3CCZ3V808Kl4i15+Yd
IgID/UB43H/0HEp1rM5lbj882aTbP0aX1UIN0TF41sq2w633b6iNf1O08EHQPu0hdMEwndJ5s4JU
Hwi78ikQOQETL4BStiZgebjO7d2oJwSG/pyoBZISHoExkTrmzbRUokxKDiD3x1AXAU1RPL1Nod20
X/Yft/rIbdQruIzUJSdRijq5lsWQciom/RRDz+AOhfqeO2G0EIZGOuGnGAsuTor8w7WK8ClWBuoM
uxt9HPNCSvpqhHoNXJ2EZ+OYHLS+i4DRJTiMuv6rtyneVTgTDebHfCGCX0pmOVofI/2Wmbzpq8Gq
8JSC8fQd/YYfO1dYB4uhpURRCuxMHmjdp7f4nnYdbIEy+sFFHZ3PoxvAy72XBXbbP+kHiTUm76vN
gvnPVu2XyTrESv8B3SCCe4BscyPIcZo+3KE35/ya6e4HGqoCmeBJzwB+xex2VvjJvNuSDqsqOgte
8OdaXhioNC+IlmtLdwdblmVqGcDrLHCxXp1MN6ibnRu6yIbwI8SWcGaeTinBXSlxYz6AkR/p3CBQ
jhCEH0+vtg8zO8drs3r0MDyk8F0pc+vl4eYtVRIIN+2XWHsLbgK8QIL5/TDAAe48gyk03yBSIwaN
PO0SYa0YjWFkNdNITtl31RBI3Ga4woa22HwB4+05BYXleT/RksFK0nNacIn6HCfbAL7v/ykWuOkX
cDg6+kubeHKAC5lA0w1gZWRwNyqpAu2xCxvzEd7WzXoEkqF8+akkPe2dY+h8PrhjGSj1UbjS0PxO
JbCYf8tDJBwvYwNZq4E4iEYTkPuuhjr+8OQ3tfxzi07yjOZ+fukg1tm4CtxKpe2wWpxh0XeX0EGO
PC5PF4tDj5jzXZhLf+/ANvdKtezZ9Hf6Z95M4G8gn+hLqw6YFkYh+V/VzlwnOYFAco8CcMSlRStU
LXVnu+MlV4aU2l9jOqXF/7ti1yaSUnLg1ETUeVzkEH4qBbsinmGmULVkZHBbsb8B9Flsk8qis5Ww
lOwpucFPgOlAjTOCLrV4FrGDrkoY8WN9fe+QzRldza3tb9G4whzHjalQk22eW5PtHQBvhpfxqoDn
lZMsI30z5pPO3zdBs/LJgijQKxM8/CMJQuUnjaggvAYvMO1oxbqX4ZLM3qxHbdKhYrkBGy+zWAow
uzzaANFxPDIVldr9xBWWjfZ/Mi833PCHlhBmQhfthwTbknx9HBKbAp8MxCgh+jPSPPHDl76FssfE
MU/QUY+DnhTCyjmkGq8aDvjelsKKv8DcoP4bS9NEScTNriS/bKeEU5DzqSTlsBnyUciEhTyQMr9y
PQRzhv7c2rlmah/xtdwrLx/A1J5LDAd9K2PWK1a1Ph20mzuw+bhU467Wp3UYUHguxuhQ216+kYsQ
AhcJR8nYDUPU4IMzdRssASSsPEhq2h95Mst8hZoaJ+vSpfBXSCc0rYJDVjg3Zg4R2rLzifPQpsjE
btEGvgIb+d8Q6R90w0n7XS+W+xtFoQ4vgz8OG1rkFZvf7nR1kXJCTBwYRjhsGunzpZG9UOp2Eb9c
hulwCuGaWhNTUbiQl/EDaIzYFox+fcE4krdnPnfbNB9IDt3aNmyX7fj/0QHB4m7bDJX1K6WuB43K
zZqhU3Yp36z84wz5G62IDi4WIRVco6qSwHdUmxEdBbZFhttlPbh3E6svTIxU+89grqwS1JLthCp9
x0dJv5TzC/msIwdWnzKTwf4nLbvAZYsTitIq6jtuOPW862U6Hs6MZs+Gru+TgYbMKuEbdqYgKt98
in5tO7YF2BgOMZ2rx4xJOTc6nqHOpfbqUjLhPQDo8+N4NqenuPshQ+2KuiiqE7Siqw0h9BtOAcY6
Jjlmnj7dY1b4WKEYR3C2mgXIYBxiHt4DLMEbEio22dX8NwmFRhCj5EXJkGDBbzTOAG2goYX64Zs5
/Asc+ffEbCIUFV79u5h2UV/6s9EImmWzC0rw8lEawVWJ/Wn8NN85LgSFRAZK8+/ZLe9mwRLqCOhb
4zR39Hs2zy/GTBhtkBYAabZqAm17EUKv8Fl7oDY73EoCkL7gwJg/LFKMtsHTyhKgDzXXENZjFIrp
MPccgc5pa+Pgs0uOPciy8Yd5nOMdiXZM7P3NwNqapHUPCsUImJgaKmo2lnjH4CbfioLmnCLti7mh
57olfrA8hPeUGMYO5hrioOx+hWP6r6j+dkb4cgVjtWzvoK69njsnzRoLNSjaRj3CBjyj2UeILyYu
qk2IrjtwrHTCpurmXk118nQMZ686JAg5w2OftUBhrH9+TYlGXSTN6CJVad+1KBcUfSM2RGgQ17pM
8zySZZ4DMK52/BfjSFiTQIstJlnFSmtS736aoJ2WQ6FuCiGhh835DW57piFF0BCh9mPIPrl7iozD
ZjiNDl+/sGtzSyZV9MEYJ8kYJgRpfl+ao6CAVcG4LolExLGJ8+D7NTUGSrNfocqjZ18HSaTcGyY6
nQe0xAx6zd91WQw+579FYS5nLKm18Y216Tnmg4a/JdODyLzuTs1wKvQ+oBT5hyLevz4TXzUwa6Fs
6h2Riiq9xnpTaEazY+3PyX9FkwTo8WmH3++FHT22Vqp5injIQJKl9urV61RPJs4zBLvoovhLn1Lw
DkPR3eVPm73WTIX0V5U9P0fS7f+dt12NVwrYV/IM6GAYKJHOnXMAXRoWyn8vX/ioj+eBRzreVCZi
9Fhl/tPxz9e3wRHBpI4VOxHha5MJ5dhuctcJACNCBc/E+jJNMjiT8oAabqP9jPtU0ay/Wd5er4SL
ZJPuy8Mq12Y9xoF4kevjD9L9aahkaIWPd7dnghchqZr1vKFfYmDfM2rMhzobiGZOm1ZALvUxZuuU
PRhRTqjVJ/is5+ZbiP+st9PRsOJW0ozIc3EJsjSIjox5sWjd8M243B762NUluKIdixtXHsVn1t+Q
NNDrEWiSt4lGUkCoMajQByOt9j46q4ZE9g6QzGGdZkcCjTCvvjXSwP9Jql7yxRzIzgNn+m1otUwZ
nlwPRuVFt3e1dgAs3chzeSzDL3gvjZHpmd3GQggyINGzcRUNjEx6VGzgk9j3z8JaVg6y+HP7lAm/
PPwmQouZZTVK9Dotp1ADl7pgpPA7Hh66ykyoG3q10xZdpPW4oxD5XAZ8fO9Kyg1C5Eo6bYUgGar2
0NpjTj1jJkNaxbEKWNTQKI6Z0iDdKadDJr9xAe7/lSCGnrLNMWebKRON7Dzffg79Va2XI384gIxg
zf9uPg3U2Q7m+zVDyb7qzQB3/O6LLpp1uyz8vxksmuhDbUzMQAW7xrAR4u+V3r9eR86lMAgkd4Ye
w/G8aslFQ/x/5T2qoxXTet+H8hxGpI4FgUuRfI37BRV3tFGJxaemMMXM+EQp8YylYNhBzqqa4jCh
I+cLb+LCSC74dpherEgQ0QqhGy0+9HPZ8BrzY3dFxiK+ZWLOhlqr81fco05XsaHm40BVYXbcsXPH
ES+qg6c4BMwT3crDe+S/W9VHpL+GTxbiwCXPzsu3ebkpFCPmpueB7XOgiB7pjZltj7BsQdHR8QDI
lABL1sWldeo7DGLTjy+7Dus3xEKiOB6ovtkZA+U4vUYzgY2Iskeac9J33B90b5PHCwoXJ32aGwSQ
Xgipa/28Hf7bL3qWX1zGN5eglb3U1UhlUFhs30q+CGWarVxQ44h0aRfMvfrPJPSi3L/3D9rr2/wo
cIoEghBjWSVdeWvgedSYRq5/c1H4n8beBFGsZ/gtNzyb2dvZ73nWEENUMYUTxl7kEFFWsfQBDp6a
EMvwaYXpPxE9hdNM9XLLhHkIudA2N9fD4XXOVFkQEJN7GPTarc0pM0UXrkYaDrcK/PjKwc9ln2co
6Uo+3yLntKyLRDYXtmZTuP3o57eTk14Llqvg8lTcRwBKUqbsvFFRJz/DhNwC8HsobSFtK4lTkrUq
e0/xyJkl5M7TktPt1BSHnfpnRTy3D7TsUKtPfik6cY+p5CD7sB19lYa+EbQfMtCK1zBsIxSKJQ6h
qhBMgIC8KaX1Ffkv/l42TxhRVRt558yRGZRaJ2tgFOYYvnQ8J0hR7Uy0yMA5ifItBGyCdYNWiJjw
btfZ9wRgd8bs1Gy7yNbUrcI4jM8TJCSfLDNw0c7SJSGOjmQZ2GyH1NV20mHW4Ihydx8oTWEXDYTg
sXqBuqN3j3Wyi9jrCEkrvGTharINYkMuKISxmPHHIiEK25TAhzgGdqfBTJ23xXishRH7cdxAQTME
a5oE/yUHfhqjytgJDhCJM3f3M01/rkxMYzUyK1NZSJpqep7h2FCUmYsAGYDAVT/m3cG5yu6Oku2F
Zbaa7boWm3eOXD01EBRhvHtsZ18K9XpTAD6lJyGj98McubeyLuXcMtvlHJCMSDvktN+2zbVdRvg8
u1AoQYbfnVsAXOMcIg/7JOM0E9lRjloIDIMnjmm0EH47396TR11NkbQCw+VfcnvNmmA9zTMwISgu
AQHROkBr7pFxLzg7sT4P92pF7El4MW48gaBgs/VRkqjIy61nW++1AcWoZCKRjRloolUkOBHMVpqM
SvV4NG9yAPSYJC3P/chKGOXrvwA9B21i+w+/1SM0txeUO0Nvjv76/+nOb7tvNfHnSSLDwfvjPHJn
1+23LI4g2GBiqyFh9vxKIWz8Ynue3rdWay9X6ms0lxNMMtG8bSZRo9UgqfIjsLvotnDrvODni/sz
qwwFVQd0LXC3L6I/znT+YU1yGEWe4EThbe9EYN0bRw7qhzbs8NhxZe20ZGnKfYU+XrYkbvwpsbcd
sqb+WWe3fCT8WKbJtvV7rAats7qjhHG1deE9ds/Gr9x1FXkSX+GMzZ/ExLt738KK2bPT4AV3zGcV
TGCcp5vP2OgF7H+r1x21n1vq+6FNzXbdflRsVue4FGCAf2gsZg3I8gd/eDxyJ35m1Ab5NSpkfcH0
DtiYC51VDGZHciVmI9rNXEF0KmN+1wYiB2A1xuRWsfQEZEmye3DufTasyhvOBKDtra0PVQpxhlTV
FtfgBoqkgp53GAqeGsxTpYO59Lt4Wq1G/0Qdeplr4XnSEg0GdAi5TFRarVYsI6AxNs33QORFIwqf
9JMT1cb7WD3meZNsabOs2jGrUIoJVowhnjIUiYFitol18rxB3I0K03Onm7xmZQyP9z6Vw0bwRblh
M4LCKKQOq43OMxxgW/XRBD7l6kCm0w+ypYO0R5srU5Icy7yY2RzzGKiPZcRBlKNwODT5E6d4AbtR
sDinNmOWDxzv4tkNhI65RlF9mGN5fwfg3vRk68d+QAUyhZMgrjI6g7yDUMkPtH8gGpL/X+spLlWP
Tznktfuh8UBhZCo5GYGM/ATkSvOb0djyQ/3Y0EZVrmlamy69305PUGK5l3sOn0mk/CztxBVdq5iO
xOgTN3K8DsL6B72Kz0GwDpTvHvEAhf2tUt1NR2AJTwY6SuvfN1gkN2GVaaLf1IyGD8RWPggBlcpa
0PifYkOEPJsAKFvEn8nQv1S9CUUmaW2tB0hjWIv0RbVqyy1Bz2z4p0iAXEnvJbtVIL4+QEV3kcNg
R1ZyL0ekwc3TsJEzUaoo8FIb97VSEJdnwFgfcNfTQy14jwEOqNmCfcqmWwpmzRl8xf/wRKQoFPIB
g0pULBZsQ75hZt1LIPsIFaUtHRwWHWjR9kbeYop2TfRZG3zcO4MG6wzNgK8XcZQSKqtzdoZJPXkq
l5Fa4+o1jjgBUhEFOa6e3pqxmxjFSPEsS15mVuV8xqZmA5TmUSD404jG6SgorCIKuxDav5Rdi21B
BOeL1ZuXBb6y32jBN29b1wQ6ljqkr01hF00VMZW7B0wlZOqJt3DJ/UzIb2oG8jnG2CCB1fvGcY55
sCRe6/2MbSS+wak09bc7buX7B0tpYc3EBQ+2Le3c0kwK6roDSeEq5ZK3ZJ3rOvvdqIRBU7CBPVzF
Wvts9K/iXTqjEwJpwFI5PTgXjH3u1jOmC21gMGuEEo/IwPjY/cRXAaHQ5yJzS37aXSLKKPaHx+C8
volDRtGKYYEoNVIj2Nvaw035Acfda62loF6E9Sah2eFdBrHyIXfDqO7kXRp0Af8mJ1hP2e+Sq4t2
DENbqE5NLOc/QuY3oeR5JzEj+m/alN/AaAZTS+B1M+fyG77IhdnQNeGfwASZase6wOkfbEupsNnZ
aNGMJuazumojAZV9TKBXPGAs5R+HjDu2WJouIBvf4s8EIXSx4pelPE7A6e/l8iVd9iwTczG6iMb1
Vz/oFJhzgFUxtZh1jcf4/qQEmLxIWSiSrevmpv7DLI/N0PJ4ZOhZGEo4u0+uafQElV6Yva2IPGDj
az0qHkfiqhdL8d053lFcY6GTWLE+/XuveV7tKWb9KEPfq008dERW17UxtceyS2QNeuDokaEdiBuc
e58uCGkfvp8S4okxvXUPqhNXXq2P7qHnO9IMW7+pY8uTtohn4J3ui+44CF/Z6OWdV2+cMawFISw8
0MGwsnSUxn4CBL946OitDQd3JGHITVpOPi2nrlHrwSfhjnqnlmEGmoVoFtMJjd3kbdKgUD9cSsp5
y+1x4uhkR9XJDXnlbPR87vrQwhkHdeJaqh1eE7KINs8g6VFT0/Few/Zh45J8qPOOwtGMGXcGjFo0
JCifOWcnrcHYETuaikxLuWjuo0roEyTgTdgeUsuAZXS+iWxtUT+7NCX9xNm4T50t/gv2biBe9Z7F
ncmryZCj/EESMgesyW1drwtT+sccJr2rvrr7mwcKGfb38e3SUFSrw6mcYQ4dsxfFd7dTf0FDppA8
TT44o8Ove1bF6NFnMfut+xBc9oEeMu+s5Ft5PMRb4IXg/+vZIq4z+tE3q+/S31MAgok25IdDRiYy
pSHtbgkPqbXsxSMAhqy0CUhzxrhny9iVujYgvlam99laiY2VUX/3FnKw8Q/gA4K137XTyOqa2SCm
DDf4/e2M9O87NxgddMVeNlv0mrL9sZC3A1f9HJ6MQpGkEd/D0b6+FoXECbaMlfNH/3IAtPs54c6U
G6vXF29DHQadacZHizcTWFuy960yA0oNxQ0UftAoPTzrQibBjbGrYIuC14jL1U+83Nt1kCCqeH+W
VeD+F/fWFeY9C5jkXNaT+tofvATO8XWNudcENkXIApYNp0K1eTBTECH05dAA/FrQx+I2fcPfySlD
44Nqaatg83y76Jop2LyRKI9kDQwfoCzppR6h9ziwI+ywa5Ii33myU2nHRKji0mFeo6inMUturThH
6tbFsqqFzXXtB5O1G+NpdNt7ZJupFN2H8w3s6n7300W7HsrspFfTwHa1AWQo8mqW271R8jE0FaYN
JosmpwX3l3z/4Vrz02Oju97IwrcCGDhKFGnX5RRkbe/w53SRlKigdMORt50VNJb9HrEQZbE3g/B7
7HlGb4cZxyw1YJqdNR295GAs5pG68A50rLHbARZDEuW3Sju1LmdafQop8c7b2P7l9Hy7xDT99BPc
XpNKLxSm+zyy+BiPq7XiweYkvSnokYCRe4UnGzXpOTn9XY6gCK4ZyVsnWZgOPfUcZZn09K2p3RTz
YigrAihT2g1Zd0hIjF/k8QESO420pHm4mQnAEij19UIr7ODJuw8up4/1WJ1MjeaJ53lHMmnrFVGM
YeGbl13uE2PuLU6xBnYpkm7lkDrViE1cA9Ikd7/A7bwWCXHydbyaci1T2/GiJQm5Od7tyWfbU7PB
q33kNfltBImnO69WoFIdOFbwmymagCf+zy3IHG9bPaeaaxK9bivwnU/bErDn0U8IWYPiribqrlWv
Tq/5OMViYiOia0c3Zo6FmDUrfhB0LKmKu266tcByIGS5K/1phmvUzabF7K+461YmhdEhaXOIkEzf
tWxotkjrGQTLnV+MPx3UpiW0hsrMt9Cd7N00KTwPpFEQM1T8TwaNLnTMhMq47pGNrq63Op6J7Xac
iYUeFZTHMqdd2xO5la9ujhnRqtI/ePOo7qYQ8TPwK/n5Eho7ONSqQOCe8/H1Gx+o+ntvn0M72gLK
4UTb+q4jg39rOzGxDgCRjIAYUylSzQ0viE8/CNw/zi81TFfYtMtyraOoO9a8Fo4E9cuYHpUmLauf
HqtTjwxQiW9AmII57N7TWj72mcgMswatd6seFhjw4B/fjICScXDqX+S//7YNZ5RIBdP2qKK16c6+
0QcFQW1Cgo+CuxLbOGnLGjCjjv79YlzeJHjPH4rKxSVQKbsNzgsLP4qdLNCGKV922MGDFR7C7ngC
U31X+Ew09b9u87/2duYzW43fa1kjqYcLvZ1TDNt6Z4u3UpWV7TOo1hujbmjw8s8bDT4dzfoYGzxu
q4NTlWpoMXD6R/f4I0wzyh9exJvovjiUXHmP182nVAeTzDx7PKJ1sb+1US9mCA2ehMzSOVat5P69
4X8YseqQrKaEz2JBh6D6p55UtB716jjIqlhXsqnxLg0V7/gcWTlK7WVvJHvMx3VQDL2Ky/pp67+H
NE1cCBH8AAXjekcHV4Wgq/F8gVQRClJJFQzmfEz+JAxL1DXHWoG7wg1lhlxHnoNyZzIezduczQoh
ADIHviE3G4lyQc05JohUPyvaTHQKinBn2y1/wM9gxAdZuHZ92ZqIjIio/h1UPfDkWaZdaP8n0PuE
+ox9DuuYlyh9WIqRrHaoxashavi204W25B4NErt9Nftm08/sX3PpjG1UYaD2Y9n34j2h9a+1TCc8
y/rMb1F/dZzPwWyuFLJ3c56i0tLEbCjgK66NThaqZOA4w/ckTVM2354sS6ms/idKB40dWbcFYq5f
7Yl1C9NT8rKsUqVWionc4LX4ys/OJ1Ypu/d9jTp3pPn28ZHuNakgXlp2PLVzfQxCkkaeDvWyvx00
uiMEpHcCgexSEnNtadwH7GfyaX8g4uVvJnZD5tn3kWIs+/K/QDBAxtjyUfmEv8WBvsPGQyGZhQxn
EKwJs9Qgga4nK6AatD5G4q40wJtSZrTP/zRwOu+SPjemkfgIpWvG6/cVViv8v1hmoBiMYZiEEFUi
CW5ZWTcGFZUvyYw7ah/a/1veKfWVZ+OHntoV8mabRB5TrmiipQcGywieRiEDgGz5eywjeIkzzze+
U47ajt6O5Ze99ExAVuVSM7POupC9QPpxNE8TPBCTs8y0PEqQoVcpXryJzHC1ThnlmqX6cN85Jmw7
FiJgejhfHigTzngjo0lNbFWGX/4uSamfeVnRZ2/qZzsOTcvS5k8oAKaRRFaxnVqHRZg6oVaPGC9w
jEiDkTAULJU9wlw94OGxbjHeL6EMq+08n5kmMOVWR3ndK0VftElSsZvs6dohb6ARFqEnGfxXc/tg
e4LnLsZlr7gdVcOYTDHzL+g03vFRyz2zQyoSWveZC0jGMpMpylyYbdChugHquZB6/04Uw3GKn11w
xOOJXudzt7mX5PrMvrZT5Ox/CU3TZwWGpNR78c/Dwn5ilMsuCJW3mqimNv/8XQdWjA/xqUZUx1Pw
D6dOOz/RiAlWnHuAZdcJ1MuOzEzK8NjCU1k1o7Z1nrKcWTNAMngDvX47NaY6tA0XTztpFn0Ke5sn
AoeworVUXIK0L3j+7eeoY/si+5OSYY2sXbe7JAEedr3jBblGzoq/C1IGWAfBvys8zuBWzhIHulub
2M+CJF+hCBsrss0tGrL0B2RUV6C8vX9H7sErh9d3xkKfpcS/aq2j5kqZOyozT9BgnvL0FZQ6Y/6K
FRYJwQMOdqERggIQjCrkjibQoMz8DG+SycmEiEmTBI5TresumwnoVdVZdJDD6oB21e001c6CgD6F
UXLWct13bhZZneedyq7NvjNHKzPkJGh3oa/YycEqKDlbDYBTdKZFlXtbUJA+pupTsh7W+v41GM4T
J3P5OqJJxdyzgGP6h0nrd3DZ+NF94DQKNya/tLEM/u7yh1rFUICThtcBzzqX13FJSzblQS6qinhP
TR84/NWdbcw28OuBq+BSOPgxQKqj8tK2+Iu15CXfy2Gpj0cBXbfiUYz+bacl3dKGjtLnr8cvOhzg
ts05rv4U61tYRAvND6oVWp3/kzjRODINaLqM6WsBQybxMNTp8gtBuFygym5+QUOlPb0FRYGtMbQm
B0hhjZsnqsJkJ6lgQVgLGlC6NYt/C6lRLgcRuVcz0URmFrcJEXIQ1nQhSehLi37x7nr0ChCYFhkv
fb1orizH7ywU9dE20ZmMvmDJLgZeQ8EbPz6rJhTJbMKMJDrFycwenRjaxh34l2bfXbREsP4RVAr5
XRbbUZMzeVuojgf37xfuu+lii2WC1rS4QYYsBDi5soK550dA1PU1py1lfrIxWRqzXOXLPge79X0Q
LTk+kqtQ+hv3VyxZxQD3L/2iS2HvfWBXxZTei9YDUQ3LMDcSZNTlB8stP1L420wwrGLKFlE70ACP
B3KZoNJN7Y0DLS6DAgmfF+WoplcoZHWqvG29A7STsEetHZ75YIAXSVQZKFqOe2euz8AZ4LI+zmq1
i64tOBCovJf5tfAM3lsKrAtvFxSTMarOYdtCDrhGQb8OfRdS9InabcXVdYphlXKITOfdgbPxI1hu
uJRZPXu3x8mznaTWG9m99NlFKaZMeF98mNU/E2XNRl/+7wQ4OxiXB0Ev4WpIgi3hnXJ6udrh51JG
4etI6UCg8OwLq3V5jKpoVkbcqNXfhY5BNk8itkkZXs0GQMqPuXM8NLAw2KmmCPm1cGiVOQj4x99u
SjFD2YLEv9NxantxhXU75JimLUN+aGA5+QYsXraagNQkA3ZQ7bVkOqQQKs743jZEVn5BYF/XavXT
shn7H3TmxjzvKPf/LY6mtwmhS11/r5Mg4hjCf+s1/Q2kuZhztLwhXNnaS1ExD0WTbRZ5N8a9+mGj
68gqRqOgHWx93dr/hlh47STjoIR1leOKr9yJEc80OAhz75jVEwIFTvgiwHWhiF4mG2a7yzwcc+A5
ahvDHlSsXTNzDcxebtxVJ+78cGpTtwJ7zHdkhwVsAi5oo09DGJWs5b7WYU0dP4kpHeuCLmUCq3XX
O9rHW6/EE9c+JqspT8oZ4B9uch8/MPUcN8Yg22Ley0YP9WTfQG5vZ06iJ8dpet584Eull/mRl37k
JNa5bz/1twvvpN7xSJ9edl/DfzPw30liDyus5crp+tPuBV5xuFTviJQBlLYz8xnMHgCpG+OMzpG3
d2YboLGSBH9kp0yw0uNrzOJjzGy2w7ak6aJ31KI4xOo7ZkjELiW6lMV5uvvYhnUSdxrNQObfG7lG
YAlfoZCEnMXh5yJP+DS5UsnrMtt144BDaJpfJ/DxDKNKowKHtLjtmVpRreyfMAx4TgAKW38DjVku
tH8Z5UPmvTR2C8Fz5PMnPx3nV34AGsAilZCiIM3n4Ufn9iTgl+ZKkOdQpDpAWfJBIVrrdYRju6Ld
C1V/L7HVOtfVt0xSbJvtoQkDpCY0+azYaZbVCKQk5JISC7VLX73IC7wYgngWuoZ71BMrY0rMTu1T
rrmmzGaDGd8+QE+vx4aYLrLUWoCuU76PBitHFo8SgY3toAq01s4lhBn4ZibHoAc3pSVTs2DUSHcx
730SVZPtgYxCtV+hFMnV2H7tHNmOki+9FZyHkEjsiGWrDkZxHKktF8yBSFM27hETge1T1aD0C5Y4
G0HlT78lCm8FMQc3117maDa/ivltag9z3nLG8AsvqBZb5A1S/sP+d9Zs0b17tnk7HudX166uqjUx
whDfr8tzUkltrdB2pdNttTr8k+NmcKGvI8ar1sj3CfSh8VihWzXj1/LQ0UTykVsZWFqQFOsyXCZP
ySoPZsJ2TXXvrbQOqDYmKMGmmccBHR1V7XdL7hxcEXREzH5vbLXFjksF6fVZVUnYGxiKuB629C7r
dmwyobBPesvzQah5j2kCgPJZWH56jZ/GuAuodVi3n/sDSiDXEu2iD8ux9Q265ZAjN2ehCLw6YdpO
ANqk6iC0Lx+D7lVd5gDcYMPpXTh2hxywbOnuVOrp178u54sNFH6s6N6omhmDTR6TgTxUar8Ud5j+
Sqkrh9PV2X782kYvC8tDIOuymAVBXrKbpy5hxvJUy1ZkHACz7Ib3A6aP9s2HiWmvVOF5tHJasf0L
jV0O7lxJvO7KKPTEDrwkfmfc3gJI6o8LL5i1wNmMwY8oBsvyVYeKdkAWi0v7tZx+pgXY5tAlI4+/
7dH2z3rgLXrpfvC5LyX6i3MA86+1A/9sHAbYmWbKZD6ilMbaZl7VE8s39JvLDLJTw+CWoebyRJoc
59ZMp7v7pxep7UQpimV7TTL44flSMWV3ikfoBp0i9g2aio9WohM1bWK5S9tNeVRBbhTgdWslSnJQ
EfEW92ZlXMpkPMOoQ66Eg6pUePEIqEB3ek1FsbvRwDpEbXKnJTSmCmBP+pCIwF/bEgLCSPUOAWIt
kF21IqIhLJ4olhy2VMk7UAOQwWbun60qqMhv0xZfoN+pK52bUi694lQGqnrTpNdcPytJk9ZMu3eO
Dvnv0imlZxU9k2bbZhxZo+p7g4nx6EgvAV0SHMv4fjaIjewbOy0qpXwsH0GUYzzQ+DH347A4Fo8o
cIpGLgwiU+5Ru7OSbIgNz4u5gmeP3mCieOzcLICMmr9ubTPil7zk4d4lDzgm6hU8L1fq/xONIBvP
PmT0OaxxkRE8xPOvyeEwxAH+EdenjlZ8hqzjf3wBNP12LapPn6jUpW5U+mewzd1oxKuBKup9EZQJ
U/pAVJJwAvvvTDH1TfCrmo8g37dmsLvrt/FKrPSH6hGCTBLOl2RNlsJrCjxNHSL0zknHi6ZRcw6T
aGFPMTDdQU7g9BJOgQ+5BpYp/hsteV4TPfXkgSKor4tZDqZvOtcK3Ul8d2QAHCW/spDjmpT616wq
i2pOTGkDJ8cEBqlzcjrnUVCyFdZ+qzPFXRKy10My2SKPOoQC47O60ewcML9BZdF3wfGSg/1c4oan
DhDbtcdVQh0GlazrgshQTFr2bHxaXsPUYbOgGg3l3+jeO37gyFsMppMNomTP9/RFLE6GD3O/H5Zk
v/2DH0aFv3EK00CWT3z2/6mI9i3QRxOWYphMDuMkrM2tsfwPn3ZtWHCW/DHKEogmK9KcOFtImMzD
oOovckRqftt9wfra8t1Act9bV7NHZf20Hm5yQ+oHHa+fzvHXuXJtSv+PJzJzunjF/n7pYClOPgZk
7wfnFobJTx5MhcxAN7lYWXuFQMQ4QPTdWR1RDGNBD85USZibnEXWc4rSbA1BACFGKU1DsN2mWKES
5eXTL8x9nc4/QwiIAV4KPu2f2b/swPhOal/li/cYW0X58iVysWTMBD6BfrsnEk+GxXjio07yT+6Z
XCIDqAnt3x6JVcBr4tmhtuLJNhGCHyfzIJi3E9/KddYjeKY5hjPx3GbxNRdrBd6gsxdgppsqlAPu
mlooQyzSsX22hbJVWI4alwxTk230qf0UhYfH+0V9lAbd4aznXh9gym77BhJFw8nJpaMN/fM9ticT
NcmQ1NQ1QunXtUvlvZg/0yE7dWxJ6GaSjpzfzzz2CTE3b2omNMB8RKd5nbudcpIgPBGRYZ8MM8F6
LXvVL6CRS/vShIqJmDifvGOMG9aSxelGxI8VVsqTm73aM56UiFSGY9f4EcBM8OKr6oy9BIoJubCI
1p13fyaMLhu32t19qK0BGmn564hVQaja5QD37A+bWZ5bMDk9Obt3b6wCFqqtzh5SUSLJank4otjg
nB2wDuiAQJzm9gXnOB2zRAFICG/11vYLtmwGOsQzbXFDUiP6caSl3SJBb5a2ha4Hqw4qVjSmy7CJ
XxGX5Edc1faZqxypsBr4EbLE5IvUz4dqz5dq8OecKzuS6Skl4cb5R/DPeJIevrDoZgLWktMlrdNS
NJ5FBrLnI2z5vsnjlUdXXUYP4UEARnOLfWQ+PYubJJTf4Jfq/kfi8j8VYEHfOslx2dPaMsfW8PhC
MHReAPyRNvyQPDpmoVKBtQuJLSPXzOK4wip2yjI5rJNV6fcBfI4iRxefjyQTJWfENsTXY7UvIFwR
AXUPuYLSRgMuD2qCo6/a+wmOj08EnE9VArqc1cIXnS4ArhZqxhXBMeePvHx0h+YrtpSDmjj4MyKJ
+HBUWUkEsO3oDo4/xSc5op9fibEsXA+pb69fLaQmHW7SG8GrXi6DIvfi9WflWVIacpF6CXeLwUuM
MN7n/8Brq41963iunWgGABw2GyimwzvQ/VgGDZgmQ+JerjOOtfVSe/3Ds0vFG7e+9nkbW8LdAOwt
qeamuH8fqF2gjtU8tG4jvX9iS/qO0meHiovKoaAf+oido/GRIeZ0fNq1T38WDHfgIjVumY8aJoLY
sjlYuqSr6Fbh63POAtBBtFyNUGPoHLGR/+n/VE+GGfxgtygBLovwCGaY6jmYPVrEOP9CxMzN+5ku
gNxKm7eM8Xg2xqPWj9tf5DVf+MeCK3SCgWJ6wLsfFNovIYDcXF48W/KXcFa9dSatYp6m1zogn7k7
nOGlwRZimd6tlH5HtGk3JSozDSFvjwclxvrEr5R1h8+wQulNiq17O9ha0b76fchbRXHyqEPvyj+l
qHjkUtBiGgf7c4aAKQNo70R+rYA6zEzgeXg4jXtgDoBQG5Mzu7oudgU89xiE17jXwmcD5TOLkVm2
0ATxtT6dTcXUZVfPVDJ7z0SBRP0sFBP7VLIwoOpLv0hJ63GR02tpXhL6ET947B0mdK0dBQgCx9U+
adAC5W4/oUppOBD10mCP2UW07am6hYTXHqnKLtSPmLfw74rwCFy8CokvYrMkIz4unpgtzV1LsFoI
T4NZPNWhwa7ywf+CtJoZMdSaoWaa0bvKCP+UQie+QnaLBUjBppDEhbneu6QA+UNpfwYblTzq9p6e
6LJpfQ0R19gZ7rHXmHA0EPLNB5j/VuOd+rVEb0HX4wQ9n+euciQoycM1R9kOAZFSHf+gQOVeFCyf
VbRlfoMB+J+NcY++/sZWOycNxcS+D3JVbzy94tYwUrtxTwv3NJ8xt3yp2x/h/4tPyMADrZfRPcPk
Un+RH4TAd8BcyLkPho+mHoDmQFZUFXMeMNUah3F9g81EBtbMM3DArMft8EV62SkK8NtrbsRDm2OR
biHq95336qvFsXSiOCYam3giBFdugzT014Ia3hdII29NDyQfMakKZss0spIPaCKPVb2w9SafLCim
JKfpFCKkT4UgeAlyUqO/j0zpgc+LWUo6zjq0XIN8KFsccFyTpP7MwZaUwNsj49n87iIOKIS6qtIp
z7O01m8eWssxYo5iS3/0pU20GJRnumv3exvsSovMYDmQWXMbxA2weJbOxBr7f91jdR/xHUZ6Q312
ySWUfrOvBtk+ExBXsYHlBwSCJRawoKoxvmI6pyTEUL/SIA39J3b+be/yO71GCsLmfe8W7dqdw3XC
kXyTc9TxJuwOKLYfIthl03CrfxXnA5olt5Np9Aj5+M9xEzyCizmQuPOO4mqgpYq2ElQrCsDEhSSZ
uJ2IU8UeCaDHGhHLAWqap4Pgs4oo3bAPY8UL16ODcx64Ud9d1hi0f2+aR9xd0xMW8J5r8mcwwZGx
M2/YnMHa12C40R9J1TT32hDmfA0BG6FqaVQ7DyyHAbsNzkbKYGKDn9CI6+qQ9eY3Mi+FhDou17Ea
aBysO9SGt9GP0Sz8W/t8ILCiEIH+7AkFbBfXS0jQEoPwyEkHLUf/C4scoivrsC/TtRNbf6YuqT4t
fFxUeobH5phGzyv1qSnFjgWtXuh/LappoQpugF0L3vK/IOjY+Ez3rpk6odksa2cz2QJienrSvMs1
4cPeyb0b7GC1cy2pqzbPK+3vSohWOnvfekoN8qJkVMLhj+faSS4+gy+a/Vk2EOkXtcKA8AU84Eh8
8uri3U0aPpv4rnduhQmDvlqTLFeqwWMQ+ndrEzvtvedikrRY3oerE+rbwuvXvjpmUP+DsukZT7a6
vRbY9kRwnn1iGMg7yqWLHEaAKje0HRIpOfK6Se4twSr0TP5332/642/wlVbHP+WrkbOSUtgjxfNp
nXl56fQm0r/k/ocXOSF5UkzZvYPI9ZgD2EdfE7ZRRvRwaWaPHz2P3B+xcRvJpjWBbzeln6LksBeR
gwwR73RfQgR+DkCiKRUrSUVgEZ8IQR/2lk63+hyG21BYU/M1bNqbSbe4Sun2GTbA6OkGc/bgcnto
0bOEwBzR/GNInoTHUHSqDLkDTu5wKKvXc4TVMm4RhHjBiwOFlv50HX0+j8WOxe6d3SfO7kuF6Wek
Ez7OTJl63oBXqBgFCeL3lfbE3xCz3gHa8Jsw43xsOuBU3j30arqg29NhCkCJ80XgUBQa5ZGML5Gx
TcNQUvQM0LZv/yhTGG9ZaPmTjHrwOPH1JhJ4DVqFdP9g1RCSGZv/rKsqaKauHQlmZoMijVsAOUzu
+CN6rsvE/X5powGpRYJ3bWYBawdQkR698cAJsZLHZv+GaQTVqGe0dKSqDBBXm53JzFxjbngB0N3O
MoJ7A+pXuw+IL82iF5Fh4DK34OhuHlTHr7BLk7KuN9gdpWli6KObbbPYjSDtiBufUJN5rWRBFjPP
Va+bu1IjexbyKh9I2mXCwN1yOBKzLiYT+rDwnw31hnxmYyO3s0XmnWywoaOqHa/2Tb5YYByux+53
4NDsvmpxCU5Dpw+8ztQE5ntr6tvqDWNkEG9Zy1+jPGMwS4jHJ/it4i3mAcryjHajDUwHXRgTDWlg
OYjcKwuozwhgSVstnd7G7jnU1wKfvC+R3r/WaGkcqFd/F2F2Klm6A3mIHKpt73l+IoHSW3dMpd2f
hicZKTt2r2KJqsqndVRsVMwivqvxPcJxgH4IINTyA0E2X4VF1YT9Gmoiazp4mEmKZCpnHoeLk9iS
p4oWE8J/Ecj7cD5yUJ8H4eKwJ9C0Nac62h4iGaKyRIeOF9gHMHhBoY6PZK/wLv0yfngvcaQgk6qJ
XKR7tOlcSZOGvh7LRXsvQA/0D/XLGVLusvuBq/vVy6NIJ6WCPJaIX+NECIgaPFs4VRxQ2CuWqAsl
HJ8x2xkT0CKLwc2U+sE/tgTzVr+30n+k7xkUBsUg2yIdcro3CD9noEJA8DXzNVF8wPJ7XwiJYiDh
B8JVFCE5VyVf7wau/k+mpTZ2KhMklrHPtWV3JXTVbGUJx9duyk36+uzrxDx40V6X1AXQSHeXpEmQ
0mHzQ60YOUqUGeHSmERj7D6WT8mg3Q0ORXLIJqnTQ9ThpccBGxS9E40xrJSZwXmZeA76XJ7zdeM8
xQcHSKk6IhnMjt6Ukz8WnSgv1/AM0iUeWarzHzZr6bvbXpn73BndLexI+PPG+8ObQDLef8D2zKjF
rrPq3xLfhtVWBaxxizPwqGbtvAbYaVJWoqOODfVETN7PKGc6kn/G8q+riSmYU3mhgglwqdYZIH1G
bJiNr/VXQh18xtkW5JR2q46ODtsQ5VFj1DAM8prMdMWsTEFaYvvP9RvRrqYrRZPqNQ+DC+FdevI+
mndVAJvQ83+enmv2syVYKJkTNMkFX3ANpu/ks3w6GOYogkugFZKSckzgNV7SgjNsPvCtdJtVmyHn
KV+lZwXRryskHkmIG+H1QTK9HxRU7rBcuFGRrz0yPXrY2N+iLZAhJsLsAZLqdZqL0bkLKo672Cr8
srrjiAfHooWLsXoiZbLmRtbzXO+UhoYKSarEtEynxiXe1ceN3rQhKlCWnhWcfyqcWLZwoXv2T/3Z
FtLyfT/Xo7zDf5tMYnl4XfTtTNXfYl96UrZ/T6/FRLe2MR1TUc2tEHdkxS8dJ+oKzWO85gAOZGS9
jDK9u1v9+NQU6/7yVj7TdZYk5edg2gbQNPrXD4IG5muN7HuaLzOV6wmBHJI58LimmuJ8ICMLI4tQ
edWpdNCRjKLMU8ZBPH6nAAC0iwA62muT+Xrf0Ypp+brOee5k9Jya94EHFaTmU5uwKNPfuBjkO/MQ
kRWEuQH4QI96ozXfEhwviYyiBHPhlWtHL7/hVfAO1kLBOepJlC77DEUwL0EilDCWowijuPKqsIY/
EFiHgoNs7miqQr1RtskZbHuFdXrlaJj+Bmg6gTF2cjeUhpje53gEqT5THLUtFJjr05cluk7QWknk
YUy3HeE0pBuOgvZY7d+gSzTWKtr8G5K4sBkEmtzwmlNDWpaxRMLtqWLHirvbt4cKhYetlEtzBAiS
lyKkNetQakBd141LoPm4Pj4KTmNFZK44XZXY7n6GJzOS9VQBmkO28gDSV46L3I3JhBbKSz5mAENE
58hiGpDQv9RakQj6V1zIbTqDPkqTeaWW1F94ZSGJHw9pRRoMgXolhJGfN5DS2MLZ0KpWmPRtAt1n
TKQp5Y59U/BwFH+lKSo6rW3aBO0jZ7qbHozkbXKJnRlY4wZ39FhVa7HqShX+7XMag6TvawVm8eMn
WEp1j1qniH0fiSXws7+hWR6Hq6gpbAsdlBTbqXxaHgVFCGXlwOPngipYnmJGSl65xoacOVMo5pXz
2Bz+tbP5Snmoge4pVVGX2vMZTyRadagwT04MaBlkbd7+RO4mdNdabxZTOWtnSwQh2RjkLghoRRie
kc60a4fEm1kVZ5medJ9H1HZLz9orLwjyWDhZpSQ+7aj+pLQnaOSHnRFQi0q8FvoR7sxTd2lsuVHH
XAE2rjWsT65BJOOYn9CJUhzf3TiSuE7OQ9uPifUI1xA61F0fRbQMExRTn2bYBGs0a3uL8vqxx9iH
wdwBtiO0GkQZGXBpZh4v08vTsRcZZl5cC37puh7ws7uZHh5oFA4x8lxH1FkP7HNlDoHYC16klYbU
S7QJJ1ZiJPI+M0j4U9/WUDp1o2jETWsoNTJojB6amAl1Bh0KHq8usXlVQG4AXcwyDXqZB0bN/0o9
D0T5PkT132EsEI9cddwhLwKjMjJGQKDfgwws2Do3YKvUpt14V4w6+xtt+RtybKH3USyPLFVCwkfs
EXXoe6BZRuMoQyc4kAZGMJ9mT5Jzz4nJGxSmPEV1GO7SQ6jZpgVV6QSH3tOY6/40ZVYWKM1h1JUa
B7bV1NchpJU4UPug7LagKEF4DffkxIA50otvZjiwWklr+MBxey4jW73amfHR56cHMQQw2wIPqUvT
bTZCNNtx98cqveph/RFeDed+ymfEiXyDsEMN1weLoA3dc3mOwYbzNEDs+fosgdybIacga7jFO8VR
Mnx5IOUsS3h6aUacrtotZqYEsjxoG9T1pr92EYTlNf0ypcwCtzYqpixb+vOmUdJM95r0sMINiLDJ
w+mavzRE8k2GKJYHHnG44Knw0T97pttncM1ghF5kq5+ywFBwBJ1obsu1lTsT2sHH358jPpqm6FUV
e5HZa9F6tA/7h+aLJdqPq+LuNaNDL8YcApJh6OZLIik8pxyVF/rv4Uzks87hshta13rstKAZuJTG
6Pv40lDpjXNCQRB9H56VnEzbCvTvJNcdOYKJ4eG55isCEuBBTbfpaGS+nV/osdJ8q4sOo5T9sMX+
H2aryXuFfWMHGCgx0/u9w6dDdiobJl/B0Vzu4byUxWXtGfaCtJxqTj9l7hTU/icPtImulucargFo
WwT1dddRoIsC/qU7z9aQXaW5rNvY+18Cv2KU0jzF29/8qBnRcVcvhjMG6lCchmJQHNZdWZEeO5Vr
IQtNiFH+oV3i43N8F4zwZV3mp0+xK8ALpPesOqTYjJZMndBdXS3d/SxzVt9bmuImhJECMSwOyFPE
EST5v+RWC6u0KWbk60xE2ueZobwDiqc/DsPpL9l0AZ6Zmeeo2TxN0TxVOsIj/DFzHDFlSDuA8zwU
Rr45TEVmJFcz9G6QKypWtwpEK5KfHyiTZvQvQFgV8qhmjIA0lyoZmDKgvtjveUcKOaNJRqWoUpis
39jxfXZVkuZr/TJnoPwrg4KLg9PSEvtZvrR2YnJyshCQybmqbTiun3z6tyr3PG9VLlp5BnVS72eE
k08Ti1RpxM/a10L9dIMMSe8UWS1gaHAaiBGR3HcXpZATHVylMkofVxk6xuFvtLoygOBXSZMF+JbA
Rh3s0icxqoKSHYR1bBc+U6aD8pWWTp4c1u2aUYAqhgU8qdGf4uCk7aaUmqs81b6fCteXwnOm9YEd
gYG6QSa8Es/5baeyG8XSB2RUxyIPA9wZXyTYIZk+QtUDaj+sZAKOuA/WCMVUaZjDxwwOVaBX/oNQ
ku3HtIIbyKHyve4Xs3SFY3Gh1gOJpBTSdXFcrZLwTHFDfDIKyJDUjpN8XLFrO5MMYG+s1IOJoQAB
g0ic/ZYpG8Sqxqf33YkD0imF0YDIYQnsXco07JcSRrhXR3jHZu9sAIwGkXvTAiKmYKyeuEhvLkdK
pPHfghHGP+9S+iAXVfAIJfkbi2zV5TQg15O8t6lF4K399UR0xcV1zukHl9AaQP+KzZ9F4RcmlPZ7
trklK9UxgaAkdIUzfeZisOvbrbMMjjkwVHoJIHfR7dj65ZyXkYjcKJq78M0s3UncBxxn//D/zp7z
j23Oib2mL44g0omUGf+7WVn4UzR4B7TGGym2yMrWAByvj6KYNX6aqo3NGp/Z3EFxOO2cAefVgadt
4X/T8xTE9rHJ8UipxxJVnFZ/54guhQednZd2AovHwRLzi5b3LCMtGq1+AC7nnqJQZVosDcuFk+Re
gCG69o19ag32jWueQB6dB4NfqMePGzQX9ALID4k/HZWOhzXNEdiaQpq0Qv80ZOCrfNL/XLcNzxv8
g4f5gTs5GICcq6By8Wo65rpHbctRPkxsYRYEY9D0nKQvRwlzmMKNHN3cksrWqPqOOXAu8F84lzJC
XTyVJxrFFGUnX3WqBovecuLdaaZx3xJJIOWkpbA+zT78ruWS5i63iiLDMtZbx3BdJAfQ3LBXU9aZ
b9Lcc2zQ4WBGn1vsltgqOD9ArWgOD8K04aCWbS4boUrNO8BITOgSjTBNG60m9bx9PQB+RQSH/0Al
fdjFUJ+shkc8wlOINTAmrHcjLEuSzm7xTrBTYgCKzsvBOO3ece87xa/LCXfaBUZMZIEroN4iv1O/
Kiipe0Hs62k0RIZCTDkviPVka3/en+shymv12XfTV+hTmrz6170h7QCQOq3lVp2Jf7J5KXVtHWVO
/imp1Yr+eXVpTAPG5DHqdoZIzBp84XiN3jZm/mkInn19p0H0EYyj6avgtvwB+WoQO+NCXMEkgOE6
vSZPDyJxVKCoCy1bZTKWqnD27bJsu/yhiKwNPTJsw5nLVQmqjeqBSWaTLdHjaYIfSwROQDldmTqv
wev0GDnSqGq2qc85+HOzrGlIWJYN4njkt6Mc3cGa6JJBI643eY+SKHj/a3REvouIBemUZOFIw6e9
gk2tjA0H1PAQGEVglCdPY9cTJFsoRYJmXjNDZB/o+oLI9Bc5ADralDealmJ++odtA7AOk2ZU++R1
GZLHdEGZdVFbodDhU7AxM3U0uZ1kuWQyjyNeUs1T0mSyRYCOWfmvnIfb+b3K/RH37l69kDdad9ZE
sgMP0Q1KHZSMPEfeKc4pienfrZNW3DNOe77YuNOW2+JjM5dDTj++XzPs488J+09fyQsjMFvEVHbH
W8/w+uDSWrErvrQ/9KwtiNOmFHkA3kk0v+z4nusCBa2CXi59NQY2xEvxIY1HiR/OeDBu5fHH6D4b
5wRY/eV9x4t1y5Pjn1FRnwU8fNLeSEihnz1QF4vAPcNzzE0qcs3bcOK96Xa/9l3+NtbG33KrbNxI
AxLo5ZUdNtX+zhgamcmTlLnY9ltPQiM4vGNymg5y3BIC48oTJBkBFJZimuxGIWwadBSHBt9UeOy/
KX30No5NWAfL/hJlCGZdNFTCJCyWuZuUNaR8tqPUNov5wQxEH3UKL89KLkL0gyFVTTLxO8eXtUJU
y4tonq6ceI9mb4f0a/o4TGMbz9t0E2N+/3b4PXtNZEdziZO2VMP1oO+Mc1ptiQPgiumhkClzmsHv
84QJTwcoy7Iwld8SLJ1Nptr4njxRH5zYHYnuLFpN/9Oi12ASA4J/ldmNAceCVQk5FcuV1HBOfWqO
HQFUNKBeItZ1KzCVIxffs0FD6OkD3J+xBcM/0vU3fgv+/YIns/73aJh4n+GxuA8PoNhbH9kjWAEx
8uwD4RzoKXuEDIrNxhN7Q7Q/+TZ072XnCqioRXntXmO8BSVZuWo0HJHb5ywVibbOu6QhL+DP+zRv
Sencq+GAomdfOIbG85xftCXyGZQRWPkaIZTW7SeBnONVNxHwE03CbVweV1XX3f7aCBqYwxaweE77
FGDSutVnIN6Yw6ebn7nQTRWn2OZp9KJJ1Zi4kL+74Tk00yq7RE1yOZAULWqiUmWrzJc5TKwlONSV
zvdgwjuHmA9MmZu794/GizxXRpyxPBwApdd9e7ngiaHhC3ygUM+qtLr5O5qt5IdFNUEfhTJjn+pi
gyVKUpicsHIjE2PciRrfAhLMt844k4Vdr7tffZLFIXnsHSnBEHnjHkN0VlPLLo2xjIncbP0q+2n3
Q66WFOTWyontNaOkvSDtCVoFFdD8e6j8rJmWH/LR/5iR6/YafBn3o0acBQ9O3fqSKyq1U9BAvHrF
YW4XfdQyJ7Di/x2mfl0kZeCjawpGuvBGD++ovKhJVSnV8qEjU0NQRKMQXPzlo4iAWw7i5KvKbOl/
4R4Ug8BZyRHJi54+l0A7P7uygtQ/O91il+4nOPsdtW7trWaNWzwhdYw/i5XQ6xSXb9MFJw1Q5tPh
1wPqwrdGnggfdGF9rq3PuAueF+z91BhECqlt07s/2V2kRtyjbQkY6uNEzEFqhYx66PnWibLQ/bFy
zzyQtRLKplIJQ6lnEEAfsrjhYQYdkQoqTDY1Z7Uqt9eL9rrJvQkC/NvUDV8lg2rxtEuFtHx2Q2Gf
saTOJtvacF+we3wBNDmvTM4FOpEEIyllqdCvDf4UrsDcyFpS+IDfbIlHVe8oCDPey4RyUCAaLycc
x7FHQmR3SiZjBEe9jk69O10GrnQ/ZshIZ/rhHKeSLNCN7ZPExuxOeWP1EkIxBvF2cj3ol/wEvQ7R
M+upgB+EoGxzZoYD2wk+ucU/KQ7ihTsSOH98b9eE5wxIKQsvvJcQZidob/TpLh/XscQq7hxfYi/5
0Tdspo7a+uRo/2g4LfyOdZhgiXK//G1X4EodIxPj1j7E7Y3fy9IuxtaChaqu3e2HhM/d/iAc1H47
QUYPBiR252nsQDtdjy0Up2iMDjlRO19Yo7AFHzn7J9dzlLhBeR/GM9yZYWco+xJYUfFJ/lVjup3m
kVH/DHIlGLQoyAIAsOBbKMvOFHlwOdt3xXKI3+oHjdfZ8AjFee58Hr5L0lwtm8YXi941+2bsLb+v
lZKqL5j1wOF76fW0TQf1dhDHtRaPERVb6cQU1nAbslbti31PhKPow+noLZUVNmNrL0Slc0kfOfNf
vbzdfW2pxYIIunQVLPDS6LviyWp7QOo1HdzTa1yAhCba8lWvuXP34zExGubiCYY7y1DIaXcOOn6R
C5rav/JepiXF5RX1oCCSR/MGEip45YEvwF11EsTqJisp65mzaKPBrCzxoeoAfQlEgU4m6RpSrHGV
zabiL2BMCe63ar4mmBgx3evKnn4LKBAqNomEHs+CTAcyIkWiH7V0Fv+84ymSOfngwILTWHMQgHL5
5BSPOKLzivhwwRDi1mJuZ31UsHeiPy3mzKxbFIsG/OsAc4uh4rcxfq4CRxmqzEWPfWq4y3N2PJW0
TuZrWz4UVBpMRucWdLdqg5GSSMD4JzooYLZccDY4ojXh6V+5MjDewiWk0NWcfTjlE7/gMCUTVW0l
hIhymgjIB+Prk2+9reKqDR6FIU+8Q3yQwLMQhODqEiO94Z83Vm9McNuoTP4DzMwEvotWrmhhafED
Z+LKMIEs0+Wn8JnmA59+ajtpsKgV3avaZhehkTQLNJ9wzu/OBZiduxXE+3zygbvi+GBLs9oBl3na
4pteTzb5mO2/S9zvQeLkXMuCK+SPwf8i7jUA9FN3Y2z8D8BQ94NtStz1BnBmNeCDXcIofIaRRd5E
Yaq6ZaQG8eFBmVtLK5e1zWIz9BGQLBEW6FXIRCXr6kKz/e2R+1fkpN2TltlqOrL4nIdtCbQgW+kV
atmSPpDdGvBLT3neTqDBA3Mgu8Guf72xfJgMExmmfDd9ESIu0JZX0LR/xdPP9VwgTBGNaDdJFyuy
32yJgriTQP/TFKSv9tu+KYR6kjb2wQLCUo4dIKcbyInTubABK7ypzwVOrWCDtLQkhatAYPs7XlGT
arGzbudlQt+B+Yv63+psWbJegl76Pii72GF/IwI7sFlTr3OJLH44mzMfE6fb7Lq0jwnW0NSapvOR
apv/LFKOxVkjTWeW9yn2Tn+0s88XSACmYJEwVMA0fz254q4gn4frnEp1U9d+/kA52OhmdLGPtLCX
s4u5EPSkDf3vV40oF6NR21V//hsFPBuMNBGvoUHYZL9AuUgELAELtgs4/9cqkNDKMVcs1jlVkOUg
9QfysYqS6CT6+Ywn9dcTfLDLDiq8LeMXNPae8tKs8f/Lgjf+UCPy0SQVaCfl14DMekzlS3kMdY8I
9Yel1j5JFDB30c+FOwKEj7hANSFQSTFILg5/24vyRjN6HzsTFCaPqlRAEbTY/0esRzeAY5VJIwjm
/MA7amiN6oU0Xr1dfIlawV2DgUApgzN0ifsqZAP7c4pcNfEhKcsI2IN6DG2zL/PXHedJbq/GiZii
Cqr1lVudbPAzgyvPsmCmDkRc7cTTf840JfuIsiDCdfjwle0Ugw1FjGfqtgr2GyK4/wQ6qChMoK2n
MrNn2tQn7fcLkBZ2N0/PvZnMIy+iAwAxTe+W2Koqi8PM98a+NBsbriwri01fO51FCXKj+9m4erte
MEs1+paoKokdpb3EGhu6YxPac1gnfUQsEKTOowgrrSBaZcByExaHtdteWbIr1xKwC0omq6TaTYmJ
E+vOwTjcDfVAspUii0fLzMu7jqYxhe4B+Zyq9wbkxrTybImcd1hRcl70NQZOvYzd5vAESdcsh0Ji
ijyI2UO0HsaGfdS6M9WdKVrgkedX5jaE1P2i+wZCBmbFt0f4BftuwCcP1spHDBW+AZ+HxBmsAGox
dzkxcFJ3UUTWYGyjbT0RVIc3BH4St4Jmfx8sfwnNV9vSpHIk12JKqw/v26e+X/mlBSXwvSnM3VjP
vTKYlyuVt5aFkM6HtQu4RMOh6Z5K4oSTTmu65koX4cIArBJwRuAfhVy2pgfu3wkooy9tVYfdrHTj
6q4n/elc34EcAE702ibnniU9ruocZPp7Ql5dznIikpUeFwaLBBAW0HkIR0pLBgsDDWmpqPpmBYlD
PcEtJK8ddPpOdlYYmuZD4jqdU1Noo+tQwXxNnEEKzXixd4C04HZu23BHjCLqUQYnv09l05Le3ZTT
Hf7wATnuLnHNqHatWwxoeidC5zVhCz133bEfVPOyYgUsumSebjuchLXCwzimESI9geVrCAu9rehQ
ZLWYxClQrbpTYN5mWdjB7k1o0aiMNKnZ2Y/Y4/aOWo7M9n8/7/oT9qUvXJSvVxbPuF2nMJ2Qx170
cYRreN/pjljnPZU+sXPHgsVWO3QMhFU52KvmO44EMv01AKB6QrD3jZU605u2vTjam1xNXTQ9tDFr
tQYJDDtxJ2hp/EJYE3u9ofLBpn3k9c1N/1tNxifACMC7Rp3b/Oh2OuBwp0XAsREAC2fBdIQT1Ou9
Jq8G84Ft/iilnaMAWaFOM4wHJK6TQKViHNvKkkgMZVTuvQgGkzXbw1uTyMpXl66yU7PqgHEvaj+E
TvCS0Mk6FIpT1/iCiCxl/ER1iqz0vEn60PW3o0m02kA0xSWucKMcbAVis4ov9p9CHDq+2KWLSJ7b
NE2BiYsEwt+S5bTR472zRBdKxiu7l2Mv1Av2mga5pQHCdvmSIeSkwVzbVEBnSNOLqHsbJoy+mRpz
FBFZH/ohnAlKAziJoP9D/c06Y0t7oGaKK237EzThrxpEhLMO3Lj/am8z/tOifeBU6MecK7TaQkOe
CkwWgfAgYF9kXo31rrjutjeKN/o1jDSdDqvYh+u8B5zq0Ql18DVEw+aJjBh7OtKAlwhVtauwowWw
o21ZdF/7j6ncznm0q0R4cSjmeke+pSjHxL8wyQ4dPQMcyCqdZY2Jeb3TIOP4zVQGmm0vuwCaUJ/n
pCpD2U1E8dQUw0BK7h2z2L1XP72MgfMmvFkJMdJ6tJwL08nyPav6MN4Q6jFHM3oudFnNbip0MwMQ
j+sLFNp6M4zro0wQE+JQ/O/+gb2VOR0RQg2rG1phpmAnGEe8Rzy4nwM+K8U7Aokax+XWhZLkMhHE
8AYYhMLwHGdj8WQW8rVXHlXkz6NyPcWo0abUxk5JqN46iUZWXZIUPvIIgEmHiHgLINlzILddmejQ
q7RYRhaJGAJ29NSZhfh4r7RzsmkQ3RF/Wp2+Z3JKsP00XCA3ql5DqsHra6DWDD8NIo988Fb1B1JG
Jdimm6Bp7SZuBMmR3mXW8zZw+hKvwWmkmHBKqHVozP0GSUvGdl2vcRmQcyFcAnitfRxb+zQ6Pl0m
IGAsT5kAmrwLu6icnOmr/RJpe4uSO8E9j8T+ygE+2AROPHgg+FWdTl34kGqOSjFsgAueDJ+D+RVY
qayya8ixc8DHNnNW2HtTKVeCXfx7EjXqn5LgO04LHFbKattfxKiV7Xc/2YPCysclCDPmA8uBQiBO
ZN6qJAxNOxlByBZc4fsFv/K0mqIwzqvtzY8SOjYpEkRKZjBuJdHYQM/1+qh7yY+jSJyHgADF9v0e
8Fwyt32lfythloqxiH9awjGaKNF2xcevMiTs949Fl0/63YaOVIxqbcCzMO+3zvhfBUmtTyLaFSNr
CsVUmwm1GT9e8/Zls7OIvxM8YGhEe3GbnFDL+K2aLGBf75ByYRrY7WIEExmk8DBQhg69BPWa/0wr
ltoyGPEMtYjvazpHGtvOHCbxNwxhcszbGFv9CSz6coZUWWFiyUnZ5eiueoYLny8ubJNXoPg7dAwy
ItRmjlYsfaWPeEPppguRKO5AzTUS+6YU5GU/6dBnwTthqBRK2ZzqacvCCNERsKv+F5SDtHfJJPWL
2hnhZmZx8vZTqMQADGetq84EaEttFbnPzrWOkw9hSSvIrHAb7ozT4caYllmI2NDqeidV/kwKgS7R
/4pXiDIgP8pSqww8RMJYzi/wuTXtq6iFiYH/52V7nJ0GjNaN8HaH8u6SC686EbTfW2dTozgFHDe2
dyi3yErHSSqNTeZm11FZzTKrW0sl+feBdB5u/cgjwAVQ64vQ9dsMLxqnUEIqVFX/gymSB9KJvebl
wx9YQ2dYVv811MYujbEkn/I/Pp1zGl4FoLEmbTj+MjvGj3IK1QkILU274g4usuN5J6d1QyYTY41j
YPxLJwl8kA3DNpGkkoVb44OdrznIFGedDcuF7QxkxJCTOaGaUruVN7Yv03yScthy35FOGpRQRwUf
AGV2/poZAwyfNbFEL+UJ+OvJGbGHn/a9BV2y1InUblIY1xw+Vu7CAArKJSC4MmwPGVPaH9d4RHdv
QcmPs2GTE/ST941S/45WJQ1U5idh3/ZERxkvHkC+HGDG2AOOubVKsmNftiTch5yIeY5GytYcUPmA
+4KfZTc09GAmO7/KUG/Q5sz7zFrzO3zvNsz0ZeZCsY9vYtT3WRvOiBbwelPUzAINS/qu+ZOMhyge
4R1P9IirtmZ+mPuZLhzMVMdwuaR+XM65ECaTP50EU2sqsIpTRO5ZIC+/wzs2bgDEQyNxCCSGcbEJ
/gZceP/QCG8t/JfuT9FosJCwoe6J9tWsSzY+yBiLPXnBEkeCZi0YbO7ZC4tqQ2N+RDSLLdSPizP0
R+GhEPTIYKuQPzhc7tm0+chWc4XBDZOzlgLx1iAyEIGNUueeafZdC2b4G8ymAXJA+hSIbzNHVTVU
x/rIfkk35CKojbRZGgMM/bNufCWvOuRyFK94RRTCGv74wFjtp/vRh8U/n1Sc9Q8NBOhLhgCg9Wl1
MUT8h1weVf50Ih18z1crpob4PC+zyCBkZiRuZLWwH+ZIB5lNRgjoqd+pE8jkJIxbao4dgtkZxCSk
zwVcix9kwgN0Ta6VuGU6HACz2pOeuJfFTCV4BTce3m9f08Arl+ZGt3qVEqVz1U2yIrX4XSiVcpcA
JQ/8cwr7tS+RRaYaedvnICqR6wnJD40TiYZRf7WCtzo72sQMV7ydlN2eexMRH2ybBGexTgi8RidD
IdEu/9iBDloZqFP8/6E7r4n1eGa715POdhMt2aXefyN5+wZ53bc197GdovSMCzl1qelTxZIkv53o
1O/QRe2GMejCftrWYigxHCdu4yMRBkqUuJohWwrnXARHIdRoF6wL+EmbQO5EXhB9MsVPJU8M3dUE
OK70Sxegep+eGgAfqcjK5W+aMXw0fVtSLtV2v7rtCdZJTnKUTp3Rm15abK48LATrekgclwSCrjSE
i610zQnMP9RkeQ5tWNq6S+fZ42BfAzdH+Ro0uyhNj6S4AJYuIVHhtxqjrpaCcUYLoOhCzEWLP/c+
02rTZT2BHoBCG+zq15IFDnaBmdpZa01Z8h2zWEw9xsnKu6cjosBYMbojh2ZPs9QUVRSZSl7A8+3B
Ijj/2jF3MfZiN4WleOtogehra15HMdhPtkI6Y9oTroarC0Tnoj/qwFN57pelXH8Ql6wEH4UqaiTh
3fCS6/AxdKAQJXO1l+CstPSVh4YumAxIEzkRwRSlQ8Tr0plLkE5WyVTI48BPQIwQMewkz3W5TIAB
F1QueCQhmGvvuzi75OqjhL6lY5kkoMf55TjXVsB6jloy9tApmlSaobIvqj3oRgGD19ANTaDdn03g
RhPYLgjAptaLW4185hHyicJ+D1rpu7EZ5unowa4TqoQTlQ9GgrLLjkDRVbK/8C4pmhZ4O7DJfB0X
emeONoQloGjvNHKqzHZntVf0rhVXNnmh5Btpv1C1jT73IWy+MnaPD1RbH+dX0NI5mHDfssWfL0nW
2GiEEAhUL8T/HsLgC3GYYBQki8FyOzocRXbzb571z9PpqYnqqiYF7NG61s0zkUuNqHHZTjCUopqL
E2oBrAYWAWJwkQ5xt93Y/t9sGHtauh0QI1rV7sJxgRfViRYPEjGVUONaGjKKLEJnbh5gbkpRQgi+
FqpCfJRPAtzYEXDOS415gSTfafAdh7zSpWXCTzv6NIUcg81tONFfnC/8L+AM/DHjPVW1OgaaDw3+
CHH+0uMo6XFBfpR6d2uXfE6vOTpH3aSDtxoxb4uUYydtG/TOHJlESuClwuqVzlbNHCrSTPoJD1Lf
jmCPAh6YCLwg56gI72DhItLpstRJEb8Tnzjz5wmiY3rPzXs9usrfoEyBynNfni3uyZpS2bglfmZr
8j0pLCLdqZICe8q2MEWppiI1YgZ+BRmCzcW5zdkmMAEMx45JzwWj0RblNKQPmIimKS4GNodQYVnW
Ha+9nrKiLEpl+2d65triTC+oMWN4s4VqjaLrlhkWCRcOhK43zKLANr8ol70w8HWoSq0/nHPi7J8T
hjS9Lk96YpULwuYbCWiIU1/sV0ZysfSSAMHMee/iA+Kma7Re/0MiyAd7jXDcrSSJqZfyG7U5WdGh
PUaOznoS5FvkiBEKKPf+9kh3LhSohnQxAy3eon9W2cZSebwR+Q97vKxpt1lD13Gtzq/a4OmhfkqF
k0KNyPWulXkO3+oOrYx6J8ZikSaoZNxc+R165y2Vgk/OtPQTiGq6ud1Q/QxT1bt7vczumn46l+wF
34cT11Wid3vzp4y6dPjl7cw8A/jFXi1oklcOhET+2x8K3r1Rl0DxH/5Fvxmg77jQ9mF07prC3fVo
RUiaBLMFEPtxKD9aJRBw1uqo1c/k84XbMF+zEzOUy/kcJyKwfr25TCWmkYRQb5GTsxzPdzERkxE9
/uO15Hvnu1Hmbxr1WeZGJeWVPW73+PYHIPB5p7567AH4oERxwbd1k6gRRrWRoA6xhNF5LqKR2d+B
WLfkdxkFmFU2Cnicu3+ucTvzueSorgOo/AMW7pp8xLeFEE4u3SC12mNuKoZkUTDRGhMVVibLcYnf
uCa1+m7xZlhEexsmilrzeeZjHuwqh2iO+zoOD+Afdlep8zyiuQIOTt+KAd8RTGEJKXuDx62p744k
ZIK/1N/GCfmYBPOFrbxtHCEyidCzn8qmOFah6RVYnke3PRu3lGB8WUzMuw16+U/yvv9aFXC2ijyF
ILtfClH9Q2KLeAgi48rt++nJO63kojVB3iUr4t8G4LEXW9TqYhwDtVOpXZydExHG2Oq/p+r4VLe+
1+7WWPNBA2f4zfkkP/tVgK+KklNpNZeyva/DYHM18xvUue5Q53x2RyUWNCOgu8ZKYE93QfbkvZ64
V3OayMNjVlGVLwcbNU/GxSGE0GFR4l7nltVFgki4/aYrUhyvRh+kljeZrd8ayJXtKMq+D6EJEOFt
Z6x2lFNZ6qdcpVqjD6UjsXWAVSTEVKwiZ6BOE54T69lS9cIepry1xLbEc+PwO2K+cyMSq2VdacM8
90tzruVMNb3HWuitDt1f9Lj2g+/e3iN7Lyjkw9fUIC29achd8cX06wMybs4mD5rfJRpZOreZm4LZ
LnIDSkBlyXhGZa0T7Hft5jcZ5e42VdvFuDqzHj6i3vFIHBdznNJSj2wq56BmuSPiSrImCso5lRYC
hPSlowpMzyDT/8nI/h6xNsRUqNneAviYtpsAjWK+72n+wQaY11QkMobMYfywbqb4DePDE6r7z75Q
GiYLoOvJPeBwY2Dp60LwI2gwEydvp+NFzoVL9iBdSJYhUqIV3nRAcQzlndazoFewO246sbAtM4zT
uZgfXazXWCAtASy+/+/8jRdFGXI/2Shl7JmfTbjxUP5O7i5Kt0owqDkw+h2Ol7PFXI09gk8NHWe9
UvM+TaZEL23HNW1K621egP+sHZmi1nMahXgdY/0ag1C6GDMQ+3X3JAmSjms315IPXzQuISyZiRg8
5p+OspiWGiXGkqDXGGeB72BNCijfGqxnsiMjlF0re9Fav4i8qVUy9XyrM1WqBkB86ERpxodtb+w8
lVyECnnIOW77vwoXVSgOfj4FOOUpid/WBgr2ZlKJYVE7Ek+sq3nYit9J9Mt8dr7lguX+rMAy3aN2
FkXrVuof8OfdMbn98jg2elpMBlW4fi8Mb0Lss5DhspCmNkt/ya+L0Nv26tx3iE3jt9neQCTAuV1r
g9wb6dffJmPB9/CoNh0oHBDY6zuE2CZuE5J7kVvGHgNdKaVEO5ep4xY/C3MVWOKqB0KOEq6elatD
wcm7VmRk2pZP6n6Jfal+mf+UQYiug/NdpWYe1Yp8bCkeMTsQujITF5Nd1x6gFhONMh/a1nPC8hCW
wkAEpOqLR6YokYVkqCshw4fmHiOwGBHIg8l8HPIKcgUg76CH/itz4C/PXEJksppOsvpN41Kd/3FB
HSZdX6vT8Xy70R2Kmnb3wwZv2zrI22PSmo5viu7J16SztZwf+7gAyqUUDffZTk+pDrXAQ9Ah5PhD
LEgbPon+BnBI24dm8B4gnQqmtrpJ3vWTNXykyr2MexGyrSbO0POjlAT1LbvtY1S2d+alccTXt9t3
FEwQPYuq2EJK2N8x57Y09NWgxPNolgWmJ1bbPQtMMX751PLc7hU/FKiFTz1UCDRsj7FFTEO/HMbn
CLi2i07OQRmCpw/FGwv9Xh/KxUog6mXRapLUbKEz0Y9TMQ83OFLOCQhJfrtw5AFSFDf8rvTtTOyw
mhU6X44cvGNL9ta8Xkcu2DMy/WXQE2L1aAGteuFYSjS2k9I5WdwZ+gaFqCIZi2/FryR4ERS0QQUF
0SgE1nPBr2Y+RaFB5IBJvGPO5PvKGO90L5S/OB6kn7RYDxAWUyp6ljIg1S1yqQcolW+FCkbVQlLS
8lbdxXEyg2ZhhQE5IVzbimjUcm9ugUVoOYfoXnt05iY7iULQ9wtl7Ioxak8y8CkmQM66nGwqDZo2
i7lkhobfCgfVFSH8h8nBJJ5VpKUF2cfA170ujUO8Js06DZqme0BxOoL6L4Q5IoUG+FsdnwNN5xWi
wUx2jEybuPVhFFz7Z4t9GOJOHi67rQuFnZgy699jY55MtY3ouXr3o+9Ea2+z43iE8xntf765xNrp
wU3d4rP6fWHRmMGK1OiMo6KVj2BgfRzjcJRWC0PofP/cSOTRekiDJwYsJ9cS/TyWzckFJuFkrmVV
3Wo6LOgNfWdRPpQ6T2jb3LKb8rpJWwMaJ1w5L0AZp6s9YYLTCJjhKRt6NhEu3LNOxVU3tNrsV74o
g7ZAHcxTKc49QfD0eRfm2RNHCWqqoPMGpoMFLfV6Tkaie2wyCDibdVGqB78Edvg5KjulTxx74uDl
I/Em4Km3Nk+no2ekILwMiH03lXh58Gv9Y1n3DL6NeikQzeX/81arVmxkzsm9U2lb3qybAjibKLeu
ZqLQZVBcmFFV0xZW3uf3qzcjQ/cvGpaiM8rcDpye8jJxqiAxXGgNl62HRUFI8jzpl1GqLpmi6rmg
1bnSLgb/ekSzPGqSHOWQ9Mr5qXk2jiG8Ip64OfY2A/nyb9B9lRKc2SXEUEPyuu8BOXW6bVNmgvo1
mQDfTCS3/TsSyIGegohjp2F6cXLBIe8Nw1qua1+ZJ5Up1LaldD53A5Imtk/+55XWN1nqXDClbOTU
lWkn1yfqkGuqJkljJIlLU4RBhvmFCpQLmZyLIlSpoZSnYk/l6GpM+mQFhOk4AitFcwPpodUycTxT
QwoaxLi1zYLFP3EIoL+v1ccdnv1j0LZwn0lduLD2jHluV57WBSTbykxWliVngLAFUu8Rz0XXUzyk
Awp0kQd431h+GPYuVDzI4ZuJi0LI1WbGlpt0sYW948PoHODMOuMOHM4tcOmCoyKbLmIboDOdqTsB
6VVs6glo7ZnhlhrSRoeYhTsR59xY+VQFy/mLC7dQ3yXryyysidrghTcFXtFEKUP9cu77fD8TF5Ts
c3t4zvHbkuFxTCLvKJj/RhJos5iQzoeqRxxOhKu7HSYQ28gcvvEDEtnyPGS3Mx7VFMsCUdTU89Bn
9v2EbvKTZnGn8fX07yyy0XAjg1UJS8cUuW7KVg/k/Xcz0d0bFsxBF69XMPsmTAcl+3jgLGLHJC/L
YxXoui6pyvokM3gMF3SBAGkN3Gg0lykncEJqjqm+LcKPtk2CWNDe41I/9NxHJ8o8DBLnu1iINgHB
QvXl4AToPipeeVdZeP2gMstbYQ7eqwukDt/IhYPVzZ6s5yGVCVwEmK5t4HJ2LJAnr2IGzKmNUt5j
FL/Y6aZQcJENl90VJx28Cm00FoAevo8rY3e+01dPoOI66EFv8+9kK7PVpzaa1q370YG4Fhw88AIa
zjesDT8NbG7kwuipORf3YYBDNXBzw7db6OhEX4pSjKA8yAh7blRDNqWj5g4tiMEbhV/EqRp2VT70
jo27/+cL+9bIp+k9IJRW7lZTzqetNjxFQ52Su8/NilhZrAFoRjoJj0jS9VnCyDXHAdeJ5FA5SlE1
nnVlBxQ1tE7lS5CU0MjmOw3ehq3P3ihbPUYaFPgpnY9hTk4TqqP+Zs+0JsJ/hsflP8mZma15Pt0y
SiY4yW5+FYqibwaULAO/Tke+Q3lpYPJ6cQcJ2+9lmmHJhHSsaFX9Cx4JyUbjYawwWqYSJXKn7+mB
+7m9mz2ybPurSDtIHPUOXDT0LAab+dySdqFR9v5t3mkbMMzWgXJCE6AyQmroH0+jYHMRz9prCC6e
AyuwszoqydggI/MeLIH+trD57z/HJtEdUakPCNes4gf3V+BZWwiWB7M8BLH8W+TivvyJqeCiQFGi
/yypwV97P0KxopaVry+OAi1o25XBj6unReDbKjWf2q40qKR7ukmAZjqNPJDufUu9xuJXmN+Aqmfj
gokepUvGlkiWcAzZXvW1b3knSEKncA6DuFSX7EnaLP0zbnK/4kkPPzorLrG09LYNaERh7fBWLDnj
QNuifocBtISLbc8YzNnuFJkNZKiTX5+1W7oFtR2iNK6tHf0yYIQzJijYJdtk0fRv9UHN64d/urbv
q8TQcC7EYTiqQc7mWvZYw1qZCCpBeOW+/2gOGrZ6OKowaGQHEwgmLUkbu53YSPRasng13sJFuLOs
PaO6VHiPT2k1Bc5LnJQEOI+Ppj/eMp/60oDJoskF9bsArib99fXlyNlyje43u323G0RZczLTZfrE
jso/d8zPDOKIlQRt4zyFVXHySLx8J9r/NtefsPakNExpOR932aG5AL3uJkJejnWcUAX1RWwWYI0W
bjnvWCHErewrR8plBgs9fYU/KVEM5fXQuB23TqBm7h6F6Cu+J/3jJGmAxlaKF1hgSS35HV71IQAJ
dQ3TJc3odLLX54OGwyfA7pjSIm6vHj9Rcj+dnbwpCYm6fi5kYWVw3U20xO1JXt04pfswRJtSSJoP
wvt7smZvZR6DZVmUU+9h3oLuQLYELJcx22Cenm0fMV/fctgjgZtRFfQweZ5nrlRhv2Er+XJfLViW
mzZPd2G6NJl0PJSBxLSXi4wMMhQB59jRfL/3b013J8oewEc+GtOE+XVJ8xN3k2pr6h53F7B6W2IV
mGo8wN9+o13vPN27veYUTaGLSbcBCYkmOez8UjbTGpvV265W2f6E0mCzMVHzDKlaYlzKAXJkQvJi
ZvyYu9y3SgPlhcr8PdMjkETAYHnFoBn3J5Yj0Bwj7ANv6iWE/G/FIsgMs8gUTiGMvJy2DsJzveud
fkuz9xDY4KbQbq77eqL1bGPsO/9VqSxE5MrILYTLTwEcjm5v73wxEsyjqj7n7pP4DSvdGBc55UTY
wZvtbYX5kbUdBNU1iJxWmk/8FL896JCAWhbScq8+JcaywOetd82S+51vzFKIOjtFuGm4OpxDwwBA
RUC0fTKTxds8H9eYdXYkAGED2xPkqp4CtjZAffy1ysqGbjbjBWtWEpFkt4zAFgpOLCwb/Vlr+Cv5
yoaEQet2RL0fFiMWJxf/IKG5i0bRwrBoqh1BwsErnyq9oRCjVkoJA07xFNo6E8f9z/o6PUjRQKuZ
lCI3gf45XUzSvKimN/2SJ1ZnU8DDdGeSVJsnWMmFSfw4rMRKnoYQQaQlZXtJb5TfhAVGilVmQYOu
M67JF2wUtmRZFYCmP3TUVUfbBWwb8klLUZEwI85tX1cVv/LjrIM24agdET4dU+psg4gkPHETMIwi
9T8K9CAdXHeby+7QVoyQ1nz95yHkkSIl1Y2g3QmqNZzv0bDlQcxdgMIplCbAndm4hy55SFOvZu+d
AawFQTzITdQgtAXwLLd9dSSjlXZ2PHhXbXx9c1zu/1ONp/V3+psZrMuNA/wgXfXm2KU84bDt9nDl
ifIz/lF8jDd5V0GUuniFY8n++pUQE6lu5cad7hMX45tWBE0EYecsC3+5volTfEu01xrjBGnTwNTG
SFHPDNdtB5okd2jor84n2C/eGxbvPTi1G5MOwKJGCl6q5L7onOBQImbS6aWRZAoTaG0W+2zZnxeu
4xbtEAwt25S8d/mZuY0yUlmOAOiyVZLjxu9GSKtEjz187wkzPsazrrU18ZQ0+C7r1eHk9MGvWiKc
eGrww0rt228jmjq6pYegrQfCGkbCdHPpYVYNVai0HtycAKJ8gy9WEG6VzIdvwv8uWQ4qgMRdIeFH
P/hPaZUHR7Kglv8j5jS33mK8Mpx/LeS0JD3UFlXjK5m7yukUTl6TGlgkzuChsPjdZI7/44yGye38
b2ERfEF1cLWcVHPTF5Dj8lzOpT0rzlQIDo4rgGNX6lg5l8lfmdAbW9+0f58C92JweE6OZVFtn44u
yfjVFLED6F8gY/6r13u1S+GMStdiN8XUh41tA3Gpf9DkPv1XdJQlFz5CT+Xgx1Om9DyGdoaQ0FxW
04xHRmvbQXQiyhwG2zYILTZ+Bf6E1fllE9VWD8/l11rZVTsREDbjr4VPYWT8LNPF4lmXZGX1ZV/y
dQI2abK1zs8oM6FMqCEEjkdYHbqhGtiqFIG2lEBZ1jf9iL+/tkeu7Te2iqXM9feHbYIUSafn4hvN
X4A0RAdgMFiQmRDbE6+MYN1AwUCw36DO2jUA9o1vTqxuDPdpA+wz+AMa1HkqIRs920tq5pBLpdlH
6t2E+ykNBAjoSsISMZ40BAjFskLKvibUfZAPHVHJ4ANsz+kPHesD/KmpR4KO5bCJSn4szVxr1puN
Eqvz+tT1g8hJeBPb+0UirCdXA9ptwdvLPOJp/1Uay5BiARC0uk7qbGRkaXdRyo3kxjxGCsBQJDz4
TcfCM85iN3G4TNQbZc52FsdvMQTD6i7WSUt/8i+igkvWJuWDvD/NxNBnDl+D3xGAsr7Z1jyWZQMF
jFv47ViXmvpmTlkBZfDXjrKhsaoQJfFT/hsl9stnu20RU9+ZjYjsMgH3zbg1cRip93ID6F//6Cn9
GYp+ZpLlh7P2SomPW0aPsSnwqL3yAw/P76J3c/aA5doti/pP1v7WCevR85xdBHMCEhIQdEukc1ap
3WxvQTJpE0oYxDH9crSPm1l6SrNX9auN4TKAc3RULh057loxIdm8/BnmPaOYByULHwkZpGfEu1us
3HkOE++QrfKPcDCg+tB1DHR68gcnwdAvyvbdh7oMnHfU8suf0NWz7ohbf2jAwPvgM4laUCZsCGMp
eiCgLccMiBE+38ECVzWwzJVgUIZl6nXKLqxNFHqs1IV/P7HvE7UzeFb11odhDSfLEm/uRgSjy9fy
wiVAvUQmbMpjWJWQ4JY0MAyx4ztSiPQukbgKhafIqzx4rmiD7XXQF4R4n7ieTXljtK01b+t5yV5q
mgHvN6h24n2eAkh6Jlk1C0O/jxtWAvlKhy39WfQvOcPEMBbspzXq3cbIA8XwcfgnDxl654oM39tF
u32lf8qiHw3ROhcBP6PQJJD61eR3HmZmp5ST1wcju5mr6FBUKcX+sQo4KxMxBC8ep1Yll2lM0xub
U5/rcKsXIoWA5LhvxlhKkghgAue31YlFA8hOsGBz82dgYHZdxT1rGzCbZueDwHgILAYEMtYiejnG
cmjqmmSNay+KWPPMe6HiKQhH85hN2abHz3seAjE+rvOTH3Xf1qScMtqqmJl6DJ7ubQtojRGfzZsi
kB3EAdLwSnbJBVkA9kKDOaW58l3kxTXrIiXps8+PFFsIZqOXGTRgKdEz/AeiU3Fp8VgThQ2UGxju
+v/9IQMSUGhM6ggrcxsrGGYnWWRUek3TYILCKXUPC817OUJhZUxCeSchdHKnbwMlHRnwW/oR7K76
vAHq2Qihbv69nHesl1/koJMds2WIQ2ly4cTppaSDfgz2ugUQ+aqx/CrVOP5u8HTkgqeT3ybAfo+J
IBx2h5NJPd5+xFZVvRP2y/gbpMnCQW8GGFp2AgXKpqRAX8hC0KGhiCwmxUtyaj0g4Mgq+ux6s8Ja
dB/x+Tc3UrdLi8fJ9wsVFZAVdy8YibpUcisSJtcks+3lo0FPPm86OlfPeD9sQqOXh61bSi6pVQn7
iMtANJmS5mPDfIIrhXhQJcRDM+PaYfsUOzBBCzL3lx8bcZYSzBUx24wUbNBJmNvbbzSK5Hvp29wq
EIs/jjlE/fvEUtqQXJIUDe6qkIxCZii7gX24tGLSsxAosdyCMBXtx7j9o1DIQZbKAP8mPw2Hoc7d
jQJh5JeOiZv8Lq9edfoNXHa9LqwYWQbGxBZzJCJNpXkCVgTONOv37fJS5Gv2yDfFQJKOVFlayD4P
Hz6ewWpik6W5+xIuy8boAujGuUSqIvnYAxblZbHxPt5UtyBvdcM7i+teAWOqpSJBhe0FlC7TSViZ
kZ0hcs/eZd6gNlJqdrgVWovVyrumzPPbyXgp3Qc2wFCGe19yXIHvDHGcd//OkgpMsYL0bWOVvYOE
HWBq5I1ln0O41K95Hpu/yqH7hkRv+r5GNr/Uv7K9XwPgHh+b/ORdEjPBybxuysfsvQKJS/CYBX0y
G0IH530RRXbZFh0DpRAuPBCMptkLYWcIZdqblc+OJBe1l7QYTqSdg+elc2nkmhloaezc6RLvqlom
KDWtmV855ueAGneAaD2VuH/9FO1z/IKAlVxTgQK3VaIKKjvwizjz68BLWsu3euxCJivsLkQECr5E
Z3HDiI3sYzh3yTCu3g8sMWTkjOKgWagSwLYdSLldrUhIHYoK5fqcvAcDPF5Any9E48E97I1Q4QTH
y/rs69cWURDhUHjnn31wbxfOQJcA0/J2x0WGPtfdc/E71s42be040MYPIEUH1O13QJ94ygmHHwFk
Zb6VQrnVrQJPT8B/PP+t1DyId4KNQDuyw/Q6E5mhguq/ZbQUKNzHPDZVOx1XEwGMBCxkBAUtI4ZW
BFkqbkZipYdOrrSP2XNVmFAtdamTG1babGa2FmzdBySSoGmRuXdhww9Oo0H7I5P37ydVSdX8ul7T
vJa9VN0MoVxtq2TCndCM4dV4supQ5/crtp3aGSoktweAOIA+fN/uXNO+0RZNO5S/BT7jAcjwOUrO
vPJM6bXROoJ3NJKcmXCK+qIdLJpABp1J4BgMInUnQ+Kli01cMY77CnNqJJ7WZ3av+nkWtETtIbEl
DCxH0x/vrKRnXNa0h4YXvgV1gCIEEvCs6Z/ZqyFC21uAXubg+QcHuchyDtBpFOComQ1Ou74x0TgM
ENb8siq8mB1So74wIOzd28+VEGgVj810zM5bsaXSB6dq3QW/Co/9zzRWmqhVy5rEd8wZ9BGe5kkg
FHcQr7Zchix8AeSQegdGoL4DfkkGKFyEVKQAwf2XblUcdYLzvLkUtbfdanEulF56o7tRBm/BhIrP
dd3T07ALqky1Um63b+15F+sCLQp0Y0N3dWAB0OSrNcjvPuZaU81AoQBJC0W64P/dm9e5iLbPMAkx
KEwsdJBV+Yekq6Cg3RkqSLApyYhvkW2Q7McCOVtDOOVT1ZtJBH6VIu6kE2wnl9MUdHTjZkbN5Xmf
1wKvE1MTxgYUFPIb656iEAOmhZCKfsIN3tuUbPeV1RCCmyT1nOqEpPXpVeIbTIpyG5l5vJ8ChRY0
fhnhdS9fFwQMC734H5AB7PxOD0dtvQr3GmC6z4FJ4ehUpmhWPSaIvf9qgibxrmx94RHdOOqCC4xz
diTMmVQGfi97puOka//x6AnMXSJZnCEPqixwN9gegVi3r2uimS603sWfC1HVp1aXl9rGUQX18NMr
yfkLNnAFnu8xXctm3VFgpgP3FSGi7pH9NmUJNgVRUe5x9/fUEGsreBqvhp377JfsIMBuwXlj7y6+
XP17lsfcE1/pf5DMc+p7hw1F3CPEkcFhmjBQOaeepptkO3Z5ltf0tyOZNw80SkSxX/AreFDAy7w/
jaALCQjxE9kca3WgOfYdticIauktBOaBRfoniiFojQxc50aKfwk48ec36CZ+g0gX8GImbSCUucU9
S6/gxSM0jCk76kU1MOEljfmxIrJa0ov2FaQa0fVH1mseY2DgXX2gP+fA0+rRabveuj2bPcYMT2Ke
B5bKCpNJkC8qjQaSJVFT9Zuv10xy/cXXsfZRO0JwJiHKDholmuewTNQlnswG2u1NOUkgKfgwm1c9
jd49EAXf5QKg1jdyN18E6BZr0RuZEYlPytaTi1WKiihXEvXfa3V7+yvcbZEUu+SNZ4Nl1zD7IKvS
RIJyjUnQATwn3bm/fyQsuxTHbkIAWwzotbsFypNauJ5c6lg7YwoZH8kwBRoII47mAJIlZNj9GjhK
4V0Gsv1ddU5lXq3DcfAnZ5GRifB3/53w+rLcYiH9I/8T1q8eP53iuzEcxWz7Rq6C/zHVDG8FSGyf
ZPMjxGRpxK02ubtV/Kq/2IFK6nhyymOMw7fJlGOlNo/aDkXfOPwLHsAWUrGGyICwzYbMYISYvO7p
+hPlAzx0l6L5RNtJaZiVFy86PkMy4/0nspatMg0ma3nLtUlXtcvXmDQLn7xUsETdpIDD+yhvpiS6
aCdeRljp3N0m3FoifPdEQXe8TQ/S5jwdCW6vM3g+q3u60bi+GotKK66dKq8BLyEERkFLjtiTfDo/
6BvhdLWsDqBgB4Gy1D6Z2WftSVXX135BBuAQwjSk06ZYzgFrdRcUSmIfaCeHBuKAUJ0hrq6AK0gW
YVyDdOaTVrSQQTwHChRa/GC8imBqcmT+pnPsyHr0JoYt11bKgcLY1iMcq/TbD9W9FWrnZmib//gd
kumGDhancBkxlwTvDaBMkBFkSq6lDAH2xL7ZM9knxIfgVbKTMLeLuLz4wzMOLGZU4GfInwiEDvFh
pUYQv5DXlfIBdhNNE4cOaJ8Z8IHzqvmbmXFwFqd6t1BbBzBRApJqm6bMWxJ/QjRbePfUJusJaMw4
SFhgloYjkCsveCoMn6pyYPzbRENvKDSDTvZkqTawMNE4tLFFsf7geWS2yQWc6vEuQO4vFdrWpK46
E9AoLLL6mNsTMwf9BvnA4NfJGych4KYSfRw0Etu/H7EhiJ9jQKTkQ1N904E7b6BC705Ezh/+nlmY
hKameXaahyQ56vte+lS+cN3YfZGuxkog6FVbhPbLZl1jivsCeBr5whfudJI9pygXcl0YCk/lEnOl
T2Lnpwne+wxttJv67T6Z6Fk69WJAAGAG/P6FiBCJNmu4a0/uTe8grUBZyDp4q19wRsqfjHIkai1J
/qoiVsUU3bomT9Wjdii4Nrg2So04guFgyq86Z8/ppIYpzJmnPX6Nv9RV4TRJKLt0YgTQkKfubM7Q
bu6RwtaWvXB7cZRhO6gsQJrnRUrzQP7MkDvxiGfZXdYol33wvZJnW4DIAn7m7chhsrLRmG/5O546
NxOzUQxaQYROZq+g4Z50jCSApIvfzPd9fwZcwa2jnx6Z+zbB3+EXRZeg6C6WSpPBTzv7j3XvnnFT
KAvDc+vG1Jgpsw6bQr/T1u/cdrxgRKBgORTAD2nseSMa1JP8q7Cr5oMQt8IhNQWydgNZIJjj9lv2
0slysTJCBQ70ilnSdojx6aEdRzuUfZDit4mU+wgTu6e0HkK7nUVcIvJFBEVwiYhqgE9neWFnucB1
vJ64gPhh4mXvRrUW9s4S1kRpP7JnxLfz7uDux425UusgxJNPsJzXPil8EEJ1uq6NARDEudTd2j8r
r4XPX6n9BdnShOwFxPztlB44hAiGop2sFCdA2IOTyaaGoIQzOojwu1NuLRXlitQTkkcO+8z70so8
aa+4RA7PUFqCSf6TqUsVfDrKZGuJ3CW7I58U+A5j79Y8qwb3fwsMGERQfx9JAnq80pNXOD7sePRm
A0AouiybPu8xkVDFHQNnRUejrc4o3mGTA7MtPYMfE2Kv0Je1em+pNhnkRYaZo2hA4UNtTvp7ttOm
p0nF3RRVoJf35F/kDPU4Rf3Q3UVlNLYmq2+sMw+WjCcNuDSIyQs0NORjlt40IIKNDIrdzurpvSvh
OdEq/dc/mDTA86MtlVpwVExXLAYhpCTV2XzFmNQ991uPPBcZu4zX1gp/joI+ic0RmcVXgz1FC+yF
ORlnCpktjE7xw8Nt7B3Jkz25uJSliTM8SKnfODuLnUExwmMKHipM2sutfrKZbW78D+/siLrUhYUj
hbIp63JxEW17QVx6Tmjn13PFvRklOuljMWNvr480bNGQPkBYy43mB6yR7JSS6M+OhnAAmA7JqNbd
ZRQHM2m6A0S/7bLmDVRlsIqFtRc6yfcGcaJnuTejlVTjY6EOqsAoj8egaJVovnXyjsHxQgaouURy
HJ7G0daVKR42qyxrTOPGvhPMCFmK7MX9ty5tSZJYW8h85y6W7Sevok0ZMFicqSmjFEqKDhCFOXuM
yfNK4roRMpNgG+tiNu9PJQPPlJo5Ygp8UEcg8CI69XrF9gMY43yV8Yv5p8MdE0yv2rMuoZoUioEE
aaeJAH7CCj9OGlCVbXdHaTkEXdj6azRoyk+9VFA+LpNCx/WMR4trcNrZS/dyztBkC58M6pPJ+SLC
9UnWE2QTzYhvg9a+M84763pApAFibRtkT7Jh19x/3ui8Ey3MQDBoHhvWXVCEB7mjYt+T+n4EUYiP
V+6UGbfFXmS53hvQLxXKvJtUjvPTk1+UbbgGRI+IRnc47FG0WPV6TBN4QyMUcTXP0RtQjRHcRGQK
IOLsJbOBk4d6kqt9RQRD6UwyXTGs3bvXOjVZTQsw7W0afppgpXduh0FnIrV/szR7+OYc9+eqh0Df
XCdNV7aBaJXajkOi8XR6SrWTqkeRuIB3lf0ONj1HEa0OrsZEG3MQ/+OdMHvCuzyCcoJxVeRJDsYd
9DCJ+GRMaD5kKCL20XQWIO0j1AcztH0oD6xDppH29vtlf/V/WfmwdcVxs9Lsfw4bYpl055NydMVi
hH3s1Y+/jXOWlrKY/fhuoaMYMblHCDjv/zLp8FEcM6HeMGve1lhZ6QHTj7zksKU4XJpE4zQkhxn4
ktZTalmjZOO8QbC30OdZmBZQmxPhxB/tfYU39DVxNdJwCB9tXh4Q+UvGxHsAhZ+SLcHGHFVvFy52
AnXRjEPipxZ9d7f2a8ijRSbwon6EK4+p+7mCUWn2ubMUYkMmC0GzQwUu9hUKKiCO5npKS4odlqPO
++DZ24+Sqmh0BcwcNPIPzsXktwIZpMaLi78rpVc6QWvWCkvcghxnjoS7+S06zdtrJVKR3idyyKv2
WZ9LkBMY8PWfrK++fEehuZs2PaOE1wqMcYdeMQar4BoME21JDdnSe+p+SYxXagotmT2auOXHgVFU
NkrGgqW+Kf8Iu4QMSLxAX6tR+jLetLX79YL9kPHM5m1Q5Ts8uA9JAvP3ilsuXfLz9PHJH3acTbjV
cSTri6djHDk1WFzRN/Svsy5FC2wUddGQw68/kSgpUg8gHhpg62slV4HOjMSFryve+9yyOQYe13YZ
CdUt+93hdLOWqek1cTi+hXA67qwCq4A/qMA48uM3I9VKXmMlimHyTMEvReycTd6XxH9+JaxhR1An
PevcNkSwAQhBCJ8uM4sbo3bFo23PIxfW+54LpUQTFus6TlSNiwt83NkP3XEOdPDlBRy0EjwB+as8
eafkMiFMIxiF+qpJ0l/XChQAqeT1PbmFbKl1PkpYM3jaOlJAwKgGn2Yzg6WadabhjXOj+JUXwXY8
LbsKovHJyjxQqgWNXohaWVNgSxMl+xFdD+UJdKiI0HEKnnxbSBy9bmr6OB9RKJyH9aYnqT3IVn2v
W25pbzW5xtY06djHkF6U9RMaUQ9ftVAuUpGWjNbRzbfFwrHpQ3slbEWNXnYOyn2U/GS5a67u4nan
frnN4hddRDW4wXdFFFvBgNc3zp+RznP+Jj0GfCN+/qsyb5Yp/+r423RRlvkGZ2v+ODPyD4MiktYF
51cNL9WtT6wCS0rDi85+ts+WhSsLan+DE512BYSOGJ0ozuQv2zt/kh2Tqjun2wOWPqYVIHh/DE0b
wYWwXhsEW0IV/p8HFuShRk2VHHc6dtIvoqK5vKGp3D5TBpveezmopE9EENoW0LPIHDoJcwHUUcYE
OLUhXNQW6IQ+WN03+WSUlctDfpmahPhV4FGAKIRyel02NM9zoAGGeBcJKWU1SOC1gRu6mucN/Hta
V5wS7DWUL8DgOBUca9cDMnVEXm2KOZ/0fPs7B3+vWtgk5GD0Np5xxayaVpeh47vsxfgiF7H/fMG7
JJLaGWeUziATqhdlRkakXBM9v11eTGfoOyUEKdQP8nuRJdEObvjloVLvdb4zxDa7CEY07g6qYyC/
CXasvEZcCi8xhYcZJ/Y5qnxv1klw9VqsB9ewHi1mF/HzSM4hRTsLjmXYAhG8QULIyGMoiMXi5YgR
fX47qdtrJhfJHAsk+XNymgVOHtqmAVHOE9l4uvTCWbmnT1UdJOV46d+tkDiH1KnrGV/wo/IjvcDz
pTfyq3qbxpu8jiO3to0Yvr0nTNZnw352omspR91BgFsZv3+gQSeA4SLUlb/6u7e2OP5BPIrSESlL
vQ1E8tg1KU7z9mB1N51pixlcSxj6HDnek6cSMKg7dpdbNbTzQ3S+1yjf8iwlZcICY9EpISIOyQi+
r3qaAnarLn7cP+Tl7P7T2OGuR9C+LSO6nNpD9Gf0RvuAJgLXWayoAbVsyV+yffuHM83l8VcWHlL9
dDokDaKP22S/5fzoV/Vv9viFPqGGRQuCdlOkM6ly2+80SUCP8dqUfizARLwqmSHEI6ztxVl8VKK0
N70ZUnZ9MCC8dkmpJFeRXQtyRHd3uRkim3ny1OWK8pHXLxT45P2lW4ZBGcNpPwlkBKLarEe6Zl27
jRfyUBJto1VkBFzimNE266q7fcSIuNTffBaKN8HCrZNSJ5m8rrWeBUIHYcEgzZSImuxwD9+jpHht
IB4d3XU7iYQuFTeLEmjvh16sGH1wlVUmaDSqARprb4ZAXCUiyqotORV7h8f3WeDHjKC4nPIpj/E2
saoi5g7jP19YuM/CTrkebYcFGzMFzu2LCE3G9gKvPJ2f4im7IVD6TOBaiTg0Uynjf6EearcdbCtj
BbyP06Cueq9dUVo4m70Opbp6TIQ3CEc3ORIhcA17XZbmYHFEWCmGg1YEelBc/Bs0MaPHA4qB/T0s
aZxV7n/NkSpX5kwQQAzEkUuodW3jLlpsuWI2Giy3I3IyHmvGADf6Q3X+15S+6vXTRgqfMvyLHByV
LN8ev0dVy6CcEr6+WjMuwSFtSl6SQ+DjuRYRgw7+OtK64UM/leszlcgvkFbbc+1w2f8SDRZgoyp6
UyfVgNyMqne5WDHje7lkh6vi3o7dKWG5eCoOuN6BOu5/ez/YYQE4MZw3GGzkOqER6/XI+84SoAK0
2FxCcZ+TfdFwBbP/FOL0BhZISUXSxWDUlb91btzXRnn53kR6FzoOt6ClSiS99M8twtedJy108mBB
YpW7IbRFJwGG2otvsVixVG0BzdlExitaSn4jwV6GSCsGkY4r4T5tQbK5cCrYvxofO6/CD1+sb1oP
GjP4mbTTMu6vlbdS8px524WuWOXinfd+qGFF29/PmaxGLr36EzjUP5mz9lJNzVeQPAW3pB0RRIkP
ln+WkneRyMpxQYV3GBX0wHBcgcCc8kDkH87wj5VKSrKLlfq25yWHJISVv6bpMVc6ofkpD7UOiQ+h
CARiIju9jov1BoHhFsSk0nmP+m9i4tYQi7A7hZIyfwtbpThLzoWB7nRQGs4XhkYAyr2RpiLY+KhG
BTaST4NcNEWWJ9Iuo4B15FbJXqfbevVRNA/xOmska9hx1T3hJtqzE90J70ePTe8731jkZP9+rJpR
IHLDnlJq/llS3R2bfPXnB+3sS6J43JOnRvjfMM7v6qzOAb/fynAJ8Nb/KwMhrUyhyoLJMyHKmubl
+5h1Wl8/tTsORJxnbFSZjKtbXJKCsL3BPaczIWNTyj0nws7frzZ3don/Je/8+nj5eepefm/WvuLP
A4cEfySEOBZXUAhCA9Gf1J/fqBsfiIl6M3IrxMdSRdHT2GHnT2S+H5th5oD0Y6MumaANFx/pQu3d
LV/gvXJIW2yrbm9Xnnrg5SS6M2ZGD+TZjoeAryJ/JRbYNo9d/GaW2D6kM9A3qilXz/1pTagj1d8t
x4LS6zJBui5ae9VOgAX//dEMCIEJ0Yq/tY2ODes93gjTE8PIfkOx0ybuLMagbqwJm8przIe0OXew
wocohP9AeXGhcdxpq5GUmz2LvLZ4CEUe0w7bgmLeLAPo/fuxJ6UlePyxtFayCTmjRICSzeI+G1u6
DxmWsTswtH2Kun/cY03KqhGfMbEUXf0JwUDa+5EPltsjLPNo+cLPnPFXPwYVl6nTO5dwY2fGDPE9
s1orHX842yEHaWBFNEuVcfKp40MkvdyKSVuLL9+90lzacBMXbBLLoOyfFIlqWexmqosQOEu4XCH7
I2uKzXnTLIdQmxh615jx4S07n+WklclP0yjmnozFa2o3An98fMotnjHPq5v+9rXaPCrpmw/X8khY
NKzMLkIKhSNWysFFpAkGILuDn2bgkicDxLfalL+gip7UKEfZVtTdATAXMbkUxYpF1e6yAaE00NZq
xg97EXfMKtHKUo7CjoUwfmxobun+ADNTY+VaA+tT161Uu/o7/RQeBpAcbkrVL82C/Zj0Eqto0vvG
dG8zjKaD8MhSBr5jxIanynR7cWDjXe0tiMINkRl8Y+QU1nL4Xg56ovN8OS3gi12ZJo57XfIGqlyl
57FzI4pnR4wyEr9hMzqp/3S7mOt4gm3pP39YV/WNgxtJopzZtgvkeeEdNX89MxggOy5hz8SE+epW
h6HM/DuUHK9FCLdcm+2iuz30JaIYn+2xoIN55SfPaeqGwcuHoB5ips+0gVAhHOTUXVE57Xi+9MA4
8mEi/QmAYfbIWyzq3Af+ZLVK+ive9jZEL3TXbesNHedGMqBZ7tsyrHqYrlB/kyXubTVyFSXpHc0R
8K+SBvKU314EVh6F/zCJx3oGQuklMBRh3CqqVXWEtn7dLrhaug62KXnBxR0J9GGEzJkl1R0SMhZg
kt5fBTYYCc73KR/ihOeOuY0SbPNFiTePRruygNXsFecWgOv81VkGq79UpzKpH61PoqKoN8zNs5KQ
IbG3LK5N0taWxTPCaUBR0EEuUG3BJEcglo+T657LzIm1AH0784zRFUtXWvkOgHqj7CCXEPhF0VNv
72VDWWeUWKyCGp5RzsA3Bpn2Y7HEM9MW2gCFeEcFpxGJIa2UVFr6Mm+eVdRnUNed2aSgnqpaYjLT
lso845c3flXqjdnD7ngCVt1leYGHITPfYWb5YdJH3/ghu1B19LKC7TXCL6BaE1GjQP5QDzy1XsYN
wa4FaMGzkGyCsGvc2M2VR2/xsvi75UnZxjFEY3/egXIk5BGfJQLEDLacuAPyEE5cHaaVBCXJf2Uc
5qiwm4/X0l2w2b8aZ8v36ZZlmU+uyEG/Su9DPZ6n6XXs2zM0+PzmhMS17dB9X9+ZyOXR2++k1Wux
8lUH5vlqjjcuvszZWULyT476ctGYxE2SJq4fi3DeENyr6iu+hlB+N1T3+zCXwH6z6Lx92ihCBdVJ
taKJMU6WcY8vFfAAETo+2aYn9mVm0EzhTuxmLecg0A7+QAH6OPvKh5wG7Qxn4B8Netr3f/X0RCVi
4tCYgHg9tn6u/2AongfuPf8Raw3IBgG7H1dGVksv5qcj5HqxrM+2dZONBZvIjouEzjrxdJ+zRppe
R9XF2GfGv16xOpOrGyDaGvcwk9/fAhkf3IxRdL2RJ1zzyezrIhy6IdFLd0KiZPQsJnE+3U1uXzIh
9X7j4m26oMXVzOS4RoHn8DbWslkxo64izSIBGYtrvMY2cGLwoHeog6Ko33t5srT2K7SsTGjvXEiU
P6WS/ANTYwjwVffphaK2uLN0mv5aVn3gzHloUJhLOx3hPds3uBtduE8CafGbGtLAX0frd3wlnxiH
jVeQVS0iEiX5PQ6w8pju1EgaHky2/3KRPZjsMD0DGt0/dChrNs3qdmNIvEtgkmazUnv1mKMr6Mbg
MHVlHB3x+z9q2VqE6jE0Hdpvw9Pc01COn7TtyzBptlvwI9yWbtTwh8Wxc8poRfiWnwyc3HSWI2b4
Q/M/r0CNNdEFWHReK1GTybvOpqgWblA7XCUZTDEdBjnDLtt3X+KwXZLwDfA894m3B0lks/tG2Sye
TXBpr2dMIxKXv7VA9lCdgblLrKpD3Uvmmx0vdUV0XRq+Y25DDi8gXwtuECDqIfIv+6qbYLJ89L62
Zk5Q2kc41mPJ7YZzSrIJ8wA0aKldN7KJ5qIPQ5aD1bYerke7VlIZu9JojK07vTHpFYve9MySwr8X
8FPLYUzB7Us/TzDpBARYdB+3bby9L8gDQUUaMYbyBirOUgUqXwk6xyAavvSEgVNjG9VQqEWwWdqF
Q+ODn+G0e0EU3dOxEPfFtLxg8oH9T+88t6jYckFN4HEFtPjVSQSRd/Mh9BvvjPU6IpYPb+ljexFK
SON5oU/ihWhVXUDBdj9nW7CF7HZnf+6l9tiJMGYphoD9a9VssVtG0Help2nh3dwRgLN4g2X5wTTO
sNuriPTw3FhiSIuHplgO+6EomDp4m/yHxDC1a+JFDjYwXc+NNve8ATI9HARB88A7kjznU38hb4cV
GFMZzwQpJO88ZGF+lx5mi18SCgNtpr6f1PqxacF2h8iEBQjAkpOSbrdVoqSQJNTz2YULJ+zD4lHj
6lbsJownNb6OjWdprh4GTlE2zWnrLf8tJPK+HTWvn7NDPZQbFFaHHImbBrTrFTtYsNIklNQzCkKx
C3zfoU8T0d0ezWCXINOIiAR6A///Ig73n0utnW1jDqaO1SjdDEbVp9futk8kH2WSMFZmuZ+66QDs
3YsIMbJAp41LFbrqBJUJaCbluf1IFx1/pPHDFquyai0MlKdbJjbGG2Qhzar1AJ2rXYtLB+w9u8pn
j0Vx9RmwkdxkWxdif80MsALq4280gVPTDMe7FErBBUklbr+9U9Te3wgHnurkPVni+k/ZXUr/RdsX
yvni+rn4Yzv+FQub9+8cLfKXH9aMwWhzOQOdg/HgphDNlts5xeFMW5dnCGgUzkEHWHJUZkTfYkSH
UMrwfsrrfEbaiuBRkv+4p8UOnwpoSyd/+Ui7d4mgFOfI+4tzFUjvAQ4HNshxMUNePSIuaP5b01p/
W8gVlJLFWtM8gepT3tNyVOlXMrBWGCUltywmUJVNWuSEv8FCNpjtV3PKXZa2WpE56JrT30XvOrAG
205Xc506PQuajT7/cBVooNin/UTVEVIz0WwnRswMqLEfo3uHjt3uCZz3KVgqgMB2EXIpOTPR6g/n
RCZDIRa1XwO36wIM7flC6Ds1TxuPOv4zw+76907N14wPyLIcHzj8Y1EhIR5WJ3osiGXTK+w9jHbv
bAqNTbq97yeZrvM2UTCy6/nNMC+jX9k9SBDah5wJAXh28DevPpE8V7K69TI12mmWhJqra0h2lSzY
k2tdCYr5zDN1ftVGhhuwujoQFaWmr7RazNv3BR8vyYA0LbMfpMYnj1m1qodgtNjx4NsCyV/GMoK1
e18cTCchD8FS5I3Be6RFi7z0GHWm9K2gZUx4/8azvvrM5q/VxbWuLGet8LGZQc9rTa4JvP54nt3C
nvfwfhPts2lXpbPPU0NlTswgOiEZ/C2TwVDOcrDTkTHTRXfUT3UmIgzBy5ec6SuMA9NjVanyKPj2
bXFzYhgTrL8VbW5ulvH7/PWRxRK2YXLFQWI697m5UqrkUfSWtSFRd7Jj2xpbM6aJTvKPLRvlJnAf
ahQ5NXdJcj2ADIGiLCvOFlP7JaoTu9ZOvN7I9OU3+VtPARiVyvcpciC3O/7FA6LuHu+O0iUKKOa5
GIqM9kFLnZCw7bfGQrWa4BE+VpVUKMGW5ZTyXnu7pfARuGj8jt5xCyNgceWC7kB8qv6h07mkTaU8
tI0A9WirfAFVJIrw5SrpTsXD97+ArCRnXpmKecTsxY9U7kaCGZz0aXSb6c4vJFR3/zNCKQzuuTlj
adAqT1WJhQdrn89b266KWfAq7R18K5zlsOUl7g2KJoNrSsjWRFv217Wf+jSEbJbuZVJveDGAX5cD
sTFOQEMJzHWMbRlh7ef0Qbqj/70QBmfMzIfo4AmF2TjK9dQQcCnRg9APfIuEuq7edbqSZQIeVhSB
9MEZnHUHqRT1gw0JIN+WV67inUkdkELietGTKuwKYC3/tD3mvA23y5uS5Xw9uXwf7txxBWo5e/oc
UP3Tu1F6A6iKVeo4mwVAGJiaTmjo3b2ORJYFkW0wGWdereb+who9hCbVo1ojCMTZDfAtuBBaUEd5
6TiZ4YwhjISCPGloRCaOTQwnnHTKEDH3TAyIo/ovZADa3ZNi5N8kgQP/sLqhXduQwtWvxFlmWShn
voJDp3TPOqfxT+KZ5Vp/mEkidSZ8DM4/LhaZhGwuxGDNpLsCRerrWC6gR+qBT0bCzRPSLpEkyHwl
TvOGdmBM2TfR98Bh91w7557GOwqNsC2jBUWeDOf7CUxl/AHa/dyVjwoixZwfydgxISiwPkRajjO/
Ga90tc8fOCFapfFfzfA6+2txlIXY7tc02y/6Wf4qOZTdglpmjsgLMgBWQl5zKx0NtdIFoKx8T06l
9fKpeTw9ShxafmkvrnRzSoYwkqN1DM1Vffpio07WL+A9T7UkFSPnHdIooUGlRWqE9f63hluCu6KK
om2t3L7FTcCWkCuu2Y24BVH/gXXPyq47muIQ9F0Ukyz82Tt9+pEK/xfsfeNIL7rJl5S/+mXpoJp5
iZ8au07kArrDpaNy+Zweu3h59x3L21aGpzGFhttA2q8oDHdyMDg+bu71tAlCL2fmMcEbd7VLhwtD
v/TqIoTOPEAd/tUnV+RH5GDlaYSfrvObKY8Goug4+PgsqUQsRBghXisR83eLDGMfXNEy2P7BMRWR
NRYFC1ph0MyuFSKfjNXVvUCJOkJiRZoFmA203O0YPH1Omfb+2q10D3985Pgdi5cyRpQO8ywTnSuV
8tFII+K6eVdIlbDdOtlWoU7QR1dsl+z5aVfprhrwBX+w4HoSZpR63rRTO4dIrSnv7z4ydNcvqfiz
r/so32zy2dPN7dUynwIYdkg9xEOvnE3LmIeLl8lZ1e4j3jrRzLhO2JMv4JkA/dYycFHOVTOtePJ7
t3KYdPe6pREPT8XctFE0jvLqUb4WQVg3ay95VTSiOu1WcgXvMsNCcxQWbp7ww6lGv2UeWNVbH9ls
wuiFVGZQihAoytiKQklpjKnJtdmxNg1HPdG/sTUq/poTOdkb5KStwYJ+dmwRDdp+hHffguMEhEj9
yFgkp3SldX7hb1UsR7bNPTTyfk/jHkvcnbn2MZ4Yoy6Nqp6AhOPGqEdN52C3vHpkpOAgWmi4Fypw
djClXu85ZIDm6WzKMNxkQ72oVaAAnwcpX522pIhb3P0YN0PiTLm7IJMGkifLXbgvbbD14N4Okjy0
+FLgKaS//4Lzq+uH2w6wtsj2Iv364MBdIZawd3WI3rYMCfKFsPFFZ2BNe1tjIG1vvehWayNvwrve
fHQVlMNGMJ4J8wIPxgAgDCkCT1AA9ru0IiPYGhXQe9oBhkyc4cjuzRgCJtvIW5hi6y0f0lrGNlqj
dgOOBFn2obSCpDJEBzpIFsMOnnX1A3AV4D8VWdvyz+SNCMLRRAZ97ctYW4bv6uCh3X+i3Go8zrxc
qEewBgOXA+Zlh+jTZo77VDYQWFYBSQgklmGZxzLbvx5jI1EOPeO+2F546nhuCiaYW+CyURoucebS
LkWVECzdYoYVoH4PBsy1FK1Vttq/9F4zXHPuZKAkVtmvzNASpj2w3VMyOwm/R84VNiaBdZ0+eUhQ
CckUI1vciZwXdeJMdGKZBcOmmCHkguVUfIli5X7wlRAuSNpiIUUU9BQ3YFptvYWl5I7epVrTr4F7
sDqM7xPiM/jsoPLXNUlu5g+yfv85iFkJ5Ydmz38fOzxbeDhIBzhoNmhK4y1s4MIi15lZOL98pmUk
NH99B4tD/9Wb02G1dFXOf3bkUyREF5f7fgh09CyBEiQj8q9LCrun0NdkKhRuGSmj2DjOK3tSLAYb
asMfeuM3jimVeF4AIsQlxBcwjiIlpxqfvAiM7coBlk/87/KrXCdyAhtRnWhcd7WH7Wt+v/+GESJW
QxCAlLIOqTIls7DikNPJ6i9jjs7xXV05OhEQofAZHltVA44hB9R4PZVwuONrojjwbV2qaFlFVC5X
3TBGgjGBk5GQwrJWdcgtDi+xexz3VOOmlYOWfrXSQN67I/URGQjtO/ftQWd6XW3zO+h1bq+RBrw+
djida5DRr/rMfbyoA0CVFnHeYJP5rNXm6SYnJsyRUNwHKAk/40eyRq+3NJaDiHaskHMwXy01jAsr
Y3QOGU1m6XnIX7JplVaczQvwwb8JEE4GhGj1+UZDHe0nE9UbDnZCaaa5gSsHngHQGiZXPcXX+qOY
ZOoAq50TijU48g6FX4SrTrWG86SlOeDiqGA8MWv8I0GAiOFJCiGCAVs54QJM6x06mfPJxxVxqr9V
Zt8K3Evv/egnxKYvYF4dR2hGUW5FlUZJlKLzeyqpWrDOxgGwqvPHR2bSUtHlqZvDnXMdZ6oS0Bs5
vQv67o7UoWAVj21mJ+lL8Fn2mDDUuJsQEXSGMZjjvelowSFDkST9aamETS5eP634caJ2lh9qpac2
RVjWU0w/9QfHyHeATgAk1wtlrl+D17VQ9we4RL6i6RIDxkW/8ENbpfVNEIKEHs9rdwwmidwOwFyf
hupK8m2Y+wjUKswalQAyL8mlXdbrYIZ3dVkruZco1qgz3xBYgtWrqQAX7VL6bhILpwq6HZY6s3Jm
aj/58MSOEVFLwg8AfLjknxuAbXbKAimcB+wimybblMZLZPPQbT79xNuyi/htiQ/ko+iPy6xqZweP
CE21bWJIennIcwgNYJjYeADN0gXlHyoCmhY4INRk/9FYUecfWlZ3C7DghYdr5m64tMM+OuUFb9v5
7rZNGTLco+9AjMY8d7TqqsJA5YeGBgy3EWNz5dpYpsgi9YQd92KehhJ+EULRXseIgsXMDzCtu8o5
f9BLC3ISeOf643t5aiwQOKl2PjH+cby0aoLgiaUVMk7veVM853DVWRU8inwZY1rROD/H15F8ij4V
rRZKzEJUsZVZ7cMCAMfVaxL9SLs+X6Dw8SmajTFJUNzQttrvleQ4L0ow847Z92CYvZxsqPJWYdmC
/cqTsvIasG9NjZxDalwDZ9/SdycavhpxNVjK4km/5FDrFDbYHg1pHUvNGLk1ov0zKqZWdDf8kB5o
61AKu905G9DUioSBOkaLP+1lYOwDW/Cp7kcpWT/yIqwMaOEhiZrjVwO4SOH8VLevzX0nHrWRRkKN
khBt0QN24+sKiZ5dyRn1S05SEBTfQPtbrRjZL883wmZVr8bP3KY0UQizgut/XwuHpQnnI5H9crAG
2oFFqDEJDZPDNuvV7mqdkbogaQSgkl3k5pRKW1DvgEATg8SLKb3Awm4rwKrH4La3jr0m8uL9PbZ2
7II96YycemceDtYIK4InilLOYNDEuWDxSkYOtojYHeU6gwK11rtG/PPPzCPp+ovqK7TUhzlk2/KY
I1NDxwZyvEJegz4rpENOVxdFdiX4k7bWCWqPDtvrUlAg9XUJcoBsl55mp5n/hzquo6YNei3dTjhA
Sq+Yy7mRDm7vSfsHmYmQOPpbiKqfWOjjCGRHdhT0EsFxx3Ysyg2y1PMEZgad+r2KRhtPQ0Q7PTlT
p32y9K0QnNdZtiCBgmSTfJo5m+bcT/2jWvKS4wDyXxF/dICdgLNh+raXG5H1d+cL6cgarDzjCLDM
tBh+xWvfVUIewOwVTK1+ypCaJTzGqSbby+uBTAGw8Jz45NIKVTEqUHoLlOPbfIKR1ofTwQv6tCTj
v0J5nxc0qBMtodRqZPpLcSVzg9+MGjzwgo9lAdK/+5cD8I4O4M0OtAV4G+ZRNRqX2vIzBc2mk5UM
7TZOSGCHg2GjI4KxVGALaZJMGh6whOLDUPq0fyOcuEgNHHpKSbH0pH84gjYqmMq7lry2ubBxpmtY
1eUvPkiVzkexJ8o7Nnvb+Hf2ar4XPJvDVo66DfR08TZVcJKc8gxtXK0mMlxQRD0FlRUITnCDUn0k
UoSprWiieGTqwDqh547UtyB86E6AYP55xA/Ya7MqMSBG62pWXrQ10uwYHPySovSaR2+Ivr3hTpGo
F4aoRqDXxzHPiqrW710hs1FNUnC9l6nAigsF9mG5j8qJMXbqIo1i1VpsBsAusNeG7dE0bw0mSu2G
hX7OpNDWU3kntBKw/pusKJ6ZcL7+8RSUoCHDuntr4cBd5K5a4Tz86gf6RdeQ5k0RyNVK/SDHMvho
kl/Np0Yr5zR1mG0grcuYsOrlpMY3nFSy4+1c98EvWsbzagz09ziI3t4WfIm+vT3BF/ZQFlgiG8Rc
GJbLRGT/a4ChihxvWvcWNcjIHTfIr+cv94ofq/+QqCQY9kdkxd/rD8xK5lBdjoi6zRgVm0GEooyw
sPS3ZhAba6WpAfkj4jjEOryH4Fef9qFSy1BDwg6AJ461Udk2vrT1ljJyDVhR97ZzBz52w7XWkl0J
wf8tRR4bEjdo8t2hvlPWtq2MUlNb3ehR2hLm17moIzdW2GbHcabhhlQeLJitYHtEp2uvsdFeA6Nq
d2Vm0uCnM/+zulFdorfYquJ/N7xjZVGIO0LdiMlAKiWBkg2yuyUch2Wd8MsPz1M8T7QjAgPkgLl1
as3V0mNwZ42aEiEyMj/l7txNMAPDu1NDF9ACO5c8LyKddrrvzeL0QNn2zwlWyPsJh88ia9+Pi1eb
6J9+CpzDvxOiOZHGvJQdylcWnzEKCNFdEhouQ4HKujjhz0D8ja2aJjOnqi1vA3x/3wumo3ed7vvq
oobqzSZozewM25CH2wxEOHGyHrzGWzUTHyu7rfeG30K6wPt8lzU6Ft3VSADG+wDHegNEmGNEzwH9
Jf9Wm+ZtYsM5YGOEJnqRhAfCnyeB0wz67OC5FisPpA/5GQy17ySWKCCpuNhZrIisdwYtH76ICuYU
+2tcnljQJGuAv6Mcnppg0/Vb+uaOHkCbiSmT9lnOGBHI2YG+mLd08u/dYCpz/eWXjGutddwvK/Et
Jealb6akPczR8yqmKxjpOJrGjN9nOEeMCX17F1YjfrOXuTa3UgGFeutAbg5tgnR9Zp6VyWwdrJpM
c2tPXow5Dy23AmgoMj0vTla6xxmuRycHlM/Sz76D6XW9MghbHgq+mgoZFjlkXrkhgElCurw+l3y1
RAfYdnvnkF1IuXhoCD5MRwt4KAKV5x6TcnyW7Adj+odV7te/jhZdD6NFSUD7O3Z9yeVAIXDmzDQI
g8pWvdpnjiDx26drpKxDbcMBADlJ0wBir1qpHBnPJ99uvopwgn5VD6lRYeJqvpodDkBHwhw7F+bH
Pt3gk011enSCsMBOsRhpwBjJKDF76JNnf7hx7C0oOxr9/DEhcyIJaesP+Cs5zQB2lbBFMBXRXhAw
SToMlxJ8UjqVyPGsxEGeZgH4d1TzBkFRaiJ6mpmVrp/pZocFWAIPKeaqTRBQSDDnCYIEA6JmIeSy
/Wv7lGJsM8RdoFLhs3HwtvP/4NCT7eG3lU4y6kNAWTeGdKSIpV0zPzCA28Ob6AsjgKRJ9qp/6kfJ
w5zEuHXrsP2tRtAq0L6vUpAEFufmqA2/0Hk+I85fPG9/BmCqo2/KbquO9+p0gNIHw0iD5gYD8LIz
BU5DUlgoRZY9uCGTwnPwI4jFLhSQQyRBZcz3b5/jxb9PDypf4AmloGCClcKXQtOlG/013F6X9qe2
pHzoA4IXlfQs9sJ/L1m8Hf11+tfIrH3jYgFj4uemal3mTk+CSyC5TQ6/7wU4xfxCR1EiWOOWwrU7
yyJJ6L4e7p6fnRACC4bR6Io4lxD4Ga9OcpN4F8EcSDQwSunnWrW8fUkvC/bqOn30hqQvSBc9RN2s
DGvrDr/d1QPlKlrrfCBi70nzId1PxRpLxkBDADQ2HvO25Bx3sWKdJNET9RNfOPpwxqJU8QnHC6cC
RYFbbSsa2c+RXvTcrE8sawdRjjLSUfVHBUrf5AwpbuiW1X8hOP5Fsrh1wad/aA98y80xYCvAJqC0
NXA6z5lN9Mqw1cTmrXCuc+U2kwWtnYgUQnWoZOTFz/cGQOkkjFXPH+ZIGDVzB35Owt8CRu174fuM
ev2sOzZ/Y/z7e+v5e/MEa/O5mZPy8/mKRDzJhti9sFHrtYvPa1S8x+wDX8LFQ5LsXQUEatUUx49L
INHgy2jKGh6lEDpIaNRw/eQWUcIt7nQ7X/B7c9Ra3Mg1TM6/jZvB2uDJDAG8F87SGnM5RRDRGl3a
ZO9+I1BrLb8AEi3bfbXQxBNQnaWcLF2gQcyf16AvGaP4sH9mT4y1/IYHEqIu07rRsjcwGtf5EIz4
0qaBDUSwoFAviYB7umjGYNS8MYMhc4KTE6TjezuoJgYRld/zGBBqCtwK7PWYMLu6BvtT89EtUplh
lNCVXg2+VVwP3Y9ZRSqWIdVhzlXyuFGm4LXrvvZ421ZyKgw35kK4ZMebIQDnhu8/nToKKm1wdftW
2IY2xmjf+1OENzxeIq7buKcxxbE5C+ZmT1+VlDdk0zfGi4AtwtptzJLz0n/bU5TppT4pCAqlO1Jv
8K9hDUo5Yy7lTTYmV8NiA4H/47Rr2uZJARqDtWM4iPZ/LAjhFYEygKlCANjMko9i11+54HTrpSdn
tWDNXWILTkxY+JZ8rwYtnnmFOe3mhIAZKwoZlsXbDtAWQ/CLLIN9xjbpFK+jz6sYL27FU+WiIsi9
k4n2+VYNTEprkRtRN+2CTrIO93XCtfXxAzCoIoWm/V1NJ6UDLFx/jF1DUaWZ535tEhuCZ5uus6Nf
E2q/XD4cRSP2uDNJAYXlyrtukFlRkc3caQ2RGPTF4XxvbTN4x744bs8pfbqnAyfIZjKgTzCDlTC8
Jw2Txoh/oSwOUf4UF4MfWs97jnyrJGs93YAXm921Pt9DvOOLUpzDD7aofY4DvDmpiwlM+3789K5u
rrWnsPQ8sgWl/OiKDp7+YEQ4F4Kivn9ifvJDRiZ/Lq6mt84DGS4x6VWIGkE3UB9jOBmuYowLi/+Z
DnCly6fnwF6vhgIuDjVL5m539eZjW2r9H6SxQWrX4HnwcxVSc1oIRyPpHVqFI2jQJb6oKCbXQk8k
E/ARuDOx5OpxcD6OJQ5ookh2z+bDOb7pKQB0QEpQMz5b/kADFY85dr33fzEw4Fu5lIVziTEojGwz
lXLAnje0cn779QITKJqulvq697aDLFQNdfsm6N3OY1f0OAnEKd4aVJXPI+E39uWTtzYt0O5bZRj0
s4AXtvHTbtSDNdF7KZLQWKXFF0ERtkIehPX/BJ/DqedzigL9MgFXQZtRT1SYgUWcImdsBtsmEHxo
EHwc82kHDhG+UdU92LUmwIDGgUSouvQpSDcebXPeUCjUIaljvAg9tLjKk4R8gCR+rzfXFpOZnbmJ
g7HeJj6vBPpdb1zCLavyLX3eHhi9Vr9QZu4YXmiOcVlvTB24oFiR1Nc2poO4t5B2kTi0kIm6cgK2
/uYg6TXtqunF7afGCn2i+TEOqJ2v/20QWqpjrrPh8nRW8AXw4SWT/nmGU4++Cq3uYu4/NYmWM3Lq
nnf+1Ib9rqIdiAY9vjfDLUQtddE47bBE+47gWh3IACiyX/bb6APw7YeDUJJfq1cEBC/4u0h5YcRZ
7xu5Q6xUw9fKC++bGqEfZYbMMkJGZPBmq7192JaRII9Z35ahrJD73eW0rXJ6Eu6Mnp/cPDHol0Ih
n4aCRnVegCaifJrgedajtabH8C8ABjV6Yqy1hPY2tlQo1MS4ubwOECXZPTdJPUdDSkvc2SH9aBWj
lejYwja3sF/z0joei5zpLnb+zMYE8HUkxk1xqq4bWWM6nvnwPdEW1yAClFojQNJ9xQoIMhfY/T87
SgdBltA60VzoMXI9Tc1P4T9JNcx3XPd/ik25YyLFFQX5qSZGZBPFDD3Aj95hLncC27wCiQAxs5kx
VrYlyKqeBRjNiySm8ueuZCzgN+L/obu1X9S/5Rq9RukXgVbTvqsWf2FGp305TMxBvntaFMXgiDZW
LAUCBhL1HEYhthN+knf45odEGQE6A6YKrWxTyr/denJI+f10HPc/dpvPGl/mC0yUmkz+mhmihoLA
qs+Czfzws6SzY2O9nB0KWclgCF8ZxaTV5hMpeisoMbVwLwJbLmwtMrlgjpbrw6DqmWhSW0Q99Png
Nc1hpN/Vh5o7DMF1+74FrEE+V1O/DLe4XY9XrLoqlApI5yUrNemCieZ5HIvFuYvEa6o8ICewJOaM
2t7fXj7izc0ORPFiTelat/XO7RCRNDq0KHKeCXBYFSfGB1DujPgXvwxoANRxrBN9GendTAdCC62t
oub1dfNi1BB7FObUK4zqi3O+HEvdrcFTBGmPbCoLbi6q10aNirDmOepV6x/6srz3014JVWhIBr4J
qQuJBB2Lkg240S/C1SyI395vNpBGeprHSrRH+K8WdWbjNjDcor6zP1K4jCaSQ31UaFoqICvaCqxX
ou/Ka/a8GPgaI6Sh514hYm1/v2q22fCCoX6tkjwmhOtR3s4MOt3fJruTjYnspBhGHw7k5QSDM2qC
a1eTjQyGP6JoLmothms+OMIN91AdyW73pglg8DfA4I/AAu4pZYqPAL0bMA0V3ua7l9ILzCG5lCwl
22yYeawahL54cdWsXwtEIecu4kNk7WEicKPBpKweeVwEmhSW5YiDZQ1TrCap6xIZoocm85leXlAv
b6YeUinzXco6vjIQGulvfQ1U5SdBU0LDAXSjD6Slo9Td6ewBZQ3Hpl0kvbhubliDl+7XF10cee6X
eNhzwT98EWo3bHc3VqGE2pXwFRxBWwhKKg+V+TinZByVDzs7mNYQx1hvh4Nj3llkdoe01thvp+0y
H0PearZyI/s9IYnSVPyiMNyC33d71KVNDJhxPOTuQ0358vS6BzgB+JduzlJXv3euoHWudCISajzv
dl9s8HI/Tszt7cyrGW1WgbYdr4HnAIHsOxJlFPCkcRQVD1NgzR1rkv/xhsm62uRY2iFLxtPeR1uq
SoJ2sPCM23CCqo/9AhA4XN1vvYTJdFI0XO9txq067K9n3SDOgghJJ+1pZPxQ5uWXGyACwkQ/bkn6
WqygIsWDKvHRUIBuw+IYjZ2kxUaR2GVcnqLmd/GawFzn7+PiYDfSe7Aj/ZjLmX99zO+Od7csYAFy
W2ptfU5kiGO/4H7zdVwWy/JW8AGzk3JV2OSi8yVf66qUJhbkPYVJ3f6Jm+x41cpOSHjgVTJVGcWV
OJ0JKAOzosXUwNqUAnlPUE6YGNE+EgWBynGxdxSJi8hPndj74Xw1y4HxHUfntJuQRKM8p2HiiJb3
pQrSMDb/oPoEmUNO4Weugw7foPRlnll62cefutr7pAL8EEGxDIGniCmZ3WpHtDJH6UMAdFW+iJaZ
QE94jK3P3CgfE/LpiOnGCyo360g+4J6UStyItlKiSKn3wEPdeCarXA9bv66pCieXKJ5iOche0AuT
1xcp5o/p3gKVAs27IHNdOJRWmdZ5alXw3hBO0SHxgYyN6BTgNhyUs4YamzpENRWAfdwJ98PAOUtY
aHD/Rmwg1rkT6Up/NIq5l4075gMjmOo5XjicStXQRcB9DdJeGfau39OQngAlSxeC9JfAJYTU5DbH
LLZKHTSPcNqk7ahCrIsOp3/+XNciZq4Zb8/GynGhWgkn5KdHXgbH285f7ZV9bi18d+JOWoCW0AAD
1DJsRk0neU8HJFPMkmXgDYWs0fy8/aQHyEudQcMwjpgg3w1o5ohRlWySpD3THJwwlT6slqpgzzHD
oWNHNcokOL2N8wjQWuPe4kjK5qDsaxEEQgQNH2mjJbUrs+DHVLTAhhQI4xkFB7EKl20NAbNdkf+C
dSm7FnqiKNuf/y/7yATTQqpeeYD5I+B0eLs9rEINaaTDcTMfEs029yjaPGl42uBnxgvWUvKkJR5W
WeCe8o246huQCH6tgbX5iCrPeMdaIaBBt5MztAqGpCLXe6tHleoXGw5tUhlXgHrvceengLc0AZUe
hIZW5de23ubBvEjHBpEh+sj3FKJsuQnCmqireSMK0BM4+5RchN1WMb0eTebgfA44bystpypFr7E4
9ZS6gJgWDeSrHVUFavJjwoQojaBY+5qmXN9b0a5KJeWMsZ51z8WUIYHHDHkdrLMUZfwAl3ihD1Ls
vlsr8cVOrvG4C/GoELpWCJyXDeuSJTDLMiQiJqeSmWvQvpqcmalWmIDZQO15I+RDYnLyZoSZfpln
Sx8P4ma2UDrI4rvdGUFP5C9pTe/MERo13wvuDJW8PNh/yyHUA/Syw59yid1GOoBRozVrItI0TmoY
tOboPtRYsxkMjdTCwP9miz3NIUrmoHbrR3DPcftf3Jrf/CaDH9KZht/OL3yzyLpUwb2nG9DYr1cB
8RpMlNDYTa54ArgcxiRb2C3xwcZoJQZVdUmrK+FkEqZoEr808UlG/ZJUM9n2M3REfgxMgNwoQLb8
cNL6ui4URBqEQ0bOquyUhXyYibSh8MPgd8xKJaYqMEUDsk44S2tH7MLHWeBQtsrGL1yPlMyyx+p7
Dy3ifHJNEoQvqi6KmjunVh/ziPxN9rkDaHYA+gslv3z0fimUNMO7BXRSbnKI7kBbkKskEGWbad9E
yUBNvNQMXOAUrd5OVANnbNXuBaH3TNL1SCnPNaO43exJmRKcr5+o3LXvJ9Q1AvUMx+cPWBQzWKDN
gi0t6TpH4kZWqxCMhYswgXn3XPvdoMITyROvlwyHkayNSoedsc77DH7g4FyzAP6+oKBhd7Ucl/zM
65nkF2Nw+0Yii22WDUaFHHjV18mBsh4dJy7JrPHCw8+hH2jAkZXWG1m1R6LsmIPgnG2o57ZT9kE2
5vbfKD0DjSSVfXgGBJ1o2y8nyiD7zY5THzl7ZEqVOzTfhJ+R66dy65abqHHGuSGwEC1xM0uJYrAz
70AC4NvXKn7rTFdAcQ4yRfWpU3c+xnv8e6fORt2latwP875yWgiBlcQCWdXTqDXjplwxdoc6Py60
YNrwZIDMX5UshafPxLU8Nq8P/Hpwqw5iOLysRZZbUzdk76F7kzAaeJso9zRIsiTrOGghivOp9xeu
42w190AmK5/OjQKYU3Ai7boTF2bWXpI05RLkyCGGJmIfTc6yZNs3A0eFNGRD2fdrmN9TiXuIPzWu
W5Eiju5GH1KY3hjYSgx33wt4uDAKmY/h2FLH27ENziPBzS1GRkE26qdP8CH8DBjdDgHCJ7EJW/xK
lIgkn9nq+pshKMie8XxvRhZUGHyePIhR9P3C30cQ0E1SiS8WA+6sYuWiQTdUf3VKPvCBYfHWlPyE
sP3YVTCbSsedzYKDqH0DIei89UP1Vgi+Q0vnL97TdhyTeQ6Mr7ApzyCy1ur+Zh9AJhbR6P4fQUAn
gKKZv5jggfKpjBjZ5A2ALdokRY3Y2DRPYsGu0oWP5Jim6iDkbzdLIb/yMsvNKMnFeVFIFJtIFOGo
TVGaYatLGDEWWrV8z7zNfPk/YEcA5/YT6u8g93UEapyzoMlYtnX1MLRQcWXIeYgsWCZS39cOC9uA
1tbtErnsaiS/Yr9/AGQFxEbOLvRP5hr8RUVuulzUNOVgQyhi5RdczrHrY/lCEx4ZWUgL4VWbZ0u/
r/kYDp+WHhjhR2ayXX7FPBXOC/jKSo1c0KAlLjghLUs24yBsmYFpUOqQcj0Y5JqC4w89W/cC3kWT
Vm9BojSvEX8grvkyDEt+dfNMMCAq6XtssYIvl0LQ06Ravm2ZuH9Qb3Na33oqx1Yjf3iXHtutWdPr
h+e8y1GgntnBDlisD3sHH14/WgqKnrSQBHItXVaRRztGZyCvsMF0CMfQ87415FSYKDDnE4ciZbSM
fRoueeCvDhm6wigckY3S/Yi+BC0+pP+Pe6FDkU5oDkbt7EeYahpuctS2x2ttMObktEfckFhYYf/j
cLnOe+YFwNkMVd03bLkx9HaRd+/vdhYb07zTtkKkxKavjU0ap3/i3CPS0/GrCYZ3GBJBS4u8P8cV
t2cg1GgI7O5NULORFQeDvyvTnHQiPQF1q7wywyanHNcy9VMvYCJZKqhM3mFWjK9vJy71//rd8tnF
YXwpNPQt/cN5DQKNBPw7ptPmb2e0KhJpL83Hcbuasz/flOFIEKyIo7cn+nzwwMF7IdUoAGDFMY7A
lt1nABlr5oQphFSirUlw24Ep6DRnxA5SdrLyLovXpQBlGU5Lrru2t8gubDNufE1Vg+xFS2df+j7D
jNDo2saTWZjV40rvbew+44qhtjL5FsZFMz8Q3susnCPi4bXsFK7Mx7rqCr8ti1+SOHfvTgnIbICA
9IVtVzkbU7t7gXZw4sbDE1wGwIgi96RyPWnTqYH6A9CRpipz+YLGQql84bcUzqsK7UPK6oT0uFDw
2NmiugAHcNQCg9V8GXcuE+D5s5KrUVjhOIRKRJXk+yeaPt1c+F/+Odfk1HS0+Ozkxbcq30DLUUcD
42sw4uLlE2R56h2q59fwAU697U42wY8ytsQZOkB+6zylenW8uvOc1mhIftbiFwP8Qn4Zqkp13306
ram/xn+vs4QguQVWnIsGXBX4PDu/IbOKe+vDCSEPFIBcMiGx3MvwgX6casdumTslAA8Yjf+s1rKt
2KA3u3UCI0L3N0WJhaCymXK8Z5BMTE29d5+OW6tBOjOMuwOdC1s9uCFxDdmLGdxoT41Vgz4QD0hS
bciSThjmXlkOvSMpjZ5EAr12ZdKsg0X310EB52B+P3AcZYLlRF8t7iP+o9ix0sQnXtrBmj08TVOV
qaLVUUdiEeT12WusIibmtZrgyebGXC+yVf8awpID4Cwua6oBJ1LGbq3Av7XDGwX3o0QrM0m5Eto8
feeQEFhIwMRyGpqDzSC/LFedPjuBZaNmtOfv3Trj5CjV2wGbuqxPior9NqSNVXFeCieWhjva37h8
E53IqwhWOHYShl2AnhMMCAOG/nHoCZdXmtSEbr0DtHGj2m4wi6QK4XxPX3acuprA2AN+FlsW/cqe
u7mX6NH6MYelIBpIz7z8z/E80DqfW9PUc0yr/uORYSjzzhqtdrMU9vqXeHCHmwOnrVHU85eKCznB
AEqER2514CuzA/1XXT/tJr0oG9quyUSDc3kUAz/O8D+ZMsUvcWvkBziJpJiv0tP5eAU5G+EXgq94
ghdVV7D3uyeaGcOKtMt9yfJrk1e/T4wA3Ro0pM2ql4gdy8RoPx+m/rpdaqn7P/zhVyYGut6e5tRb
vUaaN1cDcfEd8d/fhiturL+jvMkdOB2UY3zsluCm8/7mt1GPJIMQGy6cd4rwn0/T7AEXvZ8Nd7Nw
S6wdPGLJP7FtT18LfF4JRAz0sp9CLQDYWW1UrnqLxqZtKWlAQYP/8CKlpRn45rbPV45etMRi9cMB
rA4ADwcVvfJn9MhoeIN6+PvnEYbkRRrP7i0FMXnkGzwkjaI7e2P3B1iSZV31XsDQeXceUJC7Q/Kp
xtiw2F9AibjXzYg0zXTU2Kiy1yFrXP2ozWBqRPZCH0JBv4+hEGB3E0H4Xo8A9Q60GE593YgPBIv1
WYTJo8dKBa6SE/sVXYuNYSnY/qcCWZqZadD2/dlsl72AQSzOJDlAebseoMkT5rDFXhlMlbAKvsrF
gdbkmEfEobvWkq9GKAghzjKQ83nV5Fvtb2iEqef45TEUyMEkHFZmMv7Y/BE64019HKWNVkUFwSzT
v/U4zMfCJ3IeaGF0H3QeO8zn6sYq6LMcFaSEWbYB0x0kTbsxDhGwyAcSaOA1QsoZPyhqrRmnIYjd
PKAIpHxVbkT6O4ZyX+YrNL2vErjK04bt13iVhLwbZleq4krLMsj2+lV8EU8kOe0aEaGVxZmkVcmM
Kx8z8lZQT0T0raZyNZOnxr7MsGbRf29/d/tqaU8JvpmzFOlZnroTHByEg6C7cMFofM5AMsfVPr72
ASFfC6c+QvyOcH0vN20okHJwOveE6zc/AZ02gwoxjIFlJ9qeqT+568KfCywv7lNNwnHQgiCx/yvH
+hXfUzj5DZELfXaO/E4a/3SMmujnat6YX4h3vaOxjo2T9ZktG+wrnbpKRToLe4YgVguK5yu97gcY
LuHRVR/rRPzV4ba8XX9vUSO3w3zPz5URkN0JyTVqAZISrLOyhv79f46zEyAIaiYUVvTsKBX8Opmb
VuDIkRSsN2ckgaO8xwAkFv6Dg50URqyHk+fs2tUKyglgpr3EKUHtQ1xxPYni5fUuWlhiZfGTspI1
9RzVrwutKy1rPBmLRppdfKOuKZfTj/k2YHcyxHgxnC3+twmPnoXkc0v8fz0tPYLMhAA/W+BTao/P
toYjMEnlPfhrRYjhkDMQPsLfgrMeCwaxBJY4BPmrnaOv+dDDi6PXu11YtKGLpHb/WE56VAtLZpQc
pB05upVjBY9UkjiKS+Xa5eHN/soAgqiVLv0OxFxiG0BUAvYipMR/tH1DnDoJt79jFq1BYoC0dCSG
b/7RolVDnFUnjqhM8EQG2Ht/sRXgLYHYGplhNY+LKpHMxwe0wD0yPxsqji9O/tTOSSmWr/fpUR1i
W3dqPp+X25k/wZZ/KLegOd4LrSOZEuJT2s4mc4gE0UY1zKMQEO+lxP4zIeP0ZgB4QmjO/fDOhL6Y
ab5ykWUBhLetqUY2XRkNKx3/M+r2STi5LMt0fT+xB1s9wLCYb4KWHMapb6SKQyfXiwJMPFn4vAcv
VqqfzFW4rCwrxlKF3jmNs9eeDShLFPDq4W0DrpyOw3tLncApF9UIhgd6dd6Z8Vx0khcrYDrLkaM1
+3QvwNZ+GPRUDnMb8L0AYrQ8iYhCX6DGcCi1BHXv+Et+24f6c+qSGGq6quJWXJTTt8KrdO3xCYI4
O/GLfnT4uZvSzYkhLp5+6vjHvxyyH7MHivuuxDIuTZe2u61k+HfU8VRAh1gCZ1zONU28lvLQ/Dpm
xWRzCT8Du4UQYL5rngXCRrFy7sFykkOuqyZUChND+viEuMosDRLK06kHr22+en0a3LuGk9DfKXyp
erX+It7bnA5dpBF4qV5r1aQbDJIHzbnlFrzdJ2nOz9Ne6wizHfbrsbvOAU//SL+vRToK8Na0CR0T
qpTXGDNBdHMdmjgvl9sy4DL2jF28N4asy8GnDJwkUUqNirMUH5H0LUu8x7MLn04/jRn9cpFOB0L8
o8XMmxgy1USBpnUfyUq/CdnGbzonRFvfeRxo04iN4W6uj3w6UW40fmSP0wFbcfFi3csgHZjt60zJ
e8XibSha3QK8kwTpbDAqqKPXzEwMpCFPiV2JVprK5vV+xHeyQSdUoCILn3arVhiw8Gzmziwpo9+X
rPEA7ZKK4slMOXwMyOG2UVW2zbcHYSkV/vtt3D/o7HmmmkqdHMOquhXflaCKxuNvHv8sYxTan6e2
SkvqE4klEW7ZDfB7x1WgKGO3HNRoM/U/Z9F/idY+WY1OV3ScsNmieYRZYs2Nvi5WkQg20udmkPLv
xgrJJ0HmA2nC3jmeIKs/jdv70Pui91SVQNYGTdcT2uWiFf6UIxWVJfa/rXUoyVtfOnBJKacLEShq
WS5XbTMAk/gwkzv33VlgssgXOM96J2M+YUqoU2QVZl1ncngp+upIHU97qHRcc2Q6/PyxMYk4Mssm
QpzbyWOC9MZEL7axTH3b18NZbVCkQnviaxcUKgI7gM6FH8U+DN7H5E5H05y9ACpOKgAYjo+V2mU+
ZnrS9rpcHyBZW+O7JOcLbpuK0JyZuDEbx9Oq/rcjiLoUXN56MmNQdR65J+mZJ/7PyyW/nIKGQNq4
L1Piks3LfEELlF76/AkVm8NVxUZXQDw5c+YFiMzG6Ad2VhsF9Ql8Y81wSAvi6PRTCAI6n3N+aPLJ
XydzN2i9mUU16l15eTmoEwUmRFj9Yn+Yytt7BYNM428QTfEsT66uW5AlSki5f9xIpSrM+02cZxOe
F91QlbwsYgde7y6VohflQCRoIzW/WCPYfLJpMmlUvqWJ3/qwnPBdc8wW2H8xGc6KYOc9D+Vbi2Ef
93Fpo7YU4NAUbCcl40X3zcOwIE91A2q/pNoaehFm2oSJB5AndTGDNSisDRqKd7V2LwgFVDqRpr4d
cyyxM9Ydra1yPu9TQFMHCZPD2WMe46JZHH1OErGSAecmt+PgZiggmZLjD2ewPpMAhKvDjI8k062a
IV0F4wbaR2W45K/Y2Y/YMHYYtcCVsZ24Po1O75uDZGWI7OjaEV52iRCXvFqsGBLvngG9Tz6J0ziA
qsEk9WZe6mgzLqHPPGFeV9WuwZUP1riUbghmFV9m7+3DO7UQzpp1KVKfW7xmNICL9S04TlQNvATo
fvcKdl5ZnLUvDb/ZMGnDfng851S51UdjTyiLsTnmSV4eE91mx2nP8nvtY3+fmt9QBmUYcLEDyl6b
DC4onRVrlaGquRvIZMGQc5Fx7ZZHs+/vrSrViDeLVryX9gsy5lTqDCS0FqoSUP1i5ryHomqU1nOk
nRpZSyEwCaRimLgqY9adYagBlDadrK3/GyMimlad6BaCgM1dVAYwvXZvlf0AQKFqsKW491oTQxi8
BP0+VHlBQxDSd0RTqSHXSH0L5xuqgEHeiWmpz5XyLOUXoWJgkNVD4Ooeaz6obgX1gxyYwxljTpex
OrIsICTWOolYqCVnndWsandj0iShsKlar4Cac5JOLYLJDoPn+Bz1u3a5zgvPKh5NG6q2+Er9lrbN
E1hhr79WBVEPphPJTDiEcrHOp7UOwb7AqNMTlu8gPf3f6+32uDkt6uLC/7dosnoXip3ebA7O5gZN
XBdSVdKDk4cntgXq2j+0k6UFlOGtKYnS6ABd1IC2YLJxC4gczz+pGPNqPfuifPNrWrt19mThwHVC
dbFDJlZLdRvuTQu/UECXDyUDVrX6VkRrYEOedkUWt7hDwxEzk/LHJVH2eaTir84/Y3ahB7GWR7Uz
Y20QLwHdWFdk0yc2boc8LjgTmxTatmrBIJ2tbPI2/DCnAbK0ldFgxXznsN1oNoJfFveZ9fWT/hsQ
EmaPtqYMI4dTD7IcBzhecq8WDG7gk2jitc/ehxFGNtndp5qZDJlwwgO2gev8uF0Sw2B14p7gp6pP
JVCM3J2N6O9ATKAIXh7+iaY+Blag/8im3WFeEeU04JjV5jQ2wI+redtBWHmr+m7oauYA517zgIw9
FfEHRdtnvdLQLCFGMc/BxRKzQtkzZPTaRLhCaeOiiOhI3hmk408Z6KNg6caJTH8jrdnMcPKeSB7U
1An8RSxDIiOGVJKZHH9ND00HAsGLXImqsVM10hk1cg2RONzMSUJfaSFAe7uf8vowZgGoxZEWCJHv
cEw+wv4jQV+Aq5Sm8ghK0ra+pIR12tQ5ISiWch8Q2/BsSYIBIskR40JiZjWmCMZ5BOROnVNjXp1+
lUHUoMZFgTmjE7QA5NFvfL2FkA0i3SG5GL5PkzAXzuoPjUlyAOUiTOAU5vXZHNu63BR1qoFaV92M
hn3c5FswGJ4O8HxnsyKExZs7Ltp5L37KI+faF+w+1VJ/F7jX941XVJ37PexphYD8GSmJUFsvK7GW
DODOmRE1Z9Gyir561IciPbU2Wrqnaeo/2wQf+rqyrky8ZrQDzuvO64e7BEtWX+FkH2nc1ElOQ9wR
DHyfSjyf3zt6njVgiP+wDgAPJ2fwYVe5FmjKEfnRJOPeMX00VFhzWrqs4ztfNAPZgbCzit7fCFur
GpbzPuWmZIeWnUphm6JTEarV2XFoF0CB7m7OlL6xwzTOvaUEOrTI4fC402sBTpi0q0xvmyPAV/vV
8l7QPcFZj1B+rW2T2WLh7la82zQZFN1TmAlDAkhLPqryEOYfa2CYT03oJrW3ea66cMXQxdYD1iPv
huzuQhosubOytotzwG6JYULobRra2EsizMdLagZyTXtqv5/k6CFRte0m71F9C8m2i2x8JDrP0vaT
EJSTLAbkadWHMGgv140MFgUkHU7DLul3wRd5ScX4hedysNiWutUNNtdVkgFb9SKOwytSIqxooAtt
HKdeOrunVNz3zg5ygGv0bQ9wqkhBTe8qZ0n+6IfrExQUs/ZirBkks7xFWpdXs5qT8JVX52jjOC6F
EB15ZURymyf+WsHRDfhZFfZ9tnRLJOO8pvUVQOBbnb7uhfnlhrhfXx/N3vi0ASyax0qb4A/Oe0P8
10JuZenHEdHqQPf1nsvv2sLH4x9N/32AHFUizgaL0ItwWQz/WpGFJkfSUrx2ybP/7zJxLxIjKD4Q
0G2jskU0+DHPJJQ/IEMSYFTFjrnRZSCRHb810bqsz+bUfECxdADSrmG3qel9ZaWH3fip54ynHJUA
WWjJJY2ih0I5RMlAIw2bO4S7YVLsWhaXlftrQA2tUal+46e9Ez636wE3TaWnO+XbdT1jSzSGDFUW
R7WtU6trI+KhDXrc6EMrciPaCosZ6ixyoomYeYS0n2O4FmE/TDZ90fyPMhOj4uTK2DajsVJGegUi
7vASzlk0yzd1bjEl/cHqOZTdJ3Fzkm9EEIIsleC1uKMb2NEvXvyCKi3QkSVfEXFa7HanelnipC8I
ptiDu5BVnW51br9iw2/V0R6TEDv8rHSLH5eentgy+tvnHxsSBfPS5/XPNGV/oDO95g8kjxiGeW8N
FAznheQdEuY+nauZWyJBWjbZY4hpSzWLzxnNMRMHMIELqEiLFkt1kxmAijcr8VNLk3JTGxPlCYrV
mHusszD6p5DGRh1qAY6qEuDMEchJye5Godu+S/Np+mxhX0IqcVJLvEIcBRDZaKNzqjbnQbjv9Dqd
BUuCaKgtnO7z+mZcf9knhSWq1+6rpnr0E3PAYFetsQ2uLL4sAyDpJ0/7MBPlU7OMOTxwsfHqtnq3
JZsZSfGYiQwz6GuPWcovYnhU8s3kiWO4pUXC5BRVSN0czlwtk8BMOhdSQ76zVKogHdH2upQKP71N
/R4VPBfiR7HzfWuqn4acLLd/hwzT/1eYtXZ3SPM+8D+/KmgFrwXd5EdTpDemN1gKb+lQ8wtCVlsv
Q962XzQrWBhgh2GO2lIH+WI/mhIoh1UKsPE3AT2VMGsLOxipNnoSLGlZMWGe6pgn5i6DjGZATIN9
wgnNVHsz5DwfI9pV/NmclfEFPbx3vl4V2hKgjfqugecSe0/LZCeQ9+SpfK2SEPEQkKtIB7T0fklx
9SWxnMvedy5e5iw+MiwZTgXbS5YLz+hH6urlytMSuoR8AaeLmWIH3dz26iV1H8OcJD7KJpLm9vkm
xzG1t/v9/mbrcLeU4/fPRlSl40DBQldJ0nFk6KQE3BPkRSEzQUafAhhw1GEzhr7TdVMBGF5nvz/N
/w7bSel5E7tp3rENaGvbHJodMme/sA5MVHntD2TANb9ik0kCSagX/zvOul6HY5ayPp31DWEH4FxD
K+4ncOP93VVOvDpO5lQaLyTQT6NnK5o8FpUmUJCukFV6U6c0pUgUanFR3vCfYa64joWs6/A138E3
H0Q0OpuR/bAPMn0zYHbpj+4w5ghFe6TYDVqi0mCKX24RI/g3JHeGl94j6HBUz8gNB8GHhHJsIwXD
yAwbpNLboVm2jmyDM3e0XYS58l75agepH/rW5IkOUejnI6U/ac8OVhhE2EqgKd5api11baRGh4Gq
MuuppZn8OEW8gSv5yZ3+uIUe6GWc0GBQQRLsXEHP1bCPWPVZZKf2nxjqCx1sqw5T4YD4CkVWs9nr
8mWrAXyG13fQ7v1nDyguRmzXc6eMMcygPpoESvL54J7uVwmDgJYzI7Qp0nW1UiwVPbybR8GH/oVF
1aubWYMuerJfHk92SEVo/AONyzQyB5DFBRJxWpb87uKKpmT9ny5+PmLaMpzmpaStWNj1tXSZPbvV
wYP6YrpqbTTDRra3HOihEnAu3TMWC9jWciJW6T1qliFCHDUOwjc9aZ6ZCmwZYu6ZeL7O1HIhNIVw
43xfW4tyWXX9QisgWBnnLouctTGzu3eHXtOBrtIcR4DPfQpqMfGAz5PcGBXeCEZhiQSPAg59PYVf
tildQFEoB5EGS7XlB7PLN/1bFK7d8GwbaF/AFJaRu0+MYZtJ+c2Vm2v6CmXdIJPAneSS/F3H79AK
zpuy2IYB90IbSrbEgGd+ySgKNCVdL5wWR3NNbvHZPoZj99jbXdsgO5GN1tYGnhXfI5dIkcVsvlZN
tGcqbqxLoS+woIXLU6nwIgc6VFG/9Iv1IcGrJxiutl57/OxhPHRVd9iezbWWSI+eRd1leP6EapBc
t5cfGosaPgMnn1K9hg+MZwhDclb6fbbGq3OsUAZXFZmsbcnWbA8AvkFCKLqUsltbLwGR6o9elOoG
iHKZK5KyE9AYTsKyhST1YdBe6p0ynVLgQX++bZNzurQpx+w0Briysd5/qaVSfWHn+ZfC3p04ac0v
63GEVZeS3efr7WqZWyEGHjUoeEAxzPlZFA6yCoZsVUuRWzLp+oKalmMuA9kqhIh+tMIdEickpZlm
Xpk4H4dDRH1kgv9eKAvyAD/PY9eMV62TGDA58GjB8DZGzMKegMDdlwGUgXvTFgsk94kB/D0lY/lI
oKoOZ5QwrS81/oS5hN9pWlaWi/oWa1Lb81DSoUxIFbn2S75gFsUj/21etS4aeusJ0GEMtis5xOg6
qUWb7zXe1Q0L2dkmnNFyRFzN0er50QMgUpjLLkMCjRIGhy7ssbH18vES4MASG91HO0A+cj0Elgjr
JcDU3HVes0G2MjZsPuzvGEEwR7LIP1TSojJ9JueDPlTnb8aO4QnXZOCmsoaePYHZMfz9EwNm+VUu
7e2b+K6F0izdc7XJ/35uY1ZBWHi7WRWYCrG1dxgH/SvYWdg+CCTg2I4v3CFNRmVI0NxVOdQBCVOi
EwG3MrzBb8sTRm7Fn/wZTgwBtjs4mx7o7xNcoFJDYaJPOn87cWXir22yWOPzD3YBKFUcSNUMT+o6
AAQlo2Oq6IFRQARJbL/5xi9aMGYFgOfD8TELmablXohaY6O91o3Bfevwx+yRJDQukQMAUOOLmuK3
I14GVszVbXr44qZ7NDeCb91c8Dm0ZuWPjFQzz+DdUJm/dd3o32CQ30LugvBgEoCbUqFCGKwygB+Y
/UwGjJvJSEThd8OrG2qdOnXnaMoVtk6oX+h3i6p40+HX1Y6O9BqIu9X2pDSx/OZkGwGsg9l8NXB5
tbPiHTh1KqovHcC+u4UewowZs7mANA5HuomiOZudc8WM7t1O1BBquBxglU5eJ8HFXW3JbkeEEoIz
zsOdUfluzaBKK/N8E+tkhAPLxHbFi8R67QbxTY4Gp+Ky3ZaLKG4VUNZHozFypTdr07ehLVAN6ID1
luKS+pn0CWc9PFoeiJHcsQnEdsFtlK3prJ75z5luXS1W4bcBlz4bPOITgXoz/Sk0F4zURsrT+9xc
95V6FmyjWugKKjMYDi9okIICO3nfMavdS/I6ZUtc6jCHBlcWwdNW3LSS8CHL2d6f94iqIiVFYt14
C07alfe5HFvYanZWlEzKsv5F2Agj9Db5cSks6SIuaHySTyBs7Vjyuov7NxynIv78Bi8015B1g4QZ
0vHTdH4Y3vzqBOuCsSF6iUorM1rLHtW7y4QHnE0ZUu6IEJazYoml/m82W/0LMzivTX0YQaOaF5t9
zA3U1NpHvK9COu7beGxstS0NNdnd8pjwx3TpzQTaB8VGqnyECq3vQm8Uxr0YmmdX6e6shHeVw0Rv
U2aKKO9XBaUgj9aMSFqPWxyX4MTL39W318HAmqBWSEwVMINCpyh0kYVzYhhE5ZLjgmbTSwVhkscF
qyC/A1l/8xt2CZxh6Rsz8VYWKQ2imYnKpiVpVUXryNSstUoksmDnzDRqcMW51GJ6rpx01NjNaZeA
TJ2YXmpghNpU5WecvnFrM4h2rVXKVDl2GnkTWXOzcS4dnYVNJdbwAdhIPcYn7aJu/ZK6acxgOVPw
MFA2u1jKMpfJcpCZz0kuw3Ph9m67e7iKA813VPZ2pmJ+4eB1NgwvnTJQKxsm6tnBaRO0ayptVPbN
sHDkfTVGzb5m/vLZkfooNakuwxOksazpcI3JPtA/xSGlB2nc/MCnxViwnbH+2GYzLTx6fqa9WlKZ
EHOCuAX16dCmSY0IQm/K6I3mV8uC2BpVlRM/Z/QBuutoAC5IwcYyHwhvIZY2zwa3TQeaNmOzkSBQ
r78vf80kLjQWsRgBaWIxYyCCmPfOSbNa2XCTaiwEZQUbVMPuJxBxPPerK68OOIEEsj81WN388h+1
B6EoMkIlfkY50fSsm1O5sY/Rji7p5I93GtnpdOhbSWq9DqNitk69nhTGhf1J6azVeQecj2+Bt02B
OmDjmLiy+u/RtWXra7SBE3kZQz/jMXhFPzmKHj4CbgxxM9zl0SOiqhaUe2iwgUZ3Qofi950R7nE+
GMf1nRNvhKbYxz+fSC5fn3RWPgAR3WqkDuUiFojNJQDCzgqrJRoYauAN1uU8zML9vcAmDGuzSdG9
Gk9fCXsM3WA713c+lEfCuKsWAUkBXKhbw9RNffB/S9UVYuNQ5oSk6xVAzT7h99Fnq/cycKbl42fi
u2afDTcsdUN02KtkJSdnwsbCnNsnnotKVlx3tOwFAY2lCvLtZUQRVeGCu7j/kDDebL7k2kcnKmKp
XbouuEVJHF9h09Ale24gSXqHeGXfD+QRar668R8luvc/v/Bk+MSxZNgjaOw/CcQ8UB0H8dy3pOh5
5i6uE4EDLk1sYQlr1f6IEcvXOXe0HfNyNdveyb8DSXZfSmlhKR9ESAWJX2inVxi0+gFPhmxR8ee4
Uf4827BNtwixJuqfnJ1/cETJA8zPAcZ3OB3nc+U8DlwwXKNyxcEtW89xUzVwBDDkxaU2iqSoj/qP
nPlvpzRKD4WrGqq+ENOGBoGPFMyk89JGY0JojI4Dx6AippyYC4d9yShxuowQOghsmX4VVJ7EEmSu
gMohx41MJ7KzR+7Fjfk02caQQiv5m3JrGpKlyv2OP3RWwR9ei3uvBFsGeoffqxssYc8rQj3yLlj2
gPnjfXhZ4y51V2YMQ4D5frZZlBR45E+MytGFpVIwTjqqIveFM5lQ8iyVODMCL0Y5v977XdcDsINZ
PfySd1KBzumDIKfnLsuQKV2/IEnQ3Jh9JAYr6O/ww302c7I4a3EwUGtBuU4utvt9vC+znuTwdwDH
K2HVPa4+3mhGKtYCLUMOEq9ye2eLtDH2hnHgfvKpdDml17dOpavPP2MCU9RhvAiIjYsmbKRebqMv
/xldtny2yUw6iQmxjMb7faNlLePN5pQ/unBh6jAsQtOZnbeGro3h3IIfEAEsh704UyZDijzeWGqR
Pv8LfLMON1U8L3NJ93SG3ZIqvwF41y0bv+UlpsuWueaeY6a99W7oI8nB9pmoTChV6w+KLFJ1jNhd
6FVDMMJXAdD9K3w1/8J6JZvThIs78HX0GEboFI99uwL41KnXx+GaNIOdvb4lJpFtRof4vXyHILeg
Gv1iQux3tmu8xxZvrELQ7bICbUOd/EhCCIvFqw/uKZHi7oZ+rqIpB14VS92h23AgFpI9p7mxfDrk
xgdufUMHjEGoK93KcebMvuzilXSat4hZJ4TAVZlb26fSnDzuZhrmdr6F+B5gnrKpBDwWR3ZKXFr3
F63FLxUK58PYsAUI12BcTKteofJQpWejhqXJW5nw6si+Uj29e5exNAZDaTME3JwsxidVtuvFbT+/
e7EO2IzXTiqTLOQynrxl4qFpMFVzF5N0D1RRbk4EeuGVWNXVMsPy8k4eOS1vt1Fj1XuXCz5xNuX0
ZTJARRemI73eca6T550HGOaQdxG8j6z1RKlJsBDeWpFQl3Z89nTrnWZ1tkU6C7SgYPMoHuWx+a8A
iJn2q9rWBk8A8J32Qr3tu0syEH6kd1Kwd70iUq3UjV+DiTy15gvkH7zyemEcbxUDfjOTD6Bpz/BY
t/JUxAvkp+UlTafFkQrcS8ts59VX6fddQl6c7bP+mvvNSox43dPWSE7zHw3ktxpBFf0Tf8VnaVXn
l3fN1tZGi3PF3jYh0OUd7anK+k3T1XP1o2yEWgOcBepEWFvHVKc/WJ6qlUoHZT+2UHAifJGEb+v6
5Hnxe6zt0xMDynx9ezd1aq/4nD6rEHXdc1OrqLUWq4Vji+vqsiwbR6IpEgTC2Uu7Xtgk+32Klj3f
iwOkT/HOgRX+UKpiSo4WLV++G7gGU+xBmnGDnT8yNeuRND5By3sRjVruNNpl1mtByxzbgdZwgBTF
KYKs8y8Jaw0s0g7m/9tP1N+sAh/NOONl9XMeUK6CC6hWAXHH1S9Pbhu5smWPFhz8hLj7g8Jh3OkU
sgZBjciMSLlxkaOb7Oz8VGuDh19x7Fp9kmTrht2O8uIm76Q1hRvoCgcYkKCsKwKzRCou2L5OiEXi
3710Il18p5/1Fmqz5hob62H1UZCRVLMaOZm5uArz3b/Vdxs+hMFWVTVvC0s8WOvfJBW7vuPbI+FZ
T1lHvIfR19TAFZPNIeqtQ91rSnXw5Ye2AryBnjTD4EyX+Ou4pmwyFqPIXVak+K+pYSCRAdM+XFyV
R8c5YcBU3/igNJspEtdODaXAQfDTS8izII3iCeZmaPkCKLqU2pfH0RpbK7g6fJ2QhqL0uq3bddrd
B9CC5n3WOy2DNH78Lnah5XnaiVFju8PVIk2EGs7VsjdF7VKkHeRXjca3vMQ/hNLjxYXi1Pi1/EBr
bdhSN/lNHCcL56CNeWimtldoZO1Iurs+GZ/I0p4Uks2MxUMM5XaD9aATl0chAeSguWT2jjlWPH7L
Bo2ETMzRheMLAWKvcaw7ldPA/3CJoOD52JP8Kv/1oUYtC7Ngs5FdCvreUBKL2OJokOFCdz/9Y2PA
2gHr/BevX9Vxj/d5fxlOa72uiTcMegcPT+M8uTF6zSdb7tQ9VsSw+71MnKsH7hO3gEjSebuD8T56
aQ5FiSDVck+5xqTEoUaCA2ygTrWTsE6uy/lvSqLA3UoET2BRXPAlhj927WRp0pnH2e/QhSWRH+NX
HkeCMi3Geo0LccItz2YdpO4uaLHjt+GpPihjCPgQc8DW3TfHpgHHoY+Uy2PML4odZq+w7izPsO+r
05pDX4BdpDOyGAlESVM2ru5/egK3eRgaTufSB59o8WnVUd4qdJqbFLkoAXDFmmP1FC0+T+v8/bmO
0wfuDkM1BaTxlwtcxED+LQYbive6df7P2U4doXYYGkid3Qe4XFfZ9FPMqpw5XLMcifurQ6C45kFk
nWr6L7gsEph7tyuvLoyt5wVEPE4M1DTqpusVSsHo0VZrbCtuPYsi7oMtAaHNONXkIibfbk+MqWtd
7/wth+8ejd9QrhDYh9vtVPgWYwhwGm+fw5713JOKqlS+bpMyAgYoLAFLbedXZQDViBFze3rm93vV
tCkkrQqQgTCkYXA6hnDuSFuHCy9D7XXOsBYGY35n9d0Iq+H8RhqifW2Fix76RiHz+MrEGMkuQ55w
NswgTmRCIBROV5kHOiIvnNOeJXs7s24jt7g/3UJFaKN8kfDU7SGgnj9HOx13PUZ/StXMAg3HC8Rc
81DVcfpcXkyZYco0vyUzRGHINWWxAMjiljZ4d+FE4YomkNCew1Kkrf+AMqmtlvfxjNJLU7ov74UL
7DwsHcDg/DuJMkahkH0L4rtm5rAbJAGEkHh4nBi1wa4tMF+TDfpjjfnMhhqzAZG4l7bPW5fLTtYB
JRhc8Efg1tDIvMsXCr/AOjglLHQlC/GvQ6CWli3soOeFCEDJVtRFhEVdm5NrRYLL/jbjoDwYLuvn
zhEDi4Jq46PA0BP17LZRef2ZsKfBRxki+Lm279YSOvpByKD8cQJ83RVivU86yppyOAbiFsvOVXtr
qfrYrsqM0rC5lI6jWWUov8VkDK3C9CGbMomQC5KFlcxR3/Q/DrivzcfptZP2QYi0pNHABSi9Tc4+
2/9h44i7TaN1P8LK84HbVmhvc22H3z4LbtykRTYg5KAbFKltT5QOZequ99PvHVXyE6nHzPM21jL+
eJVnUUy874gVlb9YfHpvWY2fxDq5I0MiWQT9/Fsw3ERC7if+Qpc01o8M05MaeEIiiha2IM7rb/gW
1bB6NWeAwFPtc6C9Eao8tEqRfx/HofFIzmDTsLrLYzTs+58jBSg2lEuu/G5kUraGI5GslNvRtjE6
wCcgqaRVcjYO3v3gzmFB8RTtrZASfMWtuukUCE6mJZ0vkvBYWpMvHKVTdEyvpfu1MynTMrVV5UKm
AdOl/wKFTQu6RbhZ6Gi4DjorI4jsls5VRhmYlT/DpnQbU2Mwj1M/jefGrFfF/jZnkGrh+XsOpNri
KPKRPIXgsU/3UiDKH0eBRXGYXRIr/xU6zgjEbyueMpBrAOkhhwk4lk1pWI16+Tj5sonAvJewvL+t
zvtGfIvzN6Y0XVugA3NdkHi35NUwS/MZGvGLaoLUBtQeibmDg/ibIKayJajWQIaaIkQtyFJG0uEY
9iQljtUVks+7F9rO6zB/+Gr1UmdftHqrYs84ocAeOfsIROBaSDv5mACkubYueMY1dz1EuyYVoGTw
ZPJIL/v21MiaXbaQntDG1UsK0HjJWwia+Y1/QVBh5+xbm3TddzXHfz9lUSO8ptj5p5eYO0CvblcK
My7B5dv1cwnUP9/Tl3+C7vx40cYofapdlflBGWoYFQEE1yhSg/TwdxdPnsRPPZxg1EUk3+/w40uv
jiTmHMCWvkRPMLauWJe2ztv7G9++q8D/UL4tXtN38AQbotbU6JAd7zG4aauO3SMwYr4KJH3R/oFV
0JzTNc3RuNDNajhnxUyo9sD0lro/pH6KVc7LwwehwAFeZBEM7+JxZ9CiSnS5quLKGSNfJRj/m4Dl
ECFzQgixEdheAC0VBA9skM1WJThfLKj2LIo72wimiIM6zJq0YVL7tsLJiQqK+E/QZwXIc5CqafAm
e05hblCjpzTytJBORzKw5iCNaWVZi2LrAgC9+kH//Mp+/jYL82oP2OLzArYT0bCDSdBfuWb+Pwl4
iVSxiSX3zy+w3t39bWo/WOxypsfTF431H3T8pJPDRucpEzj30wcH2I/Bo8Dh4+8uCs8/9IIkn48M
xupIP7rTZz1MlWQw3LGPIaZ5ZGKUCatsTb2ZEEbFtIb25CZS9sTrUCJ7UMJ+jcP47Bucr9MtH+Sz
kzaFx69XeJ9RU3/d2w8Krp1rE4EHEkd6P440bHPU8ABZrH3Qtz1d9HFlT2UUcYDHfcjDiILTskgL
GTYIabgB/WFLO5ZLzCTkfD2rMt9b7SRr3KwWCtOtWJnF5Zahs1cQR0dhDN3Wa7Vh8+LxG1YDqd+X
XEMM/DSE4IrV2mwIhcKXe3r4ByOximbhbyKu0KFDX3apnHdMbJPpHEcWvQSgMNNAssFF4LomgRhY
YSFXvV6TXfW2aR9lRbZu2SvO8kaqMZJXXBhjkGzseEDlOqBNr52spAHKHMgnFGF9d+C8d42r4E32
xQ65wxkanB7XCRawOFhMPCGs3sjWY5vDOZbpnDL+oycKwjX1P8c5ER9vhhjQKpkPTfdDjN88Imfq
QvwPXdll2yYM3WROpfKjngQKTO1tf1494ad0recBia6I+0MdrTdCMsRMp1cfQhDikU0RAxEYJo4q
c7TL3u9mPoUqSzpqR4u1ClXN49dLR69d+0ctFADCPB3zhmIK5LmLKdrATTWaspgEeCFM9zH+Din7
6u1Zjv3qmMN80pJU+2LVw5bE75T8buE++x3wmM8CeXax4XPcsBCJVa0zgRYzsP4x5ZyitrKGfeNS
4Pyp/6pSkB6JABCO4JJ1+DG/rSoHp6YpimOIMK6ObCuO/Hze2d342m7Z2JstkbgGV4vS2QTStGbd
CZDUYRYFXnb23BPPOT4EFtXRNc9iwo0g4emWlPA3ryf+TCKSIwPm5f7jyS4fXmzUn2J7Xcilksdw
GJuiZ8RrDPzayJGI/fskIfWLr4NNVwkKqMURyCcW9x6y+8R6FaPFqpNyJ9zX/KniW0m010zH67pu
8vCxDhZHLC14rmvqsMQZvjyG8CDiMWi2LMKsMjBYs4CVS7Q/BuDBsnlaup/d90lZLrQsx5JNvlPF
aInwoza0696LF8XqO18xL4s96a/v4vCafuDBQP9vdc42+kJdn+VAaFBlmkNgpHI5rKF0VtPJ5CIk
xDtOQ+5WONNKR4dYN09iiCDVP/WI8Zm9Ut4IRE5/ji9LP14iOo+9mxYoUaMj4tOiTRByEdNke/vp
UGqGuK5JlnmOeWHSP26G+sXmBH4Fn/1iQg2W0xQVAs+wPYkVq1F5+twE49eolbyZm0PMh4pSSIBq
EzRJniQ5XxXe+ktTTa3DfHH39Bo3UbLA89HNpYvlqhSsuRuyH6tTQAQ/5Es1HH5c45AnKpxxGu4F
lrQkmz6GIyWUOVA3DMeTFT7wurrbicNziLiEKlT8ufiEmxlHVw8Dm1qQO5qom5ZMuhnM1wTsA2yG
nC+a4DY7v9FVuVLR2fTcUkTiKXY9WRbm5qRw6pmU3tOgh8aFBfuunAaAhVyuZzRhiDMZ6bm04a2d
UXgDX53PjRW+U0PSt/jmcySc5+Ot9/reQKoxCjqvI+tTXdJb4dEqks/vaUOhEsxPwHFlZ/m70RYi
rAGBAD7e1ZwC1vMdi2RStoyw2+ezGjR0JMd0f/acR01uNh742TE3Ms5JbPTBMbZ+/K/cIgUGkA4W
TTs3QUnOSC3VqpwZYoUeFrOlSsjQ9tcuk+DAd0Ngl0qNVdB1+l6JoGAieGRfyYIh2fdCG/TZsGOi
QL34nkUP48BgjnLPUepli5ug8UTyqnJBhcVwYCOBMnPvoVMNvit0VC7ap/DJWdbQkuBPpu9FPepw
m9d7hk7LKncyG2+QsmijFlNBSp/caUamBv6c5ESemtqdYIX9NAIEW3Ou/GoXuiqElhjFNzZp+FLK
JBk2cXgra0BCkabcqSe5ILISxTFL8UwVxV/PXwcqBFg60VnT+MK9IftQl99hETviAY0tC1FNODWi
zsN6X3IINPxpG0vCpNZstgHjlPWph9HS1wTzZf5wmiPBNRK7NnaBCQTmoj01aXSB2SL2LtWjcsNx
nRJFt6A/uyiGLD7DuSyl/qWUeqafk28U8LN14SSWvgH96Z2ioBuTu5SvnOEkXTR7Xn/dnjCq1W+k
Rokp+D7CcbLGEXznoipVgJOt8REFFMc9KVNfiznQdbGY5Zal/PD4t0VXRI2sGWwAAFrgjSeNCFuI
j8HEpNlWrXdmXffYsTtJRaRZ2Cuc27KIvWcmzOCn8C8bjgUImtpOLtQmQ5895Xuv6drCVsf+iEYS
fgeC+IvNaP0JsdyHyQDiv9vH2cZNXpb3tkFuejXhdDW+th96L9+3PTzstgLMCIfZgF1RWRoVFA7e
XSlgYLeXKPRmakNsrFj58XtjxwWvMGxEnieq8YNf/W+cfQCJVcXat8ZNItBtJd6yA/HZzuZ5IGSr
wUJsC7mXTREYOSycn5O+w2agaHe+xB+iovL1DCIgffyP/mjVR4zjwvGf/6dflR6Y2BWlazQ+wA+1
38XainiyEhhOB1NI9pPHEHJ08nzXB6nqGbZcCm/A+WmBjnvSSGhRrNS+/5RVgXnsKhlOwDVexKKB
3ZMWfdazxVOfGSTjc2cqR+DnFoNlaGVP5mUpRR8NK4hvYL//5ILjkFo+rMIfjVZqNpQhTiZROMmc
btFU3ctDwuYEhA9uiBA+R+DqHF8IuAGB8BMuCcnpYRIIhtAYxfxsKMQzy5e8JQ9EeRg1awwOKDiX
naM2Xq4H2CwWMI/7T9zz42glxK9lTSqmE7fOD+ikiHWbTJ4wYZ/grt2kPIEDa6m+C/g03oCRgDOm
f20GQR7cSm/TY+B8K67UNYcHvAFFgpa+ixzgwZ3TXGd7IngGQrsWZR/9goqMuD+DUbdnXaHBEcJn
k+eUnFQhozsmsGLRZxrIm3AHaKUaFrEYadFKtrlps1UCJOTTHlhzfXWmRBAy4YIfsAeCkwXogZSh
e3w9niMQD7SJaRPN2PHDLD9zWSalXftQcvnr0duPDHDXNsvFU8kw649ri0GFCxqRY0D359R4Zpfj
l+4xvESCqm5y6TLiM1fdsMH6apkvZKUZBT10lf065uSvvnjzt+Th80tSJD6slw8C+9T0HKzlBhhZ
YZmku3jnpdYEzOWOuqd+25G1z2/i28/hqqaTrSpFlz7eZwmDVCeO2UYh/9wGGfJpt4SqMFQ2sSzC
9Z1Vt2lRCoRB5mhRJgd2vOsLnUK7KUh02dgc2K2/kVmrSRC0W0Ic2ZqcYCfztnL08jKYLzJj+tXW
o5CKfp0slDxJv9yWqpaBYtgwmYhLF79nf4Ux9ZXWFZjJ4h2FeRG4EtybxHycgh8xeiGJwxY68OSA
WMF56GpC76L/WCf8fRu8oQtBNQMM9dySMP5MbI/3MGWSG4dCKgyCNz8fKLwPpaZAdxffiXXSVawz
x/r0M8koIZbHqaPUn8xyxWjGcZE1b2kz0mdy4H8nV+kAkIKfMTW6hIi5ITdahE3k42Fdu0rLW7wX
t0EuWNdMgBl8+AZy3aLoIird/DonPzGTFG780aTkI2Vr0M7LTHkJtz7SHArD3QC1YoyFbUS1Mamp
Fk/Cw3YAZRDY2iU3ICORUbqZoNuY9YFqOKH995apeYRWQtQA+bVNsfucNtyaaXAWtvPHYHMvhn/a
lKVJhubipH+h4LnwLAly1QUZoWr3Pm/s/tNkVFJrChCXgnRQBPBsfI7A9SWkXKbZgyz2ax4MXYsf
P3X0b6IrSzIeI1PHzZwB+S2g4wfrA0m32JKd0Ql9EiAc3tJRsfMN7ljemXmqZLKJtSC2f0fsvpCj
6LEppTlqKF2WauVTIeByygGeV00XXtcfB4Aoy/aUhG/QPONN9WhfaoeLNQ3IPopoPwiWd9j7WSUe
T4+uRizsb1bY60jKtv3szr02MCCAyQ7jniM/NJjyCGm2DJjWBbDSq6IDoKKCOHcwqJpUEy1XMK2k
67PAj5LvaUZ7Vbu2HUgV1jerRWoemAPbDcc2Pdh8nF5eW7kE5bBS+mk4YQ8IKAmvQwMXvwyAXsFR
qM8CkaCcGBbq3YQRPFmtoyijhrqEbdWIdE+1WUzT+Nt+1dzQ6qrmlP3uU3mvI1pCM02g2UacC/Xt
elHXhgNG5Y4Wd5mrwnS+mCi+BQEqR6un4i2fg497RyXcsNV9GdkbGIi8ul6hsQtMrIM/cY1a4LkM
5jrLMtou5UTOcHACO1sKrAEyRH4tUy0yUWxz5i/kQ5ntn/ejIy/pzHfmqMaUL6KOw3ZnDIWV6VOT
Mlcsj8oiUxTVgNe6nNdVIYil7+AGG15e7o8E2W8IzFbxHnzwZu02mFEK3LGqNOJQ21b83cMi2itx
jFSsXdPmH+hcu2y0BhObst7egp7Ru885530exdpUzUhheYJtUg8xMF6e1dCCMRNaqBsFulnZsOwo
RBukSM0l4IDvsNCuwMZ7+yb/V2TpqanXD9Htq3KZCUQSdiJ+4Q4XxTf4a+RpPoX0nEst3cW4Y2ih
jYf6l9yiV52rRIg22WoPxk5yApFrBmGkDFD/ZoxkhLZB25MKkxx2BJw+Qj7j3E5rjj0WnwQFh88D
995bwK+fhyvh+oA6xEGDE8MetV2P7AXJfWOxFW4eUVteLk+tBVXcDguJV1m48FepG7dY4hBmoPnG
heDzk2X6it1gUEzM2VdCBU010CkYa0yUoYOBGLS7uItQHNa/ev1w28M5ROQvZ6RYDPJjpt/+1cPU
XEE+HW1IoQ3UpmFjNFqHNVZGJB7ffZisa727oI71BOQ8Q0OTkKaFyEIKdEzThwF+gPW2NdyVkrLV
V/7PjfxNtMEXYBJDTZMFTgrRRT6d2Yvj5XHycAB5gJEqwFiptGD/i1gOo/P/E0fogBwjJr+j7X18
6pGZac+1nCHAMleXFc+bREstyqpP9l703MrOjE54TRfDTZEZX1VN6cpvYTPA+dleiGbMmdmlloRG
w3DUFfAaATqBc3mzCw1cDjX7nSTn+nQK4iNiV7I2lGyMtWvk6rKJN4OvHc3rVAvtCB64n68oJms0
oKppSmBOTp/0T9y0S3C5WASTODkhK99ml9lOiSnXyw0AnqPA9R4FonU/mMoSjT4zwG9eiqSWgVH1
wI7PaUiMdJCYys6gXJqBVy8/KKlUurOSMtrwBElgk6ijRmv9Oh83QsR7k7deLTENb4d3cH1KeaMj
E/IaQTAfUdu6Le/ei+Us+gIfoq74g5rCppZa/z6VhMPmX8EDqDrGNV89HhT7tK/N6tZnoBgutV60
keEzTyzAib3LlZvd2ZhCH45kXevAZJ2kt0G4TfEFjQJtMPRBs+Gcbd3rOzNLDXm/F7Yl7+v1bM2L
J59P9utEF5vbjqDjKnLqdWxd2W2McrduL+MgNCjMns/t7DCnXw3r8rY5jX5L6q1J646AACtE0318
3BAjlGTNjB6KcNhCIMxraOVpOr6d8lMPlXMXWo1q+F6LO/ndABGeHS7J1/MATOf/EUTpYio37gE5
jjh8xKTWC6I01+7cpyhoq7IBXvqlvHe2mstrwn5RMYF8QBWhZAYFSEct8fEX9BGIz/H1jnOQFWJk
qT5mmSJVVV3RRkWJdkqLyC/9H7cFcJB4pVEHqBhuCM8Z6A1xwjckrmDm2qiy9tO2LPcnyjmfR+9B
UhhI+yA9TCW8h2hW5J8+akpNEJvM2rSWyekqIpZT7dSZazDH9TasXyy6xYLHdWZkce0BU7s9UIbi
FGG2ko94mPLHuhoJXJUyV6flTftHA3qqMB0XB3wLTOOI2Xm88hhrPnAk8w++28Fh5ySggrwxEdu3
izz6Ac55JKUbLOlJ8GwdBNx7UP0gB8rFlSnU5JZXSZrxecgDXZNU38HLhO/nbi82MpmpqBhIlZtu
4iKSQfukIEyQWJDe+LYFpimKZ1QREaoHRzoFIRjqkX8bas6l2U9RsfUUXc7E8mKt5tVxYIzoCtJU
4iDX8I8OPltQItFBR6Agg6RJLBju7w05io646jql3cVtnJgbkuKI6AxeVtlbW+TqeEYboXpgRDjg
6ZLnafHWk3LRML8YXhejp7Fh3L1z92kQK6OHhj/+k1YYyUJZjZy+AaqCZDhLs8IMKrB62Nx63ggW
mx3f8fGLNIafiUZyjFiUoGkwQHrEPISvSrx7iKIGHuIZU+/Ln8SMZPV2PUHUbGX6NsWVqGS+jTZY
HhNvnEGArQB5FazUwA+WzpN8pzM2/BS0fOAWmoodsxtnq4iGLL1Y+E+mj96+mdhZ6C9Nkesb8joR
R3+VdTyxM3OXyhNfNmaW4siQb0jXKZoovDMWYF480LTxQ5+VvV7OCvR84CRPct0FMwlqXBjIVTc5
Nzt6R/WGfSLvAjk/xK6VV23c3chEH0+t5FF2WJZ5Or76prHqWxOzaIjFz9leaMqq5/QWFJD0DxzT
f2hbIhJdSwnKWjlKZAzYRIK/f8aKbkp4aYAbFFZ9E75uIy2fduqokM8A79at5wZwy53c+8EE9LFQ
YgkfU77akYP8S4W2fcUITkRVYLDXX/9QmgFuWk260KcBv+XuqXAfywo8VILla9xRlnVtCu1qCf3n
4k92KVXiF9eEmM3bT/BzPh86um4as19FDdip5WBnSRSWfQ3ZdnACLHglz4UdKSba6FjoWkZlOozp
waNHZJdyBqJI9fqR6AwKn7dwLMsvvn8LNjHHGa24kpTxUsuL8PKEdsaKQemN/jxhhn5z/V9CNQHg
i2RdTKsETKJZiP8BcJLQNqP+uZtWVGhevxIjKxddjD+xE6TqOcbeMu5vaNOCiwCQPzhpKfXnfTRr
hfXvKIbgntT6EZg8H25QWynOFDerx3yxi/HiqX8nyEjyR8S7j+qcVdie5H4T76YaPun2IEtTCdau
lQLoVRg+xL1lpHwaxjafbWQGzEP5/i7JoZkQYe5vfP6xAgETT9T4EXsGvGVY5fTu/iPRgmYgeWJK
bNKrrLgeuqDEctuvEu4eZCel1GiWJVbXENFZCwsVPrIC6UDK7uD0VAHOZtmQHJJv0JNjcycZASjv
n4IJxXiyQifQOlns3TBMXq7P8BJZPFXPgh9MJe80UOnQ0NNJD+PYm7MkTEVmVRrNwpQo8j0b23pQ
lERJafGN+s7afCRSxpGfCypqk4IM857Iz5eaemW3qsQX+KlmU8P25Wvxe7bQnzJfccrdNh9inVdt
t7fGrb3jYm5r3pwI4z5Udr70z/MmqRoNW+PEjuSHZeFDSOmaZOO+d8O14aOHS1IZf7YT6FM+Rddq
8xngAHAlwENZxSl4dJqxQnnyXZai5adnQtPEp7s09XLU4KuUs2gI9Hdi6EyvctJGkjPFSQm7Rj8C
LOeMsUi9maTR+uJGVUfb5Q9U79/h5McbtRXjBpK4jPbHVw2Xc8MlJQiXvEIvQ3gw8wQbpAfiR8p0
fkzNeI0yAI75yjdunuzty+I+uhzXUU67/++vCrqoSvg+T+Z5yZshqf3gUVtp7I+GjMCqCSaT2cHB
01oIkME9gpBLGKXOJmKj0cWOaXw0OYRunr3eql6a2RmpzYEjvRwtuVQQdf0UBKBikXV2kiGFx6EN
YVbvnCPQGpNeuTXEkqNA/NOBFotR3rpOqotw+UVVtZObtRa1g3tPnLEZ45FhmU/aiGGqMyZK3uCF
yo8UOhJ5L8TcQpFM1Uf4w2JJPneXt2CPSrZiK5uRRmBtG9gNYUstLNJWMraD0H2xFV1wiVC+rNY9
WP34A4ehEubAtl6JOr+5v493jBfOIlnqoayFUU+AQ8YlDm1OH7Yg5qZj/MLyWyyaj0lJJYlXLAMZ
Ic7urmmErdxjipFOeqZTgAE9WRbeapAUrwVRx+Nmiz0QBZvs0EMQAQla+TZ5AymJBdd/PPKqFFZg
uWypDjgA+MeVCq5mQxLTCQpDZgaOkkI4hZLXwVdpa4DJgGvhTxti55z1tBAf5SGiPDaHiVkvZCG2
8qnyJu4FLWqA+Dx8nHEvx8+P5sRI5id4US3MHVuniXm4AGu9pGat8pQJfk7PA8ds7899HVrQy3zf
vi3ZxaM+XS8pVMUJs/qLN9LPi++o3oWreAe+HbWn27WejXntf331etokwi8CSuvDAj3p+ZMM1Cgr
d29hUDtm39P0R1tdnmct+pQZHjBCOUTiNvqL+vVaIJJd+2baYxuUWfhk+2BKNzOYi2x9wlazI0SF
SAT6ktGl0azxBGB0A4r8om4BWRG1g7ekPpQBJ5ihAaspmmIAV1Ktizfzygsh4+fzv7jpK8+eqs9N
qGe0uThOlbG0s4K5TeANp1nZddtofX5lHZdE9WrpalwkgP8q+EwBqujVTxUI5SjGJSZn1NM7cMNK
zua0A2U6PDjuCBlA4H40MICGY3kkaqxwFiLBebA5XdnpSsMILYmqQHCE+SHy3uaqRvvquHdyJ6a5
VyYDgUDubRGjUZ5pwhGb+ePIHB9dI47+hCUZdfsJoGbwepxNZuniECFfBHpSAw65gOiO0prrlmo2
OV6IDViScYiRBprezfNtryfIfn+jUuTCsaJVh1tBGOjLW+Y1eObicA//pxtQRkhER46qkKkw2mrx
94xL1mLq7kDCJHcJsMSAInFLdEuXH+ywrZiTYEuXu0P0xkn//1spRIZ50F3nDNGfyeepgRuQ1i9H
Tts63kR28Hr7TT8ogiF1SKO8GqrxWh0FctCT/5XivVCW4r7ZE6aQnztJfoZ1BcpaX9wgb6h9cG5W
E0mr6L9l8O6ZvRtIJKEEcp4yMvusJyNBQptL6DhOaWkpzHEiAZGMPbCC1gH3OkFI6d1mKaXeXaaK
3qzA3mU9YSaIk2d8mOgnOFKdlj+orhRe7vB/TLs8RxfvUAdqTwmrHFI+csIEs649Nn6hy2KjHags
F9DnKlHh/FFaQUSFjThPdL48+9rOCQJsKslmCWWzhYmC9U1KfpzNvHyd/+LIMcEOqXIwT2l2oF9j
CD/m5Rg3V6ci+oH0Mv17tAH1Hg157E8Bc9tSp9vAQAn1wH77P6qT8ZoqA/SAPbxfa509vzphpj/Q
YXjuxi6Tz9ZUCDtrTzszhTMNpuwBWH0e/J5mI1HOUIiV2Tm3sgH7nFk7XxLsrGJSKnQuCggOVEdK
bqXJMs64kzmChEmJYhxhmEYWjLp/mjPAiINuJ4PMnjDNYGH359zJ0eyTnJ6RmP+L7zYh2LhVFKkO
PtskSmdlvA77jE1vu8aUzUFoaBtg4CrsjhM6s9J93c8Ea87uD3OZTfaL0CVcyrf3LkXB6yb7F2Sv
ZAGnFXqeUt+rwBDqGMF4hJO7ggOSrau+Rqg2estHHraUYGwtkqca/uHs890WIFrD4tXJJBVeURXW
6zL9fn6s39RIPj+S9KQ4r0hSOqP8VFJG6smW/Qumbv3HILIQLhj6kC1HcKWqIJviylSr6gq26mjg
B02Wnv32mOUWY7LqLHTMMxOVq6sDgPEwf4PPlVaUUyLRhyxw5mJve+wd6MelhyJORqrCL5hAE6AR
RWyPAlQHOsddQ+yDRdcq+gWMFchYZvfbj+qKl9VPWfLHSRr3xRq2FQsNB3BEE2IH2LBkjvOb16Ri
rK0h8KaYSiYW+Mv4KqIMBb/5JRhcBq5POh09xMGeqXIUjAaRM8ZFkXZJP2TEW7/4xkkBWkmIgZ2B
ROHbhXRLzHGnc5EN36QbKfn/Hz502wEYL+H69/02sls8jjLWrLIW4AJiOOAY84jBm6LFMUfqbXJa
34lIz2Pqxsuo8BmjUX2d8A7DU/Fxz9IRbDIBIFHMMTMKDCx4NdVoW9L/7r8D2GEZunAtasMBG02+
JRrnXtMMhAYC5U4qYPZ1n+VLt5UPovbklpCWjQG2fJ6t2sClwSBAG3Bd0OCzRqFzuyezGrfYxC4z
e3KFaM9H9QSwsHDmXgXK0+mI+5GTDD7jIGeLa52FbapFQT+kc6z6qPhz/C/6J6WLHqvQBbATAPis
hHIT1v9RouoP+S12Mqy/+mBhfUR3GA53J+5n5j2y7XPEk7b8P1vP6P+QV2DJ23c8uoCrkFHaTqRt
PkgtMCOa6/uIxvG2FfHdLe4d3b/NfBVma6iZ9R5z1P5gddZafwnyKYuD2/XL/Lz956tIES21qwWF
YY2tOVL56SQFpajv2+jRRiR7cvXkDUlSMdUSS/g9SKneSqYE1r9Mm6Y9z/37oEhiHW8ihgXvzomm
8H2e+gavEQ6qcZUvuHm8eI0XQEoY3alaXDMzdPBcnn33SE+fRNkwCVrwGbYMcO0sg9fBqFlw/86j
QYZ1LymiOzU8KHN7gPpjKgeCY9SNwCUqPfP8pLNPAFCWnGjedt1JE4ablDBh3Hcsrk8Q7D1Xijv4
ZVZPjWz6YTnoI9To3w7Qwk0wjfT3t2gOXXYpaSr4VLZkq+a2l9DosygJBHlZheH0y8IjtLy4Y6ww
+9x+lAlaykAEiOCq1Edw5WujksNQg0b4LExHKlSpiFclBL5ZyVpAUL4wkR66QfjBA8dVkIgVmptu
7/dcqYXIA22oB1JC+HONlVSLxEdmWRTwP1qOadGhXMGC7H6CziUAdTCINyXftKBqYsm09bwM3Ose
x/iEqAb0sa/RnrmFXJkS0AtBA3hcSzcZNNpcgev7r4oP9jVUrPuQQksAJ8/gFv+5mcmq/0ovVLOS
wHxSqhN/2l2O+Fu39dLaQtsfbIlvCL9Y7ZS7E/HrsoIgof/7/Jb3V0cXjVmu8v67pWaSjnBsTlUl
6OZSqTBLJfb8fbFN/cGyX1KInbeoN+VFOavOX+NjD1+PBSRZqxr35QcwS1CXBzqN+1SZrTM9LhmT
GZRd65/OvBP+cQSYcplo3L24BusZU/w20ns37EfaOdr2bZUtl+76gryPHerqk0sCChdlyzpfb1Qt
18qx3KeTmV2k83dd/roQqCpBQL4boE8AglgbdYgXZEZLjFxrVPP3iOmt7bcdB2yN0r9q+KkN/hJr
uQCqWqeFQsTFsnkyq1Oqv4Yk+jBJ/2TZdymCeOjPH1TdDKCPDPHoYhXCinqJ2xL5TUptWEQDE3se
NsO2ffv8MdbAzOydQj99R014f8QcZGfaG4dKZtud3NJJWPw7afxx9Mb4UO6wnVXXPVnPAamgRx+O
GKtS1pHMMdiQyHex1sLRzu6AWLYJ7SQHrX801z27urkIsKfsW0v45D/xS0A575ao9Zbgv4VVxYau
yp3VbPTAp5gVUezxJiK4lNf0Kmb7Key5TYwA1YKxUhIKIWqTFz7Sm2WbyVaLMJkp+qFy9fgGDizE
CJ1P8aX/blfiWFouQBPIVawjTuHfBpw8fn2hJGfswbsRH0ECYxS7pf/6SSHN+KD7GBWfexZVOlPJ
GLQkpWLSE+kg0Jq3WYdySiRmNltOnEgorX+gztgXck586E2VGMUXKVfGU7rsoqCxYqE7urII6hha
VrOGZmP/G87walR9oqI4YTeeFbcdfxk8CikOkZ5K5NVaWj8vGUZ8b1z6dBeP+VWKUy1+h2Xv9yLu
LDFXXLOgZ3sODzU90EOLp4w/tgWuSbEF826QbUekTFkQNiPpxculDKY0cNlVH68UTL43JT7wJiQ6
GiRyK2rGryOwD+wy9fs/Y1rgAHLx6DkM/kpMR1HN8zz6nMb3u5+IH3zmLLbQ3jHEgO2hbafeBW9I
DqULxAVNS36cjtJpO96SyE9p3PKpHCWj11QOACc8xhcaTvv1XPcVF8hr5j2fC1NlVXiJKeTjjdHW
4B24LExYLAMgIsrGfGy3Puaxx1AnULl/HkF9EuA4A8ySE5/ZdbScHKoqR7dwRAZmGcT9YiGJ2E9S
NkatRFmf+O0ueSjWaMMvM9zOpoCd6bwdGa9ITWIuV2M764LyKWroNIAJRjLGNrDEmjEIYprZWF+d
YwmNvd7yMtg5lG0HUt+f+R18rOPykGmeOdUDLarDT0Yj/1B1WVHbyt5iBRTExgqVF7qE8byGp/9I
TJvnnlLttdFjLljehAB+A30SwBsKknUdAqww8JpmWikEEH0IA1xQC2vY0A81brc0mGRFaaJnGzum
ft6x5HRwCrIk3pWwCTBPKrq4ymgLs1jlQXvQrulkV40SGwprsYqNFcGbEMwoOi8sj8T6lWGejstF
uaBg9lpKrMYNVjELNlGCiX8c7Cxpca24lXq9qhglckRjaJp+KdJCuwEwbw+DtcbA/mCceCNRqOne
tq0RMxOZr1yeV7fSGGkgXQwscwJQcTGU/dIqExFSySywYUDgX1BhIZaj6GmhkQtiswf7IRiNGCFm
FU9hrxX+iuelXnyVJw7ylcIlmADSuHdoYtCYRan5dwCj9rhGpVeclHwd444SELqaLfnH+eJYM4Qg
EvtVkXSdoxM4x3fWG+Y6Gy1IhsRiuArVSizOb4YcRMSGpQ8WWKbBvdN4RVUwjkrr0ff8pyTTogox
LbA+k0KBuys7qWKIAVnMEPNQsvc58ql+GfnkqX/aawMiOgxe9U1gtFYD9sO0dY4KH1tGN3Zu/5aX
L5nsyJiEBBW+sDz7lBsaWkIpFPktt+7URA7JDljxjXl/suFXnKw3p9EdNqn2xPSKsKxOsvOacgvO
Ki7Elv62gk42TCgWzZnRt3Oja97p+RvEfuyYKjI8PoVg0/BId3ENzyeB4JqxRUVV6IBNWzpzEE3Z
neB51cFKM4YicXeMBHQtR+xWYhaEb6hEjYgnbEjtbW9wLcf9JNhbaL/gMTI8/GsCdVlcgxQ3wHfU
0DqUbbxXdzJUcPDwIWcea4of7+jrU8tQ1aaRGWhFFCgxh/DdsMBEzVpwsXxV2BVHr0MfnBFfSxob
MnDSs/Pwx24FcxDa12KOxHijT+s9wZlTjo0567jYnsMd2aziIEqSRfDjfnOQIuVfjv69UYz0AvkE
IEpH6ra8mhiG0XP2LHWuo6NQZWh/uQHe7Bpd0o6a+4Rf/VXQDztcCH/HyXceyQgZq4bGbR3G9EfF
zjcm46lsKMChXEd8U7pvDjUptzVOqMFCtSx2An11iZiuDPfPskkXyrAb2lgveKsAaQKmS6QTGPHT
LIz0J3ZFSZOGNvE1aWHD6f4hcCupDwQj4J04lmFtjJYnS2T20ysYJRAIhXTHE6NF+FyIGUWHcfMM
4F7tozdaTUmBVgy01HAuXKuCJ9Lgw/p3n0kVA9fAK1qPw9f1urz2D816kvQ3/Va5sj7nV4QqQPJK
NNmaT4VwEE77Kc2sBjTvMzzxFtgj1Yn2gshlUNM8p3Hrs8p0JTJU0oGyoIx6e5zcFT5BsumhmvDH
q/Canu00w7CissSqnYYoYHin/OuJOk7vW497d+/PPqGccY8OF20NmOgFSrXAy9WkqUCip6W+5JqQ
8ZmGFfuGJjpu0+mFids/nFS0Daz5T7xtTj6K7HYSaf1fHwZ1GRJM7xDkSCDzfaGQ1HoQvaY7c/bL
IyIScqvp6o0FrTFyq9EAIXTaCe7x3hotf7+eiz0WDfe7TS0Qw2fQKkslZ+HcBEbDXU4+1+zasbIT
2mDQhO46b6nRhx53S+yyi2y8tA27ACH2RR2jZoc1ElygOEiaN+N5NVfYXfFPrzBG9n5rzfcRKY0j
duEpi+a4+PzF1dTmkGqx4XnavKBQ/2RX6apEJWitQOv2oz4EGYdDGoziAReIFRLrFakbINJGMWog
/AjiM9a62GLnA13+EbkOHaXyiPhCOE7K6bMeajiy3qGVuppL0Xutr+3VGFeSyv2pcSfL+Mm4mJZi
XVmEDMG8vacmqPxUp6i6+KiX0GMTto4IAySDkt99lxXDQoggHLLgv3dsSaVLdNF3GBaJBYdBF3iH
H/ZJ/47Ax9N2VkU5Pb5B2BKSYc7NAmnTAK2Uh4gkHjOr2uO3Jc+y4JHp8+yMxpq8kgeeN5AfVBBk
p9tbugsms+7XR68frt+UsWQNKkFzvXynZyIDlBkC4TuYT4DRreC2rjnDV6HzEDygXzIocZ69K4Ng
3SrhylL8KAZCFOjq/oLQpChNr523ipndwZlPnJUV9wnsT6qMNxO/CdF/mSLczNkPtZvz7Ykt5IPc
gfGJPhtr2dt3KkPJFnf1hVjg23FhvKt6qu+rqwGeonmv37Q7MrZjfR88nCli09z0aS0V6F3wWh83
gVxXKNE8L9Xkla1Zu9/cY4g6/WvUaja1U9BdTj8e9CXTxQuuDLhT48a5HbNGblQKUtwbBNHNOY55
jc1Mpp9mOfe4AA3cXmxGja+DilHKdu45IP7ByY6fq7b/Z7TCtuVTik68aN/Pz/IoC+W57zGOUsd3
VBT4G7fpfSbJADzdrKTLGP9IVzkJPq2HnCFw6r5xA1baYEQfIRGkU2pGN6UY/CiIyewZz2i8uzZ7
zCOthAQCuiD15d+YXQ/xMg24RVao/2o8UjqXzmOyrn9w9zwlcfyRuyd3NBLpewQsWbHnTgPcleFa
bqTjzF6MLgIYat58OBcabruWjNo0mmOKHxTlMbPm11bmsnTHbf77fgUZQP8Jxyi4ypvIlCp/Dj3k
Q7hkY7Hi/KKoe5fs5NKfGceatp0fPmFz1ANz445u1UAUmf8NIUomUiBS8p6rctmKz8vDzdwcwgAG
3tMoulE+JAB5BlETV34tmeYPc2cbtFmSw9KpIAYsYbvh7sgNiYamUymwYCOKWLiqknThGAQHlYrN
DTN7YBrk5KNJzIN78nyVqHGHDBiX5TujxjV/qsXgKWsU8i3g321FPAau7dj4BDuecpQvaFMOHbSn
UAIzpsx+z8B3U9fFT0Jt9A/JWnSIyAKsCfjMPRUOJuFVhCQaxleDNgfdCvBbDKdJpqKbUKm2oVXa
paNvAMa3F/uFSV8t4WsWapJ5TwH95YEqyooMARZK7pGtRqnKM61r1AVtkdf8bZe70OYA6xUZNh3d
ZLJTv50iLdwED7DVM5au+7IXlTyPYr4NK8bfYvWgxC/e+jbK5xQK7ZlWcqFfvzEQK7Lq3I7qKf2T
4bInpzdcTKZRWQX7w4Lp2fGddXGz+RlhVK9g+ZI84Q34AV772NJRTEtmCGzxVgAyJVHsksznLgPr
0o1k8U1Zci721PVtzm+4a4fIHy+C6Srewadd69t8WaTsrOTDr4/6EPW6hK39EXMKoKsDL9sDlRYq
W7MtnMrfGazFjPsQus0OkKF5y+I02kpKP80muxwwrsKmHNOU/PyfRCGIctbrc04ChYBZ87KrulZR
e1/CsBnRsFjRfoQvPCdATLRL/w3p0F9w/p2wxUuEzTyH7JTIdXSk/tAzFPCPrlRJKEmDV6+Yoloz
P4U085oU5TqSutxxKBqAvM0e+mkHqnrJfPXVU+mD2QswvDiJxtzvhiqyOJvSL5TbFZytXys0XVja
QPcvih30Hs6Z0pp2q3YHW0+Td/LNwv80HjYyPdZ5O5UxWwN2GGntSbIL9GG736eeaiDWgXcRiZJg
TXYtbrMBN+3wmC/VWKySzVcOEYwbz9d5yCnyfFZYtjgMhPYDZsjBvTSRMHxe0JOncIi3rxFB6EMS
xO/+UNaLDU03DkhkRhY9nq2HtI62b+pnS52n8egXjRxQMCOe9EsWvtnd6S4SdnPm/xYgdWDOPbP+
v7MjPLC1LaDcUPWOhvpvPn3kMmFWiIpEtR2hsQftMAJCe7mLg9ux7PPQtuT6eVAlv/CRuCbpoX9X
YL4AVcSKYElvQfsJKVXSL4Ft9USLU6zAS12Xq1acL/tHXP4NNxjHGXckM4Y4esLGLJPiYocYPtOg
EEqqxrGc2p1qvqU+tsDFk6khPQuJAsTiZPWxVPYkPPbmDuCaKdM0TJQzuAg5T3K0p2WY6V26IPcL
OLA1J00w46Am9QeaTpOEaAES4Q7pdw7fN8CLvIqz4A1bFIev8MEeDG06P7dlvkJYyfMtE4WrjEg2
yK1b0on3tu9kPZXde3ojB5MAcT19M0xezsSSzOBcbx7f2LKSq5eyGTIaZTfU9yfbfZdOXcw35Dp6
7P7jiCXd+pgVJdHgzbDVeKxWp9JVYFWjamH8OlGQQc9TnWse1AWNWZ1eAsO8TozsVbqB3kKbOU4g
VOmMlFRqq4BJUEAn9vJv/+WRchGFpHrXtKYfUedpjSpZx9hkz4cBUK4kf2XOLoMP60LgCs8EkjzB
mH7G2rtlQUy9a1G9w72y8FosEfESzoyHrAH+r3fFF1sVxWVXoCNLgCkwO9eTvrBnZ4HZQ69/5IT6
yQoqmN8MnZr4XbgU06UuMkb0ANVdIkkYty8AUBpenZRpN/HmE0/cVl/MmEYs1IICNBfcU+EYC7a/
Wv1Ual3m6h5Dr8lpj6hj146VtTbcKvarq4dLg0weyXppN+p2415+JlF+IPOseNiJTyfE/GXUmKIF
W3LrElhNH2FSymMFTwOz4pOXwIOwBPnJSWEVTxB6+jl9Kz611/pNu93gUr8HHnAzrGk+MwHx9enR
8Yq/GDtCt0VKOulwSDZBAmKykQSkQYJ+xBvjVwMn1uDhf2XLeWTpxXoOcfQbgzDefhKDSPvJ0aT2
r+J94bS0hXwJeEUXK7VpH2Mdk7V1Oa60EWt67b4HM9eOL8cnotLuLhh1AanKFQQKbff7beN45sbS
KPHijd0iFYL8dsV+HrCkrmmsemcg+8GZ08n/v8jPMXTh4Dg5NWg1m4ZFUfisiyopwYKSJr1A5wM+
U1nyS0lQS1Z6VZlunfyQmDkzlXJYt9lozrwThQqyLdB6kbfBs4YDpNHgytg3Q/YBweMm1fiobXmW
YSTZvmFWQCeifThLojuVLfIGvc730aNVq6h0KCveNOYQ1XJGWNC5EEyhV1+VETForlAFpNfnVp02
jd1+6S3lJxcv08DtKvgHZQwetavr0TbmifCNaAQkNL5nTIabRkp45lmB3kEGhSV3Jvgbzre1JjRA
3CQ3QVUCHWDaNbX/R5d49NEPPw2zXuUyvF03SAaiE5xsWPvoxo0JHlG6QUgDn9XFJESSo5p9GEB2
Dk2g7xoxZJVznRIRKdpCVQjaE+9vCLePSCmwK5A6oPLBYEWCPcjZb/QuX1k0TseWsl78qa7fweii
n1p/uZRoPg29mGgKPZ/4C003nP1rAjLwjDwdEX5TomN0VfhC6BL5IRh0kvYGvJli3XZGw3OlHpxY
RGmTKm+/N82sQWqri5nOsJ8+gHpe2xNqhMo+wp9w0nAXaMbXSbQ7SfbUf2lOIeZ2CM17IjRVOPU6
Z8J1IzaEr7MFC5giT3J46Z7rccUju/Ytb+obvIba09U4ii6bbz0J7rzZ0wwcNtI+BO3npGWrh+w6
7ODZb5Jo/aE+HNc1soxysto2Mpta9mPptSZVCLdPnQjSx0HIF1ujpqNk57s1yINlFCp+ykT7yOgq
8XC/bVdMHAXR8ZgT4lifgDsnW1na87dfWqUhpjGAmtL3LWvGqfnKXAz/ebtme0AfLBE6F/0MEpL+
S1vCFt440r1E6RP3pMrYhucPVo+RBB7fG8YJcK41FElnwRL7uWAGQ4P91QwZflF6VMTaeC9UXZx1
tU8m1UQ+p5V6y+MxUN1MdwGX5Ska5IxaKRh3CSP5W7gnYxkVEmg4Qap6ae2eR5JXIV/oPo/wmyec
4f9jvLjo7ywfntuHEwJ/b9CmMQaaKZKjPukLqchkveNQ7jfeNOLOhk38iQ1pq9ont+1v1XQ3IUcN
QOwWovRjHjMbOK8sjHMpmlHDMnV3ZHull8ayuDjlLF9/COAJFhGm5bwbf0d4cYydriZwcULWLXFH
M6eoNpNYwHUebV85QyUapi3UjqDEmbJFfui7I3mUoj8r68aADgm49bEauAf8r9RmFRtOX+HkWgBx
9Dq2m/56HOm7OboLG8D54zQhKEDfmO/GjhyYQSVJEbvRyAjIJbNlg61LGj2/wMBgbNzjfOt9JJ9H
/ZHloQDValhyl3NhmactA0UQ2DFmxhAlSpLgAn/pbcq+q33oOc0i4UpaDXKJhAK8E8DDNqH6aqlN
l/tjk5bgzef7UpnX1epbOuvK3Na143wsabpnUJxVXYLeY14PkH75MT+9tUpIwRV4DwpggCcrxy6N
ofq7zq2tLobUtx/6yCQPM9PzVD2oxs7iKGBWnRRN1VSqQ96HlCuIwboz8nKWWfoKZA3jPrpZW3at
jVrG6+8JSlBwLkWJbl2AvWNE7IFqoz4Qq5ixPl6WgQqPME9x2bslaksNSqxNBwQjiDrbSCOvfntG
4UPko588u5fu7OJ+ncO07lPTBXvnbFinIvheiqbWL9Y0LepMsWlmfPrMid3HehJPzDrMPnvlxIL7
573R+Wx17xbWvVw1OOLSOPbddOJV6tNeN6O5eWDsfwLmK7As/yXT09lu1oud3GodYMYnGrkHIbN0
H1puXqbEtrTCGXspr3veiI5gQq7jISVngjgkCt2FngpEtRhfjqFgrfPoRfbw9vSFlz5CQ/Y5jKml
4JsSO/Lly88+JhfGKoVqrkt3HDMCWLpZ+E3Me6j9murOF1OtK+n6SpXWkmQ1UzNe6A0gyvOEcoVL
QFQjQE3L6ieLXSG7CW9lOu+/Nn9S6nob8rKmAS/QDgwZ3e1g93shrOX86mQcfXAoAiViRzkmTVo/
DXgJUFZVwB6IkZoml8oj03oqpTp2XON7rQvXz5lzk1wh5HIQxp+UqwJOANYdka2lU+C2dWqaiH3N
5vWx3fIWSiiTZJzOU/TYUe/QkOf7gUTh/MKq+6hXhIOv21L+WLQ3D+8t7LnyK0tPjpY0o3Sw8HyO
w76jyJNSLuA5tUmva41MZW/+dq3T2/4YcRK2WZ0FL38WXV+ZmE1zmT6Zj1gguq9DIKSzduIKxHY3
5IETfXKtXH0Yk+Bkk0lGWTEBlBBEdIIxcEKhNU+9h7EevsJCHnlCz4d5foxjGVAUwEPw1aoPaOHw
qs6N8FRTAmDtd5P+3cuJHX6NhJvp+JWaKqle/6rTAzdNdxYNqUAv99w9UFcw3HwAvSXHwmeGdPri
Hi0+BJSogKfbyTemS5Jk0xQQYl7+7jkiqa+SHEYPpzqEH7cQHC+WJmTqHkiZ1QnB0vW6jDi+wFJj
QFtT9Yi5GjETnLUftg8UP/4m7e2YS6RE5Y8kZGwIcOEf0UkKfaj3PlfdQNizd7aKM0ME0L5aiCm5
AMteIEBrWioUK/3WwGivZ+u/bMFJySzQPLCMPUiFnrdzyN3R4gmRuHQQWFGrCXH70boWsIScK/+0
GKewZByKDm2s3TfZVkx8KCflrnRCZvg0oxILyV3QChXjX2VnH4gROYxxO4soZ8l2MrXdVNimGTTD
+Ysvvit4B9o6jQ9H3TDLsQSq08yN5M/ySOIOtxna4xWIJ4UszbR0tpmWkg/jHmmYECaz+WUB5OZZ
X/C64aI7qYEVmk126BzqGUulIcEvcvItGFQiW4nBICxXh7l9x6J9H7x9v0svA6GBQP7qVa2CkGh0
MhzQijqu33TfLWVgUhCc9AhtU6J7byp4w43PqGH0+SLfKSWxQdDT7BcjB3vT7QWWcs3yYehOx295
0/XqbUb+FqLWSqN6VahrUIAO3iBj6t3t+ordvsZUpfpaW75Zef8KB1EAZpc4HFZZr+9hEOpikxxC
QoOJAqSAyve+yEw1En6ARJ0XafYMJHrLxVIbDMb61mFpPfhCeFvAChlMXVSYAv4aqaEJFnttrdS6
wXaTueBCfUJ8PMrdWtC/VHUCoaxDbdCACrgMA7bqvzR/oyeT0EHXNod4IZ0MkvglBMgQtiG5ioNn
x2VYIR9dmvBYdXQhCgR3oUdWE3JXBzmUv9EppalpyIJYCK1lhQ9XtX6g16rB4j4lRp3khggPsRZZ
4E7JbqCGPm69mg6ZpGjRJ5MAGJCyITCbPCUsTJfMwl+ccUe1QGon6xZ8IeaL+Rxpa+jW/E1TJOvJ
b+3mQLZ7bGgOE9FU402F3tTPRI7hvkq7sYuNHfg5mt+y9Hfh9R5yqd0C0lq/xcF10tZDXNZBfy++
AB4YYmrufeTWfBIFkVaFjPWP8hW9MXrBcI9ivBNKirIKLEtD5sQLHpeyiIkXLz+pEZuU51597ohG
a8Wzk2OqF1wbSEeGNBV0gchsdBWPClHF8qKuTqgPmQ93jU94JOOZv2FDYghmIMMvkhJe6sJblhxI
VjUKwoP2fC0lEWPmrDTSHyR47VODL5efpt0nwhKIbpIANXjkygjXmcPe+F4gZcdPCCopr/HuNEP2
L8toGSphXtDG0wqU3Q6LwFtXuL0Rqrcki9JnKR4CY5xBjWXXO6tLIA4qtScyb+tMOtz6thg3an/x
KTnf2xctHOyjrdr12reJySbaMCbdznnITdonU/D0w/peM0ioilfak4OBt42dAORND7yZY9/uV88Q
z59VhF8QW6fIXakhJRU/hSqPFyU8MYifUv3ocvKR4/jibM/ttn2Q9mfAbiU5dhAXaNBybCpOkKNL
0XxZIArnbUbXJ3ZRRIu5mRXm0V2nh5vQ3NHl6+2unnd0Q/10oNMjyfahYGxU3qxJcB2ECeFaYPYA
QNHaZRGbqnZYcCOBME2Th88E+5QYun+t4Wr1gGngyL/MnhlxchCwXeSFvPzkKOD+zs2EO6f9fCWi
OIusS0DASyWUPS4HDWkRWYh7pj6Q7BgOvXlX440x+m7rBUf5yxxiGytTXpLZWCNFhKQq+H6ZsQiQ
2dhqJZDmUPaFtLNYfkVIrh3sb+4FTQ9vDpcqGn340p5s6YQCHP8NLFPJ2ZqTqeGhHsw+ezL91pKy
XAXpZjLZCMO+hTstfLd55KVhtGb1nHODixN6tVGEh5XBUG2lLUpBPsOJU18FYZKLmCNJGLMC9H1B
SM22aQICd/+aPFdeoNttMadKDQZ6C/NTAzSb+b9Uf0TaZObjXpXEBQUvD7rVIUXP4/NU+SGimTTQ
kicaGZZiTJVzdnZf45MvNNvr2Ao3n9vsCq9biP092gYnl09mjsUiGWWjr1fiNmJLANUEumocEk95
C+zDy7dF0LVzg8D4pVAw5dQWs8L/S6KSsTlQUl0j6naxfQRtKIHHvzhAgSZO4TXruTuMSs+xn8Ou
dnblYxvMpeKcyqQuYRVRw+UJvuyhl+MiWZ4tc54umUIa8VNYzCdCK4wfjI5/i0wWLLp/kEVsodge
cfywgW1om8wHI7UpZ6mbUkxAYXPyFY7hWR1ZKCu/SRoLogrP+6xkm1FylS9W/KZps8snvNgIS89c
qLiNpk9wkDSn0WMt+0MKoCnIXG72wBYN/HgM48nD57jpZH03D6sVqRAr8nMto5P0y1U8jTkjzg52
WaL9zYF8SEfQleugKA7jhFLi/zZlw5MGodlEJluIsUQD77f1SWSxhGaHZ416Wx0HaVdXyF3JmEHo
VafbyUnUnQ7zBke/IVexx0GdTu2ySWdb8EhplzfSI9WUC7a6Tn8JeK1k/8qUEUZNlCSsArtvRF2D
pvb6jCSpokxr0TDppKuQ2IjvO/tiFz9pT3LMenR4iv/4qMJALlxHTOdSj7hrVNEV6zKNs2RZR7NH
IKULz+Sq28Q7W/5ROHF18sTMo8YrA1Bd2VsrooGd4XseIU7bgG232HYQ0ePiM/GghCasF/IdOqrF
gjWpILpDLuGdlVZ8QF40h8/IB8aVV5LLUwzBuFOjeiytOSZ6b48xBV34nNhv+bWp5zKkWWmUlt98
R0BDcTnKzdMHghI7hZaVyR3e/Wq/40PnFMm7pgtmyZCHd7OnvMtyl55TwR9KDSzYiZmYjhh8+brC
Mpy4cylq/+jMCjdZqJIvsu1TPCQnN0kDi/5HEOpExk1jOTYhv3poyCa45lkgVJ6H0wcXwFryYzqU
4pxkm1NzTnbqA4AfE6JlaiPb035SzTCVxM2F/Im6rBZ3YtZ+R29knWUnAT45ACfxqUzCZ4GIBB9t
E5KoGlh+YieaE1uwPLNCUMD5lx+FfH3+8mG1FhaaMtVyBgNg0bNciyogvnIFXPJ4s1ZILiE9mhUx
33En1ESQ0rowiapfbGF2zL+BC9IerGGPYcLt52nba0x54mrYXOhUte6nJtvEuh2dNmxhLpQZllK1
TuCsueqx1IUb/n5A96o+DzD5Wqq7udh/lViRDyaZDHZp4gKT2fX0VEEHxpkS7O6JLc8PKQE21T37
yDlVJwIB/AexYzhBz0Q6gzOaIFfhPV/c2yu3niR8bwMfXd9RVtJqU+hGNoxA+rpqvBkXOaUEJkX5
b8BGAHXL+09Rxkz0cdwcWF5atBJw3PoW+jk6K4Cpsd5klI2AAHzHxaW1b1C4bVKAMFfFsU0dRlrN
OFQ4D4bfRhr1sTvppDDcPEaCPiHsQ7TiXhUeq+tVJxb6n0UQ/DXwFw8dL5v9Aojtx6XO9HvWhpeb
mPy0wUiW4+cpceUA2tqp4fYljKQXOO6UNuOn4ag1DxMN81D/T8oVZhUyRsNDZ4Aii98F1a8Scz80
y81DVG4dp5zrR36pATzxrPbeFsa+sJg2GAqoQkPN3v8x2+Ja5939TTiJZKWhbVXmr0T06arNI24+
xU3cUSfQYLqml9yIErpuCHZEFRzMVLPRtra7e9ftQR4rW1mVUorFooN/LaaDqzOa/YeqiExD6bcx
9LF+1L9fU4uiNW5Jb8Vn7sh5KMe1ySbcWRvA570CNaRRf8Tu5W1f0tIUi7MUtMU3NG4GG6efKleo
3Qr9NUF+MTYo7AQ8I8eGdFgZtXaUYo4p42cI7zmBll6bHNd2dZIDs7w/5ryEy2x89vrk/uvZQYp8
pnEvKLbFOD6rCTuDjBflahF0ZsHuM3+VbdPP0C04b26lxvfnd+hdH6Wx6YSWSBqXbIN8+wgXptUy
KeHfWuNyKRrvle9pVel/z1tJvplc1Brnje9iMfjeRhXkl5v/cN9p1MbG4/HGQLaF9V4NnfJHrjrx
YCZSBw7cLtRfAuAOkLgfgtIHbK+u6Kv6xID1z/9JUujdayMtF8+026qkuBBs1XyQKynIxNlWU+dp
fn8mrFtVs7nB1h1LbRnh0nMNhAqsrj8NA5rxJ52xEymRGiXRFwtSb3wNA6YYFNIJ1xf83v15X1Zu
6YPkQLZVOoV1mBUufCRnfnQSPuTzwHOQe4kTb2zrblPyqNE9y1qr4QJUenVOpIIeRBzn3/a61Jfj
j4JCzF3qC748sQULS7iKtxx79tCx11NS6TLAC9cv+wbJWioyY/sjraINEo8Jj1GQTqrmrVJ7e3Ll
0FCgt3DMONlXaxuxdwe2a2Ar8Lv1Ho5+x/T0kExsRk9K1tantoJN5aBwoz9hXWRvORdKxhe+dSxT
kaBcGr7V02BzSOWq/BJA+wE3Nggj6krtWzkWiAW+bRNHkUq8f1R75J46TvBpd5HMrV+2y/enrdDM
L+ahh8CIrBTxz7vJ085tpx0s+USyqZ28fQeNLtr/FQ+MDN7wFiV48oAWNHh2m2QN2TzibFNktuW6
JqfpgKr1FixfduESMXObJFY+MK7jP95gs3h1yecw3IGplREn/oYNPUl5Ji9wtYtDu6i9/z73M029
iTVpcx4UUKsugB5aUQBfB8EIitExnLNJx+7jauF0XnhGPCZfYBaOz73sOrIEiU8zPOpyYAOo/6RT
gFe+voablh9u1LHq9Eo/q1QDZpFzVo2K1YWRI/os3U89tZDd8XxSANwCJ9siOBW4juQNCjCnkxG8
UXtEKLwUtdsVpvURzdFJv6ca7S6JRvWEUvgE1ImOKcXVgU22B/Vil1Cx59tNrYUSnlX3+Z/en+Wn
qE4IP0A28aFEm3jr2Q19g5umP7In0Rq78LKHqxVMPswpSx3uI6typhuzRx7an6A4wsmCaQcAsKAs
+l4MH1Gd3RK1eqPxsb3ROgdBYrCQYB/AHe4RWbZToKnDeUktLibRSob5AoIU+qFydabW1Q4hoOuV
kh+K1WIrgivU8vl9nnpzekMaHLDDj6y7QF2BUxpTIliENOCf78HC5hoD5qrdYM90MvOHFXxk/rOJ
1iquyhiiwTXsUlfILk/wo4nNytsxMC9AxRAw3ZTPkRma5IGFMY5Iaw/e5WJO9FkanCexhyW/6S82
/hKSZ63W2JU/d2+f53HYwb4DzVeniGgZ1poTYHVicd4+W3PFYyqJbChQAhvshMR0PAeHbLdGio8/
f37mXJpxBpN6tXdW34rPakmKpkWv4tCuNn67rE7q/sta4ndQyN0vAg5bf7tHLYk/lpAnHX4ZZAa3
3FM+FojCAKyYG2RlCys8m+7sjsDJGlgPMNQL7+FDLkw/00X6CVvzhgtL/vImKxHII6GohRHUpoGa
OwV9iuZGQrrxGNEwvbk46PSqoJbiduXD6Fpqg1BO0Fc2loy44yUa9FGdHSylP729fTmwbd/bQaR6
Tf6wS9AZ36E8y8RkwYTZYSdd/ZvHDRAhRit7Ub32zc5nbvRjxH8jCD8bVKB+sopuSzLSrKqG7nIw
I1UfuAJc+7TsLmGysI7V5XPqS9f9Rr44zWU11X7Y+H3n6ZvqE2D53j8WQR6b5+KCtwN/jjqHT69c
Y5rkOaa4H9vcp5ITTi4HpHO8Wfwj6mJnKpQ3fmLpPJObgPO8yn1OPzd1xoPvVdEiReCX5D6DDmdC
mcxgy3s+Huu746Gqxw00EJHMqPDWX+3AmW2WAGmF0eQrHliiiv+16G1S2ibMICmVw+MTLQ0Dur9u
bVXhzP5bFVHgV5Ac2crsYiq5Ef94kPE3JUu73TE2FGRYPo/Whbm4NrYwm3TJNuauD0ZZAZuGOOgW
mxLMQV5I+wVsd6DVo5wjZYlu6oIZnVcQQ+YwJrHLQs8EgvFmX00TP2qLhT7Lw8V7OpGyUJFiP+kQ
BiN3g35zSThaq4y93PsPvGLXixGryaBOSmVfm5nuUNvUaIMLkA2480pjMHc6YczsPSdKlJLyBJS0
8m+KlStcet1NxCXE0rMEj+i67aLcAv+o/2mPiYu8kbRWYizx+cTpiK3uwol3sVO0HtwS3ftmCfrm
LOthPDZdGNdPyTzwoELoDC7RA9Bz4GRctaWTbP0iKua8KZyKoAUlZ9LnC5smssXY7OruUFPUvotm
yi3G37WfT3xrFcPcFZuRwlxONOnK0nIk9z3XMKl/a9LzI2psV6LhRT/CCcxwQfjjcHr0hCTiTky9
/anGC5p3HGfqnGu3yM04k8LFqKQfnblflt0q4VcdXsHZEfPErgOQzOqYCbkktRcqcDlssVBqrdo6
j2iPn0YGW46B+JDXeqpl0Zn7AnNgQ1JR8bKrbF6ebXIZ3TAQGxxxJOGuYLctss962Bw2mD4WjuCY
nNJqtyScjKrz0h6hHjTADSsPBRBK1L9a3G/xCFCpVXSRbuofbtqiSNQ/jZ8oJ53lI+xe9s0r1HfY
NLSbdcJF0Kq32HZbv10audQwPI1LBBhKGtdKRhlC/mlsZ+huMTFkf9NtUYUJ95kd1K86o+1KuDwv
Y0GTbcAj5e0IJrsr02UHux/gBC2c2omAUGB/gWmjMuBSPHqS58DESja3O506VRVbVCTN1zroSANW
20hFOA4P4nWmITIlyAzCDh5x2rwHcXXq1XW1SyJMs3ZqPnj1giU5kv3nKSeME1vdeOb4WjDQeW8x
IgmqEx0X+pMqroc6AVODcOlVtCmUlegmMSvVrb/CwoQe9PVolwRWG7d00J/OE/WsMQxQXCZEXdzV
DVRPGbaNFwgLuF4EmWPcuvNPMnOXwLaqxUhCI5ecDW9oztza0g2+D74Ba0TR6Yx3K90ILABue0Mc
jfqHrntGafyYjtTPDYP7VkT3vyj8pV3czlFcQ1fm1ZkfMdhbqpVKRwXYOGnx63v/7nkqXMtXwpaw
UhL0f52AoCZPgaS10P4o3l8SzSD4lJ2zKIiDCD10ZNuNx6f00BvVJK6Dm/mK6mRpPYV2CndC+uPc
iEcCmHaav4CiZDP+cXfGDv+IxI6faPTIPMOUCaXx11PmHcjyx4jCkEIz/10zpRJt3dVpGruM/pFD
em4RZ9lFj5H7AfvXztzC7CidW2fW+Acbb/pSU6jCuQ5sTc4q2FgiEgG98z74JIeG5uz+8jbWPwq4
QzXjjzptxH8KmK2t/DkwC4K/jO9aFuRjLiqa66sYvm9mH4PVqdOrKceUGy3k9RWuREa5weceedKz
wdjC1PT/wqfGJCUP6s2zR39GdMee9i0uu8kLRVtMS+eeCFHrSIwK0C+TO9BRqhmbaVR0dY1Cw4gd
yGDYdbGvYdw+vrpClGOZLcQVyOBJxGtt/rVAuKoW8yRJMCpt17wNof26vCo1GvcalfKqINREoDrx
yjCZsmnLAWq146hOD9GgOqnWa43sPrJz0PBECxokApU7u5/srf2dZCVy4kdSsSZFsCd+AzBwFwCW
ZWTd9wglusnrmVjznaG8BwywuAhyBreeyRppJstPENw2usfPWFUXyx5nfKhG5Tfi1PY0owwHrD6x
MYcvJgY4HA0kd8HQAI9BdVSd3Se54xII+LcXywxjhXDCaKpGfBNgm+e8f6mm5JGhq2xThW6SRkbo
tYI41/CMawnYL6hE8e7sNrS/wnHLVlsJHSJXWMTpKTqc+2/SNu9M9vbPpujQ7QqFst3f2Q3kkyC0
2AGjgVdHhpm3RTj8/5nb62bdIsQid4iLQXIslQ3DldD60JK1lMPXnSWO9+FJ3ZxCYFyFaudom1xA
NzLEqjnL+8dSUf0HnoE7YlrdQsdL5Y26/magqjjLTgnEuRV6Lu1brEQG2k2oz6STGY5rPdPaVsqu
IISJRYBJuwNq+10d2Ceea8OxrFyfIWAx3gN9uP4+kaLrFQkZutYpFK7n7uiZHJK8+VTYxsgrGijl
YH5Y6OATpb5ZBVftgMYw0RyUI9sM5BeRjQwS/6KJjmhDQrzUmOfgXhSZ6w2/JaXlIwrQos9it88J
tUBiKj7QJFVXjuvgY4lgd/0QGxZ7LtYirp1uLlEb81WJcgtFu7w8+vVm7Cnc1RkiHakpD3PMSehL
kn+riGtVHpmGueCuLvVNMH+PGEvDqRiArKvAazgUwZSSUVZ7nTQmDraRYSEgV4HGgHJW/jWdN1aG
w2TZQh7yMd57DqXtKlp5j3PN5Ki+eCMcA6fDpWfLIUqS3j5cyZzsTmb5casRiUjJFnaqmgMc93JD
iYO69RULnL1qzadb3eotaXMd3DvGwiX0R3YztTZvqOZNVUUhaBktqid6gOrzj50xo8lXu1Bs+Mp/
eziTw5n3oqWH93cUspQB2A7LPNxfnnhbSd/XZjQ0oupBgJnI8bUJHLyFE8Bn9tfJzXymlS40wFHn
drevPIjrZv/TCupT/7l8pFBavSDQkN5gV0hj2VrA+Td6fQ8zUmOQyCIyUXLOMy9jut8nL96v6R7z
YXWpSx49XEl/RwwwT2PYDpcZj+Lmpux4Z/6i3pE0q4lYV6JFes0DaIIw3lv5lSUcTOTvtdX7WuPf
74E61h+gZsf/brFX3zMD0ZhfYoGwR2bdT9CptuiZOHiED6+jlYSrky1u+UhpA1PS/XuVScCtqpqW
bSrBBff+JLTc03UZNNqPvITTy9oRU9AoBbUarNg2MLYW0za6763TiMRRSCcS7MtZtbdTJ27Z7AZ+
3p6dwcjuexJRvlfJxg+nLhVuyxKrkj2HNqysmRFgPLpWR9M44ow8o9qiQOkqnOJH0FNqlIJVeTs1
9QeDsFQydHhi2aG3BTBUIoR7ve/BukLuZidLINWxonFpnWdaJ4EwnQ3xykmYXCpvnMEEkQWFrT8v
XBlSPwJod0AjhcQ6TaVs0A/WnW0ETUC87iyjuBeBKaimvV1J3/wweqPKAlwVtVIJkMyaOV8icdaN
ZvElNWTPRvyFn1tmgxvEiDpNBSWrK+pRk7JXjZcdYb6swOXWeyurgvkn/zN5pFoxmYheK03SQ0ra
3Z9NOuqh7csCMerT8vokhlXQT9258T9AyoH80lfh9NLjeRXF00NK5eU0u3ececGpYfpI8rtQUs/1
HA+xKXk/0PislcwytG6cZn8LqBgSufKJutz52kcqtYPOdTJE7bNaMHJaDU7pWFvjSW3i+acG3pNd
/MpY+Wvp9nJcS7UJip7tMlVNXLved/WFyAz6Y4Frdv3urD7tG20NGo8u1vcswVAk5CnM79HHaL5s
F1GVIOcTmXROgs+1kMR/35cUhVpUmClzZZLFRcW2Ps3i81Mckx4eMPudyBfJ6fJsXIRiHA2bnVdt
HAC1O8KVbEFanOzAbfQL2GbMzSCQ23aCe2kEIWihU5vqgbhRpcSH3j5O+90LCVT1l120crYjk7z2
a7QP3Ez8xAajvEUO1WZHeaqNH5oawol+6Pz+61tN+b3EwSmn1uj6/X7zKeP5jCGhbp34sijuSjEa
PriF8RFNH7TFyjR4OJHGRoOno2Ab/8tfSoT2tk63CEL0WO1h4te0sz1IDDe7bguAR17pjfpyt3/B
fI0jY37HEU25S4cfmgsOsVxNT3Ikx8teSOJNLexizh90NvFfaT61BOLm44bpTTlHkKG6x8NOpGyt
VQfLHqcCY4leNJiqSxmWLH4mLWjB8v7Xc1aEesI13PeiQ1lOnC4VzlqDcVk8hmTrdE7ik6Ki2ZVO
7qIvIqzHPOTrt4m2wi+ssWKyUBdS7gA9PEzTQTV63afs8aexradaN99wBwkA7wv26z5QuIcKWwo+
UzHMthzef80GUkbrZiJDdPV0ateQ4myXAyqsE8DvKgIXZH9SgJ45q2o2dkuZQVLtwHtDHnnErzjt
r9+3ctkmDCodW+hTYl+OsfRhf93bd1fdE5hmOvgSCvj/8xmO1YMRYthm4pjipDPTZXkI9yUnEpV2
OKDv6sTRKT6My40uCwpOJXIF4Xucea0l9ew3yi1hBV1aezjgUVr5Epdq/I+L2bQwZP4FqIX8371Q
k6cOH02oiO1OtTqLzcEPeQIlmXgU1iIvfltjWPmEdIaywt70XQQKPt+HUeZdeSqHkbUQhDEarURx
nz/IQ/7x64nz8WPGP16F4DSMNtpVUauviGotrnL6RUQHL8Hf/Z1S4LQHnSP6RD3m4FRmg/GOE41O
OUTbvlEfsWsA2V55HVHSKNlaPGJz1o6bxsu+886ji4423SfxlYUYBF7YXR8ouuK/j0C5kbYYQ8VQ
2Me5wuJnUMjyUsleFJ7ggWd+ADBBDj0P4HJ2/fvcXVP1fpPxcnW4zYxyYCzH07MpeeM2kNMpe58s
+GIitqRUBpbC6Eu7GqSSM/QPiXh5RwQ+bOM9auV41Jl7rzekdSAbXjsbDmaZyuR5zzzB5BYHma9m
6G4ZJBS2GwPnyEwDHSvVJVuNJTB0gpLxmGKQOUxG+b/yVJWaI3iQUjBqLB85bPfBg4LrfH4CE7HH
if2lquThcIeXQ9VKP0NFLmlV3/VeHNhv19uYw+ULyIBrCj0/kLvSlBFLbhl9at7qE/LBHAnYTNPp
G6cOU4QxPfTpowshfnC4GBvnLqad+iv7lPONSGmFzewlHxFizOWpVq9jjzt5dZPS7mMXS2L71iQD
8RpwCHGVU/7iUv6fwS2YgEaoinuR7tpK5SJR97Fd8cUg7qjojCrgfWpInlUi6r8EkMTdo+7ZC03d
EUUuYLZ6lqcjHwZMIUNmW5xBr4YXyBQal+fPKp9xS44ZK9NUYuFXPJJx4AoA2Begam5WW5T9vk9g
kSqAdmGMCnmXaXBxnGqTdQp9bqNwtW+tnsCesu12zC5BB0Ne3ZeJP0tx8hbHEu62einFjb47UlPg
77DE75J9/ty0muE5WkL5cllD7nS0LZCEYlKuoB8Wc/qrq2CGEQgzH8kpR2IkwwOCeSi9uls+PnwR
EXObCjeccDMCsHD0pxgp1PrDPOelCr5QmQFH4KTWS9xCMft7VAHHgF33rUV6qH42bJJGx4EDbYWw
dfFpAtJM7gd96lFitVzFrvoS0I551btZkdiNbnrcOd5EhecUVU+SC6c8+0QWgLHIWIrSWVoOdVcY
WLXBoqmQxkYY+56NozhgPLvP3vmDX8qyiXI9oFWX5VcV6MQzypS1IEi9ItJQC9g1W7zEdSJdRnxJ
LpAMaJ9v2N+C5yvRuHbdvNvJVhPW0DALOWmxl4FsUv9LiZdByV4u/vftsRMJ47PGEkkKuHgLHrkt
uBY+QTB9alu+kObafNOcC5t9NMtSQYKOSjPpoN45VXH+1R8xRUguYWcWRlUfKxdSN8dPng60qf6e
VOO6xNE9hPvyJQ77EK8y1LkEll6X2Gu0yiMvVIBmXET3KUn188p1xJJeaCt+Ct871LxMRr3FhlY1
QPzYXRmdZ34TlTgBYZXZVv56RT4j+u89Gjr3EgxbMZiaLyfNVVVtPvNp6VRoOMxiM84Xq8tKnls3
blmBKx+QYM4cJBQn5Oak2AjfVY3deeGzZIIXMsDV68CrQAKrJDeQIBMNEubqvIYsshYPly4I+1xg
gDXiPmAjuyGi8U9OU1v7SlOzHuKfx/5EAujF7AuEcqjDsbU9vQV1Y6UWBry7/rbJmpk5nA2Th1mK
Ox+qJ0rdQ6XUPH5639VnBSj+HQVryqBbTBmr0uOuCLe14an7gUGE+GhKEwUfkv439x1CyhZBg7FA
pi74wkRR4fsvNyqmtWYanimC5TSuzdtqf2cWOlqUPbzRf9RSaEzYK7f4CnX5WCAmoBO4Co9hcmP8
Wk1EbH41ByftuKA8RmsajdOr3Oeeo82bHp5yWUkX1tsAOVobndp+OFX31LSUArxfNFpd/W2uA5sG
Au1oFUqSI494JBWof1YSP961nLwZQn1u+iGtmQ5Eet01o8chVmxJooOSNOM23GGGtTYX+7v9CT7J
n765BYgOhDCrz+w0FgJ2S7EuD/y/QAyBOkslAvRMKAXWHWqaw8VNV9KiWKIvhD6nb90dYeSF1UpA
XKK3PQ7fRSsXSzXRiQsfPDYsnq+/K700BnSDQd0oNfh0Uc83rQk3TnEGgetZCC1mF4DO0RpNHukv
zX4S7gSrqYxqzU4CGWUJdz8fpp9LSy9YB80/Gm/5+ZslegsiG9nfcA/OluZOhATlqU/50UmWLibR
SebJUxwSjvDE6DOUX3OcOJ0qYxguLpO/pFSpAxKNWMol/vjQr1suGSp072F7YI2XcvxeSkuCCQA7
5l4gffWNgpnmRL0XlKI2dMRZ9gTsrRjIpaKs1FSNpe17AQAMRaCWe8aOUJ/ERz2741rbgjvdWUu7
AklK5+QwdIrh7Os24Gio3zsMmIOl2pe5cLolBXbeqVecVoF63M1fC+tcXINcaRe3UU1ZNLYaq2Kt
gEmM/rvztW6eRsVszi1iCTxZEOCEkoSQtUzS+D6CLnLkBrGms/JeA3igERu7bZQF744PdpH8PYDc
msvCA93FDBauttdmfNS+U/oLdJ6hzVK0VsNv7SyRfpMBArqxkeM+WdP/hDwO5QR54eqZLzFkOVwI
jA7M9hA8KAMqHsN3DhOUP4Wf+3yYgqctb5aDfN16rcBppPi7G3nfWFOpvEg0/f+lPHP2FkwKsI1F
XK8DeFKa0vw5njLiuErfBO3WLYKNtgfyXyg8YwDXlIryQ9WfVT5DsSr7kb9kWeK6LSkW0DNf7yTx
s/+6eort7ZTep2rGxTRpE9qrLLwYytDIqkimldTsEvYE8IIx0LfCM3FTUHqL4Ifg6jgzpzWJm8Qj
ZttPw95OYSu7SdGG+w4YldP62EhlDdok12a8LyvRGXNAz97HWiAgoqhiarZxh7/dBXXpi4Y3gVGu
IPCfm9043jpUQTFq2Q7Jjdj/ZocsaqyBAfu7GHP+vWfPUhfQyaQKBVpRDxiE5bZwiXBu6j5yas4Y
sqWqp/hPLF1oeFBk+8XyYrCOYJffXvsn8bJ9HDKQ7PDV+ZdRWYnmr2fmc80/6K3zRREh5qMHqUCw
+8vzHdD7eBy3MWaMoCS/l5c/A2CmgMG+zqOAIoUQF2/Ys5Xfz6JkwqSQRnHAbbtO5Ff7YydLipbL
qKZAkaicI/vpXSjDm/mJPq8oI6wlg7fUxog+ksgJSNj3ADWz8MabVgz8oKLl5kKNGkptolPABG7n
kbSLVaz3LVlCFjMNqxLn6p2cEdRDs+/SpHJZbs/O5gw9vKd3HUN8nkzm0eF+yIGQsooJNOVCBi6X
BjKCAfHrb1SGV761ZFNGfAJ9wVGCnsFjvgJrQxIzuCj1bE7SDQ8AAuRRb6QaZ/43Vm+klhwZNjKI
pm1LxQSqOCGx5E4UhCazsQ+epRdWtADCvoqk4GVVGIPDuHOHGcmF3CpCC/LPq/ul0kelIcOCewPr
UhKn0qBukLqxP8wUVrM0XUEQFDYzBZ6so84IXejydaFSAaIQEkvKrqTki0utATSE7SB/h/gRnS3M
lOvcfZ/Muh6cydl1XfGp4idAOjj6OtqOfO+uIN0zE38JdCcGszx7BUowgmqn53SIOxu4EHRUOxLJ
/d9hdzl+gPPWkmapeJNWvzVrfWnoapz7D20jUVNB39jO8GuACYXgNDw+VNNt6WuxdCadFcBj2868
jtkdhNcmSGmFKUdfmYJLBPOtQg9CrKH81TntoR/Xz23KpnBi9fRiTFPDVCXdBV0H2GUHEXcdlhoh
+rlshZU+es8cpy+r928R9BlSlLwERrIjsAIS8yD0sJbUHmERAwgjsekcP6S3mLyYMPOcVLCVaUe0
EsYnJNDI24q7sXK6nxR1VXhA3fS+Z5OCJuaKX7KUaEi7OavDOej4uM4okyb3Te+Lalizgv24M9+7
pcTPAiEAFTcEiyB+yktZdmWd4SFMv8AU7utWVMGK8sJfPsS+MdnziUVi2gQIlspWGjiGpZUDV3os
z59UWqioqy1AJZLYKgHvlW2/6B95o7dypSdiDreuhqFV7Gbfyezlzv8qzNT8uCpsIVmiI+zMbtat
cRzJZcvq7wEppQ/8eEncYpqGpmpghooMu/HUxbktgR4zLMJSgiPZPYCO5/57aBDGzZgv19OpDZEx
LZ3kdHRMclONayT/sIeFcZlkDKLsrIzWvuaBjOVs8Np4QQR0B2nQtWD7NdVjJoj+QUkVgz4ibiWj
hTzbaNcB2//nRNnHwIuFYfGK+iXTv1QztcS36BWCF3HCz9NFPDCZwo3gDVzccTB5381UDiHGlw7u
JvN/82dUzv0q00q9bPdyvrRaw4MGOKPJ+pp+YZ9Mt4e7KcNYYAaidRLmBxVUPIDL6RU9rezGu1hA
ELeB7dQ9/dRBcJbEc5gJgWpHBXAkIe4BFbE36k0o4+c6QGltkJXwi8zAZXbltmpUY7JdIyZ7ohEw
uUDMPlTq9c/GzFU14IQKt9z3PDjMXmNuwB+Vrfv3w/qdjPzyG0cgiqVEKHmp/LvHOiE3OzTIqcqs
SJXqeog6TA1WiM/u92tpYd3vPPbaMokDZq1MXdU8o4eTH+HQbYUBPKqWNEquI6PvXDgCm6EpDb/H
SuZQ3N0uQ5nF9zLB2bp3TMycUPwT6fGBYxQouVbLK7CxHbWGb3m+VrlbcC8URVYuXP1hKJQVql3X
o7Z4wgZlO5N4PvWlkNMSqHxHrmIhTbN21IRLCOscX4c4z0FrRXe14qwE4unbUwg8QiWu50fyq5dp
GddDBpVIOZcevnggIj2WcDviFDeGCC53y4sBGN5ARKrU53X791+NEoJd3GWLIwL2cKw7IYQqWUsm
avIy6/qJsvpZ5WG7sdCVX422yOSPjyo5ruWWEXB0xqaf3ZsaFUumnj50iIW6EyCnkHf+mJ8sUnfT
YnXvFbZFpxAz54CbqIUAbjiD17NzL5lQ5ovVyTO5zaVVKewuHDQOqwC/sZSvutdd1r02kkqVLI4K
7N7BgfSnzA5kccsWabeESqKNfVSju8gVmxY+s38FIdi4a80euzdCKqgVlX0iDJwvPGU57VXbdIsf
YLGv7nYiYQuAuCilT9fs7/NnoeAAPg1A22KCFpJR2CvFaUocHVJdsTpE9LBNOhF5lAdyGkSu87YP
cYVTFebWSyaV0kmD7X4fyrW9dbs3BmHIbFcRhAL78gfAL9ymdgEJHQMWx+W4kbThuCW4M71q7EnS
Lz8E047cmPobRBbsbGFHKAGvKxIVAPUCUUwJYh+1i87PZIh5k7U4QlYfAWDPJuS2CAMym9/ZiIWK
QpAB9bIUhJ0zOoc0leUW1jhvpzb6D7jSACDWLQSf2S6uDD28S0NogXa1xHDNS48BoC6/KpOeLKFA
JvndqcvizcadwYXzFt3f/Xnnni/eKJGYyaNpz6RY72T5u0uMZCF/KIDlmFNDlF0uvjZx6pZ8yfrS
p8EUzbSw0rO8nuKdWlydkyMCswzHM3ULsctnhXpxewlgeAKa4drpi5uplx/js54aobFiRmmt9h7P
1qo/pLkWTl0N/OERuLlre5gQPoA0jAC5A/lXywpwPbV2Qa3XuqxjkP4hcx+lOiGPCFFyxlx7q+Ki
fi7QITia236T++zepJi4bMWbU9wSmevbGGQnhthKpyFOt4xmSK8ECGYU5CXceAh4Ty2JqNqVMuNt
b7ig6H7V31c4KQziGwO+7AUPY5B2T7Fm4JGoCAe/F+rYQifX74Zw86AosuGxzdEsedyrMaUBLaep
hO1XdcgSK2QZEvbY+zC945YRs3AJu/E8tTcM2FLi/ExLFq3xLvanrinfwQwMqN1kUKJvsOTUxzpl
aPEr4tqAxhny8CetmNYob/lKXlYQvi9dFq1aTm+Wuepj5tdmgEB0gqCo4O4n5ZQHN4ak4QCtD3IH
fG2irYB9GVUYxXVKHM6Z2OKuiRqRkZPYblQudAfDwpSnKvNr4ANskjjOXUWjcsO/BJiWJ/tQQ3kX
2nyPvTAtj+6/XUmYAGnasWaAAy9qjalZAIFJ+sYwX5sD25qxtFXNFX/2T3Si7LEPV4e9OhfFWXjZ
tXafvhRgq52lbbyPrF3A8zNhBLnthJP95I0VuXt1jaLbgknr5s3QL0FQDYh/N7foWRhukACV2N1q
HbaZORkzqP0M9AyuULRHO4b6+51+bLqDhIImnmp3kIFzvMSnHU0qEtP5E9wbEEEp62MPHz95B5PK
/eBc0/OQqYWoW+RqdE8WKgrKeUpH7CWQNJKeUsS5qcLixfMK2yNbXK24BXQI2GQmXiWddjIw16q7
hzVgcW5r2vbAxMp7edTYtVOl9JPCetcjM5RAYmWposBrAmOEFqwplXDzWQqPQjqm2qAnORQq3rsf
zI9VBwqkxkZsWednJQQXS0GpgOUfCnqUSHXmFW/v+QE3zsw7ONRUsloZ38uGp8pgBDbBm8FCx7XO
ebDcgrhWRHZPvmDKBwmaaLNFkTImIcWt/4mpPNu9DjPOzX7xuSgU0KQwSOvpzEtM4D6J4RRuXY8T
tmlN2BwsVqxardbgNjRun1Y/8Xd11fUJasqjaBHiTfabCC7N+z8SjCtFDQX/4v087DaQtQK80xpO
F/N+5VHPHvm9QCqIzBfpYdaVTe3WklScGUpVWXCZZ0YB/rTKM7ERvY/hgUEoVj8AOReXHEUBZoHQ
r2MPmucCIkl28GcN6o5NrjyRQ/mv3A7ZDs9nwN8zqllx9hbsnhQfgztAt0oEdSYvhxaW5WDg7VTp
swNAgUPd4Gtm9xd0SfOzgOYU372YbGPqHCfCfZwy1QmvseOuTHeIeiFoOV35dMvUTFPKSK9yNEIt
wIHabkVmIoMIJzsQnCWXXUbTITl7DaxTVcZeFoeymtE9qXjmlS8he0ExVTVT8wirqmTE6xJaId3W
qpm8FGRS4oNgKaSsNPWmn4J1laJDByiTusMXtRHFcFJ6aAe9CUiF8hZ0UVudx7ceLhngnFCFtPgt
2Qz3z8+53FXuDNJNTVm/rV72Ll+/kB959g8W3I6DumBVNuOEdNhUQp9/IhfZtjCsP9sf6pmfqUCV
nEHqAXSzYmFR/Cm0UcNbWmgVAGvdC/WVcY9TwtC3yQGLrpFNSlhtlqZcCJKomWG8gvCzZVzn29Mf
9WNAkabvwpWNd/MNwE9Fh78pddefFxJ8FNPKACfFDgbArvfJJiKxNA8eBROFO/QfzZ0hLSl5sx7U
AgTYaERVNFve6USBQtuyMl42X6oYTaAxUPzCmf0/cxD/2tr9rUHP+LJYCopqX8BKUvg1Z/oIgqOq
Y+WXoXmv0AyJBS7VK4/DUvYqY8YfBeXN0nQNYTCYjSUCsP4HV0yk9U3HncGWQe4a2gF8xAKTAFkC
Rox2Mzbjl7qem1qoB/LAKvmjdmWduqy7+nwtAlHKGtWFqiSiA+VoovIu/TfpwUcZ4bLTQU3T9MhC
mKqslzj5LuUEwd8Ay2oQuEDcTdHcE3WuPFcOwm2GI0bHyAwL9kL3ZGKhJpbGD+oOBm+ofAOc6DuJ
rH0ZtILRgcTxxI9+ru2URZaxSJr9W2VIUkhHyHTef611zafiQkzYM0RUAX/7DX+9nmsRlagvz5l2
ES47YKRBcFwFIwNh4/9AdzeMX35e5rNsHBEO+lrQU4rj/bz6sKIMBc9bYLCxTWceqnwGt80xXoAX
QBTqdZBL6jFnYQ5m+4r9QuJa1ha0ey31B//BMxrnUQgtob+0CgKgUZqrB91ASoc+ecFaJITYX4We
1OJ3vqIhSh4cOjkO6coOBaBTQxwWdpB5VkLOr/BhkC90qri3+pjF/9AU7oglEl9l/SPlURrOzewD
fPoILJy0/ZAClezTMn8JQToOQQeohb+Pjc+BlYvROL35B+oGM6TbTpcixDD0FNylZhAhl0n54scZ
c1c3QPFtnphgoIWZc97KSF5kqOWWeaAv2UUDgGD6gp0zDg0eBUq4obQHKHHLqRNC7zaWL3KDO5CA
OGE8sTHqFavtMCNtSQ30Yv9boKuOnnU1qVSEDKj3axCrue0P4AfJdZhYF50JGBP327mOw9mZktUF
F35mfp69OFqXwpe29BkgwGMHnN6mlOoItOE5FW3COFSi/t2Ir8Y4dhA1GZ0pEGaUOkCQmVZNavj0
794UTMw5JuuVlCotjRsyon3ncCcDLAV7yOPzjbb2N7TDYMxgTDJnbeIuMcIMShNgob4aLdQG0wKr
zoEtFTcpEsQ1p6+IYAZOSqdms9OEdTadRfNStjMwsTzTHEJnVvHfH652Cd17EA139qMONRgP95nv
zeiLh6Vr6m2lfkjQ+XfMhr/yFjPlYGaNnAvknudp4qx4H8tB2ImWLk5eFmarhUCNHAijhZKR4Mmz
6kYJr4xQrCQELd59Dakbi5qH5ZvoezoRSSOlrUSJDJoT+/Ylc5SjG8LJOIQo0rCx1RvVgant0xvL
246Sr/6NP7j5nY712InMezqaqaHvr/J2JS13OsbqEgtEePbBkO9V0/cg7vE8Ygtjpng+K2GzdEPB
FN0Q0OzaTshwXJkekktfSPL3C5BJqCsTT908SY8hoULL0L0ufqdF4vO/iIa6JGHciWUPHIh26jXJ
u29F6OvNZRxe17VVy1A8spf7GV9GbEL51yPsRm2JfQzMNVcvhCcuun5boTSLpsZrqxG0RKQ8KXTi
9oNXIARCd455iwJDWVuersmq1mvoUlZlS64957K+iY2YUT36tbn++UTNLCF0C/aGFV3VQPYdV8T/
JyIsSwoZ6t/YZfRVOC3WDG+ZBptm4d8aA6vkGxEZUbWsZi9C7G4bBVjUSCv6ipo5+G7XHuWlptJo
JzZDuVJfW1GRoCB2aqgMPEraxqnbybgr5MHJ7snEpkIuU++/URCHUhmDTLchxxMmNydQj6Vol5vC
GoSpckd07UYAl+JBRBaA6cZeVAI3imRjMjFUmejyE5QO7V9F6uGSrSwuRf2yVdyTmZ5CNkg1YJKs
Hx3HP+605CnJxhPd9kbDo3R+VMswko7qX1yJRsIxiYOehKMQY8E9VrRxU65FNvJait0GjLgWENce
sIf2Qmt3PSlXxuzVkRJXliMk6s+uWt/1ZVdsiT1FhP4B1zLG6apiT0Dl9yfy+AsxoMXKC69OIqQX
4KihkfYgbAZrIE7J5jSZmlmImSdfYvDIxFaD1lxZzSjxMngIrRDBmh/J9NEcNYcBGm8177ZnwMsI
gUsPKe+ooeYlAbDXjHvgXZ7vJWK1a17moNJXtouyoGZifPkHaa2d2ipr7/lwXJsmNfHPoig784Xd
tSjXHMagEhtRhFZJKtxdF7lcuTx1mOwFTXWo48myAFjtO9kSEsDYoYXwicnIaUbw4vZOFV5+d7Lr
7yIVhTTfFjjPWStM4x1DnWC+RO1PGXDWB8OXKSfHV0L7q5diAk81OqXTwOzdwlXauazImJ0mPsuM
bDzRDpnL2bLvJOfN8s1Cqp8LgklgPr1ToyCl+WeNsKS19VkeQvD1TEqnolMBPflsBIniDLw0YVFB
0X1Kq3pVw2Kx/c1JHnFds8nP1QN2Cns6xhGsHYQQ3Dx7w/ea4VbwLtrnNNm6ncP9AR0AbhLcXu7p
vFAT5LUrZAB4uAO+nA6Sn2+5ycm8R5O+tyOssNOFcXZ+z4zfxiZeMzyvdvwGnmHHuhv0ouv681Um
7rUeasqlJLhtcXSlWUXRLXpkaah4nvfs3HwKhwUHdmkjjmS+QbAHqYip/G1jNE5VwAC07rpqc0Ue
6EFL/tU4njsHnKPrWNt4qMrf0Vj+/zcwf4x6F2HemddynJFFUnF681suChqBmFDv6P4uQ6krUXjh
VstHq46VsHMdc7iP0chzZeGbBdphmXeXrwNukBAzl1mIorrnSD6ph2BYytTemYjVInmJNItZZQn1
UmOx3pfKIwZotSy6ufaMFcynqvl+flaLxrS0fr8EEq3+AEoDjXoaf/wicYOxb8NfFoMm6g++tE0+
NeodoJqdtzsAQYBzmgTOhvBQnLnmypx1o4IIBAD132YvlmoiLwgD2vMFpQc3zfrKm6vQTwHYF5PG
6qULPgllAW5q/XJKC0eIAxHtgumk0ULfJTVify9EOhWvGOTrvjKJzPSGtL9zmK4pYd169M4t5a4a
P5x+iprDAgDQjgpRslpp4j1dJUvxLVzM48L9NzGBrmCfL/WeREsN5lN0QjfeNLxk5RJ22AOig2oq
AjGYCtNRME/1KucuDwHKt8VGeGu70ozr9l1uixcnO8E4ttBBd6cZVUote6c60S7KU0FenVmANX4v
Crm/jTrbEQdrRHmVPN6jZzyIwDM9oSPWaImi4DCxnZ1NY5U+MP/zRA6ILRxrR01ab58Dr2YTq4+W
ZXScw819hCpU90t9RzvaSGkrfe7fphaJW/pygo1NqIS3OJdWQKBneWb9CK/2+unWDIHsz0GIWHbL
Y7hdvthDNrF3AUgGTpBnNAi0kPiwI90WTxmpZfHzIcgLkCV6/op6EziDNQ9Xf57IlnQ2eSrgtU+8
x9yGE7q7Bs05hPdKBY3Q1vmB3XOz1aprPXVWmSdxdih2Ldfh2BsqpkmN8xwEMInUK7VVL8h05NPc
ZD4S8jg3O+FcVxKvwrWkkny1KDNC+zWhrUKSfhKVJBsIFJ5wVqZq3f0UkBDahCPsBGFR1f6yzsQw
uSip3BMHMeQrze0B509Qae4+od5QDm/+e8HT/jJ+HEvAJoxNi7LNXCozjiikO4E7n4Bhj8dV6Nhj
KuvmeZerxKHdkACz8gaX52FPqjAVjQ454k5awj/L0/0HIqVeTqaC4J3xbEFVhZ0ElIL0dwDM0b9e
3sg4209gAhm7qcAC7+qM+olN1c/pCZH5f6E8OrcodEAmYRdbIO3TT798E6T6KBKUm8caYYRQncT2
Dtoovwh/h5ye4F9DWy2fVk6a77JVpnuoCa97f3DM12fxSiYBoMaUmmt1dye7Qe0KEFCLzuxHabZZ
YL51q8vnpSc3G17bSwDfGrrC1FlXWgnXT0IjMZJ88/+DkF3ce6XNRKtdr6HQv5fOUitfGBYa07Ss
JkAfpNt1y35c7HUmaxd5UiTjulNttjc6d5i+Y29ASnBX8R1aWOiv8KpWjEEr5fKhdO0T+sgNLkvL
QvgDWxziQJNdIO//KC2+zXTxIONLFU6hkHhBv86TU8t7QR+2kpJ9ZR8DUevdg2fOtT4VJrRLtuyz
DqyZYo7AdT24uDd3Nh/ONsuW3eZ2/tBZIbTYrqBEtBxOb0zuF3+LyKRaVuje+wMpf0ym+OeVxp/q
V+Jp18Yqx9ioditLdjuC62eGiCGy/H3YusQFJt78eJhGdUX9o3q3qso8ykUycnS5FOpajWBsNkm+
y2lJw8qnuGrIqegb6BRVJaVDWVIvV6+V0pW0Qd4NNcyRMvJe9/6DHuBN44jJ1vTQIEoAefvCr3FU
rsuNk5ZMeRq8SYA62bb1Mt84Npkve5gdnOipCdKLggkN9zuxzx0HtO0j+TBwY9WIszCQi7U9c2ec
I6Ie/UMkvrV54PU0esM3S/asUt3LcjAqSr4gYaPndZqx4T0yaeMUrTMLPNl6I+7UNjzjBRnj79SX
MVcsYE0Knze1MwxAP3aiEVeOb3pth8tnjv79cqnZx3wiDQGvbiZcYNc0oUEmuLGU+utP7nLMuViF
5TbjziT70kC/Uqf9VImKfcliWUqdIQODCvusWHMsNpgMo2dJHSgWind/tfdy+NVUxh9lSsKyx81G
MqO28SXjNxDp4Auqa298nxV2Fz5i+NhrySkwXF/TjZlOpGgpxKqneYWW5kNi7xzX7ZRnstuimkyn
La4H1Y4NjEAno+qWueJ7/2JNDc0jsnKm142BrWrtbAOPqr/zKSeblGhZ+d1yXhG1ZoKLoVO+4Ve6
dZI5RZ9BvQp8svZRhnWQWuzgbK0UN735Zeme4ijkuHC/8DdazgvIQLqUCk5FPfroRwZth5dpYOVh
7MwnXsME60EjKyyAVdOfgW9RwVwVnsfIv7kClB0TSZtWWtKjqKYsQRUpPaeoEKyEY3pvRT/h0Pvb
Jq1Yz6K7uUojttEKBsu0J5Vz56vwq86ed+DpaKF39PySCtUGcM1U4hx29ezleMwRbYQaDWm5wlXC
mLMeq6PHIj2B7FjLJiC35s0Ff2vT3Kdkoy+Cg5arZc6gilR2CtXmYGp5MiwMHKImaLQhixi2NgQ4
HBHA/zLxc7X/ghtPuAFZ2QKm03cns8a897eXRGfpg6EbJwIfDrwh11vnZ4PSiRnw235aT/ug7mZB
EYPtBiqTGsiNNr1YGX3EZ8sNCRFUPycBJIn5oOo7YLDUSv++J4dJhygYeh+ZphFweIBlmLujnjzv
ohFS3Oh0DQhTpzYN8YKtgzZorCawRvhohyQ/IBqCpoYHx5iqc9UCg1hQrtAZFgkN/HTZthwR695e
t0jpVj78k6U1cDwcOKWwN0CUKu4E98V12ImQ9Aett9xjLWTTFNTW6yJiOPyqiBxtE9zeZgxpVr5H
Z9z7vuCkz+tophu+p7AoIROmtWWxYVGJf5dBjGjE1w+sSXnvwrW15OlP5MibtH8Ve6ImbdaJsbG5
MrxnW5RrAGjWCDdx5HouW7MQo9UpAS+Dc+npxrwsC318wSq66TukO2z5jMhu8ABd0bQZ1PRmSegz
0hoxU8B1+9m9cnQNlZ7trTe5ouzpxIyHOw8RMvs0C0xbAfxLGY65xyF7hT28UqnIVWr+jf/KSra9
M4bS1Qlsm6ur2FmPm7VOwlK1gKPsCwLcOsabHO/lLkUk6nznUgLp+aG1jkBOUy3cO22EFTglgwJY
KpK1SBlfqK3mAZFlR1e1Xuhxlaw0C6DQczFqTfCrTTOwv0MNZDAzjsBh3dEf+97zptezKZwnVaTU
5Iw5RLLlUKO0ATSvUtQfrv//Xu2yL7Kt01ywSzXTKoYBcntBHp53Tf0qW9BeUTTKNUPehieuCufD
W8Hjgn9ruHcxgVKTJda3hCtQU+dhilOo8rHqGQk4BvbbyNFIjZ9q+iGUbjR2kJDrzGpGg5owe12d
mVNNWOoCqpffXnvkFNimFt7F1rVz/Y++t7mp54872W38GBVyyHosm04NnPuq8n5ftW0IHxLJ8WxK
Cf4EeSbO25/FZctY2/QrlVI75G/zbveB1S54RdB0WBbjh0ye/4pqxyvyR5TccaSQoeqZM/sH8PR5
DDWvrBnBADISnXjvdH6yQbz4QDVFJPjDD6ecAwLCSzrb2ebQgXGLT/sRCFx+UH9g6jvP+fx5Mqdx
JwI52UFrWl1GqrnIjwJo6cbFUQjbJtdMeCbR7/ICGjJf4bl59xro8+nOdVYnrRuWJeSeH8pdRnRq
X1GCUduIOMMeegTytPiVjAk48dh4tmrWsXVw8BaEdIJimKsFVbbifuKR/6MkiwGYOsY+dhWg7htj
tO9OMnsDBxvHB+rCRuqB5WvEn8kPqr5tp/N/tgUzmK3oTpOXnSKGeGNfSjEbpcUG43/a5ibhdJw3
tecLhVJfrHDj3SHEzpBOYQV3AqU2945oQHhEWyuYBjHXjIH+J6Po/z+pRJEubTpJHAjhUstC64HD
gQ0/qZGz5yUImaMq8MvPLx1YkmTKU87TCwzxuaOCEfDvTDM2jbv0d0qmOFiN9hhVl7YRVshw7TsV
GSdIPrzeVsuH2MbPyJM8c6zcvhzpmEzb0umyyYorSalqz0P++o/11W/bP0cJHggjPw2+x4SFWIYV
YMZHJ59ejNAI0Mukt4ezgEeFRGKlxBDRPhatcRYutrx7+mC+KoTznL7w+x0bxR3jDabgbL7hLXWD
KGX/knIY4q3j7IluwymM+Msd9o8M+MfyuqDOkyaUSjJSL82cFpq5FNMFDRvVY8oS7RavHpxF7zeW
NGa7DIYhiuvojcNtktTb8f9e9d6uwDaFKvKnR6rcE5fNz0RhPoWzqYJb8YywqzFcZ67XfDaaJDzh
j7OEqLycvW6WNsgsa7lCUn8z6YyPe4Mz9XF8k9GIlinvL6cLPHBI8ht8JYyEPPfNqF+8MoJ3eIfm
8jGeqKCymelHOhbAuGkf8zun+xfnUxpfGFBREyk1dgyJESD8Mbh3QOEQHkkbcnkbQJVKI7k7Mdqb
dZ+JO4+uTHbqHnRDTdG6KvWyD4NR37plHunAUoztoLEWkeNMYsz14KqFbORUTQw3aM3CX+mWsRo9
u4j6xTHQ9IkDlNx3BlW+4oFZ4vxEtUNL6xOS/wPowKdwT29ynZK0o/3H/mUkuGoTpJBVr+1003Zw
r2h+hx7yR0UHFz6ja7RMF328Zg8bn4TPGcAdSD7sjYL1bIKsS/s/Hm+h46I4LIS3bR4JGSMNK8y7
csk0e5EzdW/ZXUEcCk85544/Sd7vBTLb++SO0KXOwwR4Pe9iz+rKZjxIdMqyUPqkFViA/DQnI6i6
QEnauo+dddThzNK0u+8S9pYGWGOwZ8Cfe1siYZx7OrU3Fc7FJpFMS/KZlRU3Jr6Kd3/wdZ6JSpso
ijusvmFivgXzrcwfoX9OpXYtZPHNBTo9ueygMfvQdOYsSbhBQVzwbf379H02QsxHQkluKOpdk3ac
laaSzjtLSkRTrAN8Bw3+oK4N77xO9U3hNMBjZA1fnKl7ewvo6e4aduxM1XrxXPTRxQMpHHue7Y+E
hT28VQTA/ijlSLxYvzFTngIOTinVyValIAtoJU9EcuskmbdS2NER2q9aTQn4pF8tzeEser/mJ9Nb
Kqr7NfLldLTsg3gG/qCuqNlpvw8hH2ETps5d7h1zgTpgQJw4xPzsH/sE+PTziuQz07HBqoGTm7X5
5i20KioBnmU7VVfAMCpiBxrQjTUr3TmTYX6uvfpq1QntfBaRFtVcD5zEBaFTvU/vCcvgicTy0llD
cC9mJSVCfGKu1uAyCQ5KK60Gf5Zm34NDYRr6GrFT0PvkEti3o2i5a5RkrEuxVQztuxPUNJIZsv89
1uDdXaKo9oStPUBwFraYuwsqb2zYnkIGHpEOX0okIzorXJ10XskNyDNvB/a+VB8uzHK/VUCvWRNM
o0x+RbSNdeJW0jjatWNqIyYJppzCVz/MYSpdXLG9DDuG+drWOQqWoa9zw5ngy5+yBhBWneEfmk/f
rGv2KDUv+Y3aGJdVP334h+UNEBIzfVZNITndhX/MIpUxsrSTEXB5ViVfAtu0tgpZ9Bf8+WIpsaK4
7VlZ3RbikPZ3z7t0h2xrNF+i94pXh5+oJIpqECvSUigsM3GRnsfhfIyYJOBSVljHLy3p3zezoYJR
t5C5TTKj/o1FjnPoCf+D2Ep0P/at0UTDfhVV1w9YQTMInp3ypFZKiF7huT0VubxlDi8FKKN20kJB
eh+UiDyE7p4k+iGurBY2U3iBujlF09aNNSuTtzYOtIxG6D75QN1yT86/tfo+hsRxGAAV4qgxbrTX
pVFoZ5FeY4qTpHxxC4fuF5MfpupdcoOhjgALJVX7OECimuAY6K+NGBmlvXa8IyfBh8asidC+SXK5
BJPFmMV2EN39SwqLl0WC3G0ToIFTADCqQAse34dW//zkf6cSSQa17lbUnad83Whiy+VahbStwKMT
Ot37KLaQKccZfk0kGHmN4KOWy1kwwvnxndeWm2yDGhK6b30Rb++Fa0+Cr2ae9gsI2Xy4ClezNkQM
kr5y2nICYMWmDmRXuXVIckHA63J5KYnDy488H6tU48rtwRw2xTED+LLoNLc89JHGoEn65NxJI4n5
Kbwp1U6SAN46Azyba7H8FfMUZwVAT+Vz0IMk+hS9J5v9otFf7LHoy8wPOwVecKTKtnzsW5sIu3ie
CZi5tgsZDu+2rhx92TgcexBlxZRGn1OTARmvCCCmqP0kemu5qnSYXfQqqf9CE9O7Esneb0sEDR29
0xa+nCRW5II/l6LLOgTxK9FRIy/cMbDPECLtxQSxaaxq+NYOg0cbfpoZ9D23UrZgDpEHQPD+Sh6p
g5gH3vVzYSWl9xvLgXIvFQwHBQb8J41aWZUjKlvO4mgctF5Cuw9v4+KxuQozgbfauKY8BhMIQhXl
IO9asIkU31wsR5p4m8npSx503sRePmWJ51Wvdb3OH97z7ePI4qQSZ/YsC374CTbEv3KaixzbGL1/
SXArx9JqdO9U1evfbDzBz9z4OkYBbnBSKIdrA5MdhnZKfgUCiPW7GNAs+yvtN3ofWPWdXCwzogZE
5olonL+brbotwXPTSvhgpTPoD8J0JvNJO5W3cn6Fgx/0XLl+XcFkmWBMmxhxyy7QCWMpABzRBy5+
/RkztVHCvTHwTHYUu1+r9BFTKrn9Fc1qHFMUAkOVhHIENzSGCYOgC66WlbQs+aPgi0/zuNGmxcwN
TqRaeBleUyVwfRQYP+Em153Zlb3uz3mOOvRG/GGxr9TA85TD50y+828Qrlvgudf4cRMFnVLv5/R5
tSvMfYV2rY8VFnDXVU160tpq1H2FtlT/MxU3iFmwsp/GQQNfskdguyVpB03U+qCNxIIMoSx/wpOo
Ury74W6/KMKK1zPXeriSVpHEbhOk250Dkgfyjh2mr5d93bwz5rHUTlt0NbR0vAyEMOcSItuip8r1
M9YSmmy1SYfELlDR883C040dNFbvQy5O1rzOtEy45xduaHiTpqQBRYMFZ+UDbk4tdzVAWg26mUfi
kdBsgFfyi/qdBFRx1AQ0NLZico5OzjsMx6Awj4yPzs3KVX9J0pNTRq52wB0bh5o1u8ikiqn+LyGa
FxEDeyZ6MqPmT6KvPDJNpiT1Epifgl+d5DMwj6iVgkxp53JM087y4msieFm9jinVtw+8OtChiW3X
cF46mEXujuySPvZL9Cus3YixaqeUH7F5mqFZiOIIcVom5F3hn9JqCcgY9CEQfwl/2cOC56pp+WXw
G0QFhqbX6WRXNRL4289Tfks7KE7nXUjSEQqVEY72IA0Ko+0vwTi2ajBKXU3ZzrQi1iggkrnLfe+4
9j1QSJHR2QAebHQx9uUm5+yOIxsf4XUublMjSs/0b+wW+twgw+41aKIeWRM+4Omo/4Qe8+fBfyx+
HRXC7vWXSuUTln18Q1XYHTKIxVj2iZy5cxzQmpStm9fNStSaApMNQvA9bir/xDTdLnDIq7prYwkr
Hsw0IpN48nvIRUb4Vi5+SwmwjGDJf6x8j4ipr6pEr8FWGoFstp1fOP/6Y0O/4MOrkgnX0nrhlju7
tJ2WDpYy2teQMC5xPLPIzLwy/LfagYAZFH+B6q6qAKwciK+/lnt5yQyOM1e1NepnfDqx8u/S8M+D
z8jQJNytV9db52IUdY0EKfoLCTL1xpE3ShqjLGzk9YNnqdFUu7ZDjCj1EopfW/43f9cTQDUsxIl6
o2jIZROfCO8u8pAxSlUyPka1MgjemaydYJXHWoI1j7gRuDFFR8iFxUhljfkghrdIums7Wz85HwJ5
653uTTlGm5hjBtuGzS02UPjk4Cpfb6CtJSa2y+9dXzbTx1WHqalIUF26IJElFR6Dr8wwyNtg1eH2
dn7AkYy5nZ0D7uiON7xG4HFJzBl9ShK3Er3PKtfe2It+E9eWTjTNzw9eG71zi+wzeJlm7qKtJJB/
Jxfw2Pge14N7OllR2j6c6p4+8D5Yux2qrHah1VENe9lLB6Kl2aXf8svdshcXtXB5U/TFvZviFISm
iAgoB1vwUpslmgtGzm0XfeP8CbHhUty4HA6WpCYD9lwa32PElCdn5vuRLG9x8N/MCoaXHrd1UXhc
xuvbDt8PH7M7zR001uPhreIyzXhOhhMCZ78qmS/M0VRava8FVrygVyUsGF61iuT80WX+AZz1SFtI
koUG8h1mw4eFB/7dpXKJWhRTcuJCyuC4fQzLPuP7f/inC7FqeBQIPlApchE24t00N98zEXWqO4lT
01zg9hMIxzTBza2SDKNnZdDVv6KUHzfucKR5FjY6sn6mIz3UxUM69hwsq4JwdxKJXHQGBD60C+BH
RoODtDwpJDERx4ocZzroIHUNwBb6//WhNZe6dp+lKEd3B6DexLCP83LZntgRrU1jufUkxNUhQZYp
nV9Ek8Idf4OmSqLYK7EvF0UVk+55sFlzuk476/9yshOnbQM43cFJ6bAnMywm2wnthAEPBWgLU+Rp
S1VOZTv06QZ+U2W3ty7ufMHZnwfrwkUtRkdNjZ901Z2gC6fRlGz6hakcwjkmm0JVdXPpOM7ATBbo
hSjC2jOFHP71cSFXHDT7QwiDjfOe7KwydHADCquiFujUT7fi6UGIdwA1BmOZys/sss5lkzQft5AZ
jOW1iwklZC/2xltczR0gnWhenJrGZ1B4YNJemhxbvtKtoI3XEgelqA4NeArUZ7f52UfGXCsV0If4
orj5e/YssRU3pk/pD6ddbvT/bggXxnuRc8ZHC88hIkeeq7btr5tuw3OkwJJUQmdY8E4J31iIta7l
rXaDzYDP3Rf47gY0Tr+xq/0530QJuhuPs7Afj9FN8VOm1Wz5Ad9kl8ShXersW4eo5H7zFRXHPaGn
suhK4NbHHMclw8OidYg1ncCIhgGEsqV+aOoDzh7aeT1f+eVGDSq61PNmpLSbytCenmahwP3ssUjt
2rD7naHri61kB5gQH9DG4sdepy42XiGZmNMQYzduPtT6yGcORk5CttttyXcZZRL/N1u5IcE9s+fk
DXPXnGTIEwBHDxU064+bOrusqSBxy2be+dYb1UxjgBYjsBtDvg7v9cglqXHgwRiFvWdFrpz4PzYx
J4gpmN84XFf/hG1D762JNOcAE+73yx4Z2dK8Y23R8+rhtK1Bn9wklLuSdWnjtecO+QAEwpGgnF2X
96YE7VAAhxz8noKVBpOl1MFntVMXBNS0sUAKlzSlKkMOGOexZ56o/PgRZP/S5MMUE2eCkRGQY/eH
OOj0ZmrxclHXb58pf5hIeeYU5c3wRe5gyp83O/DVjjyb2UxRh1uC2DjBOQpr2L1UsqlQbg9tf6j3
p7r/YplnR4pj6uwaGiAeVrjD0RXxzlOvPjhOpYzsyEQ+Yh9zlnwlsC3BAzRUs2ZHVvovO0rIwzp9
Igx7YjHPvy/wPzaAZy1yo+SQ71p4/vyuZskxNpWD23Ka5vAqio4Kc0uzdN4/gqdnkPHY7CCHFi3W
p4jBYMm2ym1+Am7OgpaV2vSeL+oKe5ANFoNL2oRchIAvwsxswoctCSuslfYo7JdVcSmvKaIFiDQw
oZio/7AtsTpUuB734+NwZCMm6/mChYsNswLjfSTkScV7CqlFQOnBliaQCPfZICemtAqYiijH79/P
JrjM+ldIyZzhtbWU9s6nX4wjzVEQ0VytASM9Th9t2poxbstMIDDAXfJKkvnz1Zyw+eqibCl80Yze
AjuY0T9PpnpRbqnnoEcWhi4tKkvi15Cgvw6Z9V7pAeo+ydCImByB4r5WmhobsrvGp2jMG6KnMhhF
/XtPBEOad4MSVO969R22fFKrlx0fthY0byCskuCTQmezXFhyVCP4XIDQnSCmZ1o/MzFFM8SBmLD0
PbxKW1Jo68aHZVoBJXUS1E0Q0ltlO8goZXcnXgq4NW1RkuShbqzs9LPIUYA6u/MrYg6u/DxAfSlp
dSO1VGlDjNYkV9PmgkyWvRfH2B4ZmZJrcNSwLT9QcneotP/vwmU3JSlUOOuMn8eu37tr5O6VwXps
W7RgGFtV4ajEXQR4PeqoteETIFL8fvMWMGouqoagAkBmilAgF0he6vp5a+pItDtpAYlgV0TmqJPq
q+XtnG+9VGtVaMHx1avLXm8MXknKdkIc/edzlFhcE+qEZmvj6U2NOFmfjFYu6n00GqQdjXnO9YG9
aMPsxMLvg/fGeZ8BaKwftsYkEZKrU84ACzBo2FUdVpkEv7W/PhvoAZySqaRuPlZj98tmSDDACSqy
NCev1S+GXNCRQVvBT76ePJqqsgQJfGJY3G9njRYJjyHu7wFWDqHkVzueObhXmw1SjXB3RwMA5tK1
dwQIboU/rGDqTrzOwIvGGCgqgJbpIT2ycmB4ER7QtygbD1/bnCtw4uwr1r52tR7k/Iv2UF5ZLGav
JofvaCe5V37lGsWXeqwgJCnRV6e8eXQk5SKldhF7dUQD7YSPTBfRY2oeVsUS3CDb63D5lOSPsE8c
Oh2LbLINq44+SdERfs5uQaqqMi4VzAvXCp4cTzL/XNeLpg5ESBnXqV+DFr1f0ab/zAB9M/k0wRqY
4KKuCdmWVCyqrDedHT8D4tIMnJjR1YbrmdI2s+Gs8SbNcw2D0wuyNbW3tX1VReFNJ2pHtnp9GE3A
CBeGJ+umpW6EpAKVi585NAktAVvtms/P33kgiiNDxBQEyBwDeUn/fJqrCPpNi0B9Ttc3Tw/dLDAt
pF5TSHau7+ZbBAIzw/U8eEhsIWUhED+Es4Ioqazb5la2KlLB4OWoApHlidTMBWFRvXaOVAvpKDjy
PfkQdlnXyxzYdTp3URMqoXY8vRLxPRUQBvH1W/z58sllEO26RhjMa2oyT7rRN/kNyGuilrqT1iLS
mbDgy15rMVxzBuhxGnpkUmygC5fa41PqKADk/Q1Ipo+YNuHHqN3GXIsX+Q7xb54iXNrTmEnjGn6A
PfXAzgRwASsgn+AyFHfJWLhbexHfHEePdVXqzHTU1v5xnLEmlU9Ghm85Zxpcg/+EuNaYevhFq4Ou
aa4x/7hB45o0quaiFm+gdBuzQWdrx8AYTodg2EAmSQn/ziXTqwAd+mLR6zqkrAINJujx6/wB9Bvp
BmEMwTR1BCjoKcQsKtt9I+dif8hUab/Q5wLC3/45fx2VPRCbNRc0gKb57dOOytKfM+r1JKhExROd
GOSMeD2Ql2kZecP1xWHR/Doac0pZFtdbYqoNPojUPRvFkSH7p/wMkJhO+9WyEvek8p4q1FL45CE8
Tl1YOSpVWekPHmKjF9596gsFfV/1Q7PrG+fJri4EmfrqodQyeEHXBCxPBf2bfh/OE0byMTevWHL4
dFBEdK2jA4IhP2X92vMPCOMx2koT61qMZQGvmHbhGB9zFOS5AB08DOhEgP5FKOBYFXxF9378yZD3
YoF+FWMoA+zclXEFcHfPosN/IzAk+zWNXK0O0PfhJSh/e9kU3U24FWbEOik+ZRsMLKjxZcc1tEs8
Ymtoy6w/mx+VQEHyIONf1XGoYYWzUCMeQoT5eFOx6rP3tny1LOHmg4i0O4lbRjdosxcPIZLq3EaT
aC7X8Z3hnsRmHjZuTFVJky6NH651dOhVf/1xscbeESYZdiM+N6+LUQ5Q9OG5WENbOcM5YCEJUGCM
W1OuvYwejSjqYRLSRf1NFB0pHBhPPCUVirhDWo84d8gl1LJrxwOT7zp8UNZlS0v5yy2+R0A5JNPy
G6eCZbY1rKA2G3rgn+X8G1bkfhpWfT9sF/k/VCJiDELXIPBllCQPPZ24dA41ZXbbqNSKziy0MX2C
L1hqVWN0v6yas4PsJLPwt4z1Bi/gdnq54fZgbS2GedFrxFcIQpz/RJuYoJyP/71pKQs74VsiRh+L
o66SmGwjOHyK9MXf2lQ1IKG/EJm/NJnveY7GADWj7THleufciJ7oKzpZ7CdoUZ4ysqO3zxAW4wby
4HEJNtM+pPM+edR3K2JJzd++7YwSMLqerD3W1ZT+ayueqn1ZYdqWMeH/ESHGHKCy6VY2LS6KTRcO
fLWCUYUorxAi4VeJk1EqXFQRaBtPONoudXGQGorLxsFluRfwhjhTJPux2qU96R4QSU06PfJCQwL0
KKzwxTyRNSiUZCb/P5mZuDbjabFQuMlazSAUghXNFSuIY72CuETzXIm4G0L/HyoiGenbjRVCWjDD
bTwKJ7LLxO8E1iq0yNBrMNpTFvfgQsYriEHceHGEDpvX6QLL+b2ZSQCWpNBBlbENhWxaw6jTbHM9
ruG76eCNY1HdXaXAde70yfoN5GL6vOudzSvwLzV4XxIEk79FsmnK6wTF+MVMFUGxDzGforTKN0Ld
66fGpfCPkV/J//rZhdW40ZfNYPBLDwf6GHo6krfqtBWR46FlGLa4M/TJjnl1MPWTDY+65HOFeLL+
nsfp6jG09vMnSwur9WGVdaTiwUL0YHoHpEbHSJGWns8Pb7hr78RnvGFrurSs5NI58h6rNvnrQz+s
nWSfSqDrGf2XF6rtLwq5wLcsg9epsOyhLCKBSO3cdQPjuF4lBzqGK0VSJNoaJo4eGe3ekuhDHkN0
NLkDE37oXO1jcFhPNBZRGXk9dDiRmY3B72Svch8lrlDy0XlPQnbXXfKw6oP9rSfqrHKlcSznDYtx
frxMWfbM394e7iUSwqyzAGLcGYdYItzqlW+GyVI3EFDWhXTBF6rUx/AqxWzjzK1udWzKZwwsGb+9
K5xvGp9I+m7l17YZmxdG+A1RLKs8wMoiuarqdF7mWgB57TIy3SnTsn/nF1JVSkY3cxvVBeaUXEET
ilYzJc4Q6LMAWkgyEjyw+06Iv12dmRkvK3fo1x7aMK/lN6P7iYbcdXCAd/MI437p99LWxPR8avlL
dtwuuNIq/cYsK7lkpiw6tUETk3f8Oxn7kOqiarimjPJv/Bmt2JAGyUpXdc0KYZPnzlpwtHB/NZWR
rDhuxeLogt0+gVe8x7/uakDFaVWY1ms2yO2LU5+Qq6FNoFDwZ7L19CxZtZC2cJMv1+UYxkfqBIfH
ahMsnIYO6cvPH/dSTSOlQXd706dAsGGTayKq3Wx7Qgw9SepmBSsV9VKwDUjffAWKQx5tOGRWzEhS
pl/2ZJOWHookemxfd/4BioMYte2IxILEtJYAvRaMbimx4noHmgAB8pp0OJZvJJWTXBZJcvLQmmK6
kcIcIoXNJxu5fJQ6iilDW5WGSywFZLPLdi8I4aiaefeptO+Cqs8WHLG8vyYuHSMIkKBhMLvSpG4n
4TaJe7dsjTFlh36ZzMCASzWE46QI660XJDc2uPfEAOfN3cQlqs+S7SdKpiezM8aaSBCj2cpBqpK/
/hzbGEHD62GZYlGA1+Us+CPUpJ0AS+tlzVMcC/wAM0yn+ibrg8h57Wn0ICbkpPhI5vimHxGwBOod
zQzRaVluSmj2LYt1MXRoVHk98FrRpidmlZqYfWQld0yIQ2zJ8ted8ITXoSjnj3LUemaqxGKRRFuR
ei0/muiOtfbO0+Z0TmORK+ENu3swAsFJ76ugTP6hSnGRPoQjFE7UfH8RW8QcRnHkq04Ci9AgzcCI
U3t8JClpjn5IxT5KLjupbgwSz0wonjqEqIjOXbjxCAQD/pmXhTCtRpsMQrKXlq5BGt00VwkaaA5Y
hz34RKdOGS99w7hcbyjNKhVDJkf+uulaRkvOUFrCihHcMhGxJYPrvGEe+mq4ZHXQd8GhC4narr2/
JpzWKowL/iNffurQLHLINUU9HGT19H6UpeLgYgq3KEyn4HbrhxDyfJTNBkvkgHalh8QVD2X1gEIW
mA24HfzDkERxMI5ARzShnFqjaq4g0gTTgxy3H1OwdIbMek36jAJc31XLGu/YDXj4O+UW9gaMm68u
oDelYCXTYBH+D5z2gHpzSTX9gyQ8J85QOA9Q0KXlLIeXqMitwuftIxCl0+mJuO6D+mvn3UucIr62
ipHXjzdAiN/T1ZvUsinu2RMNaifLCzTqf54tGPlLaPCeSDMwvMy63RuaNZpcCt3WPQc9xt5P39i6
EpUl8wxhiqf2HiqNAhX6K7I6nscss4b9fnWgniOPYmI2qyWcsE4MjDhoJ89YU/0AnE2V3eGLoZKU
dOLEbEz4rNizEPKvq7P48yd/GN0h6C2NePX1TRGcBS7A/WaqF0tMajoXdVE0ccBTrGAbRLoysW6v
DQMJalL7dsQVmELLiEn7s/8a11Bln1plPJeakJW57wcYX5HEWBWcDJyVZXv57TGBWRzR6BfIbo8c
m3Ss+rpCR78NW8mbYzAjAXnn/oLh9D60rcQxaMTJwH+t6WXzPM2op+dGh+fTS1cJE5vWwDr7a7/N
oX9evgZ8ibulzvVdRxWrdud8bxl+U88g8uNW4bYZbwLXWfpS+nre5i+qV6pjVjFIU/s4xHVmYzUA
H1JjTNzWbZDlXz/wUDsBAWvwtn+jslxBBxcHr8YzvOleRrj5z74Y6D0O6ps1xKOPi7bAOC/1tA4u
BJjdTViIpGguxoQ0TMmn7djj2O2Ks3cCMmEx/aRvEsIKI7CWToojRobJg+ssxH+6W3gFbPHKR8b+
xcn9MuP/MOzbMYTPMiTFuoWyrYKQiw9DzB7VdZDrucsGhsIH/Y4OzgxjaHfIF/SKWqP/PyfTERUH
K7VCUKMCPl5Tq3arWiRF7nuTlIn2qdpSIZaiGoQtJ2qbXQ8Ux8TqEyJQGkf8XSbBwY2E8kWcFAN0
hgmnGlrLoEzkbq+iXAHgiDAxJmmckM/7LUfFCjcQZgwiw232JZzGxzr+OuE6OcnPXxrxgWIKvTbM
7E7h1nn9AkPrN4l87UJwzEOagqt8w35M/cwPwBBDxE20Ex74tpwswTsCpNe7+sw6f2mZwdzllpce
UYHNn2l78XCsoq97q4U7/jVq73vghZ49DmZ1d8bnw4meTOJSWvP/Re+SckpGyNU4Z4mT/nRJQ2q6
bUO3KYrFUnyNmdXAP9ylG80LtMpqCdKudDGkjypWhjaBXPSdEHQuqiWYKQLwbDvmXwN+3TVvHFGO
B/lD1ogsYt8wD2u1w4PkFQPAurEYym+8DZX93cA767KKjPpKQoutEIUWCxjFV473yKruYpqOohVU
j4TPDk23TrAIYCjqdl+ca3WaOq6HmbvghLD5gVCvuvSilybSjWmmedeKWKmWLec/MK2cG2vxnrXZ
WbMseRtgwKDvwwHPmc7e6SATSQwshDGnROu8hJvuZmZ7lCPCoWOWIl9LdelUQwVgZpYTTz9ADrq8
fJiZTsMYOYgBZpdKBUg8W4ekSLG1KHtX2TN3sbIe734Z6Q+5fZKeAJ0lkCdcE4zBiIJJJQBxXgyl
6J6hxTQGzV7xgQdDRVo/o++XCEjCOYjFZ++VDHfSgGPZUFskx22KJFpYUPjeFIUA0+nai/op7Ot3
vbeXn/BzNHlzYr0+3HcfbOLASIiS1TUfwWihIMQorfBJLXT7f+sOnHMSP+CeZgF/A3tIJ/bU0cot
LQZIBNeJvSbMP0JlaThpXy1UngmkSjI9Xe131Uzl+GIYkbv/H8W4SdC4qEgUeAj4PZig7Rlmop7S
QHqkHu4V/6+OKieQrGFwfickHPtzgxsfXUWmVfxlAwtD/026MFNwW/9+VsLyJTXHi20rkXlPVjam
5w2qAyRn7rvsimv407VR7+ibmfM8C/eKzdiYqdHFFXR79tGNJMSuM3haXlZV7I4kM/Ju1FLIE0n+
M0wn9WqGpPBW4pBVA0lQ0dfvxwVXWDHFrt6qqxwvjwYQ7CM/VCNDNkmstOOBn9pt3+oIqFv2+j0n
GswTaSHbyFoUbqiB98RUXDhHdcpUW8/IaLP3/mdllCDdlGzWp/q1l0xvcqpYsCwQCZlEBq1hBqFJ
fyPoQDf5f4D8HGyPPUaBWLoIN86fOXAWWIfTYWviffjmnmAeyHtvJok8CN7KDvk/Lg/6gyEcE+aI
DLteq2wCHIdMv+WkdIkDDh0cZ6Tb++kWqOCNMQu7SGpC5B3e8NGlTDnLS/YrMI/U7quahBc1Soqv
Ha6zo4ubpM9CshJKPaWCdiAx9QAjqcIiIXsHQnQ0H514Vt5KoKKEZmyvdqAkDZpjHFfFw3Agahow
GlCK76O7V/1PIEEzeDwNZQj/Do2YrxSrG5qjeQjp0yFirgJEhbPAd9RuKq9kfPFOo45xBMDxpCWT
qFWCL6jWMQBqnD8qPyOm8Wt2UiM9upwUCheAaRw2b8YxxwC0WKmHEp1QWEQT/jZ1x8ZylRKDALTE
PYVHmByDGmAK9nFHWWGBPwRe6BXbuAzkDKR8v1F3SPehoQ7acW2tfTT9EbMmAuKEx4Vh74CGpTZY
qTvRbTF2uvUzFzsojS14bYMdm4KOD/znQ03kFTF6EB+Anog0iG+bLWUEZWKczkjDmAfJupWmeg/2
olFk+TFCRgufPXCF6pU3fyoAE5OugcnQdFJdl/Ud73GtpId6v5+Qv4Bjjgksbzmd21heqSq5SEIM
LUyeDk8OVcwJTnU7o9QZIHRAU3FsZk0fuH3uYRqsiT5Ly8HgwMkoZmLSujY6leI7Z9k7scawJ44P
orh4zPsCQ438g62C9mbtgDUd5eVgB7wcaP2pw5cjvmHxHz7qwC+zwZgXFTlzZYvy8sLhCzMcFU2+
LrSmeRXUqcSxEMxJM/7tBCA13dCXBTbi55uQB+qC9aawU9INPZLQ0udBPFZ/3EikK4c3twu3pEMN
bJuvIVdwXf9obyswzIdBII0ofy2FGmVs4ZWraVliC+CVzqBV4vacw0xZKT40ic+0oazNopWBCnGF
kIsYOjECDERzrX/V4Mn9XJWs5BCQ/C+M65fnvz6818telBAZ9cJVs2ZqP/Py+k6Pox+8123TwRoQ
8uiyRTd43xO/dFNK4fnRYGBbBF0Rs9ziLghgYL7TA9HnkKH06d3jQJVyF3sSXqvv0Zfss+8tcT8Y
MO44HBK/Oa7hvEr+DoYrW17063V/5OY9BMMRkgl5nbrpEARUcDE21JzBZemsViwKbXIz8pONXgwi
K5I2aj62IZKLYs4qFeVZZj9UBDL7Y9B/TsXW4D22R1doCyJu2Q5MCxw5KTHYG3psvYHCiC4oaQQa
57bzpuqa+faJ1DkogP5yyL3Oj7L6EDo10x4X3vjpkLFCeyEt0iEMEHq8LDxsAeVDpJBNpiK8Z4VJ
A0HiWgT6jUuKEUVeqaVRnU02ZuBmq+FB2vKpM3XuQNV05/jablONmvRn2ccSIwaIEdxZU9F2RNzw
wPexocepB5ZlfEp6UoL5iVFcmrb5o9t4nCCNmNA7G9gP2CipAQC/gqiemFyz7FkZ56BITXVpCGfV
m7zC38wNGE/fuauRDmouhwHpbef24T8HlOZOJW3AdGpkv3BZCnq9+1D9EKCw+CrnUN+661sRN4Ju
BMZ7p2/eIK1UYK02k3CKYYXy2f5kbuT8YPk2Zyl+bIgAHzvHgLiwjJ/Li+hSw9gF8smiHSl/yqqF
i8jm0s97mMcXz07g3nm7Zf58kNHKM0D2EY1DYAYM+BJgZPwqA4/2kfRoKkveRsE/DH/FhhT9KIAH
8iLF3n6vFUj39J9+96FUFYCdEB7H3lJY2IWN/fP5RHl5u3BB79z8Zs/fUsOQPC/n/VaMx5bEuDTH
+sjNzucwZxalluZpF/JzK1umpcqbBIYYM4LUn71WJa32u7evWYnFbMsKx7gXajEtQm9DbPOszQmo
7uXyQLqxhNLnFFhlLKQdM4TtcSxKFI3HZmi0IuEXBSOdJ30xYnCDqC9muAhYs5Ta3Vc0nRRvwVDN
sQio7ZvMjKuXA9VbPOdQz/pEwm1FtgxEGK8vtuIZ1I0gagvyBiyKCY8uJXuZdVu02kh2c4UeK0qX
yqpMKZAe5yl4Uv8R6IjoRaOZzWPJqOIqECDrZv4Rl+8Mh6M9PTv9FKM9tJonAKnDBnRqL3zyROIV
2jS+1f0qpqs6XdtRJ9Qy0y0S7QDbhhf77B1a8Cdif+f0PIXExRi2ndmtROPKjkHtak/7vZ/ZhaP0
mhsLmQbhmtv12XQwyxCrmKpn+FLQs2GxNRvNk1MMScek5D/N0op5hKVc11tn04vJdOubvfNwsHvz
w2qJxtkL/IwdtTngn00zkdW2ugjO/aYpUk0p++J+jTdYiNACwQ6U6hJ4v26bsX74iqnvIMJ5Pmvl
z+IW42/bPWxhzrnmnFsfyAkHqQCdvuMS7ZBUdt54qMFi3QtCpuLlBJHWv7x9/r0bSeuEUcH0pirX
JzCksVqOgJEzF3RntbblEr4GCVh4AJcAgPEYPy1POFoFreHP2kubSY7Gi1NK/iBWVrkgTm7WHKQz
xcMa+ZJZaKUdHR0kao3fLAH7/ss8khrE9zZkLSocLUh9fwzpJzM/CZsB3kTNbVciVg5mrHBJ3Rm5
8FIqI7gpji55fyd4NJrbv5j1ksTc1NLjaH0vHmlK0yJ06qvgvfvLOJMMSepGU0w+j4e3LkrmYjO1
hAT4oWCJOVXMwtS+XHEEta/q4J9lnM95WSKFyhKhglXONWjfoEJ7v7NOIBHTlarSo8fmWWnvJTnv
aJDdUf2kUizYeMGVTiiZa2Slt2RqfMD2RBCM1HfQ/ammPQ1vWo7rexit6aNLyY+e/Sfj5s7CzT+F
tw500abFNGnUB/LIZCp6T6g1/+GzOi3793Ukvz7ln1odG/DCNBHIdbVa4xeewWECJOcy78Cyie2R
jzdIapajjK38PI1TgCY9cf2FopfKJ7uXafcmnFpLpF47D2iU8o372JG3JEEstaNxnDFQioW7ZGcu
a1Af2oKrqoQB9ethzmdJp07FbvHi1FmCvuwRZFYurhaFmGbUBweUZscldHRIHoqlxx8hwE63Xfs8
CV8ctAgD+BZ1z4lGg4qJkW+DuW13U7+FhleH7MGOw8WzchELcJKnsO9DfqpuRXOAOmNASsjmcSWM
Agss7JH2D91c25zuV/t45yN4bXWCGOXNDfz3jZqf3jJNh3FbiOv180JDKBTp/Yd2CRxl8Zi40nAK
bOumQ7rBocnKX3z3qpDfCfx/0S8hhhRlefRw/yrE5Ri66d7aL18Yo1xU9T50cZbHKGX63l/JNrPE
fqyChZe0Mq0FjTjblfBX3TwPHAzxDklE7m/SB2Zg43+//2schAN9i3gG8625ZQFnQD3Np+I8mJvk
qphjTsBGR3bZjcj5CxZ0t1P15d8fpJ1GwO+F6TylHhWObADqTnjCjUJ+gZEhQbSX7hc/MHiNpdfV
XpQcLj/5uaYWjIfpyQsFsO4fbEhc3V3zJxKZ0ZzldAn0YPEGYFtRemBLa+kbFOqP4SpUvQHpkx8A
gftuyR5LM+/pl/hjpb8V6SZBAcGMoch8G8+KkV3hAbRGXSsJLHJ2vIm9SOrcaiY/HwwVPzK4Z+23
pdBTFN+rhfGt+diExOSd4rikB+Cc6740tNhgXCTK3lDI2C6UclkpGhHcRISwe0HTU5Nf1Y5vpEHw
/U53Lkpkyjb5K7PvYmiiLXzoLHmDOdf0xVcqKhJn6pOXFrDjE5qWA1o9avM40TvhX8YH68XNh4zN
n80VcMRAzk2UWVYFFG2sPStt44BuUtAQGmGNd3LGdL4LcpznYoVtcWc8YDdgvkTfNTsd+jMUrXTZ
d/qi0V5qs0UT1wTdemnDvdMlTzYBNWZhYcYUwuc/2H1tvYcp6ip5gaYVyGN1wMGKjZ6wAHhwWn72
+ahyRVmm8AToOpWGjrxlRynkgXJn104eNQ3aCBVz7AavLdNIIjORsmw+zvk2gFZA1nf+djMOpczK
PneJnuGpcqTF4z5yMHy/mCbbkoN/My6JV9NNcb6D8nSo7ROxUQuvmBt/jTlmEUSRAfT1M1FgLga9
vdaEBBwn0GZF/Tn3/77nfvk3Drjz6GhY6XRMUfdrz3q1NTpjbrqbENVTUmG7pdZ/fxB0bdsRrM7d
gNNCqjtUqocwNK9ZnZJ7njFSmGs/NtyuYguHmdOrXYE7Ur/4aiXvYcxeI3O8r4xG5T8C+VBN7UW1
W9WJa4Xsfw9Q59YTwmDP/3Eed79x5pnMl610oDJLym+COBDWiNHoAPJDU486gwuRzQ5YUanObRdm
vcZc0FSCpUdkH+F9qtbOcw72nK64zKG3+YDfZUfJANhiv9fjmNhMCeJp3+/ovwgtl79S4uxjXgBh
Xz9An1lnWnIYVnoxl4WWzlOP3iKCQLUgtzmC1HH9JDbXq6tCIKJrg3vhRTP7DwWsd6+D7bfHnBtj
z9SnALlhZ5MABbQ7BmRQhOAmtkl14v66/5QSM5EPcVN9wDMqkl8eqr1cBVuTEplZJGCDFih1Iohv
kJH3ejkk7fNcNxPYRG63hioHusiFRdBbsQ4zMeQlwPbu/S8JbWRjiswLri0H92eQ31YDSguZDqfm
4lXyacak1TrbaoRDMn2MqSGqxljU/GVet56X4tqwU2ZVsSTMXuFBT5IWvKJQ3EztT1n22y/RdIsp
yfhdJEzkicnN1ld+MIWYzu29nNlQl3J9GjCLFeZCumsqWAWgw1kEiqMJbccm/Jc9saIPNfxeSsTc
cLIpAURK5rj9RkBRHF/vt2vOQSWynEsZYpYTvXLOlYW2Oh7oEhuv4ZctbQ2uaUUELF/wrACIzZs/
TG3dF0PFywgV+Cdon1uXxMI+Y7Gh8yz7GerbAIQD6TEfJoTWC6cvZm59V8WqeE/unwVj1M+DX9ss
qOXE6V65z5N0OnDg4OZCWTDkC/AtcSJr6CyD0CksJN39eugsH2vQooMGf5GaVNWKARi56dz2oUJs
yN0kX/Kx18iI9uVn6BE2V/wsZRbbn9ZZ02D+HthOMkS/sTAvIr7ndV+93EB7vC6wq1GM42sWaHSU
A1kDCXjUBMMQQfm6GApeT5JHMR4rFIkc3Lcl54eqm4WRlwai9BP7NmJQrK1qGA8yuTLhx9cbWLxO
4wxQzZ/hKoCYYbGC+Ow6ab2Qbzx5lmaBfARUtDfrofvmaUtQx9bsGrfg9iEHoFQPt3gBPyCF/rl5
dpxoGzuPpRgKEh7VI7fV4I7hyVj87YPhluYxqnS0AkcsHQsAp1nkesWXvIaFhlhutLmN2QgKnPDW
e/N7sEFYobWG5nO7kx0+M29uCEyLntfGGBS9VAZfydTSZygIlUc4bSLEwK+DCofiwx00rgjToYTu
LMNH/HiO5ivi+drhEWwb5aMyaV9FXWgYjUrS9H5FUvzvI3+bmP2km1HYOTrGDFhkYO87TfQtKtRP
cGEUcgrvat7M2gZBY2KWNMzk0k1Y+0XXir6rvYL/NSK5mjZfNljmxwBOW0Ie8EUanfbRnr7pzT6N
o4jc+hQ5foFcQe8AXkRNOLkhixsL+7fMZ48qAan36HIKYuK02f6rD/PKl3BlvntT2ruX1Z3jiq7f
1mf2/2mJBvmMcyGYsAVEa6g6lMdSnyYHgfNCDNzmuXAMXfztV0oxhdKCYE6j63bpBWzhqWxXru+2
NnVcpww3Aim3wSojEAGIZJoQgyOIwmBhOnMYloTsYB+7oxNf/T//cRPtOQSrmdDR+APsXPQsmFjC
rwBjzJhIWBfKm7Sv8Uqm6tz/agojpHkTaEnuRTtPMqQ3xZ61jUT11sStzXEVo5Ehi6UFz2fETNqc
Szadaej+pN3nijxECupYiLZhYof+p7pZaoJKuEJ1XdNG3y6BTG2Sh5cdb6F4Zh4p11jHUCfLlBAy
t5axAWvJkTic7qCZlbg310OfhxRJvq5s/lrIPS5pWIPfpEutzcUSyZWeMC5WmwSHyX01SvHha6aP
6w8PABt2eD6kdc9HG4KMWy5dLQ/YnHUxG5YD7xV1xr1SSE7u9CdirYY1FnLmt/cMOtOlg2MSh5re
hvWDQ5znXowo4hXOciHtY3GKUW+DOMPrODtE+h+i5oefMrMF/JkEzJogGB2TjI2qmgx/pp8IOlHR
ZU+dx1tFssKwEn1YGRQee00x82nnbnM2nY5k86GljT3YLGALpb26IO1YWPbYMO23YAmu7ZcuVvF9
Csp/OjzSpNTTfB7U6B/eLlWIEZIwiR/67LcdCF0JH1Vz1kjexaShxO5v1ukG2tDREn11EfHQKX2/
uBCoCNgdUTckI7XDZzlHuv+PswPElvdiWxPffizBLd0/RbEPCHdAG0OaKWf2Q4hYPkL6We8f6a7X
NfhH7t7xuEIkLL3n5XxNIRjZvkVBKmWUdOO171n8vg4jNbLB507M3KdL8G1GlZGQiaCLRe2sWSbI
SXjYrJ0wwW5viok770WaWRJlrp0CZODzJWKPjDw48gaEbTfQSiTs0N2WzeO75p+Ee6S3/S+nxJtm
3V+hKgjd2fe2xtDXafBh2vZ46MvfpmCvaZND+0dnmupc145/CIj+iOi0emTzInKDVudZilMA6S7Z
oA1y+oSAJfDzq8U+xG8r89yl44uhEbTtIER+Rz78hgJn+xJXJ0Qn1V1vZ61WGQrDEnJfKJEn6fjC
HqN4cxit+LWq6BA5YtqXqU9F2+BgYxGlPBfmoN5/WlABkcPLvRUBRlWQPHcuMOnM25Od3fQRxOZn
38Q/csWe98VwMTHF+88wqgrBbfqqc6Jcz25jBvMRZS6AAUHWWkJE61bQP9r8PYOLwC6TZCf2sIMG
70+2MeJAopla5OAfGLZYWmQ4HAVUPs+xmeK+FLszxAc0XFtJj1OCGnhZ2hbwM3jdWWjbZxrzwAFC
nq7W+9zBBjgy0sRBUfjmwcSchA7QsGWE/BJWTSGHRo1m27t62M1WKMGNnuOneg7nDebsNJ6uK017
NtEL/4Jja4kwWyqRSa+/+PK/3Ioz3yXNhCMVwK43iG812XgZ97LS3vRx18UzYjhfYZRC5LJURObs
YGSdqgHruwb5vhRLyUDp+uXAGF9YMmSmdGDaBVO9DF98RraK9cixpr0hWvIdB9b4/tXui7sjR9yG
q/pI0pW696z7+DWx4tRsy8p/9d1OcLY8lBH3wZHILxgSoCE6IRDQUCgFPc8Gy9RsjZ4vh/UT+dOK
WdTC6G3C+lrUaDiMDUBnC2UmezMFjFdnt5570OKcWxiqboY/lKkzhwOJzF1mDUs6B//xJuQYpseJ
dNyPQ7ClV8qlxTml4tZCcPRc8WtBJWGGsGxRCzRwAhcW7stD7Gqo9ua7dEXCdQ5FSqVeqj63wc/E
+h0uVE9O7RXuEK9Fa3QHud+uCKrbYOQzJ9bwBQJRGaDP0q+BYIYKySgYiyXyUzUnRIWuZo8/3kxH
WX4cEaDNzDu0vS7TBqDctCWyyiqlgHqf0qMWbjikh+XT4yENeDQ/hUUAHkyb4Zf7LNAsi4IrPdE0
aBgDj4FFTubqhQh0JoMlOIZpqPl+dJPGNMs+D7bSgN/Exhj3gtgAO7fyPFiq9jI+luOPiaZpkcpU
bcyrv4JvPpUbdJdlPOkqSIE5Y2B40pZaArjLuAw4NTv/H20IHPEElD+cXOlSjPMSEXB6fJOmWNA4
YFhMSFysLFzedXUfkrDW+4WPhQcRxOwKp9cfSVLvqX3eioPSElfG//1wX9pmiQaBC3/AngiV9qbx
ny7RbFxaS1UX7Y3WqvGiwoZvaJY9vWL8mSr9Gvv2LiFA28TRPdp9WZAiM2GzpvfGEYXW9y1oaSx4
tapCbt3y5L2h0FJ5rGrJ2Q3v4nUFuogvt4ern1780v+LULjHbaYcvT+ZGKPRLgULDSkVJjz8r4SK
9iLorZ1hIm3ggaZgFpoagcyxwADPI+dOg/i+n62lqwhzjHw07Ctmd2J8PNUxoaAqqPl4gWLDL3vt
AVgSj4IWmWj4uDMPitVzu8gzJ2VrVUOoR1InDe682Wy4h0IX30MyA6qF6nfK8cusGmvDgWt9GCw7
fksRWCkhP+9eS3LzKOF76i8PcF+253rELiRk89D9EnpmqGEeZEmptp8+BIfaKfQdxAOyFdH+A62B
hYigyIQESl4QmqWItVm6QprH37X8YtiweWy1u0Bmowtn5isCEtHrAo234WP1YbKtSbytK/ZI/Frn
UkRCC9nTU/mP/41A5WmxJszSti+kX4A43cwe1fujKh99jHk8y1Ie51snnHBhqFkOriirq8B6ozSx
xsIDNbyVXbGmtXiISgLSVW60O578e1rHcc0Q2DR3rP/sGtXdqkLBUjyAHNXe7BERtYCwbugkKKaS
hpKl4BJ1G+uzxIL4TrJUKTDviNl5SMO849VPmoG08fLz3nMONFGe6VdIDaDG1EZV7xqjQgWa3v5b
alcIpqgBrhhd91SOzH/AFy67l0rOnCeUaz6OlbQ/1o9KQLgL2gm/cilwhFsFpki+UVWPS8Wo4YGb
FY7euy00KSc7fQspzU7QUFZgU0jz+zKVJhdJq4qH/CgbYbrLK91l8/MhW+3yd5mR+tKZwCv/Ic67
vNNa+n8NWUs4IzWAXDRcTHsR7E1JB9kVLWCnImdGyAg3WXTxhx2pCDzIPYLw/TguYoMN25leOEqb
Xlg/LR/37+HJcBqu/9Itr/ws/Gy7DrA1IQgHasbz73voBfsMdvaTZlMtm/pRyeU9AXKcX9RFcQVx
efOzS3OIgqdvPTWJGjq8wZM5YKFoPIoyKfY72CcfuviXFIGoc1bdaUkFEbBzsKoKlm2yvTdP+u1k
nwxRnpSTy3XRz7AQdI3kvPiI6bVBD8IMJoHs0Yziu9z4ddWMa0KdNULjf+7lN/+6CT2nBnnO5zsU
vFt6bwyrLUf+SwBMkOTB44lthjQRYqluJD0uM4DrAKeWIziFpTsRA1a/deK+AjJt1+2tQl9QfYpe
0w5zOrqNacrW8N4gfy8nbKYoStokhNK3cLP3j+thWoec2ertrxjDYB9MhsFUdIOD4AJrU3oX3Hzw
ZG0bDfJKSEKi0RjKoLl0vas6YxFTGwENpgPcWXaO3EyQGL4Z9gom9WhyJicisbfQaH+zUdLCvHBp
kky0aY1WnwJLbVbMQyGowdAamZv29mcMy9iFgLX6sbw1g/JkofYJ1o0ZdCdR8lfTJYkfBP9fPF+i
k4gK5PTNE5b26o0JYBWpPs25cQcse1yNDfW77vh3O3Y0KG9O+5okoI11offTMRAddnlO5Xdl5sZy
g0mMmQO0FYpKcWUaSsp2oWPZQVxg/G0UGzmmPtyN2FNigJ/EXpLy/ntM0YGDHDx7OwMo8nHd1LoG
ecXcJY0TUklr/h0EZUd6KvyyVLnfuXNQ5b2/99PxFMyybT15iFihWg7vkGQUi/l6HeD/PP2ABMaw
3daaPLWlj2N4O7TGX5PlvxHMKEAi5PJHxKvm7clPbXvMs7y1jIOdr4nMo/kR2QQOj5hVGbJNV4EE
+CynSK1YzEZg11Jy2sHUSVw6VoxliJec5XVMWes43mXR5ZuzM/ZTW2g3pp21IHZMI0G/swToqp4P
7/9Ql14Lz7xqskWZKCsWb5rBn6NYwrdP+8nJrza2mxIzwla2OcTSNJIJyjR55YUuZ3jCP9wcM9Kx
Xh3qExWkjm7zK7/YE1wuHq7ebUn4KIgT3dBIf7uSEbIOkSbUDotOT1lZLX8gHJqu3fWzuztGCK1r
/KbfeTMov2eDjPJwoBlzgNB4Vxhk2yevuFMeRpFtEEHErX5ope8IsCWE93cUzJSwew1Nhf84XDA7
EvrXB0WsZQULoyzA9o7DjZqQzPUtMX3vZQMTVe3eyFOI0oYRrFgrNaNqdmN0Nzv3C+Q8eQo+dby6
uiCoCl63jedph/qrIy1FO3tKDeGlRwhxJdGfeZLAkakGM6c10yl8nezNyXgf1crT/me2q5NqFq/z
WepDCgRZIkHBW7wkjPNjl4nifn99OVDpBBS6iegUQDldl9I5C3HrBn7TGV9laJy0nNmg/Wso59Yk
aBm5FgX8xnUoDkzlzecmcnbzv40n/ai7GRPdaTmDtmRd76k3LsxpmIBmrrkuFnzGTlpM+Ystwu7M
diG2WVfF+mcpqLfIUWRqrPDfNtGtpHzVaXtJHo0jrw+ImcZG1arktuqOcnpLKuz/jjGp3NG4grDS
1urjo3VIr9b1V27jDSPnpLi2q4VesptyKry2DxDtYkuZ/hoB94N+6sEqC47nsGhYP8JbkwIPcyaY
gXJraW4HekDPQ9uN0vqTosj2+NrlSS0u6Ljhv+xd4+4EfexEDh/HRqu4UQFV0jOG6Ebuot57cu6V
FzItfjCNxwt/psHv+bx/0FJTdnnFhq4DdjR09QUgeHC5SIIp1P28dKLnSt8mckRJ+botRsNT/dzs
R2zdyCQhVCJP1RE1yIrsCtFrloksydBX1Y8fX1nycq31BHRMjYelHlCa269D0jNNlBFaH6MbgtLI
ogl44+xpR0LlS35Ddm+NZF7/jgxaVxRah5t6Z1ssodLb4BC226dGkuJiXK+fe4HE+PVvvWMe+YkL
cJIEp9fFLrvEE9pAMH9zKkQB80OqvZQnFmqowFDTRUpr4wYnORllCYVknMkJSNrTxSNaAiFpEFi3
kFX4YTOJMjgKwrO6Bydp4HYiyObvbIeNi9ZVECMEWv8f9+uFQIkv4+8yhAe2C2M7SphckntWqFLA
C5d1avvsIQYfPe/V9lTDJbSUG1kwJfqYKG/KAnXunJCYDZaIyHF7SeBVdc1KAGbFydm+Z9PGTP9d
ItKyEdPLIDa3uNZ2WrKvgwutm4YOGChcsOD/fdQCYXViu6EywPpyNA54oGZJnIuAZJ/LQjLW2Mw1
S2GqTzdthi3HL3joaWQsH3BDrOITUndb3bve1VysAw9Ep3ZBCc3rft0pTh4R7zjlkMufdPZy0L6E
p27zwqf2FAMhu/tojIJwMulO4UVc/JgmEIHW74/WyOtaxDbgyqxhUy6XggLsGhqO7FSSKp84S7+p
6eh1myRqMcqgPSpHHQxAs1zWS89hcH7lUASC4UY6qr55gWQPjkPw0u4w/S0WgVGZIkvhGFeUm4BW
6JNJyvosb36Op4NNXItOAdriYHcyG+ZV1Ep6cAAaQ9a9Hz6k+EgQc4GKVTjHPbPFMapoL/zk77lV
uSu2WZnbfPD/YViP4oqLJPzezwcNGHFcheDuNs/4N7VHKFHKEQKpQq2kqvzpEXAp4ohgpFiybjhx
KBm64HKCneoNTvdvqr1J3YhlxGz9JGtTx7Vvhaw3r0v2jtdipZG7yyQoAGqeafoYTveii+r5sE1W
frynKyvY00nJ5KKLwSQ5rNNHeOxEohZbKovne4eg3P9i4vNEecW+2Sd3D0AzqJXG7HaFFo65bW4B
3o7W2Byn7y+W1KzRWX7LCkMnfpEHRIkL6eKtD3AzdtP7655r2nF+idjGtc1CTxBB6/cXD89LVVAc
ILC2js8Tpg3PT88o/UayFkK1AH5UR+bYX9oB1fCBxEF07whN4ifjD0IJ5duunlosEpj0n0VwNGJA
c/L//mEASKYR+WSft0JFwBYhckRhnIy7ZxxPzRzpptv8msLGiTRDyv7BAnYZ5kOOddcDZlILBvbS
azbIpHAdcLu6KbJN9W7t4ghj8KGGB7O/iQi/cTt5ZIPo/1oYquahweAk421pmCCjf0fop46Yuc6q
DusmXCX/wca13K2ydyL6/IbQwz5VscysOJ7KUrHNe/GLsttY2fgghMRq8XOg4d7kWOpwHtdkGE3a
td92JRd4sDvYmUyMW8i03T/AsBO9otYJ6ZAfUjM82Gz74rLLitqw5m4IemUgB9NSddhpSVXxb6yn
U9ca/WBU3xQYkt0+VVApGvULemQTV3XzE0C59y580dou/u6+KoU7gNYbC+kmvVSRNVFRyAgDmQw3
C1GgbPVTnPORP3FDnSdZTZGNFwmC0Lhl1o05jBus6KChOOAamohtUxyk8hSsvXhHxShMG4/SszF3
zqjs+ssSY9hmhnOFf1zGin4fr0YOq46Gaf2kBzpQOQT9ICLnSd6+QQ9bZAC5QY8PO4KzlUMdVmwY
FUtPzAkOXN0Z7D1AsjjW95YeIcqAhLhz3VBvPWeyJPgrEIGn4cCqgHVajGMg7JmJSJFZhzO3cxri
t+s9soIiRNYwhCA49/KHxXleTW5dsTrcEv7hBccnR4QIVoOm3XPcUWPSwIq6FeEkZ73XeC7poy4d
6OoF1m/BvmKxWjcGIfFQ8wnTKGpEjZr9bRW9x2fLDyc8sLjt7QP66DSpuo/LSaPVaa/Mm7pWZLSJ
zSCPmCxFm/EO2Ykgehyg4lnlbQ0GF7TVa18aoEVLJmqFj22osVR1C4C9gE4cRJeaiVdD3Zhc8sw3
d/kR3oErcMg8KpL3QEx8c2FvTd2QFtsV7RmG9K5Usg5n//CDuCY/srhFBCwYTTrrlbWC0PLmV5KS
isE5JrJESYDhGuXt37xUBz1QqmwigQ0ixI/FqUZUWo0fYaj92mRRxgkT9mfQg2b5wEA8oG/Rn2Su
RpZSuINqxwYPpNd0oMZfIzuJJ+y06bQgNBh5HV0F4Khhy08SdwVKNQ3/kYJrCRDt7LZyAeH0YlxP
9Kn4eMN4OWoU7bzbSerIlJsMSwoD71ZRI+3VBcVUzAurokzfYHW2lh394zBHXzkAlBVuBshtQlc+
lnfU2jPgUoPatPXyc2VsKxwPqqwP2TdqG1paZYEGjF5vB3eR+BZ9HSarBd+f/6CSD+vTcGMsFWlL
iJ8l3QZF7dnlqVoOmsZPhMnHpaYUXBY32XyuCI3nPnpht9WhZW3ilIzRxlz4zX7QKFrtAAwDgLa0
xPa9YA+NVEJCTGwFCgQSOZG/0vGvX/pANf3Kn0hmDHI1aIFbXeXHVls+Ea91ti4LAtjYEvEtwh+H
FFp8Huy57WgUMGVhRVQZVC3kypLt6LRB3AQbeFP7gZaSHHFhRGHEyhU7gBZpYYjV3X/TzsQ9TGwD
rDVhYj9JmjyF3m9MjiEnkJ5N4DrUjL/tOQ7Re3orOg2LSmt6iwD4jwcWNAZybgj3mmRdUZTFaTEw
kz6D2f4Hlpg+3dzunby7tYAYhnfWuU6CMliY7AsWvdFDbLp4vQi3bnOnAPLH902QAbCiwovfdqq0
BR/cwbtXm6cWDISO4K71K3Nx45J/nJwo0GJThV3eglkqYI7GoLxbX28xnBzuao4eypu+AGSCP6E/
tN42LAKY7Mx80RPgzN8zDFCgQX7prbM3jIPnFssYr5ytLO1i1BRoHS0ZaEfnsLZgdgyrp+Jy0dOS
TJPczICtX64LKBckKlgrvhMIY2Reiiv2vwXJjewVPEUazYJpSC32RpuiY4oIe5NluSKw6wPOBzcc
D9S40mMPji7e1htGiQ6DAXAoaIu9JkHp7aD/0qgGn4aFIc5saKysIFRAOY60dHvLGbIBFvLk767F
/GAKmCwVg7/6d+hPabZlVo1UJdFAuEMOoEosWGqvfh1FqbLLZx3WRu/MNlLvds4UXAq+Xyd1KolV
q/ZCS3mp3Bg0pEJbJTCMR7Vp5TbN79/zTmv6UzWRIHVgyTyWl/l+lnYU5wwXWauCA7VIh7BDTGG5
ct79UNl7mtHuv2CuZFhfT2sPfk6zv0gh3VuNBkVJa/nQAF/jFwyIp3+e2df8NLg0jRVxmKQKCrvc
hFA4znaIee+UmOlBB0M6cwP7l90fDITqpoIotpQYtDVvcVwtJazKeznoB4k2vILL/yCmukuoOhh8
TsMcaCCyMMoMqMZEiT93dsEzD/HmenndcZA4USvihGddtxJrFbfRIQyb69mjUqdmXz622RrN1EG9
mBZZ37xCnwrXTnbLyM7D9Qa1i980J1F8dBqmQl20Ld1qGYePsXrFTu72kF0RyPIFIV7kONejXSzZ
T59h6SaxWACBvCgZya0qbACo4HJPenLau+f5mqvGAJvUS/jDQNojGaOO53bLEvlntDBUKDoYrC2A
6gxAkCMpixM7v7GuTT68D2SIGI5L6UQ7/2vV/OnCFI85JoWgFFFi9dc154/MlGFafRjgwFaDm0NJ
/skFOIMk0rfwOpwTWUKL7pZUIUQ4lM7F27zZ9K9iuE5VXWZXhas54DoLzppe6vLsCp3NQahz+QJP
Kf6W89PGQ/7fD4Bmv9hKPcBDWUOjtL4vk/HIabD6fI0SLSI+zgGrIsK+z3fYu/Qsu6KddDWfnt3e
LOiG3G7TRyQNtKNB631el7KVLKL4w+lWTHSWyqiUYg5UmMr2qBolhFy/sFsAGzede/CObnuDOHKc
0j29y8vcDVBi80kJdUN89TtbUVmj/Nnm3jyWSIQcOFTiE9fEb//330vrN77YJPA9IyUSlsDfBC47
tupTvxMhr2ecma+8S2oYEXOBKZRgV3BNhyWfQBpbqX012gPm9aYUXUoFr4+CCfUlbvCNDydjTQvY
m1XJakQ7tY67brieOf7r2Xs0m5AfrSXXwmoy+wffeWz4QUJYqysiENETQeixcOaAyA7yxlh/T1ZA
7tkPAG3aelQJaUNonLCp35+ymJ4GT3WgACvQIzEyYM8C7enuyN1LYd9L571uvd+QINKtcYTiY6v0
c85vIqbExTNDW3GzYlM3KpQGyAP4j44HA4YpuKmTdiLUYoMrCasSYPKec+o8W1bYEvv2kqPWZhtg
xG4fiJNOLFj3GJTaDYPooARhs7aKKgb+z0KxHI7DusIrxq39XVHoIR+cCb3cgHmdMs5Sbk+OOaGt
eKSOoVOqXBnkqju2EwNBSRD8wV5AVKpbF+i9gQg11WRCuagWcdqc+IQ3ZZRwheOE5UDkak1oiWB0
u+aDDiGU20fsZwntBJETakuwdLm2xwxSo7U5EjVKM17wuEejGgXL3Ztn9EJDyxBauIrle2QfNsUe
VIAI09dUJSLp7FtUsrFDH4AB+3H5LNrkY6d4WVNbS6K1dcP6XGfRy4mvJJlHLRPLbx/ltqvIg6BW
m3SMHFm5Kf2avM2tPOUcYLbfr00LyPERUlygUcG1kEHfsZvGpiP7UXGjQVNWXlM4TncmM1/oeIMd
+wLz+oVVmwo8tFY1R0dMTSx9S8AS+LYnJRldrf1kNdnkMRLo9Dcs8NPq+CfOH89W19BwR4VUHs13
Jm2erHicrD6HdxAe/tSFOYXypFkU54e0ybQSDM9a415uyUmlqfrEcafJ8hssJeDi4UXXkZl3LEKK
Px5tqetJiADFBdum73cRsub/0scQJUxd9IntjEOj55rl4zj+XjkEuWDc4hDYIVW58MnGCWPAI8DH
ucayHGCQvYCDwFbZHDfhP6dRqO6ikxaeKTI6dw4Thpw0QbUAQj165YBlcszm2H89qkyrIaYByQ9p
N7OobMaM/kYOUSB6K5uNnzjdFJbeFSY0gI51VpsEZ9MT4xmSIz6B4NngPLy8aEMa+TYmeApS5abC
4CO4AMKDv8vFzz9hPfUsmDNRPNwXD1LT9c2B8Z7folzXNiVIUwJXvKtP32YUUbqj+oJXcf9fO2Wx
E56anijShY1RZg8kc2qzh2LQ8vScaMvhgrsqGPIQHWuFglGJfSfdxMDyD+q8po/vEmRvWNLJirPY
psS++v7Dc5yOzf0auNSAAY1zQwPkCyjnU4fDUijxdEB10R7T6AL/vjW/VCyAu2tbCi/8qIWdtx94
dSC0UGyJJwKby6QlZSIsxRHBLRPnuait5RlW+6VZPTDfXuwsQWNLsnEmeqA2ygzp782EX/hLi/S1
Fwpi22nmcb8k43i1XQbbKWn4QpjXVWQUnJqT2ByjlIXhvyIB0hmntUG7oxellyCmZtasFkQbPc1G
44l+d9DI+axE6mHeCr9WThsOP3xGZczOtRS1UAbANX7lF5KF8eTi5z6rneHVKUsz4fCQzpUpZASk
/i8IjURLyiXLWFFY5Q3vjhwCgr72kxyGv9+sYH6BgL96Qi8ILACOXl3D+6O3k3UCBxzSydaF1pUj
8EoAvX2xxn7U+KNoscFLpU93xpbhVFXS061fjHhIywLw3tSsw13uACp85YvknGFqCFGF4q8Vfpy8
Iu87FYaY5fEYNy5NuEv/Wb5Fd3jThP4b/imFPwi0snix4nblak+Ma3Xp6AaWZa8HxWJsV1k2cL97
GPfd62vEThzm1DEJxEN60vmomRqVfbWcUuMmydT1msYx5TWeOCgW5UfJsKxzlbZFtUanGSMK1VoS
ahlKEt3HTXm+A4BhKLAGatNC7+TO67XKTee7BXzermjrwbZjcItHGCtayZSdCmLxyfIIai8ArvQY
J1lI8PD3SMmyttDd2O58BGyC9IZScrVJlhgqetT8BWrKPLTAuhpMlFr8FM2N+IlS9gixF6GBWpKi
NTDVtB7QRPUlnLUYQS0hIJc0boTfsNI6D+JlwL0ra5JJRPDqvzGd75BEy5rRg9pAq+skgyt/jc1a
RV8OMHe/H3lsQeTUsv5Tbu87ds+SHTULibI8K7ajRmPsepnmYPA0r5SD29sZlhrjn5XhkDtzoicT
zSB3J2OYD0ODo2Xe7nA0o3VJTIzNvbRZswmz24HJG1mATPpG1Sy7IhAquffO8OIe1vf5aA/qyRQE
tX6BD2BUSMrsN7nq4WHQSAW3Pk7oH6DXn3cyTsC6tFevmjqs707XMj+EmKbhq/jF9VUez36E+r5l
AY8j7zq4bPIWfRvOkbb2PST8Hq+zP5JIJwbcuxVtUfVxvIm45SvlzT/F+Q7E7a0OP/W3j1Tuoxup
lRirCSqncS2BPF9UmnPJ89eAUiYaH1e5XBBhzvd9/M8+ERQ0gzb9snh0x1z7fmm/a5l9WAJBmNoD
mQOH9fHa1LuPCLuXl5s3cEnmkwitman/qkyNbyLFo6K+HX+8zcmNXRYwpPKEKfpGcewp/iajCxYf
6ogz3pFyRJ1irsBz/9WSeyluxUppf8GpMYJpapAy+611F1VOUZGowGLN4AfbC+ViD1S/xmKKM8wW
F1FNv7W7CKhQUFBSluCSLLgads7OHr2UKlyZXBkLXzgnFIicU/ZnpL60WVxwFy9W7jo/T0JNUjvE
arf7Ju653P5Eg/N5A2+tM3d8L9vrr6nNvOd9zPkKgOa6R7yoTbIgN6Vo+2VJ2T5Eryg7Umcx/0ts
AEC6XpTGGGtc1du7i9nzkc6npWUSyuD7VEJHTL6O/y58WyASvgWZDUzbeIrPGZg6w4X16v6gyCHz
Pg784DCrWyOlk6Bzb0YIgexBJ8Q5KtFhcPLrQrGEIhyY4AGnGqErdLxKQVQ3uJyRMhxe4AqFV+gH
iD5mSCGIYrwMpF6wrviYdkPG/DZ4ea6HdAZdKj9bgHhSx3y5WKdeGpdYpiNFejaTzy+IYYrsultz
DmB+tBSUoC0XElclCb/6h7LjG7dFNJkuHB/q0yaB7xX60H3GCjvEpShYXtqaFWJfMLsB58ot2mSr
aLZwQEumjj4CZskN+IwSQ9N1PTWzQ4NYtNiJSp/6GfjIESwtBMmgfAoyrpIj2N/kfA3L6my9z1hu
zT+pPgD1n1sEU3m/BlxKWC1okiGyfMQQ53mHkUVKKpkQ+V/wu1JrnHXwILQToAiBs2ECrkU5vAX0
gmZwIpDwyaAOn/XcK//X2jbC3jOeE5vX0+v+TNQxFxrUgIrOpoOUBzcPDvrRbVcIvCKjLYw6ttQm
VqEG7mt2TtyNL685Wl3G4xApX+CBTjq/MWhfFjLKJHNRbpbuCjpmWRrTtk8RegpSe6+l9HXDS0Mh
bVyD4rBKN1VuJVgkU3eNwIyDShz9DtTGGqb6FzRIDPw3hivK+ORaH4rSbKZDWIkVQf6vB2UY5+kh
lQAv6g3EWLWP73tl1XA9el3c8j1Bc0hr2ZkODV2NEGQY/cj8ZSNSwbArEYvHxaDnToGICJyVXoYX
BynqKmBTISqVOHksfEajE2+DU1hHjFKToHLXwGjcrl2Cnmf1dVkG4pHrEP1BYplemDE577skVKqb
yHUVi/wGF18+8NCnOvA6gelDKvm8ERb6pXxA3IBgIxDfm/pV9a/z9GspqK6cX7H+RBZqCNpX6jtQ
5x+vraBw3rFNNdMnEC0MGa2QBFhDhTXbTzb88M/hrsHdO0ivhMX/sdY+3o7eRmHuZ5ZnZ6hvztNb
fZVSIjrAFCSD32iiH7/deyVVT0P7v2szpMmy96wDCXD+t046zrkZ0DhMExsmeMq11PsDRO8WY0Ox
7s7iIuAz2AujDm1STlpDSaB4h0rPidW9vLmXUrupO8PVrZKhK8n23S1DJsMKROG/LwoIPLTLsbkf
xg7XbbDVa50cwKVl1GGvdAj1e81BCGz4R+LmoTh2u2rPusfuhCLNQ9bjdR5hre1n4JBgGBo1GXvf
IwjAh1VOsDGB2arsoLhHICvnWiG/N5+A7xgpMP9HFLBOWVNRfXhCycvfR0uTO1xFzd86UNWXaDST
RMfo/d8YWQKJeFYzcTi3Ys4HTvm++mBQijT/Z6girWlM+4i85s2g3g3QacxpDxdDkYFIZrKShrXB
WaJhg0lJKbot6godsy7GnSAk+0sI8puNR6sW/bLcbu0GMYSlOo98Aarpd3qW7bUdhDhGxcCflS5/
r8tjgmdavvT8bLRSRYumtrwW91iAI0uyTDH9FVWMMxQJj8EoG3jMBMUhTWfW2Q7mbHy1yCoFVNcA
isbJXcGB5IZFc133YEMeKiNklH1x+5QWYaqxCabN3tvkyrVH6V7cGGmrXLMnt3tVxX41jcOHTwhB
gjbnvvu5Y8dNuYQ5q+hSUPYItR5bYgHlH2maWwGP6CWrc0xzyHsf+R81RuUZ0Sg/4UajPC8L92+E
zeSZVZjtEN3iD9ePxYMvhEf6Ie+RXdmaxLLPhH0Evy+SagUSr5i46JkVb2JrYPoTSzBcdwHSymiO
Lda7L2k0sqDZwJkLuOX7MWVgfl3mfs4HuOeEexIL48k0iEUM20Hl3dzH9ALzQqeIfFLRu//kC6XF
XXk3GkuUTHyhO5HMUQlvm5KFPsOKSOwkTv2gVTvkmbnAkTUF6gqbha54JQnQnD9PYc/2F40g0LSQ
QuRv3Z2uHppHR7g0C/2SaOhfM8fAnnZ38UW8sWmwctH9kvlgGwBY9Om/iiq/xxSLKCIe1j4BsXrM
HUCX70f/Lmnx2ZirWtRqD/xhPzGKhKC2NbhVaG3WlKhK1Ea407eXqoyytRpWnyc4OVsPd4dQpvIv
0Hjmy9JIacqjR/Sr554fDuhooaC5kgyyevwYG8LzDBCGoWUUtv3vsuB68KCA45hHi2/qPAjrL++9
yIESMnOdFrPF4Z3kpvPkAl80KZCbsKWhYTYvMlmH9x4N7nkMju2o94cMJBSsKWiqlkA2kuEOXK1M
veujOC0KsEvEkNS71s7VWyJnPXtZGiQfk7K5nNn2bWvvN//B72vbut1HuLI2Meog/AysZMxzj3ew
GotcYxJd8n7jQqPEY5WNeBj0+662S/rKNj/kwN0UdZH7m7PWeowif/0LP26fi48xt6U2n0UF8T/z
Rx21mMd5/otXHdY44B0kmeEyXgCsvjuqq5t76Bhbjd874qrhJ/Fy9eU8AfZRcgoYqWZTawhnPYR4
cFIPwKEL4CwaVWTqEZtxTxryBF+I6zPdlCIIbdXiZrihrsX6xKYdO810Y3Lu4vHd5Rm4LE27YRis
OT3T7c7leLoGLx0iNl7dtJWAcZLxzLsm+G1gUUV7dmMnCKNktVnDWdrhZWm72XuJK6WFfX6fNjlH
69Fs9Z1GM7KX8//ihV/TVtmUH5iyhwq8LHVVNHX1QtjdNYn3Z2WZO7bKaXsm/OKX0jv7NWAyagL4
ZInBYVC67qtBJ8na3x2qdNBmhL9Qkqnilm2/hSlAEo+tWZPXalpNpKdYRfdHUCxrTki7dY5r+Vwe
YnwFx3BN/QuL0BJ8VgDPnLN4ODh+J87XJJPrglJ+XEW6hhq+kRh5QohHJmRgd36VkUz1D5dWLtZk
JbjM6lKX8PoFgbpX4otYoV2i/thPN3NUiPrjr7CV2yg3DA0txpNPOqtJu08hCLyrL6ND9Q2HqPNp
GwGbCrWYkzJBXZ4yDsMPnvKS3gFCbg5Y5sT6XMrxLrZSFfpK1uDh2JV4fbr7nf2K1ZmxlvtdwDw2
zZLQ4q/mCKA3/KuIJ8ghuXRHLGC/QTPtYP27ZwEDffx0BoiASE2RR49at9eWTWXZE0+vspfE02+k
uE2KAmZUMgWD0yQTWHT5yPgb0A6LNCJ+UM0evcC83awlrXdS6XYJTNBrmhHYJAnaEPTwyssL139Y
IoB+Plxa/cq0CYrYc3AWo2yXMurZ44Cvd13nemln5d3ixwsfAcrtW+oGcGuEmFxOj/PkeHNfUgqA
ak3esL96uWRDYyr+WKjTwWEqx/5rDVPZEIO8Ajgb/ziUEAQEy9kMAfvHcBKbCYLtYFBkF2rsAQjv
2UcSdBM8sHymsOss4w7MK6+J0JpN95BJH1myRxfx0yxPA4MfzBOCSJkyGmBojU5QuJkXpOzpMa10
GUXmPg4rlS0+st9MBNSRlLliGlDnIEFTppB/gkEb2Aoc/qIZIQJGMHDNPxYAX7ZlM1nROpDgnH63
nTWnbQ+njSV+eeIIxuoGO4oKH00AoRTg4Ir3B8y40fZDbZfsM0L0RMhd2+5QsCo2MthmkN+f/21a
JvCdwU6iYe8YsW29hR4CaMDLJ5IrWQvSfxGkN7MWqiJAcHcTyeN0m5nSFCeaDZcGWhD/teNC23+F
999ninDjw+xmDKi9+GwLikzOAn5Qpm8ZRuIZcHwQvSjU4bk6FdBl+V0+r0JKVN/UQpYldgNPl+jn
CG6xJxn/pifvVErzFfOj1SMIsELNLLSijZYLPWGUPpO8kiq5uStiJq2T52oRFf76WzCGe51VZJWJ
hes9ElMVKpZ/frlv63Sht/mmOXUAyRRw53aUuZui1Mwnhk4YoF8Oe0XnowVb93UhR0Uylr1o8In/
ljXBaAi0tv1eeS9/q0PBOpattKfevlgO7EhtIzAFicviSMtSu9cumdHYiayeFhZI6AVtx9kD1PM1
Q9azV0w7M1y7jj0YNV89iQX9MKepT7QavH9pDOm8suogrLiOuj3UXRqn876a5zP4mJ7zE46FkPgK
st2RmsdIZkJMk/+Oy1m6HYTXuFpt2BrX9kzQdvbx9doqs36v6cyp9O4fnDMsH0sEZT+TYQDliOmX
16ZpPWopTTkbWT+XNusabVQjhrgiF3yJJpir3NLIu+Z37AGYsQPLDCddqQ+eXOwx2vAnCZ/mLLd5
AJ4cHiLzIE55+kcCfV1c/ETAkXVq06Xq+rA+KwQlaRlFkA4p0+u141fObT9kcPJ1UMvIeH1XP9w7
xXR0Z2aaJqphOmFCW0MRv2uB+TeiIjxtypaZ3eMAH6DE0nEkUcdJXP1uVh9p+bNwuw4axqnng7hy
HpMLt3J7S9Ug17fdq0nIs1y6GHcX1EFtr7srCPHnkMKVPWVpuVEFqr0yAi3ypwlSExJt+OWVF/av
PYzBYpPoZG5a/LqwQFu+5upUKDy09yQ/Jy99goyAUcYBe1y2HkPmm0LGWJPbgOdVDp7ZmSgwvqjv
rS4KKhmN+ErT0eykxEaXH9bpWUm8eZ3XL1fW7E8OMsNNZLaK6TYo8nZp+/ByeJv4+TDL2pwGdGet
xDV0nPIQphnuw0AuIOzbys5ytth3hSfr0mVQRcBvz+0FbBthcDbOoodV8Ku0XAcdImdJ5bqCVefm
0iUVD4hJ6pGYriIjXSAdNziTUrKxhmb7lBZQQwcYXHW6vpQfRSMjH7vOQXP8VqcIRn2KVoGmhkvS
ODG9rPj8Ts/BguQuYC1+IkRBZjVwvDxY9Ga3qnLDS2xDWl8sioDuYKLkj9YIBWQ3T7jApN4JSyJ/
QAcyD5mn77JMwbmUu7guTrYQVfDX4/xuehsjiTbCKEmbRushkSOAIecKc0NpWKMk0dlpjok4ech6
lakliFAB+p35vYkL6XcNHAH+C3vmMbvy0C+zfKvOzEngPRiC4pU/mbkNcJYkSYh2nDzxBKJ41gmu
jj89+orrYvNjQ+glQY6XeqfF3bSA3B7QA3EVT//HvGYSAdN9J3Uk7Afmr7Eb4Krrk2afz2ezu9Iz
7O7SrDxan81P7zUWAeSjyDF4fwc/Kwu39qIcEDqcsSCA1fOLQDmUwSQ3y2NyQdYWriNh8FuxEQvG
HinoiDg3j94Xilt0Jb6sWe5QOILym9wvbXwhdVWtXjspA+0S5YVJuWzSWJZWwVgHo/LKa29HdoXQ
lM46pq8SQOsZyBFQwKR1qQIiz+0yg+mvwpfsiE/wUn7GlkhNI0FBnL2iAnPpf4Z9eiqoDY3YmRs+
/JKMtVZ1tMpfGIkGOhmEf7FCVps3IICts6Z1WAvgWS6tj990rCeUqlAPTKFC+AiAqf8jM0YDZUsh
5rrKdjbkgClg2Zk0QBBMc8/2zBwqoLLPQ1YAqg+uYjHytoIl+0zfvUbFHrNPxEuv2zF+AATof0I/
mHNiG9Mj/WX1TPFtuw4EbEpCfZXUXfEMXuBfAP9svFzcZVxtQzURLSrfaDM77KVzdUk3u+0vXC1S
LkMKIasy3QUTdauzdEpC73RcvsFFDwgvOaLCJdJIHFpeMpqhFwUA13/EKQa9fkXXHQSgd64JSG3k
SIdj2pO5zm/tJL65RA6mUsOOBd19SF58wNw3k3Z6HVzYcMuxLK/XqMHI/2KKMHxvRkrsb0DfR86m
UurLdeDs62vt1/o+k9Bb0zOABABAYO+Ez/QSYlboSJ7E87++ho0j5jN1c0FFWQ7s80hJMDlOLnK1
OkG0TXsAneLPX7R2/7Z2LEX1jgVMV90Jfbt+PWsjTs3srE4AuxJWurl1yVNQthcLEM9uzMleacTv
xjmKa3u+Q1pESZb9c9oWZNeth7RVm2qxNYgVfAXRZRaE5A9XkV9suaYWQrIZMBcbSe0P/gmodkHW
y+fMJpv7xKB3kBhUZlJdCig15ZnaNcRiGcD4mmKmpkAPu2X+ZyH+EM0HWQUcEVDqDO4cEDx08/nF
DCAfbQ7EmLb7czcBaE9ElAAT/8O18v4JhlIPRLnAWGdEs45wwAgV9PrReIMIQYCSwcDBcv5gm8iO
0oTO0TuPf0O5pN/kTErbVsOM6bohGMJzjTqvsKxCty9JDN7zgqs+fGlwA9fr/7k8iSZsSZPsC9KW
lC7cq+S9lcydDgNsX88wgPUQAhqNah6frV89boI4niF4dpiao0Zxll86aTaxvcrFTOu5BAmCUpGl
vyf5HbtNqDZo5kYvRPxanGUKqQ0LwBf3Pz10x82YrGupz+2FycvN+4c0FZIjff0xK7XF5cZxgrpp
25UeaA3m52mEmMaQV6TqZAGcVgOx4KsrgaN3pe4YXSWZdU5jut+Nj3etSbfg9QxjYBLFW/K5Xt1Y
mPfDIo8XsvsMDGtP3dVJYLK6raLGCWcaeFfshKlp/t33QkuZ4dKucxxBgxeLM+TE1m0GZj/aJ8xy
k4rnTvenBSLIgWXq1GKLAwZDlkAaRrxbGwBwU+ZSiiNfJwk0Yr7btjvi9m/s6kBZesKWTgeYB3fF
niqQFvOaFiPkuYy8C9HgeFRpHQUSGur6TWUM1WntDiw93yLyJybOSp63GuRw+FBROMRJIqPNP60K
9zAOQELmnJVNa6sPRJjyb95MWBl0QO/YNHKX/wyZuyd3iNhhS6iIGmWR3j98pb/4mAoq6V9LfyBb
br91oq5GLaMBWzrhLeLmXinwEJ0DB3Oms2ENde3SQUbvjufvFnwoIShWqVuvL+Dqw20Aai1b6OSw
uqYNcF7W8nm5z/jJhT+jggNgP/5c0heFioiu9aIOATqO0v/AlTYUyvJoKS6d169BeRo+uGi+g5fp
E7sUjmX0j7dTO/9gRsUyImEVnGgbdusiq2mGjIygN3N+plsz/EHHiTayYk3RU74Lda7Ar3LNxnZg
Syi0JMyHFF+p8B5+qNNX679KnFDKI9ZdIlzsKXAqkb0/DWNp8wM044LjoMGamxI01VS7VJTnwgq4
Zdlm2N0qQQlPLPQ9kuJ9aJmf4+MOpg9X81EqDOoVwR1t+vcC4ET14iilz6hWJkNVktIxCfdhpN00
bzsnZJEEkOgMYzhhMPnrpt6ArES2t5D4ignr/yfib4KhOdEflZIidT3nRhaYgZ08wG1llNmXwobI
bLTPwzS7kWJ7tBB9CXuuhMJkfwoZr0oKoVHHeEXVWw7q/t8q3vyX4BFB3Zws8Q985pQmW/EuG5eZ
ygZSeM5ItpMg8BKuLjIYuGh55z6DkUrnNWjBFEP0iSbEcT7tFz/m7dQmvzSWMov2a2fMDQijbrn4
8skqM1eHhzJobQAV+I2BPM4cCM70/Qi19ahVXb0lofhBqRUKi/Khnv5JINXYJ7gBkhzGjY6M8VwK
x0iiqQBMgp95xkhN6DDHu2LSPIqrFoqxGQqsrYRXqMDzCwl2vyQox8VqBitbHvAY9Wf9Ck2ioTZq
DpCaKh5C61sPVToOorfJ141KVo8mYayNdIgjAos40zmwg40hhOBl+j8Rz6bngVIgoU0WcWcHCRip
2z9Sb0eVDlavPZCy5pZspGZ5FXKdOBqHsxXPX/mrqJ4ApE/SKYNSPUJVlST9ZFvQiIkwQmVMSLgd
G627TLtPBUotR2Cd2gPfp2TVmB8xBynKQc08TpqsGmoh7RP0JkHfGhgW3LI21VvMaCBXuOUIGPB3
znZPylNrWrzaRTMKH0eumCnZgwS0VXqIiMjp43+OolnEMAu5QRSEe4kJvMucTBw23sI3X/EkhW1Q
21iSA2SYSMhy4udhCKZwvU1bmN+5P9n8oN7FnaK+ZBHaCCJ5Sz664Lt93UHplSKphPAmNEGxI6Fv
VZtLVlE3URJfwgNEuCW5XPlYnAeQXz8L1Itmx5CJw1ynPl8QAyNw71di6kT6UiPwtHr+iQl6nb7X
U4vcj+JC0n6w7WvkrN1q6y5bN9DJCUMvBPZcLJpYjFIL8haY3OZ4tdEnEejCe1SJ3nCNXy1x8sQs
ISQFF73H6DXNGw5HqV/XIjIDmoxxwh0z0gqsXQnOsiWLaXewoA5meksvPPM9M+RSYo6JOe22cCng
CLAIvMZ4a5fPniYUXfXdRE+Oqg9lGMlAzAE8xx9LcYRprh1k8D+oobsP+k+ag9CWERfhgapPziYb
OXwCQXyKc8scI8QQzPN9bi1jWerLFXf9pCeHF/4BnNTcfsj6nFfgodkjfs777tUUo6DriZgiYa4m
Yj/2rjACWNaXJSL6GqC8r2Op1/wEA1ZWbsP313tCbiaohw36t3wlNWnmWmbtBZtQITy7PQEtsek5
QBkONwhxDG6hdvoei5kaq/FwiN1hWKmE583GSt/kIU3i6Puu3lAybdd9cwMX7qt+ws282m6GiaMs
QNLJsr0EhwDvhIaABw8reBp8bXrmIen2RmGRhUZbCQNmd35ZSxAQ6UHRvw/U8zx9hEpvv+jAstMy
NW8UJj8ykKn449BHIi+Wvn842Ypld08ljm40h8gXyTlr7L7AUc8o7A1g7UP54m+21wPElm7RYpDT
1miO+Hnfccg7zk2LPfndPqIFEUX684MEDBw4sj7PxALulkUtTo4Y3UZwZSR55AxHnHuAFBObx12V
TnOyG7RGYxJc7Lm1YkI3uMok9PBKFQwQTVzqXc+k20cuMP626bK1e2NGUwOjq6SAqbisdh1i9UdB
wvCiVlsgqPiJZ5PRUqVqgOqTNxheNU9SM2ieWHVAuv0ZF/ISaJZwrE4X4Yc+wrTPk+19KpdI5Zry
06B4pMAnjpzfNv85JmL477f/MN8JCXV5dVI1LwqR4nZwRQhe+ny7UnsTITLrsl0yzaLejK2Ame3E
wqXQpNQHENrfEj1PACGUGW0rUOUp3SCBmfqDe1zdhFDztcXUHcjyFTS/UYtPzt4KGiInS5++akoE
eIEWxhMaPVeZmt7m8yuPe1gt2uZwhwta9yKVf8mpiwgyZ8AnFZ6KA6Cyy1k9aUQfkJvviNT9Ek2N
w+fwW3d5ppV0Yw/06vsRruamtNU0GSUlRdtRwOyYL9GhGSYRDElfswYiNirZNuJ5SdlIRMK/F5T8
bj4LBu//TY/0r5hHq/1fK+FK/hvOC730YIsOjOr0z7gULGVcx5tSd/Aacy5DnkF8mJNiS+qAgB8x
7p600ebGh1N6Zx/PF0aIw4f1N6eW05WnxGskNPuGCR5CyyEH/bD+XXDC9Ih3uAm5WYzP7wkkM06D
gB+1S0CE7uRLkHIPFJ02MPXcnR0x5f9NqMq+oRvzhQGG1P9eBGGK0OegXG1+43YfnEBC+MYy9uHx
7QuqlY1ffmGpLNaxo5+WMB9CdWoOV/9QhKZDqlYNuecKMqPvw3iRKhtOnZ2Zi7iHhe6r+SEZ7m3I
TBlebW1amFrcONg3fSiwEtRGLGo8NgjlwqPwhpNYTyyiKA8sg0KvdSDydBh1lriMSoEEao0G1C6z
eBxjtSHcrPl3CNPeP8IGkh6lQB4w8QiJE0av6eRpGtUPEAz8zVZA+x+yyVo6Q7nrVqnQ1wekot4D
XiMB41L5aub/cGgWyvWWv/p6G+npd7I22k2I89Iv+fD9MzEv2ILKpMrBS6JmQ76ySGMI7eqUz9K2
bHakq0J35Ocbz63tBMA7b0ry5GnG+A9xyVam6wQwCIylssjJklfeF0AWckU7bX8AMNUltOzbem8Z
CBz6PQT1BiaYRy8jQowj3ThX5YBt0nTY7F/UvOeQSbMvFG0mUoNhF64uzRwbQIDIVZ4FV5/g7qKi
WJSDZfmBn6NORB7pk+ZcRjrxA6LBlvhCqYc6wgvN9PqDTR074BwWjEBhY8QkT3DjXvRJf1Hpx/8U
EEDg9eZ4ncj/SNfShQ/VUUsgtVZ+YGN5DFoUqZ/ga+tx435z+tLSONhEBNVoE5L5xO/VyGBbzdxo
9mwHZKp3qsNmpUmMXNP7L7nBDZxFvLFQF6EcLxVLROOTV7LdkcZ7Qdz+L5gjB6CTYqn/8V3eF7db
scXF5/SUl3Q3aNPAzIRcYO59xVhTJYW8BEDILViTzrOkPue0fz8ctLkelsafTNcEEkH+77LOd4MN
njdPhYD/tLhUvv9cN3TLlj4w6l8VNcxeCIdNGWfsZIyit0YRYSQZ3+a0bLq3HIYRL/VPdARIKOTW
duuFzqc/EalVjDZy91nQ89uxVAe5APLDjkOAYnqx2jg2S/vdndj3b5LsFCmCtzIY8rRKfW5F3N3j
KuKrkkGnBWzVygJETsnDjteTMOjc6TRV+sON5iGx72BXi7v5nb0tcOdmi/7/cDALzqZvlbvAImyC
BZlTpk74UdOL808hf2ELZzHLJaQohrF5QWw9enLJSN1Fl4/WWY0yZKAQ2VZxyfL06kNCu6BnvsSX
Znzla5LSWBH2GTSwQTwSMtdj13wO/8ylFFOypWpme+n74HH7SNEA376e2p99ND4a/de1pCOHa4PW
IOB5zP2WDY9Xobqyqs9ICCXQvPjaB+vyNdAOcd6bcQnq4H09w9O9+YdN/eK0ttTxTbPsr2gBEsI4
oJbEUyPOUs+MZ/iqLtb4k7E8T9VDpQPNgy7jNkWQfylo8lOBxtPgrbbIJVVIkQawg2mHsF7tWm1W
uBPsB9I335tppjngP4SInlv35UKhNJoB8/mIoGIjQa8qcl7rC6CoaN5d064M9M7wqxaEH9xpbMIp
1o5hDtzyiidvrbRCtrVXrdtRjv6/5Fc5ONLgLr88bsnWDLg2lVLBMjwLLVFrKZ0CGALg9DDrOb9x
ADFehf4XPFFkTPcrVr6hxTFgj6Xxt96QOjriCTY8S3H3hu33/lBn6YlU/HXWJCQ8Rn7Ds2EG5RIq
SCo86DVpFHKJwOSNOL5I0COzLNaaXbg4UuRMveICUEPeVZSR2+FIvA2XoFT66K+vGFjffy0Od2JW
4Qf5TqDekHrzItIlUtr0Xr5Qdmnk6okMh2sCH2HbcPb1IuObMYX7KD+AD7HwCue8xorfVPiwjF2i
2Wj80uk/auRkNosbEE52gnaH9d1j4VwHKFekV8zYuRoWe7gEY28nS9IZhmy/uhwo9gSFqcYiBk4V
78V/hmz4ZaPheFEqyX7pxN6oCJHAXDPo59XfQEvlcBZajJvFcHalyJggvcrfQJDPJOHh7AKot+BI
x7Rz59wm3Tn/4ZyhuUJRl0imC8XWj7/bj0Q0EOSv7TIy8cjlrtlckHP0c7q1SZhVs+xO8qRN9BRW
dZkztZCni1wvqNLLz7/Ertq/ASjsGvxOdpTmYO+zDZffqwO/atVZZjFm6qmKD93b/KPMThShpy8d
K0R70UfYQKw8wHqJ8Afiz/OlgxUrBWmzYm90kfwYmPecJg2jhSUFaOX6hw1aOzd/mzpsNWTMQslr
YRX7zwq/K98Dlkr7/qFIugz/hkY1By8MkzAqrsZYfTrJXYqdeMLHFVX+LecNQBe2HjuCmX1iCIxn
A95THBvhiuTlGGtNFPjZcSSTUWT190/jCOz19gYBkmsS+oMWBA3UV2mrAshQk4RCyKX2cXB8hRUS
/+M3tgPK7xjndBvAO3BSNbzjx8Zlm7i9UgVvyjeDQt4bBEdbYBm2CoxifF/TYH0lXvDsMyaqhp7X
/sKbO9eQj2GHseJdNkMpSzadYjSiMM0ataBP73IQiazE7dVrJG1dT3XyPdyOtXQ9TNIbLsw/lh03
14gTxWUPcFQjHRXJMkgQm7cEzL8BCpuoGGys5F1A8/4vocELefmAVP2tCPwQSlOX0+2H6ufHpGKD
YR5ywiah77mgM/YN9WpUKAADh5JoEqTcdFVdcvm7sg0gxMsnj9MKoqcLk0WeJbhbA4CT4fw75ikD
9G6Y1k+rck8VIUaJpyYkSln1OLG7xxDzy0JOb+jC2GRNcNBJB1behonhoXE8Cra+sQ4w1FXjsmH8
fXue4+3YTGGUO5ohb8LloR8c6cNhw4KrZSvkPShiQNYuR0/DlACOBqkQfCinxhkMbF8M7SkUWgVm
3q4Kqm1OgekRgEpwAPhuHEMcmBPHaZej0ciepjLHmT84F2s34+Od6YBqjMRJhqy9F3u8sN+cY8sN
gDSiE4/z3lOZdlCMSlwkArSdAqsxHje74ZWbendTudwWmLw0pv7n2BIqpbOsVOliut3xAeXebcn2
3zIFx2vn7IYQdGk30nlb9E1Dy/7flICNFvOjiEFTUuiuYu2gZDYqwBQdw6KFvJ4ru6KoBIpHOIG7
XaY2AjQSNCFgahvvSxJGgPhocoOYMTxsermpgNyZABqiYjQuOfENsHmDpSoLA6KOoGbrVekH426l
K6UlGttpbIk2SGLqb5UCSjxRi1E6G3lFBTWAKiUI53Q327Sb5hGTNINix0yqvTkEpEhp/US2s68a
hkAlrLJRmwkaffV+NFJ/pj+PvxGkJ9jIZe+0b3gSyK1KDWge8r8J0oKAa0UVEs1y8VYbJST0LMhi
+Pp3OD/IXy/pxXUk0cedjS9lR/SiCp4SnyDImlqE64A/rXs+UEZ5hzIyRn9LfuYLbr5XE3dMBC6J
u7jvb1m3ZNrVw7UMsscy9SdnrbbUbJwIuf29nSvMtpCv7UCrRred4d65HNMjXpRwWA+3bhVqPEa+
l0otomN7wTd15Eronq/dt+XvMbqrnGw2DdbuIf06YcMaI8J0geLNT/xb1dYC8Pme/VXJ9obv8MHd
oFQy2t2UUj3V4b5zOs8eqk9Qa5IAh5OwL4wxx5uJwWLcfxAtZM60Acgj4i3myOdbgRxWH6I3oVn5
DyAQmmeAzBDK7qqKCjDqI+ET9B8aBJowtfnDiSonn65e+b1QLmnj4c8XxA2OT02jxsljXaODkQCV
0ERfs/wqnq49zVqeB52EQMsJSRUl13GeJA4J/vmJ6HFui7tuLIPV1ZjBJTMaK10F1UmhlmxxsKVv
22Emmp8NjOumbfh7U92jlCV9bjqvuEgeFf7lHMTMOzB05fwNoLqA6RV9z9aRcckgfx1+6X0056zy
8AHcN4CwuJNzssf8zEt9E+JFoxvmiSa2LRm6osRz+93fIuycLYfKIcD3hdWvR4UtNkK96z2ynSCr
WcDtkl/q5BzdUs4zPgOH3rpoU+pAtIipoXzJgGXjK4a9pOqQ/f5VB7HWXZ+1LKGtlgCN/h/hNT2X
18YT8H6Iwd4gkhpRfmLcADnV9ss4TZPm/S0IyCiov8hVRYPhOpOr/V9h2yBcOHLwKD7x0g8XCmb6
RxYL0Gk83rFSnBjobKIGb9mgWKGAl6HDX3blZ/zGxA/RhuqQn7hS3skfxn7nsKXQEfb6FgmGpqDo
7EtPioHcaxx+JZGQy63U2xRroJ84Y8LCF1VV9o/NGMQgmOvKyalIDXKXzAWFKS6ZGbl3Lo7f5Ce9
cMCsJg0yVp51qzcCNY2SENmbZM+u5T+ASl87xI6gFQxOdo/+i9duI6m3egu9wO0uGL9fKhuVdT8M
0Fx2YStn2xHwhcWJUNNeaXFkMUG92rVvneKCOEqIMstAWDXIDEU34QOEPtOM7yxSuUh9g8/76e7h
/o23eBOM7kxFEaf2nGoHtrt9+93SAnRtIL9uuct337YyVqvyaThnAH4byosR+j/eIrljukwcfn5x
iyoIMqmQOPD2TpsdIcVwJKpJRSteeCTibmDJQ6k8NrhXwLq2jsz8IpL79aNoYhiZNurb7sch+RB3
sNlOvJvk9uAj9T8zJE/dpwfkvAPgmZPmXli9mbSmCh/2Ch1IHwkcDaMtP08mDlBQfkFrIZeZ0PiQ
3vgd761xozuEWue/FMspn0W216p25sxJS7jeBPqzqaB9ayYo2LFId8bdQyrGxZsoxIdmGG0vjUen
cTtPyw6xaTyPRmC5bWwBgbYLQtUSUxplRuTt37OmwXVC0jSQP63i0P4NKexcF3HvKgy1gwPFVp2n
SinML3nd0gMWiYNM6rpuKxvgciR6J9l7hwOUiMzRZht9R9wHSd+x1CIdbgpwlT5+5ZKEEdhrcJKF
VP/dj6GUARtMBFvJ8sC9bZOVgUYfgQbWhbNhdvcScZi9tcUOxB0mxVSlZ+2a5fAfhKNdwFPdwATo
B4qGJYjz8gqgoJPQpsIjV6PqJI9FAZyzJmGRgVrrWEfRwd6YhLTZ/Wj1viaakZo3qEzPpNpncJxT
xCQh2ZlB+2FMqmIA3fNiiwzkoLIuM9C9xAc9OKurFSXjevd739gZEdydFhdgOYKYl8D0YKM5Jjqb
hyVuRiPO5YbNDXsoF/r3A6XsF0UUHcbSronRHXnc7ttEJchvDm5hudQtGnXc1CEnlXtrsAD6L/xg
hJbv1VykZVGwEF9ttw1zZ5ffVxICQJcteb7IcaGI7rqSTdLAYvqsSI6a4/Xfq105+fIyvzpIeb1A
eIAoCJ5Fr8h+69UD94Z7yCiXWShhq9MquVB2OyeCErIrYamN7zDwZZAvAdr/LlQ/vaWY+n7p25Nu
WfxIst0JYFtrgkLg4FN32cthTAyNrdswecpRre370/F5qd3bnv6QGNc+KOkUVjiunQ74n5q+YWt/
dX8DM2R9Wfg2LkbF/VhHzx76N2S+4OJ/QiQiUN6tSWIXWcbCzlxCF50dtwnk39R0fByAta4CvmpD
CAwExPDUAu9xVTvR6aUEvIVKcyqbyNVvsR8WXbrjYZ9OEROWdJ0Bvup8r18IbLY8uuaBFXSSeXk8
/Z9T7xE3JsKU5s7hMl7bZc4LCYctnPW/9i7G/gr99tBQuYAbJGqPhuouwnzbT0AXXAMi8KisJsbO
cLTwzOSEQ5wdG24K0DmQGYKdO64gsL7YMvvIUUQaotPiKRGgeohrXvjVnj0OhEI13gJeZflX1KmC
G2o6FX+BLQFpoUVcDzEg0jjiUf6Pg/EwQZ5pTBizWqmxD8UehKPL55jiT9QTvkFDoRutmVf2Z078
haTq8Di3BzmXhFwvhj8zdEKcCy6i1zpxnNdyHpZB8NzX8ymNWRen6g96sXJuTqdVP7pgdj/xtOxc
lJvGmCZ2YaUYQIqGavH1tkICZaCsR912QTPDrFWUjLdrqL1JUIle5JiFfWUi4GKB5A1swcbOgFwy
yefUgNv6Rnq2F6mXI/zQS572xcqQd5ST3aor1PEifWPa14yVpjvomSMdE6bPkSB4qaHW9ViAuvpX
Fp/cAm3KntjdD2MchFpiUGvn+T8FIVT6TA9LA/B3tR1X9g5EVlRWhTydBHT/ccdMgDRGuQ1MzdlK
o3PLLQVR5Okp33VurlRmaL2VubcpJ8/svpHTnVPu7qF2NM4n5jp4NqzQTF/sBag/6OXR4pKzzRsh
SyYJCOwjiO/vw4kLiKgXv1w8uqfBWhOMh7yGzvGuCqrVnh5NzyZCvKpQiNWu7NSdEFPqXjqA7EPk
3Xq+D/N2rjLOCqCl3cfUyicVArYqeZWmJJxtZyHrUBTKauxOllHK+mLb3kGGf6uiV4CWCcD6r6sz
nWsdfAXhZa0+eAwHx7QutXR1zOrrPz/bXWhFTjSWI7FJWgnRC9Qn5YG4mWhT4Ah0NuqSvy7TJWjr
Kir1RgNMcMhY02KtUiozw9j39EcwpY6efebKy2rTR3kk3xWicISwHfdO/AtOJK5rqOQzVul9jxwd
dGJYABP3ydR4NZC6IUell/SmZI4CvzNiZxPTTJ5/5O61nzuB8zfckT3ClUiuxKjpej6eJrG5gxi9
ekMZXuBro1Yu5mwgKBBgS5kjApbeRDavWeRbVABQ/3343kGuSzvu0Bugvw8Xx10ZCdc7Qr4s9UdO
/3VOMP7D3cnjNVtQAKWsOhI6w3qmBLUr/xJPN52WNhVejS2u3bVyZjx+7juxG5d/L6VqGb0VFsHy
Pw6Muw26pwrJjhMYUyFucms6yvc6lSLKNKph8cH8nUY94iKoJkL/1wgp9ItVSLTy+XYdT2+lT4VI
cqUg/SkbJ3gkQmso1NP8ASXGNooboLejkKxHvIQ08odR9lRansRcQzImHQ3abqDH+fnV1rLNhXi0
k1F65vaGACcrem2suYY8NamD9MaQLcPj21CGVkZvm5UVmqwufjq1EJEQNt8DX+dxSu4mQ6S7N+zM
clM0o9NOIjwBbtrrIdaxTVqnJ6t+rXwhfMc2KylmzTMACc91e5lSXzxwYrrhO41e2DxU/9iE5Oa8
b/aCrySBvwBPQF9hEVAFAhjBLQYCBlLkUtQdBzrJvwf4eTNb4nDp1SB0BRHYjTIMX7HYvJt4G7sb
bn0iuWz4fhleWjkva4eQOW/mm3UoHKaLDUaOTG2Vjlx9Z6kUW5JybUfy5sJbMtcrHQsqoFFPyV9e
IaKKRnCG+/4sjaokjRMaW5bTwtHCFt2UvX3MuR395NmPryN+y66s4AzRX/pwYVt1Z8qEsU5/loZF
OPklp9TtuQtOXScoKeL+278rYOIHj/2cXfjjbxWRu47a1rJYdt5AGA1XSUX7472gX3dc7sTnl3Ac
1CVfLJJJRoHIoB/dt4cT7CuL1Mc21BgNIBcBLivLDeGfXBOXE+uhA9+gesZWXsNFsrbGfAbvwWDB
TWlstwc02FmECTFeI8t82a1WGnL5V8hN/j4a4RC7RGnDAwid++lnCYh6A12OhRS1b2aviO6/70if
8UHoZp3AmT0lDfvWQ3Tzr8TYXCONabogtlwP279hzISfCBQV34j2f5ZtgOWKAuR8Lth1mW9oMyVg
Bxm7DDUT8duILMOgC4zGFC3143YhBR23TcMp+SvZmH6WXnGBoUWAh+2h+1CJJ2ikgOBPMHToB6GD
ICvtrfk/HU18weW9RrGCfJSBj14GkhAJnKIw4HTuvriBsmYj4F2bQCdaNPNru+NOnnHrt7VdWV7K
lfYUVCK8udQC8zFCbKVgb7838HCaAlIOYQuCi1u7pCUDaUWxTHvipOd76VBQtWlw1IoWvX6LFtxq
rC02f4UJ4+kMSymvFSsAOX5cnSIPeap1IH1nxvxO89oVhVynHJc4AUblxMBR0zbxslZXhV32a4rK
IqkzR53rOi9/lczu+nDxPnSHrBPmVInCTjKxdlENwjfpDYuTFWmmUpUqlM6U3wZE9dlVHuGDAgiX
pzhOf48Nem05Zztr7A3wVZpZ9vgkLx4yLltZWomVt/4bYPRM/NvBS9SAvjYZ8mT0UCDSTXJ5RXza
w8ep7HZsNTCEtPYfjnId4Kak1u/pHpRMqHk1LYyLSa1r86mc+HSZKI51VZY52si7VRq9Ggn/7ILC
GBaUJVGNHbEP7eaeRWS2foMjQIldPfqZz7IKnJyMSeZ14qbjnnEa5e8aHTbZ7VpCRBzENzWV1vpg
U9VvryRv4Yv4Jr8Z3jvgYpakCD1XwOY5axetbTLfj1c0OMaSRuwCwSqfZvKei+cmwle8SArjgxtH
NFl7xeELoAuJ5IELnxkRAsJnYdkAWgROxYcGoKUpkaet+JG7n6d0fxwNDJjhucoNP4+MOtVdTPH1
wdjg8ebTahFepjlIYSk9OTQzLIsGEtxuYmM4zRFWX0We8HX/5ectziNZIYwaTHL8SkDZzWlu76cU
kkNPzrbT3NwhnPZLOJM8CSwafKXpY1WvyABJ3GvzE9mFNNDLyopS2+a5esdeA/uMcIDwYtuzAp1K
oL/o2UsTwTxGXrSlKAD4E7kmC7PGrswADXnby5seqniCNVKAIOQ9PDjaGpkMaLRJmd4L+KQJCPZF
Fmg2nxoleySreR6gOtf7IY2959z3EWapKUp1j4pCWACmlgb228BNpK+QLh80NRbP61NJbKcRl/ij
qcEd6cSmm7Gu7aprgGA8a1mf6K+qrOYJnjHCQ2H5aZJC7p3yMUPXpfFXcstr1igfuOgyiviE6qtE
sdwF0U1VQFZjoxirMEIGRr9harlUX0m2VP7tils4apfpmUwfdpSkrd//lwOLLP2MNKPx2vASrSpr
DR50won4pUAiwfbSc7nxzRJMIouoPQO9BuVMabDWegOIGNy1CcCcie2xIBdK/aST/gDyheIsFDG9
/gifUByK6NlgAeYVBgZrMHP8VI9tytMLdkxiD9EDMf3Lc3tb3koo58Tj6VisdnhUM9WPz5VRQnFK
SzlSsV6PWJ3JA276DlXzZoukWh8752Ab5NUct5LmZeZuYnCPkO8GrnPcXMxFNF2qjdDhEfyuR726
n1A3ndGEd+ArjJClm5fbw1ILCW+73Rl/+qK0Tgf5Fa+ZGf1HZWQH4tonX4o6n3bEslD7UacSOwvq
45g5oCWTrvje3LyXQVoyHZekidGVrx05P9V3PhBmEMsjy6UZAnd4xn6NiQU/MigYzI38f+w1Ba/Y
LVEh920r9Vgl/39mwKo/mK0r5ISXH90h3pAecK3tMFo+X2Ngezo7a3XnN6NRMtAhkzS7Mb/V9yXS
gkdpeHHF96T/lwDcmL6tVdYmvR/6LOnL3XYVHxOKjeCAyFm0t/hBRGjQ9VTeU4Dy0j+1wmbXBORO
NVuPnZuDWn2bHkmsB6Wt6oGlfaNGzPoSsgxKVmzHRaKdpG0CVPsVaTkyOMoe6xgGyNSdzrRvjAfv
kccGf6rQNPKHzg6uyN/97LFmoh18VWyr8pAFO6GCiGxELp5lBbaIDQJypxSfBictcO9SkuCskYiR
xoDR3zpyoTUEN4nYpWzPtZ52bq1mXGYAYybKFMLm1rkIMg1IyD06Z0U+aRgaGejPzToWHxYCwydI
QbD/L714am0D+AEbYjY8/xwMbfLH6rE1BQDNBxqpXQ6U9UhwVevU3nGniAtJf0GUCOmc4Qf6pvLR
LohGeDGB6WtqsOFBA8vLGgC+2luh93cr8ANvLOhfGR1rPgjrM6+1bAq3/dLecHA1BjWTMH5qqeTK
HHoA9hG4cbeHqQ3eAlwIFKGZiT/d1GYPisu4KrpZJOZRo/RQ3sae456Xpb4ZAXzhkGA1vm/mWiGu
3hdykm4j9ZHppNsQSr2hzO8+YbbDNpKNCr3KSxk0GZXk7ogzco7f8u/sehZcxvA5aPIFC5SMhBZM
kmibmAQw6aFpYtgPSK1/eHCsUJNIP7WuiKHsTYR0Kcl4qjDq5kIgz8Ps7d4s/TySlymXST+fykyZ
xdvQXMAUQB5idAKty1P7iWAsACSv6YUeXKCRQcf6px23UXZWaW//65W3jLnIEVKpzbfqBUA7hjrm
SWmK0UnhcAvCVuN25KHs4SQiO7TlZ9npLo+QAtuog+6vVYjkBgYeQCe9rGja2xtEiXWPpA6eWklv
2nshHVvoHDiyM/J2I0CB1chP6A0kbhm/rROmM8zef2bi+XsfpRCcDSGqprBj31nhFcGkDa0J6522
CNgaWfQn26stTKhnCM1ob2FYTlRKKiTYoOGVsHC01uvjokstTqE2b/lApjHBdvxfUiGdaOS2ZGAl
VPZaY5nFAwJt6T/VJYZa3QRfEISLnaRD83RFvz3MYSjK9AXFkgmp+s16JppGL7MFGeYFXqMlXQQS
LJovgGzmd1QLAVU5/+kQMGY/6wpY5AAoMxWe37lK7VAl6+N3rqtldNwQxdpU/iFsC9ZnC16iQiQC
/A5ToEGYUlHQ9emkIbj/RIkLIVsrhcBlIC+wRp7pFwh3376qCcPJ14MnqxaaWjXrskXLIe4ZZmL0
ik028Mjz/5/f0R2O1P6zyzsahSz0TmdEmWl2wAaM7rGaFKiFuY6zfgvjkNNYolPtQie9D3LDfwP6
n9LG6kvC921qN00UTVu800DhVUZUpnDKcSqtGuuFU+db1d4dqhWn/+476byZBDtIdfnPkKK04E1+
+3qrg27Xy1dQReKaGC6wbYsAHNo8Dk9imm5HDjmd2OqOogTEv2i5pb/AXrWsSjX9svuAD/uDSu0G
l9WcLKq8k+nSxghvbq6pNdEkf3OEFfD7d1qDeqKH/EChkIVqk3qvoR0lnqC3dm38zO2GRmaSB1DW
LE+Nv1lck9A4JngeFv7tkFmJvuRQBE6iQ4Gx6euSTCfSYWuQ6Uf2T3YeeEqQDvL1quaErnE+xutN
WIJWtRLHk4QR9N68ne8wJbEQdch63ytHIWOwsPIrXzttOx51Fx5F8khOKuaYT9TEyFgsC21PqDQK
Kn9oCEozc/x+rj3LQy7JmYUPpUFsslD2nQyvmHL0MUQtqKlED4ta46t1eCKnm+4Eo4Rpgp2csQ+p
c/HitkkCJ1TDJo6vrhDxpi861+Hx8xDQ0dUPnTQ6NV+oLBV347h9yt9CZN75RZEqYcDXMTh1fhdL
sFb6iJiJOdCBz+2vgA2N0kITi2oQwmLgt98UzyDYGFoJDOH3jvr5BPPjME1LQ85JbIRc1ddxF8HO
72I/rr78enp4Vw9ddXwiO/xcPQ5IbLYlSeNQ15M/8ZpKYL5VKrBRhmYZn4inGRKEaFp/I6MhuKIG
ZluKtg/ApB66SJXPqmAbZny640cLJXJTmGAFBWcAQBS5ynMg7RMDstMkDTC1c5x8NOtIdcxNCCja
q6WZQs4EG6n0/7k6rdu77zHnZy/RY67LEmbhxg8OG50F4kmEMJydrc1RO7ewI10UE25WpCLtCUjf
TKkeW+F3f2PCP1YN3Ky0z/3uA+KEncbBvN77mvR/saR8+2XOhiSQ/Ek6cJ0jodMFTgQsWslPrgwL
fwsRsvYfnVDn1Hf5TMFqdeeHQPL+EfkxBwa3XOLE3NDXakLTwiJvzQJ2b1J1xkq3DDvXr0z1Ah5R
bFgnkczkW7nNBbZ5py/KRKkTNqdUZWjafcj32+1HZRL4Zj67jrmfplHI6mznBpbXKNzCxqHj2au7
NHoWNIYNJocyQ150z4z1voLKRxKfkN/7lpPy2x+j0jfzh1vRa+HJb3jEdXg/N52k7ly3xfnnVwtL
/gzp+RbffWDvh+kHyq2pDHrCJV8UaymPsFxxlzdOkOCAG7Iv3I1XxIhEx+OyhVMokB93AN7OzR3x
0fGZngDG0RsdkBtdxoJXgQVOcP5KpkC3HgGc3heUEl+MTkZSus3lJvk95GTTsArNjmAwSnVLMvf8
ogFFiXdVj63YBr9bpLuVxi9MrIfjrMpccJ71eaQHVQQivI1bAjl2FLKc72W2jdGpSvf1l80mTKdU
S8Mmhxb7PXBBoPOLtWiPRK6jjgyVsnH8HBdq0icPSAYaPPTynfPkZnQfWEBquWRUUhm0tzpYiNko
rERr0ZU5jFXC49py9I3c1ILYkjGur0KgthGaOv2piJDawpXzV7nCzy2dOZ2lq5pk6kC55boJn05r
u0uYo/TvVTJyxIuzbmwI9tmeFiGZ8tM7/qJGL1ynENGzCihInTcA8b8s1ZTR6Y/XgcXyYzNis+QQ
thptE+Zljpp3hVCtJljbwUQU9Diou8GSR0KM1KwY1WYXYvf/c+pq/W1THJbMpWRPAJ/yrA2OuV1X
qW3rZcCBlIeeNYlN0qSY80613f6qu7bxDMxycbpq0d+TqnGSAMO8cWuVGVoBFahRlIbHYyw8avJR
wpPGQmoWImts2zNlg0/g0pysTDd7sxBndg5eP0teNIuMyQ0+YNwC4ZnOmKLCFNlMf3VAko2Z2Oy8
pcK8VCk74H/wgxXFng4sb5NjfMxEiESRK4j10JDf/5F4PvxbiD7Cw0y2aDNCRTUEKvucfZraAtxh
6h9ccachxjBvohkmcvyEgDeDA8Psf1yNIWurUoanBdFpxlbwf/n/Hz5LdP/hL5crFplnwtMBeXp3
qgbQaAy+eQkwBsYmpe2RTBnkeWrpEfyo77Zx5kDFz+7U2nwTkHsatqcakntaWNu0ssvT/Uh0vcrx
BapOsq/oPv/xGD2XCVMSaGuRzbQ31Gi4tczqGxkyvktg+dMXn8InPW+RF8+BUPjgbb32XaL8be5f
ghrt+/Fujk71Wkwp2MkrMiElZQM8bpfuoWthwMladzNQkl47i4OSWpt8uucUyN/D3NHkq+OmiIiV
RCh/V0TBT5nt4kCAOfGcDeHHUBpiMi6yHkpoyLVHNMa9iZsV28s4rIXWZF8i7fsjWdfIT6RrkeIO
vy7Pf37HtpDnge5NHKBCbErTHZzEc0y/KKRcoKfGMCjk013gig6IDyKnhEnWnD+5XPZ9g43TEwxy
7M88wk58iV1HU3fqSrwXSRvuh1I1EcO2HYHTQtnoPWST9AttO/6uvaqPSDNALSHDXdqqTjzeQ9Nj
BzYaZFaPazbNFLAo9E5fQm+pAEes86QNEpxTxmK4we3TIB4ZZgMucWvbRlap6oIWdb3yQTx9FD8/
tnGdt2rl1DabvqZjQl6fbuWld6DQcwF2TjpdGecqLMt3mm1oT8qwwy/3QQXlz9PuajIye5fcArA9
uHzsSOfoRCx6oKdFBOuYZtgPYZlSU7x65zd6Oq7Nl56Uxr47g2LvXPaptmH6iPGqSmJmZWMKGTKT
xDCq18zCadL91h13fk4EcDJ1u0r3kY9EH9IxWRrknHlnxSdN0qUfEh4MrA1FJKNF0N+/mhmiCZUY
xEyKGVX8l5DjCXo1UBTJsMKlsrOqkUuceI2aN/xJwBO4wLvztg+rEV+RApDSPzd9XDlsACFYjGWm
S0iV9W2TcEKvANR+nEOgioD9yhr9pl7ooU1UNouVLW7iMqPp+quh+LEKdWflzPMWpnDaYfYwC9F+
0cWu57XPE8plFb5tpQr0Me3bxmXydSh2boI1M4ZHV4yHti+lIWPJ4vdf5WeZLCad96kNIiJp+RIo
mq3Wic4ZxzUqNIbtTSOFgc85N1nRAfug2IE4LlRBZlM/iuHbwKwx5JDyzfWJV37S/MVm0EFm1zMt
EWD05V9sS4DBSLy+aI3Tp+NOFyh4ejIIvkfUKDoW3cSXZUjuQOXYqHIlPaZu7Gpthe39FfwK5ZUZ
pvKYajM/AOGXzbKLy1XcWIXarU+msC0Yhf4gouuFUJlLnpy+MBxkFRMirWYHcRaPaiXchr8Wlwtk
sDddI1hcc2XFkTOZwCfrv86TAUIGdA9Vdi5CqmPksHWwi05DF4FrZrs48vuvtHQ8wdkGGBy+JE0/
64ej/WRsUUsp2gxtLbLFlcTwlu8v8C6nvGZpv3BfftTSDH4pELT+0pPBBhuMhBfO93MrsVaNYtC6
4RqHkXSVrFKC5IJBW9q564hs7YXXE6LZ0TwklEO6rsF3Omv0DSyo1HeEL/ZgZoHQfPCoH2HmvQxw
Ac/Pmr0C/WK1GiB9DCPOFraAPPAjZs2hJ7cFaQXLdhn7ozIbFRQD9PCBGebpIuCQ8oQhVCzboESi
tOzz2rMHimLhD6of0GgU8Coe464wynHa7XUCIoTc4+nkVBSN0SPhr8nnZlFwb+SyRw3RlzUbauwP
NfRHfvXJ9qEDDLB++L6nO8Nni67DW4yps+tf5aU9Wbas3j7hwMgdzDu8tAXMy7OGsEeSY8QbJAcm
GCZsvIkbWwNdG6FVntYLKvZKwWTAjG4unckghagqo+yh5AX2R93wF97DwNK2NOYdPL+g1V0hD0P+
59Pp54eJcPJkpEsZJH565d74X9EuXeNt5waktERQE2ZhgeAD8eggxZbepnkqwMRiH+a+Pxg+Pum6
gGgTV/yYQaPGzF+jubonXFM1GVnOjBRqzRahJrp/T0tCi2SQXJBRr4zSinyOKLxhL/jvtOunGOpe
MZRkETKwkNVRt7aHaOTM5z+2aK517pv62npChx+OrDFgQvJsDoxOE2cAq3mI76PsE6z8FSvCnTD+
D1kFkPqul3rWyxkwnlKwNRWor0cWuTOfpHfc3XkKyh8kxLqRhHSiAXBNFoeRkVy49GB1TAcyOlie
m8B4V+yPmxVhv0zfDOXj/G8Hh8c+95krIitjmcbXyrYVU3cDG4HKFjQhYrATsiGMDrsXmyK5msZX
tmaoNFszcnAsxPSnZ/D9RCIYHCrXccGFAFQ6f1OFeDnmCaIEKz92PUafr7RXzX/VyX/ugcY91XLh
+iydK+/BbaHlufDKwBvixr4RkAqGqoF555LuCQBnfprZU+GoIcE9NVD27LyUpPI4DJctlA/2O6wc
FWxg5ukjpZWR718laWi8fcWvLMckM5IYUbmYnv+RxJ4FLf/Bp13a5bsXl0Q1/Di5UknkpN5ska40
CPGKPyqFgM+SqMEbwH0Z9C4NVKjEw6OTJGpQJMNgGPs84GyRHqdiCd5RNqY5thdx/VpQ3zr8Agj9
XEsk7HP/dcZDawJOyRLBOkcX8oQAzlvsXIjBv2jff1G18XjlaoaoKRqgvH6fCtYEpa5+DJqpSJ1Q
w774J22oKNX1EgTZemWNY32aGE2SIAG/DqpACSVmjtxFUnrNBJDgPbYrQp1Y31zTxvNsVw2AqsqN
UhASynQxVCAzfWhOid6rMHqiQH5vYB0yBfwAxjoCg/qLOJ0PJ/wTt7RCqhXxZTBrCfmW1MNYe80j
4HE8nmcx0Do0tcSAA2HcjazhmDEoEmxD5WZ4uTXXBGRwyPBW3/uW8HGL9tI8tpVw69C5RLOGGbyu
vcdGgYgAkpB9DDi9ZQqy0WUBWmMCDOhttPbOmlrnUYGTuciBjaSaRBizIpdeTh/fgPxviHJOxXOD
u/6jOdM2JyW49yuIZtXcrdwvig2lCUGaolNMiMi78sDGGOVn1H7n7/exjIF0vuIVJDDJZpOy6nZx
xvtO090NHwI9qyNjS4vNftB3d3T3ELW7bBHNr3vtUHOQblqjEIoevMqGjzGfob8cNpjAStjuw9JF
CD7GfFSLplk6xh/54qQuu8TCA1GQEc/VeHMtNZYM34UtPiIU6p7gJQwLE9YtvAbwUChLDg1/38wH
OEZAwqIFBps1HhUPZlmOh3ck/IrD1L6Pa6bjwr3JrpVI/bT1DeY+duGV9Ah9QI2Q6Z1Fr/9obETZ
bZk7YtxnLWoh2Lsi8nHc1aoOPm3+xPo5KOIgVdTfgwkxtqGo6jCjmdNjIkRCHXAGCt7D210TTD1m
JZCcHtUU7a9nu+W69H2bTwwtWO9byVq0r1J1qupfGoTSyLkmrkJBqe1izBWbXoIEHL9srq7yWhNL
n2EfHgVi85tcaNKAPOoXpVF4ZJTIfqRTBtaciwM0dTWHN9//gxoDAtWQ6Dsxe7S0CXCmUjcc81RR
sp5VLQdp+Hhjyn/7+qTezH90LGJurSJfpFv7oAV6jJmBSgsz5DMWMWA95BJlLws+tkZVPYEqFesp
SeGzcR+6t9qog8EgVlLBUv0brEbKA77W2Vl12f6xMAYLbv3Yu7ixcWlsh8tgKwfhNV741lNfmjgn
j8J/nF++RsgkXPxnHX1DRKVY7PbmnBjGK2tPu9zyi/t/tGnXKn44TcJ4+N1ojoC3QesAjAOxHXk/
Q0VBkHNMi5kycwFTHF378s1QQZ7YtabxaQMrkMealEFOHl7kbRz9FztnZWKu5jjG0tHhOHvhdN8N
ZLPmYi8++Cba9wJ7AXCculnGzteipGtF/Rk9SD1e+wLkaIHkfRabBL44nazmpdG0oFnh5kPYK0YR
iAzBgmarkY3IHJDeq3dvhB3i6OXsfBJD/679KpMEBV9fgykxwDz7Urx1mEpqQ68jEw00dVESe0Uu
t2Fwakjq2zOnXS2LNmTGyug/Kl90p+JYcoNpSy+PJxlDp7zPbqGIBZp6AoXocuR+BGXLN+vv07nZ
yjqpptJE+TJqEckuNW+kc1hvzOPzwOtjgLsg1dioLrbs17f/5qPcCP7uvAMYBPJxxkRuuVLtRU6U
3NlND2faRmqIOEz6zCVxHH4dIb2ikHLS/my7cgiSf+ZAvCyipjpraWHW1Pcm0tNXYDUeHF2IKKL4
L1tEvoQMkiihUB4yUIbbj+eHEbf+P9MameIXjozwkGoATccvm0781e2TSOb5TZJxs141qqDYJ36b
br1NcaYCrMN6s/DTm2V1LEVhz9eH1OFqggrh5MIchjBC6h/d4LoolBh9LmW7Vg5Dl4Mqb6ic/ywS
mdzb9HK02EXutSOZGU8nHW5E1N1O0gcRtfeNt325Wv5NXvPVA0m2IU0AbJNLZgQc6FbMr9ecsuhf
3G4F1ANHzffxGeUlp62/0akaY/+lUGhL6R2SMM6olAQFw2P5IDyAQxUbN2fJ1R6HCq5NObPrBmOd
4D7Zqn0ZnQEwjvZau1OSgH4SOEB+gXZm/KHVKa/xokeV7B/+lo/16Mp69z/WKIOSFGyuHNLySLLm
VJ774B6BC6cgZt/QHU9juJjieTMWUHNv8fsDIpzy6MtAgAgsWNS1MYX3wv2cAYkfAIXZbhSivcEx
0EbaSUi8co8jcKjBIMUfNlc9LkHCAMDQu7b3FJZID32Nf8UTAKepIIYUvLEUCSPbPnfwCFvMJCtH
GS9pA3G+j5xpUeADUipD1lgDJSaX65QuYO4CnxdWCmU8nVn4YaydEgarufKd7LF8i7VcT2UY+TgC
uSmahg97MmjmNa2JaD87vvi2ZeNO5/LRoOz6cRKWIRvSr2hXTLqNwuBz30pkvdi6azMDG17ZWGvj
L0nZksYVKpmcx603VHoHvKaqdqZianG8THEayRKdmFOXcXSbOPWvX6J1xOvEfUJWs3vv7dRZRfrd
YI8I6VXfgjJzw8kec4aGIPI3AHP5XEnLY7dJm521LQ7ZOWNml58ABU7hnLxk56k1Ju8ZOqvRNbIb
YwHnekNBkjgrCtcvyf7JgS66LBK4SqdhrPZTemyQl5T/6W8Fq+kuvQBVuP+QDTZTZErFTquJUgua
YQlqXttnpLuuM33ZKi9dPc4MzazI5p+b1Cczncz9erwDyBImtYwkAQRn/CUWs3ZZQWQYYwnN2MyK
MP2A8GQMyjSZTVAWEb6mIN4fLglTKMCDILOe9GUeKX9e1omMVRu5de/kMMfWwaA3MYA0qF2wtQGH
ZgjydBB3kIqgwKGbGPPTLvOxJ/FWtKR23tZH3fl8lnfDIJ1X0uS8i7YtWdvj+dnocAw06Nnw2E0g
EFB9l38ukXZ7SZcYOasIz5ZlJ6uTADSEjxZbziXxd/46tvrDrnVC+k+M7MYcX0rUVg4dUkBAX/hA
/q4X/qE1wcn4phCnYYbbl1N/TB6FnR1hyQQA3UETrJRFo50E6HCfKsHCCbl4jdkoR6sSwiTZx5d1
w+BrRfRB+4NmYHe3Sp5o4nXHJG6g1pdzmgr/cS9Kpch7Xmqdj0cZqvIghil7ST9v2pK5GkuwGXGQ
h2hLo1FQpN418YDmmo4+tYoBqm8idtOyNm6im9Oi3Qy68nnv5fLx38viRkOobtZLMoZt8F+mh1J/
B8flHAGn88Ynx+XfWr4a2VRc9u6vtlAXDcbuhyG6zpblO+jldqlmSzNHBL5bomYJWRDbQcWhS4bR
gV/SH/MSCqDMfpIIZ1iJS8aomT3QbwUpq8d14VwonlI6PR9iKnpZveBghMOzOhtfUeoyTJN189HA
nTHQjLMsU7DnG7rUbE8QV2eEXejOlOT+gbAvO07RDB6nnKnCdc2EI2+R0DOWvPRmA/eXLC/OW9fW
8BRJnCvu5N9mReezKWLzy015mmlCfVxYHw/EaxbQF2atE49bKpL90oMCYgZQN7Wc4/KAFWKq/yL/
WuhaiI7KtItTLawufAxX6jUofgyDrVwaF+BTi4ZXixBAOHl839mv67jrfRpDJuJ34JgAGE+oyOuH
1jf4SpcC74MWYMqIkr8hlBXKsMON8vGAKRuaKDtH0I+E0n7847WxXRbd30khiSAJeoU0y7s5VYy7
t7vqpQO6Eust6RRBIYBaAPX9Acw7MiH2/PyL7e2I8s8OfU4iQ9kg32kXrtcWdrZvrK9a7oqSqtiy
UBBT0+r8K3XC/kKeFMQsfuxEJcUCVFrFfLx0P5Vk7/cUFveFLVIkHvTXyLETdKv0P1yvUBhii5CO
1khMuj45oiKPP7UMHoLV93QvHEIIONcctqt3frcsr/wfiC7suk6bUejXGCpHCjHxnpQvVqmSovHh
iwpxMZGkmXHWAV4rQshgibB56k3jt9IiW3if8AH25wy+ZDOMM51+wcsAQGqpm7vZ9lBjt4F51qj2
T7pAe6tvbhEdqTifuSxIXTMqbD0dWC8OvU3ll+x0HIzrQgi5MN7RsD6rSQeQEBChADtapBva+HSK
dbB+eilts7qpyTxALTNdZ1VKMyG6yCmtij8iD780fCkEebuNs4MmplDrkavj5VqlOXbEtrVu6wws
tg/mrKiDM7SZ7alQia2sC2cxz+vzQFq19XX1sSdacfrmSnA2HFv1IJsVhmKpJ+47PS0oEil3+FWv
Z+x+PiHie5NdRWXMLWa5NlXx6FdtNJULBS3/Fld61PDxAYrepsKL5nyTqFKpmPB/jJEizOCyKave
49aj3QCEAAwc3l9MM0EY62RVUtSxq7Q7WsXTahePYTcGSXOt4vB4L0OAt7xUDFqolUHtqpEQLLLw
N5qchylUAYL2wnuN7jd1DItvCUdzx66UdmWCVUz/Fre8AcE9zXFtJXvIw5S1g5K7SEDy/WMmaHpz
DVnH4JJ9MAIUbNUupvlNFDQ1VCz1BLxoUrc0v+Hz9PlARWlYkELIRk/w+b51BdHN5Gs7yHwR5LE2
5cpKJLPjwtLOMLzFcZekUl8cJGt28ZnWipFlQ0ygLiWgprLWjtGjvJoGjF2DZMJaiidvX0SUeuDK
UXAX1b6z/LFIBC1obBNcmuCPP2eCjXzEiNrdwh/eivdRmdFNTaFhTSPWrCQTa2d/ePFk/WryIzmI
oEA94ZCH7e70q8z1E/wY1dLN43I5BmQppjP6veW31dtDXkR59ATbn5126aqx/1np8nvNZNSK2C3M
UN6qzev7h3sa+YYNapz66pfaKJJKXySa3VXgs4FqPtu7u5FAZ9+vjy65R9joZxt1IKTdnHc8Q5A4
IM7L/sqJtmuYtv9qWyG4gRf0D6l60V0F7zSDy9a828YGCIJS+cAKwyeMpAxc7Iqo/xpf4iKPpJxH
LBnl7cOpRtoQgqbsv96HtzLPx9PI/zy6Guc8mZRBto/Jpn09My7h/kRz2mu1v6gUbFsbv3w8NoaH
fwLGmva67MP6VGRWwgMPgfDpaC+dZhPvD+CgkVmoF3B+ZhgeA1628NxmQknPPzHhLi0B33CSiN3L
3c83KtIkF9fciDNI32lETKJgj+NAb++t3/18gy+v+Hnqu7cA7Uguv8+P25cOX18GbVKupSnesXRQ
X3PoOeN6kfRmMVCsP7wNL4Mfzx6jz67mRCduV/OjX3FlwTGfG8Vugy0MlgZXLAmY+E6Mpfs9KPIv
W/Qi+4tL+UQtWZa8a+kue1a90hO5176B57YUWXOyrijJTIvViYhGioD9yOQzgAWJMVJAk3hkHtcX
9DcEiCo42FK7KWip+XxcdAfMEcY5mjOtlwBB9yhm1JJ0q19CMdcwzZ+Dh/Pf7mb0khga6+FNpYQe
6wO5OilvX4mC79yevvvkozAZJa5Bguq60nD+ct4g++hcKDNTiMJRY9TyKkIakFb8txJRC3A9P0TU
99hc678NJsbtQZSCDhyBU/5MtflnYESOKGRtuj5qEZBX2dpoCYrAUfJ5dL7yg9lapkKZFdsmZKQv
EcRLPrv81oc+OCOIrnejp8a18UuuHXke1DVI6hJhnmXoy2pXvu4zQHFwZO7RgRJdcPLqxEcrFHKY
WItVLGUzaLsjCkbUbBHt7arUjkRqySa3/SpH1p3W7y3QVz3G8D2xJmU6zjbnnXrUtq4/nb1TJ/Dh
9N6DZQr0j8KpJGcuNhopj4JH29HfpntsHrcEoJsOejO//5+4G8JEQ/RZUSdRsuUXWEwB36ec6mUv
BeTsvE0WsUer65N7KBePaoBezIokOiqYJ0sFLiT8bZRs4VSufPEWI/hlgW8vyafOSmAC6dK1rn1h
JdHxcJcEc2Wqvq4zjGFYBeQrFtt/w4aeKkfibuOkxbqnjgaLdUWIxpbwlmBEY85XItuMREfJ54zv
tKw74S2cyTlRxveL02xH7E6g+oZ4vJHpmfB72MSwjdH8k9bOIxQ1SvkQNDxSlhU/0zCcWLIyyPix
uiSaiStg7jFIWiTa5ksJxroDTvGniiuaJHn1tWXHiqFu0gbySEA62gQSh5rspgG+fUj59/A3M5pX
laFQ9egMc4ONTvbtSIgsD/3kdqKGNg2RGLsy6F60ZLScpQSXpqqqMx9+AEurQvC4af4l1Hd3GfKH
3n9FGJpnizLS2vSHRrnKPRZztiAID6HfgHKXkvV+60+bzsYIq9uquBNfE3diLhZfmoth4WHgB0nE
3XVrPmIefSwYNC4lqfwfRt0RGZg8FZCtMGDkbUO2wiAqfonftPsdsn/Rqmw6juRcui0rZnAdbyyJ
4+UVAyROUwlZPlTcfrkhjyhtRA0I6jyMVnP7sDqurqKLNqvf122hjYy1qIJOHapIcx+9IDF7KknA
FdmCiGF+JYxMkksMbcVVNossKsF1BNx+9wVEx1NOJQm+sISwO1nVYiU6t99ClUGh6INbRQW+A85s
apeeLkEFq8fyCmZY0i7sg/juGBoKTNI2GMES35UecpHLgIL5DhHEbOpieXlH1l5B92SHQ1HLo42L
gT258LPnW+k393uG9rSbTqgioNS2W+/DXpvZ/C86rz6AtbMKB9Nl90D9Cz9K4qHI9FqLY85kd737
nk+gitjfK5VMn0i+nANmZJYbUaVmu9I0xKGXoHQcaFPiWnWyxqrynB7dUzWsTpWl/M0472FDbiuZ
8m6BmObOh5xWVLbBJcTSGIapd4UhnHrmNRXoF8SURl3jwip8HTaEDn7SdOqFhXY8kmO72/Mxkb/H
Dch4BsiUCDRSVG6lApkmsUd3Kf/G9tSqIRTVMXJp/7kCh+xfhEFizG17e79jnQve0C8Qg22cwSzT
abc5iNXm0Wc3b5QSGvq8gFNvsqtdnxbONsKSt/pruFhNv1AkCrhFNl/SW+R1UrxZTCKTUg9QFGoE
lpTPmhA8jPmrMwf6m1h5v0EuIU2fY3fIba7u510ll5xeJ+p5l6ky/Hzng6wJq76Nx6rO67RQgojV
+n8/gqMH52Z802hHcY0UKnK8iW80DPAaviR+nIRL9Jpr/ZhUoXa8PDSUCBkmHfNATKE5t2WCwipb
c8w772vPdcDL2Nq1U7PjQo9sMob+tjylKUrb23Zt0vJ9MLqkMBhw1CaVFSKSZdWm9teqNBdtewVi
AAlFrWsY/IKGkGO/md4z645quyazsgIdFnJYyMCtyEx59c2vTBC6xYxgfhPYv070zDafNl+fxJHO
GjuYH2hpdfUTxEqEVMQElmq6a/XjbhJ35MuU9QNhfsfO93/9nkhv/4uUmjYT6Ey/RbbTVP9xDls6
9mFu11CAg8DfQqEV4D75lU6ywxjXZJ37ZpZpei8nTPr3xf8eL36nK/G8/PEUAXgjRr79wmXHF4oH
eH2buQa4X2fwyt0PXb278r3lc6tAj0UnSTwpT7f9nVGCCf3FHfEZg3UCl4UddT0RcIYDBmaC9M0/
Dl5Css3NmxhM16aZnRKq8goEwKY76hD1HwessSC1iDduJ6mOm8O3nsaTqjOo+4rytueirTU7IRVN
bsb9PybI7OlZlVlNCf2HGnmXRIyqrWHl88hScxfnnimbvaOTJGJaS0ndIq+/vH3vwNWa8f1khvFo
kIkezoglVvAp9YA/IY1IUHnmhtWfNEsop3RD+3IN87vOzG6YLPE6ONWsh62LPgXSHmVV1QvW0xQR
hkKUuqxKocDeLcn1X76imRhujkRRYBR780KzTuc0/hRnUyR81R1C0W81+3qWcyXOw4ugGkVcoqwN
wIXIfLsnETAnM8j2ZcZ4f4CRifNtbcvfHnYDtReGbZoKjhaD7eI2G8ll65tadA7O3Hpd+SIdmEFD
fhfvMr5CZSS8BHd4Pkn2qjUs+ve0BCYKcvKj2ezTY3jPtSVTTHSKbN0bRTRpjsYoVHSa8BU9cyXd
p/TGqL8YvaqiQA6I8mmrWB8UrKKByeo1S8O23zQD3EJfRG0fBNyAK9HR5hjc7a35FNS16jQBom60
AmwZCY5BUBCKwxEPrNa/6JFFP1vB/8wJt+GFKC9vvwSzyALtS/HzQcWB8/a1/hBZHuD/ow3Odebp
MPEraah7H596+vAvCIi+0mtg844FBj5mlJBnvjClIjObpgBxkCxum9kB1hXrUzRyTNrq8I7IAa8f
+fbdFfYw2ks2t9XuWbjrEB600Zo0TiNNGPuzMPigdYCo+7XQ5tpJk3RzoaB8Og9d7k0Cr3yCsEsD
egwsyJpGJWxBR7c3fQJbRNz/v9IYWA6vhdbAtg2d0tX2o2kTSyD9Lx8nHAv2Hij7NSHK+9gyMmUI
m7Y9FkKUWTm4afaynmTvo40ge5rdx4qW5SKBjRzaNTfjHbTIJLi/+K+5U2Fz/JJOAUy5KsCZa4fn
OOB02q1hlvzskiLTgzznAuiKtnqkcCFXqx6O4KIThrQk+73QeGl3ZmxfQ9mxKnVu0ewvAvBISolj
2YS4ecbpLQuQnKz9CbmQA1Fvv9pOrieR6ok7iZ9LHAXTPW4F84nCN0ZkinhRWPv4b3EOZ43hUVUR
wC8pfuA6b/OavB3OC2M0UvARrVC1BnPTzI7wlaRpxNw1ymgwvVDuQqu70XgijuQloD+DCYaqde57
IOb6wDUOy2yuWp7sRil8YGLPM9yVpe35S13uvdMlaqJK0us38YKXOeqUcbHWBTn0v+xvZx41L5D4
56LW8X9hMLKZmOjsFGHOj0tBy1LemBlHuDFz3N+AGQRyyf9FqWrsgYfChgHBLsbZu8ue3/Abvi5H
SxHpp9FDXFcDk/DcDBq23CmlTEhzOPZOCp8ysHAeS7zsTe4ZRt0UiH1lbJPUOH7/Xts4p7U6aPa/
sb4EvDZhpiDTOtLe5QtHZlnQmsAIAAFNKqUEL25g+ZAXT9cMImo/e6VZbASS5Za0YFsvTNFRx3qY
p99ih1KjUM5Stw4esfo+hrIT+glx04Rrmg6wcJtQlPD8Xv9+2HYVRtFKpN9pq8L43UL9Jkh+bkVS
JdZ82vWg6bAxEO6YcLa4MeaNQ7b5g6SWWgTKJmUPN3HResJFz3G8TlBsmYJ6zzy/sXJTFOGF9p+m
/6L2YEC2tUxpEP3Wn4k/jzH74he5Ykx2XWfdmgGSJWghpUAXw7Kfq1MN8Et8XvwAwokt5T2lPmEJ
fS8XD3dasWSf1sn3JQ296V2bMwDDSLVBEzU9gPs1YDPcWwvaM46t+UIR+VbGem7iOUeMKSz5TapZ
fL6Mbi202IsEdRZkCKbvAY3+uwbDsG4QibdC4ooW0Qri3nhX22NUctp1++KJiyDoBOineE8QYmlK
rp8+GNlcsSb+pQT5+yM58bKILP4eBrsgXz51YHO3oz19UxugbvulGBpyaAuApTsv4E1O6jy9cO+O
lsWGzRj7jVPns/8Ibg1zIpU9R9+daVkIvA2C6wo8In0uO+SS4HlzrvMVeV5xi0zIWNWsMv8hJ1wr
xbVSmx/YcaXqd17Cd3yfYKStkX0Y9v8HSec7Ihp69n/0WPHZat7lbv1cpRLTyFqKmkNYb74uD092
LGEMKKaPZOuSXSpa/gJ1F4LBcGuju3HEBYNo1YBIDtu93Tf/GuHV9aWPdjm5Wy/wpVGQAHlsYoNX
QLm71sd8wC9jO1+u35CYsYi456K1HThESstxVMt0IAlaWKbIwzpTe451gaRy6AyHTBt5PFjjvsoJ
Pff+GUv232/mI5wmLij0ikuntnICqrtPfqgC2lrJbm/+5W6oOAOP5VuyiIpCaFQiSPFzlp8l6o8l
VJYMFNDFjEtqni95iOuRHYEFfza2HaG1nw2RDWRLXyMBbZlhlEmcpN38GaKGhho/a5ToztJUxqaE
wZpXs38heAH+hoEnFBuFq897IcXkdfLVSdApn5FNE/sTAiIXfsRqlq0xpp3LhZvrULVYxI1q4cQv
ZI9g2qn+iX0lhzBGH1oXyrWtTNilkiPr0rS7lTa01Z2ewOhR1qiAULOBGDI9p+or2iWCuBPvZUiZ
mrnurrc7/rKhDqS95Svc9PKFNaAFJ5efjvCKWFFSd2zVhG/DZDYY7YPIkOxrxg8fx8keYdj3vH8r
pJzWLjG/NMXVvpDntS/JZ6wPS9Vel5isL1gGm1OO/62O0dL6CBmkqUB8aexP3vEVpRAr2+w5Bohy
Xg1+GvYb0A6kHmEm/2MH63cwVymtDRnZWhpafmosg9FxwDMKA5kfiE1C2WPIQGAIRjMTjaSQVKpR
Ra14V5bKFfB7opTWux/aLc3K5pf/w9nVOdluuH34s8E7zzfir7ros0rx3jYeZV7oqxdM09vi5Txj
oGiWBiE++yZhDB3KeMsWG+3OKyZbLVPiyWUazy3FI508cb4qnpws19jLXc2nzWTTZ25ENGBgZaud
7vtGX5U0X1NcU1OEsm8mWhbU5RQgkuybfLO34CiYeyzeFMLMt46JTPlDTlFsAyyZQZLdXmgotiv/
x+C1peRXDbh13tBluHB6wjKgmuTnbmG7EEoR8QJDH9Ws5JZOh9tXrUA60Z9V6wU5+9k5SpfSZbym
RbbkLTfToYcchZdfrwInG1yGLn8OpCacSXe1fvJMrelyyJOWQoobC0cNHgNeeCm0VdJtogn8j2Pz
sMey4tLWmtE+EWGYVw2nZh+SmVB0aS75pZ59VBa+b9kJw/1KxbQUGGRn3sXXfSft7GL3u1NYfLvJ
iIgrJcjCx5mopzIMXVHmhSwz8M8Wa3CmPFQ7NIJqqJX+AffJ4jXtKyVLNmo8yoezydzCcFACYkbi
UsIqbJFkUKSZ04NlHTU1tNhXoFmDzjEFM87gXE+r20n5J0qQymkl2TKgIaP+3sOucMqD6TyTT2Ii
98Wp/Zw+Tt7z4ZKzMTQikqjmoihOpsx2H2SvkEEkmnkERssuiZJKjEAS0dnY+7HN5BMK9Q7wZ38z
3n+mFJq882TMKKSSZ3lRjkc1m6RrS/siczMwVW0ghJjm4gLbm9O5HaGSEccn1Lo4oF8e2iQIIRId
dLEZ3Xz+wqte6hyi/BxeLnH7uSoM3hIErTGjokcffQUR8QRHtLZOh0of8DGDOiRqiLJf6Ee7HIXY
QksuJilSfJmbC+H/7x8BvSPC98iWGT0ZS9NUPHg9f540lli5/TAEfPNIMvwb/z+D+MZvbOnW+uu5
vgZupsLLwJZo0c1ECbRrBfa6AZjDVcYruL5Qkh4UI3fTldaJppa9oClhkIKpsiN8bIQ+j6KW45X8
irou4SqdkpByUgTu9dVBGcZ+t0hz7d962wj4XiJu7DlXqJK/qfpaKWO90c+q2Ubk6l+45UgqQ1O8
tSGZ6aZvfX3CjAXKhjh6DBssZPozFLYob1V4jbCKauEs0yCauI7ifO1fP5qMxD2LORCp08nBwY4F
vRcEuSTqnsq5hc2niFVbHIc2gXgFzyML921vXQZRSXmtRbaj2p2UTpJZNVRGnU71CcxVUqvNj8id
LHab5oBnh+9yd3XkTX4gufYYPuQwugS/YpIoL6v0ebqFQcioPhECf2IzRG5O/WsY3W4BPBXSkPz5
FZubzVSvyWoLWKFkYKaWpa0v6zkUjgUF81ZLBL+cW/hV809mBpbYfJ8IKrR3L0oOArpOnSgdeNuR
epFes//FwOBPw3yUQdO2W33Gl93xevvd7t5BHD/BDKdYvXFhhgRwcGtdQ7eM1ieJxBTdFrZe+JhH
xz0BDoRJkL2lFsJhVmgpke9gq5GJJJ8Bxp9KaA9U85uPBUEZOnZFzLDNZy2lpfjiNOSG0wZMw6mj
5wwO/XZpGbulGGyWOflo5KWNBZnS32+Jv3drCQwJGmjxlONNmzcPruF2VoElUiOQbKxeqipUf0HQ
j4pzJP0IuB9NCzHz3zEi14Z9qLJ/1KXKpAII0M2v2Gm9Jn+3FYLrCvTVhaTdKYzISMeb/WOtDmD2
zPajr900PEiyCFEmnDpobt984Y2Q9tkGJGgvIc5mmj5peTPElKXPV4rBu2Kx0UzwcVPdG7CqVO7K
/l/4Dd0N/ekyP3POx/dbSDZvZXaaSuXhMZyIMahVU309gOjzU7WNoHpb1DEmMzawWpHER6iXmJ4p
3ToonqcJU7uQswE7YUE8iS7PlycNcSjg1wUwpYnNb6hS4NpQEYRA1XKRQ/gn9bVcQ8bUOVZ0gmr/
ZlTTIVyHy60ES4TangHYMMdkhEtEnOvjxJ2oxX5iVlqoMlvyXLHGhH0RbLkJrp2j6NEwyv3icDwx
XhCQMpVtSG0u8W4D1w2n8guzGbMRvoQBZStxoDINMB/VWrqI47S4JXoUbG2apq2h5Bg/zOA2UzGC
0Xg8t5XQdbjyHviA6EuWEIJxV/A5KmxQ6Vk76ohGQ+XjQIAUEsk6FFCl6gqEfW7ebJEhtFUW0VRg
kN/O+Sl5X4NrxRBOmKfaPHXw6fX14cfngXNp4tX17tPCAo+OT39s1i4XVMoOkv9q8+j5uT/CxSxa
uNauSlnXKxlLIlJYVIM9lQ17a9382wSKIMg+jMzI8yM384Sc4jj97mdugYGZqZWtRAH6euuUiPNm
WQ3lM6AYY80zP1IT7ue7gzoHuUZjLPwCfJ2JTK2hiHQpIBpnj/G+hbJzCgvu2Y1IbgvoaVA3bwpR
3Dc59Kh8QoH89bbO/nxjpJgqo4UlNlDMTemt2G64ld6q2leHMh5vzjyd4XcjUPLUDGnGuO9b6t/k
0QBB9vvPSPhqaTXob4BCzetOmL3Izkal3lVquEQ4WUdxRDSyLjIeGHlYSvwczWLuJ05tCo1uPm71
8w6zIW4VuxOaNwIexdRK6SchuB3O/cd79PC8rwfGxnyjxYzqAOFMQ3e0tlSb+qzz2VlG59YQ+g0i
yM3fTqarKJqhSxOiPe754UwM9CqMcXDXV1ZADZ9iORvL3fEhCD0gtcuYKIRFF2fd/Uk7KmY43Cpx
dEkSaWIhYHE7zkQHitQsrPAGS/d4ru0CYKaowjnQFY+6kmG5g9kAMS/OB7eMXcfIVRan7e8u/5iT
Z2MUdolG/HHYA2HhiCFh148fXwORMtRflSdJ59olMhQBC83RVlxkHFWBpyXmCatbQCyzFiVIynjE
2ICEX0F8t3s5oIJjJLkv4GSTZEazXQFp0aEuof2uoOX4xjLq4omRH820J8hvwi5u5kKThGPp/mfn
fBBHqioqJy4vR73Lwd4FRuA8dFQgmUoV1VfAgGAHh30o5i9BdTSj+6ufaJPKv8g3WDpRxnXHd2m1
M/6n94fn3vwCwj2pbk8LnYa1ub0zfspFaIU6cZBOzsQq5M/7vneXsLtfKlF/v4KQGquSz1gu0jRE
RjsSLx2omeByfzPSfKw2yB7cB3eXmIGbDrw4yhC4fURXP3JfPmHNyZTs8tOASmNCXDhoLSNSNplp
LwfxBG/N4nZavaguZnqFxoRIHSKtyit+pn0sFF8lAK5zIPZTBF7UM842V15H4yMxBVBjc/cUr7wl
zqXVJkZSqGsgwOD08wxcMtqnU8CDHKdVzTExD47eh5OH/90JT6Z8hUP2tY05Mg8FtATAPQEmqjsC
oDG2tXKHYJp2/onsY4f4lIeA7HY5qJi952capHshp5m2TtwxLGt5H/tUcQnHyC3JScEeCzx8PCsm
+zXK36Qft9Hei4mN3rE/LGpxkvYqtGOIfvujiABN77ynO8W3SvTYOWuqfM2bmO+rCBWv8NnPmcPX
T1tirhL/qxyv/gZXPMYcnCnJDyyUPXz2yz8NewcLVokiiU7LV+ivesnRjaQiibVN2mscwP/7t6PO
SgjLhwRVeUuwQJ0XAqrEwq/kSZGLQkwdz2OVZV2PheoApvnLNd/v8rOVb25jSVy6HZ5zliP5ClaT
wvSPzwxY9606H4bSKHSMpkriDda05zWjjMxYV5s2YJUg2uoORQGuvHZZj7TN656F4PhlBseCzONg
U4DbjPdTM0cuSRwf5Xh2j0h8L4l9S/oZsFSZ3Pehq8Q24iAIgxGXQ7vixN05uYfpWDXeb3ySuT3T
4d8xiqH3xdvLjmaz+B3YseVFQQKaUKyRK24IYmo+5XQ+2SQpPACfM7ZOhnj5jXVDIX4r/xckktsd
iOUNC+IRWClfwb6o9avCMHMK0gtalVC0SZlqF6qFfgBD5dRrCBlvqfQcLX5lBjG6dSe/lm2NpRyf
UI+oOhLKPrMoHWyY5HdbO2OKk1T8YgarARcEc3o4gf3q3EGsHK6zhbySfbU9zItmu3De29M9yM0V
fscXHPiu3pt5HBH9m3rDiMf+3kyniVfx1IRL0I7MnDKjky7XiXizRC6WRMVqoxDcmzSev5/N5enn
VWOyFavgED5xs3QT3xf2L75LMWp8s8PGaBQR8D9vGqq8YvyzrloDsLAavQjZOPqO2k+e6cEHW0Oe
Jrm4csgEW/uohxuQ9CcQSIP9+TTbK6B3VbeqWE8mfaSSguxmHRuUvR6g8AllL81rPXiJv+ObC4k/
8xr4wzHGAEXPklT7++4j3zgcCHET9hePOmwOuhZZ4CusjGyN9iUMDOl1opz4TRvE3FmTlDmllGcm
U4iKPJ3eSBd7FXkvFD+tvZE8lGYk+riH8T9L5yEchpNL3QVY5/HhPEWM9UBnkcZ7PHzTbadgwD/R
6TcIq3WzfvVYMGdFqjM5tq8GgWiV7/WozFiEzNxp0xYNdus/b3BGevTktprDNT0Jvn8Wk2iPK3o7
8VQJK3KzNpl9l3aK5ePGw/4EsfM0NEidHQYpOU718oRAQ1Cv/IlYKEmXUTKaVMIHKh5e4A62Vc78
kEH6jzZlKz3RuaWb73e7AYx52hbExDP+ZgwaSlx3Idd1uiDfYqvkgvcAEQlad/sR5RPNe0DBIdEQ
70RTSNEsn0V2QBkRENSJ7U5HBAr2gbzlhwX4LOsj53Exn5LfSpxezY/Ofy1aiYpMxETJbUBhcmUj
qWKJ0LjXjgVBzoJXU7aTs9KHnIiyKhQcvWwFPaSKh1Fb7nAiER1OCHhQU+folPp8OkvSsZ9SNfRX
SaYvXMYHFbD88gqkTj18ThDuaCBDR5wS5DsdNnv/rmdRyzrVQXoEZg88WouePXdtOGk9/iD1UIio
I5+MVw0QtGG97Jq2pADuxGe8HzrDO/c6uQ2qNuoKWGIN/rKFrApKPlwOTALO1lYGrIhr07IB6oGO
HdGBtdmDvlU1s2b3QjY6vBLl18hs9YfuvDilTSFqX/F+YVPBECkMlGYWvgMTz6I/bbALTlSLhY12
3KjkyrBUpF86O2QycsE3p0f/ZqCFy6pXBq9ygyBdBlFH3VhTzanxa9DdsKHdA1mnI4yP0kIplpgM
UH829p7UagHhLpD1mXXLJCAYxGT6vPGGfacvfkKQGtHPnzJGVcNE4YWjF88Su5dGjRFWXCrBZpx6
z9moA2EMLE63f97h52yQIX6AY10daGKbt9ZOk1kte7MyF4UXxoF1DIDJc2yIucmUHOnP+nkHpJ5z
VKnL19C9JVMlO+PjSELS6D08goHEbNHaB35iFsQj8wvHL+vchQn6K9GmG4C37UK/fMs+YLRUh5ZA
o7gdzBsgajjfSsIR9Wv+q+B/0vzk+enjrg84LYYp7BU5SjtSUStSZ8zKfucZ3EzkxDwU3QZi6Bbs
n/ZJLcd/xWpt8CqGfDZykTL8GM/2l94dsynS66EPlBXKEKFPNEmPjH4FtLx1BlxqEqPt8JAn274+
NRnKFfSEIEoORHnzlK/k4eJqOTd21/KAoBZ6F8f5HHjV7yuC+E9TGHjx0GBtHgMvkAYwpSeiJ2B8
4hfhhwLVnm+g3P1Pnu3Ur5gwiQ9LkUqL7HmSQE+olqrRFBBcZGqksUG61fiEMqv2J71fxgoOvmTV
ZA/1ORusQ+hdlTCIwjRRfaSwBNkenGxohi+u+5BwVzXQUBAPUC1SVlP+FtCnLRmFo97/x/dSBw3A
bxY2X671C5PbL11Al/SsZe5QsrIm2/8OfKunSsW5r0DXTfQDfjYt6S9LX3nURJS0rAeqWaV1IUuA
fZxf1XHywITEdmVypn2NnuKdRIl/BZW6+0fSTRiVbNyGTB5ylhXsxbhJY56KMjKNDwzJQ9tjV4gY
TQQN3cI2z967GdTk4FfcOIzjJer05F63p8L9sbJnzaOVmeVY6xEmI6DhhIWc1ve3cxXq8sSZ0IPJ
k2rP8A/d9P+1flu1Kmp9jqV/S/aCMBJ+Q6V7HosFk6H8sC0Za4yAznobkM6a54eqNs6mO1fE//bH
PD7ea2nHjuL/kDUOluoe8FtOI62K1ywcTkZXXLZCfCjJamRaax4jk10uaHAoauXk7gplr6ag+nsS
tkavd/J0uDyOuvorRTWKg6fGm8eUyeZmJxyK8thd+LMVOAjGvJu1pb1DNibhH/ushboJXyelfN/J
QkSEBuRE3k0bCDXU39p0OrRaLetNtgBY4keyL5Yw3S1+fXagTvSlCBk4OrTHbHe48dwzvBegfbaq
hG62jlTql45Iq58xBWpmSmZNgp3c7jFWEJ3ZohbGZfb5J3vYVG5WqMl6fCMm4x/bDtmQdQPSgayB
P0EDuwiZ/phGEZRIOnHJKtchtcSX1q406DtBxbj4RXMDyuHyTDS2R7VyyOeqWru2lm1BPon1jfbC
ND/8eO9nMJzQ8/iybxlQ3T2JizYNOAqKGMfdEgW/wR8FgoSMuuI0Ei68Wxw5j1DnlxW8LfIA2op9
FPw2PV/O6AIkjiODBRTAMnQAF/CJukMziSp96xYlxrRhzTarKD4D111LMCSHMzcENYNWoE93MFf7
rtUmoHwyTjW6w1bDkfvtdSvNX7H1+rqpDXFdXAars+5PQTXcL5afLHZ6FBzKWEKiYInwhiy0hNJc
hFQHpsI1JNJQHKU5bJIX+ZsXDj1KUR7kRcLY81NzcyYcqX6xe4I87vflyVURjp4Bkfj+uZmyBHxu
IKzW2FWO91DTa7INAByBQ9rBrVkg+PhkJnzfcaVYJuKxQFSu4BzXvF5wcyDyLyR8EnVZbQP0N8lD
JWVQ2FyM4rxtV1s/UC8EnxaTgBhawLkqVvOpwIg+0SVDMwhVKxANVOw6ubUWGzwkBfUQ351haGZp
VKkMnW+X/ygMWGlrNww6wRmZ5qA77Sp7px53rSCfPQUUxcY/bu0aakIwiCvz9VoSRi2XIQ7C9sOm
4dpMNeDKM+hA/0oguv6kaAKZPEgiVca+y6PqCbVs4LWPIus90L8/GmNNwyVFeod7k1VtyIqR0YQo
urzBvL/igSMNYoz05K9CKAQ3CKMNAbg270iGlanFlXBr19dF2vZlPb5EeWI1rsmZG9L1r6gDDt0d
yCNAL3RPy7xbCY3LaoU1otC/NyPjz7XU8bp3lc6tC9lkJcK1P96LBqLx95Z89pRQzZVG6ACJFAS8
wZSpe7aEsRadJ3Ld4nAgVf5HhZuTw4GUSgm0iXOe0+2GDbvqsbbn/wt3gpxlLsmR3Y+Ewun1Nr1C
WD8QC+4asiU6VoCuR6/2QksSRdPmac2EL+GAXoFDoV0W3+fBWa0I8oeXgIkGsMyhHvdlZbM3wnS/
qvsiF8YLTcL5pZLMQQtVXieRbQ4QA1goUfJIKgpG1jssrY3YJHyAYD8vtpiCQzK/AcnXtvllGPRI
lQd5gQcGIZfzU5WjGmRSx5smcBCMKjlpdqtXj4lJyLlU2EJ4pToiWirzvKeWY/j9AVLWyWOV/fKi
szvcpsgGhpR1Gs0LIm9aWptxJauYcWL3zs4rfGTeAD94yp+HT1/iquOH64Xp3NKwI2jtzdCAZ3Vc
ykgMs0NGZvz8KqNkV8tG1GfjJmG61hZc3+4Tt5+UxwX718NYhzW0kidn/hWZ+bG6QYEY28seAVi8
bZRsko/UKBX7aXj8TR7kTKU68SiWy5anA4b/e/nE8ydMpOuuE07Zl2c17HDv7L6BIg1TbW+u5Rff
nJiCYP3fheuyCWEJkQ9JR+2Q4vMc4ka1+hkhdTZ0EizHk+fhITzonxtruvIsYVsUB1TDw8Hei6d5
DFohj39xCVAlIZtNJco3xhgx9hVmEygOUORcyhxwox7ZgKN5xWZPJf/Dzsg0i0EeF6rcoDF4r0fl
JmHgDG7wF92TvwvsR3XQv4E8B/4LGo9j3cwndsKt/Mi85C3cCzsDNLwq27RxRrwAITqUcUN1XwI6
w3DAjhuHIIcvFQWdHK3TRwUX9Qf1RQer4gCMRFxwaFVIr6F4V32N6pdcKB8FVHsuH8E+o3ojMF7j
x5Voj69TVNb+/b1886LHLB7UG5BnGC5n2g5Psfr21aFS4plaEASnzH86d8oukiVUlYp/yKzpsxUX
Fj+Kz0YSMW8/fcTbnatQqXBU2mRssoPPb+Z/TrCRrATdox/MRBN9Hqr+xVIYoGGp4Pe437aqcldJ
DfaJ0VzaKLtMHnOV+5JTc+fUgz2SVSUcb11zLE36PYZoQpUE1InZKzFQJ0UE71ibLnHaHQSvcP64
1W86i0s8NjtH7z1QK9/08Vk8UCP86vGbvE/dJDLWL2qBioHdhSXARaXfkS0TWS8UBxF8637UsMoA
62IyYMxsbvqEeX3va2KQdT8iZWAvDP6KTThHrHegh/eCYg3+AMaw+h2kj3DVOGyiIczvWJYsQBxI
oh7V0Xrd1dpp/UiaKxHZ3krUz9jHuHA57484YER7u3GLl9seFkzqsLQ2AIVZ5dyryP94jLtm2O2c
XWyxCfzxG6PLJdB/BBEHhCfnPBqQSmLYzsRmHglgqs9aHmkWC3MVP6Wim+36qMVtFJiTJA6oLx5o
PaQLsllPF4Mr4lPq8jI1+Sy/TmurYPZtebPRD5XClIGloypUrYWK2b/a+BXK7nZs/mf6+ewz3ap1
2vJeCAwxSROIQFUNZI0gnEttZmWFUX9bHtrY1r0pX60yZ6iMBl0xxbATi9IJJtaaLveLFjdrC0jy
kBH1nb2t+LjkFt1oqP2Uw3EkCkpK8oKvwo9qiw3up/CX5SyUmG+IzIi0vO3rrOTf+rjg04YOPJxC
QWrmWymMnVsW6ix3XrDKliku1bsKYFyjQXTVD3XfHwvjplzkSGi2g502KzjzO/hForzB3s6ZLX8N
aFwEHVmDtRHikPVFK1b/xSAAuMoFgvtAuw8OpRqb953TzLHmlaRlWc7shRQLnnWC3CoR5v3ygkb7
F8XVLWvdMr6889oiT10qvmdc/I8ZXxR3HC8c5quqLeobCtT8qJ5Kuka2QhBlf/8jIux454R9oXhr
0PX53r9f9/FotxAPuEIezTAu4cSMMxycW3s5aCm8BWgWTRWRkjYqqz0NO2TeuGEQaltrTT1woSxQ
3l7XI8ZJaB+QLjI1BquXskmx5v2vglqHhc1wPK2x4wfTsfeMZbjdFRKmNWjb/5IezRQax0XagaUp
y+sA80jB5/X2uj7BeGLNRHknoEFTI1NyUtODFhaVWCbP1FUjln9tmoLXMsu38ErmbawPjncuZzCJ
aRbuFkd7pDCCxJdiXFKZn4Ohbkg2dgWwyzqEuNDHoMApyboprST+A6oBP8RRae9Icd9hKdNFmcpc
3Jtwn+OazALEBbSARmdj6IpqqFYgnGhvzG4cLMLSIqieyBpWGYXQ0mL6hI9Qk5wNGExubUTfIeRd
Cz3AJfRqGTd3FkimMwHq/G6k7U7FoIjF78xLKhJs3LvTkDqrnIUwhwufLthkQMyx0qUJ4phTq0la
mJ+k0fqy5hoylOo2cADN5OuhtJk2HgKW9VT0pKrqSeSZwmdTsk7zLuN3NePMuyxRieBxZFdTFSg1
YnuTWd0L1rHbgbD+sqaej6Tnpvr3yIEueWA7ElIuJKV1X4dgFWe5eH8twniKHMe8pnOE60fdqasZ
NlVSIbnLVR2FJ9fNZgttPiRMRF5VNPyCtxIdsZrEtNJZ2LHbYsGjeZJvTsdtR1U1ZKXTsyY4wBLq
U1887H5jw8PZMn9bs19zjEeO9fzNVQTZaLmRbLMjQnqeR4X64DnkqokV4n2UklNJALlL8hitDwmk
gYcuwE3o5SS/CwR00RbqctP6YGUYT50NtdPPfSS5IFN3Dn2y8BOSbjpENaISgr+VbwAzftLqBd6r
44k9z6nVDDsRiXp7NS/cUrrUlaldQty5E52uvRhCXdaZ9VVCPzE1dxSis77T2YwiU7kqkJQR87JW
Dy4UEN5ceYs1IjdVccjmIDcRN8n4wLYsBsXm4YNQs7FlsooEOxY7i/25/VmKKTfvq8UpqUz27MnK
ux59TBvumyFnO16PfB4SqPbNJ2KJWZUbbFp24DbWx2cOkQelafElilymI0+eVXCkqVxfx6moTGnA
6gJxMgiX0DxKUy4UrtyDOm/uIT4Q/og5Dl5ixZHynlCszmkmOlBcCXAeqGc8e6Y72dxUNpjnMzmO
IpdtSzAAujytfwqIBGO2yh73no1YP5OMhR4kKpJCPGhBLGC+DQmMn9WiP3tJV1aaFI3JEL/ClfY/
4TvomidSQrBQZS/mMuv9KTy4aA+iN6/sJiJpZ/ih9/VJeluOPxZnTB8NopfL6iGPQDGkJ0Gu0F5y
f8DlvBTNCSatKTu9a0GF08Q3SG1+y5Vzv/LNWxT5syZh1iGBbHqtZviMIUDHczOidOcL8xflkHv+
Rfzvdi3qXbraPfogri93xCRErPlc0nxK6wdsH+gZYf5Uujny27iPd0RyqlYhYWYxbO1KOOa28XA7
nvoNoZ0Lx3GCGUQaDo/dvzqgf+Rwl5voK3eL6v/KaqQnIJmSsa5n37RDfiea/Oq0LiGF0DVWWJdb
qWYTpx1nOVXqF1n5kr4HeFAo7Jogsf2qsdUaE/a1J9ZdtZXFKqtObBPCLrPC0hGmDj8XyBzZ6eN5
WWUGnd+BH1QsV1yTpfxOAngy9s4RdxmvotMTQ2MIG/anb5WtawacReAaRJwzNflAdMtvodjCbcfk
v2HGP0XbqP5Y8kRfPKbh9N4OWTbCI1tk5pnnFV5+PDBx4rTpkYw6qk2QcfS8Gx+zBj8wL9M12NCK
8Dazezio3b08NG9KHKth43rNruTWCb4Gdpz4afs4bDIgsuqKv1koq5WIuNxgyLVbUVXIARSy39l8
qTLSKwtPMydgPtprSTf7Jb/7GKq1ajEmanxuFdaolUyxhGXyqZLU40puoK9nNq6hcxUY8Wic8uvd
CR5HNp7aRDFpQyGF0pJumt9s1sodXI0kMr5GG/o22GiArqZ2He47bA9n4I1StqUtZtod3LlTQsIR
afHgGCW7pryi//nMcBQIvxF/3KQqkdzUj7wUg9KLuUjFmwKkZSuLATG16eKYvctWtebFN2D1mf67
Y8TAKJscTBW0EY6mnxzOcbpH47IaoZnLrVpn9Krbp4aOQ+Wb+2ymnhFOnzIAqX4InLbxmCWtspjE
p5hKB/RcWKIg//M4rp+fU7H9/151CS7uWsFwjK35UrftDd7c9nvoquyZyqZoMn4rUDpu5Tv354rJ
r5Qur/+BcbtWd/ec/rcpqJHGCrSYXV9NCFGGgzhJgpBu12LRILCIhgTpdOopsEX1Mm7/2i8lBjN6
ibNODJG5u2D8gySOm3Xcl+xuEzOUjaR9UXsqCfF8akWU+JP5L31/PR7Bi+2f2283zjPSlHWDlSeS
6pv1FDRPPeLXSOaB6HVv8Ud8ZKa8DAUZYG6G9Y5JZydQeD5buMHs02hRlOlGAwj50WrPU2j2k0ms
CL3z7XYnbJ2eYvhYoC5EGDa6Ydavu1FKgoJ8F4k+aB/hBQWN1oMOB85oz20GXT13svQwmWIwEeyg
ph3eAH1DDXnBfKRE/pnI/sZzVkenjBF+1zI7J9pm6aAehSV/mEBwJiJgm2FULrY9B/uwPliii9xZ
a1Ro5wzrgvVsfi48Rl+syMGN2o2Te4HyZaNY9YFz1g+nkADfRzdwdguA7bJxfLeLfShjDuvEmZHc
53/T9AOtRm6WURQT6lqnc/QNj37i6cBOZe4rn4yXB0/T8dw+B8KyonUESS+Kr3e7SlfrmcVOiist
tSMt12UWnXmxnC3h9AdVufaktRRkOA2bYFy7hva27J4sEsIlZbV7qHg+Tpwm1mijTGtziWm2wRfB
Lora5vNNVu6+aqBlDiTvK9mPSIBofAb+RW8hUIPXty8PmlvLD6v9di2p9hx0+CTTlRbpliWtPqTl
0qb2bvW/Kd01bM45oF1+JtNKZ5NPlhHNZvL374+eEeI2/F2a9/wYzm8mRcDispIt5G2i4Qi1poJx
sp7bN391Jk9oEijQygyJdjTRnjDSe0CiZhUjtSbEF3huXS9HpRX4cB0QSLbIQKYBvtgVB4TL/5Lx
zZL9qDc4isjdm4ZxHqb8QnHHEuxjxFsOAyJTAlwyQ85n38KwG6wp2aKF/u8MnBF6IbOByKFB7sFn
nt+o61GGX3maAsyADjbr+w7lw3WorQznOUW5xvTn54a5AbmlHVdObhCyAR4O/6MKHb52EaCP25bN
IqFyluDFZhqFVMOT58xzGqX9ahwJuyKL8EyOvEFj/mXo9lLVc8OY4i8eZMpnrPihn9TCdEY3oWxp
b+aiiylnbUklN3y7+5y+mwdtUUGtiCdclBa3cYFGpaHFihsjxVCyVaZ368U4vWvkQq0wAJpFC30M
NFkSKLUP1er/Wzoh+JobWBZdPvLMosLuQTllR9Z1TWeqCiMRLjUYFDbqngbeGghY8KXsZ1whMo55
n4ViCaE0hhOn8ME0qt8A8xVUtUypWapZDIoa7NFLdBCBl1OBxDWN0FW4yPnbQq1fxwaQxpOT7juS
pyFTb7rMERBb6dYEMEBjhjgitCtleYNoTw01L3C4c0Vqm2pGK3N4bPuDHO0zz31FM4jndg0yeXQq
HwLqRqy1AzfvDw4K2OmTAoptLsqohPU9sHuD3PsHDIwkUawqgk1ENGHz+VAaiJ7bQyzJG+g9b9X4
GLbMCO083nhblso3KDc9uQs7TzqWAPMU1Ynjl2WrYqufie7YZ2YhTV/yi8XiEHA/DaxCdf5lU2bg
q+GMn/24HNdZfGy/zCM6NSuBxj/nobexnBzPKVm+Ol/fXjdz/nD4sc4jGeMfrDNf4RZho8Ysunrt
fgDwB3Zc8nMCuEoiO4ABbqk6wXNWMAI80qNxZ9on9EPCzSaXTuaZageCygO+kk7mMA8Z4oqUhPhx
90gMyrq/vbZyD4aIipfy86Pi3KnKuGTyaty0W1A1R7KszRsLJMC3gcOb0RAULpVYeRzExvkIzwEI
El/B775KKAuF1olMoo13Nh2T0O2DGSP+OgGIBH+4FF4oFPDskxQwfMjyRGavg8JfTrrLykciqYB5
lXyuAhUsIMWHsqYMbjhcmXDH/dsHwiOYUBxcVCwkodNwBTU8eagGLKHGmElxgr+ig57zrVYPw/jf
Zaq+XdooBh6KVCQRzlHM3SHQc+BMa7oVy6NQitUGmnPKHGqhyN2uKUM/9UDDkibdlrSv4dpzkeQx
ZCdvAifPVet/oxdMafbSzM44qFbGk7KVBf7w9nhkcu5N/BszdhnUXWxnbol/lmOTGQllent+souL
rHlNiQI1Lee+rtxuJPNS3r5UqS8Zu4USKgqCBeuaGEbp5krdE+gBdmreFIbn3daMCI3tFmCRx8dA
ENA+8fBGNpB1CJZaMWVidkIdtmAeiPs2pg4bxDW3GoVfLdN/8Mll2d+rEDzAEFJx8UJMf/picyhy
7qXGcVS+P3gvCb26fO2xG/toOKCHq05JyKwnUkSdigIwHbr5mwcH9GG4dmnBaIGffOGddlV0bzJ+
1GEqbpxWzROrjDOTi+ydWAiUYvmg3KGRszcLgOZh7mAv95HyceKc0Zu8nMJSaMBMCq+MmeVO5RNm
+E+0w+6ulkgzPOjRE86fmVeDX+Ac080MIrPp84DR6VGfKwbdSAx+K48SiUNhf2IplhiJl9ulIY4l
Pf6YCL9kCq+DPHttJDkhAB94FcWopx+SogDe9wYy0cRKKCT2QRnZMlgWyEod5i/7UMXMl/6AoZYA
UkIMjn4h/8uBEogEraEp76BI+QDLw450dHSY7GTD70rS042t4WuHxuRSaCsWoIeEe2pU6ssylozU
uPnODTOI9Tv5qS4PpnzhrQkhojkTvpqv5LRMIEF+WHe76pEZAS376mLz7UhkUtxi6fdvutmfapxR
X+ku2v4amkoDZ9SVsUd7BK7AT5HwssvyTiSibN5Bf5oQHsor2vlN5wjZxiSxamTM6Vnh0/Ai/hBO
XSkxvqSPsGbho+/XflXPXDVTfFNg4TwCEgwWvgf9FrAxPvPquZ3MQTJoqvlHmzItOxrcCiic5Boy
eO1AS6ao9VTabt6zXktbS8SOKhl6+hV8vHZv+1gmmo6k2RkzFeHg0OmHlG+qBhNWbXQxq1omrlw1
l08cSbBcGphfHU5qGNOldA+sjzKZcf3K7yxB5pSVbPLa71KGF3ed/5pv7o3EjTyLBjXBE15Hjpz0
+oHmc7rbsGy716zkStnhhpU9IgpJssvlstuF4K6Gx7IMHhW7bUEnFPO6gTw0QZ8mpbKRKCojr28c
siu6zS/3BcvEXZIffq67pKkzFGLfj3dNb4odgp/vk7IyEX9oeDkRAxjRr9uZrRaMkM1JPiVtxSEs
JRbNUflmH7Edk1J4qo8tccy4tXgu5StUI/jpXkXhfL8RQMkyT6/z4RCPlNpxBbPMSXrtCwGxDY35
Ic6SNp8m+FGJaGpZ1Pylk+XnyeQUYh9sQJx5C2P7CkEknsm2oelr2sRL7oiTed6VmjNIZYSZkLGd
ZIbzh+f0Aw/72c7ZzsEF4rx5dBoS97Xzwpx5v7RXWMDMTocZpP79qR/kJKbRLOLgpyA+KM2IZ6KE
D4UyqUp8YtGIiQoxF00q4orjDckdp0dpzG2ZCNH4wB9eoWSHTCfuZeHnfGU223WnWB+ntzJSmlyI
vdoEPCap5QROQcSjh7lZLKOlHuu8Wncw4ukTV3zHfyh6aocdqOzeJA0x69w+UCuUX30QYTQhaBlW
Mkreaw3N29Ua8jnXARzzjB8Q+BXqgXiOwNrD0cewirAA+9EanBtFuHnhxYduK1Tys2fjQBKNeea/
GGHAO+Wezq1O0c/n80lskNO8hrcfC5Wt52LZuC/dUuLUN1cEvbZI/9iwC63eFeyEt55aYDXreSfx
j/jcv/bwrzUxeHKKB91fNVUfgXNVag7bcDPq8rOGDhCJRzCyYNunH+WqACEeEldazUJz7oWz1fXZ
m93lkAJX/p1UnapSFohO6sxAtnqTjtgGlalRTP/n8wLKxQDE+SfDyzpVpejzg+Hs6JlNbK9vjL98
dT9kCdZgVRTdLHCx7/9m4uzHxGYP/9Wn6G8V1IfIc4Lqa9SYkNRZ80LUSnZTrh/HqK+BZKabrG1C
SfhCCZZrg5HK2B9VH9wqX2M8UysjeTHCRnWVXygx6taZwU8pFRjDWRJSA30gs+WxpGuYdoxwFjpz
67910OYHczV7lDYLAk08X5Zd/KHPqsbf/0zUS2RF+omQ5apUTT2M0M06XAgUtF8w60KTrX8x9KbQ
YlgTbv6Dw2sNUnoWJ7DSKzSfjskW3uyaK/25qz72dHrn7b7ZKVw/ohE6foNQyYh0JGRT10itSXkF
CdqJfxuKu6Z1iiKXj0tjIOFjoIc8aCwwvkcF6FQqbSEPxH821ZqZyINqlbTNm/HlFilhzaJWf9tt
MHtpaPe8shfXP6i1S0kLMIPgl5a44E8IsC0GC6C0xc2qLkcCoVhH/jg+bURu0zchSx7FvALbG1bi
J05++YohdUqwqpBmvi4FPEZCiuB554jky07931EthegVD18CgS+ocnF56c6GlsEJD/0PuZO/sIiD
TWFkkY/G6irMW5JME44E7Tb7ZGSE9N7cgDAtcV7djCGmNg7hvtuy9x53VQXvcRe7impVVbVTyPmF
KFSptY/ZMYR2G1eGTtgW20O8mv80WllAB86CZQqYI8JChAUIgte76lWknTgQBuOASg/9Ml9C9Sgd
DOaY1MR5iuGwwyJOGMTk3OFwvqqwGVf5BiO68NGpt07899mWhZLhLVQxeQfcUdgrEb0eypZ+4cKG
yXgwN1rftyvi2hi4AEDYYNUZh2BO0XzG7yMI87kqiRh2Er26C01E/KJEVN0n1I6f99mJ61QaDBu3
bejLEFTNcTobmBnnxwuTUogYJ1nm+8J218KGs4Mz2fLTE852XpaLvaJWyEUN72V1J/ZjnKADXE8T
lllR5roppDQJgA7D8s8oFlj2mAkS99XR7EWOuaYWpB2T25ASBtIqA7Rftcw1qq09OuN9fgz2cl6C
nZjj2En3eaLlk0qd6SqJa1F64MhhD7ThU03D6Vr38CsVrYfpw3RTnBh/kxTidRNOPz9Byo8IAKaJ
mbipRWeeKN68ckxR+H5RtdMYEAIo0AAEX9SRvvltRpZE3N41wxX2FZ89IGgeA+a0mgHZlGXFh/lx
FbgSH/A188KV8sYBcjCcD4MrFTNgAsVt/F/95WzfyBqkxoRiFgxX07jglkrIrMQNSHmlWvzM9BCj
qPrCD3AhMPyiCOWBSDC/dEdq24KlyoKuL8YzkebaX11m+Ng57aC3fnQCnwN3rLeMxGMsWcWMYwX0
qMGwfRbwa8yNNjVgbDMTV97tJGkj9mlpPHjJhzVI5x7HBBFilFo4kxGc/bH4pZv8Y8pN4DisAGCb
yuVoF15WnjlN11WpfdFo2u0k2Iik9Pol/U4LpSYIADaBslXyS6oEfcsuXyXuwCvRTNE5cFNDuJk0
rwi49qX7l4fE/ohab7b/Y8fCLeyTxhmrhMl7Hhc3A+N/K4iXkj8+vxuVzPP8yRsEvwPvGDWQdo4r
G9jh4Ew96s0uO5Itw6yiW2eKOVH6nCazDvRL+dK2YUrlLM5v1B4fm2NW5SysMVNujQV48ZwNjURi
YfRmLJzSIWayetsHuO5190AWMr4Vi/dNoxwIu8iWCPhEUEqi+7ZswCQ9bNOo+4cFUPkBjlGHhLXY
rq6TMzbFBtWztO3HaqG/fcsjI5T+bnrNBNk8qo3WHyRfaXN9bnvZHM0OncoR/nLAgPKUk+rKZUYH
HU8gfKc2X2GqUH99+Yrvj2dZW5V0jyuMDuMBpZT+c/3orrshGkpkqaunz9HToE7F8hcw1uZPW5u3
vHJ+jImD3ZMmmQNgVTFJRVeDVtpIF6OXUKrpInTFYbhiOw6sda0lN2+KCDi8CrkpDLwp4cvGFRJ6
N+y4uqmUHkDh10vvZLv7YzQsYlUAnE3rEfdyGMQXWxj5DJB00sIOe5drgCTUzUtL5G9SnTC7jsKw
anbI76sfoDO8nx9EhFfx8St5a5/YPY2ZpYUslZTKDLEzqxy73R0Q0FJpMVGn67jjN7mfRHoxQHBQ
8+y7XFxQQQEBXPdYcWDCKciHuHo8TcLJtvGcp+HA5h3dunCN3YoeWN4btSp/wNPgioSb31ZMCjrm
4a8kL8S1wkw5sWXztb/Rrwr8TPdo7BCfmJeTopAflWVPtccRILay4O25e5sKEpNe4XrQwza88keU
Ko8/bG46l4D/y0bDkEYLBGs3pTDb9516ePwneihzKtd+loQ857FWZGEpfEkPtQ13YyHMvpuP3KBt
MSGkD4Nr4W1hge69FMHlVeY+0nh2A/5vw5Sa713TKgxCHL95kfGZrFvSbftyc25c4URYKJaw3qoD
jyDVPomY0ZgVih6GsoECAqEjN71q8F820V1Wv14d7f2R7Qel3gjgzkLahhqPAgWkOOWf70WsGcnt
MDWzOZgpytpzLSO2ecQ/oPu20d5ClPJocjbssg6o2cBqbk9cXXk/J7i5JTcfY0egG/dQpqiN/8OM
VUWV1pnYplQcMumJIDVlaf1KlUhm55rnMtO27FuwmYRQOxLwhVGb/Dk/lrTt60W7rbQD8OEqarbX
g7XMAvrS7G8jk6F1+9z+tRRXEEwO9yUtxDmMqaf2ns7v3TkeycmHzWUqmdfDjOzYrgOpMs84cKM/
WwHQuQ55juYFp944JwZvDaVlkLAf/r6qqPCJbl3yFB9rBrHQisBChsRx7G+gAFNJALsapq+AOFzo
xqxV8XAHII+xqZEpb3NAs8uKXqcnLcryAas2fWrsCQH77DO3oYXEc7JfdEYxEIO5NRm94+m5VmBD
bRy1jwgk1K6ODyh6XwezXK49LwEQqD0K6ashda+rm9+khoXqNqfsPMo0MQP2z5VajL85NMK1T7+o
hzWMHzMvG9JeZTzUx5SkXJOBslwTN+EcjM8lj+UXe3uKR0StzwWKwQ+Ro2qyBvb1Q69NJ3lbTiRH
3UMzu3GLjQNHKgKGFZkQDALzNq5YxquB62TYrN2pULIuU2RijDQigFpA28oxtzYxev1H7zzUmxSW
8yT5D7KSmyF4SUDRq6pY/0M3rDhKWn1I79cFUPmvhWeoMkzUBmtOovuqxKbwqcURqU8QAtUxQ+TP
179HOn73gGYJQ+Edlivnv5Xqc+ja1bFSe/R5XqYJcku8YDc/o1hh99ZjrP5Wr/p/b0x3TCgGO9L0
sS6rPz0lHMcTrEAlNn6fynQCXBP0SJuFEMy+9i6+7xgS6/aOTmbzriUBeVCLCQEkXvv6+wmd7YWG
+S64EnAJ5kDvUz5/wzhL2UH34oaTXQvpQyflLOA9Oh9uDEioVK2/zg9TxTtl/ANS2SkPhGIBXow2
hymq+0d+Xww1o/2k0OpYYAFcUdYH5GZtTuDLeg8LlIAMHlwt90NL6Zb0XGoTB7W1p+VR/JtoxOpN
gtw7j3v05QmasG2XxEXwzrpbmG7mbFVCIuNZ3i2rh/iYJaStXdExX90cZTRJqCbhOfPEG0ebw3Dd
gGVQ0NVk/aFxuFhXepUdYMVgmEEBTCK0KUl79Hda9VKRfqU4bxNmMWP7AlrD11TYxE6mWCBr41QE
jINYOTX48xCsWzNuRTTxshgF/qrve8rKUVb9PjAOXhwghfqPyKXMb2HTeP+1EGCEzZgHKW1zjc11
Oy9T2RHATgW/HUqe6rtKs+7wicDvYC3bXv09SAY7QVpwtd3Ei766dUxnSkhMJEul42SI62z/vPY4
gQiqb/4qVBm1Su3ck+TRhQu1P0MxBAXnZssYo9dhsjLM0d+UfBZmQ4/TqhiQEKPAk4qqnxUTGI+G
a1AOXvvtHps04vLwfavpnstfD7V7FxJqg7OJpTUbwVxSE+DYgaqHw/GuKPmpRU/Pz+XU+lXMJXh+
By9t4AUTWizrYHuU2Zwem0Bie6bRZXol2svqupmL5AKYpxywcl6jJ7GhK/dZZNPUm3FpOvoTX6NK
e385nEGVBudUkUXDXoPi4MwJzj0hv25vCgkSMMWRq5DILdJZbRxbkTA01FoYWuY78VCpMOiymPmJ
OsO+qL64IzmO/hFfXvfqVFSz/zBwCti5kRoCA9eRrOwZANFwxLHIql1W0nl9UUHRVVymf1Bve+J+
hNqoU2ihzmfG5DcHXq3IWI8bZHj1H/pwnK44OzmQZTqfFRm/3nYsIh2kJ2Yg3A/YYWjded7UNoDJ
7S1GTz5S/aEQm8R+IKCoinG4TkO+WwYQt3MAyn82XStGszKnKQlBhAyUF+Lc1a99huGaLU1ssPRB
G1OZoCha/OSK5VwjkuYslxrIBH+QOsm8x2nRz9WUCLJB75HtAYyMBugmA+9e1TS0taKOrMOjsBvO
ANXU1UDAs8Ue7pPFZr+5jrtuGNvQ6V04uvSZqLlHNV/wvmDP5dXwGSNs0xlJnvnpEH5xcbBCq31t
6wCeOKv+2th/6Z7DiFjcZPZ0mDGPDcSn6Vi1fmmOq22jACGXru8j7QcrtFBL0F+adQ4MIcEz+Off
Hd73K1DS9tLWwltwyz6AWnjRfmBrXu1wHQTsdg+m221dHHkNDBV322Q0MdeII2SO0kpM81c4+JlV
bBSYKmSkcM92yw0WWIcrxB1FIzW7tZQZQXJH7ZqG7NYvf660KM6CYvIyDqQ5enxD+l4dYB8/z8Mv
ACWr9bFIcuCKsFUxDq4p8nNSY6Lz6rrohMu7EYleDOCOqEhFxA08AZYejgreRfOKk+cVyLzsd/PY
NzlXFo8DQaZN34q0sMyRAsT+qs63T17yNNs58V9CjYZn7v+RbDQffWxZQPxvpy8BMxe53wAQcRL5
tCm7bWo+lfmGFKAL2HhnZn1KG4+do3Hr01Fxu0oAx1iMuzhwsZlQ7LRFLxHB76KHzmyXpo02ZwIM
3zTaKlUzbuTAHNJjtesAzwgnh19azc73/dHIa03ssoEp48rF3CVom0FCM7kSWdLdLSqTMGTVxA0U
+XSiYyRGVtfasmkCN6vLCgC8hDj3opyysZ+iYtOsaL95asdXRALA6Y2VvRmlx76282oo7Mh6SQGh
m+KGp/7bA3NZncQCV5I2X0+Cum2povRY+b4n8/8RPGmnAQ9aKpg0IkhkWHbeHDMHxZbAgzOinHK6
XBN0Cffi4OtRYMy/9Zu5Qao8AEddHpAV10f0+uImlsvtscK/K5QYYnB1r18oaVxpLp97I4nMB4T5
O91BxGJQIT57rZmdqCopXX/TRyDQ0aIhlrx0Yr5sBGt2/QQHREn8Pb1YyqpNwt0YjAv9TJytam1i
fLMI4MWtrlKElGhTFgz4ETvnwTbN6ben/ts6wZCPs4OIl3t/tOiIvSQGJPNyjR7D+nLch/lVeNWD
v6mLIQzx69V/wy9aXi+MPGCKwHnHQixK2TqrXMkAOTGICr7Dza1h22O/Zd5o+NvzIRfbzTvUCvhY
JgDEfFENvfhOZEmbXt3UAYw5vBryWBcGWm6kMoiIwzjQb4KgO3J0p2BiMWleKvWOE6GCD8cCVTiO
SCFKjXeWmw5dmE9LsNQ4btMAuZowEwu4NmzVeQ4No8j9yi+yuODOiLDwtHSs0tJ+m9UaHsZ/kQgZ
/rAs5u/+SuS/cXseSQYeuRuYH67iGb2xOfyDxYj+fujOP4XmR0Yl9TgDB/lK1CMpdtb9Kosi1Rsk
CnojHu9XRH1r/SF+IpP7j5icAmaVcu4OrMbC6K8cDXQ3Ltpq/wflysLzL9as93HRmKBJ1SSlcP5e
AzFSP+fW5uJVSeOB5qn8k3d0MmWN17fEmiQxoWNZzmN0Ve/y/wUI//rFqcxj0fHtJrdA790nDG8m
qvgp/4eifdRArl8P1jVhmX0HokpJn9/871grzfInKCvFN7ETKsKbrY4S5r9DUDKndyPYx6WSwN6I
/rdBpF9G6RgaS2F0BLzxGydVJ5fQ5rbA+qk1tSV0tsxfCU0P41h1wRvAWq1yUdURTOcV/4HhK5v2
8F1dTWtMVzH1LdletRbuiMyNtGyxqD9o0FGKNeYnbhM5WIZ7qI3U6mraYuTjHqVMt7LkbILl5E1F
XLgr/Lpv0VhYLPz4T5BhLiNjqM7KMDaTJnCbPef+dnyjvE1JTIMv4j+6a91XD9LM8qaSU0Z/f6mo
M0JkV/cnLLBTWN+ks5Ct4OA08wONyJ2ReSZJN3gJciKHz2abT480lmrdDDkLeoO/7+Cyizhyq4Lt
aEOEqXoXdLVcajdXnfrt2UEGOIQxMLg5xov8MUaKdw7fbUhb7ed4brabM33kiNVSm10+hqW4JlEm
kNkOszIK0hwAp8T4bmLIcynqwbEBGvP99Xuxpqpesj/g8bu65DMRxO7YK8I299iHPTGOvFQsQqOO
Mb3Ibrj4dO3VyT1/8Trx2zzZr2mQi0P/hQEnEXxy3jxxPk7gRJlFJGisc4D6mJa+xvGv7hzVIryZ
c4x+mMd5iQIciVF6XmN+jjXY2LcI+gDRqQf0vfJG71lQNRpuaCqsEKdBXu47jdhuK7AHq6vmjA8P
qJ61FF6acKRY6fTQvAaGrUuzU6DiC8cTqPDUmsEm1pf5uWqsWfD7+IaKgxTb7BPv7tQHvCvbWOvW
QHpLPUy/ZZ/C6K6vYOCk/CChOvGCmzmg+ovwfwAXyEIxxXbjuDXEwKhFnURfq3x225n86ENDM5BL
WW7n6XaAgSGdzir9dfBaxOq9KkUpE/0R6NTudtaqPgwDIfW+wwHtNtGYVgNwwka+SDMEPxoeIopk
7vLBcOkLPL6vZYPuNhE/swC2y4h1u6+QGQCuGQn7R1finLs6JSKqoOGZh/N36uviFOax+ClxrCgv
Oa9yDKBjcpvd/xb1/0B3OK0I5fnQasJDldwYQDNcMsA7+Zgx3V1iAvSc3ziatDHw16eg5SDJyS3M
XpN2+ThW/NJH9P+FC/9IzKVTa+id7RHKffNErlmiFgIOcsNSZjVo+83eZnHdlac1nh2hJTheEANU
zgK+73lG+nwYN1ToM95iRuEdKO6dLMOf7CJNRCyqYzHqbOMkWsy32ud10+LXhxi7bXnJiCmlHUAK
aRXlZXJtMN4GZPwpiqQTBBBWtYwtyeX2HdFUFSkOVMImYqKV4xmYGioaBsQ8/5clZAxvSI4hNL+E
GDYgylK+Vxm8corjLirWY/1I1sHlBg/r8p2PtqVBbC3bWgcrHt6Mxcsdr+L/BFS6nY9aI0kF5SHn
UtjYUC5Mt1HlLzHayZyjOxK6IE4/KST0f5f19yu7dTHPrzkNcStcJtYoxxNSk5yiDGBNBWKlhIp1
nBGRMtf+bXwC/dYJP5CiGXpsBzqF7x+NfKklJc7YL/u9dqxwo+JEdOsNxWm/1dCxROxotRTJp7M9
63Nb5OxTdJizMpegYfyeuJZKDyQp6EYTCqqV9hLW9Z4fPSX9aiQh5nN5w9OKLhMjTMl63zvj/N3H
7xWbrrOabeGeQZbl6TvrY+7N5YCNBXM42xmTNuq2U3u2wFSeEq/Y4Vu3+HELwB7EVr0yHGwEYwed
D3pgdkcYcx4Mt4VI4t14kKDjh90+0fSqTpTaXbks2jBaWEwLYoKffAQEKG+yCkA2Ulb7aNJSFQ0d
I7DFdt5zFLS7x0Y9YQLUKRxU1h5AXMmXB18y81PnL2l5pWW1tY+itVOmuTR7okJtQK6tjuEL2SqU
TfG7yZCLY9Z9GjLER9EzT+MY0BRQRCo0BgjWYGcdrYWKfm6FE5b2Lw/agJplWnZobwliKBtz8yLN
C1BhqFy883Yx8Tms06GBP5lWPV7nJ5+vyUfjG2PEHjbBeZo+LIfAxTDpDA625EoQytrfqS2J7VuL
kG1gNV4HV+hfZf8vCJZz6zZCRqyl8s94AW6cIgKqZmPnoYmJtsMz/aJTLrKfps52+pZPVxSjJcjp
aGSzIbtItcVK4YX/JUSWVWDQTZvPDUfr6KSInTAhwCYmPRFdjMc5SsQiZFRnJiDUpRyL8LlYW6BC
5pVZuxZ9zyzb0b9J8Ai/oKn04u6Bfe0XGxsMOVZF0PdelXkh0dEfwvxMMY7tQVHB9I4mUb6bf+Kn
gWHvoxzu2EzwkCj0at3KqhgbtI0njlPXXbkIsEdLeAxMc5F8HeaQlbxPmhMSIIvBw+VpAu/qzNrJ
nmSMyR0DjBADUy++YZIJtk0JosEtka6mi3Clt8FmAuWi8fRwKmvGRxfRnTZ12TO2Heu08wxCGwZ4
qKJkz8HeRXAaY4TkLnzYlCt7ykYb+O6OIIavsJ6LIm7jpA9y84EJaEvwRv2I1M3vgdksqeG41Yxs
T+VaOw0cdP2/zUpXgyLAA7NOx45t5SWfNZyXhD6B8OCP3dO2pRFL7oYeo9pDC+2XBU0Tepg+al5M
7xm5/rmuublkQYV3R50JoZkLRyNY8pZ5VwelF4RAiqiUl7WGomDts6ooNpx3dtkQ0LbQrccwbAfI
lF3QdmZ4TT8uS7ewgkZUYrqAxaA0r+p5cXAmCrye/AwmGiMn6CKpFkbxAIDSzAW6rC1Dfs/okB73
MwQjJ36L3Q8TiXn84SZxH+MrEKokp/xitvQBBzIXzPaXNY0Fpw6ZrbEOcapSY/DYtoYoMVy04OVx
yc2zrdu4Dh4ynyDLUsnCJz0uzsli2XlF1PSUSx7c2K19GSrnwbznjwKLyLFA/niTlwiqaWAIhpfu
LvgSMd0kkFQPnhfoFz9yqeGDBzMIcu488So3i3z0XG1mxbQAQDVdVT87B32x6Y2XwwAhqZCrc5Z7
ICcBMO9Ianx9tn7lf3LSnoCIHQc8XA+1cZEBTHcVvfGO+ysv5JAty++EDmipAZwNr5DKEFULf0V5
xN/ie1zZCHZ+/hHNYOh4RZJU+bTT2EGVlhJ2MxncIGP1IdSICSAPmWqUUh+gfwBI4fDxwbr8/Kw3
dnY2HZnFyZBBvns8iRkBLkxxQldUyxdmQOngyG4trgOJoLbt5IgVX7nTnB5pKJTKYlH5toG+nIEG
hlb50rfSQS0JUt3hVkat0zp+gOFcfvKQZmiraLzK8DHnSx/Yh97eBUA8JKeqqWOEI+ZIjqFWe2Pt
faV5gdTygBW1OVqmHOVp2a8BAO1FlT8GWMeIz3D+PeI6/590RtpGdXnKbG2j9ipKXZ0EuXAwt6pw
nBkUcrwYU9hag9kRPUp2pxnWv2zLvk9C2zRqnIBD51agZ2DtXhEiwOdzUptMOFDbWZufS5e8lso4
UnsbMehnCnJSnqHWWY8H6Qq1rZX9m3rBRhzcNs7nVHMlaWDvMOsJY8PAil4OBk1IYWcpLOTJIS+d
IMuNNyWJO0lAcTwY+Q1aB5p15gG6dyXwFlTvKo1hDZKAt8yYqSxuqGYHCaNPgXdvnIxpwi9Ihzdm
sEXZtGgsBNZeW696PfUDkAf6LV6GwFbCWuWwAzmrx38upRYC7jBfFdsqB6Qn86IQQcVWbdsGs6d6
4aKUSjkr4pXhJuQu8pXglnRvY8fJ2LKKvZFtacXsmTP4eeIiqjOQcVJwtzPkmVai5zvnmBnPLhRD
2pPxUxvcJ2yYKg6/uFiCAiP4ieuMlRwwxUfqSWuACLM14EAPO0rSWlaqEpOWDDjkcw13xiY9D5jO
2LsQRyt2Wv7ouL208gWaVuzeYE0cN9VUAQeKxUfl9yORT9VsouFEPXiX4fnULflQsgPNlxZFY3el
v/hkZaXGS2F7h9zJiKvdkButpNk/n7AYPu9nT3xGuey75MxIp63eZ6UKAL7e5IuLq8qLd1aB8mdL
/U1TBsftOsKRADgxv60cI9YJN0Hf75AkHT1Czbv1H7/nTEijptwPh0ufEuO7SCPBjSAN1LkPh/OO
iABx6N43gafQu26lOryATxAj83AQNNcxfE1KK//F2XG9rkdIg65uDvJuceScItkfencsDc3EfKRz
XTme6m/5cuEq9Q8Z1dBWSrknqc3jcC8M1h5SNGoaH8M/JYxhw7FOMwHXgzQOAuELtPSrZ83LBL4X
A2t8Wt4SJjMPRFHWtclxwKwz//E1WNQcHK3iSAyHcXYMmcvvnsCj4O4Su4VovjSos4GFi344taQB
mG+1APKtCbNIg81G4QfSFgoJgYtiBN8vrcfFKemaa0aQt0ON121rE+rn9EvVigCGMahcXHL++alH
/xfXApl3qbV9o16IVglgUOA+UB5h30l+fnmrQx4G2Na51VPk5bfNhuFiG1ZKa29gFttqcUYjfwC8
MN9GMf0bHG4+lQqCcDv95pfWsXqziqjev73EZfPd7M1YIWB4N/IBKpJu1dkX3ltTR1VJwDbKN48P
DrLUawDGdqQKL9hUQGEeWd3oUZj/rdEwbu/3Dfdqe4um1f8OBW5B6a2kDqj6YA3FijKhhIEkKPuV
/fgX3eYm8+P+zQ0iihgBqIWkj6xUy5f11USD9gYvyQCI62o7sJjFkCi8SeqKX6bUBJCzVqAnw/1G
NG6r9lL6sIyLs5K9SayxLL6iAMCnN9mkabHc8JK0VhU/2mI1Jr283HtvIjFNqtiCT31ERbD+B5Tb
6ISyYaNkczgevozMvNy1005l6vXB0cTzzMBY9vsct2aHN6g1NC7IbBj+uJPoSpw3GcgqXU2lqTGR
qkBXPYGlshZ5QW9p48PcyM1/mSbvmg3REH+IUNWyrZHhOqDGIZwv37NOTIBUQQXPKfd2kCBfznOx
G/wkWrZxwipCszFccnewq0UpGzybVQKcfaoBQchD1+wzoIl955H0Cy5iqn8U3Gu2G5R5lkAveDrg
90cwGWMx/XN8dPy6cuGlibPjQE2j7YaO+cmTZcNrNilmijGhrw82QKLHshvGwL0rJGDlEndvcPxH
yUmbMZz6wwWCnlHQ1lQVU7+vvZgefdnC5uh4J8vRj5Cn8MqpJnx5Uk3uVy6j6AlWftJnVQaHjqnX
ea8nVlg9U3hGDpbSPS+Zv3rlopjqDlQDfm8nu0Rj56mMMUjnbyKIP6H3pPgYLxYglsBHxctBYSzz
J/gMJ7HMnaHM+F47xEyaBiygX/utnkNFatqY5NfLjIHdkRvSUkLcHPhjWa+EK74Jb2eKcxTFMGIb
nHitrcNkW7zGPxvdjr71cvxXstKv/7K3bFMV6+6qq5mLzfmxH7OgRnmDedNg1MJROMutR3T935Kh
U3/sJ1p/dKai2arp4U98JibHqdZF6axYB6ewu69DIZzykk+8JJ76R02Sx84MBcKyNapdi1Z0L4es
vVbTHkxXd/Yqo9s9clRvtQlkadm4HzkIEMq3eBSaHt2R0gIp/EUtIMVDsIBayPk0BYn2mOu6Lxb9
nuPOpxwq5qbVh0yoqMiAm13CF2C8k9BP3+G9b2WLhPWqPuYQR2jnpvRNMTSZR9k28MNvPe5cRQC/
UqkxRdhaOMJdTITEAZQa5bC6WWOX4TQcmDJ1WG1SRiWf919RRrooDKArSEVzvKcfyPNeTDXAwDf2
XJMap5M3QFsiIUC13iY7SR4rj6p+F+LmfTPdAkrbj1Tc5LYdJCSfz1NQvK9LTvkOM9KI0aR/Hafb
H1atyovJDDSeur5SYeH+6LylSAjvgKI3ohDy18MBPnNzusCmTFUZbkNd2ewVMWRVN+h10aPifldJ
KXrOTXPOry1KfEThG9xxyt8+SHGUa8djnlZJEsE5QF+KWBKsekUJbw0SyAFHat0cbhnzL3RyW3lw
xjDKYGwBTDFa6uRWbYv77GwBbYAdPCwyz2zbHJbwoSTrB65Q1jvYBYQ8RPV18vfI3BM43/4l5NO7
2naeOn4zO3ZMzzKpePHIgWZZQjd6r7YYvf2LUTkT7IgNN6Y6FNYLAuNC1B95wLaDtq3liezZOtHL
FJIadJ+xcObX5Q18SUfhGV52AdkdSuG3mrRgX0Hj1xtWpcpVvUoiUb+e9lo1mUcK24nPF7GsqGE+
Ar3jEPkGMRQXqUFaRY55hwdFGaJgdEcGR/EGv2zEsWPnic2+J1wA9iXRZyCs9KCoFhyrObBbHGYs
XK+MNHXU5qlxKjjHmaz0ysDjFpVIRnDqAALF73hBC2+Ymmy5HUzwA8DAuucjvG6xUGhhF8xABgUB
J7fQZXTzR+9VnxcTd0ODAsQhPlDah9azcRDj3DQUA68FzR5uh3DV5JsHjysB+87yfHWXZM2ZXaEH
0+6Fa63MoorX6TSl5UJ4g2WRvEbTgFQW/aD2qn2uewIIu3rcOHIiDynZDdgMkUluywh2nlISJePU
pPFFBZd1kiaRwWN8AiFSkoG+Rv3iiA5IwryUjANstvSg8HzJWyQyAa4eh8uGJKp9XQ3Py70IEw4A
Z0sOHb4KY7+BvQEujT4wBRQYnxU+J02APGQXUAiJ1VYdiPmomdqMkdauflvl4WiBSu9OzMws4NLb
rjDHDHsxMiSIMIul2lOXzXqljy4xAzueUI0zIr7h1YxduhteL9YzAP9D5Rg/s9kSptoInRqOpKus
yrIReNS3/5ylscklhMgeNXqBfjwBA6vV3rZOt/SOowZFsk72BHp+ggwi/AxZlYp5tHPr9KVJqOAa
mzCITKf2MkwB0HS9+1NILyAm7AIOq/Tfgq/2TF/Xh3048SgxKpUj7+o7nl0tC0o1x0K5+BR0LwZw
J0Riz39sifPdF2fKR23JR5IjIvV1eqBiDXGsk5uUzchULL+QNOIP4OvtTb8rFA6hDeex1fleMErj
NmnYqRwnaYismI50z9UN87WCSxDHHcHEJAfOQ0RyHXVzxvnxg7IjcApXRQt93tRtQjcTNOF0AbMa
6p3QyMgw6Ylrl8U9WgAEEzC32q6FkS5+iWIlB0jj+tWd9lSJx/uF3pq9x4bmQJ9gAfM8G+gUmRsV
OE3odZHa0p9dG1V5CQlnjp57zmuelRYOYkqk0ugkuO6XwUBPLCsTjgqkplqtpYeFbOY+wd4XdkIg
WEB37DaRU2KY6fOhZC3Dm4v7dt0cUXOwK9OK2+4LsrOHUtzvSc3K54Gkf6oXHD8B9ZXILtQxWbSG
4vurSmAtD7HKA3x/k65XAp/cIswSmLodKSaeBnJhYGzwRqmggnTyWbZ7ZfMTB1AmUIebIaklkwCP
GOW+IUDK/vX8qAudMyUsE3sAFOtr3w14mcjE5DVjNNVwipZBCa1a45VLIyd/M8/fmKGQpq73WtXd
MZTvkMeoANojGeZhVtxP8n40dYMgqx/dRDF3NYTaRLtN+k9qAFRDbdzdwtWCG4vN1db74GiqE3Bj
WST+yGTYfHBJFp9w7gzs4sU5YPrSgh70MdF4C309zS5SnYQ9wRsSTDG4LACo4OcjRzZyN0nbteuS
/mPSoo+fLcAp1Quh2RCP29DW2ywjWM99jePi1OmWKbcfD7RTHT04dy4cmoOGFwM07zkkCygrGezH
jS5v8EYCHf89lxtQjdX5rkq2U2n/jGcvjsdVdFeIvhOJB+iIYG7m2w6H8MjIq8YH+81Z4Nj4/RT7
E2BB6zx/kSQtC5KBSnA7sNI4uOoPxhIeZIDXaOVDPjNQdlKceOI4ue6zn/NqxU1UFKnKAcGeDi8C
2zI6t2IlpzKDvmVaT1qhf1cerysVJWj15IjA0z59utvH7QkPB2V2/FFwKTq7zGqcBJvgpdo/J8Yx
4cHDISf9/z228QNIrIKe6J0UXDSvUPbbnu+Ecrs0ABfncjSX1Vj9BJ6SUuRbOX0YDVLhQs9dzewJ
T/ceX1R5e5FaNjLOmNDWUr5OGwNd/eIF7GEqPabkom8wwwrzmTsQTKZ3gob3lBdMfkZbGKfmkBln
Z2HQOCIU/dHeljon+6d4ESYHNFDmRDZ3PCvi2f+sknevF4DKO7S/LxW85C0D1q0ziL8FEvEPPO60
CnX5I+RrlXhk1Ed7X3bfCx2FIkS4JUliNgeTG8vKx1HI/ap2Gel2tQ8SIgNh9SQz+/bSePaeJCjw
cdKVP5/WinQBUFzoqdz9k+tNbfJASIWbIqgwRTmmWaDeAdBkfSaJvCwa4jO96ZOS+JKKv/MTCzsB
+ev/z9BCEBsHSZOQ0Gx/ygA/fUh3bWL4MsFadvFzIaLFC/C8r7mC+laeED9Ocn+0xCdtiyMNaAZ8
BqC18fOox/233bGmE59HxZCRbHhOcfNIBDJi4MUM091oHRPggj+OxWG+DJFuHwsHHHvGfWNHEzwl
lfGPxHMsLS9yySc/cax0hUF7HBJikruiXruXrKnFpIXyFSDvOqnFyKiEvXmAW4Yr6+galIAvqL8p
Hf1gxRVtyiXy4dB6eNjLGB2+yl/pUMXHKObRa5BM2BvBh1JQK3FG0/5A6DBDsz4/VYKmOl/YULsN
Ifjw2leYVeltbguwXPGAST/hpOv72H3VEobtvo3AjdQ0hNz+J+YV+VDbaoFVpV9GUzfHJlz2lBmo
bDX5Y3sFC7fKwPv/0o5hXOubpy92EG4u3+xxv+ZZq870zd8zaVbDjzqK+sqBVcjNBvhMg7fCQfUx
f09APycx5WKOg8j73+rccvK/5Sx/5hn+SWdC+hE3em5BatldgIwAYXuCe0S++5Lmk7sP+vLZNSbZ
fF+PGKJCUEUITRbNSkbOrQ3LKSa627gFrjN1b65glnAHR99mWhCi4tP/oREASxugGKokjFUtuUnO
balD3gevfz9cEKeJfDHW/l3W+EefzFVAuMAIzKAQ08m77oATIM99PZUVPn3+RkjTzGYRJ6UGZR2R
WAUumG04zX2ukWaI0eLoO9DybTA0Ok2RrSC0z3D5T+iXJnxEITYuZKOtLsw+UpQxtzmdk0W638Vl
DSGzvqQuzABMrTb7hlHoGgAa1BO+wzar84asMJ18gfHI2XqtlNyx+PY/AkM5OvzUxtOPJOMI+QIJ
k97DJvxIQ3eoNIrAhQ9Sb5iucYWnQJUlysu9UIbTl+ahnU4EC5dSYm5RNaNdvxQuu8xTxay91JjS
opF+Y7UrNOVhMjFeff9zE0KMc7dKYXStvgHCPPBZDI9O6ZpEkmMmACnL8JOtvunHjyzPmFa2ft6q
xMp2nhtNq8M7wTXOyf9X+9LZPOaRjxBFIkxMRpxd3anOVNeQpI1Z6/zdgvow/mGMnUhcbx87NwCN
W0UZFSltqTCRBEhLf9ts04vvSG+wXBcx2Ai3ZeOlgAzpwkHZ4EjDYALzHNOsfpOvaN7oKyzGJK5e
9rFTrchpeoI6tzvj7Mxo5/NotlHd8EbRQAdB2/UrqQZ4Nhtl9XbBvl2AdzIA4dh8iWovQ+T5cGTE
/WlxJM8zYYY3KUrRsU6OqFaXBZE2nqi9dxwFfv7BvGgOs6y/okTQyR5oIou/Tm0pQmr2dos72eC+
IhD5U3nsh/eAKgiZMkICNmbxtIRaFjsw0L7fDN6M97jsS0O5gatOXD29hn4X/pHrfhbJd3ygtHv9
hraLPPSu20V8eCvM7N+oy10NDU3ewAnsvaooZOzk7Umb571KNHrltD3D5YE5elhn4bmx/M+TPckp
8s54ZG+mhVa/PhmI5k95bgFmyjtoaYGBsqyJIbTKqIwybyJET4xNtlmxSGMWTt/GYnVIbtyOtDJY
VyrqF21f5gvdN+sgrUUh9Ujwey85+399T9+U6prKEhRSQ7qDFR2mIPY4iIUBYa5QzI3fogaw9ZuV
QgSGt+m7sY4sPAtZAJADUqDqULRRwIJleOYcdyHzBsUMyTTLyySYePTc9mQoqBfJTLnk0X8+RqLV
rt3SqOlkW4R0e7k+EPc8XrM8cX52MtyFTrNKfsITM6v1Oj1Uzq2rw6jXfNP+wha5VouIwNxIabad
U/xDp9cwHHCGHRUx9j18QvLzc2/C7NsMdQpTmCRxi239QIeVkrIUFg34C2zhYHNvkzFdwit3KfWT
b7Fq5lCUB5g9QA+UnKwYj6kWFMvB528t9uDZIHNVEB1HpzJjOtDarloxuE9CWj7kuxxHMFl47Kvz
J/J/NVgYv3e7y4wkZCrrvWCv9qh48tSVwm1TxsVIxlcwIIQDOXpKGSTvvWWw1ifoQHe02Am6R0lW
w1hjmRzn/nsddwYNt9NHgN46vn9CbaiCrf57Rtb5L+vO5eMhI2r13DSnTaou0DhP1EN6RGC5fVs0
jpI2J9khGYbjOyVkJghCQeHTY2GVcYPIrh9CLrwt7DzACY/Qi327Fnps56scKPDdgnuhXFxIMdAl
60pYj9OKk8DK8+ZmT6jasPyDz1TxL9cSDuoO0HnK27nXFrpIqjLDg91DFRCkIGEXSTBXJNXo3IN5
my6N/Jhb6TxRzLaI2wM77MatFRCNjFGg209VzrlDfEpXHjGUJ+CvzDtouHHaaoO1ZQg8bhd61VlG
ydd8gk+2p8TLbOJof7rZEQeyE/BkYvl5+x/gtcuvOMnymFt0kEDw3uJtw0K2W+9JCmUGuykCib/i
9hyfh8rh9KruMnzxdYtHobHhwrR0pl9ZniLMtAndxxZcnp/3YJhJxEyTebLCWNmRKf2y/bNzDdjw
WCAaCSLaUsPwknmXGzs+s4yRxBeUhg7kn3uVd/34cDyQW93aGUp0ychHOgRNe7V5ELiYC+tUCcc1
CKW+gE5Zj10yzigMp3AlNlPyJCQSzVtUjohkYGg5wiw9PMjPKx7jB/mOKUM996kxN+TcaffNeXRW
hWke/D5JDzJqMX1aQX0XWF7YbegFDCxbIxuz1uF8AB2y7D2x6KrXcOc6FKy66bSCB7HwtsHuQDUG
p0avh0nu1r7dAG4ulEbibraekM+G5cdjIBITjQ8GYJIqge5kT1132bwh+7j1hZgl9Ch3qo6+1hOm
cSdKF17+0mKnPTrPdKz8TXxLZ0vPpUGSDrWvbTHA2MiSv3Js8XrhrWpt6/Yl1IEzMWWN/R0FhiMM
16hocpinTYpNgzmamliH4Bqu0KWoyeiQOKhkZVZVQNd7JCzgqNENFGCEBjKWwVIumRrMsbJvHuyM
O61w5tkHcB9CSrBDaj5os0TFWOlmOGPYr/NGVhifpG7bk3ciXzo+7bYS+SxhOYmOdC2LR/0eq2f0
MgkV2idUEOmKBnXxgIGvaNoljDnjc79a54jYmXVp8vkVz4FlzV5H+lOqSbwgsvvRp0IQRrnGfeI7
XhFNCriZzJy3Im0vg6jhxezJ2wE4l5HUJ4BL4vVf6fk/J0WFlqpT5FissSRT+4U7n9cBqc6ycOQx
F8A2YIHYslyE2jTL2+ToQSSPsVqk0OGEFjf9zEofZf436mgtQcBtbhITTqiOTaMLlW/W98BTQejR
yPAJw+Ix5IgeBqvPqmWW2sGft1mYM1DZzvUcL0Ts+IC1h2rTwh5Zl0ASfhl6W0GEn3A2ghTvyK2k
/gyX+XUG8E6gSOFy8bjwZ2efhWR6HRqwhU8LvpmHz8ukTU0NnwoY9rIty8caBPLniqf99kgv3s/P
DiQpa6G84yCSbpRjRxKDJLHuGK2gfc1WzYKncSpGfnhtmW9rPxstDnIiiNErW/+9l6JyINhvYB3h
OwjQK1hAx0ZmppGgZrV4vKYVWnfGRp5zKoC851lHBXhA/O7BG8oASRkajbF2CcSi+OQPiqAqdDg/
BGEvVBWZNAu5o/+W0/JwBObpWy2x8zHjhnVeGFukO9Qpg9z9N4Ul3LbNHlLt2KP4BSLc1CThBfpF
XeLmfG37mvKT1QXx47G40afmGM5SuFxhOnJ8QacjLtBEbMnqBwmfdCsWeidBpy60qNCvvH8UWqz9
7JLeam8Grd0koF0UwAZGqw9I3Y8L6eHFez9X96tQzbcjK5bvOcM+14603UAD/bn3T6aHSONV0QlQ
f+LyU2RhG2r5Rl8ery5AmbYbrSKDsh4LRiE99YVd9/vWMREMXP7COgcSgyKeSMJQK8fFuMuh5EFM
G8M+6DFQfHv+Eb2f7uX6/WVwelwKpve298Sh7dn9zEQ6j9LLCNXQHq2tJygNVrgj10neM89ALAD1
jTwUWcBVpQdxbZuqIkzesiwYegjjVLcA17mITN0fd7Jh+8XCIM72rROK5GiZGfdS42YXIW8O7wIq
rvH7zxSL8i1497zvqmgHegRVF28ZRaZlUoq1e1lk5iX19aexZPc8mHjrqW2JeSZ0hCSVWKnv/ptK
TZJbD+YViBRFDCsYZaHqb8ey1x5pHP7iQA+4QuWTuDnO2zElNnknog8BlVMZi6UO3oRtLnYPRRNb
2rcy0QYVtgfvngkZO+lyI97MCbmbpxp/15RfmVT2ju3bNEyFa9v+9RptV0al8u9MZlf/diw88qsa
rcF3lbpWiyCl+zmxjXCbYkWtnXz080IM15Fcyp21scCeia+gNBks1IQRtRi9P7uscZfX4tarBv3M
MWqf5dqdiOWzwcQwgcj98ulNGuET36fnvoc8ugE5hlL5J9T3TX789zuZBuBIpDKJgGqT+xsqNkTP
fwTZVUa4vdUInAJ9AZuCFrPV7jFyxcLAFJ2bb31lrF3EdRCVQP6k7OX5X/hMIwRw82+GHijZEY8e
jvmQWFIdETeoVwCWjDc1kN5z0honJqlLRVZwtVLx9utTrwVj/4B1ysge0oVavIOcZlzcW0/DsguL
7UAdF68X+/McRfHtaO62//n2ir+x/5JA+s/fVU+F3CdfGrBWtdr7C60+W1I0o/9W9C90Cv3NJ+Jl
oKYE8w2b01D+h2qKH8C5TjDM6RsQ/RXTdpoY/WU4TXy7DNuvlxqugHPtx6w32CGHWmUzYSfK7VLO
GR3/hkol2CmaDH45FusL1Ig2JVIfHAqHhUAB7MIvBFI9mQhCQH3pqXMIulXUSc/lyV8NyhyHHvMy
YMsuFbwnEmWNwL7c+K4QieW75r1I9l2FsMkBzmedZDklJDMAQ52LbOkRHciHXfMPwwMru9gGELXN
L5Xx1NCFWW/bPCT7ArwBb9e6QrKxw9lMtCqgvTGSDP1qvumyyp1xuiWa73GJ/uyO/OpghrDNPU9g
ZQfNpixFErP7jzgU/7oSAVmvIwjgLJaG43gMbTn4ltskMEC+1He95f6vBN9Nujr1SRjS5osdrS9G
inMpCTZii5ZpmgTAeNq2GFpdIiUzX7yBuQ83rv+DrCz2JKFZCz9fzWfI07Or+G0lKhekK5595gBW
vKMSRt1JkfCrHJ9eaY5rqIdE8RAfUPXwzw6NP4IufmAiUp4/SoPXJX8mBFvlocdhQOZOInN/06Oo
+KihcnwmDVdX9JrKwxaSpeyZNyAc8Mv+75DYjhjjeEjAOoYaDaIRqHUln1K7xRBvH0J8EyxWFvi2
kiQx/IsL2S4cFxNUGtNHKmobcq+T2aUtGjUmL9Z6qIWQMuC5hDpU1UguNbLYA/fhsxTeY/z5At3u
FKj/F5TsBblnwTBQVLDLNzbFmVnIGmV0Fsbl6E1ma8KI3YUfStAeyg1MEY1Jmg3cNMTDqXbvPBog
Ys3jWJRm8JNSjdFyby2oQngc9KTO6z+ZB/xzwn9sUpRZ64RIjYVPkGmwAZ4uQzyo7vTSrtcotM4+
zMTzwqo0a46Ej8JmHIJs7YqUQMl+U1XH01S6o4we5DGT+BsHbhBFSdB30oUFD17HSUZOHqSjXU9w
2rQhdJa77OkKq/yKHNzICgn56nyK1KbSE2R6ZZoZhiFBtJo5nk6zhqwjwZosbVnkdGdtR9t3ioN/
lzJt7W9fMJxPJlfzArNxBWvSMv4HN2Ww6WdBCGNqMzRq2JWKDg+A2qup6es/PpqjezKeqBABKKQk
LhxtpbPaeqgROp3bcN2Sl2v8mtFzPgytbAhOq7tIzoVrYT1EEWQ0xHFEF8lptA2bycONvUh31oV9
jGGwfc3p0xe2i5JNTFX4trKgzocOpBf4kDUJM+ckk9/Pxe5sm9GulNxptMYvCgSB/KwnaDzD81nu
ZooksOkMVJP6bQ8xr8FiN+dxxvORglXUxqjUYjOmqtxltmitOLBKxNOHds7TyVJOWWlgwbPc3Q69
yx6ded8LBlPKlAdlufR7F3wAMuy1XoXJGUj6P7UCsgcu3WGnh5cuEaFzjCMb4SpOdomGxRON9OM3
zktWEal2aunAQp2P47bBmBn1xDRK0RULd1PeG8Y4mW8ZOJ3Slmt3FUvoKurmb36vp2JWwgvLyFe7
2tld1qTOsNvw5yRPsp+saN0XBrl/Ff9H7/qxs++FW4L75XPCTRKcz8xDwV0iYhtwa6tIgNF7/mOV
nQwcXdmR+rjuR4fo40TTo11hOrLcfDoO9Un4dFOirmURN/c83GEttq78LMJVpm3skO9+SB+OUeuc
IePlA4xEAp5eJMMSsckaA1SEVhm6VWPHHae9+FcITpObwJ4x4qIqSc7+0i1e/OO8h6Xkyq4esYJc
HOgICheZRvWqn003Dph7l5s02A83K3Lfh9kcjOaaIA19UZHMKUUkQYEw9gD79ra2HUHH4u4t3b94
5tdAbVDFIPr8aKWi6mm97A7e/G8ev/JkHTTPskbBDR0eDEgXo+QP/r1irti7lzx/C1VKgO+FOr3D
h+jlyvUBC72lOx3V67Ogqfccl54Y8OK7q143cs2UUH3GLciMF2uQhs8bzlBDjQUeJh42mDQ8pONN
gS+byZoC02PcGZqufkz1YtzfFGnD3m21DgyAX6FIPXZ8JR8z4+E9Hj1AUwdvAVP2U8qHP0zI7uBY
vh6xORc9vIIJAAMwzMzeBK5od+xwQGYqoVIyNvq8gtfsOlL5PdvZMWxQnMkitVO6hu8Cm6Z5D1Q9
AB+jOjQli8E/ocxXQpbegdj/9SyRJVzvH1Y0b95x5uTzroP1uHCeGNFBTt71LNllgD4tCo1EsolU
ie3fl5aVH30kRKnXJWeyHht9pzvTso9fr819uDMvLzvcgIR/VVzIch3wIVXHZAPRW62jQWgOtBIo
bNpJyfedj/K+p+N5H7yXumqHNQ7qlJTu64i7rCUmnA43LKa6e620dPoF2IPpg+dVyAyjI5FzTJVO
bKi7SH8yiD5sEnjZq0YPTu+6olTKQ5as7rF5r2awvQWLffe5112Qqn/nIccvTG+1ucyV2yqGB7xH
dqlMn74x5J0yOL73BTtjxouU/oB3PQVIV6HsajqfBzFbkvusMbgWyoThtVSche8RYLXZyO6WXbUF
zS7lbz8EMz0P/kWgXudxWXKm0ecsOKad/7Z0lAE/DpHoUVOUfbqAfAoGQct4b10Vz4vyYUyCnT3E
GcIGVJEQqp4wNOxolk1S0jB9UnqCcTpkGyeLDwRl0i3av5z/K5TsPZL5v4fRtHdLWuaYWkgeG0Lw
oSfJF0mWZ7jhtubJYytA4qJzHHrvoEhOY/K+J50eClWGWHfEM/+zaz/93qtehucyDOkeQLai1/IY
HLD4yi0XRPs5kqZ5hK05/zRgZpYiFD9M6ixEcG9QCdJHneM4HLCDuOB/O23Qjzir+OhV7wrwFl0s
8mJT8WAST3TX7mY8LrYMQE+C1TWNgJ9L26QJzweDJOsLSp3o5Sz0V8UpUuA0gT97uXIoPGj0RAJ5
/z2Lxn9nG+DjQGUnUO++aFNfmfd1fX5dWjh+LT++7aQs7aE88oU+JNBocbuA5DgQqiRjqkVpMcHd
COYL2GGds7RH4NHxUKN3zRjZ5oo05bUvY+Tceqq1PmoLrLE1NZ9mF1hfVX53WCaDotut+bxj7l+D
f21P3GgEVv73WbyZKZb2jA90xPixYVRgtki48mE+LmxAWOae5pDgErFk4bC+I6XFm6bvJ49KNrpr
JG1CZThtZI8GpfaOc7KyGuCxfjz/q8KTX5kwt2A2n1VMQeAFRqPscIbmg+RE7/SULINWa6kHnWOm
iwBEIf+Jxq6maJ2ewuXJpoxVmEV5LmfYmtf5OlXvZy2DYUO88adHZxmW0HohNa2zRe4j+iGIZ8ID
2JgUGGb9AvC7OUukBWhlZ1FEQwDRWr9q5wSVbPioWJ3iFDSLSF42B5kH3I5nXdXKGHAfb7BioYom
lJdxC526GZFM/9lT58tiYlFIoPs+ZAD0TYny1RA4rITC0B+WvuN6+l9TsP4Z/8lvY5/MBQSu4cM4
ifbbSnIiR0/S7vMVha56weD2TNTPg8h8qlRpGtuTCxRfF7uDJvbP+1m8JCOraN98ep2u8U+N5MNi
hWN56YHM+PGFi6XHVCTcX631eQkNO0BOPs189hIrycwGlHP3eupLovBHyhWlwmfdaqyVKDOA4oL6
b34fEoX26owUGgZqwBq2QZjtoAhAxcd6zr2D/a/5AufzVWozYxrLNChqplbL+HcwzKm57odJ5Xiz
E4XiXrDr1vDLdVn5eTY+Rv+XfBPpT8lMS09Id1n4JjBPzgU7CqgOqVvYV3lyUPOixRL2cYW7QVqo
hWjvLyEbPc6VlEIELeWMeD6GX2XxD/JWMZLUDv+Lsyi+Q2GwutyPw4L2zg5UAnKR8BanB+HYXD2T
jgLN2Z2nS+drAKFWvTpVZa7n/wZ67nqHUHx558v1DCgKqWuf8U9PsiPxSlTU58hMcbUQArrUhC3A
698tadQEDwBqO9lxrrJtNrxSQW0yAE16NJ1NF6zkHe7KBUQEE5sG+sYGkO7Kwz7IBBLycRGRNQQh
r23RDWTX33K57IyqucoGo7ZaMqpJhMit9AsPc/DWAzz+z2/lQR8iha24pfo5u2AY36/XPb0C+4w2
RnzPGHKx/tIJApbpaXi2AusGrlpXjJAMMKz7EBlXwV8BX7N9dkuKJ3SFRksmNUl2sTgNiIYceDLo
zocGm3SiU+HT69W3HQmqDuvjvMbTM9306nnp/xMVLYhkyZrNIPH049EtOZwXY1bxDDR6557AWjff
olsYTla92DOFHdxEpYs6ohffgbwTNq+inyS7KwFVAaky8XHF9viPONjB2MSxOK/ulpmoKxkxB25+
TMaZ/pDQNob2Q5E143xLP+8U0gvyeJpvxym86ueNdfefstcXwGZov1yAECppQ8F022mbA+akeVJj
z1WMmjT3/R935E2CSHU4LT0TzTMVPlswiHZTcA1lPF0XNd8/KE7tA6RbuGQjso2rrDjyLwrceG/H
07R1ZkiU82f0PcTFG3wqS5mq1l2YGF66oi+zfBfAeXw8mXF0ZsfWKGT0d47I4AQ0t2rrHZ5omWJo
Nc6tDjHSoZE7GTUHa4E4B8nlTsRqL75rIPJBvBbiI4QR5IPFvRLWRRAkDnyhfvvIrIlFbxVqrXRk
3PAqODtaB9L5doTnh04VDHJ7UQ6io0czRSrbpEcZZjMAoHd+kQecvRYyLlz+7XTXeqqPTEJEloN4
E7BNFhZ9GdAkOWXeo9DNeyu98Nkrp/9QNU1LUkeSNq/JmZMiHIS64+RlIU5UpeZaXi4jrrc6mUsM
xcRZ/Ea+s8XW9Sj9znjFVGIz6EMJyL850RuREfgEjHXMUEBpu3cicVhPDcrkiPSwLbXGi4kBaxks
9KH0WkoKljygXngX7npow+01baRXRZzF011Vjf6sn+oYkqmQLt33zjYUiwRHZj2vNmRHuIw+60nT
Lmd4a7ysu8OMYshxJI/1twiehaKqx7PxtT1JbEmVdaSyV4yNmr8qxegcynOHKKYWtXQ1EaTMUm4f
hqbsF+BMAcYQg+ve0Whz1Sx/X8TFvtmCAbwI2AZ3H6X/baQLWLrnlgordBFXh6ZSvMxdorTwV0wU
644htwrdji5yQlyPN3BZlKWWrIS+TTia3XxyvPidHjWTjF86l0ktvu8cIMr8D7h0LHCNF04WhCOJ
jWktSPLAAK/zkHPYjQ+Rz/6oJXOpujXui8SGMf8Lf4e8ljflklq9CljTNfySH9O/Ngf30CQKWvui
Fy4u5sX4RmIwJMJc/+gjWOHZWSnz108nHdbeT99TocFqLbIGTd+4bb86nE7klyFXsIQBgkqRPziJ
cTu9qJhz9z10zYEwHl7WY7+1M+tORLeDE5Um2Vgk4yrZ33+16fjZWoDHvSOl3he/qu7lQWrmdJ+S
NhIJYMsnV6PkWHOvNWXs33vt+vRP/vumI8FDyEEbR1xRNBBN/TQfrsAEqZJ+BAgo0EEOTpEkjQnX
KfXc7UVYbJ6F2sq0/gfaQpSlZNCA2w9PDBC1YCO/6eFpJXdTncMM+ahUcr7msDb+fO44d1I5bXOi
/6seoXTTwyOfdGJBW5sEvNP8G2qN2bg+yYFdA2kkPcxt20rd88N8gaj2lGI6X4aF1+3Hsfg2YqbT
HGkwYkPe6EGBd/zqFD6PkrfO+VGq1yaTqeVlLbfAB9GxO9SEtuFxa3vN7trIY4DiAFtHuf6BSEGw
gOk367hHjV7DWHo/1tRygS1ztrr+F6nv/c41RG+TOESbAhrbluConlYdpFk5MFkT69BppBWKyyzl
Tkf+RJUEUPB+khgYSprMeLiwfixLEcAQN31YOOoFnh1X3yZQFiIEarWA0I9encbGqB15SJmf9KPm
gY/RDxr+6ZvC5fI8b13K5DPjxy+Z1OuTyg6y7ngZPLd3/4Mb7lEcpuxyyBiOaz4KGbxqGDlW3hdN
aQRCA9smtDFEDobGYs2C5nZuTtDEJZVSEH57ZBsopDFm6HdtKeVqLb50V0XVBAPsSjM2eD1um2ed
oI+IX+6Lwd5iwlOgHVD+tdY8j2tYKw6zwzyCrd133SDJGHPIHwgD2O2i2DyyftGsq3pJvwaD/OWu
/DrMMVTRJJaR+HkCllbwMv7So8nK1+vrlvUMLhVVz4zSBmlCRv32sYZ8Ki/4LMXdNnHYFlA2tMwm
T+vW/Ci46o/pA6Kxnob36Wm3HsFvAhgPcMmHZ5O5gzpcDpugpXwOCcBBDDgMcdSDcyE3ZOV9/Izf
FFl6AXsccqg86Xinydxrh87PcCuvb2XejyUYF1R6YLiX87IxQO8+Sc9YWGpV5qwjZMDi4oBbHxnP
oo9dgP8fGqqNcLr/IV6+KeKIJ3V9ZEkxcM3Xl0jtd/lx7EE97MhPeEGfJ3P64aW21mg1VmlX4b6I
mtzJ/1rVt+4A+iNCyerOE+lWIbmHRxrbJEWSHST8tYaHhbSlzNRz3MB5CkmOmm0yVE59LnRHFNTp
KfRLZGDq5F8hHIV1sC7ZYxsswoY6IyMrzGLGr/bYWIn9hxNT2r3bhbJAmfBlYs7KAGU+yOBNau8f
lbpcyY2kAWOVxTCDsfWghcR9VCfEjEMBLUzf4vWarpFLPIgDugFKgAfwd97Uno/Emz/6okRQvX0G
G2rFUG86HzbjEGkf9LTIwhY2B1sJNZZQEzElPtTIIJmvhLBlUiDse9tjnLdlNStu5KrMeBxnXjsz
tbVTfYGOEXAfZDIgStm+FfPxilMkjVTLM3XSzUB7o4WY2ggJNiENMEqxfzhwrQBdYg6MWZBfeGGz
7XHw7xGw146KrCPPt9LPFXrC14oSsQS2UstTmXjumAyDJ4EE6HHcwbI4pzDbQRodF+PFm1krZPe6
fysKXIJXLbiaQoU3kYHZGWMGCxWqEJXA0DPBByjQcU08cNUtCKTY5AcCYmrkXYV6jjbMY7hqz9DG
+84/K1YyQrrgutNDfH/yMaJh6K9ycSdK4V5Ig3cNX0YWF9T8rV9W/fKxXc8CB1+aKVjEuPc9pQO6
JVmnWWtx3Wv7yh+2AuOczpyQ9SPw48gdVCP6F0Fo9rIpli1wb7Co3BTx4wi6rRF+Hb6rZmKmXm2S
5mY7XKV03kACc0OVw6ZSnEjhi7ocxxTr898J5dxdbE1mKByG+QqbwjcQFNRFF9LJGadgTjpuqU31
/dhC5Rq6/SC02Ul5lTO/Gp4KNHtnDZTnbQeWsY1qEsmdppOzXZOHrJloZUCvFpwRG6CrPrrFNh5n
YckdZslq5ZFYfswPLlXIvQuyhwrSQAnLEV5GU1oeKR2br85Eq7iAEx9E4/2DeK9rKm9a0qbArFEu
atbrofvhOKYRe2edI4mEpt8Ii8gqaYBdCwZT/wfgSz2C6EEQwAlELwt2xroSAmFz5EBeiQk3ltwh
WWHJDS5RLK1ZTk8yP8WMHFCtIjjev+JVSS+09dEAksg3c2Xox8ZsmCTgmbI1nYdHBRDKbj0Yc2F4
tLHYuiMaXu/WbQ20t0+OqXnkan/74+7yft9sWX63FGbRpLh20S2dqLWQlTjD70+/sO/I2/QC+piM
3s8mixJfw+KcnygxO7UZRyEUwINDvnAmHJegGfUZ4Kds7zlX9nCw5sspdI3YCl/GuE7tXvxqK8oE
rKoUuL2rf5p7bYaHnhJ3Fex/be7NjlClxAz2SkrpfuKLtLWHd7pArAyOPGFuYVPfuJR1dJ79PIT5
rJxL5B+DRGreds7b2b1/emuJPZgOcRBTt0QS9bin0UdLZglulgvQGi/9hNP1szlV86F3jme3AD9m
pLG545eV2k9XOC06Ie6EBPcR8jbrGp+x5bkXfmIk8dMymlWLzVZAYMgjmYXNx3hZnIaw8ziVAopd
i73VXKyoFM26S4bVlGMG+zZedEElzAY/FNN6JvCacr5/X1h8PuOzDe1eykifpZXjbxB6w3ho8B1m
X9YsOu1AgC/ZnsfoSv7kXTnHe4rktidSLVAWQHL9sykuAKE/N+uhyTpiU1wFoldyQarGoqoSAFH1
yb66JDlSsDpOldWRqM00INjjQMq58neRZF9wQcvYiVO/6KU2YlR8vNMGYoqGsJow2xAXBlogZ6T9
PHZcHnVo5MSD7Iokf9RahWikXcDVkeZEzL+AI+Xzu7l8tgDjp4B7DMN2MRwIKfNgHLeFtxGzYMPo
cjzaDd6/WbuOENuvRmYHX6m+dFWsAm4tSVAcHKN+3z0nm6hcGgFH6Hcg+vk8HA0PNOByttBNWYYp
jUY/AW03w8/lZ5bteIVXVgbmRDn0QncELM2b51qRkGN5xRcJN1qNL8sE//TwKM183FIGfTmMASvJ
DAPlAgAy3nQTsLlJ1DRx0TqRhJTWNlnsJWmpoozHQuN0QsSvPziDUrc+XUDrhlaBobssg0fbY3gF
0SlVnvCER9t/N/AZDQZQjxO+80DQIhe6m05GTBH+IY3jGt32ypTSLDc+/vTpY1JIlRrrDrdBRwSU
khDj3lf68tT7WPDO+VOKUu3KRHm2XD6mVKCiXEM2YF6hyqGQjMvNq4tT8Z4s9GYuH0+faSDxY0vS
m098+/tDIs5D7t87a62cIFQNR1bj3XtIT+v10HOApJ7SVBqK8YkcWDjO4n2vOG6engsJbkcXRWTJ
m3hVFNhmwvFeMd0Xh3sq5jCme+zFN75zo8Larly71g+8U0auhuKdfKn2j/yibtBiz7xpzSrTwLee
uLPaRNJMB+jUgBU3yyUebCki/tBvMOT4LqnlFHzvntx2JAxTtM9fKY6cqHclu8DKnz3Z52zLdnon
Fwo3ywH31Hbm7dtFpbTXYq3tZe6u7eWueNEeEwOt5HgX7WLYYZQ4k3oPZrr+iJhzWWmif0o19pUx
tiG4kPUTJzrvnYXosGRl0xiEgg2w6qUIwcWxO79EvI3zrZk6H7ltx3G6DmM51LK7xmw/hCVWYaYz
5yrFc5wjoAQLvEljDz4MzObP1YDvQtc5ZSy1tnZrAs8nfNy8sleaRJJo/E6gqVPIDvqN/+6PgDN1
ZtSDM0YyuNbJ8RQ0G6O83z4e5JmSoyGXK/JCvDTIOJ1QHHFUQ9mw3dRnTivYwMBn7TiQO9JG6Wji
CvN2oKF2pnzJfRk0VDe2oOV+3OyIAy+3unWxA8ML1GO/PDj+Xi/mbP8ndchRdAr3CMeyCc/TUZsb
oac/NjqH+ExxcmkRfioXD0LYRYketzk/bu5Y/LVH/6dsaPy7mEArGgl2RVuoAZgn9JtgK5qX8Ozm
UmHXisZ2ZG5B9HWusnAZ0kfoLzx7CTI8HKzkZCXyuHAvsEdtf6h+mrK4IOed2ylE3NRBuHmII0g1
t7hWF6Dve0c7S7E5QyPwHF5uNcPuUJNniQ3c2ccYBrpd1Bcq0nxcX9iMbKlW12bAmvUWfgnqs4Ov
nIbD/nX8SAtDeSxP3RdXEuwyLXFBPkkmJuqCKAg3NHrNRO5KAvwuwwItktor2s6ByqXuk4ZJ7PX8
pfZm/g+mdrRv10WYFq1l7zY8jFHTVovmhHuH73wzCWV5bmzKwWOZAQSpNZOFmdqu53BxdHL6etff
9By+0M+wCwYrTSK1we6ynt9oSvXxuvFSwlkgUI7serk3Zophsi2wfyvN+ik37u1VwoKFwfb+HFRB
mryL9p3jReHSYOlGHVrL9OPjLBwKholXNipwGhn875eGhpGoki62dfGOXAU6aWxK410fnKFgxa45
EKXbhlyJGUxMiLRkUF4MqykvgWDIY7zMaN2ZHW2/INrafQFbQxfVByhvLGi2AOa34AgeDQoK8vg+
Ux+FKT/JFRSZRP+TvOP6SVHgC1B9bdUsEZbH6+YGX4b6g3dsE5OiG3KyOyMWvzceUR/42fwo6INP
DyBnC/SpggpBwqj+G5i2tuIP37k0xIiep4iqfeR9Ze6keAtkhRFaCfk0DbjxvkeZHnMSPbhTZjpB
RFF0GZQNRl+4LLf9BTRc4LWmQo7AMjDYlGjZ/UVm9+X9IuNp0vqFLmQy7lF4tksWygxjDiMxA9tY
ZzH4FJV4PXZFNGc0kG9X3IHNUC/zHNmGUepP4mYLcTvpb0ERBNR66nWa5Xi+7HfVcRC+TT1nJomr
eIN/IUhsqgKTFTNiAYFNeswRAQcNEBYT8ASOO46lTqV/Ni+v8RZxktycHCgXUFzIp2mPKFxzt2i6
KY86PB4BYcPAmrj61JLs8+7YkdxVK8RmPwDUGrF+yxsfhyv9ywgMT7zBAs8ic/p5D6Dyi7+Z0CoX
ClKOqej77o8ZjhJEj66kmK0Rhv6KJv6tuoM1GRQdaHxrcOFWpkXTsbERtiLukIT+R0zEIQyQufSZ
VORKhipqnA0ndCjbJRBZuLFhzzMqTEIS3RsKZeR3qtj88jCvPxsMbw9slKnVDSSzeMiUjaoMsq9h
uinNtRjbx05H94qifKSxkuarUVzhRh0tRXL4bEaS8uVBgb9ws82UWv4sm/L1PduFhjBNlca6pdhl
FdlqF8jPN0QDwx/qdKnDWCMEfoe0ExPkQLI+2/riDHbj9ZnnT6KOSPMiRdBCoTfvy9N049AU7y9y
IMgMj/JO36qTjaCFSwaQ7YkfZeAdNKPERtRcWiPANY87In/fOwJNkIIQ7QFK/PKaKoHJkI5JEMqm
v8JkITkQXVe2p9Xay5UnTz+swmuBw08kZBuMFx823iv3gs+BFCbImxwDKQEAqBmyTWK8uE3YC7s3
G4u0Phbh+BxURhFZvbDEJS1/XQyK76QortyuFasOeKAtJeLbb977CekKt83IbNLuujGNpkfWvmtj
NZ+qVwSgfEhv1ZP4lGy4y5USneLlpds+jl3yGz/hzCl88e0e3gvVYXOKwSaJ6E6+1oNqfDwZ8n7o
dG85J8kPK3/op8lhxut42iWKb2lHGWmjHB7mbTmm0J63s9HOqekQ5lN18pvjtr6ohocplROHhi7+
a6RK5fR3Hu4CURLzJ14EEBTFHo7EiqHjNjBC4xCJ+v8WwnL/biWZnJe0MKrNdU3s+T/MyCiB71Md
vuS3iEO0QmjdJUTAgScGWCDcwpaE16U4hdMUFDqWEWTb+KUaPCIYVSY7L9p1vFAtaskOup84mWsS
y1DNXMux+VHib2Gs2fo7U4QMHrEqU5292GaN/m972i9dOx82m0qEznrSpx788gOVfkX/hIVfL0fu
qcCUSyBRWcRjUZgsU0n0qbFFJ+VTbQtOJhMA3vE55pX8ah5AsyJ0xTQQ9kzwOs1tD45Vc8vJTLxs
cWk9I5OPzyQHbqehqY33jOSmWCjXkEb6jcIRR5+YpAgO5H7cWEurPmOfFGR2MlSSRf6Z4+h8WxeM
w1EQFcPQXJKLTAkMFxATpJSUnfVoltF45ooy2FLGnBw/aki2UaEHVko7Z5wKThkU3bCcZi3Dz81z
5kLxVX1+bZkSGmJP04L9K2Y5LmONg8S5tAiKqRc47KhH6vpHJhb1ik8PFQJMw7ynyQ2NdwjBEcg2
2r4A0pgZ8n6JJz+pWmX9IcXu009PbrYUNEoIco9GjRFgg2Mlm+olyjs53EFWZaiJn2g9mBum68iu
SWixj/BpJa8ZrHWrCbRH6x3Jkyx66le0qcHt4gzr7FMTFNKPtVdi8WidZi2dfHeF/wnBU55YbHdt
q1oHgw+22Syoyo/39xAWIExYWsbzp90patPRNYQ6/UM760kvjB2Z4594ioZYqYH3XIq/zq5uV+6L
LARD91RKRWTUoW7/QZlJZ35vlBibJUUFHYTlUZX7I4UCNk7F+w2nVWKRhWK/RyKMPYpp7UL70fzK
WKHxWnYdZhP8xNvi39K3tT/zkY3srIFOERQECn2Id4T2AIzibPRpMuWc6Ii0hdsiRaXhBKMbrfbj
/IWIsW5cFJSBC7L7TIy8hAlGeu+cEuHLv1tCAFjvaDPerCtoFUpzT4uTuEBGgqNgZQyRU8pw3szq
eOWWCj/72SUVuftJ9p8aEmU8eOeCnVOjy8IUqwCQoFq0EZof29YO+IF6HZGlYUT6H+buRNwh5d3B
c+YEDIo5/TeurY5Ls/QOspfK77tNHoLKlEjDIN5q25qHqzuqvTO1Yc3iJ0YU+1GJNXx0my6ZgwXD
FpLOM/FP35GGai2zpNiWr3C7TK/dqKGmD98iuwCrtYw1aNP+8XoFEviBQJQS/2LsNM+ynTdsBDt0
RJGD9Vogs258KGl4DNfQ+s5AT6D4lwcxXId6Wls2la+rcEcLIezTPtbY1x2MmQYKp4XHhVvyHWZK
HQmC+Zliya/6iYS6DEDTewfJDHu0eqlucU/PcLVrM/2LOCmqilmBjR32WisbvECRxRnGKWGFAZCQ
Y9MhUXPvvbBehWSM4OV82JGBBInyGDcZh14ydZYpjXNszyju7Hy31ogBaAJX6M8YJD40PNt2rQ/j
EZi8xYmojCTPH5M8YXqF68ubZl197JMT6lfGVvNJJNeBBnCaqmu3zPRXHRYEinnq3FpZfxO89KT5
Oriedr7YLILgFf7VMX4HADnOtGeQPnbq4/5M0RGulsKSwrnaqaLowLgEILcFz5dh50aX3IiG1jdu
gxRq3tTRF0mFbUaSnFThBa0Y7zFd8dQR0ElVWo5fE0KXO9lS9UZ2f9wJX81k0ht+GFL2Z/pZEB7l
w3Xgw024IjwdDIMKkMrc3KMOTs4m7J89ek6ist3qnDGFlbolexiu1vdzoRI6UUvuJs0aNDmCJ7U7
8lpDzOZkm0Z0hJgATikHcYXa8Yj8nyFa22r//lPXQBJTkw6wBbcX6y+H6qKKAjVqnro7ZgR2X2Zt
PdQQuejXQiPzEsNndC5McfE8smc5/YKlwDt+q9u57hzDzSSMOG0JKYSp5VLqUhbCO90Jte8rRthA
P4h4BPLgEFNZqkrbAHoElrXIaXtTWduaIFNyJh+BsXIwrYJYTWuh3wPZLX6fsOeZWVec4oMZYWeS
GqduxjTvwU0UQMm97M+mJGE8+Qm0qCr4quWt2vdbd8cX9cyqHnQ+mEwCG1kiiTWYWVE1r3bGnIUg
oJS300EoB6pZYQU7hiznbDdIWS3fOgRUL3S/YvJJAL9vyqZwMC+X/QkVTjjNKklbsZ9vSLq2n9JP
5FzkRgSt090fv+vQdzlSaoY8cPlwDy1diRZwra53hbCmFHq46+E/hwqm08dWpriL5HehSXjxFI0n
tuGUW63RUB/YzwjcyRNNQw0GoCF2lw2Wvtsw1R9Axzacqc+UivC5qesF6DRHODLen5gtg6Sfn+oh
VUpuWDdShDBKu6Gj/l3s8oGYOirhXYjPECFLse4UaVnHoReDT1LsLLxqdfBYJdWDbtJD0MalhnfN
h1gfru7AR+lTn25Hcu/K/cNaO6dLf0RvlCdLD7Tate/gJ4zO9fCy6VKFsig+HIwC+0jETCE9A0z8
nXy8eTWS+zR5470BoVGosZ1H9aAkHL5UGfMnfidxeki42RExtc22+XfdQ4vnGsyNhP5pGMqFijU6
/Y/T71R16XJifelX6r8uAQ87Ae36ZPdPivcZd0VKWnYwDmDFULY3Me0+AfXq0tTbVPKvT2GLdwGq
FxLV+94MzaLUUyoGG7fvIEXL1RkHEeOMDiai4ghcwn4HjKtUUvNBt4K/YQ0kRoM1vjavyZe+oSLX
GX3G9E1Q6Mg+sufweFR/XB0ULMdAs+ikrb/J6DuxMr3yWtcyRJAph5IvJAkzisHYo5qbes2ZV04U
bKWU9iTXzqfBEhDnjfivOHuSovRgNN4tUhR+3ytvD1i9kQGAGUeVLXfjOpDqxWmdGbbIlhRFn/E4
nqymfCrPxG+322szk0mAnTWBNqfcSuA6e+XOwzrAspGD8Z5Hx5P80DzZZWnXsm214rxuWpGqlw9a
86HYd5ijJI39T09dD+t5DU3c2vUrwfOVXYUDt3CPsnh4omzVRFLVVUii8K7B5L4+VM9GYzZcV3Mp
EALsybSd9uj7PLl1BZzaXe0yS9gHMj4aSTDnel1Vg9kM6YAcSamNIQA5dGTG/71NJh4NmHww1j6L
LspYMTUu66Y6eDiaIuid5yZV6NvmhHPrDG3RFjP8sffn16SydrYGPjh4gTtg/3CGgyfM020O9oes
mohpjUL6xx9X0Or9ycX5TnvGeB4czs0BEpmAqzyyGND5OsHylmBoYAXzvlt9SsbNpLiz1DdB3Lu9
hPGr3ZsQBr53O3DigFLS6NAUf05gq6AVBffXPJYRbRQW5THaxaAIOJKEF+fnuxBLuzR2PfTupWSE
IjN7IDgWKdeGgmMKIu/PjqHViLJly1v2xTWlzLEHEFdEvVyr/6T+Mxu80RgDTVFx2XEPf3PQOX6m
T0llacgXJLxHv7mdYD9GuYYtvzR1JTBhz1+hO1Auml3K1SbYd4dS/y/kwoCBduLvqeD1z7zbZWd9
EEFuyUrGyJ/eNf51Uf3mK50wB1NFZYxxfvUkCW/4Egt2RGD/tY/v2hNnoqJaFQbgJK1ZukQkIc7J
HPARk3729K7vk1YOn6ShJipDvAftT2Hg/1Ra4VecaVOOKljSsaJski9Vk91hBQyHI+BbMjciWBci
yKZdVb5KSRSIYmOPg3AWxRqqbSmthgNOjWgrFehNmNJHU7cFa/amNCPP/uFKDLL6mhuU7em0DoGP
Hv5AuL8RLL79NEnfmAhNe3BQf56gXZM3Sr8sG8vJ1wd5fqK+h2QwClatkSY/yNjqLU/04C0I3GxU
1TSHuYIF8JSg/FiyT1m2+tpmW/3XlN49ImMAJL5z24Zu3DjIOB+MHcut18Ut67TBwh2Blv1zskBo
sVKoZPXKt2Cxa0c0ywtCd+IhBQacv+wQspO3Z/u6cvTkpdKhSQrmEPaS0Ky3vq8cuaVu/auKN4AT
9MgSpvkVqlywiBBGKOr0rKRerroJ7vzzMdwQtQMXIgCzP99iOddUPDqYT7MliaivqngVSZNDS1yJ
CrQdizMNsbhnrcSObOBnOc8JcDM3p9qO4ydR2/Cu11+3NULPtGh8RiY4KAVpW/YstYpHN8CpUM8H
XLRhQU53btBgWwji6MjFMIq+C6MxSjnQi0K8Zry/nW1HXd3Dmm9RSUcEQ9oIvGocNqwHNR4Alamv
ZR8grQURawFKrAzY0QoCrBwx6CBeIZz58wJYXjsmdBsWGlwfQynMx5tKmzPBSv0A0hBsL18nH8/c
SBYaI4gfuUTPbMGH+f7L10q6lnTBkYqGcIff0pzww1z7OzXHqwgNAD1UcXELVWiBAOkBfyDogb1T
SWlsQJOSo6/FPswl39lH81J+lwyw3E3qHfcr8KtwHQfAcyUYfAvf9SJVpdGzKgSTASBUdCtGjhYJ
qghR5yDrXxZ/Y3OJ08tH/rkEUont2aYXGj6XSXF62XNoqh9csGGnmYr13vJZKppRBzgs5j8n9+sy
JaXMb1IloHts3/TLBy10Qp3V9iK/3emZa1RWke81bgu8GVqDNgbX54D9yf2NONPixhD8BgyF87HL
lwo1yNRUoqfHwRWYfQm/0iQR/awUchUpAOK91yB44QAiSpK+sxm66ZVsvMxvOMZ9adIwrjzI4Izs
7kaNlCiPlN42JdtIq00Xb6w/s/9mjBI34O+/cxSyQYW1rFDZfrHkHN/jeFYEQYxb2TnCnZR3Aixh
X4mp7mE+R8/UFtKwl0Q7TbAmbsar8Z71Cq33veuExkq9YtRExDRki9vhYfxlenoa7A/ayATw6FtY
SLxu+siZolRHamkn+zkRN9tG/RcCXeR17AhyUhqO/pICpG33wn61DySFI/L6q0tcLpcD72I2W74t
x3GH5XFf/jl7AEfT7IJ2rueDsB7U5hL2CvkbPlp88PJSHPQmVcMSYmJ6hr6e05NgoBxSyyYJrEL8
sezvBLsK5ktBptZl15SBJ15dBqQHGeInukktmZObzZSuSD+RDYK0SweVvLdF/DiE1qagTptpbDAz
6txzDu2GYsu7alvo48TmhFLBfKcultOLBHOZJTgH5vb9SwJLRPDbu8Z+tlIe+r/dJFcF80D0g7Pw
P25b/wRDPBHzW/WzH86hEH/1M1ETv2NRJfMdHQY5VPHvI6Qz3/35WrjmrIJWFYGPEW+pusd3DsMA
8kmbOO/nLcxuIDWgn3MXJdaiKWb+Zy0TJJnVnhskBFmtux3gYE+nB3TugXsXb6d+cxewcIc+1kE8
jQZV7m8Xq3t+EQJ9vhp2yCI8x8A9Dv+iThfcDL85HTR0XV9zDXiHyj91ZHy+HW11WrBU6agRN4vZ
Jnro4cyMwenCjHj1Ss4sjA+vaVY8EWi6b51Z9eXgtt0JsHGodyNpsTtasARBO3JksTEVwXHRcZpL
Q8lNjoQfnz/M/H/18htgJvf9PiMeDy4SXFRtNgOvm5yc/Yxxx3W899hdMQQ5ovt0OeELLBEqlsBo
yJ/vcPN3wQrSSfhrCkaSZ9XG5ivP2uGt6ziQhJsJczzL/b+fF12XgrFNkecigUd5wRgjT6dCs0oQ
QnmWjn/5Kj91T1jJYhI0gO0KrR8WNH1WEH1ZPrnZkXoomXbsg4X14ulPchxbwF6yQW3NFqez0Z9C
Sf45UB8FkFMvMnqjzGcD4x/VUgCUtyzAs4Lb5ArVFalLhprETqyNPR1SRDDHXF01b4jWCXa0f+j4
D47hkwkR4x84qcBA1hnTXvgUPkj2McW5A7ms61zhsD2MpSeuqJy7k9BPBY5HHwi1Ev327uGEIqLb
21iChaWRqybJZMwwGwFGgI4+xzxbznAtqg2/2yMT0uNyhnFnQXgg5r2aiPn062dRSVuXAMhUBov0
eWsfCVsddN/j+7T3XPHT3oRGWML8zWKaluOFWpiPbGFh5iopFBUEqF3CfHDU+5jeR2WLREgJoxrr
shiuS9XzX340+Kr/i4sWqt4GD4PuQXLsVrZqn6Xil33D0xTNhInlMjywFXRbNSPC5UVqfZLaqmsC
gIcqez0Od0Og/PGPGyDDQer/nCu7I6gjfj+yV3z1BM1RYyLcCRbkZ8OfwrqeJj2uHR0u+SDw3ynb
g85hF1VS68SKio2/rlAL7sMoSzv2rM2gd4kc3Vsk2V6qQsorlz4oNOfCDS0t5RT9fepy1+IG0oF0
prsrnzdCnb6TIL/51fdt6yVZ/62xPp56TM12HiTUoW+HwLQbr2gBq5htQswJUjVwRkl+nVv35e7+
2UKBumIJRtmOU/xGtdrpzWnGggt6xPhW5WXeY3mboa1QMZ/UqBHUXM1xqmwiV3Uqa5nH4qUzW0zG
7taP6eU54Ptx6ntcO/wO+v1cWY7ie7B4N9HXlMYavPpws5me5lBT73Ml2eZsJVu9N8gVlambikQv
SEmYEn04d9zcWdQPjoqeqmUQZV89OlUgCRyLuzEve09vlgD8h4VHWYBorf11I9W+lJjfT5KfPs3A
FWpeJRfQCm8LiPiMQw5jF0NIZqsOXLJui5xw783QTK8UQCSLLINFHS1fesHbDIteXa8GZ3oAHNBG
JkdtrKbFpA47Dq8hVCIrOu7XgFC56tmJ0FlOfgo+SH040aMYG+8Th8QA1rZCI1BdE06oRG2pDgNo
p/RZE25vrUXAokNBMyE7kNHTiC0TqXbmFLr6QffI3jLexD9QJg3SV7x7YJ0lFfA/y3uxobQ7yqu2
Lms07cpTkNDY7FjoMW/UjGChLM6G8eP8wRIP2oe0+zv+3trcdKGITHPNME+iQFPlMaW1LnSWwrup
7vXEtpEvkqpNHsbynZaHbOxQim1JsBz9bFwndqQVN6TJ1v9q6if8yx2AOKj8SdDyMMI/Z5XSEroG
Apg7DzVgcvCic3xD3Yx4voA66zDJvjxoLO3unah+tcmzYC+Gnfrf8rJ5J00xKcG/mZoz2H9K5vdU
OdqdkW+6MVlRVnUXiJWd2n7OE0AHgaQ8khdzuHZ0Yifzx+5Ag12XeFVTO9PNIMmnJU8jce95QJ/f
pTBOGNfwgrtvYYodTtVKL4dCdnGnpO5SwsNQl3KsIebGlHGa2LyXc18SStexgYohBzBpi3MPEvIT
GkdXc6L4GkZxJy/8KcIU63frl/Lf+UbX3Fl7drOf/7uV3taNuBJgY7t/yO/vaRX8XDg8/dFAADCm
rRSx89SAtWKUPxmC7wYyoF2qrfJ0NTRQLjgj8h2JgOCEusxUAIdECcxe2Z+UDv3UHDGl8juF16jc
kTDGyQyqQeD0x0azKDrERsMOkAYxe7foz3S99uFzIu7qCyE+xrJgkUwkYT6q+3mt1zwPSFBlPo1j
P43Psdr5NJdb47l2YWIMLv85PfUAEHkF8+Jhovf80xm60x97L3IerafgVOxAdlRMmbv4dlJ/cZPV
JxegqlMDDQMLizDPWZQwfCuRp/469m7oKeCnmWb35CtM0CYHRbUBrzIu6FXECS+7PsyALjwAC6BH
A94gwGjp97ZwKW/r3X+YrMBIzzGPi2WpKHdehiLip5FJ9YDNEyogWJlbee+ZhsORspH2MsDsUz0h
eoko1EoBw0TbNAXMY2ZVGLDxYxV02nbNll/tFw4Zdy3wV5kalrw8MXpe+YWz6nCEHfGes/4UXLo5
cWo4V7dpKwNnBECtVenz1IsO/TNj0B81lEQbIazYFWn9d02YIpbR+Df29bvZ1/Ryk4SEOpj4zeG8
oVlaW4TiCWRiTZyHP5AcKdvFq456JnPH5uJb1hqD5tzbbmGCNOHqhzfZ+X4L4kuZty6MdFxKDryx
XOmnh8jQsRqSw611KJ6/mU88u/Kf/ZiEziiNzCtIZFkiMxFy99jCvB+ruxQRCg6R9qyQ2ybMiYeb
DVHqw5a2jfMWxSKb2RbYz/EjeFBcUuIRspqhKUTKXmqpahrXkrKXvTvkXfnE9BcJHQXPu/3+cuj1
BliqAG7wHpWYOlNb/2QuCx3bYj6z4ZeuE3FE7ZQQEg5jh/+77iDMCIq8Mzb8KSTiQSdgGy4aFAtY
qUyAmu+XPAkMDu5o8VTq9Q9SvGXLkfnr4LpMD73SlgZF3bBDpbMykzjuRGWD0daBQNDt1uBgSpVd
3rwxWEoWvxQKFeg3giQ1eQ66kKDjtJItH16hANdCyb2LAbIWUSkzHuMhb5f7vuZrhqfy9YnVegNj
f/iOR27oEJ1ufzYXT3InWC0cvpB/Ekqng6o16WXzkreLkaEYbZ8PCMASMNM/OACikyNPn7Hu8hB7
vgz3vn1kRFeJuFyZc8lAwvBYa0spUu++WqtXYSmr043VTt4viL9denxlbPE3OXs+ydM4m5aUD7av
UqcMaVjiXL+beg9OEcS78RpB4jeQz7NtebOpCbY60rznbYQIg3xdt5AuEsqzM/G/qIvC02T+b4SB
kuFT7P/JfRSAEWlNZsh6j1jkTCUsqZ5PUDNuZnxz6SS8JldnLNo5UViI8gDY0C0ClAbbSE6MENMv
4Rx7lal4DUtZzx0tsbChGBtFA1CwyJNPol7+TveFDavNxyAeANFk6ECfEvdgevtwAAonsoDhzLLm
puUZz1GqV+eZtVUH+bQzL4RUiCNoPDQz15TFupLKXt5EpuDf1e/aGG+vWym+G5ujPzbfvswedvZb
3PkrzLlgNRvKLzOm4K9/4QnM/3g/ijiNrqqZNuDiDKrvb9WNy/K9MVL/dbcQz+Y7dclXv+59zHhJ
AFJ2O/kC6sTmRGRgL0b0gLL4u5+SOub/sge2jwG3CWse/U542YDF589eiQDZoCOpzCRZD8CNqOi+
elfUaQ1NIXgKGG/7hWJ4/YTkMCZxLkbPLDrJlnJ9lIKNGLZOj9BExlZ1epv6mwDVqT0sAfaFRvjt
bpUvmnfexSWHSzLt9QeC9fj+XBG06FJJn18L/KkMTQNYwua5sdEKkJ7NO2LWEsHWldIkDnlF8brJ
02J+Eq87xorJ1SLo3HEMLYsQYjeLpMOb6MhMkTTJPoPZjeTbD+LwqbVGaEZNC/1vWMNslh2Jw8Kn
mE2UC8VzAd4u5254xMTsDDxCqvBRP1cFdjKW3JHYG4AUIo93sxVzg2SXivFiLqiQxJNdHnbe9oXD
7NBbZm9LDw/Kzs5LdgOo6E2TsrDTuFLUgr810SaCZcelvUKU1rX5w18t0VyzsbguIZ6RRQV9mRQ5
+Ge9Xj2nVQBUrmWwmDFO68p0vycXTwPQOJmHLz2UopGg6chRn6kRXrnLc7r7KUdoXywX3W/MjRCO
9ScPcEpA/2zi9CApYKOdjrrVLsHfk6yqWwtN1+WNrJvzWYLk2EIsN6R9y7uhGvbFyLLfrz+Ggegu
96kg5WwYCjZAMn0S2UTgb5gl2vwbeXuE5gMDnfdJ01neKyTKY8dnU3A+tlhel+yzpC9TuDMvn6mQ
GKrLTaIl4fPmdqmwS4Zcaf+e+woaSdQOoA19JcBNkpZBuMmcuvnLiUR5IBMFKBXLuVKG91YXcmyp
yaYFyNmLBo4zXHbUZDKZws3X3bCwa1EAwkVofkODCacmKx8ntqK5tQMsfU7AJv7FfTBcV06OQJv7
AIXUwTUCw+KU5ed+D8GNR/cWT1XAwRW0w31/bQvTqLEFwWRbxTrpJkB1XekcDB4NlpDps6+BWrrk
XB3rKtVVXrJhfZJDAkgwMiWzW1D2MTzFAu+2xFnnknOIr2EZbBO9GWWtJDnhRtKqGfI8Xb23je2t
SoXvN0l8NvjXaJgctq9b5wXBwqqxVhBtcuNwVamPYqUbVbQAht+g3OKgqBszUNjga1FSb4g2h3XM
XK5GLr5H9jlWqaxI9ws54GnkRkCcv9+jChcfAcSvEIOZTri3f83rP6RuXoWvfFiYSpPqKg2TbLVJ
ee2CROrHcDskRM6wLdXJPNdm7dg7a6GFSM5nnq3tuJwungu1Dj7ZlquzmC6R+paOhbm8AYuaEFTk
s5IyZUXc6OPnUWdyvHWsCO7cXgOWdk9CKokfeGbaw+lawY4R/U3unM3iNaoHGVs5kjR7ZNVc+A2p
+F/UUDNg/0K5Ed248IpzPNIylNGRYJ0rKdq4v2XNInQnJXcjlS/J1Yc0aC//9jmzCEkawmeP4t1w
z1CuWsPIPoMnDUqbEBo867UN9WyxEG8v+FqV8UhxV5lVPONUKMavRfaJd1zpfNBuPDSGKfoj9KTz
ZIcO/SX202eVZYgGuwAoo2Ru0uYGevrd+pAO/jH9rj/M0RzJpS2Ak0erQNQN5B0tkYy9Z3tONi+U
tE4tM1rC9QS467BsAFG3Tbvl0Jhyu2K5wHb4Vg4Bbm1HtH1eqvdm1AfO0+3iHMyaoXfwacbU1acF
gWv+glXXm5Wcurwq0aMTMrMwSSk1OQOxo7isJqWtn2nImL2ZVKzwVg0p3+MMWm3OHJwBthUQgv8w
Al/kAiqB82xNIQmQuxR3mgrMWgdMis8C8pl0cyZE5tac/1samGPCN9+gvYc1SSv4LRMvKNId0/HO
gXGpCGlToZBIP8Z1uIGm1HwIxpONuDPFGTvxFWX3fELv1bUM1lzDKtRpLsKRLF/HLs+IBn9yp+Ah
Q40pQaQR4KkPVoCzqNnkmiMjYkXbdgrO87UiIuPDaQxt4o8FN/FCsLvQTAT0roqj7cVm6gDNbBwm
8teibE5fegsGWT7OBk3kn79HW78C2911jVXDgbD2m/o1Ns69EPgwEY7u3Uii1E5Ax3dZXXceqieo
mvaVo31l/2YGawBUtVvInqj4awZ2HLP6D6kaz+YsusoqvyTO45VR6DaW3mo0mL7qXPR1RWE1JIZX
mK4nVvtNHPYUT2xi1LyvzepPytOIIswgJAIK38MbER04yg1LwMDBMVbGpST7vMPZQZXUom38KfBe
y20bb0m6jJqI/HLZDl4gExabiLeyQ/W580ItXj+Cedn/6WYtXjyOdtxgX2lUldCcD40qowb6PoIG
iAC1A/crJaG2B1YP1v7QyD5BQFgcLl0/4tC15/ckxNKnsPoxJ0ZOw3zM2sINH5kCA9DOdm9P8X1Z
nHwBJGPW+kJEo1L58VnN8h+7Q2lte+WcUMmr4UEdEhYbzsJS/g3Qd9nqkdUCmF0mm7pzZoJ1fMYe
InTCdDPsA6WLqUolVjblX5dyo9kcl7hvsSHsaOffCpk0NBq+F2zFaL8fjQRTSnUUJhIcc1sO/fjK
u0frFfjpWnLqM1EdFkn7mo1poGC+s/WN1+j3LJ65UGQorCjx1DK9KzWxiecBfyO+nhMqzSDh6pcj
PXX3v4kWA/UsC85Or6asRbkV0TZw2tHXF7TTT6vaqOyif00VaGnfkGzft31N0FX0+3fTv33c1Kzy
MWQ/BR3fmvG5O6zNq0Cd5oOOYRhzV3kWCBs2YMre7l1RQ1nAtsheyTNlYsu1lgfWUyWOIBwwFqOv
v9cdFouL39WUSWAYrbkrS2G3xlqO/TSAOJsXuyMKbrSWXNCab7QYAdf88uT6Y9/xCTtNhs3WDn9y
isZ9eMD6v3vcWpY8QWWmBDA5YR8vsJCPNvz0cdmlbshyU/2+qwDODEXgf3WldAzuyv6iiTxREWPj
RNi5GBdCCf693/nJkVzD6t0yy4IdFpDR5n3mt1R24a909DcnTjSIs4d69JkclCSTl4ZimK83J2Y8
PaV5UAufQ4dYmOYAeFF8UI+VkAtj4zO5iRjpaX7qrGBaqXkOcFDXNWIxdeFQ7OeIsoEbigsT3VIA
2+424PmB8M76RrTeBBOHxEquAMCBk58XRYdCbg5huzgKGR3qNhF5Re4AEaaU2FBOLCfRpy5qIHJK
wr6aW8ljnGYHBY/NnJyS88iMkYrtsy5DWOFt+nMh25PXbXE0BdLWG33GE00nkZ1X4cJSSuxWaNlJ
htMZI3Yhi+aJufQKpf1NvwMu1eU/D434V/61oJvGmYL/4CL3kJXftivL8wugfa6lFUYkvqRd9Yao
3npjA85L+iL4H957VyifNHZLGbDcfNpZnJ/JyS0AvAuSkPExMGT5P/UmgQtQmuhpVVem5z/1L/RY
dVAd7izqa23ZAi7b6ppV969y9JA7To/DEoAoLywd20dltf57me59SwpcB2puOMNKrbJGF3Vr41iR
jl618thsb7JrR5u/TyzHCxnDZ1+dBZJ+GUVo7lDR5eaK8ztMBylaidSiNLBNXILgEm76HDEARZpH
++sjBb0/V0RPJ259We52QrKBFrrs/oB4xCFMNSh7kuvmWwmc4OLuvjS3cF22cAVnOk4GGzzL8uZ4
m7ZY1BqiQMOOWjKjLxK4wXnk9WCnzg4btBltVETiQ350ZCxwxA6sY5zFD66Q4QJNqHiuFg44fHV1
cbym5hd1u+KtF03YyeQiEZiWGYoJSQ2fWJnhlwz/am3B96Xc6II58UXs5gXMopawNtu3zo3XvLgG
ZQiDIcLXjtnLx4HrV/WJjnPhgrmbqNsGGVx1mFVj0rx+6TXsvwdRGnVc5KQOALK96ITQqskmoEC7
75tmgZHkM2++yexgVa4Q8fik/F08atsnUKgaMcbv7oKHlhI/zx1of+B91WNOt9m/NGYDYkbUgU+t
lW7TXg0uMwRIpiVqA2gLc1qhOR0vwAKQA5yA4NIb38WO1dozqztRXn24Fvs5jWrl/ykLBiDcpDcB
m/c9oeJ/QBnc4W+i0HYHt8ntscS/SB0ocdZzBc70Y1xlMrmA0meObJEuQ4DbuZ5R5U+Z2RxdQKKD
j1gd1LbV3lJkl6pVEkGmIGN5pNCeZ8ktwyYH2619JCap7O2dNLwsHu8dQHjAQdldUToR9qUAhQ5V
kboJMX9xZo8MPzC+N34e2EcMM5A/hwQ4oUlxLhPCrNB5wWEp8PBrBpFOagumClS0qlmyJtMpW3HI
eM7iz2OFdyOXQr9PHjjKneF5owxvV7VhM9rh72t7xYXywONWJTNXPgIwazvESNbiyYaA93DqM0kl
fM6Wxb6xWhO2gV5bAwQ0hyeHI2pESFaX5iKDFMZ7okXO4ag8wv2hh//O8qRaRGMUa9qGSOJ+Fm/w
lGocqtWxFZTsmrdYllqzzSnngar5bkEzNcslJ3wUzouTA8RLRX0HOJJDANUESAvcYrxmxz75Nrb8
eBi2KYlHdOmpJdfpY8vXwyqciwnGCfXVmB2P9mZ3wbc+MaONtzWJDufSOdSc6zWAOg+IYfNYSULj
YLcqTdQHmx4fJCmYl+4/toPCv9kFB7ODSrRrxk3DYn/9BEUuvRO0l/phx4PP7vP3J/MjszvOO+4/
3mBNOOshQFEJUMLINrkoVjh3uwFZkKWkVqxNElgFyAent47vzUwO8USB7dLWyyrVT24XgktOOmKa
+Rj2u4ETZVnz4AVqz44ZsEg1bp09lOQeg2E2W1P9lRhFQ3cUt2jHHjEt2wwNJq3DDQ83iJBQRB5r
b2g2c8twxhgOWJkNW6SHPi0lI8kyOQHB6emLXa5F3BtATx+3M6uvg8XjIB66Pdxg756vRsoWCyeY
UwiAZyUZvZ7yM/ortSb4ZxFufr50nppDYcidY7f/8Wq18rap1QrBRFKudGMd85Rf7nnamPZo2KTh
Om3DqZpekEc77yA4wiEfDrVjMg/LaFnn28YwIPQhgp+7W89EgB5q3EATSa7jkDpZmTL5KBZuAmmB
xSFco7LqMiPifJaBgDbuamArtC3qanH7rMA3C/QlkpPApPdEYaYiLExfAIyXRJqPDiiKIvmQKtWu
RPPAYEMrS0sWXajNpFmmq7kELXQGiHfXkUjZ8kRudFUszLdImaTjGMSOsRcO+fjU6QwBY9k+JUjz
IsG9qvqEzCFKKhhOSKwBYUbGZmJEXKSNDi7teB8WE3qvn5n8MUGkZsOUodBamQ33SY7S4PjRuD+h
ukbQMcAkyrDnsQC78kzqqWR4nQa94ZiNG+4HYLFBrwXnRrc1T8Y5yCAn8D4b8LwQDZJBMuSfuZds
rhjBwdyxClJZ8Tqehp0jKu1jtBqbD9jGGW9LjpFE5GRwRoiX5LdWEgDuho7xOIbEhXOgRSgVRI09
h4x6lDCE1XTPJQSIeyW3swUKVuqab+ZAQAjShuJNzJpnHcJNrg+9y5Q5ffYVv6Xoa+c6zKXMg2rd
PUCj2cd4pvxZQL/jAvwdNTiMFg6Z8OJWyoeP7nZxXHvlTVO7irkDslptU2k1he/I7c0pKBaxp4qr
uq9Ui35i6vZLXdgzT8in0oPIfZ84O0VgmPYx0G9G59MnzCwBqaxfYjaalWUdbalhNDfhJiygmVZL
QXU7JRkWqFDZuWXc2yKfZsgGt/xkFSuyAToxtePAss+fxMD0D5rfhj9MUlPd6Yiz23jc/ucmiDuD
2t3hP/sdlBSv3RGFGKXdHMIlYjT/9z4kYkPeEWuLRK0FVvCHAmT8nFboIjN0s84IlFwibJ+cvvYF
lyMqpkmXJTfJPOLG0jMIdbizGSExXuknS96dD94nHqBILMkF/iHfj9av8h6wrFTfL6XTOwLMgXCi
o3gdFZNjFYgpBR45/oXH8A5Oay0Hd8xEkxfxwCI1pAW2dpfxXh1jiIXeyaD+PAjyY9a+xdxFXLIv
rd5SrMuFCTpG0MSO17865T/56PlfALCz/XlyRZ3K6dXct/JufWYS2kKizucF5xc4nNVcREEocspQ
lnuRdkx7r3AWkpnBpp4zTl/av/oHm6AD1T9JCqkOt90J93Z+OUSt0YWm74qlXvtV08l7pKjI49kI
HH5PHM4uoAzHfeBz2iyOzHP7+iJ4YNCCI//Zrm+x0+bi9kDcIYiA1mWYe8IagO5cfJ45F24UbPXJ
JjeldLGTaB+dFa3P6KM2D0sLYHtmnX4+yieNL91SEorQdNqzxjB2PuI7hIxOBwn1Ss2c2+jY+4QQ
yS5E7wTZuhzwcO2Kq1Rm5gW92gjv5wm7B53ip41d4SLCniKYGpfNOQQpnkfUsAboHFwh1RY/iJ71
1g4pZlgpLsXKv46/K5yKz478YVWPBQa8tKRR+N8TUPZ0orsG3HE7qSJ1xkY7i8lGXAhNdvGTIPI2
92D8vsT0aoWqmfst3zdgUUcg3BwxvS3q+oVaAItSvd7qzQuCVl3WwxoK5PCGNQLK/Q4atHDvqGPW
yj2ZCViC0I/NXMawLacZisXZV/B2IUl2TAcWx/kj6rDfCkArOhMDv/u8o3XeAdn9284I+v6nbh/v
WUfqFNqAOJct2Riu8lsn5oaWwblnvEvI3259YSq9YirNqVBdJWa/QtwzJC3isHfbvVOG6xKrflV/
rQbp4DOHIbfQF5HwG+Sifja4NHMj9yU0TSm45ImjzcIQbsK0CgCg42c5WPIzo9xwfSSjqIRYPAIM
ZuMSENSlcTNk03iUOQpPiugBPcZ6nyq1ZRycKJU4LOS5QMTNoEajuVRN3gEHBlZ5iOv34DqiYKYl
M/IVwj6mrFcbnQULKGeeOYjHurL2QworUVqdjWndAHfCb0REhz0vsJT9CrI1N1Lyd6XF7SRbR8MX
4yWruWVXhaxzDkHBbGjAEPppcXa18NTnR7GutDWQHRUBNGfFxOPUC0ktC9kZRuj1BTsrZnFAgYqt
DJyf9vqv8tZgcuJuiCtpU0DyIccqadhbX7kWiP1nPeWHeezB2o3V5cNvoPYEz0SCxBLo4gtyZggn
xt4YiVBrj8lnc2NFAz6yOEuglcbAlsK7Qk2kwHwN/CYjIdhx6NvHLkUPynk2mLVszJGUa45Ta0bJ
0Hl4BcpvmpNmf6hXbwAUnLf7sta6spg3hEBdcrEA7xwY+omUMTP4Bg7fotouQ8/1QiwYdFnX+oFd
U2jyGtAnutTQSw3JerRATNKxODNNWRvrICLrjvGCG+11Lky+iU8t66x9OEFOzkva1FxXcVI/2w4R
nm/A+tk+rEp4QcBjkK69EDdU4diAv2+7fzw3nKoH9dbPFyewrWpCHvg4F+g/Ltmhyq/jcZGsd5oj
F0IgwjnyvIq5FcgwVTlXm1Vonfayd2iih5gO3v0X0b2z8LaMglrikRlX5vUQSy0A3dDZ598QQEG/
eGoayrVv5/vo/GQlaMn6v3QdOQktCmCGPo6cp9ps+QtzGLuR93zzVEw5/3jn+pqawOcozecENCN4
KBVYZjXevceoTKBuACxCnsygkEsUgRTwIGAAmzBG9wIdwFPtBQDW7yypGeBL/l1XPYXtaEII+gyI
hUpDufsUgQmDmIz4T07c2rOck/X+x6fFJ2ELDlmGsTublt4wM29SbONRwLihV1EOZZujRQ4Da0cv
xKq0Yn8FwdWmxMf9OLvHqQVSQW0+QEfPltcH2upkqrnF97wmiQyqK7SYb+l3kv2/t5WD83EYjpvg
5cbU0UE+FBODoYeTEiY1acy09MfElg/HZucCVNqS5Zf5TmedSd+iNFJb3OfKUUPOMEwYrCUMK+cx
6G6uiFPVPeH3pAxMrGJ0znIJoVLgHVnxQbqIuxcfs2RBSARAbojmX+E+muFEEnAskp+BkAXZ8t3K
Ypg30MYoWeMkWhuYRhGtaxnjEWr0tMZKXC0eXYgweqNMsWgZrxjNckhohhWvjTpWRpUhECSsoSch
MT4O/y2P2rQbZfoTUFCgfgZXgG4vGDZ/X1o5piBPOgisfiqCB8wMgAbXhRt/LkEALxQ6r6SuRxYU
AbLjWqLz2JISy9PvOox1r8YtKMOJ0/NnNNqdNRr74vPOB3Vvh0mAjtrQEglhqeiIvMUwECT7Xbbx
IMGthrt+I4BIdamNsxVtuq9OwCnJ35c9Y/Svtuq4FuMMaaoJZEnc1wVRVeDTAqKW9iX0x2vKQWNc
3wW9MtVnQp5vv9QYWz/LKrmD0fTbmTka1sKDchyZaHoVevilj5Vn0S275dkZWZbplZaLOMA0IJX4
7nrL6gVauO9r8bp/I1JvMHjHQgm/XuzBx796fucJKHun8wWN5rVSu1XZE0znshJsDZ0q5CVhNm3D
VUkZ0w35F9en13PMqE+I3kj/Vw1l/IA3cEDOMLmMefFK7Q3cxoz4qjHYlP6G+StqSl32h+19hWXG
gBWPIkBG+iyTlG1h8MTyQObQSEeq3n1wuHyBvxlRrbN4K2SXhh9vFFIexQjU+oLLzsukRggBQg+X
Hckn0ZxxA0UWscwh7YfJCPJ9g9bNXa8boWoAI5WN+JXfg6w19uNcnNsYwWuy4bFs559CeykO+0dn
3au8zyyZW9rVWXalZN5K8I+bxmBNvydDo3OYZsKX0oCPz5BZ/PJi0WVAlmE8Y+IFGIBLII5yFsMZ
WaAroqwwcl+MD3iEoZ+7D6yXTGMpbphr1+gNaXMtec3DIA8Cy8rt0xE58hWJ4mM/JUCqiLY0meFI
h9j5w5MElgN+zjrEHH3FO2PqzV7prSPPALsI79dp4eY0vcelQb/mHhlTqfAEbOpVdzO0omzDWPu8
JXzLLE5Vy6H08T3o+fyDVAnHOzTUWGXBzR/1xDFfrKRyZrU0fdvOUrZWMyjeXNW7poUAtCMCddXd
RaI+7wk1dB4z2VlgLTaP4GwewAuf2zozTUAyjhipH537FrCJ5uJh34iJTegsrA0U7mBzVlH9IIcn
jBb5vlbi2kOGeR5MqgkEH3asGq4mCfn6fG87Du97zDGW2/otE2Ha5dNAgMvQirTMcba5/JX3v5Af
4MCJS5k+NeFNmqhqaUNjg7QPR4bbBFIkClAeGNC3cnntGPCydR+cxAZ6bfbI4s15myfJQW/7zwQ6
aOHa2tOyocSPQ2RUYHUx5tOEr8YTjxAWmw1hK1Pa7NhOySZWnW6cJ6WuA8ECuWHwTDHDNeSzJ7p+
iKfJMSHrTJZfO9e8dQwzYAVprW8dsvMaCYHDTwlx0iHQgO3ny1EGO731O3V9E69nqSgSGfdGy9Eg
SXIF6JodilFH8TwYCMb0KGULCh9fHudLlhuRUyofJiiHKG8R5MRTn/6UoJzzAnHWeuhBqxAQ36f7
vXwDi3tuvG0dj/mh3hJXcwcaPMTF8WJkXj8hXzXoS4Db+L9cBZiKFQcTKPAwbkj0+Lpskw6z3RPL
aD0QFMd8iwtWZLNP/fNJY2f9hv/3XqDweXl0kcl/j8xIRsMFPGdWq7t+EyOJ4wAJh7ZT8U++7yzw
ZIwOIhjvL8MNKz5ThhbanHoHXTZeKRqw5r1KaXLLKGutkMc5EJHvgeRYnKAyAmpHjt538AiRWIgq
o99KJWgzlvjKIWQWVMl0FIZkFQoymb7UKA9BXHS+ZvR0oXLvTk7RhaTcdRSkjGwRR+VsVlLa/AYz
7DJfYgLMFkzPAeNv9hdIKBWQm18dThMd9+6oHF09+iL22sQXLB7LC70StiDm/ouQ6dpo4fFsg94U
5KVfAYZ8fYKmJQuFA+s/2M5872SjD8yeExJ9J62kj4q8olNfCKMZ361wxUloPaEwzpGR7oIbwaH4
Au4E39PpFAF3RUss5W45WsWLHeLok+WoIqG98jiDUIr3fCJDZJC/5rZu8t7V0/hHptYCYxUPwDxT
axPB6GLRr/FSOzbgI6FfYrbYGaXEtOqGN/x8ZIejT7Hp546V46Xj7SEY8/3pPDRQHduba/0OkkTC
sm0CHWfwbv2g+fTQLgPCE7T0SMJawkcyfMGp6iLR3cfkB/zYxiEEz1eDypzhKB9E0Q5Fi+EoJXto
ae2Q3fGcG8goMd4RrGg7pw/7FA2OX95G2dWh1G/BhUUDRC/gg473YtXzJk83vmA6mXUf2AhICIZn
SASsPNm23tIpgT61y2tQXO1fDFtTxDb5Fi7D65ZBs82QIsumMIRhtTQ1z77D3Gtq18gOhzdQ1dt/
drOMttJTCK+EqlcqQHGBqTU42fYmDT8YWBVCqnkTk8u7O7CZ8QpxfVddZEjdAA2XMgixtLFcxbrb
VNLV5lcZjZZCL72xM2i8KY5Sd8j22O+oJf6+AbPuAjprK+ywFzmFJT1DDIQQIY5mBQ8LlXnlxj9B
4bdk72JnYvd2CFqQt0j+Hf/UhFoWWuvBdS4n1LrIn9ZTJ46UhN2veaSiGaazsQ7vInPVEP2DO9m6
Lhvs3ZjtYuE468LLwuzFiaNq8ITl0qbJylFZGR9yPDi4ffMK80po9N9YMVHzOPqN9TnGAVS2vUm8
PXo9E9An8Oy7zPOipJqHM8bDpcSGXzBe74e6NbemDKHaybptrDpWdOyephuqiNcB+Mqw3osWI55p
IVgYtJjLCk56jL50O4Jk3TZMFpP4oYaPKyUlxmcpGPIAjAC8gSSNXIWIODyF9QXteE53I3+pRMRM
haxfrDnXZ2k4TMt0e+bDiosd6oqNB5iXdkChdwdcO9UuvVrP5vgAxRZWdUqWkIWuQHiOhsrZ6EKa
p6Qpj8ngSnEtM3pfV/L6FJ9lhAU0119XbEAuCq+fIUnFFe1L7+SQAVBa8l8hq3mQpW9gd9slwdyq
liohSRFP3vAnMCcUYcPWE0GwYm5SxQZbgytyX3R8+OnM/k4XQlfIg20+Mm3x3czPfXKploR8kj3u
DaMnWIqqj57PFiWZRNfOKOjfdR2w+C347+fK8DUAiil1Si0BpzRPlDYT7n3LyUjbrPctrxdpfYMR
bqwqeqnKy3q5CLP2yC4azMyDLysuknoN19HoZzNkdkHEl1QUikEGZW6xoAlm4VyTgKqE1Ej3Alws
DUYmtQ+BMl5zBJ0P1XmGWpZaGZsZEgLEuplW37bdbLesKUWCYOY9FYmkvWXk7VqFQBmBTgSyQRJP
Tc2mesJznND+UIwfp+YBFlR/5F6vicdoM2KUGxV6omfq/4qIqi/eXqNMnLgFCOLGjDc7JV7AA08I
fs6/q3vBxo2Z+fQ1WZytBg6m9S57KNpJNR6h7sYbOtroyMcNif6S5IQ87z6TGB49ZH5Z5zoDkLpC
diFj1cqbyOLkxY5elr2V9h1tJTZ9Dl2eTyyVSUAtLQETYp0PKtVvHy0FHDQ1SZEnrLqQFXB+pDHp
l4D0us4/EUa3wsYtQP/PDQd2F+H9uBLFef1W/31vxWsvUrbhBBrbCG+iL3bTjGSV/yhMnxp6aOrl
Q45erBS9W4StmmVvAIXZMbyoq3i0hCL3G56AUXXyJrqNqiiJOLVEe45QT2WldkqY+YPTp0hdJw1f
CDGb/NAKenUkzdE9H+Z0TkiIQ/Ph3JbGH/PtZk+IS93eG3t6bVX2Mf5LMt0jFeT8HaxygUUVPoTE
3n2TBBA12a8tWTT/S9qtwb6W9Yy42HtO8/FcH087+HcP1Nm6qzNIeDxvWfrA42ebnISeiyVLmeRq
ppUb8SZN859CQfbAaoSi9j5rWFj4xIuHlcZzBSRyc08iQlTSMCrd3ufo9ylBgQkSkmg4mj6smqCd
9RoPjoXqtEuLpF8PK3kEeJJ40td2/scx2J/OIJaH7UCW0E/nVQyLXEZ5puG/bgLvXTzlTf7ZJLAs
6kNOzsHEWwd/CYfhzfeOun4vNx36o7h72IXz9MYv1MyUgB1OMbwUKfEx77lUYGH/c9okqTgc9QPl
NEwdvbcjp6n5EWi9BmlIVtZrilFVHsWpnOFkggnXb6FtMtXm3rrXZ946dfUfrjAqoMgZISDnFHiT
Pc535BaDT+1HaGo0cQ3dXrwmr1bUDF2bQNUQRKB6srGTkBz+3h/++4XP4JLmO76c9lyrypb1L8NH
GMne3k72X9r/LlDh4ZmTqNAFZND4kTqDH6jNnqXwDnZJybKD8wktxTUuQyLgXLa/GxzSLE4BzHHR
IVr5eNrKciu8X4r2rsD3xa4gJLJoAmcjjg8eWTg7G394sZ8dGO5Wa5MB3s7UmUNfQg70jYnyOPu9
nSzBQ8Yj4Brzsicdj498ap/5JIii9kZyaM3PoWNZK7eJfCyEBA3uf3HjOR499/0yZOFkGBEngfFv
SdWuQooxTq/X2cf5kx3cv8WkCTvdWL4FTp47fzHdBGRojaUvKd6mtPTyJRnU8OuDA09Ue0aAE319
LHCzCiJkciSdRJYGxw8ZNJyLE9Dl2ptDD/jieCMmzmw0KcXEjPyk+5StyADT2ezWk1p3P4KZheEM
4AnED6FeN4UYXdLGqdhal+vuLaqsmr/47V1Jq8GblO6NId180T0oixSNoPKYQYMNSWGfcJSHkamc
Q0dMMx/3a2J0lbqcAj4DlEH1781K/qLqQtXMaaj9kpdJ5ugiIKJwB2LSxtBu4nh7DYaGKyzBu2bU
Bw2jVs17Y4ArCKVQSShYhAvD4sHdwUrwNo+H5GktTw67O2jHXs0B93lCI6WFAsufsr8WVZQI3MwP
/FTMLNVULcvJbkyZIIk3t/WDUvRoa4LyWVBfv81lDO2zODrk6Aw5VKvHKOBb1tdnfuKqQRoPUfwy
zZJA/9es4/BLE5tzqSYlHKdonHC8twseyiYroD/1wtUpk2NM0mVK7ALT7utesaWWTkqBKvP7vc1b
vxc3QEadKL/IsaV95149j8TfrkmDoYo77AdyKzIs8WLqHI/p7hlv2j+ih1K2K20GdXn0HsnmBRXB
tlu8p5xwC3xC/s6Ik5lXdW+nljjghjxekhhrd+RZmG64HdgSUOZPCulY2M76UYIPKAymKblLxaYP
ow09Yik7I5DzpYXOaNeAM0CRaq29ULMsbexeDQQB20sGaizNwEF5j5g6iLlFzRgkKjsmUCKR4jlx
2mX8ESue+G9mpt5gLYwINPo4OJsYdlzd/smLgmxzkEscus7V1dgyLnAYO7DhqqlXOPizft0FI9Z6
kEZzB8ThndcgZqZOSx4iYz9UystWmZIz2tL5qVc414jYm0x7Q2IS4Fr8CgWtM2AFacpfN5D+JIWV
GVDeTa9t3yJ3Tfm+9MhAbw4if1Yx0L10a8c8hwam+2GsyKPVn0CGf3m2dEcB7Y9TzOHesB40eTnM
LWOTZrh9ZSOcDTmLS/UqrBXAkWRQAMOMA0G+g68UFahmJoA3gB3KZXEAIQtZqOEVH8Xs++Ozfhg9
J5QOANlm53BlcaUfE1pGLa5+QPW59Ps4YKYIWYjyp9jBTdtWBSXjuNZClxl+Yc5qAPtLdIXWpNL8
VxnzZW7cQlU8+sULW6mPiDsxnzNGGKWQsicXtWi0ixRuZYbIZCZiITY3ClfXOW3EAqWBTU3OOhHI
v8CNak3ONYO46ZLFuO1tavhmpLkMc9/w6fEeAltE8SNOeZWbgNeQtcHhKwSv7Av8nfjcOeRyOYxM
7/GTW+KBdKJdioJQ8rtqziQN0tOsfULQlAomBIIbvm/pb1Vt2PoCNm0OboeQhaeAtbCzw/xyN7IY
x3DvnxRvuj75AyQaXxOBxxCimw6jcft51HqSohTzRqq+wagkC8XKRJTCfPfnZkxdjj+hVFV6M2kH
twO5dmNkMoRYZeNTq0y30alcbzu7moVcL9OcnFvqXzq6nBxPnnBJegUqhhiXTIh0qDTFBw07NIOT
k1YFpW7Co+a3IOC+AF+5aDLonuSGM3wyXrtmtWxz8hZnnPTN0xPfabZq0UjaF9h6zNIfUYWGHnJf
hYC3VCWLCVtP6b72LYQ+emSW/WVhTXCZWKac+dEyhOHLdWKWN56/6ZU/Sjl59k/Bh+t1epSPFjsn
yZs9oMG2ja39k1nDryIspv9htZiGCcJSiEXwzEGxQqNJCKMo0TKpxe7L1Ly/9YZ3nHlA+d2CfBSQ
4t+O/S0kcLjPkCU+aDaSn1k1n8MROwHjs7GnmGsucUNCz115FNL4bG+6ZEHVfbQXL96ZJXq6EVQa
8X0HoCOGAyxSFhiQknDwJm3EKT80lAeEEg8qoQGyEs0E98+DDzRQ0peDuWsqpq4jqTKZLwc7l+JY
/0bbckuvZbWkj76Q31fBBLRY0eJsI+cHsRZeTsRXen0RMBGQ907IQPrG9Dvi0er7aK45T/2CQfMb
QdL9x4axele8lEIRtl3LgtSDhCTbGB7Y8TtCxqvyzer2C7Tom/2xRZo25bz/KA0GbGYbJ9/XToe9
VFSl/FcryVlO/K/UTs7gYS7Yzx3VLeQ9gOrGwn8SeVCO/DD7BrAUtwbvGml2iGCpRRaRboIu0Mxf
37xOVWQ61yvU/BKnhg+WYt1079iz2xekGqK2kmwZUXeiNPKgwaapM9+PXt0XgnqRsC+hDLqgvoZf
km76hbLFSU8Ouh6yhnA9Ey7D3/Sc6VZ8OidPhdZLnXH7f3Aqo2BIKLKO6KgJHOLOEr7I2eEhY8yB
5SlRjlXcpG1b5S8hogF8rvx7dhV9wMzdrtXRFj9NkW5shuijJs52FpLFBEWC3ufo/48osQwW+nEf
YniQ+XK6zxBlG9xIB/CD8qxdFCCreXmyVw+BoQYqNkXCVg3RZ3z9zFn5pUtrWcbZpPibd8e6pn++
YhQURL5211iZ0+VOlgexe5bZ05pwzu+64wpaf3ivspEPo/AcWR3/3IYGWtvF3gRZJMJrEiCfCx0g
F9bOTkC6jZtGy985XzX8dP3RRa7qET5+BIMG6menQJd+2/BGm1EK1WRsaqtL7qOX2GyLTyBv9I/J
4VL7vX+msR8i7LxMdu2KWwm6JGw18t+SUpdA3ww5fho4xDwfOY2GshOR2ZNxiP07zzphBxjbJb6H
bCykvb6yR0/LaDR4x1plmfzerj87Bw/nrTRhAnV0V0mC1pmGhnEnwmaJnv0x32IxKs2jsPR/R3gh
GO3k4QJrioFEK8E6MRh9anWS5DgWgjV5y92Mjw2NZ2wHtIHBY7GIWkxEAZPZFYFEg5u9IbPynDxx
YKzqNvMZWR9EHBoP5mmubvt91JvWQ6iMkh6UZMOvOSAghGFwWPG8FL4IhwK7+eBzqLguRSwSiUbU
wpblm0Rolg0/3CKZGuV7Xkj+/1nSGwpvOcNLTsDKm/KL8TDcOvzGdF8afcpcqkVdR40dOwQzODa8
f7EVURLGnv6LVBQ5jUbf2CKggCUrGWCqbgzR8oxYvdOC+T+5GSVUnp9EGR1ErgDIC6PIS3IpGp7L
CGkfKvIKW7VxDPxxF3AB5tPdjqjmbJ5IfF1A6wI0jZdXxtzLY4i6ubpGvmZ4c8hC/xqkGXJ/6dwR
jHASVIrSGhuEuS+cjo0Nn61REIZYD4KTxxgiNB3MRiDEbgtlbOZVaM+Xu6W4K2emGHDOuT13jnzx
crhE3Kxm39k+hrr3wV1ZoCfuJKAbWwP8pQSgw156P2jf3gaW5IXk55tvN0f6MydhU1UHrLHm9qYL
uu3PL5XMozSDpINcI5QsySnfla3Zwv38N1FnFV/Wi3RVbmKXev+U1gcGNcIM2YENEFwv50c3BSJW
MCDxvOl7HucnAebFdM36mSgKmYbSHoqf+feDiOFbWdSvnavOO/P/ES2OC0sbbg3A7DTko7qZ4dki
fTuKtRphW7CDqMatD11HJ2EiwFkiGS7vKcquPJ3x2t1Bj9s7RUZx8KDieBZl6VIzhmzrl6YgOnjx
OVR9TqD7blyrT77G1EwT67ghNXlDUaj99xYX2rD2XPWtHvikxA40Zt7gCqSSWdYnysZKraA0eC1V
nmZnkfbqa47cIUSCZwu52X/hwgMdJSf61UkGMI2DWFyiWvB4CBdt4F3k0A/xRukQqvY9FM92833Z
tFm7/lzv/C8VOAKMECg+Ormgt4UKh/SiDx7MIVpt8FBtpBFs5eDNOx13kU2nWiz/eXy5WRbFBFQE
tBE+tShVMjacR8rS/j4peyc6+v+XyEWFFt5CLw9DIsbxBQdCBG+8eckid9iFhDtyKoEnt1EaGjr9
tC9FmD7jJTZOMv1fcut3bD1wgPGvywe9D6U1eGhZRdOx2TkwbOIlTg5ZYZZwMT5JiqRga4SqxSTx
TwDC4eaYzRMxwwcy5woUqk2jbACj7atDrb1XmdECgztkOrvQrAlBEC8e+y0JdvmoWVr6R0u1zND9
qWyKeb2foQUX3msJsSpZzB9XZEkkIrgc8cedmwKADbiHRRbjDB7ugmtxV8aoCDkGV+ZzkoYu8yJL
dI+Qto54wSuWkuvompiOnVEIx/ebBbL41Vns3Ibf5cGf4cICtMwaFumKor4QUw7/JDUDCJ8LjYB1
h/s0q1U7EFaELCLt/aBuuIufB+ifJy19NUFGFCwn+rB7Z9wcMNom722cfJeKL/g9+K/hO+2EZv4v
nwVdGvQvUzFJG+gbtV1sdUjqLJz43DXMtwkQnLbDicTefiitwXDwQUArIYJSSHVvwaOCoKgAi43Q
H+IDUFi1OW5jBad4XsGc5zvqHPFgthyDJCrMfeApyEaXP9qXlhFqEgBI+ixux0LzQSrdr/TE3C4k
AcHU2233zW2Ai+99FKDLdFcng6429w/dX9fP01Axj0i77L2dGHgTaCjMLh0XxBgMZS4Cz+UhIDAx
nKUR3TIpK/Da2PjwPHqLqXlWyTWcFJ3YRcm0qFgr8Uv8n3+rt/crhVIkPPAxKOXlinIOKJUl5PFm
j96mD9vMM9uoWOyFk4j8SwSYqSWXgsDyCDfXYfaFBGfEqDVmcYC9FsWII5bZnjlUjCuSD/EM2oIb
7wW7l3SIiFkKlDfu1dAkTyPOKmpoV6UdDETlJNOPJabCH3f3aG182OF1C1rOU8zSjGbvkGDRYTkp
qQGnR8/R8Y2oTo/HbmhtPkEugba7axU71R6n56c3bOup3owO4UPs0i6j54G7gcnj0NEuNvtUkAmA
WKldYdiHYHXy6J0+CEMQPdv6X/FAvfeJKOx9NdfjuV2WK/dU/h8WSx/HO+XDd0Ui+IMwQE5yn88W
dDQBhD6UsRk1cF7tHgLeLrlGLrFILVXEOG5o3cbCu04oSPT5m5HjFWdvxhtsIeX3uzn6I+vkYK0L
qlyFA5zB0aTYQd3qZGWZinBOUBFYPT2O4awCxMbQhsY0RCKaP2TunEcnqvBJMAXnAW+eVtILwjtR
7wkAAvxVT/nBQ29BB11ZCcLHEJdRYLwcQrYwk+6TDqKwm0iUDjOclNLLYsuontSCU6AbRF0Zse0J
bW8mDiNVBdBkaA9qqEBwz1knYoPiRGJbIHEHWVaJIMyF9nOYQYKuIvU16TSynVQ6xDVAg4CzcK2i
leDne3GeC5un4SIyIZlycIU9zM+xgPA1m7CziH04Dm5egM3Y2nPjAx92wHr1UxMyOuuO/w1otZtY
tPx2i8AANOE8Hh8FRMOf570VOvY6D6xWWl7Y0a0oYBap3UejNZXnUY/EUridtewLx1O0VTHJ7P1P
EuxO7lJWObY5/EpAWyoyblE0cHaMYZyi6Ug7XBeYIOQKI6611+zoeT/OcR0Q1UIJ2Kw+w3c/q2RB
qskjTpKLnPWJUMruQN6Llr6axOQhqvZ4DaUUnX/ieYynDe6Xnn7HDCrf7R2f04lO3BtRTfKpj9bV
OuRAYMUvU+E/qrB08cJSzVEncq7s78/UhJRJmOSkcxx4r9FgNSEreok/daSwAVoY0iCKEY5RqorC
FptG4eqsG962gqURbpT2+SGoFgPQ4pKmb1XJTKRLQgWnpz3SjdNzOyytxzkFQHNnYUoO1+jmhQvz
lGME3yQR4jNpFdW+aCGzfuVFDOeYRoqtEwk7z1cDLMSCrAwO6ykIS7Bpat0Sdtwz9L61/YQw8BeG
ZeBwiVF26qInSbD40Ol21wP05eeKm7a25wUbgwl0SO6QvG2Q3VXKjwPvK/m0ja6Fx1ZsabwirAXD
ZMIY4Ym++F7IFaDI6ozDZR+Gz3HHGPU+jLFgZ2p/dZk/qjHE3LDOT+3U1+Bg+YIzAvw5vNx8HX56
GmuMAYqO+T6nqCsHQvWmqE3dxGshwz1WzWcdix4qVmNkgvbaJhFQhS2kDtxXbGG8IlipDhg5PyYH
9sAq8YzO1kKo0CvozdN+jLcHXZtsONjwKEh9NalcPhQIg6lyRay7X+hypLUWs4aEMCi8bk8DVNl0
7kUHa0jREb+D7sf/Uyzd0qdvRNHUGsTB9vHIHw+STGCpSENTeW8qC5d4vr0VU7pjzT58rAA02A4H
ORuAy9NrPFFYTeB67B8cgIhaxGN3Bp6+pWGfVKW2MtJurIbmSqCVjHbGQEhUOBqkCaTRBMqTtgvo
9L38vy3or8G69L9EDfKKXoF4S/FKPGtXNkY8YeUELEN05YCy2iLd0UKiVa5zs+SAf0xVNnTYbIGt
qNXgXsYgmBXNyleDe9UAXGlIJOVP1r/1h5gtt6RBtKxUpsZly/3XIbYtRvx9yvWVuZu/IosXQSJX
oDIJUhYRD8geS//fCzzLVWnEdkUVz5zOeDinoxTkBrXWrmrSPpkGVLGhAzEr3xFmUZRnGR4tqyBY
1doO8OR91GfjJbmFV4tJLqvAhlGZELpnxUuTJp+CHW2UqzjGiG9YQ215/C+6ip0qa9BRwdiKYaog
eA375PAdelBnDqpq8nVbTSdPgBruLhMQLsoujTE6+1Cwc9nZw4BTlFns2So9lDjqs7Y161aeiiDa
Cl46PPzvGlo6/GpZYNfBdtA2lfYve3PxgH0E3GYTO22JR4TJqE47rxT2uLSmurTJGcKoGP8Pgkjd
Wa7EUqGcCPCKGh4eTsWicdYENImWz0tU5sgj3g/7GOV2WBc1OZNDekxcT+0EuXIUso/rUB0Tgt66
M+9UIm3ntzyS7YMwb6WH0Z/8OSRKBHouVHVsjPy8Cp5ka08ZKgmXCXjsxZpCbu0K5f/MfkBUWDF4
rKKCn3dqm2L0XDvYkCmNhC5fvwQQnzj/Wu2HsVxHdykjEoDCKKBgbBIOXSEXBiutnI+kGe68jWiK
oYv1Bcp/v/MVQK3wZwVLMXj47/fpCW6CvF2wbeA6kdWvJEwHFqa5H6ShxEwKmIQzRgZdH9HexhHT
zsk+eSzaQM30B42Gt016fmbtcFG0U9z5xWzOvlYdoznC3zlKNOZK4UC9O4kPi0wI1hRIvSSbaRfJ
w/gex9fiCj/RzODkjL3PDvVNfzDboitk9B7qyrOy01hbGC1aB0cEThJ3BcgB9zv1xGu+/6YlDV+R
oa9cZkhJ1viC4EmlB3H3CGho4orszLEPNx5VsZw5SQ+hjBJBGQcucRsVIqNTrQiMv/4VTEjGUKAb
XIpsFreWifxLWPM7Q8IoUX7wADA4aoZJ+p6GYlvAaQee0P17aoSHGFzHW/eTbE6HS06E8DDUaABt
NJ20G/6IPYdqgGLdU4kxJnv3Tt1I1oIgre1CHckuAxcNvrgjvPIFwN4/0AG/PR0zzvcMwdIkDNdM
6b5iMnaIqFsz3ssMUxJRu4AZIKjeMqU23fW+yKqq93s6rvlUsT9f6yzuUOnHl+02huFMQORYBx1m
fJQt3366agyyZmY+prKP3xL291CAWO3rJ9OcjrO5D7sKT0j814bdgbiMsB9mgZKcJi9mJWqaJ7MO
Zkv6L1Elpy9v5zY8qglIYeVYtC1dhCvV7ayaZQOW2963OHYRwv2wVXlJHVted3Iaa0k6yWk3jdEd
82ahjHJqErRiyW+TRHLXh5It+VKAkCgxvBxYtfxYrF85leswRE2iFRnrzQ9ORmjkWwqtYY9gMYyI
vi6O8EI69ye2218f+X6HOmoCe74jziKpfUR8cWsI+bnnhI2ogg2K/bgPoLZv6YWBO1JKkefc+yxa
632jNTZt51CzFRg0y7vd0D12TO44rpcX2AOFUFYeWyDI6qhoIs9eXpZLAoQ0txtkhjvwQkPnZfCu
ieSizv4xPGYG2AoQM4WHudoxSmE6/b5hKlQv2MMLXSSrA8QpcnzJv/HN4hR3imvgD4ztFmyzxdcb
la97dLjjuTc2mgDHlu7yJfAk6pZRzgNTgncWrEsfLifUHQ0me4CpSuktcJf0Yob51YuSZrl84v8k
1EjPqIW/Mizlrt0qTr2UsqRf6a2RfOb+NyS5QX0shAX8Fa2PD6xhTxipKmvzyK6q6VjjrWS3Vj97
s98JOu3RWvLt2CQlAC4op03oh5iX7UcliTDGEVP9uXm7x0H7yh6tTyp4wW08ccHa9vCHS2OyK6l1
YrLGdasjnOgt5kl2NF/FjpqbXv4ZzuHh4yrrfUQf6vkXE6rFyigzVbCurXqyktlnYl38itp4qJ8S
NHx9ZKEH63f+WvaJgYVEWUJ6qRt7sijdWFPHzsw0cOXSdHe16jW6HEn4fRTtkJoZB/Mm9x5Y1o49
0413CFYXytrLH4ksExPy/nzsu2LSud3I0/IEu0CtcDlKz3NzuxdZA1XC8PzCgl2gxEysMfea7GaT
75oIih4axFz+JX+vCE5oPfnUIINnHgBRjbTht0ZRLD38OQ/RPbsG6DzAL3lgLLFrlxKq2so9H8ZK
xAN+7aDA+20TvhrCzIg+mpceAW/WtBoi/DW9AfnKqy+ip3U4gJXp1dRrxY7ZKC9aWhrojk4kQvj4
IfOEp3spqyP6M/Y7XTqLr2kGMmRQaXJ3ind5jgBzyn3HGy4bSlUN2ZORWKHeFcxxOBvTP3q8yISf
HHlp5sfMhCNCloAuV1+56oc6NvUohjXl75kwTG8bHA5hUITATM5llffUPu8GdaE3VeFdFwcUC3We
xLg0yDhAyKtZ5fAWhWwhbR3crtYeWymOlO7xWEXmL7rbH8bbHY3rsG3vAEISMx5Bpqt6RZ4FHHYE
mRkLEJmTys+Usu1tSIpcfNm6vqa2ymoJC/4bAxsQ7jeVQftGEtUK8aecVE49UZqDmJuOp/GvHMSA
6TK0vIOhr45Lp5yfdtogH2r7J2zuex0E4nBXqeLmoo4UTg7PYzGf5Q1t7WMhpQR65JdbW46a+sBc
uCtYW9yXgY+pnp5jo0Z1skSk2xGiJGZNm213ABfhlPNeL22pl06ODpp/df+NX4+ZebEDCNpvR6lB
d9EFF6Tv5hGevEd2sY9c3+AIrciUmolE+UbPmryOQaNPJJEi9VN9UcYBGLo5RwBaEO54pBV7dqVC
SbNO2JlpTHZ/7/Q2+cLd7mLd5rVTF9TIraPkXLIxAqCPN9lbsBJ0jTPzJp1sGiA0JjxNd6Sv+pP2
U+QfhrFXohXM+Gn5aH16o2YsZeSmtn3K3wwfjZ+3amDrnChMPENRW2GQpjbGljup7ZNEEwae36+2
dBHUuShZWhoxn7SZFBOv91DWC+qMUzoamv5tav59aqxkLplDW59wVghitbG+90S3zIxLIe+RMpNH
vcRoJlkejiR6Me/uYv2ULerFybIcIT4NR2dk/5m0aLubhe3FfMFfx0622Q+Sg/kgUGzC0RMRzmw+
l9Jm7xIVRVS6pGyIq3PcZR07I7U5BQbikgwCykNz67Wf15bTswirhwX+ufqp1Pp8WCgx+e42rNxW
x3bPc6OMvHeyzTkq18WYArF/hkPEsNGvIBellDkoxLeDVwkr+7CZEUxs7VkhdVv7zDTmr7u3P8Sg
7s8PObWq3fYIjGZD394DBFR7NZUZRT2G0vi0Wsc3tXecS2AhWYR9y9MTI67MF6lmkNHlqDASS8/4
9H0W7AMe6iZYljd9kh2fxhVz+LQg7ss5IyBBHpEFIrLyYZDNX0RCX1So3h2u/Ae/U5478SIT1Nwx
hdej25J2DlB/IcvlFlDxAo7XQ8g6/ZmMvVEeTrAApOe/tBJuHmksTRak1oAIkB2SbjduhHIo8JIm
yKVMvivx1d5ES0/qchzOizbx79Ltk9Ak90M35lqOEar4kg2lBXElLPsRNrO80Wrmcx/DpkhKk451
QAXg5pZLa/TbfN3Gz8RBdv39nC+cNpRzYSU7xw6FBvmy2pfWMV3yN8w8bFEDPmAiJ0OGRtGgCwkC
9WMt8Ul4bXBzVl30kuMC0wJeoQt13kE5zYPaLUKlWryres3qqY5qjkURCKuGDBwlH5symdx5YEK1
+V7l1SsLGEXSQKpIuRS4PTkzyxAGaWqO11g+tHDFYPTq/K5pcVja61EkYFNUd8DrNJogdtr7VWUL
gpeIrTgdEY2j6BFg83n6/K7MwFAbsWEWX6e6GR49AJ7jBSlIPRdQ2IJ0SoR7IPtJOMhp7irOG58s
O1oSN0RcE9HVUxFhDx5yUYYXObzE1MBZ/CIWn6rDLtiHMaWaIeslFPMRD7zmfJYDKg8MikMaZYFr
xa3PV2voml/lrbgh1XphnjofQnzXgN0R0aZDOKBJaeuSWXdISmYNKIzANLJugHMp67xsVzFV1S/T
rqDzs7xJ1xrPWGmKKiHXSb1IT2+Rekxb65Wv1k8D5mbOonyD1UAOQ3zeBhGnIDyd+mR98V1rL6AM
WK0s9h2H21XfjFtdMjWV28NF6Sr9giv7fV9H/9LfInJiQYyIS81XidnpdZ6r2P1LYR1pIfroLcRF
vh160SqW7KoNWmgTkpEkNaXZURGBbGYiNJRU2U5KqOX9yyZ9EgIxAGvnjPVI0uoMDep9rk8yWrwY
2AvgXb9NImFvxW6qp+H9E6HacjGZdvFYTPD+IosPhk3pyIr7PmGAxoeJET28Q7PqwZQq2yTkPrR8
ic1KcvwQw28ovPe3FNS6pdPa9MUruSSQt7o6KM6sMFrcewg1xrlVlPRDPvWabh4rshUxRJKxsn6S
7++VuXyxAMWbktKg5u+HHWP6uqPUoQu00jgD0VoRt5UMM+Oh2ZHvSCVOWxTYg5B/6kD/J+U+mJ6x
Jz4XPkOJxn7vw6bJ3OJdC+/HdZTuR7lnka/mWhKYAdQqJSw4No22JaXJyjhPD7jDCobMYhDWJX7z
twHiQ9pTJ1iqfY8co8LUOyyODki2O7tiEd3BUNNhiTYy43YGiZEdbpio+MDfELYz6crRyH7HycOI
tEwfbRCqza3k4cV2gBPoyHNAy+0BSbug8knhry1vRWdf8kbHE0k6G22H2YiLCm/IzM2Bd53Cr9OU
Fg0QfEWdvXsK1ppYTr/hrHPPJT6uhw+9hyMPZGJzPXLfEnQTQA0sdRYT0LjTDS0vVtppt9cYm0+Q
5wmOXDcMW+dhwbtserk0bUa0nOCgYJtUJEJktq4DiDPKethOQf/vjWyWB9oP+K4MFFewstSJECs7
Qp+lZzty5WztHG+Wm0ONSgdYc3x9s3DMFXxrChnsSh1qzk1nk6+dfyEXShDdzWcp/TrZ06k8qH0U
fDxLZD3ZzbLpYfjSx8Ya9LL1BoexfUhVOg685IwrrVHOUnizbpxCxJuDjYZtTv7SzgA3e+ZDQWj7
FA3ZDjzdY9k0pn5SPQB2UJD07j6ZA3DokRXBNcF+9NKwoMVqdshkOsFdQDS0KfgtBaUWn5JqB/oV
UurapuFzq6cDTiwr0hZ92iPxdnjmbNkVK1J2bPIxhbbVMdYeLGhv0PRLWkPUhgRc7q7vRTKquIpF
NgcSFMyuOt16lsL3mW8Zw7jcdmtlt6ymDi4WeHQ/Kn6SDCvMhITzTGDyh4pJFvGYjfNBH5D3/zfo
fieS2B77IjO3HgBqiYhLE5dbTXYGPPWmZAbCzmhJOafnCbqsAB8CeCyM5+iIK8m6WyzinRFNFAQC
/49HUvHV3FeBJcdM+Eox+aQC3KsKLrpGzxkzBo/oiCdjQxp/erPMkjDx2h/0eXPFwriRmYRQG/vC
9LKOqj10u9HRFHf/wCcNIR0sgnyk48FVLWwH5DmjJTjbGyIhLggM0PoFoDtD/aEZUKP9fHjySqHC
UVb7MjH/uB5HuKxo28O11HMOwHazxBBmooX8OTwsKmPNZQAHc7T193eFPsr/FZvtUY8AokZqVai8
7nDqP9+DGv536tXPFwRWa3kIcoL7DpvecCLep7IeF2xXYrjGqWyNPZrb9RrjlModPsUm8SmV8r8O
7dBKpKuHisinQQ2PObwG6BVSNCZnxxwUFD5JYr1Bnkat6sv4XaaZwldFo8fal8qKH5OXMXjFWFUh
0KCucZytpNAbEg7JVbhEQ05fsPGMyLZ5RYgrfl0fKs6w3e4D2dcLuq5XTTlcG8KJAWtz2DRzrxCt
UX1RLsEcyjMibEXlVZM7oLfFyLRU7crwkFMZpPJOzH+GlXLFT7QibbW6mDiaok/3+TTI6WMCxiuz
MKJ3zoGlWXM4UuRH2oYe5yVDvm6NYHere7sSqN1Zfno2NcLtgY3Nh7x11DHvA/GG1RSeNxzs/sZf
syCyebAISyUJ5mAAhlNfx+DnmbU1Yz3zAfXyet1KHlON8rsVmWe5Mdd3a65Syex3WIO7CWqP6s5g
v/2IIU0Kl1LahirBta1KhWD8ZvvpT7eXRXBbF+/bZbHRXfrK9/VQGPDGoUCpVcpecsf27Ioa0NN8
6Cr3y+WXS1bRMk5HHmrBYjjgfNgzImlGXY1AogUuTihzUxlUy7edbIA3OG6TT5ANExZwbzSwbgL9
O6TW7MyJTCTANVdYQHUyOCJT7uATTy/7eresybnSPhWegyKtvVbibkhpwCU4RYxcHK52gZu7kg+S
rMKtQCybiKD2Uw1FPOrCK/nvY2aeF6Gma5BTf0yNr58UijY/ll26DW3k/w1YdvpEV80Ce16pjVgN
GbXM6dbSQN4bH5pU+vyaRYDUkTqdkj+Ve5EtQztgghc7+p0OeGFAsbTUclCQUx625ZfphI2clNOs
K4ncValvBua+8lRnpwtQ0747rJrD6PERJWsKd8SMq0MFzYyPVRdhAOYa26eONjSFjsl0W2UjPTII
JcE22gEEXvF/GKRXHbyYzsJTZOQYoTj0IWC4rdBHiKQywA8ocbtOqeIQkaeKfqF1xf9Sp9EP9c65
SohqtgwK14nLxhr+m2mHy9ygZeCXqAtLkbkgMW1jJN+bgJ0807Q1b87EvmroEd/4fB1D5G7oZ/MZ
hrI6Sn2/QxRXJXiNqMQopuo6K1ipHPxP+lUE7uHWbn30rVw8Hg0zKalIxVBI2u0w8PXSCroNA2Ie
ILyLZ185dwwKGgrtfoayuq+JgLcuJ9EKyr3Fh+ueI/UpjxRLjn1C1KpLA+xnolqllTtteF3QEAvk
2phTkgB9zf9GvPW0SrapBNdYaTCAWYE3PqvxJGbjKflj8oIyty96RTpS0Mc6Y6vpNkmJJsYCaiGM
OVgvA81U1SDAH8iWQ8Y5nElBEn68maEU9AmOSFA6GfnOV+5lUmGmjwTil1m/FjBMZXlNGUuYnj38
royYgCiOVnOeIBNCA4Jgm8r8sJbGltSguMiPa3kxTZ94+o5Z4jIuPH5Tk7qiF2ZYG2jWDg1baZpY
jWIbQJ+6syBwhbQW1TgrQ9wd0hphfBd6174vz5pxNmxXlX37n6q51N/Ao8TBfU2Dpvqm5Gm6wwtI
3hQlC0KB4Dm6wQEIUJIVB7tfBeX28Izhs5zEoKgU5xov6DBOqOkqtq4IaUhA2YUYP1MwEQ2GrzKP
znFsbw7eDhwZoc8y6949OHylAZaq0AgWe/6yPhKHcqec4LnMJFYYL3Lm95lCAhQieru9mmex+Q6c
T+5dd4RGZiRnq4m4F5bz/kPP++a8t0MPL9goP/NdAMichLOtTJRNMvEKxkttFBIoWEcoUJAaJv9K
/jVR/qlLci1817poruxu/nvHXMoKiCP2LdeuoB4/p1aZ5YZCcGkPDVvUA1E1a79AwKxRz4OF4I5B
EwqIvkfbz612R6LeKTQdmGbpjgwQXwlEoVDVY71ViH4ILt4JafEZyKfIzhtb3MAJht7YhXtE3ltI
Ayc3JAXZ/rOoIibwUjqn1tj2lmW1nP99kDqqr1y1N2cNs0HqaXH16KLRTtpzNqM2irLLaEWVSk7E
ARCZBoSx/U6kw93sAz49/L0tqFibueC5fnMl+5V8jOty+qVOLZmqQBNbT3eIyaCcjJKArHO6Nk7A
kO8VcUkoocQeNWTQ6sNZ+PQhkMR5lshgybCI4U2D1ky59xzfZo8qj6gsKz2/spFcwAK684reV7XV
0zGrF0kB0QmnhGaRwZkF7oslMSVaC0vw0C9XTizKiiCvw9Al8ZMTTkT4rtxXQJpkFj4O7f7gG7I3
A8703tZOxMHy83aPXxtpqRpSTpSVNRgR1O5B62DMqmcMhl+RmhHBRHbQBIyxdE5UaD7oulFIejez
sj/RuyBDqMLzTCMQDxFSKImvGlB6/wr1eK0DAzC2hK4h/hx+pQfQec14wMMUyERZ+uvk4zQoChhq
rTDv4GqfceIWCmKY+Am3NnV4sa9WOOosS9RMYNK0H1t0ziT49/4qlW97txPdfTigqLYwkTx7cp82
9I/O9wDcE7SicX2PzxbezMgBKKTXozT7vUg8gXDaVeflmloNiUUn0CZBiz3Eg1d7yfbaaER02ebl
yai3gXLiGkCLU2U+Qm5iUIH8ZBADtvDacXpRI4IdUrEYRLUbgk8CBNOGzemfSv1ix1ai6Rt1eAV7
QuuEnptPI0PzJ4BXI7b8msVLZFVzCK0XV3uyu+e9y5EoEfCx96m/ouUlznTl5RxnM2oMTZNyRyH3
EZILGdrp1vYkWiDZqABSY1U+gPhImQY3StLolOAdK/QdLP3UxQPg0Dz9990m9NwMo779C3ukcXKd
FFBcE5zCEoQbjBitcfbfYN9X5kZ/u6avDeRLsWEXnffad1y5uuYkvb0d4Px5kVSxpgNDbR186hKY
WmrOlo57itPawUGJndKv/Eh1l+s3y4imp1Vq+SJKPlj+6NbmYPOab6clktN/jcTVqNH3h1y5jMN6
iJEpQe5NCHxvSClx2VR9pLJ8QhOLlfJNX96MG3JIWMRF5OmrCa1FNniV8OE0DzYBAN8uQsN/UPPg
21AsSmY6ckPktZob82ZAcOEvZ2TDJIjay1/Wt2cPwTS8gZTORlYlkfKlk37syv/GxhdhPVHAWavn
+Eb1baKwgs9WpJp3YazJ8kzDt9kx55qloPFrFnG0VQL1v9CGqlynSorcQ/y/ULj7Y2pEeuoh4xdT
pvK4OgYtmhSBXP82AhJXtYy/JakJktovnFptWAXN+02jgNKoA01PPpmRrGoOFUobonWDC8gD9mWL
jODF862sBhTwY+8UJMxFWw0Du2P+Dpv0a9ZKUPRaP6g6htLGCgPbJo+JEBRujiXSQgOhrseG+V6/
KAqL4XJY7UJR/g4qKQBv7ZRfAsF1ONLgw1prHBa3HkXN0a71+B/Y+R7WtSfP5bJs2cty7OlG0zCz
PArbJYRaPSDyAjsoB0xvlW3oUXaW+l3w50QtYvE7ULG3Ri+VcXRCZ28LNtb92OW8ogDJOxyVrtE4
hspTMpJja2eoywVCrI7kUWQiIv4r1WkORygMVA/rHU9MuHq8Ai0wrrT+GPx8cLaXKYRTz9ew1rO9
uEltybx2cmZ0ruJTih8m1fyJr3xkJedZfjQkXCDyT5lAvfhx4d70GKJ4aTm35lSacXMhH+p6xmH1
MmnAMbtIQifox1VZIP6ak7ym96J0518+bXsn28jny7xSF8JlHVMMdj1dsxMvcTbSXI1suZA+1u36
4ScK9Qgx9GH5QeStXDituXric/xHLXHi00cvDwUmlmt2gCffGoOJrKSGRwgajwV0880sGuWD4jVZ
KiYv6WQgKK4M9cXYG/tQu1+RZZWFlsWl6JVwO0e79pcJ+IdMOmoEvW3fHM+XGBdp4P+SQigBe29u
mjmONhNApLnox0fyPdhSeShb+n0CSIxpckdmi2xcugACgQp9o4eYEWVX1Be63GdQwaT4Wjle8++D
qe6B2vjxax7jsTv7reX3Li5hrYSToIbMIdZJrWy+cOIw7kz5c4zhQrwVA+GgR74vjGFRecCDUAz8
5jnViCezWKvYMguAK0O04L5rwAO1iU9KjcX9qCBSBT/6q4z5h+HUVuInFoNq5yLMJ892eg7F2kS1
SfpgmM7dmBZyzXxH+PPDWcxKyQnJ5qPkfHTZGs2nL5/Gy6Nb4Kff0hZ08i76Ia8eyVfPKszYopli
ORNvkJkGADk97/zYE6RI/gOP2+ViB7KU0aXsNM4Fy2f3or/nxkXCaIExaAzLKu38pe4JJYZud8tZ
jEtadpB06WUUNiCQ9PomIQ+9mD4llV5WeT+5qseR0qBPEqJ40FI2mFbo5ejRa83CirSwtREH93pz
MrBeqhMnLbVl6lAsFHMeaTNgwp0koxfdsuscDq/jaoUi3BMhIr19VEfbAgF0lsY0mpeKHgZdBzon
1b8jvheaRcjjAhgtZ0GwD5khZ5Xs2kfdQARq6+LQPi+aCeLJkkIkSnbQAEg0LE4HKhgHgiZXJEPO
t5KzFkQojenj5tt9DYj4z4Ps278z/xktK/d/L0JFEXByisyQI3mtX3fO/ZtcctBNH44FWlM5i0RG
/UuKEMvWsDp59wwthu380syBhcqziI2hNVmDiFsa5qT1oCxhqm2QU2jse00jMzhNX64Ks0yi6yDy
+rT5yUpvl3Ea7+UOPa9EU7TJl48IaU0S1ca6DC9PYdacUoZkBCESKpAFtyEvL23fn4Bsfq9HenYG
wPm8Oz3I6wbMvp5B0CPe0sUiQRqxlW/YQd36beFwkuAOkovOAWLRIzmHBJgoNpT0njcWecnGBFC6
nIcpnjXIOcr4IFgcwD+vEm8PbR68zRvXgVh8pX3B4k0cjnVFTAay72GhdyfhCS3zJL885TS3D3ij
EhYgGe19ehELAQYLDMNL9hlCCvQOtv2tjsXXI2j8s+ix417bcAr98w6wENtAYJSWS0XDYi27jcV9
5Rf1lINEKAqDKTVwdPvrUUzRKyR5DcMBqARSEfvrtszMTiE5ce2Gw2ULWOX69vW4aELIhSNg65RE
DOs2zPlSi9E9QgzaJ1kbeRV4A/oxPG6StXV4veW+x8EJGPGrmtPQR8BDxlvrx9/jlES5fLOk5hs/
3e+I376IcOQ7yFaF4xprdXHQfzIf5NXUdssrzLJUrCVqJafVMN4po/gT0f10DMz2x6gQ792zdbmK
PeX9FeufFnrc/UKivPitNhfKOnHf2M5SIdmsKbVJ93lfhSXsDQj9d5uxIMDH1BX4+2LThH09212P
+JrPD+ljO2ufQlOU/HNiIoTUvGZ2SJA/7zTwWljy1O4oE+ulwFSCDA78sw2YuomyNDl+jdvECCIr
zMDL1XvfueLiD4W8f/a7F/2NVwztNFqg3fp3xFrMCQ7eVN037hlyaJMd/xNwsQDPhbe+6CLed+d+
ef4CYT88XYbveQ85f+APUZdW3fBzCBt17LmmrZ47/tJR8vcWdVep54ReQcCNuLmCjZzkpM3JJzxo
wzJ/2UXtU6et1JgI6Sp5kvd9AXNN5HQctwZ6K+Wl5QWl+xWFvT0ugrp9i8CgMzvcSmref+bdZwOl
+1nchqltHeZlGmZmQR/ilyss9480OdmiOPsv2fnt6O6+de+PV51YrnPwMYek/OlaCb2N+j3k2awo
t+4OPjF6WpQdwOo4pD/a2SxSCrw368R0Njm+J8Abv9cKKTbRqwQOIVppNkZWtIZwV3E6QdQtZ6G1
naxwRKt+n+sDFv/vV0XseG3kFafNH7FrrQ4Ym45RHckz6XeSZqPtekv22Q7psDZ5KuIFul2sBGPO
ghe2YSPmirzPPxv6WCWno7ARScrWNM5+lwh48kWfhKzxM6lnHExEB8brieXcNsoaAUUhtMtMwcJm
IXA5feFu0V2ipadgzxxBZAL6LbmovaTAPf2BgNE0LgFGCIi146DEMob+7Tnk9/BfvHx6/rXr+/1Y
F5B+PAS08V+GOJhrb/LlUw/bmG1IKe+fhhgXRh970reGhGaXG9UDZEodOLtZX+LhM4ABaReA9ftU
vnMVUyQDE9jgaudjjb7gbtuClEOBpEQ0KCkgYG8KAj0s2iYXIiDtuxa4VOs7eh90RvTicjfi63mO
oFqrm839Dd186wc13GfT9whkZK7k9bMTU+5B33WCud0yzCc1u1H5YvhrO7CH4j9I3mVR0KBiAXVX
tJFb+7cHqoYi285AYsyh9UH5/wYIH63d0S6p6FwrLkGBbsQWI1/mAccHXqasno8jIklV3XUCY9+R
vVWNjcUVwnxIW35JYx2nSL5hxYgtC652g7sWoyN9ySleuGZp013D96PHNrj4tPgsiZ1zSnTxEk9z
iywxNhSrdtcEbKjTFBATGMwTH9yUSVYCXi6SXAexhQvfHSbMP8p0JCjeJRnNAdaWINxl42XO4bOu
6FIsvrCd1EdW3frgX8aVWGMI4YPR4c5oJqrAxV7sOzQB8cg9LoUJt+jT4/FVUtARBuPw222QN0y5
fyKyHCKRYYunuCaZ/W4bGVYY43evxBSOov/A0+0KYjtbXxTxjA1WN4UFfCvbkU9GUrbSOm+ifyre
O02e2jCsnsaEU8qu0bIfqHwXveO7rrhno9mf/Abf8zLbvE5gtnRhL465QLtSnrcOPmshFR6VNEf1
xvAURUSOohjltPl9aSE5t3wsZ/LN3FJ2MXvsavDSh9r0Swrh3bKCNtFCASa8x0nH9X3Zp6lqnUPx
Cz6jb+F/Qo9MtTI/yd4uM8U5tzv7O+UwplFG0yve0sv7UTGkNZhzHnnk4TgQDwcO//4ASKQmHVGc
WzYrCAyLQifw2fnEvaNStqiXvmh4D5T4Or4QZJEZ+aPyM5nd36IB52gZiR5pWwWUR9DhwME7VZZO
MfYYTPHv2t07Xc2uqDAqw+OCs5gTjB8rOqWwupm7+WMX3k3tPdLawvdPWDzpBhnfd1g/AXSSwqM/
MadZfKvEO37l16MuRRozplHvKbHyP+cebEp3xJQZe889vAX/LK6dSWG892fxi9eEx0ACXJZgE35Y
8rkN5//brkqO6ouj6FojJeJTjebkZ9OfaeX1e4aYCAitMV6hFBlsQ3SNTCUUlBvnsIw54KkcPEfu
MgQWfPV8wnd3Gp5vFN1ASBPYpsSqtUPt3NlGD/RM5XZ/PBOwknwHyU2G5gD4r80mZkdQIxHDNZ0f
bWObf2p9OuT2XIOzPzfZFNc2M5Dyi8GN1UvlNl/RcAiVpjIdaqJmU7f1PQW8nhs9AFWrfzByXN/t
ceSLZfuXo5/69PTyPATJS2CUYUFhUabpOZx4ErmC8pt18Fa/FrhcSvVBwRto+sraqfZu0p8ScQ1w
TanJ/dkJBr9eRzoDPy0KYkFY4wx48RWas/NmqgyDtQHdmvgqt8wMF5YMAJYPV3ea+Mw9bvDtZ/p5
bnGJGLQ33JQJ6+GPMMy1vSCbueo7BHy33xXJqHZIOCClci3w7Bj+yqqjT1bUgrJ+5FGt0z1Dv8i6
eoJUmbm0MhzJozzu4qr+nKwEOER/RRr/9VPb300Vfzu9ot0X78MhE7LEDL8RK2QTFzELKpbp2mJy
3KDxQ1yb5r0U0nd19N4YI30Aj7nefhUUmB0swmPfEgw6kJSII01YY2jmgVoSv59mh6WpY4M0VSQW
HLtGCvVPy8sqqu3iik/XbBYEdSNm85fbw0u7lfg1aT8f4oiBc7jLVdLJjM1/o1gakdjoMtclHtgI
dPj3VduH918BgQBaYGJdWjBqdJpj6MURteW7RuFWhKxsWgL1tWHToFw6WWTCDr0jIV6MUi6XSF0M
3xaVIUGZlV+J5t8O7qlai3BTAoIpuXxd37NO370OkwCDStorS+IjamHVSGBHJHWfRI7p+JjnAMAh
lGIYPfA+WD1/KzN85B7oOle/mR1mC74svkZoEY0UNc73L3HGELs1MCiZzfwzPNE3L3DbISdupFIT
1OldJXKPMpgO5h5XdQu7G5ERvFcJ4K4kFQzMX7tSF4r7pgLwlfcFrn0W9Jfg8PhGHCQXA82hUQyW
ztdI4wRkbmCiscUqzvY/jgYACSxBW8TjZ16N5bWq2Y5IVgoGNFb7Mo+9m6UR/GlwAkIe3+pyprU3
QpkD6AhFJIxw6xnZXx6vb0tyCYDqcm5Erp0vu1e1R4B0i0PAEwj6waNTT4rPSkEqP+UfzdLkFqt2
1BudZ8x9kPyCMio22uhVZjc2Xm4Cm0UN9dUHzrg0SoXfe52DcTH6sA2B5yKArEKWOxmmrMl/bhKX
oqv4vLZjCD/nUjDKl79kVeYV9wW3RXgOtSOlIP3K62UfVotqH+/TNz9PIEud8Vd7cEWyY9O5/WoB
Izp5Wi8zuVYNKRD3mxaDr9R3yFuapuLcrqmOE8veOOb3KzZa7saXsnYpAmYWcefFng3aXTtNldlM
ac7UJUsBMKnv0AhmfPDgaNnsiQ2hIraMoEKdOReUA8WMJYxHb+9FaBwOy1cut0KeNr9gKzLxNuCE
kt9AaotA3a6gM7S9W8jf/Veh0hsboHqGH8fR4WiZwgNynmTVzBCNanVdk6fs5sbGfl9Lkblpbl5a
3u9DxL26ENPpf3HiDTE1D+x5jX1PC2MBTNa+HT8IB9U+dBIFSGfsNmOo9m43okEeYpNooDwz8nvJ
fvBGAUB9xWnYGrg+l6DkcfSgG+yqD2747gtYmMLHIg4TQad2a4P2wA5e7KcQHRAdlEwIA9HkXOG0
OeG/lCYyxQD1mVlk3ZiX5FBuAhfJ5vHR9/nM+/xumQAyNyH5Hj72Iw+jB5yfaHKp7V4s4LgHzlKn
IbVZcCsX5y69qNpIYIjhpJuSmUdRzpEUwaaIsVVmxuXSGFsptNJUcRo7Ka2axoWe0LVQ3COpqfYk
kFuoPA96t0FJFnCZdQCy2vnf33R8fATZMGywwDRI3bmyv2SPTLyDFVoNF8v5UDT1vipUdJgtjFyY
EWDrbqcCQlJD4wjGdsNchXYiVhFYCXRwF948Ab79JJKHPhRlOu3yvQgxtKqLgFBpsf0e0FCMfTmx
8DScitE1ijkOieZY7vDOlKt1H5Tew+WUvE3EpoN4WeNUDweN8RZGqoOSbKKP5r68PYdjU2KChP6V
JklAwEF+aWaqN5AV+N8z4zQN2kKvQfi0YuOkDvPKVKfu68N0lp4YG51RV0rbWkwPRunSpoijb/O2
ZCeVUVMMEjsRObOzb8mLRo0/iW2W4M3GYI8NMu/DxI5SfJRYVBtO/CiZna8L/F2OQFoE2mPZFknN
Thb3ufw60JiRnUo1fuL6yXkzZ1S6fRF5hsuArXphXiHpuO+NXc5HrpgDC6tC8URvsh3QNL8n8ytK
/6W4MYWy7BHhLQalteNyX9jKxRivXmD6VXeCYF6GzGAGGGTPw9KB+ljWePPdhGDX9ywj11dvfbSD
1FeOcZX9utkYPV4akpGMQ2q90YXhjDfd6gc6Her1I2RhFmwhMYchZKmBxwGdGNyKAF6DthFyls0p
jPQoq8DIpfqtvhcW9z68Ceo4CL1A4AXHPEke0xVhQNkTVddiH7Wwh0kEZRsAbwNnun4+KCLXVH6d
c+c2+6zqrOcwh92lcK2LXb2HQX+nDhEc8CpasMEP5ai1olrlFiR160yhfnkpuKpXHssnv9Jp9b9z
4jNsXzYqhKM8oBs2kSKYOjMK9G0Jf+Nxn3PwyL+z3TpvD3fsYdZ5Y9peqsGz4cSFoffi01waGJxO
EZVQ4dpDdfPUbA/lIHV8FfEq0GHs/Ovt2i/I0s0+nisOME35XqIjFUrqJGkuZjAnEXS1WBiDNWYt
967KYFY7eRGueHs0OktX57AIus95/ZF/vPCciEk6TLeQ3eM+MlTWkIBTdVjQzCplA1ywCUoaMHQD
vBadsV9qdxnhIvsrcvuCoUX6PF7Kwp9elgYwRkymk56l+pXbwBsiSrvmckcAi9UQoR1JlLHTQ2p9
oMW20aAjyxRt/gv4vvzkIS4eF8ywV/gDVGwNHINENRoaWE0Pe3aKwFLwnpuHdqY5h/mGQL49pfrG
938+ifHVwSMuKWrdqqaOPLKXltJGzmcolw0tug2NYejKBn5Mu39/nsWtBJCRTgkRP6lwp9LKJNmV
7ChwOn4UiJgcvgS1XiJJtsbzvH/afLxpJnR+geAwZj1i+3Ftiz0YDMS+32zzjROuYtBYIpq/1Hj2
N6kO3PaLHfUu1KqHe7MTOTclmyxaOasGH9z3PKo7DbDUC4JkAweruVcw17s+wILmhpq+qpCmz3h7
PKFauSSg1b1qsSqveb2vkjRPPGNPKMntG0pPr3XlV92i2PKYMRusozDVCbMYWClZrqajRlzrMTjZ
s1Psl8Cqu8DIqXmA+RMOs0hEQfR1VGgellytW5MZpnCAqYrgCuddlfm/3xMeNCaebm4VNVPPA8q6
FLuFD2Cotio0W7nUml5DMzi1Ue96/4bOrRGDgKlH/7YqW1rW9l9liYVLviOfWo9fZxMFuy39AW9v
60vZTCWV+nd5PJRyyN9XOeMnNNYPyZM9NyDCZgBmq5eC2K/j3IrjSgQ9EWTUeDmJIJW8GqWP6W5o
T/1QMT/27go0AIXC5g+Rz3C/Lzy1rd7ykKnZBEBkZmfj76+W2MOydl4csgB44HHs2WSRDbrIyI7L
JCZBnzA48wnAFfdfDYqvqNkiWFfbrEq+2NacU0vrR/I0AqAf+BM3qLU6zOXseb20VZslFnyX76s8
L6OK7M5BWpVAnNY59eCFwIdTV8n5awVRwvm4UL5F37bkyBkxYqdS9DUcbWdspXwgX64Y09w/8ULV
AZ/cIeNeoNR92mr/PXGYUp/Nypr5V5lhkAyWOJFGzMQqWFFjd0XW2HBLf9yVaxmxH6isHsecJTAt
30KMCYOIHrMZCQJVh68edN2wLi/NOQlCZvUzWjoz79hd4mFzEVj6HE2Ymg4nu5fQSTu9KZjxBe5+
5YsP2BmD+69ihJ2GaQSFWCP6I5UA//yZaB9x95nVshD+BG/LQkj+CeQY5HHFVaISubA0epjuxfca
8ZLHQMhWGUAXBh13p5vTXCqhgreYCl4CpkvkUWzQUKYVmiz5/jopeec1fjeis6Z2aqy1w3HFkCIF
4c9CG7dJqnrROvytLQYbUFTK4dowyv/+kHZiT4eVj+J11dM4T0rxJT/G7ZaLycFbd0VOUaIWjQcE
FpR84AhjQ7ar2iaiAlAFt0Nu2MOokBq6f47SmGkFnu0ApEHSqobbgFhDyTi5KVy9bBpMCNy2NeSc
c9AFLywAZMk+A0hBUXeyaA3AlMx++3cJm4YAIqBhfn+2MzcSE9Hp4na6IyZ2URWyCpBQrgzM5Im1
rjzdTey+89Gdf/tH/WnpAc/4F0wCEDYmSJ/Tc0LVmcXJoRmNTJ4HrpVCb8A9obxKq7tgMVMKPXDY
g9dZzuBRkpXOOAG2WY+3GdPliDEmfFIGDCxy9nQnk32nl3Cox0OPMkQ7LoRoGeTwXZb+LVCmdtBB
CYle/KFBJPMVPiSZAm3Aavr/l3IqgtV76PxzM2phIInRmAGSfXx18LnliNS3fIXMBRucA0vhY+9s
cSeWo03TMy05aRUtFos4CHZApoL63UJjXY8q7ARLZtHCDuM/d8AUR6KW4LPq7Q7hGoWQ57JOSAc1
YLZK9w42m3Pb10Waqm3+p2h7yraCdGldmUKPScaYo0FIiaOMEGjh1FLUO5KI8Vm5RuaonzvFby0O
hUtzZlzSAJOLwzQDqSsdftEF6ZJJaWW0R9ICMmlWUjvSN7o27A6aIYIMZ3+NjFOfBHMIiNnQ5CCv
ytEntgfc8oz5pMiXzyPk746ZmZ0LR6eipqUEUfj7DQYGWHXCe5GVSE6HhOdlIsWSmpivAGNfuEAN
8P84M+Dq6Vzn9UXV6wZbukP3K78W7hoXPiZQdQLIoA5MbW+zV/FseLioxrRzDYNV7riq6KPCT61/
FFxrdCId9PF92vjMS8pTBzwKl1b9gUxl1GBTSpUthrz6RGHSHRw++CAW6XiZyKmz+oHcrZTsiUUt
INSjvfgTgHSEZoVtjR+yJUqdpZod+moq9GAWstu6Qldefi1XW7NF2XNApOAtqM7Xb0kGxrAFcqbP
x+SzQSs/kkJ6OepvayOt58hG95b2xoH55jm8HlYukIjrswCDG58hrWCIOdZ8gCa7BzcgpW7CYxDz
4j+iToR6XFxkCQcBYvkSxzvNeFU9cyyu4j4Yls9XcbooXMXzOKJhkVugQeVhRtQU3/Tni6e0fe4H
wyyaVVGeKtAXrRJVxmQiYFddS0DL3mDyPBnhQN0Qf6BIHiYS7CKna3SJkl3MZfnEK8vCRklg4IQF
J6Vg1VyjBrntDMS0MAYk1aTu+xzTgz4LxJrOb6RVH944qOrVILFToNh2wgtuencwKWEqfKtoTMf7
T6K8oVWkZXFIEgbmXOY6XHY7uSJCYtsBSU6/jLJo9WR/35s57Ni56SbZkwLhHjj2nggsQfaifFpH
BTI/4ZdeJU9Nx8VpPjMGAmCEoTrNbkSywQ83/VaUKAlvoTPAi+WN4vBN4XtSpJ3kqfM5DXCz7uj5
9EbgzFlQ/9NgYp4uQKccQbonFNtX6vjcZH1WtQo4KpbRq44ED+NpUVkvKZPjl8I8ThOSwK9mn/ek
Tlzpgn7iIYrxDh2NQ9NfKX7F9GU8m3g6U6nwNcaAW8Ip18j5qLioxo1kEk6sbf3PqQ/gcFFkacbK
1odgYOx014pasza2+kmgSazrfdQ0bqLNpVhy0hneX/t7dTNFU6CMlKUlrJ/hJRUMVn+5MnZ7//0q
pksN5BymVU+IedgIm4hQ1h3L2xUdXsPT4C7ELtGbQoztlDABLvE7j1MfWW2ykF/EOQci9VI4ZgmG
w8NkPsmj/QZDF/bJrOhwfXY6CtftfOL0pAFEV7h+jppnzQCGlFuUI1cwquvfNvKHbv4JRUg8wOVh
c7REH3Wgi7UEEI3FXEdlrdfAwGf26xJA0UGhJdpax6eOMH64G4RVI4eBv+JgEzidKBTYW6kziiff
uDe7HTF4gjVGpTayJK2Rk2Hh+HGar1+6E4T9sYJ3y04rZLVMTDkUzP1mll4cysPZUrh+fG3j9EC9
4U+dHVGF0er3N3WS5R1U4DO1gAG/uZWDnbFf0x3ZzO745ELajRx5/bPdm9LHrqGNkmbdEn+w3VEy
djyj4XhIxcwCHzE6YF+ptATWAdvX3SQPuhpauKlOOMxtof0LDJk7KujyuWNyGldXwuEBomz4mN7x
OBLlTll1UoBqZxXcnswv0JMmyGu+eqxT1bzVVS2rZphZh4TgAjLcdYPEogDe9ixDbsbN9sR1h/in
cXyLghdvg+Tlci4Jg3VDKBTECfkSKOzER9VcrzOHeg9T0v6rr1WGx8oP2zhTVGeXGEFbup0P3ikD
NwYX9MZZ1yWEkkDW57QxxH1P+AfA+CZ1Bc5/PIznTs0OEU+Ap9ocvB0ojJRhUsZvgFPCYdD99SNi
+tgvxqaqS/QhxSsq56zxwtVN0sMxVzCcuJqVdGE/X5q/5aHPHNsOeTWWZjhgk5Ts4vCPrYWEkj1I
T0eh021reZUTrWJLiYEGYf8DWUyGaUPuuN/sixka/W67g45w8a5FnnaE7OmyGsETisoVWVPURVOm
Ab5EOONcA74VF1u+umfj18c4Kup6Gb/jW+Pe0ppeLqtpW8hP4H84iSFjaTSHRoZNXz2LgXu+OGfe
ryH+xvuZYk2IXB3n33MIT8p+cvpONKISi4ViMC3RvFBJW7xecEJ0piZZ/sIbbgE5aFh0MN/9ld/y
NNldSZkXEGsUWXYknonfA17uKJT4nDhLcT1BspahGqFZgFwVvutuGpJrSgEBlQt+Yf49h6A6Un7a
iDx8E4xkiO6nMCEF1xeQcPSzb9CjsMtDZ+1RpCirLcXpkc9HE6bJdDf8MRC+bSzLODkKwH+HHVUy
b6zgta5mWCEF6Ay/xMGBrP4Ix2FOzHOkTXMNYVDcklxyfmF7+id0RZc79XHgkTYaTVBMnZdioh6A
5gXy14nt37N61u1I7UNDuQEq5ba2WNK6R6A7HhSVtRhWCPk3wqh+dfUdksmwxwyCrwf0m4Lz/R5r
0r1DOPGqWSehn0giBBQ4R1B1JyqZJh9oNvV1PrhUGzMhJkeYO6vIVFap3APx/iE2kb7XHcd54kLR
Qz00u3Vhruhhqn3tr48su/hSedYoFwyUKzt+SxdzHMit1xe71RDnC90aQoGOsZG5J26boeT/ipYW
QYWeR4Wd+GVBaGgZOeH4pigyVAgGL0PROfNBSbFdZtwHQ8EBxh8eF50jYR7UGMBN5Cl/3a2P3pAR
CnQdbhYWNbcbNiPdSE4mFlXUJoz7Sxfl8fGl4/xD+PFt84VzryBqMk1to3AXwSMWbvolgycE0NjO
J1JzmK5+qHUmhrqszLBF4vUaJP7LNRUjgqAh6T+1pFhVbeZ9zaOA8Tj6N3PT3cmgpZJln8EYsrEt
9pzmD6GdF2V+gnUb1WJK4F4m5LvwyiQIdPoyQ/8Az5EtC49T7qGTg7CTNveZToJSW98M4D+4YbMC
K5uoQM+BTa3pMj2P1bnZDfYwoDd/o2rSPU6IvqwsnL1eVFMBxhzPhCqK5yRJa5KeoqKof0CheubZ
fvHH8LuPMlapdlHQPxKUTc7aCJsctMc5+1ahPtDoTq+z4kkEEktMKfvj2f+7vD3cejo/bkAI20e0
yX/rBr1xUEZzasDtV2eE/aqnVsPIOl6Z2JVVM8OHxNGS/JOaEMNjKqasHyMiRHY+I7lMarzKuEZi
3eMbH29D2ES0t9i1dEw4Itaf6dgAt23EkoztclxmWcK7YoJJpAQrT701SbZjdXWkJt+CUEts0RY7
aMKKm+I0ZycJ6nShr/Vfha4ZAsnedv0L0YHk0ooOMVNrODLMa2Z28/2G9aaW5pP2o22mglnT/4KU
ojBR9Di3ALAjVzzu5Pp/T0Rl3nEoijVSEW3n8fdmhiREJKfhFyDlroc8RbYzcsLcV+Gua+eQmYFB
7Ee5QQPgBbsceibzBMtjgWh6cJQZpFAE4lnV8aKVArsjaF64n2TcwLg6gpcB9A2u256kb797Wo1e
PHLn7PlXS02sc7REk+WL/1LQ6iRAyIiOd9EqlD8YZE2VOI4oTH/Fw+KdIB4hBGSDEkRBCUQlq+is
c3WDEW7ZFqT/aLxrWuLkhusQNrVvbAyhk76Gtwt6KrliyBLT0BFpmTmj12Ha2bI4/zeQZl73XOTB
Al3MD+KzkNuN1d+mQnyVKaYTpiOXI3OjZYDvhEFuDt8+Q5OjhU7H1iqcJUQo1t0yu7r1hqNW/FdO
+xKcaO8Vhv+qHumywxGMcS4QL3jMcni2/ZVntZ4kVyYn27ejTSDGr/Rizn0uTk4nxV7F5ZhSDmn2
obdA60B5mkNpAYjU4W6M/uLuERAh4TjRZy1rHkC+V/0ttV69GaRaUcyl90zAmlsKs2RXrLGE8RwF
R7xntMIOkEaiSdvYwQbA/u2TwXFeP9y1hRQ/H9pur6v6anPpAKEbju+L8FS0+XZop+32eB3C3nm9
1rM9xsuUOQg37RHZ1bfgRW5dlioOnIb4ZqE38qIHmIWUoajoFaMDM9amznjHJDYBnKHA747wI22X
RF/oaG3JSyuiVLADrkmSwnukbJa7MUVSxBC37VXxMSk4wutsycccb8dV8nf9E3lPdErwAUBgilF0
W+sKrPftNZj8l+J37ElqeBbNQGF6dT6ZhOWHsC6vhWFoQvP0T7i+TeExXp1+0wBn+NxNQwinTXz2
zqdSTwgCHiuJRgl580i7jGFjNx+sbQI5XmRo2ywdHh7YyYgOgZsOm9mVDF8glpRATDEAFIJzKcKW
3AjY7YdHwUY06nyOKHIwf214GcS+TIXTYDlPSDvv0aPUWR7zb+cfWItVBg9yT0LQnPQI22kcbl63
Puic/yOtwl9SILH7rjnspY+fGHXnzlvc0Drb2GmK5lvaMA6h6b9xJmADXlKEZUaJXMljCCgPQCHE
rJHIZrceUsGNNYmENwWPHdHUEBFsupt7D00v1lNzUYMv/GKZ99+0YEgBhwkh6d54rYh5UNkxRMCd
NyyTIV0CCL3nAKL2uZz5WrqJJQNCGcXqT2cq5LbtpeEi3OnujIMLPU2J7loKkpUbSnB6XaLRq83t
FkWwUFHWe1gNAl1euCYupAaqbWs1WUHm/dyKORjvKUo7BoK4NNnLGrjrhBDR2iWZPzEN55EUJtjm
m6jGpnLtamJ5fQrTjGYC5YH5GN2R2CLaJUPcQ7KJ3wKxB1pqzXLYXTBtI6EcWlWMtaXxwbCVdMkr
djtWBiCuNdmmW1WA02stLDKRIvfuNbLT23LUzyVShnKyko5FQzKhhBOOUSYpqYWpI8453Y/JX3Qp
wuZ/USVPBvwx5hxmEMP4qt4zqGnk6CGS0oknk0VN/KneTLHdA+QzvexnfLosgTHed3aIoX7uJlbz
N0PQYkcZRmUGP6VbM6MzC1WQw/iAM8WyzsBWc05pdoqPqMOLvmqDSOzoIkmNwSYskwpAjCjU76YE
ILE5iYx5jq3glH6VtLWfZttXB2FwLZfX6MWq1n9/pv3Ej2/QAfyVh8kuPfZ62N2H5klKBBTakpJV
pjDA9iphKxSSvV1tLye9QLskQW7bXjZzBeB/ZkBv8rqzAmRdHsbRcVtPkWzbsWs8ztpS/ZgqFmG4
TjaGonDh4T6YqkEhijDu1HKcHzCQjK+ptpVA4yWFXII56P5X4ykOj2xLUiIGXgGNkkBtTjqYvUtU
ABXZn5ZjZ/r0t8hEI8TvtXj9VrpFyV3B4yg4yz8YEHxweYKa/cg64Vx82S1JCJEKyIsErW2L7Ynr
RMi6aFLSvu7xeaxEvbodaTMzDWQClAiDf1eXWk/ItyNtBuJ2iyqoOjT3vM5CwFXyYAlaQWqr5ya/
TIqwRJ8til9Sf8sBWFwwZWUfx2EqNjbhhy/O7ZeMtWRDXZMKLkLixrGEFvYceF6ylqMdyca/D7H2
+3mzfXp4MlfV6rm2mhamDwx0+NffEOYLXLGYMyQpzbmjE7AjpoNz4/O0zOya7GL+kAV1hOlhUjJp
Ac+45N0LVCcua0EKyqEnN5fTysq3QcnUtgprRE6vOPgXYouiBj3yx0k8JDAwqaz9D+6w1l4/s2bu
/0cnxVENgpyzyGO2f4i16Zdou5rA/CfrVuDVhAmhooJFaAl1ciF5UnXJ0ESEe/OS8SPFvfQj9qFT
W/vEopqI1JGF8V5t30hRHmvYGtH1cLlu13+LFPSyaYxH8ZncmkmYmq+LH6ByC9S+8zHAeLHpYBFz
NeDdCIYQZW28l6cv32mgNSr4GZBBM5heYfJ20TFyh0mT5tBlZwVzd30qoNJheh900kQECY/FzdXG
WhsoKJBtw15N+PhJsygtUJiaaJbMm7K9eQ+bMQ/DdMEMZ+TSAbZtva4GW1CSUj5LOfyvNrqT1PG1
lNkY1zWczOPnfxG3E9j38/zeIuiSnhl6cs7vLyL3upGWElxMzVn0H8Fdeb3EVHTJ9x5KsyZwhbfB
5UjSDFbXQ7PGFUqB7AZsPyI8T7xO1JlKpw6AVoI4EWnvk2LpkEnR7wu48qNG+23PTs8ueQ1pKwnk
qXIdqtfIHqZPBzrDLK0aCoC3DmBQijT76Q9P1zvYJI+DDeGqvGPjI3dKnUCo7+mMKJR0qsrB0IAQ
mTAX+HNcGrYhYMbSifXsqmg5zlRJLZ9VHnxSpQBIEm6zdw0z04ukvFdMi/pX+5vBNba+G82Cdb/n
2EZrPml9y+f/CjBDKSVmL2OqygC83YITwvFdXTwY/SxuIdw5tlz6bfShX/YlhgtFIsJz31Jmx862
YY9nhsjIy6Nb1Z5zR9w2nsTELqhY3ZIgHj+9nQKwYS4/KH/ba/xo5wMgosEZ9hlw/V9lcZbQVIVl
/moyANjOXB2Mj/L5DXMQFQLzoTnvfLptUEynFJ200gjxW54lnnxT+rynFV4A5yPISANiZJCuMqsD
IfA5q7fbx3zTlm4YTxGHJ7smXV/UqkRPNouScVpsvDuN1VTlGtYoveHPwfM81GqKeLry/czncEgF
nqBjk4215/NrGqPkKKOUpUIUNLJ6w5QzdqzQIQsuT4YLgztQvdrqX1hrXHHJPW+xLwz5+tkSUIvX
8hGCSF3Q+isedLna8qVPMKDJTwOYCnTFpazFeQCzPgNDzDGDh3pmJsfG5POFqOd/bqimy+13PyTq
cNyNFt7iXkBl669lG/W/Q/EHDDxi4weNsAWLhVUE5d7pdMl7evsZAJyd6sab/QfEwX5uVFOu7IuB
YcV0Ef5a33j0jIErnfwOamIbcBvCcCFRC0G8Y6+qbXher9fI5GN2UiJE+SIMykvJDAttBdb671ml
h1IEdv5Q0uJKyLYHXamX1Ga1gyWKrxH0Svmsh0VIOAm2Dx1SqQHv/CFEYUd/udmJzvK7DtAhUIoU
IUQYRzcOxnZtuVxNvEZDC0DstFyfg/E9epuNlWlh24fP6E20sNkCj0Xo0NIZKwxB0UhoUK+dAl+t
Ypey1NoXnLllHCGclgOME2MeNgD+d0eyqQH+FPiXCBBnJ81C63XR/1m8hJMYu6P99AiIMCFli/OJ
xokvaWJfmymyabUlGDIZhFKWWMHR3/VwbNA38K0vrUU3XzoJ10sDswTDMr/KnHmIcIX4ng8ye3KO
F/ccCQXNY+lbLaEUOoSOKONIEKv8xZzqvMWkg0ryMWDp+U5t3hAdn0vd4ACihizL4x5+V4bZCxQR
14zLEEx44MW09jMD5fuvWCA4Mo+r8E7Op9HLV3yEVFV9nmb19hBoR8ufBPie1mUU4u9ao7LyT3Yi
lTwxji6ZAmRdA5c+KBO1i+D+BVjNV34e7mcpaO2cPyMjOgXutZbWZY+911AfLY/S5aT1OjCHi/ai
gC8ACFbEisO6CqVttUiG9bxU3dcQTNl46M/iFFkonKeGQ3OQuBcecPKIOwUaWAo+mHjATd2IUiJA
j3PXumCHGpyMOsc9ufkyW8LOCrlXk0R/8mGqdMWYbrqG7iRAf9dMR91FgOJBhUGGbDQX/mKUWGiz
+sY5t8jdsulhPrQv6Ozsk5QIiXtuWPkH4GoVOyigDc+8f6E5/FWGXtmkMpEZjFwt9nm12KaQwcuZ
pJqokO0PvfH+uS2SHTQrmaDb155DwiR1Ql0uUSJ/adJHpdZX7DdWy+j3TLXVwwBJObY+oW14IPOr
/UKTeJDzRXRHaukIaBBLvI3/bngvSi6xHGOkNbdE2qCs39OEn+dOP0OM4SR+iUxAFh9kYsi388Lx
KCY6xEfuJpjjOQrkHPyQuPgE/DRIq+pryc8MSAQoxcy+LUGfvjArUT7ZpIzoxl5gibZtzBQlAQL9
y9WYaH8h34MPU1hn5xpX+wPv73z6mVQ5aGxUHcfWutWy4yfU2QvwV3P7sFWQc8HdkkQKZfdx2Hwf
3lLmKGJio13hh1gUyzb4hcFhXVmLCwNj42R2MGyabdZCYQlBuEQ4jFZBLDjxYiN8Rebm0y8Guy9/
hfQ73/qDCSJfbh10KRPoQI53AQUN7CJYOcrCg5rwr9GWK/SNuqY7NOqCaNUW2b/gOkR2zN/xNvkn
+0kboxQLJqw34W+ZptJYRxBYkKLyvKEJHTWBwxKCnMun5gkZiTIhCcJoujLeaYjyp3a9jXrD9Saq
C2N2/uqjm28qbKDNoNgMrGI0NES/3gol3wI9VbJ198t9kh85p+Rf+d167bdsnWH9TpOKZbmSi1m3
KKbfz5+O4UU5bg8GJ/HFRKh9ssdGp1L/6CsSR3pyrUC2P7S/kfXohNfY3wRs9tHuz4JOLrhiZFOv
MFaUmArH/kBQjHykeR8gBK//i4sqJK9gpDDVGAUfm/l7MXJJESxmKB8ZjXEqwXpwH56JoTUfTDJE
aIGSSCznsNG/yBVih4mxy3Ot0s3Y0tEOGHiVaseK6SIqeGGpWIR3NI3nAUpbhV0IKIIY52Llc9Qg
wQ9fq9r5gKGnjGGlmGqH7mnZv3XQJyc/a1L83/GkE/92JKHGdVf8CtOiecLni8zXKEGielbqn8fK
WDvvOzfXm9uE/kp+FpFHatRqu4MiqmXPn4mxVDq8VTUrTNczAmKrpEz/PKB9W1vKp4TVKi5dJVNi
P1NWx6vNifgImJ3xFgW4YM1/PJ9NVcFL6SHMYbPpZUFqJWep+8/EIxcMxiIprgFMzccsGGMfg0Xx
MgxjyVJ1KWz/C+QLEAhTLsZIVb2bkPx+/2RhqzPT7/Cx1wWhZzms+fEQ/ADMkOdHJeFz4XRoCcF9
9CGmitDt5rhXY9lbeNyHz3qDdMrWJFvQzec5SN+4kJxbBJkDX3yKxgpnpTq86EeJfxzw8F1IIRKk
W3quTRf15HfovLLXzyDdxYqKsdLcE5DpPa1w8oFqQoxBrHTEdWpzsaPxj2lXKOS2lPWVW7ybaonV
iPWLyE+QaPND92rUn84PCJ5lZC6RsuPq+X4WF9Y6DARBIWX2eQ6WrvbNxyAFsip1+fUdlm5IQ4vc
ynCP21UFUgJV8jOHYOMFLnbyHHQZWUtMH0P9/uccZPHlDiRXIoEIFT0eoD2HzvePsE+zQsuuYgJP
ir9r5hoUNmLVMnnPNkRQMwaElc01u7vTi0mkn2xUziZfBTnHeHoS2odX5BOcukyBnE6hiXtbb9P4
RgCT+qdlshQjdlqlAZfFAVUyIIdKD/cV49GplgpCh/otJX88Clq3pKAfKAzAjmJRpkePW0kNUPvs
TCJHbTdaKrjOxRCqH+2bcQbz+mAHsDRVIJ+j+YeBvPdkL+6pHLqcsRm/QuViD8o9Ow5EBvXN3SD6
GMD6Ch9uXW0LVNjccVziMDINNM0u0bzj3h7c2K/DXbq5DvrrlcxrdDPv23isSKcF4b/mFWzBYszm
+mAzYwLTB3faWYpDTdMSADkByjJ0OIPb59UmKVYCAU7fPWzWLzFE5hM07R7BJoyTdvIEdzlwMAvh
TdirFxwWC7rDkNrn8xUySujJJXMT+D2RUSCbggR9K1KifW46DgHEKX2HGhW0pribSRpOkuiXtpUB
sPtqYZ5Yy4KUsc0nZUJlM2WkRHmmy7akETbS/PHx3MHXKXKx/uNyTvWZMPd3iuZKZHbbwJLKmEfm
HQ7JYyJLA3J8Qeed78BbaKmeavbGTH17fmrK8Y8pcIETJubfgXqXWk8mbDU3/8ya6cjncOvDw5tY
GaWwjlYQIXaMoa9xi53LyZ7RP6fxGAe1CHO5sQJjkFfuS/XLAaLvNv/09xBC7uWehVE37uz1Hw76
eMz0V1ZGJcQaEReSCFRDppR9AAu4217DjSLsT9Lkfbqt0x2MaBHGk1HFDmOG6empGBK6Cvgqu7mu
1g/tR1M/vzv4Ma6s+VHOgG2YtuLCJrMelBY5jJK/73WAD8A5fTDWAwyKaKADRgq0SjyjWmsnKyfK
BaNbFXQF/fiabkf+OC+zEsrrlapeTQbV42orny0f4GeMkcUCVQgDkBdbXOwx93BHFtp9o7BnzxEq
ypW24jJoreP3hr573wvzxt0//pg5nKylsQEsKh9wo5TElNYd2GLV+17WiAfRfoO2TXKj2pYGrQDS
hOArsZQTE7FYFwFGbtZfr8H9W3odzFiViokmGCAqnt1ZIbzQjeuEQrlQt+vFtVMBFiGMSCexdG/P
yA3btcDdHt9AXBnMHvPfmBVZumrJo6EzdTBxUEWIWOoAvmkRfhZ6iI8r6fxe7OARof0NfxJT+Yh8
obc4qFjaOUbHIg51E0E5GGHzuQAeQOXzMmZj1FugeqO6i06+x8qUsKUWr3j5wdtadwGhZGbSbD4e
c+b2siGC2FMQrGdPPM1vAmfLV47wxRb+AHyVHA4TMiTmPsHTrcYdBqNotMsv24TKeYlK4yILSqKX
uFEV3Lbso4Hkv9cAp1DFA3gATuPhk+2ZfzG7VSLgg7Al2bY2LAGYa3Rt+5a0vnSue5jhGh498E7j
e0RaKruvG+D2G860DLeMjw6FiJqFophQw9Vqsgb2cIOul7o6fDWa6So0oDk+udzrvFonchFkAPow
OVADhpggP/cLECclq28JYd+ve+07B6NjNlaV4vw9ideBM8VoVQ8JyluubxsGnf6DL8lHbBwKa5ca
GabQ9uUh7a81/Z2rcoanmAYZXxg4E/MJ5s3s54q8b5XQ/KfMXnHTDniUMMRtS6tCUjzf64+aaibu
+nJ3f4uJBqqXZASecAF9DLu9VFNNU9xZ5oi9eaflxQLP36rVh1fIt9F0+g0k7+ZJu2jmV+gWm8MS
3iA1lk32ShW3XfxGBYMspo7fVnfX17LuUm4l1Qa8HCmRabBQ+kLa/bBAHZW/h/qMj2cpHi1VoN4p
cAc+SJVku98qRcn9/jhyOWFa8DzYvnDT+BvhNYSluYqo2Nt9S3l/OYACLNwD+HB3MJuO6jhVh1ad
eNvcrncf49253pOgu6yce42Zz7Wmee2DkRTLzPdGsZBYm+e2XGumVOncvBLXnNf2cWEMEUWrZG+U
PbkFpCGNxGVc62rTO4bYnTONC7NZ2S+ZqIHtpffMmfukhLWJ6+Tj3FFLvkzZGu/xL4HAY3Xvx9dm
V4WIou3XfSrVG9tLrkrPKlk0aXcEjHIubyx/UQUcrfdVbHR7ADFM5jPjK9st+liaXEBQniL9VOiC
ZNkpadPKpONBfSbmgzTLatOxw/uvSQAEelWiPWWZm/Q1j83u6hl1GdJ9FBoOCRX5DQo7sXFJXycK
XEZYmgAbedWwfiEQsvMx8XEcL3wbb2imdUq7KYe5SYvKjVDpe6yaNqAdu15Dn45YRCPbUmWXAtIv
3wiOOYCaWEYQ6vX3UMji3vvUG/Oe/NDOSsCEU93BiwLxh/nfQuCBHKiFSPLD2P91a97daEB8L15J
2whfs+5PMeoxjv25TpfD4tCyp7xrPyPs2flFE0RtkkuFseujbsCdnSoWyBCWxHDh6gNWNXSR4Hl6
w42wbxZQUVk8zvDgieHlb7JlJZr8Cpp0df2/+wkluDq3liZyz4v/is9a/VfijqcUBHd640KNpjpd
6UxQz/BArQWCypBBWghMqdrlvl4nPbL2YJdvv+AmeuilpOA05ov+h3Qjd13UDi2Id9TEDFMpXLEy
CieaZG+inQJTojde7LUFh/VReKMEFiYQXaEyjT2RaXmwexXd8fc4Y0Is3hOlm2E2xz9X6HlzG7LP
U9045pms2OcsFLyeDuR/C+n0VBiXJKZtf49uEF1nkQZn5N3/Y/3fxY6iRnp6ZThvfy1nnbFSAhPF
6npNBwEtSjeCO54Bv7ymbZecKkKbnEHN29/U6zVDY2nEVpjBO/afTX8U7qKqOcqRldtK9yWs1Ulc
Z2io4fCfoS6nBP1fXDnk4iH4uGr9URkuRBdldaFq/XHLqA7WlhrptRHF/JqgJQ4FLMp0K9PVoMdJ
dBrlLgqr0cvnMVeKmMVZHZ1KzBRMHrSo0GWqWSvM4J7alPpgkxw+5GH7ql2np5JUpwOOPr7qQ0/7
Oh7zA02rTjn5784bid1v1UzFWB1tc216cH5Ad0q3LEbaPt3Div1w9l/R6VydeOY8hwawi024hauT
xK1qGYQcdw1P99Bys4oq2z8p1zUIYg0usLwZqaOv52pbq9IDptUltA0yosUQCoI3/g7DzPPNFC9H
xuOubhqYFizO21cZqpZetzvbWIa6ywcFOvah+c4Aihk8CiYuW0itCaIC+x28UNbaAS5WUs+NG/cj
LqAUXTW6hsnXFG0oESe1Dh/hQTOJvfl0v+FyI8XsEqRc5CYbiHrwXw2k88PncKsbP3XR1pVFn872
3mRgBnO6T/xl4Xt4MUXQDfhi/dRCo/zxC42pwaEBoYmoZkXDYb+8arMONxQv+svNvEiRvWCn4Q6v
SMJTb8lJ9Md4M29141mSR5cku0DvnicSbuOljeTJLx6cpYluJPhka7vF7O4WfKbuKDQK0Ll42lWq
qcRDSN8/Hi+nSEUZxLjdhr5t3i8Iw0dmaRSEoI1+Homnk155Ut46hMDhPAQpHg7n9h72NO0Z8pwx
2mXrP9TGj6eE5ceWfiZOwMBSKnLEpiEct3qIBRaM7S5T5wrOolxliwSDJCO75/JECIBjvtmCk7a9
lEle/DWJZWn0KERAx5YQj/1c/09WCDqkKrE2LbkCzuX2kw2T1geVgRvW4bsV4DShzWqKBQBlisfm
fVrRcd16M37UlVOAhOntEBL6qP2B75MEbLxODgJaOUi/28boF93n/1HgYo4ajv5H+iJqnA3yGgVs
TfOa1ebgRRCpSdv6YztRH3Za97kbFA4QGgvP6Ek3dNjbZbYaTXbK58PVJWo7kNGRzuoy8UcrE0yq
SYOvPabxXG1gz75dGRWIDP/8CAuZ1vyEmTSa+N2RBc7QK2lF92so6+3Ubfej7cZSYT/YHSshdM9E
ms8hnTUhJK+2aL8zF5E4ooBngj3b/qOKPnLrZCB8kNyohaoKeGYlKGx5o/kaaqQVcrtSiurstq/l
Ejtv51V8Bu0Twx1lWzyKzvyOc3JF9EZGl7NUdiGUAvy2Wocg2QIsTUU+mTLOv/BgiHcBXvU07ENE
ww7imXzwBZ7wNXMWfNUa98mwEr9WQ1OIdKfYKICxIH15tZJ+9j1pndlZ6EbukboI6Loi+pNoPWPm
qVANTvCpGUFprEuB7qafuu6wTGSLfCH0HwNMdWO/vVH8uj+kSrn6OLV8MzuCiroEDVSV+kmFD6LT
sM/FgFiBd2J/sf6ZdBHbi0i0bOasUfJ88dGH30rX95ocnrtEzZLod0oCMNXizXUpDLPyfDfmsPcz
LWOgFhQr9H7ztcYGaNbpvSzkVD+NsBd1ouTPJ3CkIsqmT6g0YyEn4uR6ri4uKSye2AAB3OWO2aV/
FhBj6GLTRoAIVvt9Jl02uHqK2w2WG8AgzD2FoOcqm+a381wuaqJWdC7ORRqq8apWLZBx1L3aJoZK
Q8QuqZ7QG2rVV9wo86Eeex4xrGSzmGgk21IyfcECxKsQ9pKSEVEMk71/dcqHc9qD5slZE1SORiyJ
DdqBA4YPRv2PSq5KXXETE37EayQlEjVlSpgdxVEaP8qIK3BnWqS12KCnEHOjXxO3mffO/Lqc4ufF
1XM5VYWE2mNbjZUbn+J3Ti3FfK1KTr93UezJUB8Fsk/1AoKFpiIatlPquj9d2B2dTg7Kmos6TQ0B
M9bi43Kb/TliGQbd9b78q4WIHdbr35dxj7cnOl0uKMGAmJP4uWbtIbks8vtvdpryWYXdakcQeG5o
Mb0elrvZLJ8je2BUVqou+6FaEmmwkjlLOgvugr7rw2N0wnB/RD2x+asmfWFwrcLj9AAJ7BQrp17z
QPFjVbcG/YOI131sJXvM6iU35KiFdfTuPUtBUaUGV01plQxaWhEIq98GauD00dqErb6a0Jn4Ux7p
Wt8tdFG7owhdCzhMCYPJE+dlQCg8ecosLxcN7HwE0rDwHhM/T6qgF95k886BRr7lHBrTuHqU3mrU
U32U9aYlQF1hvZ3vGy0zHyQtYXeKFavBDZ+wDeUyfF28P0fK1qD4vkYUChg0eI7Ko7geOg5XgzYW
los7roUNARmMfbXSRsXKrQm4h77UlRnIA/Ivkfe4odI11OFV4hn740orzNgYaLW04x/x9uZhLxWv
UOsx7PGsASAuCMmQgW06kJt1shIiTHrp3rALQvcdvTzv+pcmOuB/vzeRQHikGeNAlVK3sFRxJrvP
KnGTuB6cb2qEKNIhHUTx02BNOECwz/doGODpt3OfBoy23+wo5MAiZsWwjnwiialqchd+K0GN9LIO
4G/RS+xxAIT7qcXn/zu3f0vZj1mDZvlF/VZgIZT+6igfsPaRuseMvlnbOXv3aADJO7/J099HuMlD
2ZLGcQfPT/jqIeYTcqXR+IQNhReDbd43CrAC7yyfJ0LgCdWZg0Xtv8Jm7AQ7WnrEh7Cz57jWtlDn
c2FI87vNRvLOYN6bFSWq3iARUq7BYHdQSIare8azqtTH+LdZ5e77f3gG8lQIRegpCdXH1CCADXzk
HOlQdOXj4ppL8b8CQB4nIkaBdZTYGxIlQpBK4aq3Jn8Rgg0i7uRPGl2n/CDCPwU1+uQgASzsqsG2
OevdtX3Fn588TAlJdI8OHaYXBtkZSnZxZd0x2afE0DDGmWyivchUBAoru9NM8+d0nH3TBAc/MU53
uVyePwE7qaiOs1GICGu2Ip2Ea9f+X7blxzMhU7yZPuIx8J75xZR9hGyJq4HLO5bK06pbwvlo489L
1cLax0558jtnYwwl03ZdGxAy+QhmIXvDYBjj9+a/9qmbd8JpmihhjqNYQKrFJAKdZrGjL1dxj5Dw
3bdXT9vE5KmS1Jlr1ubHqC8rvnBO15GYqOWg5lNln/i3ff0bdIIxKUlecKahEhFJFD67Eq9z8r+g
pexaa04QYaMv0YylNBptZ0lBSCqaijQaKIjtMPVc9haeRmGL9RTWvvl7aBcW1LGEyBPDpCa2lWcX
4GGBOPExBDfP1BjVVnqFzoaLjXCOUz9bfqmPYlUHkIkN+TjE/rfgRMN94yV0XA7Hl2hTF3B1TBBO
PFG1SgEFx3ySVSqWHt8VN+RQrEGtRHpKfJh20IyK9OlOuE30uPs1CCGBtZyL9d0y5cvJA/G+ns9P
YZ5a7ZemrHBR107rPu90bGEwh0P0Lm/2c5JuwrjzFMo1F2RbA/t/YIDgQe5qououwWs4gYK6BKy4
hcd7dbXE0inL72Syx34cIStu7dpbj+NKdPzeUpVGzr3BKVFUfS9TOS7jFxxP5YbrKAYZ6SDo6pQU
yVbc1zfUPdaNHkohhwdD5b2cFzURZkdxUE3rfegzaK3OlGPgBsOYm61rfOKXGJhB7oIYX7tJkJVi
pOO2voCQ0BY8YHYlwHg5qlfwDqfk7PU9fQ4iTlP/t0Rf7wsIs285A/Ohd9NvCTgFK2SJUXBI9AJE
2jj8cTlo0iDjmzr6KgJyfWq8Dyx4wmerDkWPo+Ea7GaHMixLecbdmlaW6O/iA69o9kHQy/j9tGJD
/kHbofOI0ugzsRTv6Q0AdkrVg3szrsNuAryNaTpwc4C5AR6774dtEhqDhyQn+GeCAV/l2/QZ65lB
0WUPG0BqicD5bitVLMbXmqgPEnpB1aALxRde1zpxv1H8gDzrsSQWctN0NmgaAKqVtiRai/rD0csD
1sEvM6QHnTpmb/rL9AldpkOpXaBOdw2osns+zhnazg7IeG1ITR/fSQhm0et4giqM9e0Cj+ctB68V
yF57l8AFTAl4mElMx3/4qKg5is4Y3vx+uHV6xZ7XoqvW7hliaKsCFy3vnVz73XLg4BG/OaciLJdB
5XCZIcODjqzJZVrESxTm9uZg8ZkpCydrxJYyZlwQbibErSVXy4VQM1YCMKR1+5UOoStzMbJKfEaW
QPlNIV27w4xT7yLDtgMnvMei1zO7YJh4q4O/y35p9p8tRT2oO5qXCDuJHpCw6wWzypzonQXy7DqM
jeC4NMfwT1Q/3ZTQub78tY8jfHIazuN53gNNYvV4h/T93sIXH+wnnEDOlf8lI0D1gRbOstaKLFhR
A/UKn45kW3IxjxnWPdU7xcn4+mnbCRwjCnxoP8bfcT+JF+fHNYE8XY/UUNtpK6VNIYVDIax/81on
HRTGwuZZh2iprmun1hEIPu1OPHbHm4KZm5aFxp/aj46QtxRBQI/PlZLIEXFzXpbF5baQP3dA0Hv6
bxqavCbL5FdQWKazQNfKPcgQnewM0FdNAU5khcB6c06LKpR8YufjhLi58ux4MCJwo0Q5xL/S6+V2
1k+0TO4K+Tk36Mq0m5Zdhqwg41EcksIsFYcn7AYSmjUKlLQ+Xd6Q4AS2SOKHEXRzGcXwfInhlFpd
HRt8CTT00XiuuOaci2Abd5iTl4aEmHSHtVNMQXY99fyRd43RyoivwFURKZf9+vqR553TRoOpSHkD
O4npkvaYe7A1FqbdtTSv36fwEIvLiE+Xi9Z+SZ3WCrvL2TwBKdaf0uP1w4ZeIIjq+ttMuA4t/R44
zYJ2y7VmJOs+rq4zW5gYCl2OZcBOFy2m2+fwf5oubqa1HI4OriPnZnzlXGfY7zFGc99s+A7D0YkQ
3uto3FbPNjf4NAr0P09VaRVPJuPcDGIVWiMJIvjLCQkbHuWWN6qyiQ0xEktc5pAvOVfvI7WCUadZ
YrtG4itHfhNoRBU6Reqx+xFfFEioUO9c2ZeGUmk0coUpnwOsYTHzjIbiytZE4+RWtA8rvY21X7SE
T6OOp3Sr3pOVKZFmsXRU1S4hwEVngj10DH3Zk3sLm0wdQHhdjriyX/4drk+Rcwj/7uEzz2KPJ3hN
Z9yjtkeUbdoW8h0R1xVg9gc/lX5K1jmK1y75E18nQWg5lczcCpJwOTJU7fJc62DI4KqGmtSraGQx
VUhnRm4MXMt6IBWDDbYrg4RjzLdUWHU9/qHWyleVqA6LxSGqSIuOBOIVeVDb5PSEBqU0tG3j1BSD
NpZuxsKWt3UhoQgstTzdEZtjVm+d0YU6DQOaTdNhdus8gbnyxPiXzW6/geKL1N2bVyMOl9N6mYrZ
xxKWMu/boh71xYqvuzLjM4F2VxDZc9S/TgS+I4RMjLDWW2vdN+rj/ZuF/VNRY1K5PYZAYwjsrdjM
NAMfIDOxhMqfiLNhZvopcyRZtf90LUHzuKDYCsNBh+em1uYi6c/5J5nTaRVPBuf+m9OL2XtG90tQ
DAA/474mttKcAM59hKE6v5xWlw9gLZR5/6PnnH3L4jkvEfpufjhcxa+77SJrcSIue1PRjoB9mDrk
nWMV4Ft8k4PdVINTmQrnggv7+S5WnH2bpJ5BhL51utzbMYa9UsQONjxNm9IXkSRQDDKO87Bk39i5
80qjpjFBfd4a3eH0XuKVb9GpsZSOUjYJNkZUdUpJrphFRXMAZO7cDUf8sbT3DXS779tiLRZ0Bymi
HS36B8I/XrPotihdFfbeZMS+RDPCCVdwy613Qoxx6d2dmuncDxVxDB5UgITg9Y9llbpWDsEc1VKb
DFn5BdilX7Pw7obxjjHVPqLWq3U01oYIN8xJcdsfi41arB3hpCQIInHCdcHGlqmbniuY1nwhpySk
ZboyKqPDg38p0QtYWcSH4iE0Gvo3M7LzQHr6HscUP6KCM5DPFfXrXi/opXq4tnFfpq+vAXunlTck
qeFNN4OjXwKmL3qyVuYwOK+6c2wN0hUfbLQhyEQfajXzPXhdkFDzI2j12Y53IKM+CTj4Mlt62EIV
P/GUKosjZhEJUqKnUwq+q2teLPF7iIEyO1eH09rsSHvKXco923UZqL4TxcZAYzfD4W1tCUWAiies
DfjkikrMy/1p958sQ6cqZ/7zPOD1r+GJ4wSCW1Jbw64ElC+NRBSoO5LWL0f4sUKDQpMo353MQLtf
wSE5Tu2cl1SNdQsoZq9NjpWm/pR3hGLvHmYplz92MfwYhwcNnwM0yyT/hWmSnplMWllzzJNHZrME
w65kUcxKwlijtG01qJH8SBBRIK2zISePqnNczjyh+H+k5Z6ocjX7skULxzhjx1O6OZTmu0c4/0YN
nEVqgCxJLWu/06/3v9Fsc+rLMeXYV4AAkLrzRUoTAj3Qi76wVU1mdbUWigryyGeeB8XzB92soNKK
yk29RjOWgjpgui/9lg+P5jNEHyn7couQ5ujo1F2s0V6QW19D0EiDJRqNs4+vCdWr7jOxSAOStz9Y
QIdNWQ1OSW5LTpmch8zDYiPi3P5JoErRDGOx8N5h+Qj7MZhF3sDvb7G86wMcfiVfFpAWRsYCnuUV
dnEJTggWXZzmgcVMNGgXhkl27VkTXyp3moDhPlGW8MzYc1ejGezJisb+0tPCJtJWsuo2qhJYcF7s
GypzM0wGc4YWywK2MPIVjUs7fwEbGRnFCRBOetlIcsHa73Ij0Mjqwko9uJ08srzhGF8gU1LIsTPt
C3OwRkdkop6MK2pZHjaLc/8Axl2zct53NnVEC1dqya1KF43HuhaVB17MMiyM5pRaX/YBie45V31N
eh5rkw/2fjI8CX/XTUAIC29qyOxqLpDMDERTTw1KFLP6VrNkWrmv6kc7TWUytPC4JHZy9jrDsg+N
UE2bf45tsdGCUU0/8Rk/othPuePbcCcrjaPkKDNmQFudYCutPJQvwlLBEZ4DeoQKxNTXdtVHBvsW
nrm4hk1Wf4OIUcSunTZlbVFyZjvVKhNZSnKH+Pf7nstRe7EDuFzHWrrJV/L2u5AkJSMAhaOWzRHe
Qjrcf1+h4Ff0ODzqdpCaXxxqj684eZutDBYR6A1PM7p0OCtGUduUHCi0qWINw+bO0NT2+dxYwm1A
CLcDfUzzgLLMat4VbFVxqqsX0NQLIptL3GAARPZ2uUBVm6TE0N7ialyXcxtva+V/7ylE9jMB4m4b
U1+Dmuy4xYPDArVvv9wmtERYzhsIXwZ5ITHHJgPQE1eqop4YJaatmxUAzDsYCFgjmZCGqVnbwPEK
cmQCeIsKV4AVawxw7+2em9x0FOZ+CNYeEOD0wqZv5I6yqrXPh4V4n63M6DO/K2xM8GY7jwDc/NIl
uhCCqOcjpTHXOFZbvr1P5tGolGJ7IvkOVnc/QfQLNXXelUkwOVn1cXvibkdQWIo7mtSBs6zB7uc6
ZU+Y4LEQtGisgf34Lfg0I6Frl4yci6B4R2YiIF1ng2q3mO3IVQK7P5Jc/4AZPgzYoIZ6d567txGH
mrl/+C7pXGuLDCLB5F4FKFHwo4qYdvsqPYHAbpgSaexCyO3Yr9LxiiUtuCi2uTGP6XnIi2V3WU9D
UysvbVAie8xLBqrXPOT3JJk+Zs13WA1T4fkgIBAWczuiUjX9aY0ucr9trgS7SJK8EiFAPpSVJBmU
Ud1FXrTlWbvpoebX+eY9iPdRg17M8DpnhGAQ3Je3AKB0DKkVqrLCjDgu6qjLmkndClANwGUURTmd
hSzy5iINTQn5PCfz05W3t0Zks/SLEkhwqpGksWsCW2xiAlPVmOe3R+Jxcg5dvEoceKMNAQSuG6/B
jLXRJ+slwEmaead7HLt/sUYDphvUzdskhvEEpfGEN583OZZ49Yg15lVLTggKyp/JY1kyZK+vNDPM
BF7FokmEAORik0AOxmfVfiizae3IWdZfIws6QreRZv0u0dGl0KrkP2vMUzz9Vp2+gzlp8cy3l09T
DTq5GTeVaJ3biOP8zfRbjGylDGgIPQL2Hp1bWOitwzUGKeWFmb1/M6adDffLaHLheSAJvx9gm9LQ
4I0ewzHFWAg4sTMqwV65+sPX3VDaKVqJ/B5kT9jsr+u/dsmy6aSW8ZtfIonjLvMtfp3bnaGPTP0I
iz020PBP6wqn9BjT1Hzr/riBJNVzdHji5P6Nhe9Bbh10gu8RxPbJzWiROc+8Af0vQP3Sxda4uteB
qfQ2ZXMp6EdgxVEVodT9L5Z7O3iVdL7Um2RECbVvwgEJZmKtORVZnebiR3Dp/G3K/sZtowRqKusC
5rZSOScyH0/i4fbCJBiW7k2p6JSGtxAjMu9C576MoC6lFPg9PYkfrSMvTpBCCj1bCIqIvAzMFVhc
tzlLZgdjXSZRrhyHEoqEq2zMSRzO+Ybk1fhLlL5ZBh8ANzzrlL0hL2CtmwsorbfutFcmSbeyA0Lp
4YYe79eACK7F9bQSM6ctb6G0OeZVhNA04G9Iv6W6gXKrzA5GPUsiaN5phg/WW3zCs8J16A4ep1a2
21XCwtP/xJe8eAT1w7uGsh97eNPeGr8lb/5awXeMENzrf4YVXlWPbR8D9hZEsBKqeqDDA6jwV0Xs
eLiE4h9gXxOoKCeGYUVuww7V54xGWRwYbRUGqmE8g29ivtspldlmTQc1IQnFYjCqRMk5IvxTLxsE
P41PWGpMBSvryVhDTDXQVhGPVWZgVGZxfw+QAe8eayTNwWF9RxhYTglRWRS0Pzrm/y8nkCTlZXqT
68aQ2WGS3L8XWCJmmr/YJuben99/MWlBMNOF4khPNQY9z2kYzvQ7EFvXimG+PAqhOsgaUHpFzV28
BoZR7h8M5jDstjXjmxFgWe+I8JjXsEUs4QlEPVVzeLVhBkLx4Q45Fsa9abU6CbEbHpRZBcp8K0Kq
T8v9H9bFj7EB96afaMfHypTMedh8jXaxIRqRcPZV9dnzrpJHZ56sn7gRdWh1C+VIhYO6DkZMHF6A
U9cRscU0xBh8EfrVH23UCM4+ZiRclkxrfJiQx563AEeu1/N5HdjCr9e0RWpjsev/McSGjE6cmgD/
wmR+VIuENH1SitwnsekydBHdGqXIrnrdGtVzHOq9yIqnCHOsFCgCML7k4d8iKgPO0HmLtGqjJUrR
UgGnvqSZI0gkVSXrQ/B8Nw1mdY2XzC5nFmlKFYSMmNwzUaVF7ZrX4PbpXFHSWcaKsUbKyKq4bwi5
3l6tcMPlFnhcpxtLt+1nwv7Vy1+PmQkIbbXtVQkgAEp1t+9jjYFLz3MVpMSBIvJnTtb502hf0IEU
0gqNbdf4qracdp3Cg9ualZ5I3ZgI8PnuMWyYoHoiIcFD7aQtnE+M4cnxVzCHBN697PJKTYG32NA4
PX/0DKnj2OlQHJEqLGCwkPjNDfpjNDBMTKMiLiW4WKyqeuB4dXrdbzU/fGa9k+9xgVLaiKwAy64X
RCQdsdRL964oEeTdTBozCfdPdr6v2L5o3SWYkRtAOCES+rizrRHIN8TpJhf6w2AhOW6uhDtKWbKq
FV46PqKVzOrToKDOxDKEKcTp8MIrxt9CeT0ErHl5CJOtE3fXO74mienIPTnjqbDE5QjC49RNKjlE
Utbl9QHQ0HUGe5fiu51P7YAk0Sgrk4kBUp1wCNXrKTzkJv1cbnCpHZwWA5hpg8iDOE5YWiIXMZdU
jD9xPkNeqslSzg7yJnw/A4pzRdUO8DdzpRdBl/X6dVMn7V33vSv+07IQZnrSjw1XxoUDv6z5/f5Z
m08iL6b3itLrFwbjeI1hkjqPMTcZu30rjbJ15OWR11aOKgQiWrOZ2XEkT1xfqBcm1K/+BeCSDVzP
9qsQTu49wI3SunGp+hTCZ8oLl3r4Z047AH/MPsyQ82tOzXanjEPSKbb/VOCjq1z29lizat1xp1iR
44KIy73+B6+ts7h4PUpw/KKG0PF0JtQnFryCuMdxudIWWbZaarE2CTUOiuTQI3fhTOxjzIJgcsPv
JlLvYklGxZ4Sp5xkNqSZrKbTIMdqBoXuwlkDV7/rQqKIxsyUkeKYQY7HZSPx7Cbrj3jJSpLLjaz/
1RQQm3wyIG/VvbcZFf813VW9AHTXX2vrGwc051l3Wkk1jj7dmaU0LB+1Kzf6g77pvpk9Ns/MeuGY
UznG4w/DucFJ1XqxWgCh3Z/asFcrsbUiSVJcHgZFxz8mGxnExeJBLcz7UqqvoRvohJqJjV0vAYVG
/skho3f3qvl0yDMD3xa9WJ2Wlloe3Ic//c4dFWlQFeFlE6uiPswvQyKMiR7SaK1cVvO+JAuPtYFH
ToYGE7sk5WQaHr7jw/bGHMRytSRPBM+bb0QKEyeTL9KPQshDfxtXUneHhwcd6uXzwDAYNkBJ8c40
UpDFQGSryVw3XY7Gu/Ae6kXb45T0YAVtUXMtQbinYTA/2tZN4xFz6gZiakljUWqfk1MRkX6HiMZh
Qq/xZ1wuCZMWwqMWNmQKIXP0X1MrsiKqeHjfsd4nOKwt2EuROgLyurh+H2kslPLdcaK+lAUQitl4
Ukvu2VG/CLiCw1hNRNjhP77uosisLeNg9EbroyzTMlQ9U5Eof7MU1hJZil90y5Kd1iW0Bgt2Xz9B
T0W1iPE/oqePGYvRcuSnmSTJqoA7PqsemcgCPQB19zJSOvDYGD6xx9sI0TvA2UiEJRXRHaVaV1FE
brhGJQpHpYj9fAeVuK+csBohYKRxHtpXzhR1NozxHnNPUC9gOINLTAXTCy+OAgEuJqnqtqNPiHuB
updOyyN3gVFP2kK3lWAgFbJj+iq3RnRmOWPaofamTbfKwLoxikBWayhUSPQc6OxgxwWwFyE37T9X
V+2cmslH/8O3Ljmw5ksBvm0wOgpp5vC5FSO+Kyc9W+lUGw3m57YL90pL3g9e0JEDmtrnoh9HCTNs
qVvrhCbdAGO/OsncCNl8dnjY+S4ytigDTeWbRfVTX6CHXPb2pUFzk/XgrdVqsVCtjx40iIKIXjs4
FcwChRDYMGHNF6rZ16xcAqnljlERoOCb001xm5l+KGwVMEE9S/1Bny6fB7DVsGtLhvK3vNPvPlKK
TN7xST2Id5RbDHMi6kn/686L1SONgCH0+gR+JUYa2F+U1Opg4mrFMgjW0N7frccCL3/trspGM44X
chWhnogAIKeWSQ60N80WD7b6V4wyHrjii+GjaZfLHRA18KXK/z9qVODUI2wPxwzGjt6mEvpX+5hj
ogZX3mbIoQpxBt1LJr0UTBjs9ZA0qJa2a3NSkFjOScbmq6rs2gMS18sFZ1Biy/vTMs1WlxhgrNBF
xMMnb4XZUCif9fDpyFFTl2e0jqJTJGTafbU9OVT9+t18McDRfhE1NNZlOflES/msr0SZwVD+wsou
HdSGyYP3yA1y0kBshD/9zYFY8amV7aOhDtmNQ6bukfL3yLNnv952GF/6zWM+ysf9XeQJf5VWay7y
yYr1B80YMMyKhX6XnD4sXbGhuCg4PWNjB1i6sR9DZs/vykoxVxzGe+TA2iSGcAEg7G1nmbxeT05J
gcvwJowINkYmjOtvVMn8DiusDcw5IQawTc8OIVpa0XxMhS6qPMQBrUBZBFKuH/iaJKnqthz/bt8G
Qzdz2wrdI9Q8svoBsZs3/MsHEO0ww4lSrTAIr/avlezWIDHArjW9HDc0qxngkjqc6a6JzYYwJB7D
bHEmlbId/d/1ns1AdECaY5ftvJnoIHCwdilsksj/xUGVwoQ2n/72O7k1xQUZnmMpYai7pwpkveDd
o/2avgBOwe2oW48HBRSkHQll6C8TYgiwO1pcz+mSGkIlvQ1CgomA1ExaQzUEsyXJk6vffdZEPNGU
kasN4qt4E71QNDdj4LRy7evmXQ3tRrpqBsZHnbcmRZSpN4NeX0gPe76EKZLuV7WdOMqVsUMZME8w
I4inFqotUvtDhlPK6vKjz9KkD4vgxqRfI44tJhkIv14Q+xxM8FvYp9O7qg66BUaX9tS3NSOfhEp8
szR1dIrIXLFIHUtpvO1cTFUqBH6qh9MrFWmHxomA5DKxocmb00o9lkgHc0LLwetG5co7rKbG4jCM
mBo52oTys+qZWZSXkzsKkE9HE6kfpt+fr/m0yDiY6dXeDLkF4IyxeFABvxgCyQfwXGhlgEiDPENd
pye4dUdCLsNd8UGe2RnQWWZFtzT5Ks/HWtuRGnlPdK+SAX/clYfLXQx+B8KgpnVuhPcR6TLk4nLZ
jXY0TWwTWf9hyfDH+3fpyBQqCYcKD5HiVqVnKT2/LTZmBWex2A05VUcRxHR+cyi0hWMayaMHPtGq
wYGGUaNLdgkFMrGwXkIrGRnYLJKEDqcyE0HdWd2HWz5bNhUTZgm3XN7Y3LVGgcEyUCdG1glDYwOC
8WmdegmcpM4a4lEK3mu2yIivsTKIjYlBn3ASWjGgS3+wOia0v0at21XsA/aaDw0sx9Fi/V9lWETy
q+iQymVtUi+mJ+mB+A4YLa8Kzbd7n5x71DX3U6YlnjydISSX3Xk5Yp92OjacnN9gA2n2V+lR1Sqw
lrDxLl7x++NDBPwA8nYFof8s1Pt4CIfbpDNoRndk5u1TFubrU26OwNsflno8if/usYi9bZs9b1K3
TRaZAZ371+JYpg045V5U9jCH8m2A74mWm1RmRlYWF5XjYQlzbjlaes9Fxl+2TfZTEXimzJQnAFBd
z07exWzQCwFeVEE73eV6MsOCZmnvl91zKWvqgHyUoTzm9uaeG96KtHhBJYPF23xSGWRGnwd+bjhc
+oHFOjM0UBKYjB4TXyNKCtEpjJ0HRvv3p2yT2+J7ndiYv3nf7wtCfP3xhSktaFFm4hH0wae0wxYn
mab3dCJnL8yNLozehxOiSp5f7CdeY1yh28LG/u9JM/feXzXHaiCYLmuemnjxkf2v83b77aCqag9j
q6l6UFzGnn7s/+CVsDDcLE8/b/NP3wPT4vrkYksaL6Ngp1d6i4CnSYT9qGZZjkQLYzJtic9TuHGK
jFd9WxSpsvSeL1IZ0WZee5je3fDexfcHg5gKliaNxm+A4GGIQqi0vl/Aoo6tLE9CYjtz+LieCqzq
LjgbTE23zkQHOJq6XWwuD7b4+/Xk215IwBvnrgxeJZfQsPCS19eGNjs9i65zpn71rHnlde+u1/y9
SgzCKg6nZL6QuoOFPL67RGe+MNj/SCMti9Urgl9TdCcH/uPHrtd+nXz90mzLfLrfA3YJUswtcTRI
MlPF41Fr/KBhq0+Lo8T0Gd6MQe9q1aX9TulxyCzjKH+kFuEzS5gbo687EUQ2YmkbhDh7HjjecoU+
JdE8kwIidbURDZdd4JzolbcH8MJmd6gwgddifC08iqHba7YwXeEqnk8UEZu++F8SwQOgVGGgm8jA
voMTtn2NT0WrtT2iEsa2zPelOlKy7mBV6QJNEMpflWLPiHH/ZQbYae1Lz1ZmwhL4Tn6f/uKfS1c4
VME5vsOQGshMi7E+OQKXVUaReB/ouLn2dpCSMbuvWdferEwhThoftljrBYWCUhNx0ISaRydcTr3w
1pLAQaelQinYG39hjjEGR6N6p2i3G9fgGQmoUYm5rCW3IPAVso5NUPGfWo9jIDqkR2NaN+8Q1UW3
FDseZZGYwvCM1+Pbeq6UCSOPI30Y+NhlVOXK30H3/clZcv95F/oDK/DuiGtPuz1ten70KWyyVPfs
pZmWBwU6/p93ODqr21hEI4wv1r/X1tWOTZOgVr1QPOrpy0mw5xNKe/MEUQl6ZBjYpPtKUtP5v6H9
B1c3du/cXbdK/ppNU2BqXqd9TdnctQPgIOTUy9waGSXOG3V24ozalHqM8quWaUSscQMz4gymNOcu
DevJHT+pTbHi19l0Z2z/doDoGlU7Ft3vNamnLnphPKosuAilNyMjYQgSg6Yn+Oop1ki9H3dz3JM3
eMB0Pc9iyzy+bi1LAxhxf6tNoopLyvYRR8R7eDToBpvZja+mWoaEGETjTEYcZ8wZsJYaWJ+yH7UY
FEPGnogdGtcvcnE9iv+XoRFQK7suiLCfmvjhQ+IY5MpQUSIPtZCSWBLCtR//60dT5nG7kcFYvzSL
UUDqMOC00Jm2P1mJktHbsgp7P9pnCvzt4hm9rs38Y0d4R8W4whl40fpzc8cMpSdoXtjEyw0vi1LY
XSBeFv/FkaeH5EWK1+ydV7F7yMH5D9C6e8mIaT2ZFRSKfa3XCUWujHmw+h+KclwhO2C5B+r6AiZB
v4GWTszoVxLy/MFoRVAMkWHhMsGorUSo+wWhHP8GSIqd0j513Md421pK64RGi3ii/GYIqHn49Sg/
2YLbA7lDYYdWa49rDEQx9efwUDGeYDPX2FBQbWgpzBojHG0r9h+j09d5B08nZCIOCO7wfLUdGJeI
gO/ySrr+Fr182H6u/8ujBQGawA/O3LWeEoY4rH6Vzy25Rh50DcqhyEsWw8PvsT/xQiMelqtphY2I
tIrmztPevIrOHDvsdW721ujI/80vLgbM4JHXHcqiw7w/YoNqnMHN0QDvcmsebUbpv+y694CelzfG
ctRchhL/qfcq/xzwTxbMKtRqBZoYc3PEWI755e5hSsC4QKvKlXVKh2lPPbG5SIhrKXycfNFuaGyT
K7Fm7+l8hb9kv2x985LocRyb34RcRo24ovdFKPL3U8hvLWjJ0sbo5PmX7cmIRM38VDtzIaXQaN9e
iMNYrfOVgzz+mz0A3YR5kql2vFFIitwAHOGEZU8zv+ZCuhLw8kMLqJrCdOZhWZEhg3BoR/bflH9i
daStShMio8ZwlV5bZCYrIrB8Ko0i7E8Fhc7IdLEjQncRmyyJH8h9htRM/e8NsU7IbLz2UIEeOuyz
fv5NPvfc01/TyIzfBOoMf2WgfmUyhlX0O7FThJCANY/ZvsGWpweXsleJ8Qx0wH7X+PS5iCPfCA/l
j/XzlNuYQZ3QAe1I4IvQ0cn8FfzM8oAXxYU8i2AAbGpla4J1yY552gBoi8QeeNI6AwWbkTrgE+VM
SzqonUtS//z03UzllGeWFVizl1HZwlM/dhb4tvnt3KYaohNeFBIe/6pe7Lvh4aWVbnW12w1aYLLB
5bP9+3ijC2V3UClReWrNmS9wTqH15PaL4WoyUsGAvcJBBs/pNOLQSY+u8UppGyKOsJNkwS727osU
ILi8j52lLEO1SudaBFMB5i1r6/50bXL4XnUWqJcgITh2U437q3k/2z1HQi8oUvNddYfoyRen+fRD
F0LC5zI5b+nAMOffQ6YBOiy80Y6xXSl8Gg2pwDXa2XiIXZDMFfS3Ajnx4Vy8XYxGPkDMCyqQHF2a
WcsrM6UiaUDNqEydWmQie3AHbqRKNsGabXYRrAyfROB7bIaCVl9B06wF4WlDB0L1RL6lVbNKdALt
qLF7BVXXzLdDp0gVAR5FyJENSWqNIr58EYlEHAvwm6Cb+e9jZZX9qwWkt28NZodDjdkxeiFOgq1O
Gh3+XGYA0P3P/zcFUqCVUfwvdFYa5nfJxgUuN/7Lb5DPqJLuBAd486IvkZLjdP4NOATsibwx7PV5
7nmgFMcUJ3Yp5D/Rn+mDHJun2dte1pzqqxLO4wdPLv4yFjkiPfC9DjKvTs0piRNMo5MFN50Qmmrf
xiX0R4ne2ImHDmAO+8lKDyZPtLWHYhdJaduZkQwKpL/xc2Agor+aaIgYAz1uMb8fPHSOGeRr4qOZ
rSLMkWbHPOzTSqM/mDhmz/858i3yIF8gNJLqer25NIXQ5oiFnBCDezFFQWEFhjC3FLniV05zFT/U
v0fQK3JZl5L4QZlqd8yfktZu95i85NX3mmbNuz4i16ZZ/M0IASRw0vsLukomM0s2SSTcNnLelnqI
UMlsEaGsJAbc6+EIJUfdxJBhyCYrNq9ErfK0JGOjqS1iDcs+r7xC2Ch0hCOY8zkRw81lEGlYU+J1
ZdMI/10jXQLY9DT26sy7BjJmPZVPIJn7BMfLP9pcLrSTr6hpmjoVzrfIBofQ0XEHHaslWh7xztoG
z0e5Q5J2Gv3py8jRu94m+ZJbrxJ4nk+wDNbvgM4osmTm4hlcSlMeRc1QGQ61NxpAFFZOv3tMHSwA
APDck5DvHOPc8d1T0gqrxfsBlR3vpQjL07mWTuMx22Spkjb40k3cw1QIZZXM0+CO611uCS7pjdnW
ai20Pykr9vvheNDAS2Ff2tBoVfnzZUFEf3Up0JbGqHugExuuUkn8uP80KMykFGr3SxNUokST2GNd
RimesBU7SBbYhGBziHHnVI88HEg70J7hDHMwCDTgXpn9+WhKyB9bffUl7hOCeZrNXRl+bcJB7hvt
8Om7ihkhrNfkYBvp8/uELkO+y25W8TxPUGwvAimU7dJSixlr3J2cmElNDEf6hd6JTkDxp0S4WltT
I93bkKiQaSbo4qOJ+6UFRcNwiFljFSXcT4uUmAJSShFkXx+0grSSGYerLKpAegiyzCpdEnx1937j
j2Sa1ww7lw1sUIkq55Bv5monl5Q/Sg60H5g+4d9mqQe0mkhPzLRooVbDr/rNWhWSF5wEQQrcHLu0
h8jpzQ/kJOKZBebuzv46GXwbARgQVI9TfxyLLy0V8UURcq9t93bFO3YPQBYMqFJ9F4UzfS7c1qLc
tKMUJvsRWzsktoEMpsEOm1/oigIVvxMTRTsxUWLfqspXDBLQOa9THHOadfCSxDKtvx7Mfqgyz4YL
ipmTd3auerZ0X3rldcB2E3Mf/1caw7Lq0dXKu0OYLDf4ydH2fUh5j8NvXduVv+eJsgdhJrDgNLRc
Ed/09XNdyFczXYMKq/z+smB50OOeqN8oyAZb1H4XrWJiupgIv5TGyYUmA/gIu5J1YrpyQKxv7jwg
knuohAt4smldJ/ahvHVKPhGnX2SApEPucJNcKmxGb97SW8it4cEQa/wMq6T5i9gdoRmcMgNOpFve
STNIKyz3FmPKRh+SOC7MGykI/zqUn7iAtYmKXIrqrQMcgrHFJSgfuV+SCa8bU9ysNfCE3uvpw9EB
PSpoN8v2BeqYKJ7wIwazN2bBKQC5ufsvm0n/EOVev2vOfJ89S93Le+JsLHF1nEjXDq4qE6vaGsm7
qagNFtHbs0J+pQqRbOQVNexJqrAtRq4OZ16CQUXzM4W+RGE/k51p9mGh+O3C/9M3BtwxFJ7JD64Q
za14F0QM0RRxoJbQYJskO5Grbk27z/5sHXGS7imAWPB2I9KnhQN06LtrVxMsU08vfO4fjQZ9JGJv
0j4XtW+ZsLvz8wS8+epMRszqYl4GAKYA11HDGdHP+HFHB8z4S/hC8kzuFyI9eJzY3VQJggEZNXaJ
s7Ldh4mbNG3bsftJpicB5zDPiS+z0r8mDFWsG+2tXfh9vlEvmJyFJxuzJXA0QgZ7zFwNP1tn5sLq
bd7EMb5l+Xr1ZLeGTbGUeQqQQlbAyrjykdxH6x54Iv9cCJO6FwDR/nmljOsdBQP1hNJ3TUR6AL2p
EPjorRFUSKPEYjz53Qo/aVkfgaEM/Qq/X05CNucKkJ3jc9cZPC9jL9mvdGj+vIjCoehM0R1/7iV9
85pk39KNfTda1RJGBNeW7JXto/vXkNj24GDre4sux27vVvq6RWmRomGmH3/z+oEwJkSizu548ed7
Wjux0s23Ii/vwtVERdtJ0MGYi8gxHCnAegiFFUN0xsuH/IxWZpkncOSqeM6/VMMsmxJG7+j4Ffbn
F1Wkm/9Z+FJ3bGOcZuKNJYa6Lbw8r3YNrUs6EbiA441ZAc3qOkbl03ebThlBs/ahLaZm3NYZmzTb
OsN+53OHMwDANLTh5thuA0LOzRqJdpTRZAKmeOVvoieB/cOI7TySmclbTouRTrrz5MJN5MbJL+VO
L09thN+jKpMrRz/P/edC+qHnK014dpYhG6VZ9qrRjctl4W/WTtwFWX7XHHwZeY6BvHKQwlomaFIb
Y3RnkglanpgwuLpBUtejw5vIpaxTz2SkvRMaAfpdMYxWpUp5P4ZMTAKeGydUXBOZI6t6tDMVnzS0
CPDUtj1ECsggq2wdwmg048ec3NaAr2r+L0fezhYgyJln5zRT3KUUVLFecvDVSWEuc1tcAsKuuagf
uKxRbQdnvpyEix6pOo3e6GqvImMkzOM2RR8n9khetwf1VkLD/+62uqnEHcO7rVFQz7QlGf8ViMYU
RZhVOQ5hbzUVcVJju4JTW28XvbAMGbQjmEle44h87nKtOOVwTR31Cp8TNCg6IMQiqL387GFkpVYb
iOoZdRTq/Y1Y1a7M9R7mM7OyZDQZotpo/ByxF0PelnSCkN9rmqSDkMX/zlP+6fGa5C2yzVDiPQsi
xlC0AefuRHwlkDJI15DepT5LGNC1MvdoT3p+mXfD7FPmhZs+4twsNnXKmmFraakmKVLPcJtMuUBb
XgJLK1Gey8Fe74pOzqjcNH1aDy38ml+IbtsDU3nYyBSZrCBKe8F3XffnjxM6BRgU4CZx5o0dMWZc
VtgBIq/EL2gb0GShONrFeQpE1Vt7Gznalqfm5qUnNB5hqf003avzRLU38UE9yKJ8nC/ZrHYTuuzs
j4nJyYzELoGp3j4sxcFC7fSbwMAhl7dEmzOZaypzwtmYStRAxP7NXtDyBRt3CCgP7TxnOC4QxOxX
JjHP3ZgYcsAcGjaSXAnqPTu04p57RwbtmIlU9QJjUI9bYWiqRQmV5uHdjOd5V2qC1HpLs7zkTmsf
4QYn9zVpXzVlzXJiRaHJgVIsR2zkgGtzNS9U4+31cSGJxtpBeqAABSJjOs/Gbi43DYTln/UDpj+Y
/WEMLmhXyQhvSp6NGw14aunXfyxDGR4TGMp3wJhD0f5OwFT3RINt7nuuQDwGX+GPQNhZqIbICZfJ
ZeDsBin7DNmRLC+fUlOA8c6EjSZrTFZCS65mW/kKPmodbkXQhKBbZ1ceQ7vkQwTTw8+wsTDsDGYS
G5qlGLG33TzVWf0EOpYBn84lvuB8ZarNfME2S3DsMzaFlr4CwVFzbx7lICtkckfdlucQ5oxSkd6c
BogGSBgue1OGW19I5e0pfA7OqilG3slXA83Cb4OIt5IAv2N4g+zAyvYNj40E792M36WF6G62O5/f
J/nqJxgeOyt4eS30N3RWcDHaZTgJWAB8EIk0EKr9r3DuKn85vVAYuilA48y/QmfIhsXltferxh18
qxFWP9+DAiWUcCtnNVe7vTp50c9KfeLfOcw1b7L3XoatKTRMnoJruecWlGyCXg5MTkNt319SlO5E
/9Q2GQ8jhauh+OUMm91CtP4F9mLs/DuRAPeFOXbJz8T9ZkfJew0llOjY+y53YBFaAFWAVlQD87bU
JHbFui3HXC2UvG7Shp0tf8rMBoARpVEjvopkgRb3Ypqh/VARNknkjqQgPvm6hhzsxZJPdEePVj4/
j7G6Hv51Vb6QEJ53g3/n75vvuIIx3Y9UpaC31CX/0D6hfoq91gtopcXTHVcp7F9xiCETVeQKoPgz
blcqTTRyhE22HeVQn/tw63f6+2kmwMxSJbl506/QU+xHxwxZhEzd3937ctRsV3BOeOjBog4q+9Kc
BePCVyKfZvdOK19rg569hr6AWBtxgEJvKtSTM1ZYHkSyPYrPySnG/ptolwnBxpKid9hNfBVtJWNq
WFlTsHF6kT4P9jcLcgq63ACwKHRM6cGAtfOJ5e+Ou77yaoEoeyB+3p8MTAksvI44KB+nHyAYJlEj
zubKVzBYNpnqQ6yfUht1zoJE3fgl9+YOiUKmYG0wFdzh8LpXOkq6ffuZvjJWqgHPELXScEecFUBh
l/F+2YaKuJVbIaZHzH3UvkJ1ni6Cgf+Z3cVNufBLnw5+WeajIRhQEE8hUV0TzKYKPpdDikOBjjYO
KPwy3d8+3jHJljVD4G0qFw2vcSLiYE22mY2ja263rq4sj7tbe5liRFjpuchP9KYmkNcuvvyBxOR0
Sc3F+YTKEGCZ6x3dF1yAhUBE/jZJXg0h68r2R1c5OEgmOzLF1wvveyPZv0yo3v0w1xooH6Mr5GA5
Jw++YqGXQf44PXUvPGJueKg2EPF9Dp0y20w/icexwPb700muI2O7A0F4/CfidwgF3Cd9z5znTBmy
2fP5W/hNUyN+itu5VghMS5uph25aghASY+IXkKv3tMkgJ5NmBxPewTNWHmc5urcEocL8c6NLQTig
UhQxiVSrXS0yAmBxcXb/dW9kso4zYA8Q3HiHJ5wKlbBUGh+NjwXTPbecDLWV0JVmlGuHVlgssc5C
2CLssEK1W6sDZJsj0mwejh4UNhNpoecNXUv36fidtapHKyXW7QMNN+KdBX/BBHcX8m09EELyFIDb
OLqPdyt8IpdbnNVvdvmZzWXn8iytzzCUa/nfT838jCtZIeJGsrXKESKWIF3BA318ZTcch0poUcDU
y2K9RHxQ3rjEwsQyGl6NtNpZAoVCe8tWf7S9FD9D1rroRKv5O0Jf72It6HSBSpWAGEVPRS1QKcE/
Aj5PtVpDnZ4CJQcVSnqqPAjNuFApgjjEEN5GJzTl3SGVQe2lEM3YOH0Uh3ImYzf3CoNGyWkCQ3UR
R3qhArZZXTUQvAri6wwJ7fobKcw7UNxdczG8lqQ7nijAE/WDnTEA2y7gNMuwmspuEKbjuKtmsvJQ
ZdzUcmgkr5rwvCtxgN0oXuVvedbPXNpneuNvAHvhkNyAWQ/NH4wzmu3xN7pOTbwkozoS0I0Rb6sr
gLMrePenMzHMRw7WIk4TEYAfiMW1fnNTXkZav1m/Ds+wWfRMQL53Q0k7+ZfpLNbl1fa89qwpClwW
KgfT4E2GrBcMYfj1snU2h/+ez6iVVQRZHYc0an0cJivMgB5FB0uWJmRjKIahuLooBL+AEPMatJWZ
cr48n1fWByFgvIGLnnnxJuwbty2BCzs+BPiUV0mGDlmTG1psgE/D9tZy6JFA4FzaBmnQD7cnnD9f
QfDHj4WHuHMtwAV55Og/dJnn18Dmf3IqSsdlBMJ+7t01leVNKM8UZhfbdFnSPpxlspZLEoO8/f7b
1GweF/aHHY6+j/VTJjQ4NDNOzUeyTrSqoAtT8FsCqdvzp6npYt4ox+V2ulUNL0GnGmc1q01GHVLg
2iswB9GLeydgYoPHbfVfWcz2JCjbYbYTtWesZCuT1MJNkRsVjWLnPOFF7Px6/9kWojnhMsOKJsy7
IzSFgFipna4HOsJfFEBfRS5gJxTXAPY7brNW6qJ7Kxi9P6YK02Fa78PRN/W4r2sOPVOIGjbxuKDq
pNsPvnM0fxe4RL5osKu1+n/wGs6HiE4fbjygSg6W5vMw/M38vx7sFyERMQqLh5AqBmgypFswXBwL
jZm2xJrHvNc2xdv7L5KmaeO3ICoAF7Zz7xKdeCWYuUwnKhqkX+DEpV2okG/kk6TCSJ954b5KG8Tm
9QXVpQ07GtOPnzMYv+9uUZ6ap6tDZ+ndlFBE/Pt6NoL2Gk0jgEQj90Gtvw5f8b3/NdVwanvcvFOv
FQZUA1PBSTv090h/KJb/eVQiDgasbCeKlxVci0SbksrkBMRkqJI0EnpwRkVx4dAeWYW2JPoLM8Uw
53mJ4ik4oTIP9BZUQlFVht9tdYk2qFkXQmSBN4XR7H3looobVxCNXoWte4g1c0gruZfCB3eWowx4
vgcSlOu7KJu+ZODDCJtM9vCm9wdt2GNjumc9VeqWyuM3baOjkEBpvJ4n2u2KhM1mNacsN3Yk2zf4
3yw16eASUKA6EXpUGyVPqkDZe9KaGaNnq+LMnvw5lqGBV/mFm7/zt0Jk7de5NHLRM7/Ixmo4cLHB
26t1fK0uz/altJxenptIpkS0C8IMA2jooXI7uY7nvHWX1g9yW3ZJdYfVkzBUvAy1kaWjE7Tnr/xc
GYUTD0SVZjgkyn7CGkaNFDok0Y8wAA77qtDD0+8dzRci+Uor95+Aevtn6ADbFJ1j4WVwLZrS0ZX6
JcYkXGyDy2RIAwM+JdCMLDz9j3WTAocNEqOtYGaKnMXEg0Ixz9dtDmZVKFFdpmf6IXiykhQoqkYN
gjs5I6vYFXY3zNxH1QHdNnWKUSeBgP7DzA4zhYn6ALAFuGmZRz9ZHVXq7nVx3DaoMUJPCSPP6eMg
hsY8mKu6QqnteV4c5A/KM7BTwoioHMRxFnvn4s6bdJdN8bhLJ8qork96PDkIlx7fOsb2YTeW3IEb
B+6wAzlOkHI+OAzCvzkGgzzx6jAMNjsBi1in7H8te1HhDGy7HO3gdENTVZLdb0t40ZbNSyyXA17g
9GaEEQpEHj4yRsxufI3D73qOxwPFNgWD+Hbca4rJwAQszSQAO7dtO01OMVS9hXmEdz86osBBmWlr
vw416xNZ/MsxQAXovzQW0oHOVEkVlwxnVcW2MAM/RRRCoL+Aj1a/degSQNJILD3MOmusAdoIgVtP
LOMuZtQYv633RvPgT0Wj/76yhcI6YD17+3d7cWMkGgNeWuUsyC/qf5KXd4TPYu1FKr5mEdBQiIag
Z0kGOiJKHd/kFIHFEHDUO012tB8VU1682UbaC7lDZzyvk84qfQY25R6Rmv93K4IsfS7ZfYO/+kWu
tCmCeZS+Ij/cB6Y/JGRuEu5wgcTXwVx0PV+7wT9p6SRVnOWigUxEwjQP5OPi6mdiJRscmeKckYFd
u/wi9V2MfmfcCQQEeguJ3RCVtefk/+HCNaaHjZLT+TtyxVd40My2p3U5Gqirmkh2xzbnnPAIpXfj
v/gqvMY/rRG3TD0bbdjcjWlmCBa+F/ALjc/j1wrSBfgNbC6orLwu33z/vBldkMN22u2JlqTZqTU+
18VbP0kareHGubVolfo1GenUv19LZHIy9y9lo54rtIwNa1Q+q7ZCP7cUmtwPgWGbJBsSosH9dC6i
27NbfGTx2z0Kwd6pXiWtYBSxF9AEnFQxuR/3kiFa/COPh/IwM4b+GN4ndt0vKWN/TpRMGcosIe/j
MJ+8OdbDR/5k3e1zfUnCDoapMLTlAuYUKbdqFMJfymLzvDGi47dKAXn9y8q2IxUg7uon9lxEwyx4
LjWEgM7Cn3QMLw+N4ISDNTb5vH9voHbanslid4wGMxXn+tya25q8Wk51j+VM5mXsj2wGfrWVQb/M
UzLZyXjyHO07gw82sk9prqw++prh2eN+eFyblpAKuGqq8/zmlz68TlU3Lfa8Xy8yU9O6xSYorJ+1
zFT/rZJKsuiRgaXguSc9E2EpchtIGa7eTMpLMabzKXgMOLUUKzTF/ZGmbybfXtUBkZvim91A3IGy
/O6XOvc9oMmGPMQaVHjePGYWNy4cdTU5TZ3vWKtJzcdVnxer9PoQZkniCm+85tNcIUeCc4hqavd4
iRcLUvFXWNSPESCGp3f7RWYClyFAo2ulqVvCY2COO36juRHD/FyM5jHk6+N0oCUPkK8kF3MFKaqx
hBZLyK9vFee/E3rpIiuW+Td6oY7SKiUirUah8i2Z2aFli7Mjos2gnsT5MmJmNDsG/dzMCHquULDt
npjDtAAyXl99/VYkV9pksY+iH6bJEhaErrJVTixGzBcsCDhEU64YFrZxQOWZPWOO9DVF2zMymex1
8Qmfo6LYk2mz2s02F5gCeZdqwt/cdsuRK6WWgvXcp0qD4+WHBfhmC8lFgzRv6KV1h2mBuD7irbHr
YMKgGZEPX7E9fETg2xLT2sCUZmU0U37jxbZGfn0QdEMCPrBvMX+O3wz84UCUxrxjXzcPfahlgZwx
PSvjsBMfQJh0ej6g9LBCkEGS34nd4Gcbp15fOvDKcL1ttLc1shXobFVCU4rju30R70PUKcxEjlgA
IO5Mh24WbOaawxma/Siab7bfIMKuisMDHjKgxmb+n3U4dEm4eA8JBmdcGEAfASPswMdBBG4oZ0oX
MLROofRMkHFdu5BJ5MlwXRQFe0T69XtbWYyymaSyl4XjWPBAxqNtf6tp/YIWz5iHdcZUn/GvP/CB
s/ahrBCmnL6i/2Mpu83rGQbib+ZuxxXPUMu0B+Aay8CRGmfysGlhy42wuD6LcX7CYEw4L24bJWw+
SWaDaA4ERO8zQIASAt9wKfExCSDEWC2Kco8OgBFnMnADyNRJWRwpaYZwQhoVRVWV03Y7FDHDuIMj
0FLPcDpjzJEKV/bwBon0049m40uLDDSRfSMOnvhCeeVBgj1IOv6ePtzvbQrDTEmYQ431um56YKVa
sKJfEGbhexyeu/V6b0bYv5dvL9ccYyxNRLfcEzlibtgPYmnI65e86dueej0b5hcN8wrBogOpXYrr
IfGgL5UO7XprRNg94cyKHR1J5BfxcpyYi4l6V3PTwISNBbNkS3kHPw6yHTDlmZhz2dpEW4pzmjV+
UWwQ3tBwXtCW5y+gsiCw5iifEgK0BMon+//cNRME1Y6FNgTSL19VIF66IKhVnLJAJEFl+uXs+qih
pRQcsFJ0QP4bgYSXPe3QJ3N3B+6VxjMM7/NzSYKgtTsZvtisIoaoqz0VruKCEPqtrzic1yo5k60F
Xm431TUQReMXmOkzBhnIJk3smqFN31iQIGeJ6E4+7Uu1N5v1BFZl+K0hE3MUiD9etVXWXtlC181y
O/XGhpxBvFIQWbVPgKYYPECEJMVbrVDMe41URovCD7ZbfZbngYXrdhlP9Tmlg7gJNMZhVICCGZ4N
thyAQZp293b+HPwJkExjNspmLCHopd0I/4kF7QMY5cuczQSiXMZyuF8mulYHojrt1wsw3dUcakrt
UYbopvlovwqdBtRyTzi+0qVJ36L2FHzKDTngpQMG5yxkpTcRFQ0GipMq93GDpmmOdXXiq+XGNPUo
QZF1y9AkyZ5UFeceoe3IV4k/o/xYQIgnZC+xhoPdbqt1T0rWXCyRTQJszhipLRCN3guBN61Rg9V0
lZN6ULbebQuO+DxnpD+vozInQ/UASur0QWyo8boxvcZCAC0zjpY0VEyqnl+tLexvofvrNBVDpTHB
tYtfdFDQXULgS5dY4y6TTp+fKH5MlBCMSQJDzPV2BUA/YVwCNLfl1ulgzg/3ucx1n46X/kqwRipN
PlT5GfndJHVmqPC+pxe3ni+MlAXVQ9v51BpLrfval60GflrRinZaNLEjAIMzZk0zvgZt8tMKZjkm
JnMcWwJvw3d3kvTyD2LYec2vF/jsHZYJ0iQlMZToNE3XnKGrkLi2V7X893nnW8JEJMhpe36W1Fuy
AgFZmMyPyhpEeafIx9UXvHUwj8njW3PvZUyNvQU2soQXdC5qBCzvR5UDb8JTF2EuuWE5ffvaLsed
XHq9Q12azJX3u65nGLz9hp9W+4h10T1ssx+1ja6owiF7pb0Gec8krpDXwAybR/ExAy71oPjYLGcl
qOHmP4IS4Et6uTrxZ+WP7RM5nO/a9lDi7Doizy4Xi88iTrxmRj28mWQJn7YdpPZE3Kh0q3zYRXvZ
3ZazA3f6KFnM2tr6f17anRvPzsHOBx3Tbxar13LWOM3JhM8MXINEveScXK1f3/4WCSHQAKjqEggr
n7qS+uWiec/gvkIxP8Dsp2dTM7Vc7QIFiEW2DsqFCuHM07lUTBdkZJUOAf7ZNeFqwgyP6wahYsLo
YbKJi9eQ5/x/+tP9QyFS27mNhbmbqhPQzzchE0P2K5NMkNQGqurv6Buu0fjrN0vM8QpZSCFm+yEJ
ZwHtgxn7JTNFiXDGL9/vp80jhZpXtbzMPIR0fcBlazaKoUeq2FQK48osmgIKdoqJxNWQUN//tRQ5
c+Alu96JBHZ/FbL8eSZcKJE+DqrYjwZtiB1iFG3FOG2OE00zG7tAN39Zv0oTNS4Xbc/T1fw0bJsf
OVHZQRWtUvocT6mpXlHg6ME3VT5AyL76MQWXe405iBkblOg+23fSLsT0qSpUtNcNb5+FJSRxMKRA
hFgrPq/QhUl/KO7bf30DDJs26mHQoeyxB0DiZH8quNqaqilvTB8cm7uWE9PqJpNS1QLxCLGljmyx
3/eGHGuBW/FCS5YVoV/MTXH2ps/yc/8bC4kmQ6SSUX9gxvn1FCDxRIEm/6GBy3UL7mwQh5qGScHu
oI7CdegBTubJJQlxXJTzGYVJbscF34W78apNh7FvslNHnWdzlG/I2/5ticSBKu01dXjAhXjPWIIh
waqpYstIEtAqOFup76wqGlPcpAyyOJpcuHc8fGNXYUc+J6y8oVm5RUQOlLPG7pIfVUtUJrFVKWx2
WRXD+KX7q2chiMh7LqRqGiKyg0HKOduirFfDmqAwmUyLJo/ZcIhuUiUF5sUOKHa6wdv21H2Qtm+5
hz4svPw+JK+lB9HLmeeGbHFiHIXMKoUzTrVTcG0Y9ug11D872ltRmtHkYAea+XeqvF8mUGqSgTiT
qGH8GJPeYZUFN6Uoa/wEYAukWj3JIu5ZdcOI1j0hS9GrABkcSkHJm+/3SuuMKWFgZIYOKqyt4ZCR
f8M+MrY07StCqEVnc7tYG0TE3qZ9KuSKN3gHU6n8MMJa9e0fB49Js6SA6qHNR5dgxonJJ+aR/qI2
cHX7BHsoVBMhfWsLC4tDLsdqWojIeTFaD4NuwW0zVFbcx8rOnDYWLw+FZXW/4xWqf1gWEdKg/lSz
jXKGlPY04SwmDG+2ZxoF6jCqrifF3o6c65bdVH+yF/fhCtf5ywufqJrUm7E7+w8qkij5s3L9gMcy
eiqexqFN++ha1YdyggpBiI+hqIwiJG/CTYUVkqg3fOiO0YnrNih5zhVLYANy9C1WfFwir8eL+C+7
Rv5GB/s0A9eN23AlZSZ5MBsfMz3tjqlddBDPWiJZ8T7IVoFFzeIyYqfMyhRc2MzLciDRmPSogzvn
h0cETv5uP+Is5vpS74KHhpgkIIEcv/4FE1eG7Cz/Xk/PdUkpY4c2YecDsgtK1xhIhRdOWNaDGnQ8
meJYr1ggMipzf0cH0bPUvdLVYhhaZvZpyGyprft9GmMqPSY6THyudFDwyBmOYKuhN+iwHCeLjn9D
/CAdJXD6/L8uyj1zPjdz36zenljAdwwoxYKPgwIhhmLG8xVntaTmVmoYP7R0298+LoROlLTzGORI
DBCEBACGRp8/gwq2jprUuVxGoKKUREiUktaVIE06Sr9+iX1ALxqytVBb2jfEXpBBpG9/uS2qwU5B
EwlrUyE495hoEaYKYwXXaAKAxhLjXXS5jPfoNn03k3RyWbXr8bSUFDuVYwITL+BMjcJ9W6W/lcxV
rh50UPyCBxGU/CLGZnq0s8T0RC/fihTrk3z7OynOnEiIZGWhMQ9X4iq8Bpky05cpf/xQfUg1z0+d
fycX0R5qFf/0iONJmCescCD+C66QeyD6SV7khw7NozGPkiZadS+QUJW5xPV7PMdoYckqrandbjJk
7fpPmO2wnjDyK/RCXXZTQKycFOUvmACbnpLfYH7seSavV/7t7BlgYJ7LAZXz9BTwmYcESWLlQkDo
0CYCcRZ6v/XL6Oo8XYP6RVH+UZKCpM1k1OCxUc/BqmRHnppzKa5mS1qV4D6bBHhPZM3vQlG3jFwJ
ggzUb36lzzoJMSlFwyVE9JgQVfGiawo/2mp1PmhGyWBG0NFzk6uGRQtWVODMurq/75TRY/moDuJo
tNBTyVvMxtmWTWi6dEQBxt7f0B1NUeOrcL5Ojl/E/DAfmCRR7Md4xSBO6ZXPuGN6IwxNzqAp65M/
CJADrQDRuokSOmfTc4fjTd6Y2W9Wjeyniby9jZ/iEFKniCFA2rZvQ0mSm8rrR4R9BbAUjzLQpyo6
okSQR1K4z7hhWtxvOtt0mGKHmP8B3KjX/qxghLntKWOOU9LrJZnrX1TIcptqwFlofP862vY1eGmc
5MlcWgjVC/nBUSsRWffBROVaxQe7DKOQKH5pKGBmyXC2lv5Ss6h1XMQ8oOBB359HdrhyDbhyTsID
xtHmX5bkUfwLvbVnfMEz7fntrL8wRjZjeSjN/2MPQ7+/TaI79+lxB0GS7zpbf2gwPD4eAgJ7aG0E
dvFoXu50ZnyDNuDfT5O8ZiG6fxxWKAhfYgE9H/JupSoV09/sAnC3hkXUvE2KNB9Prf3dC/0lw3zK
XyoHLD0gXZ3LN37Uxj9UetaZinCaPSZOa9zTHoAWYqT2BTT0RnBbZxnduyob8SVCtvvccMphroNt
68WB7lCot6ivEOTSdJ2dG93lWyAJk/Qjx5vy/f0GGna6vOQv5O6vg2U9Ls2S2b5M86OnQohh3cfB
hkVEr5nFdJdb1AlGkFxaVJj4iNY3UpoWRDIQcN4qIxmab9fa52QaPpcnqn9r5y49ejmeTNywtIUU
xsi1zrcHvIoN2RJYqcx90PFUjF6ylVjPrKxCLb3x/hFoMSit1azT+KE3E9X417r15VSjASdFhBbS
pXSv/TNs8/bbW4VW0TJ7Tvrxlgee36zPgLy+pnSXiJKrNa59FWX6sdAKm0Zk8HED2gvQIqZIYQpQ
CrpTo8m8ANlvVScRVllnX0ii7cFSFomqsEJZuZBVSxJp3qxHX507XVmCSDyui9DrC0haO/MV4YCW
RCZBgL373I/fKtqm1/6gIYaElGBynnh0g7rAhnDaloVVJcOBv6GL1aSbs6ZNIALcnbmxBmbJKLOi
CoUzgPIjaj4VHy2sKBUPJeB2S7KhaFpe+mwnW15IMyDEQUahw2mFBU5FcWbeNk01Tv4MjjKqEXEF
TlMnI+0u1KwdPcfrDakEDaCYB8wIydWEk1AtjkXU08SzHRZ6zUxSGqfcyV/JHRgWo30LW9hVEjr2
+/Kz91xgNnPPscw39MXpoMdXkiYgHn0YoFglBkhKrzlS7dNgG0D08biJodCH9y8iUJs+FDAiyMzQ
DBoQjC3lHnr1sEUdAg9z1jm80MuiLn1F6bmcoVkA0f3vQL7vuou9urqVa+2rIT6v9sgF1fMfePzY
gQ9LbuxTYfvbO8bwXBSvMFjSJdm9IcI1NzfqZk5BbnR5iaSZk1Y15r6e+3BzjwtvJP0DKmbhHB9S
Do5qpTHnKyiMBWxxFGOZ9ohxBveR7Cqy92weugPsIWTt2088ObSApfaKPOriJBODX3U0+e7WRsPF
EgdX5eZlql+FWBwxIVvj47xrWFWn8MdK1IWwEh13BpbxwxIaU3o+tJOgiUmEWsQW4FAMIo/KIsgx
DJ1w0fnGM6GRi8fOGHxTmLhxDqBi1Bg6Pe46ANBceW9h9E8bz6maf/JtI/RR7esM6PI4DheKEKDr
DVMrwRX5NqwQw5cViQDXBwO78IdL4iGmvmwa1TaaW0Yns7hHlCQvxgnuFeP0jBgGXeMNHVqPUamE
6D/smX02QUSDQiXZj5UeSH9VoDdV47IbA4wxEs3uMI9R8WUci3zAwDofla4XrLAplPANsSN2l/+b
7/7bNaf6EUupj1yJuclsmCdOlt3GGIkcKZuYXVE2XUcUZ76RvdVeaaVWFGPSY6CoOXg06pqTAKGs
hmrcx0NusZ8VmwgTcTXvTLZ4AMZzJYMl4NaXflYSsQW4IzbUqa38ZuG4EbGlvm+QIx6u72CFJVbz
JrexDyNV31NYG6qx3Yw3zYk0Igo110CjwauMCeiw5Hycgwq/HN//U9DN/P/FEBxREK0cD2qkJVem
RybY7FOyWiGNKq+EsR4GXiB9ua8Hf2JERA7dE+XlFZdRoIMBpAjZtp4EwvccUL1+vqJlWRtBUXEE
4Nm1NPlHVBVM2oYoyKNgcToLp1jP4sTnAikua6hnl1wNmUqRw4MlxwVjx3Hwpv8JIVrKwwhqAFeL
AlP2Qvg8pDYDLI3XNh4MGXkZNsZU/+BV0qj+gjWGKZj4+/iiY1KVvGDOJ82Jhv5QbhS9H2bWCmWu
ZJvEf/Bun8qjkLZMBM7V8PhXfYnFX2xIxDu5xH2fGCsqwPB4Q1nR1aH3dVGvZptTWHnc8z3LgEm1
/CDPjq9KrRkRhmu+ieM/APGZdddfyQen8FhqtjWKj8N59X7iZVilyVT/r21zrAOLFQCAkifksnK/
DKoC7dFyMKzaT20XJDtaHb1Lt1gUyOkkyhY2OrdnI8EhEEvW1E4oA8FrP9f5MnjLiYzF3eSoMa8T
i52p4w5STKV9uwAipO7CNEZDOXezog0+E+RR/EjUNGPmWHWYbSFHirgCKy49iFBOvZ/OOTLpjI23
hd/fb2LC07UxacBg5NYratoa3WX/TkUkFR259izy8OBzXrmmDlH9JMj98HB6SSboozGcLH4XF54j
q07ELvZ1utcTZHGqgtvZblpIePrMxGl0tan8x+r1cSL+PVe+5Zc+rdRpNUrq5h4ZbH8EBkxpIY8T
1nTB2hhLfpFJ6ihz+X4i+NENFo+0ItJwJrDEwzTls/cyUzgGViIOkQPug8687bv8RiOrBTGihaE2
lJliq1cvo8qFhkiDSZUT0YFw0mbdPgNIxcVBYJJZsonTl7ObBkDvl7zdMNZqo5agcbRAY2eslFMV
yFKDck7gtDb9zWmVLI/vu+pnmTRCQxie7h8XRyC1R4DW7CQ6VrVLXIGMYTz2hA1RK+3uXG+7FyqZ
p/LZI7lu2xQ7ZOTGxTja1DdZCdoi9DzxiOoGQV/dE+t1muVRoeIXUCf5rPOVBNHsSNDE2HTxjGV3
oJest5YTlsEjnHqfyXWSsWGmeGMuQixjc1++u6mOIdA7eY+KffqlRC91YTBtOyW1MtCEzbQq3kYo
uffNjPaSgjaDl2pEMgwEui5x7HmIFua82WdNBCXP34LmXXKRUb8xLZXFH28p9YizeaoGf4el2rFO
Sd+44TavEtBwBuP0jjBUVRQ8bKM43YC1B1i9MPAM2NTA9pTEdLWxP2Fre3QkXsgvalVCyU2uO3zt
ahHMGsNpwI5l1ONXrgvuIFeuqen57syGCe3GXCFSz7/Q+tykL6pUOxobuMRaqc33X/2FVx6GDxB8
DPzgePHpAoqxRqyWnoCNe+KGHNM7T4+g/Vqi+Vt/p524TMuOxHix8HlKsdEgAac6qOsSQNT+SSTG
3GlURDLoa7GTQfiSOO6BGA4oFoFSlhZ45/m6iA5iNDhIEj49Ihll4FInYwguXHnkil+Z2x0KnBf6
5F5ratkBrvPxfRPsK0tigtI/Zum0xmhkgA5YACYq6beAYQnJgb9Ye2xw3IY+Rl51wmqGPP5X4mk7
Cb2T38EtLRfvnXvd3r3yynG3j+3jNK+nJbJQLxwggxzqCv47mpcesoMYwPFwGnAkdXil9Pmr+dGy
MvQeXNgy8kwuvI9aK2HOttzL8HmkKTwnGh1OGgr1MziRV/ZdwfahZDSRe7A75NJwLBP51JwKIeUw
9aDF+n3c/iiMaK3izkl7DVehixNypg3JcrTRhqf9/tGL9Operkblbsr2nvM6GmTHh/oaPdKmFFVo
5g8hCKhvyxr9tQVmEQHVLbD+QHgeCfKbHUqpZosVPJF/e1AvpjGP/PXU+toxKlZFasij8eSOOpwT
8TlS25ZK07zjQXvl4KS+WcfSSHa5ZI0CYvZ/P2XA0DXTevZdg7ICypb6gDe1xolAXxY8qGsOjDMy
UV/XX7KzFRpNFA/lmxYFiSwazO5B5z9zh4+Te/N3OroHI/tbG8TsVgpqg7FtXbHsYWj/pZJutmWq
iPi+2tQSnQjBA8Jnrh7DA7J/Sw3rNePl0FUiuGgkuHlAqG8uy3FPu7OMw9qQvNzvzeVBcCDvN4U1
ZwHEFnBLo4iot3qU2cIdVB0fmD0BYm2DVum4AseElDpB/uRA4VfJMixcgxtbhO/0kjLVLKrT7UVO
XYM5qpRxYJWjsbPfNblhZNql5Ken7rZ15R8KL8mNXzK7Nl6d/u2SHcqNjTMFJin/4oInyZYLS0C9
FUiNHqE939sMDEtK0nSYwzuAq5Psn1RUrfWU0+9sAZ2N7YPu52G+AWUOPK2fbG2kVNK1uf3ZIm3U
QVa0c9t4RuVY0MacY2+gkVt5nWPe23HumPdEnThbn+a1NtYzpxYVNLseMOiKKYwS3vdgGYA58jsr
kssHNa62A4ZDyPfNWnHeCK5yw058n+y2maThlHhpy4ivezaNNfWwnvvl+3jSTwzQECRLavwrq9uO
YWEy8+XKIP5e/7uXIwGJ3nyAbUM0v0CqMiF1Ct+jF0KoGQqXn277qeSxye9MI91fDJjzK0XyUAKp
cUWQce4qWqJE/dF0ziiLqE3l5Fd7EKTiqWSOd3cZqnrz2yNf/CFQfRaI4pkb5XqTRwsphZmZqhwI
LXs6SrRCIgKPbLbPsBAc8ZzNF15G+8eJ6zNVxeh+x9RJraTig3G5XFkgXmxwc+Gb7TqIgkbP+jUC
m2sUb4o661txx+vcWujWNLyFc7QZOSkyACr+lTYSsfg6TF4gq3ll8lKeT8D1RAAFKJ4kNBdG7mfC
i8qlUNwGpvwLeWfJ2md3QGoIowIg7NNryQyCUmVvFz2E2s3h8Akj3e/7h8OYqaaKouexYT2Ka0I3
tnFF8FRA8qJSPCsOFarlZFapUVUB0yCrgYN/VWhi1cRgf1xztY0BF9CL5Hyg93dzdn1Hw7zBKWeJ
IKDW7W+siyoGvvmeHtsmgadhn15pc3rNjH2QwWqxDObWs6F0AqQjDYIEAu7zMepG4lpJqQbqx4eE
bl+umEkbu47JcMD7b0DxvC0i7rCkyD/064khkp2me6YpKCJzw9plQIMHKSYsLy1tlvKO/sbjAwmc
SCMSHeYoPyrGOo1vm6Dt6GG9TYXUd08MVjHp4IFzX1uf9+WX9m+ofu091xDanuRQl4+LNkU+Yjm7
jH5qMRH5wY1JNn2TYDrUIXxksyDii2Y9XN599/hkcidhu4DJ8SydL98Cy4gA0+/c7QaN0EAInoIu
fXLGvYBXLseq8m/lXPIsrct+1rE3f8yPx8VfhhdLo+YxKPn0udWyrvl0439l8S9rRMWxjwMVvOVm
yDX4yx0lfyT1O7eNQQVx3ua4zIkCNlwa2mcNcyM1Q06OYIeBvNBUnBi5E0j2bRQdqW3OLZxiE/Gt
uFW34sWtALjRTuA5EO22jkybERA4bDxYZPVZ5MVGv0CNCZuY4FtivbTVkgGIEwGLPIPNtDnN1dHM
V0t6fCmEonh5wdCOXpn6Ldf7HZIHrIglk+OCssgiG/LKdwAgL4/W/c3bf5XDb01UMjJqRXthQkfx
6AZ3SJmU86IsLhLitbAFWcnpwDae254PWovhWE0Gdgi7Zjdq9n9tfl66C4n8ss6TbOvy5mqCq7sU
ipwzA6BMy3w6AQN+dClvWfwWDfDQw2NwYAi2SZAMb7asZ9tYAIPI/Eu01lR0fX9ZavaVsdj54Q4Y
ICNA8UNBmUzfS7L8IXe6/W7ywISbWeoczLNHdCItpKKk2xx+vESWoYG7/qpCY+n9vOj5nVn7MZAt
9RehJ7Sfgd92VZuKhH4P73IKzt1UlYua4E+fjRfKY3PmrK5Gl/CdXSvD1xrqFX6t7Oilc4zR1q41
Zp323+vMOjD5ekyKmEJJH9ZSQJvITZ4aHMHC313t0CE5bkFeKPL94QiKkgtEYqSs7OdZSjRAhxvJ
2WSISStO1a7YXcYX7d4pmwvY246RFsFCCal7m+Fha2AChBtKcCnL3ufmhv9Iq+IzDEW/XoDY6IKg
2OwFQ67IHFgTVDuE4Zt0R434X88jCJddKDPl5+WebQp10NxHgue5gnxctJNxaBYdzSJTF1D5wLJ2
Rpm4VpS7TQtXARFf0aPBO27tBSYg0ooP7a69lhNURcPiOGFBJpAimoQS3LyQGrnyh5blMEuBWjDq
IESiyc+bK6awJM8qNRQyqaP3tHlAGi87Hl+6O1ErtcACM6nH17b7B7u+ZyfHDzsUVqXrYWNdLaPp
58HMwiOejNC9JODzHwwy2i/BOn7KIlEuN2s5wC067VMzl2+e+PfdWHy6SOstqLjnUS0AQFWlve01
xLPB3eR+zwG9huKbp2xCIN2tw6bQ4UGEr0zJxU8tF5X0XKq1aFJPaH2Myn582wEZoYH2zd29ZF0h
HUWYSCNSsDsZkN99lRYcxE1m9JyNX/EGyV9TUulLlZOMt7uC7ImU0JjP8Ay1K+Pp7HH4ODuut9eL
wlzsKgNJOpG6HYZlIp0lNRm37RpppW+DyjzAqPkPJOXH7U9i0lUAA4NgzCN0ACnXVHaCOHjJRXmc
7KJsCOQWEfk/LAw4N6Gdti0smTPK3NuHhvffpWrx771TbKfdQ3RhnRg25jSH5Cjgw368IwMs4UmR
stl18mdslELCtXSuE9Kt9WMKwq85ED/WOgLdsGON3yO35Utk92HP3ZUonfK88u4mipThHqd6Dz0x
Autv+U/LrgCFPTyS1JXk6OpdXC0x+HUGylbknXLaSR3J1HP44fMJqvHblPR1vaplD6T2EhU3zUEW
XFg/GBVF3NR+hm4CbFYTKgUNNEh4CQ7iyjFQtxZ2sv2ezSbfwSCbgMItqY/fZakFRMwOj9Cl9cl5
HoMLJGjx/Wr6UiiPkup7JlPxYRPHzBIDRmXNk6tcrZOEPncE3FlxM5AEFKyqQQ19Zp+fXfMjTNZ1
N6otwBkNW0Q2VKaaQ3CO5xPh3cvHnQ5FlBuX9z5PfhoPvhupq84jQrnGLG0+Xki9/AuU47Ext1ho
bV9kac8E0bm+WFtjGP5cWUZZEZ+p6biMsPSzTzp0mIoIByjvo2149JJYMC63zPhK+pooh6m/b/jj
uuVJSdNGD7Maiv2PZp/2ULZ5cQoXjo5hl2ir2XYnkak8W/Ii2MJJY1fSUPw1Lvz9TJHzTmsC2qqr
kkHAlF/Hf5soXWRCkvyDFZVZvvD1E36whCXXf1JTHg0W5e74wbNStHg3Q47Bn03mcgDwrp/8WFCx
8ttz9/M9GBibzFOzMYrWdstptt5ZRObb9Hw7qkWkuy6/uDtf5gQbXuD8C9Iui2I5eGcVI2JgRCHm
zyiyCSXRS+kQLKfN1kzHfVBZRTd54DXHrJzEtyftJQfptkEKws2uMhmJ9S8EWyUtufMoxJLLcDIR
EdUGgDJRgKnT4X4oPt2teZ9xxZ3H+7nTNtCGtO/uwmEfNjSOifQjYwaEZ4CQxx5E0E8tx+M001HY
kSIAMbXVINH9qCACoy9DTYHlTnOFn2n/fkFOLioUiEXYZykEsjx2vcOtVGw0ZZ6hSU3BK9KkQkFs
CoZ8VjtDqzdAGMEhcNZQgDvk+I1kpEDg0OAzVtYz8lBGqi6EAsvAyurTta2cJRKM2P12o8fVw4la
VSF+IDqWYHytyBf4CRMRI+zkU6TQH76VNyI9VooCirJzyIKUOg/9fdoQWJ/cXQ7hfNBiwvbkyjhA
Vb1AZJ1Ijq471L4aZNgip8mw7+F6cVgIHx0CLhACGWz0MrvvDMhcn0GFuzO+4JBBwEdsgKuwmbNo
pICVhpxp5Ii1Xmlfq7zjXURMEG9NRIthNna+ow7vGx0DrTbTj+8JP2y+B1yMeW6QQWzexJvlxVSr
bgD39Wwo/Fb6C9xuYs++PrDopGTdClPxXUiO98trwylLh3Koksv1e3sI8dWH6QgLrTim3prO9iGx
B4f9/iRiqDH3Uord7l4Ei1c0oyVGeBj8OOe5iwSRrzack60BJuKV9eBViwpzRBU5ypQYCxREb2lH
rt/FhXmWMIIbsRmVbtlUFrzwvlaLlaZXoVx9uWXJzL3Iy5RB5Dumjd3+h7qbnZ37uKln66YZCEW4
kMJ09ueOx7CRWgcKwsBbtfycK4tTcHSUshz7eKOpiEUcWXB7rWnKBcsQHxijDBcZ3BG2jfztfEGO
TAsDe38BKlv0Y31XG4ce02byGoC59oGnODg5Vu6nBzyDz5aK+pqHmMJKIMXLQhqLxYjXHnWEiXZU
ySNtI3m8OWaQGzH+T+5uT9hpFOG+022Rsuf6RQbzuoCMe7Tck+kB2PE/mHz9qAaRj92GnZvHUqvv
FOMiRnmgquVJCOqsMYj3XF2Sd7YI+Z620gZVBXVq9dpJTYA4gIMsGow2f7BumdAK0bs+rctKmD4n
R4EmXhHss6Vgd3U4so8gvl1oGNiR3arOFAtuxvyGMjHkKdheZbdxdB4uZjEk/tlbk057tYCQqNZX
DrkYEhumUrseDe2LTjeJkXPGmi1C1fWoqgp86egMz9WnWmnCUcD31MyWaG/Lw+Gjnb2YPAwSNbgi
M22yBQa2OtEJtrjPFNzgNwWMt90ueWTX6O40nOnATZBj/etXZIzXAWQ9wCCKEKPrh+EuFPJQCX8E
0f+TMtYg3vJwDPgesEywIQ/T5e7LzOTd9yFUphk++0AGfUo1vrAgXJWOcK7aVXBRNAjLwpysm1pS
3PdqpIFQrQyoHZ+PfVxZqptqES/dajqXaf1nwMdgBFv8BE6/gt0+kbJifXg5cN2P1qvb5Z0Ddecs
2kPbjif+3LNyS6UyrBSfHCczOt2ejE9hnzQbK8sfWsDZP65KI7jiWLi3l6m4LRzNcLoswsvQtOTa
9xsvJaoq+tXEv9xBX2NXFWnJPk/f5Mjw//LvOevUfN9Bq5qrmG14+2Ge5em+BfZkXlBwcrTbZiW9
vRmV8YkeqBS2v5WTKQXyGUQtaJtsRlPJYEnpN7nI72WW22TYO+8lmjOkjft/EkxiE2aiJtDPBTgK
/smBU9EO5/vWdyNbyhnG2d7YPMJCVPtwnArtsXNpF0ZyyuhHbcBldKpZF2lrMOBi4qV5a3pxR026
QB+lvcZ7e8yzXp4ncQXlVncoskbUuuVvQvlLgfQkvnz8XnixXUlx4eVACmBjBVZ/N9MkQporZIBz
abjJpfvZFeV+3OIyfEnY+3uUXX9jGLyeYAMjyoo+ElvjU4PAE6VG7rNhoeHeo6Mq7LnISDHQgcby
3vWkJNifca4xxtxaISJl+nfNPnF14qX2uNcnkMNCt7oy+LHon4E4WR3wJ+0Vpjz3DBA5cpIu6yEU
DXiv86NTDh70jhRZmvczUtQ1cpxt+xC+v9mhdsAhWGzt4mKcYmSGD1a783tsEu/0ceqjLcPfZhzk
xPyDKlnNye8KX6AZ4EnIxz4/BH2LS/WcdNngOhYlQomCXhUpZJOAZl3jrafYpqGKPqVYdwU1IG+W
P3n5AfA499LSQzD80EoGI/jObz88cDF8rZfI1r85eo7v+41UNGcorGoaCsTnESalzeJb8OLFHg2S
cb+nhX4M9o5XXApTeIFvRA4VN4JBx+rywP2vsF2TUdbLA9y+Ie8AxcTAGPDeURywxY+GO5XFZsVS
OgLQsFqXPCTy7Lwtrp2RySESD811weSjXe8hDofPfpfEa9PbWRPtxjrbiOM1o0oSSY42b2M7xwNC
PWKAPoQycvbN4TioDtXPtbsl1yIyLPcNumqmLUVT6DYuTvo7Y/DZ7V/fPQ4v6/btqRz9GyLNBRhg
iBk/VQUozMMAKiPKkmdde4kXH6kSc3ciGpgFDUKYwzpEXE9nJOazhF4zXG5nkMFw0Q+8X0/fvFJu
pryW6Y6nTrYET8wXTU2ILjrImPCP5NWYifkz37tyPz+V5n4x62Z63xajfWbjAU+XyBJPsZOiISC1
ChHNIqAD3Bw8oICSinAfOs/49a2LGLhDLvwu9pEPOPITjUFdc+yCxNO2nIks6CTnNEYNZYZfGDJ/
3fU14g2FEESy5y6w4EE2c41Y0f7vrzhgAgtQMAPtEWe6MdEPfsBxm4bYED9sz1XJIaVci5NFz2QO
bDzoq7qg7fxOzIw1fbMoreBWnquZeLB/DxT+ecXKDvkOAn2iMb5UnqXQP0bTfOQvb+M54T7u1t3D
iH/NsrosGmMIKSS1hKOcKggHYigFzEIzP0gpan1fYwmJpxKv8kGrp6nqbDs4u2k147P5TVIlKDP3
M/vm5TZZ+qiI5VlfTMsTun367YuSqVwMbpkLH3GVgL5Fg8D3NQuxTDHlzJ+bCY3RbzaZmxibGUbR
eBjiorEcLbPOE/bIBoGZ1qwLypZv8Ur6Vmap31mHLT00BgT4jaQkdF/QbFXVLCS+63dShc9rstbq
ZRM9ehB/HVPt8JwlUBCAHkLZh5iDxwHnpBc20rW6sy121eM/fyxgnrTfHXDmCLsikwzi0koMh/x8
jHI8VtMgktRu7ziGOuEurVkF9FeOZXdrz/Jh3CaEwoQuRFkYZDYGG9eawAfagkMIpcw9XwiCBkCn
4eXXZ1Tlk8qINtWlYal1vSVH2fd/oYHQfIyLLN5QxB73Nqg0Y7fteP9olMKQxjuEdL+iwCWoqdvY
9ZyHhCM9t3gTSdDKjc/szc0j8ioSCT9xplE5uq/rSjPjWYjkNYCz12Gm9HszfgMfSsNeUnCeY6NM
T0Ox7ztuVoLQhn6WTWJXYXUmc8zYnRQkOE08MGBAMaYiS9o993CJRnpjjz5+LxuKtGh3L78DGegB
48iQ1j3E7grLYgm/7pBffLDiLMW4WaF23aeyIMhWXLFEthIxBZW1qT3TvvXhlAznCcwt/l1ZjNCa
wgGf0PvIJ7IlKxIYSlmBpM5r9Hbt8+lOjfUcfz3TLffta9QPsGyEBZgWT0Ku+PyXoRTOzROnKsoQ
qPrZNr8BW0X1KKqvWH5oZ8PH0Z99HXGMVZNustfIPbqzvxLRwTFAO8Y3ZRG2gnh/pQvuSI8Z9224
qRTJjO6nEHFqLI3OL3btlzR0QEfQHPjeMTliXqt+hn+dlgOTI+PTnx2waFIHjMezIQ+Rm3S8U0mz
6KDwNsjm/q8Gzv7nBC5eaJIDLFWIpFb5GvONO7PAKFLYg1r+S+jDVVpKv2r0Z8wEsY/6906ouD2F
Kge8E/CBqsCXszP8U74ADAwjYdN9zWsRqKl1Qbr9M6wYtJVuUIRy1RmkPXNWUyVSxDDZYJOZdmd0
cfZYYlVI1GKkrb5LWt2sT2zvRi0Xzf6s6FK31sA9WoJOS7avlCId7BfwVrfcWNPV0fuxFpb0AwG/
IMWVT6KRREQJ4Asnl8FuEovQ3nvcjpJzABzgioXCaV7w6o1EmngQjpw7TKwg/jB7QuqLhGtbzFX5
MOjGIIaNs58B/qU5nlrat/ZwtXZFJrvQaccNzoV5teVB1gKD+McPK0xYZafAOky3G9p+Ob3M3OM/
DUFTN3LVqLQVms8qzs+stVx9kgl9+CGWRFubzuLOaqJnmQxN4vP9Gtdv+zIvURS+ryRb8mjlKu+D
6dK0lx7ovWQmC/5bYRGVeodbm7Z6YXoDP92Ij5dStFYbapBbhKCuT+3MNvfIN6fGjyVttRjrdpFz
MQ6+hGKAMPEAhLFkFAQGql10fBxbsr9++QAhhQxfHCJmfvPqdqNhcSSuGQ1ZlNaf4zAj1ci2TS8K
cZkO7Ybl4WI4u9dNZK8BTKqXAjBUrALsQbzCVPGf6Ayg9JzH6SagpW+Ubo+Pw/gi4Chl/0atLVYa
aTrUDlJx9uw5QqWzIVljja3k5NeLnZBQgNVs2ArXmh2wDA6xqjBfC7dcVub4zXbOMLTwikEUEh4z
MVgSkxtlxaDqQTJ4H3HaghphGWLTClPmgADLjY20cv1fLvAdncb/LBr1akXVkDyDWdRh5jQRs3ZQ
lmoriO/LbDMNrqks5wfU8ZqX6UK4RQZRNLkad88t9zPJiC2bSLG0cEBQloNTamh0xdAL6imx9yuN
OpeadOOnM40AfJspEUMCUEEvefGCBIjyb+2s9WfdS00OEV4bbxZBR5aBnS/2C8MocX/bTpnMo+ih
xRyRpK7PKmKXjNzTVC7IllwSEFrjRwplGuiARVi4EidACTg/lI7ZYFfRiGrra3po7s5JdjYJpnKh
JHJDwdJoYAWip2KuH/vOT0Ss5Z4l9oENswDa0futiHy0KUxuLO2IOXg9+yPvANSLObOtdymCh32m
lp1a6o1VdTNbtyjwWNFDBbo6YPszq6KrcvKPOka317lwh7O/EN0nPRGKOJpu3a2wJ/bhx8O6AVkz
SsRjgfXrJR+5jRZDuhkd+noUCoRgtN81IJ627EYNc4NPgNuN4sOJUahwziZPIctF+dvnTaaxuen0
6gqk0YPeDEA/i+8Dab9PA6aL1vG+mQTNE9dwWT1eHNbjPuLyCOsPyBvyKG9jGThcgBvzuzgw0pC/
cUqM5Pj7l4FY89v5mDqQyplhIrVMFsCy32+OiSzob1xqKp/2I0hmTPwm/hqwRwZh+qt1yasu68qx
gxFNGMBfCGHcmFBDcMgXayCClbQpLmTSq3vQ+AM6K9OHFLyXVV+RTaZjc50y0d5srkQvgrexN2cl
ML+FwG539X8fndwVw1zMExrRBm88A6rTD82bBRZGKXGeLjlzb8DYRck6ZUAkcpE6RbLqeOSzUs78
yNFJDbulRk53WLIDeEYl3UNk6P9B0VDjxz6mzhHlD4HA8uQdWsvNdaPdOvvhb6g+e5r7wF9A3dcr
YNY9/VVKEUvkK05lVtXqUufeZlRkmkOCw4C+Kgi5Ly8XML27oZgaNla3OQZ8kp0+zg4/Rb/bhw2I
K6qY9YZqSCk5l/lt/G3GspkmcR0YNIZQOw3FBIJxa9YRdEbZVVtP1sZAOIgYggiRNeiyejRn8qZW
iL0gdKVbPbFapnimssX69dIBwwG4OXZaydUiWVjA+wJol6Ey+rE107ZbWaqzcl+NwPtidqeNsA05
ySplaESudWv3YTXyQLLND84II+qF8PNEeZsPcgSoEtrcrx+dbfeVVgKUhWcw1u2zhKsnoeGx/Lge
Ge7UWkp9uLHfOkDhAtGGSYGgYRZTmxOFcBqBPpLB+O02UGwH3eN4iWrdEZk1aReUdC09s5kwhaRe
9zoCIC/wl4+UR6bnX6B/RsyEha3iQWHJd2lOlL3ZHB56dQZX3SzwhC+rKNquPUdyFV4HBUXJayr1
pOqXaIaMR8u+ZLJTOWd6X5Siys+kV5gu5+YdZxm3VSKG273+ro7ZUJkgS93It8aDAU+CHQpVs0zj
v3QKhTzUq9u6Ga/sdocBHhqkxbamZfN00DdeMrtTvIV4Fbz1EpavX4CFDHkz4cY0LLf7N/t1K8u8
J8t9Rb+tIGOkxQof4QeFSk6QOkPMGRnaorhAyvcn+ezphoQvC0nusQZASn2aUCAvdXZRV3gzGv8V
ch3kCWynRdHaguFZk59aJNaRjyk5QAYv4pyncyK/QEAhYEbDH4031HUVYiqC3ou9O6NUqXd4kBuW
gIUSYkJyyB2YmPqP4N4nMzqn84dhqN6iT6bEBYCWwHfTtqBautp9gvSZChU0xKsrjPXZ/HU/egNN
ndfyuOyUjctex3bDDrt/yBGJT04zJ0HXgdNYvnV2qA4VwFGk6icoihTwcU6/TQvkOHcRgjODIIvr
pvnMvdEMlZGT7m9fWuQtsW5kozUk7JfkWFCh6jTFXnGOiJAQ4kVoLz5WChQipECVFQShdv8QEAju
vLM4X9IXnEYvuBojNfZKw3AVRr+3J2CeLlJf52sXhVoJnfHcQO4lh50xUT5aDmlTyNRTsWpVCmiC
2T8p4L8kIVaUz1ZuvoyV2vmq1F0tT9Ee/lO4uBU20Mqx0qupZUCNDnXYUgV3Vr2bJWG814i4vqMP
PucuVtdTwjNhkgmOF5sfDVcMZBjVk21WOfjhUXkzsg+Ve5Gj4bC6oPHP90g4RJNihLiEioXUlzmU
FjNbb8Rh3gSIjej9Pdl8RfzreXly5l50+o3AGfwE1rEmU/hebT0acRW4nbo0RcCMWaAxNZfNRo8k
del9BjLgdTTVGVLt9gtByUDmhR6tG9JADGCOUp7i76Hacui34KaiAVK02sMr6gITqffK9kVoDKqK
/d4sFAxqH/FuFY0qachAY4La8+Wu8Y/bh+4lYZJ+Ffc/sH4mExUAehSC0+CwomTNvv2/q2X6rx8I
v8m1OBop/ql6taFHa30xJids7++nGieee4XZuijYNx0ayUVr3tqL8tXVU2SF5nQCMDWox4Ms6Jo6
BalE+UehLNZs/PG+UKI0eUtN+DyOb2JtdmAXCaJIAyBsk7o9PKz3UHjfL2tcfmFl92rcAvyUf3em
uHsC3oLAg2N6nQuHG8pMhXCDDzq2bs9+DjD/3AHV0ffcIvb6+1rtFAwUeaKBP9P5ql0tejUTzyFC
0lYud7idXwHi30uEEh2CquKSqiQ9mtJcBvcgNzjUs0grV+AbmNDYfHFYBjrjFmflz1K4Av4Ya+EJ
eUSTiZOaWAVLOd2b/qPRtrBCN+Pi/JGD0/Wsy7J7L07zR3fBUXyhuticD6C9pimJMgTA72fmd2kV
DzOjVfBSHlQNIab1f5DYNUBkEc8FbFoHLxpNzNA7lRM60ZjAEnuzPjp40V1bp8jF19dLqEpxiT8T
TI7JEPUh2uFHO1AYXdjemnTRorRRN1ZW7evKVrFTC3H1hqe3rv+3kfr9/mjqDRq8xRksbNCpd/JW
UZyj7IJ9JGs8ACXs2OfEf9Ai6IQvJHkbIQzNxqIC6O/AZAfV6BtUSuipopK3HswDexUhp/wHiNwU
xGlpRnTBjze3CHe+YNsWGnI9vIrSq2eOnYlYoQOOz92hpalV9hcNa94P5ghNJHUNeiTnxIIUKsua
iGJ25JBesFX2Mhzrb/lwrBnYsYTkNEX3M7pbq0rw3C1IqL0Vb/7SywSu7iyPrpwIkaUpIcuaTSje
yl1cQ9Kz6zPYfLdoYbqx7Hbyw+Z1EaRSfxHznXri/qK+kV5Qk2ZXR2aJx0lH3H8HXgJ2wR7MbxLx
9V2VX5WRE8MJilF7LTUBJ/9/c7NDddjw9wS+ES6IdiaT2IPlffytONO6HuUxikjL9QeIVbW7xggC
yPJ47op0OtdveTVMPJBUzL3qc4SwZtd1+YWaiE7j0Qodq32zs2JQxh5giJXfN54WJTEiHkDpVCPE
Tdf3Dobe13WzW1fxs3qPxGUgt4VEnX8GoyHHQhqqfrpuAJl0IswjOJf+K8nyl3GZTsu2r2onHj1M
AGeezXDWL3glUvzZnySfagQdB6wDJC3UCsp5+kxzGDNUE098z/GBxltgWWbiPcPJTQQQ8LKds/Gg
NUx8XWlxIqlrJo5Zjwj/aJ7HsdBlfJ9FkWtAO4DkCSQ9vhnGnX7rVZsRB4XqZXsVVm9jRHb3vUZI
HHwujTslV6OBV94yyOwT7A9ydYEO51970mIg3e4WdXNz94dgg272/8PZ7mgV/GZymztZ5nStPBRR
9sPtVVN4tx0tGQCcHOmgbiAG8QDls1XnO1uMU/u05P/yWzpiAauyBRdACj0UCEc1ugO4g3q9+8+w
lc4vZ2WmlPd7ATTsg3AjwYNtWKOZw4L2ZDMp0AyPu3cK0jgD55pz1HwxZu0J8YvoKxmZawY9Qn5p
Y8i1v0ssUi85s9jc5ucXWY79mmXD3+vttZw+YVbuJac8FO/plcVSzhNTHq48s/vNx+RLMPwWu4fi
AuUbiWZmS9dAZhX4vIF6hDyCXhh/KksNsqCySBBFQoisSLsP/OWmUsl5b+JW4YcR0tAaXJKthCU8
rRZTUb0kwKptHcmKUm/TzpjV0tvYCCyUX5LGxcrBm6WaD1FwRKYqWACC5+Wz5+G4wQZx7qnZieR5
vtgYXE4okmLTHDtHHwWjsdMCdfCb5gYu2cUN/HwLwgwvaExhNUW7+pWjvF1ODM2J21cPvaxpHE9a
caKQDiwPN8gq/Xr0Hgag6j7AmT5MDOdgWZpv3xYY021BSObJXw6r6mYvmAFxVP76GZy3UXQ5TqGi
0EQC8Kpo1Gv/jcI0Zgu2YZw95e+LqUczTjh6HM14rFCtHs2/nkGn//C7AdpvhFa9PfCJ0v5ZuQrF
+jaeoBVE/GGJsQlPFIHU+T2dX/7bNr1UbDag6/Hi9dbSOOJXkEVewMzys+smdiJXJThrjLN+dwv0
kmexRWcqJaUoEFl3AK9fI8Yu6mPNZkYg9ioqR0xFPbgh1BFs3JQe3WAmQRTVuDn/nhMIX/747W6O
s3xPxygeCQwTlFqBMUZjoJhNFzCTvs9HIoInvXlfuG/5KIxDVH6nDs5bLUVzFwkFho6zQMTMee5f
iVbIaUpZ8igmf0cpXJv/VS9RDY3CUXFphtoe2Gp6P/gGQ7ib1bQe/NoDOOW99Vtrr67QGj8UbxR/
tepeAxRs3+cJcT/dTroxWpi9CEAqfkGUt/jTttoAgqv0OdXcdxp43HF6CNMOVUWuBa0/BOc8tLnk
T/kRDVNFLOD2ndlj6u5pirwx86IVs+jh9jBYeOTU2UoWJtNscePTEVRUoesC+V0m4whPj+r+47F+
tBquwu2m1da1PB+Vp22GFFGNnvSIB3uWttiWnpDQLZzk/ecxJENktI0bx9dmbKxMDtG9khhg1ZO/
e9QPgXJzNX3TaTSTyRbiU5JfYBZWsy5DmxrJ6K0ABOjbPbvQXCmuUE4LmdwxvD+OR9CxX9GDn3uR
zz38CoFk45SGQdV2e/W1qTiG5T9UIGTB84JFJLT8BeyyDeMCuN4EBApjwbOmpq3kT3d0ZEjOq6fP
a521ykRqP1XvAYW4S8Ul+vdKPHwjWLAstoVXjkAUscKGvyJgxz0AT/ZpRpieLyROA8KdaU85krFG
QrN7H9Bmr3OJyHRVUeV+4b1me8JVO/w28I1FRikg3QIiEcWdzmRzTA/X5Ik9tXL1gfLbfgB2dXPu
8bQC23rDUerz7KI62MTZe9tTGOId92dRvYlaEm85Tvv0auTKL1uBFqO0RPDSi/baK/B2kzgbtlhC
tgAqi6GiQLAXgX646so5aHG22O/j7X+4e0J7xr3oYpHEPILEKXXJSKQ9+T8F9vHRGxe+MyRwOAr5
/JcA6yftoX3XXAUmginOjtQpzSvXFEssDhHGj6CK6VepJeATKvP8t+PSv+KYRdLdTID5Xsw/CJ/h
9nV2bLQQWROyCrB8HPy4JlFugTnIAolg/EvLRTDvwjNYcPjGclsUQs0F9moDDKQ6TVsoeKARusRt
9vvoXZ6cHlj/CzFPKLIooIrtKp8VoSGcD4N2Drw7K9uee+xgaNrqsoY6Zve94diGIlI2WpZ9a2S0
Lrp0Hru/LfFT8c2iRQxAADKfWpmuCSdidTFGfaUX+jhaRcxXtoTVGGoZC/MWARV5M+FcqpIDPCVJ
D/AyyOkE2+g23d8yZeSIAeDWJ6yr8HCORmIMwMl2O3c+ib2n1Pnb9uQd+gRNmEKk2Ngf6Uh9yrJj
YEbZzOmlk7dLcnc8ujDWHfpjLjOI62ylhkdkm+G8toFMXY5LYFfkX6uuA6x3y9Ud0zus4EvTR0m4
Nd297EQqbE+yWx0zmCQaxXHylwLosWAEadaA6+etHpwE9t39eMBNF55TN5X97lmw55vXHQj/Sf1l
QcLf7gAMDAotkmMVA43rnU7QsQmvo6X2RGUUVZdxOKnBaiKXTSWbQjTAjrGHHG26asVK4lxI2fsZ
KIxGkifFToLiYu1sR7+dSg0BhX+i1Twjqcl6/bhdTGgFqZrb7xCUlZaemVDEchFDxjndvFFzeTE/
gk8tfI4gSt9O/OUN442FoWBd30E9kH0zkyiqEDWF6TYzSdDGA3bu7ViBSSW47bAS5i89x4sfa6m8
e1wHy+blUFX8D/CrCsD3lxNuh2xni5T1lTzQqHss+ed9IzVXiiQaA3O80Bg5ZxqjIDzte8Ji+e4Q
/B5wySC8pnOkuevbhpe3tpDSbVO6KX7Gvp9nOrpLG93uhGNdHU29rqkqPDTa685xpd7CkpGp9Mvb
L779wjZOSYfGDc63epntJY7GZkSm+CW0830neZrOBfhMnNuZDu4VMduhLdeZYSXIaQZ3w/tHwR93
foynQgD76eq1/C4gGVBMnxEAkDXbjTg9iUf3WxnrANY5mo6f9u5VRTLekYW3SdnjMOYPvh9QGnO1
26jr9ERhNtt7dEFw2bi0tPkuvjjgMk7qIHNTyJnYIqofR1upSqMY55444S4Cjk1Dba9hyvKmuqAG
d8HshHUXU99Q4bIf4dKvWsb28Z8pxxlt8ijJEGOYsrIouRZa/sQCORx3iTJqrkWhvmuElPBznnWm
Hz2gW+US9hpAbhDT8QypIowweQZZuMe3AXfznKRxbn3ZBKlwiBO5kZeeKmSzCIZ93ciuerSdw7Tp
kWdkClTAwzTH7heZescZdt1FBSFOls4yyphdZUnEIo4BE1WW0qWdmT9eDGD89PJAmwtDkN7euNdH
99onFjWokO42MYo+5x/rM3tB+E6MtvxzOCEdyi6vTca3RD2k8F3/g39MaQLP7CRTH5uG2N5pkLig
HoTIJFNPViO0L4ZTt1d8UOE/lEqzjSsgjdqrf5WPM2t1tTySIvV6FpsJxHsPtBJhzTzvgw7G86pY
JxqDlnOSAlB4hk9yPfysdfuyRErgHlscynC80s9ldHyJeFjtqo97e4Xj2eByh0BA5GiFpeaKERV9
breOQvuRcJjftQCi6jBL35z9L9PGhlsqO6w69Kpw48QAJYK7bPwzJ41jC/M4GL7+s9hTeyHxguvU
KZ5/P47A/A7d747imNcHx6bQohZ69fyVKck0fyHE7yIULAjnP4dS36VA4G1WvuXIKnTH3S0+rVa5
zYR9LWzuYSkQ9efKpTwXDcayJlprrjQ7d+JWbR0F8klaviDp54Vhm9WpHHgww1R1KCwyRPXlicqt
B5OuSNekDkiEgDJY4h1+Lf590EnBZ8FF+JDSAB7GuBFEXSQ69+6hN8DEa20FO70iU5aec9SPv5hL
Mf5mo2/Aa8E04ZDA8F8Ck7tGsr5GDLlqwEqb7w/VXCI6GcheZYuHRex/qbM7xlDLscpbyMoeAyFP
1MpAZ8g5qMr5n83OmCu3Z0bIoxF1zgZ8vLmmfMLJQ+7KaBH85/anAYrg/PtLBvO9g+8LeakwShXr
LyHVZlUlNsVU8/9Vy5hs3WjcqoXMbqavhd0Z94dYRHPwI9I8SnEE5Ysfz8bkI7INChQkxWgKrQwQ
pkFj17P9qU2vaGhB0axKvtai7Dv+q02sLORf95ZQ3qjTcct0epYkiNchbOl+8xWiUTf6s7KPfELS
j1uJigiFpDKVQp2pU12ynOHH3rCKZ2x3zqkhXq2mrTu59NbAm+pVeeIMNbAhBJ62MsMjHcMYYZmj
X51q7LKhku/mK+qmGuaYwx+gNe6HWXsqYBBedtefeTpQRllc5vzEst87Br3eFR5WbtLF0UfYHD9q
rrk9resjF4fgjXbF8iGThqW8HHc8atuxQmVeXVYES+ajGQtoaNbX+x+ZFngNGiPzHp7zzMCWe8Bs
p4j+DRt/HAVB6wTTSYQ5IO0A5Ji1k+WBVghiJup8dPUH9RFWnRNZSDIZXKkqUtIpX+UH5jwdobKA
MD3ADLwORJa1gk3Xb1BHOAWRvk9zAwg/UocYVMR2vZhqep+tcCbxQZCn4qcKcvy7RCJrvYj7As73
RJ9fvc41Iy8CT03zshTPvQDMG3cHKeteddOLPjkPgA9RsbZ4lJy6S8gEKC+gphIuIgMP/3c1roZA
F4BYYJ2qIVw3Rl+r1jIGWDaAGicpu82+cNFxs1Vk39fYCwVLCFBpppvbvFSyc/jye8wK/T1vAyPI
eNdSzkiJIlcZNXakRJ7NZtVn8u+2qykI+/7Q9HKqseEZcEWadqbqWX7RKs/e/cnelTYyQUIWCnQU
Dj6PCTuySQJQz0vDcusMtiXHgig/++gZ3G83lWCvQZ25SJnSecXODVKJskSQ4WlbqafmNxfqS3Ta
CEaEKoQUF9iv+fu/9n0I3iwWS0XNcPD3wNJ61AOdGw9qb5cuoWbiLi0tzYTa6Li8MZmNdnxCtVsl
dVHfyAfjT9Ht2Ad5dFg8wcoPMPs+c3QV9cMg7jFMeGuX3pMymIb/d3aDxnYAbRvt4e1GdT2NC/gB
aPU3PzqB4NX2ayiP2FXKGsRo1P+aXPBkjPOMoRv4opyD7OnlPrds64goj9O3B3Q1J0kyvZHK2hyP
PFSEh96EAE1AbFGMGRJgOWRTfMv0be5jcPFeMK/YVvIv7NUtiYN+K/A195qek0zxrieppJN8WfEp
ulYW2C1zRtuIGaIR7KnHT2tYtLYX/i2Ue8UapKgB9tjzF+YuI85252ECTNvikFNhckllUKBk96/A
YBWK/a1HaSoG3uL/fy936+nKls7tK3lQMSLk+N4jOX+IMxH+Ka7NhGkykUzJatQkzAuYmPhVJhMC
OhgcNKHjZOCxOBRvLY3OlsZGgOsSWQaltyN2V98bDBXQB/huDNIKb+3voxw5Ul2W94biGsEBN6LW
fetZyLT7eOtNDLS8YGB6l7ehFDgiMzQCEeJSjChht1krzMz/74Srlrv1BCDLUgui94o6i0748tC/
wNvV1dF+u3NKdetun8524fKifnZNtq00pdwC5r3Qt1GSy1enpu04tyz04JlaPRawiLa4XxOWle6V
+XOWnKUaNiA66+fplCyLbOBjcIBgphk9ESPNIqov1N3gY5n+5gnuZ+8kgu5A2J3MG8wLqsY6HZby
XYrfvGcDdtf2vJbS7b8K0sOuByiTKISMt7KFvpYJUA92UsuHlnm7Act3Pu2D6c/F2sJNC9x8HWVR
pTeohafZQR4MhXteOLFfBBAT+MlP3Xf+SocursuKe8cAw7CAdNsbUDyn232EJEd/W2m9CzFEnVBS
Ca4sgEeNeEaOkmum9/dj6ze0N2ZesmVsvtSfFzmA7qyeQHA4HxrgSxZOP7pjqw9Mm048sWDQGLQQ
NOC+zuKz8Ob84IhQEbI1CLD5J1W+nzCpUEYfVttn6yl13Jal38Ncfr+KxD9QdLWXVOqWpOxFSQ5/
UdnINR2QmD1sUG17cqszInGhVCfKkjdVpTimsH4n5LfwN78dg+/hX+FR5Atln3Ds9o/2ioXVjC9Y
0fRZjA4C6+ZkKp1bjW04BM/D9CnqwKZaeE8n81QOcihU1NcJOqN9BpFYiQRWZVWaNYX+rzCAUy9G
P/IVIaLCki88OKKuchV8m0Ah4AkVcJoFZ02APmqTOhcXerorfft7v7voLc58jHtjJu8NQ+0Rg4Fd
xX1eXE9qY6A+1pGl0NJBoChYpfpjfs74Galz21RgOBzrSzuVcHAUnSrmcqU/YkrDK0SKWGWx7vXe
p2NlTeYdrHbl2D3VsGy3kjvvTRfU8I4OB6OTPKHStctptHOK6EWnIjkB0X50K51z7aqUiccBmhz/
Tndx4ynwB+WmoVD1L16Kl7t0RYbvwhYLIVYkE5ixkKqwYZRgUfLkH03sqpdZvvL+uhKfxCk2P3aT
gifZ0P9d5msoOdjagroue2+b3sDLNqTJ+eu2CPoP/df6cP67IedPhHWwluvfln13q3LoNkSsk4hf
F5njGiGCASeCcyyM1VxunSKjQkuyIQQirsuZ/tazcgwgRXBJ0/7SPEaqBWju1cclosDslYdh6Ywd
NUWoy6jKC2sUWWErIxUT915dD5K29iq98I1vOtbrN1hmsrMsju76lmF30/OUiLS/Ef/BNiCxv93D
Td3pjeEzahCblsuv+nTzR7w4eobzLwDPa8thFJheKJ5YwoKTB8dmqtQTgH6GoyOjThUegcjTqc4b
vI2IF9bImu9m364VIz0dSBdMudPn+v/uIljTQbeFm+3O0qTndhvSCSnAfxK2tZi9J+sfzF+fVM19
cJzENQUd9QwtpQHQz6COW4zLeNLerFKSMIZL14x3wvdLfToVlo5bbFJfLm/A0oPyVcYSsuajOhDi
VqmLZ52gdg2CKEelyMdfw3Mdu8PjfyMO2j8jw3ysOIwd+LZTNbTMSk06XsJGYXIiqOG33U6fxWev
mCSuPulGGUDaTDq1RK7xB9WtMzsBwk65wgbEWowyQ2363wqpsZcBLons3TXwP35S9TDblAt/1qgJ
dE+3cPUKEbf0Jh7uiaHA9kyZVjUuKfs7rwIdVs8nhAO2nNvAW/njRUlsFBkWDVbxv4vVh21MUZsl
5fMys4LpnS47w9iPYizVSWsgMaoPNHx8Im/C0GT477Jk88YRQNflUUjO0spvI6tfbM/Jig4Mx1bt
/ncREQVqNq4833ype7PMVW0OpK8l690/IAIjkNApLUbROM4gyiK8cdU54spt3KDZ2E/v6fHRw8T1
m45sOQbPyL+g1lb74Ue7X1I596BJd5ArhYuTnq9k+VhdwLrXq+H0Y+LRA9IhxcsAX4esVuF+BTHr
YNYu8C0kWaaeZPsy/aiERVpmy7gXrzJXWH/ldd9YVXobD0HnF9U1knzuuPMlsjUOCB9fkQ7VLvNs
TXG6MRWa8ZHyoY5fBiE6GLEzPa8EQx0wBCpN9i6pMYLR5gmfkOQMOQ7GcQ8Vz0LhGIWw5ocyZ8kl
uo78F/3QgWP26RkF1TVYA1ydGuAfJFLmx3dSqSeP+WddBO9DUIh4xHZlbE/cf32OHLZUaSU5263R
ZeWTMU0+OegDYNVC1AFyHCBfHFB/0ClRqZcG2GMqNM8Bmw/jJx3Z817pi+bcYVUB4XXOcCmAV4o2
/ABC+mDcxQwEDPWrVWfWHUu7rJCIo7zGLIkBWiqbFPO46h6mUtqVq2jKEHpgpO0QuxLXToe6KVVh
3f8wabsEfwxHzp/5O1siyfH9enLSDjXUMePSn7upFD36aaXQqyjsbYEtkDuNWsnj7PHuYo6TssoC
i71jFax2ue0KwXtDhM+tDVYW5W1AcJiSgZ+66hxAg6QtpkUevr5DudG8mRMw1tdzVMKNSI5CI4ZD
jrUY88TclMX1OyNFaaikRd6fBUKvxupfUcuYMGAzcYogxKCLSMc8Wg/Z3EccwCcwWyNnFyVmcspq
ferG6X6/xeIsPaJgLHPj5oSmh/vAhr/qvL/bThzGl+3w+Oc0iuyRn1uu6xqIxOTuh0wht14gPaGK
jo17Moti6cQeAkpkmfKcuQuxh3Ss4ZoQCcK5ptMrlJZWSJBVKIjeSBk+3+gz38pGn9CtSzfWxpla
7CYC6e5AqM45Th9PiZ6ZFYWzUlo9gSR02gBFI2wx1ZH1sfUrzNT0PRtL9uuUQ22FHKv6HHCuohh/
CGqjjd5leUC7XIrcvGqgS4grk6LzY+3XWsZoM9/kA0wfBnkA0cLDXZcM+lCvtcrPRBoAFT+/lsD7
kSIRfhBdhhvxOZLuOA+ldxz6+q70KTryE34t/CiTSWTXKHMLMwzluX6ZCvrhCUdxklewcX4dn+1Q
1V0O1/i/tKH3VfFCssd4dG/7C2uadQcz3ohrycLl2UCVVYfoMvrEMQdYfg05Cettjj8bAMRGw0qp
c+H9CFdsShe7ocMmnSU7frDS6KaZ2Me8dIuo+nkYD6gP9vrRwmOrmN6BfA2BDySPJ3B0hNFZoXdF
kBErHxy+IX9cCacBymCFsa4Yaev+3FQzTvk49ZOQw5i5mgquVA/zO81aaq2oV6Q1WMXkJd0Q2PHO
FE5XnL5rNck+XcR9j6z9l8JTDzorby4LcLOYpjQeHPgIPFzeiIgDgKv22/yYUu31M/Phzf/TnYU5
4QfcUiJtIybBXV8GAaMMJeBFKETi0DXOPqkCDRkevM6NUMavlojaXVnCm0mhig6JLJIfgIidiTGN
3EzKKOsYkaZG0y+74dc35bSBSfG1+vezapDPoAZoCX8Lzwo+aBh4+iI4Ka5AKVMcimMJaqH22tWM
nXJ4jPX/SI942Ep2Hhw+44Gloo/bwfRfTxTB/E8uUMidajiccHx2b543fdpdrtGpJKqppjlhYK8Y
JBWL8/U+uaFNYXkoVkFOgM33fs+/OMmz4uo/7DyVVOf4CzBeNAAu1vdQqdlen/VoQZUXceSAjybK
PKeZsYeTvw1aDetXml7BKSWDL3Ng9YgyamioneJ0D5VcgDe+qLinDoN2Gg20Da0Au1MekFXNG5Ux
rZ30zlLlhyG/dw2JAiaZN5FDn6lzqdvn0dosUz6tEqnMNjACk0eXfSrfDTG5L6dJ9REFu+jTwb/W
/N1UN2pXdxZo2QAXIc2jNkmJ0RqFlqZK/kk8QZSa+FmVzFRPZUJffrLirAKN5XFovOvpbA6uNQOl
7RWafbvXbKlx093TlzBn//ximLSCkk18eRsegbCRGmdhaGJ3EtcxCWp4YIWWURlK3Nt2hoKD+QBa
y10vT/GoX73kdjHC6Tf0rKZa83UVn2SFpcK9Qsd4jMQgOxR61s3ydFpLD/1eNFIPIZi0AxN3LWKf
FUG1r5JVN/WAJ+JEFJxJjgfn2IMiEVgMkAnxoQq2ek9KBoLRHMq83buH7+O+ePHB3wf2tWQxP/yy
Es1blmtEkfmwg5Gr2K6hIo2ICwq4cajEi5wbO4wdGd/P5KAE0hnvr+RqRA8+vofSrUlKAdHzymD0
M5EU7saf9CxViitTrbzH3/oVn8/bTIAOWjCRj/mY6uQG+oagoiidboNCFdoW75mTB3tYv+jSGKQW
jUbRwg3j5F5yoVTdD9rJW62Ag464i5Q9leV5g3lSTNyU6q8yit9YDttK6aupjzieF606mTFzb1Q/
sMf9I85kguKDS+i90P+X/+6sF3LELbkFvq3oVWV/NXgGLDm53Fl5XzLjKUgnbKARxT+rs76hoXXS
LUQ4mb0+SQ/dhFq4jHZ7xhfLeQcQ24qkgkLw8ZefaSeguYnzSit4l1c9z2OdgN9O+O9HrsypDeE/
lhZOe6P5NZinSZgYxCNK0lFZB/EDd3cgjqFyPfD41my9trUES+HCrAJIyeZhaZWvM32p5qRg3VWh
VtQJCniG6tI9hUdl+kDr6ypq818UC/vHmb6VUrnlEEWypoFMR6UcrbiTEcZv3/F+v+1UXV0L2dD7
rXT98IqTtwk7nYBTgF58JCaEKsjlgNjcr9duW2CBcLnXheD7bEjyTUWBWENsO5NdTF2ckYaMd2i/
W3hNSX/YwrR3rTlYfKnvEuB1j/mYiVlLv18h0QUmT257W3rd8keOkW5ZlGojfVPKTZg+vtyCO5MQ
RyswFb/HgPV+vIb1ea0G0WxsvoEAHLDLcJaVB24ewxVqa+mIqjOKngVAya+rCSlxRpkYDOEBCTIu
lTb7Z+2tnHcAGkv4SCDEA4KOPRBiCQSRDANKdAeCdEoA3BGLlTdO57cQQWt0NjAEWcQOf75EFBUO
kaKPj+Ii6vBoI6z4lpcxPtwN5Q3v3+hsY/z9jQelWsJLhGRYByvQgImEZ0VkPL4K971bP79wQDqT
87S4FtPZ2cw2CZeTiEtTmANtMdnIeSuMMwi0UPpYmtWNvJRmFOWnzE/ARpIyhhRFsMrG7Ap4PxvH
4dKme+mWZwxgxzmORzjefKbaPSFr+Ewoi1rExvj7PsjejveSckmorggc1mVhlLcE7CUijQSvbiUA
bNPMegvtfHqpgFjGj+rt1cwOjtDgbi7etqDvNFjLaeu+PF0NFTHTmjNf0nh/Z/zfIyonOhxet6iY
TgjwiJdGmKps56QdSfBChNCB/gKjCGz4nzkyUrrxeNj4o1h6M0V0KL9nB468bq6/WUlxoSPZtxNM
2a0E18lo/YghOiAkBcDUk2bgmaLGbfpx8ZIfxq8sV7pUrIUKbJBM4hEKEdsN/8JsYE+aD+IWZ1CT
3DwFlspvRTzNm8+Z3G1GDa+mTpR9FrVIBrsAPYSOVySPLJyEk6ljshd2Wq0H74KuGhjJlrVCLfbJ
5xW0qzvxOgGuY5WXIFm2gyzynQvV8g8SVCPOo7Sc1W2lOoII3skOO37IVPWnmiDXuszrgpm1CBXX
JVi4ND70BnWGWeHWaXhmTACtEsDnIr3ogg7VMmy6E4Ny2y/I7c7Efuph7lRbSfvrEqjom4XLst+H
a2bocx+DPfCxNY1ZlK8JfoOkAfGmpnYqlgFavh/MObwCdFYkvVFz9m0jl0QZ/BjMhgBttdRU202h
/EH4BwEPCjcfBsO/9kU3qt2LA87U2zzRYxcGBAkd0ySlAa95BChlEQQzI0om/iXUkb0IZNsO7dYa
SxKezOtaT1Nr31/sDPYAmw55pS4VMBt3BTrun/YVoC/MpoZIql5WCa9Y6mcNKS1dkIvb73410LS5
HKTjUyRkY4zxUB4gAbdXwPH5zto+qfFUy5hu6xKsQTYmxE2nfaOlHYAClPDwKkyrhnm95IV3bkS5
VeIrn0O9hexKY1frPhrs3UTdcfHPxagRoD49wClnxydSwRMMa4AjF1XdeSCAz1jG59ljjdF9FRKI
+kDATD2VYl3K9g4p/9FY5gaMBlfedj5D2wxb3XCYmPUqCG/uXABUq9OMoiat/CEFfrzG/qYg3tUt
AK0XnsdT8f5Jz0FQgjuPmXhJ4gHc0WF+l3Z08RSLVufX9uSjRz2eNXlpBQsbeOydmkvtRSbenAN0
A7d7phHGk9oTgkCmqSxG4QTLeHBFfmRyCWcsgA5JBWbi2NfwnoGuYBHUWpchc24kIEJjjQQX424O
pIosj2sYDblvbwrsrd7SGp3GRbERWGplqZThlYeYnvJqREi9kK7AHbPj/HI8B91iM3rfzv4eGRp8
Au9m4ROjVzp083FxuoYorMBmU6qErCjJoITJW4iqT238oehsH36Ys2j3ONpgXDgyN+sGZVf4OGcM
pzfui2vYPIf1Sv8WvC/XBdT4qay9o2YoEO/v56INAAKaV0FW5Bkjy121PLZewksvdINrkNMv7dDW
M1/lPVCAhvsh2SsrLP90p4MkGZrEc407UGgyMChVD9We9HfDHG/Y+pwaDNxpA5S616Um7a05zXJl
EXyuK79l+e0VMYkoe4QMj10HEdo41n1mSboR996IEy7AUxnnVBNrU8m/i/ej8V/avqFORUdqlzKR
28nSPvzMCMbyfDKlzWUp3uM3Xl89d3vJfXeX/vFd+yggATQjghGMUwSTdKu0jSEjHcv23o3Tzwdr
j8fvIxl8qDy3Ehkwyk/YAOcRzjqVXFMBqBsdyMSaXTd+GqQbp7RgqCmnYZaQVikZe9RQwtPAo3q1
fpe3PRPI64yzbd/AbRLuU6KQUdKCptV2jGHRNskJh1z+3o04OttRIw230WE62lLYYHwHCn8o/1tp
9r8aTHEqRwyQy2+EkEL0KC96y7esgpR9vxXoSsIFIHpXUiJ6GaeXdawUBArrp9uEPW9LsAFLL0ZP
gJrV9UBdfGWnAv1WYm7hP9jtgRI/5Fnk1IbM2V6UPj0xLc4oYONcIjX+WqYrv2dhDAZJQu4owFbh
gSG3tB2S5j49FTxbGmw9XySx2Doe3bLwG3daD9/fs6z4ZKUFepS2MIZVe93CM42DXxJlubhF14zy
5q+wsWvZj1ahdJyysAeS/CMLUp0qzMDOR1uAQsEvpTKOa7Iav0321+UD1B+Mx4Y6MHFTENv90EFD
m0z3usPUQ1Vgj+WPB+GYfvGf44bf+/9Ag5FYMBVWTTKifTleAeE1BkOhHblev47X7byyEezVUAvK
fMvoq6cQ0PDI0aEHDd8z5ZNPfEJqWA6CjBfd8mgWKO3m3O7V/3ewtxwICw+MhFSS304dAA95/zhM
pr5mDFU60N/BHlTCGPf1YQiez+nbULs7fGaMCtO5ZoA4uSbzTbOfn7ut+T38jotC/gHCwXrkQJkb
wgZTpwl/KfCesYZTf90ZHeWaBBA/AZNyg8o8PwuhT0VIhH8u/23DARIss5hB/JAP5+G0fOIKqI7D
pKwbx1JIvOut3/FF+i/eKIjG1mOzNxrKZF+iJ0qb0753sDyYVMxc3pI91KhAC3zHZ3bVNpRRLEPZ
S6rShJE1g/k9gsWbm2KfG8wg+uTrRBJCCm8OLnN1OD7a/msBjVmTDAqeM5FJ7MBSiLySzgh7GNsM
nADKd57Weq+Ps1viFcKc568zSVI+lqDEr4dqJGUtj8/IH4/5Awr7KAXi5Yhdj6OtUiX/IaDn5Hf0
XcI7lnMzNhC4qCVpCKRHhKhjyZLKb27QotGLsEuWw7duTB1F4DLWZRE0bYx80diQcv+Ws9JXRTq2
Mn1xKSvhnK9YlygLCPy+PtC4NelI0G8PMTD5hAmm046dwCzOwSxLrYwBQKIsmXUJrvaHXUGIfBg4
ZLbgzLPslTG7C0j9nAe5FzXGuGAcWRLQOvPApGiwLqmfa4mEFo65lyJFBiAqDMXiZg1t8p995fju
xkIBa7lcVgNNP0w2926P7hvy5M0P8Zbs/iZstD2jzaiWdRwJl4N22IAigtrfjwH1xqJ551coGAie
AfaGTX6ZqZD9clHEsyKxQgHoVhTurOPWT6zEk2CEtrqiMKw11/72wJk9oyZZMBjSjYPSZ9uCJxv9
AXDCcaZM+LrPa/oNsfrdlQbiJH6oHRgTOzGAuiOgFHGYZ03GtjST1TrMdXwRRue6vqenZu0Wh7Y2
t2ZQnR8a7k9zZnZlUGxiJhgJgjt/NOGt1ozj/fmvdzDIbXPLA4HBOx5lzrIPetHoKsRnwSvz2GGB
DpZ9O42dsXG6w1acSDsOk46pEEys0pS3HXJKtJnRNooOag7D2NjH6fP9mDaum8FKbqfJ1mjLVXwm
aXTDT67bkAa9cRiFwqBP9AXnxzU7LwWwprYiJmo6wpcdYd+Wuu0/MLFDh7s0UVtul/JVmrAJYGnm
GcMSwi6ECqk+J9QWmp/xVkez2rx2QdHADqkQNPbBVmC6BS23GSnnZ/5/Are3ByxkyykfDIvyIUz9
qaNcb6V1MIXTWbZjfPL9q8CGbHaXo2HIBMR41fSUDxfkWJ9GKGpTiB3NGP6Y0jWnwEyKyJYD/7GR
EsLoCiou4okmG4K/W5s0ZfzJY3VDDhvU3kHauN87S/bNYZw/PzfomWTN6im6igiNET+TwpMN92p/
84AYBqO0bgAzW6cKmZPHnVvK2D4sm24haK7Kk6x7jJVQQnTsK9/Wa2KD6IIaf6A1Mas7PprzmGOi
Ru/22LAz6ZN5qK1thK86g/4xsIz+QAjWNU6RhDk8vSQCT3bgTak0kRdOZ3aNQ6E5kzVfMCSC6nol
kx6qN6tnPsKIHmAcxWiSFCBM8j4/0gZQzvjVF1u9orlYN1e61BaxmSk3Z8HaquJHWX35ZwfFJC4W
F/0kZvdwRaOae3VW0L97ZHJOSYw2ODIH1CWyY7pUaB3U0Yoqqv74SwStKjTOSP5ls9YLz6D4GTBu
o8fElLnfxLcg+/Z++4sQjeJ95ymXTAn3x+t0KygL1xRaz0pilefZCRCyuocCxQqGM3jbnvQWFgFt
3X4CN8tGg1zBiECr5t9YckSf03haNJPB7VkF0kBQKTwPQ/3likPqBWuogpEhue4GWKWsRT2ngXrn
d/InDJLOgnKuBSR3eZYCt7Y6q4fpNkjmmFVvDtkuBvQmbpxa0XJIaLAoT4S91NptaP52HyR5JZtp
/9fga1+W82ez2n1RLWSbwVn0t5PpRIzrFLGrBsaIBvXOE2GNo/iqvTOGw+6FtavqnufuZNrcs1T7
il5fRZyYXi7ojeXf+JgLWv+O1dyBaXS/oiglkZwIaWCeaxkl98L7YtIO4R0WGdBx1xFI2YTMScbi
Fv/wGTDFT+dV6nPLM1OUlRpODzIoCLBaoCVLR6dMPm3xkPwLV1/aCEDfTs0DGanJkNfFPC3yyJ3T
b3EXB2xQy8FJYfutnSFhRwuWAfvKLUnh6Dh3aKtU0jJSlow4mljSPB2SYVuETGyhOT4U4kWZRxIg
uk+hO0XiP37teVf71EhBcfEv9J+5AqtcEEaAkUw1FNqUwIUGp4hZQzF7YzjzJuze2Kdk755CN6Sh
duKodf2pTy73jeFFyumYlfBpcXrUOjjX/P/2Xc4beQvCpTmEig+JBgJdxeD8QQJMBXWrOtsdBDfl
wbZA2nUUeFUfraTWqnZIG8amgcucUgQe6OfrKXDXzKWcz9nEje+Fpbo4HbZnKcIHYa+5FXeU+QR1
Zt/7BrlqVXgieRpY/+mbia1Uyna9CCZFqrWUFJHJuXSBWTG0OQJz6yp71urdlvB03QgJQ1Jw9w9L
jXX+UStLsLl78xaqX1yljpgJOu0RJ3fu5e2jBGudwcqL7uneuPX2j5To4cYwOlPFkoqIIAVwSLyS
bkfnxnNgrx2jN+1a/wATdQxrzzQnP4wWAGf7yuB0ruQI6ez/owiP1AYmDfbxVQ/nf3vGWqWuztUB
M/wpMOQErURIYRv9GUvI0zCVj3lmKKOPRpXSWhu21si2H8IEhOhT96KhElUVL/Mgrt/FJa7OULiY
sd1JBf6oP5nvvnF8LP+GDUFKzer0QW3cHoJUrbXriAQzzZMEMS68e9YWR4hFl2PgMT83FXzPxtBG
A7JB84+3LbCAUbsv9XnzlWX0Zl5ZpsSi1+UJiwd+GFQ/EQ4lPIpPULiDzwYngyLLVyFETQBAjQer
FUR1jzE9yc0iDYeTr5neI8q1G5crQq7S0bFbha7GxGLsOhEwtRq3ZPs7a6P00HF7bYH1m+qZpAXS
lXguTrY2n/ovyvgerJPM08ubgimKtJ3oZAKqJ5j6rw2WmH0RVI4si1yukhYR3qcXgfNHOVuN1w5w
cwPPwScY/AG8NQO8jqSWYsYdb/fOlF2s2YJjEgeDDCHgcRxEbPrpZSl7k0FO8+x1y/rIonqXSohe
djIKsqAtZ5J3KBcTrtCGly8bxcur2gQwfu12dzLavANnuO+pyBNcW2UhhgASgKnG5haiqTP3wP6q
kuMqGiVTE9e3zJuMWSSD+2oNi2wqWad2i76W1j3CraKgKgEsC/cvtODUC6VVkaqYSr1/lkXcfO1W
O5Cb01cTI8b7skxSLa1/JJopqv14KKPOW8u0ywS2VO4myZdm2tFvA+eXnJESvL5qOd35J0nMApbj
i2kswLbenFSQaOK47MDbvg21nc9yXR9GVdHqZ2vFklKUpanG5DGeX6rT+QdDWs9IZrUYRfhrSWyq
3FP2tM331DGfPldutAKEQh68nDOqwxPhgM8SuPq24kc+nHyV6y7vpJ3utLiltS8EDXSl64Hm4hhe
6Mqp+S3cLv0mG+EAs4wZFCM+istkGUDw4HZN74h9edSpRccr+PFNJ86fnBW7q/UEUY+RzfTXx1ek
yHRkXhuVfW+uNtuUEYq1I2UTcsYVDy2sKWyyLUKNd8QlP3VVfeReBeXgTVWHx5gfNY3lUS60458q
7Bg8HcmryiGuHvw1cPZNTGUQRQ3S3PyRFgl7gqJ6/qKJy+bqYyXwvE7Moz1MdT1g+yE/gbjowsgN
/Lk+NwhcpF6202l4a+dIwhMnZdmS2kImHnF0m11x7oV7JPmXibQ0OCUq/VCxaYioKevwsURE5kTa
NkNuuRQnv6UpEba9x7oflg60gGBZWq8TXcN5ig1Rf0rRw7GbwH1Y71FGt72u2YWFvrIo4Ola7qsq
JMaPA7enbE0fh4bvJeMIlUYkCLFdWr8YmgyRQnaMaFJwVDM8unsTjGOr+VFoRiE5DF81FWQq0aFo
JvpLxIJNRsesA8/ijJh4LJ86xU+vGe5RtPOBn44m6VK5nr9NGWynvZ35sUS7HuZ72+17zgXUzj8s
tyV77AzQ5tGEjipLCqnXfyGNIctSD3qYzsAr8W9t8PSxwN0tpXWl6XbB6IVvk5PEn0kIwyPXgdpq
QSMZYG9x66/5qmeS2svot+zLYv01j7N8U88WbapEuvVbiz/wH6R5OdaMCcn+z001gk/BCXQF6RWs
X7udXSfpz+Acl1LDu3iBI5AEaqQHM4EuS/5aUGXtEEY1c8QNwqwbvOf8ETDnCuP5D525JJu/LL/d
W7uWocLniF11co66XEF08l2S9A6TxnMhwfzs/ukzDoqfHDBAIKXZXupkPn/TWQX7YddIB9Cbbri+
yx5iLJY8skUOHwxzfbz94pFsNVNjZhBO3ePc38IVT2Qpd2Ehkk14qjz3B13Vup/F7NGCJ4aSZvHx
QGQVBN++lhn1RYEStC34pCyns4IxNay9zT8hgfg+9nQnLYXD2KZNE/i8eKnM9Arn7Jr/gjVXoaIo
aXAu+GOGwk3mNP/Wf3PZrfmyIlCnecTvKHArR2XT2l80mmme64n9WkhCDdtybZw9/7WK6wp0x6F7
3hoKFTXkVA1I6qpZspB6OQVrakzsXa65eX/vciHo5w3ZmPixU1cQ6Mhk6dnSlnmxBd0+WQ0ouSfl
T2B3ECkY2eZff5rk2n1utmV+FOmbY3UPI3nHNhm/yLSBE4gMO7VMAt43OyLaLEXOJCCiSMMxQLdB
P8MbSY9nkFSAPriKNE7LEaTB8KbyexeKJWzxOvQ2ILyjcQZ4VCUWiQqxS+qKmuRJ8WeB46qB1AaQ
KJCPF+yWb0Rj4ICpu6RotFzP77lDGaLK74YvbOYux7TZa+VMfcb/pWDAuCGHRmxZ/yg680cE00Or
1pDSZQ8IIBWEtdFRejdr8vooJnFqp1Jt4XPMiyGimeKPogz8qXQxzSszi6dJai29vwk6ODkCS3D5
9llL3OhN3ebzu6XeyRtCfz908MqYwtL2VW1OZGlwhWz12nHOCdv1HaUmjLr1CyiOmtNfC8S0xhBg
7Ak2Z1HA893vqjNdE6oDx9AH8WWLgqhfcxXsk6ShmvIx8x6Gip8jKz/Eo4R7PR8aA8sFV9Sgfe7A
k3bD+lk6J9lioPph9gu03va8z4IMDhhYEMB2t6W3L2cVF9fpnafyWG+kdV/DBA86ruVoTt1ePRH2
XRl1LgSzFaGtnktMtunmxHS1UVXYusTALR4MmfDTb5P1uurN/UcELctXH/mofWB3xh3uKZyj36Ek
HbYcUGjfPknIrNc4NULg5fCf30r8NP80+yR0z7rvLIlIpRqrszs38/GRBoKO1cbENYQ2APSL2gMB
nj1Uq4jdsh6f/QpPpv5v+Ae4bAxbltzRTuXybWvBw8060HXPILIbHk8pggBO6J/HQmlo4GD5CNB5
y87Mfnyx9SMHE0AFcNKV83UiHYl40Zk+iGVnb5GwkwsrwAI1Eg5lEX8ZhRtEiihVtCSNzFwyBrLV
URC/A0RiuyDWk0nqS1a387Xg4qHDhv0p0yFF1aaThAHRmT1AxaoZ/VrfTxA/7C8qsajtvnuTiC/6
ltQ2ffi2gDmh7VRq0ocel5uLQzGDRfb14O1nz7MoluLaSYT628Y7ALUYGDxQ36hYP9GRBRv+pqhS
/3Od1+CMP1dulJJxbaA8++jMk2P9dfn7M1GmXCse27ScRMAZl1UcUOeIt6v3KxkpB09TdEvuSmP9
KhGow9POB1y/9QFtg377Urn/FEbzg1Bsh5sYZCikU8KY4oOWaSe928Ubn7rPdO+pLN2kAyXosh/s
fS7K9rDOZC6Mkfxg/VKB/gNGqbMQPxJnL8qRhzy5tVneC/3Ra7VKDtyYPEFMNiEVOCika/ZNMNRV
tet/Twysx7DLwtevO1sa0/B9uM7qJl6Zdu9PiHc0sa7SVCx6rvUVVFAHGXhY2kvJ3HEmJYwR8h87
KsVrH7AOcMWGg1dDCvUDHaax+pqPiUPfWafaAUe11NEVpSFS4F/XIQKK80dZlzAk8kD8vTC4EKpX
hhlFufLzZ+YQUN64HqjvF+4byXVJAsIUs2jwk9SmPm/43quUDUaNQghJ+hw6sQasRi5JdY7gTBuV
PgF2gRQqqlXij4pKebwfHZtEJvWWAUkdWXJPqv0qhXGcjiShW/7Enwq4RrcVBEQhrbePvrNYib4w
osdaSKk29gA9eVXU0bYgmDm1EjCc5GtU6n7FI/zmVySJ5shp01933R9X5ic2yZ7GmVqTwpgeCo7b
S82ESN0N57ixtdtDVELFLLTUwZcxEf98bUN0ztT6Ia7jjaLfKdX8z/b9wdWyURxKcazFRFvsFGHf
EtmNywZPreNbQGY3ANUiGlEaC4A2KSeCvOBCANcr42ZnNUC+o/wdKpH63eegA4Ly3TtpJnlPqUzA
467VbiynLDnZuf8L+FyGat/RfVjEwNSjjlmiLyHIsOczgI2aHLv9+7ZgaGn+utxCswyc3ZBxFmHM
coFaedRMt/oVSTiHrY0GHN4g/0KOcu1phR3fsETf41duzGtJjc4hFASZiH1cWpO96C49AfqY+UY+
A83ORVAbxbgdVla282Hnc5T2U8hWZqmtTOsyRqleZTnvYbQbYBW5NhksO9EbddSeozaAhAaWGGtb
vtczxXzd3yu4dxcMEjClUplgxhRLC4YC8vw6qMsG/cIVVw1gfXY7Vy32LdBIfyMNTP+aDmv50C29
uuhXiaRP9lSa6vU50dTugs0WXilDCdgL6eyRofN73kqrQRKkCOBA34iESDQY/fU34iKvkB335RPs
MSjs3wMoOSI7XsNWh0zuDhwfNRWb1P7WblgP6dAPoRneP4T5vD2zoiKyzquV2gpjisXPJm9F7OnR
2lxhIhFARm9WswQQzHFItSnVQr3/cpfUf3X/FSY0nCADCn0ts4d+kTb8+7DErWh7kK3udiYJo2aK
NCT72pqB2ZZmZqbi9svw/u8+WFvwEuLJ4+GXknYvam6IObgh6TsRObK2wlGiMNKATIebCv4vQSP9
Imp4ku6TqXNXgfVUTtfp4XbU7+jPp8bM1+NEZNJ0SvedPCcFCwE624lqWCjMk0NGM4rGNKYtmYht
559lCLGU6kAIthsyw/Djec9mDJvTzNK1hOBVmtE3XDGByUgVVhyl9kP607IEeGRZgppA+XnaJwkE
JB+D5HM403tBjbnDLdRnBfsJ5N5C1rcNT47oSemFdPyPNAF66JlfAZ8OHLZss8FVJm9agMGRrEtE
sMsY8QlxgHCdr7lSVZvxpVPZlr02iY1TuvogshtKsTcqpIoxxqr4zxik5RgtldqYpFm9h9DtsSe1
Ny6VWjTYa7Cqar8aZCTKozEJuFtPWvplcuTNG7X9Fl3SCbzxFbwPlUKsVWFzdRb2+RU8z7DhzbIc
fSd7dY6dRcf3tE2hagpobh1we4dBqIKDKG8Mbmcb28W6Zwpe5/ZRzsUt2XMknF0xUzCfTgT+zECh
Gxz4m9pW+ZrT5hmBzaxsm2T7gWoPgTfY8VvxVFV2nGgCI4O5FOM3LyYqnJKGjnVXZZfwVIy1sV0P
hBR3cjz5KjedOo7/lS3Us7Lu/TJwizUTV6m7tobaBLEsLxQbbMN0pyBjDqvBLdPe4WQEpydzGS/4
HtXGDvGoodwKD7E8l22+TKTgfLOuqTBbqvYMoNqmFVQiAz8yHT7e48k6ZP3ERX5JgM/LLorQH8Jc
59kkMnpv0FFNEgV4IesCLD4yUUXyFXgaoOI3zEWhMovtpiKbZ/oWgH6mSQvnpcXt+Bbt3c0r22pK
EnCIAjBp3zpK8N/uf1O9JKMqeTWATOPw/59jUdxF3dIXZvkbQk1ZN5s6NjCQ1bGdTARw1tKpZ40q
1MtubsD/9BvYOjao2er94nFpa1SYKaUJZi5dCif20DDsOjh3OucFHqlZXVgC5UpdLzct31FUNrSi
bJn5gp3KSjrYNRJO2An2vhBEh+ik1VeXbIZ/gCpiXZ+TzrebZAg/Q1n4GCAYtjFtE52AEUqpHFVm
ZZw1FIRnbqHrLh+d+n8dWGjGuXFS1hRB18M1B7s5frdbWhB/SPwrkpTg/mOJRbhfYg3+o0dc8oEL
uChEnbqzDCVwkiZ+2r5bYArgHdGX9ftjfVIzDk886oxzWj8c91rObfJ94ZBfZGhrLHZIepTbvy7o
S67G2UG/+OwGiP+qBY2oiSLD1IUknl1OI83XQAhuAFA7udEA4LRXgjRx/M+/R1OQ1qw8fWd+yWul
oVupm8I8tQxmyfY4Av7JQn4Xlvb31fXojlurD8HfQZRDLKoQtp9X2rbJEyrpLhIX4V5K+LYqvvzB
MRH+9HLN9Trsqy97rIYbZ/JBdOTSuaEqfvhSoL9c3bMUAr/GMwKIrKqzOy4k1vW3O5gErGxtRR/e
lKLEdBG0luHzjxriJj83coMSZ/+rSHBpkVFSRawyY5AwlhTLFMX/hOiXKP9NdQVDrzhYPs0UJgKS
PsGsLD6EWDE6Q4AgIvkT5v9n2pw86Yc9B9wIwNds9NKL99otrdgcuQf/S7kRCB4148j5N8nKV1Nw
f07hCcAiEBRjrzJ0ZuYN+Rl+hVlSdgMc7qttV/abnAuVFSEn1guLrci4KbI+Mfa4l3TL2HIpTeK+
6OmIzUgnlOoGr7mhDBTYip4yGiOgosG0j9s3l8nHQWyYMphd/DgS4AQr01+pUdrEdn3JFvQXui2y
ccYKcngFVAuLC5FfN5FdsvwvC3NEPc4qaaf4eW7eUQXAKs2zhmJC1HuXWNoakQKYaaeD5Hwbl+my
F8EBYDUgT1o/PodVN9VoiwxfYn9uYI6SK/boOCfBmHfp03pYMQenjIgcuf2aQmNEZ4fD7TVznAVC
RQx19crJcjekhTaaWNsuo6lzN5bQU4ITYw9KauovqyqpxkyGTKlZx1tgUHrF8osqigRFN391Ix6O
oBk8gXet68L94ZRTweYUzIHxy70JOkyCbY0a161Dt+RYhQHMjahvgcBCAvZjC2VKPZnMcm40jvAp
i/ZllYbrwRlNjHMlPaI9edEprBnp75nXFets7F3wni6nhF2LEL+z3It5RiRlQ/YGKEQZFUf2g8K8
lo/81XmlYBHN5JWadEHZ2SsgJ+w9Zwa3+8nJ1I/sCsai0lnY7ZKcp/pbm/PkkmzrD7bVvSgqMKAB
c+yn63SVnHn+8VNxQ/VPw3CBFPx3ispcvEULVZrTrG8+s3p0QghBmPVj4F5VSRW26D2iOO7CH96c
xzKGLX6CzDZ2vmqhoXxQfJfzXNR7sO+EjkgeTcV/p4Bxx3YE3Jjsh7YxBBKp6HxyUKIQG5DcBc00
Dko+G6WfPrH4YNWF0SFj4u+HPOPYGQ/kEbg2StfsfS1xehHjNZRQXbbBfZSP3xrKzYyWIAgewl0r
Gmu3FNVQavQy1P5/DZuc4+BU8K1eFAIHxgzpuq2JOea8EAOEleDDo8D9J/c06g94vA7376FjqLsG
v0MIqpgUA++FsEYkP9yzya/4dbEkt2ipieOP0CpbkFBBAg6Pdg9gB451WUlsc/DNunUgPZ/OIrNn
PFgW0v07sigy1Y3EXtxo8vNtQ3BxfnNZ8+FSSXdYzvPitkgDv/E3+AnYHD87s7H2UkDxcoR/UMQM
6piZmyEoLMMR8iJe7s/YtHMMQwxVpVCHBGwkYjxjt0gYVxwDL+wV7g4+gobHaJPFjL/k9+YkiIQ8
YYMFsEcKmpjrfmJJ1m6Bio2XwKaFgXLIaji393XZPV0Ha+Y/LOtt8EQ3Gss8eTk0aAB1cuklHjU/
d98tPXU/WpDbJV+Pj7F5Kk5gGV9a2OpteWgSNngrKEcxFFRplLV2RBH+FjpguL+yEp2GjJzU7XYW
5m2hI5WIsuo+/zdVM7FVO75KN2CGZWDMtDRe1bLsPmxqI3amblvK/s3mMq5rv9rmZaa3bDP0WN62
7Tqje5Im3YloRRinsXs747M18KKfsnQhukVIySjdTVoee3olo4P5WgCrxbwXkWzlxR89pSGFGBkU
wh70bUmfACeqzfB++Adr91P8T5p9oTZPFDXo6cvapIASQGlMegq1M7pIum2kqkc7SMW7HV6ivMK9
bg0miCpTMdC14qONNwb3xDvja6NV2of/N8pcDWIINFDoxJrISFd4hVhpClyLvcVd0wkXx1rcYdqU
XAglBJZMtEPBB6LEMhOOgjovqSh5MFUgLXsmfdgIi4SFr6n7ifsxxtib3gZbipyMoYYd3wABMg4k
drlNrzOxmJbgcQlXYtZJo6T0mkio6e0cofriUferIgDmC7r6PaFMxkm0qiSco6v7NJl6xmn9Ft3z
L+vSHzFANSJhM/W8K8D3BmB86ZpTEOWwAMPNedGLAYpVyb0hgWd0muzOstAffCrmFnQyqzjqD4LG
+4rqgoyedYNNeUZ3DVJA1M2KMyyyeN6i6gUbgqcni8uj8xWo9JgB+ZLMtEtnDCwOjS+WYWAdhs9k
ez5p27haPELZOGAYMa/r4bEP5t0YESz/yOBEkIfOYHOSTfO42NAvgC4vLYMY9LqYGHIkwN4O3c9W
drcOIh8lRB32/C8zS/oB3I0J9Qnx52gHXlxzB6nHgfDNdrzJddXhExaRbiwbAitPlmM4qyfrs2qq
xAo6iza7cjNjhAm+Jtu365T/oaeJWlEzOJeBhMeG9gntHzQAcyGUFDmMcBV3n5US+kWlxp9wVZLo
Q6yawRJbwAa083ipbYt2FPW+ovlA2udGv2nbhtZc9mr70t1NONd0jy7cAje0VItfIG5cCBOudJRV
S6ShutdkIkS5ReBa6wnl3PgzYXTrTup298Qu8tl2Vr/uJtL41RXaO0oHLXaVmXXm/MWpz8tr50Fp
SQlpby9qJVPMCNaL8aEHBOhUoqjA2HX5JDI6KpfZjU+WUdQefHYuoyRcym/LH+mQRHmbK0VEMAKw
FVQrBXRzLKI+XNgYM0PlcgyUmdqANUvhnBAeYPeKkEuvqb2IoEsYrWJ6BOX/Hp5TMQMoovcEI31T
Jbm0yVirIWYNfd8jYQay8Flktxlc7jcu1xrxu5eW5IFkO5ymFkismH1bZajkqr5wtQXnnz6A2Nzj
1O9pSxq7KgtvQoB4yNo7bEiQLaqsNoN834amwR2FwqwfAGyCYNkrcfQEqL0ALh35oeks4uIpYmz3
f2SG6XKSHtjS2sq+gVvsypl5Ms3wDxfv6BkX2cuwfPF29aFZYlYuQrwvZW4do0ylfTV673lfwtxF
oCq/XCrQNIjy7Hc7nCc0AGcWVTxzO/ny/UX6RG/ahfbGX1hpc/yt0ZMBCGin/zCrfWf/m8hQxeYR
F0XjcneXTN3WDh3DGOHlEQhSciFuu3jaRbiyr+wM3KcD9dnIm4XpHYXb17eu+N8QRUnlxCcQpxwa
KGmSZijZNFnGdWwwbK/xUKGvSjNdHgHrfOZ+yBz9oTTNIkv8zWne1yBZdDhZ06dKbBciKpj3D9Ch
NqXaF9VFiNOE57J1/ZQRaF7WoV8LRpFu7f3MSS7BOodNzs0p1iIkFTWUIg5zraUDDU2MLzER+bG/
l8m6+PsL+rILHg2nLEs9ITv8lWk85McoBQ+isbaGVnOnrHQDAD2jSZl8SM1mCEPe1k9XeNnBukPw
JWspQ9SGyajpBPry4eetrtYRpTfAa0HoXLYlbo7QJP4Edd3Ffye4uosDu1UKyRER5d1N7QMlFYdH
E/I5U8dnUX/EghFLJR2PF8ZD7Yp7/2aXQksjdrbs596uxaWe0B94M32gyeHEX+gKxzT1VAHBBfjD
KhwDWe8KzXwbY0PYjOHjtoF4R6O3JpKb0HlL0O/SXKEhf6rRT1FQAy/aO2pR52LrZHsTsq4E5fPW
xpfquLikoW9jV5H7j45T+xIbTXSfomMZz0lrPdqHv3H7fH4QbnbJbCZlBXJccQNq1YS2rgIPZ+wh
4o43nCkgdvOkqDnzPrBygOxmNchHrFdziPHzH3z4dJdJbcQdN+VUdKVFkGwzXCC0G7iWpBBT1bfB
1nVPB70mYx0wk+gfAgAKcD/A8F88rocOck8smBlj0bSX0P67HbtC3A+PJSb2EfNTiYy+jyyP97JP
wPpKBYqC+AesyNObZ/pMXC4oOqoMMMivOfk96V4P5A8p2qUsJZvmpjbcPRu+p6h4ohxY03RPjM6O
3lPjYrkq3PdzdTU+wgRnXWdJZnNG4L4caMeQfbemiumR2PSl8N9uIIZbWwi3/klrw8q/4h+Mqk7P
yUluiz+rTiDOeAE7tp3IVAGU1AW4bwAMMevBZCc9HTNYg1/RpAXykZtldFRwpIIxtmLB9wo5g+M6
gtMKADD34yqdvItquKekxNQ5imn1MXArYBmit3xts6MJBz8qyXrp9bW7mgQZXlYXSQqLTYLRAnL9
QX3f9+kTi1JDEtYOZNinNHDpvJk9PfTtbedUFkl36Edfam62Fawdq62QYgxIcInorWNpf31iCp6V
+M13JXLm2qFzHmX7ZguKQAzggHVFi13t2u4lGJN/Mvn4zHput9o5US0TQDzYMlLz0uAJko1QWqrw
Yv80kuXV2sXVVBfktdqhTkLEYolzOg7RsWdgVAKhOzOnpHj1lPxGDylwTmjajQUd3GL8RXncC1gN
YQjnGVAs+hxJNejmoipI6xcYbzedprcfqz57VnXM7GCkiq6U5XZF/aIFbhtbr281I1fGuaEB398f
+9bl08kSzAhCsAeR9D7brCgJGbIc+XwEKSTeWESLpOkDtMxpc+MRaAAwHNS+it1NcZaR5ISGgkz2
XkIJrvbAI+why9RWrqvfqYAAXVWkUAPBDoCBAu//TKOCa4UrqQEcjiZgyU061pXYuC6QfDHpHbiA
WHLRoxh/OYOKf+q4GUJ/bcmaJBDQwwKsO6EXBaG9c8T6ajuDaQnK8rgOZuRRwixYJC5OP3zN/b0v
/AgqMzKjincTGxIUqiMNiqOP5oTD45AEB4xvGGk99kAcUQCo1cw2Y94++fGEPusB6sZg2nwTe59d
5JGPo+9NHn0xdgyiiUZwBtcDBgYxPtSc9ljsG7Vxbc/JLYID7NpV32tj3cVBhK+UZr/j1adRhRf5
kL42oJqCQtbFWdau7EmtVSQHI7iexJ3j7mARjdLhkSO9dEKADkcFu8sccWo5pF0s2PWb2vHwJ6p+
hWeKoOGE6+RnGpfw+Dz6Zw4S+gmi6a7LF10ryheyTIPwldbKfD+1lbSBdeg+2t8jfn4EFNOTeRGk
AFVo+WPBL2zUscIBBgZoBSeX3S9QN1+aDZIjFZbdU5Q19VngYD7DUhU3767e8uG91wA0MiuL4KJP
Iawm5SB8g76AEvL6ntifDuM21VfKWusqKWxZ2msEYRLEtTBd7Epbz4LfaYQbVFsyXWpO9ki19C+m
NRSLSfVS6feZ9NImLN7nX2mPGX1dfriYjSEFp09GRZk6c7r4rWjJmvFCxIbdLsqU+HcZ4hkJNlZ+
gCSx4Qn/DWH+O3QdRnBTaCj/jpj35hEWYzerbn4A7XoHFVVTQRbz21bNreQFL8wMiDMX/w4y74Pf
3ExAUi0ph72hAn7MJB1FPFC3jJX016IksUHuNPNVRvvetw1hvznmoe1yF3/08cRLGFI4Qf6oqBr7
5PPVdrz0wfG2EnRFqwfi3tbPJqkzJ0EiqfXlNPqpAl5EArh9sYr1fH3foKH9IsQE/DoCN9l93qMB
uOhMhjQ788IJreLQrD6gjRu2KxVwgwryKaZZKS82d/0OsOo8v2ERxtPtHG9OkVTBzZH/QOaVCKsb
TaF2pC2TMl8OOgfUk7tKtlI+VUi4S11UxC3Ktf9TLrMLHRYRBKkCycNrvPtoUgWKgXgUWztJfIEl
zDNy//cngCyFLbUHedPtq8UGD4+Y02lGZjqmzVa3/cGXdGZC9g2yYFSfyxY6yoW36LGo6GE22te6
C/qtDkfNZ7M+RrOo9Gpye0+HHReppcfZMa1RrQJY8mwMmGbPBzxZ9wsxzhgQhjVD3nGSzJWNZyb0
IlGPlPRjMo1PdFy8ZmRRbNKGP82ihJPMI+lzHXgBcJXOG3FZgDfjXRXt+HjGpAg0HPOKS2R21pLB
1lLRPoLy93SK5oRIAuK74P/w8igTk1leploCnujAYrnCzeHy+MK2K9zeA5tbJvl5YEKC1AKthjZH
vFduBypUNGu3wCsEbfGY/OmKlVsXM0+G6NiB+HQKCPRglmgPKe4YyYNsB74PRI3RxVKJJSkyCwQK
O5xUE9f+HUp8yh2fgdK/MJcsycLkNDdioWc2TtMO6D4edn7mKMw9gOqblnDmikFpxNtzHuwym0DK
ALdMcHgkjLbzbK6K/mhqc9bLKR+zSoCAtbsm61IhxJzXlq05gx2vDYQHACMJKbvVSn7iR610y3HI
B9FAm2ZbdwZWHCZecss8/4peAybKU8FZyM3QV1PCOzosz/myWdUjNVKbQMsGsgtlyytQFzeDaaSD
J7En4w8iheh9MnfVcVFtvkyQyTrweqDnn1bZ836sgZmETnNl+/HKiB83W8MIz4Lvv52h4iuUtL23
oam+L9GPy30Xs05prMsb0f3TymGzytMemaf3SEB+WSuoTeqyyaFiEaWzO/LoomzHMvRzUnKDwJRC
45Wv1sY6QR88HbcwmwfigdpIJtp4DkZDQEYya6tkn7fa7+dp9mpnz13Qi8+RM9xzZkSjzGvGMb4z
5N8zogIHmqRay2xQqHcl88hqOWfbFXgzm0IAgHtYM6/CF+2qsu678iDiPS19yV0valtraUmjL9D5
8hk2dtBzXA4VsAZRHGqcqfK81Thzye7y9S3fwXg9fkWhKqPCVSjgz+3Zs+ak/0xvbTSyPUdqUSke
eYex0X3JecFBhAh0lqJXcBzOc/WYHn3vUyeoEoYzXU7mYCcWbjGXqXwsDvoB/Zb98rnyqY2UyPej
gGpkaD7jNoCR7WvACRnH8zu1EAlibwixubI/TsAif9J2WR5qt6VZ9DA/J1W5hS5dCaAKSThe5Juv
W+S5N03LK2rALSX+ejfKa5qB38mX/K2SCtebh8RWqSR8TMFxY2DR+Fko6GfDIUxrg8vEz3M0gQkv
+UNNkGzotRVysdXQiHUBvoirrODbANdePJdUbbdTkFZ6nufKs4325JOju+Vvn/zXYmtcSpDm9fb/
98N3VcPtDh2Mw9o2NWXdr08SW2aJOCjrpH1AsTqM6Jq2/rHFaYNMK69s8aguDTHDkrU8VVMSAUbk
smYNmYmIXtJEar3jUevIYJDig3NhaBJp9iG1UUBDsGfPqUarDZaGBd8oTC8dmvZhWEyqaBN61rZ4
S7jb2jYBmQnSvcpUt6fp5PXAeo8nG8gU5EzaYg2fhTj4HPb2idKTd9CWw4pYakIaFFFKyfbMa7G0
tbyzP5rsbr5C1z5SluA5G3xvSQkgqanrwqSX3RrgEFcLjQGAVcvHe5eRZg3YAWG5cMC7a4V1PZn0
swDkotDhgIhKfDZCMcvWdkeF/7kVuk+W2lmUa1gi4PVdcwWdDl0vPzvCb9LItOyGFSjZ6RfblOrP
XJ4qMaHLaaZCOhBU88HSm0tMWlvRoZC1pgw4oICUjZwCJEWYwKhyzXaXTT9XDD9oEgyPj7sxvR68
56bgzBmNoh8NGBbRRGebTVtQl0j0L8hgNyQO0a7ktMCxrmZJJVw624a/5kVPA1NQrl4WmGV7Jtn5
7hRShsmaT5HDshfKBuHMUOe7zXHlUl0bStym6hJ/N1NJZp1OaUHxOWNUSV6ptNDP7BGlbG+hBl9x
ohqrwqphAE6pho5fqsZe4D1xE6mJWp/8OOEjzTl2iTvGpgJ6RvM078SEEynMEU5lBzRl7zt4HZz5
64O+H435hBX5Q17ZgLjJ0lv9bDabgM8Fpti8gWwYiVEIkkt4B1NgP82aZS/ra37rqrOsQnRAQQS/
KTBdAMqJjLfv7k3jgd2liVE4gRVIJssB1vm0WKMNsT1GVyR3EJXvJun06qIJZNCEZ1jUgHEO+4ij
OGttgb+YFa6mqp3JxJ3fwgMZ040uOzDHKRNkrEih0DjEnqjyz01Gta5WsCH4qXRGA5dWVZ2hpg4P
0StA/kSIwVnBAJixw4Rff033O06T8PgabNhHvvCCOsaaSj7F5fTH4dmHp8zHPUkmJbg+wN3EkH1t
ob7cHyNBRWMqxVxDpDiuMNx4ZvCU0Dn91YQ2vL3/qdb5pOqibYpN+D4s5aGUM3bVpY42RxK+1QLN
KwDyTlZ4+tL722AdwfyOt/EwzwzPvPuLER5YmgOjm/JSFq+JjmuVegc0BVIN3F0/tLckBSe2BEZu
trIx2Y/QDXRwmut1CGd6tOAQHIhhOp/qbPQ+UPFBHltWkKKDrbDxzjka+c1Mc5dTeXdFeRGsnGaI
hER4bR+7EQwSbR0Wyd56tK8I5nF9ZIUS4KvjNNRL4+Q30w4Qv7shA+umsvYVxg/AJz/fto9RCsrp
8kVH0MLNUctJ167evPDKgWVX/3CjWz/7Tt++LaRYcwuMgZEY++pn/Lh5shc0nJK539JDJYv70NFU
3vsoynfrF+PGjX08Sjr05byuPyUtxiz3TWCMIKzU+YTPOKXJ7whGHWxKMozokYebEhUInGMM0JlI
EKssfqqm8wYlC1dOLhwNJ9Or7KNISn/GuKBonleKV+/urVlvMYWN8A2bj1RRMkA374c97f5Yei5C
+1KndOaOCHlOHwrmbMaWtkJxZS1D37cqkm27hkZZSpCvwz3hDUGFVsw93MngbX1PnC1tQRD962M9
5er1oUNdKukI1CSQpt/KpRLDrlI/UIC9xDfeiwCmpXZgblE6KTLiC4yVCwy/aDB5NaOSHO1dbPkx
v/BatzSMtUJRNluhwdEkTjpEFGMZ73fvRaYco95gzjl0X9QPNjZScpc+VhqvfK9MB+5ML9Yh8JIC
TbtaXS4ka28MggLDPGq+LgyZzk7LpSn45tPRt28tdwrmCkST81Lcm0jzPpwLxH/fjTBfzqhpEvAr
b64q5uZb/Kd4teYsrfhe26zLVzGJhgl9Ew7exldmGpWgBpZF1uSbbhrm0lqq1H9bsnf1RDWaF+BX
P70ys7TLOnDkNDfQGbjAMN6kapo4UJhjOl6UdDfY+ciH8Q+rYU/6/1oE9hIXXZVIDRRS3RyRNr2v
WLsD6foWkDWQZ/CK2M+UdTZptyds8lIWrsdQk1tVB0C9NL0IGMhQL7S69ofQhcgC8I92o4BQEJcb
Hw6TXlsvnTcUcJux4BB4xCLfwzb3DqG8T3eba0b8pr8xHy1nbMuxO07ZVLoganV1wvx6Be485aSM
Wxw2z+eBocCXPLEJCU/QC74eI9ulTa2u5wZcBCzvAQAGi0448NJsOoWuykMh0cBMfN/x//R63PqV
1mccWU4ZRIZ3jWwNFrwd7hj+Br+hICTqCIjhO0Pje7MHCRf52nskQ99QzxWtM+RQfpcVM6JAIDST
8WR904dYSjX79K5loUtOcqT+fr/BN/jpVjQv4ldTTYLFim3NvRbvI4/IaK3ggD7OYaKJ8LgkvrKA
+d4qFsh8fmFwlDuP8HHFcAYfnvbV40ifiYVabgHUfpumUANgM+GGN/klmS2HVYiF5Ws5qiRafK8i
ouflGPvcHrsT20R9fKCRxEC+QPYbF6qou1VUvpgjXDEs/6B2fhfBT0faMYfyOMD2Wy+CpZcoBgSA
TwJ7uXdYNKDb4pR0jXfJJszL4RY9dAgLBE5BtW8HlpuaoTMeM//6x8wO88+ROExgxpTRIgGNvGrg
WPnFsoVcnH0fyk/kNC4oTKWNlf+eMGrS+Ih4m3agZhljU1z1/BHv5784YF0tq4/ew306yaqmubhC
AGObSN1Xc/LXnVtsqTcRwehK/2gH79vR6laLjLIwyCrR+x7zaBXnOZiAgT/k8CBiS+OLeM6cbluH
D1QE1UFGmPbd3C2QggSMf7Z2JQr0WAmlWi7MS3yzouJmy3sLDbd6aGBNpVafEUFxn6K4UPmS4rx1
gkqsqEih9Mv0Acwm+CCMJasVoiB7LUvqSuQm07uEscuSji5jtSiF2zI1UcECycsKXvEcEeAIOwoq
LuA3fvlxsUx6jbm1iJjgZOcLWP+//iYj9Y8oBxm2PGZWM78ns5iRoa2MEx3KSEr9id2u+00O292x
c72Vq9AYd7Qp2oG+K2SLftG9uyedVggjoC73B94wpl2Z13yEYgnGOQpMpQkNzLvT9zgBkJnWB1SU
S8y1rUlEj1Xwv/0RBJVl0++gpTY2A0qV+IllTEY5/9M0dBEgGioAnK6AM7VEiO7Ej5LsOrLLQLoV
l2QuJinZHImfGpH/RIEvgQkI/do5XIeStwUPajAzOdrnOq7kWaJ0CQU5a/p9ckh/iqxFBY/FDejI
LuIWnHc/tB2AwkZnlRiN7cKdT+u4S5/kLbOM0MlNN/hYvTIvY37YVxIJnKHYHiNkPtwI7YvMjC4M
uLRnOFezg8//xf6UWYwSsbuncaYUN3I0JtXzGQoX38ayd9QT13Af3A3hp2oXW55HlVPMmarZmF36
+GKC05dfur6HyJTPrkht1xGYEXFWgjnGMvTpEPY0oSVpHzoUzkPpiEyEQ9biC8wMbV0bakS3MY/H
d+xAXXfM6P6SagIlflfnAkTNXaNsxq5ZC2IJSJx5o0qFi7PunfGAY7cLGzpk6mhehJFxrpJDlbXj
M6tBUM6nuWYwmJgF93/A/pdYeZBdOLqa7D66hqhhpILTQf4LWNirWxU3/2i6xpxayeoT9ZsQY5//
5AOnK68V2ZiXhRkpemvItR6+feOvlR1Xd8l7DvJz5Q6WrlCRI04u4q6NlhYXTwp8W3YeYMOXNLeW
ktc8o1qSKMG1LyR/aKMOBuvm4ZcM8oMWIDS6qeknoKIwg5/zlHMhk3x0mFfehpMReVmRuS30tfqb
d/wD5cc9sUdOcm5e4tR+JJ2+rI8A7ISZwD5XvlznhNjH97e/O4+nOowtBkrmovf4beklDm73eZzA
H2q2+PBZYd9wFNf/wB5eEclgLLfusXBkxYbkXB2N4kPrv9RNHoJs8vl8aSM/LdLt5AzfvJ7FCWb1
mv8ieqFvFCnzKX+cJHXtUsoreOMbljHYxwyowyYEO7oBPf5spR2g3yUXNa97rNDQJI9lSqyHlZI5
Rn+uyOOGDjB4rsIhzzy0i9QDMfbTszpPUx1PGtVbcJL3MlWmJmakCgt/GwytdKIGlD+jtBgxCvzz
eoAGeOnaZZb8b4TxdrBgpGRZ4+5K/tBAOUvb3SXWlGTurfC59Hp+z5lYwJ78+n+xwQToRKMdiB8W
j4R3A9jY1eSBkp9w3Cr8iMv6NV1DYAVgIlGGDVdVngKLS5Laj058xvMKA1waSwTlzrL5cDxRaz6i
2baxubJwL8U6/Q7vf/lpgU8U/frh5+LopTr4+IYzuZctrgnbdztUXjEZUOvaZINXlqQaiST69ZWv
kIXztfyXHHxowy8pwiXRv8I/acx8LZqn1+gYg2cjaxqWfa31CbdiuCuBrM8//JjWpuVip4UDoSHX
f2JpavCoh3NVDx63FydLI1JnzV6LdB3SgusQ/1LoOI7L16hAG8CJlI1pvRDQPIp9Oh5Nxs00Ax+8
womrOalIwKk9zx3fZNj90DjXTwNX04mi2L9QOivG+7zEe8QUV9gMpAiReO3KADS1Hqe1XwUWXPXy
qZwh3mAtQ4ggP+vltQq2oKefcA5k/N/+uRyBetrttQqTXZbuTo9w1CGwpySnCPMjVCAD19+Tpzhc
0CJgwO625NUEewT2livhWx4i81r+o0bplxvwjkO7Ld5QRNXygLVr4LEje6b64H4npGtB49KToq6Z
54WCpFhPijIztpGPVN3o1O3DdCBrCoMwdQKE+i1wl21r94NTKuKi2kIdkeu4f8912bNWSyFDFd8n
t0zbRW8AnnAFL/ipAXdVUWMs5SHZHSWUzIMpg/kUHLaMVfAgugmYNJ5GS1PIaIkSbk/tdp0fcgyW
laaxq7kPNr5xeOOcjHDb7tFI1hByNGbRb1vX/n5mYW+Xb431qbDVRq8DkjXL1XEL/JTxXMuopDFP
8t6ESJ1Os6Gg3AUktdlg8e6a+xXj1GqTq/6qOU4BuY3loIYvyBIhdQlf9+21Qou0PAAvc1tGLj7b
r4p8WKFJWdAktV4sxuyJRoYYqVLlUYsIMEm4IoPT2Dze7IXfI6Stm5zqakpjgL9bo0LJxy/VoBBp
Hp/NiebPPyp9Lrh4Tyj+c7xUvfOstynsAl3mfFYqMPIPubZ5XIvgSZWcwJNJQ6F6AdA9QloWyjjJ
/vKBV344AXXEVsT5as0VsdWadpSAea4dtM2iy6wL2qhbzZGQm0pqpiThQ8iN9Z4V4lQIHL1KV6BR
ZzYLUfCKHBsK4MzFnn6hHMRf9LGammqGY8hSRUwzdZ2D6HlkK7q3Q/4FkVXH1aQHvRcuZR8ZUzwg
7e7SaR3j2q18oNblVr5zL4+Ogb1IWabxHOMiH/HFK89xS7Ga8tVnbAEnKCOz+U1LubCCDangr6WV
a1CVxklnvJ2gDE7vh6tOS5vCxXWySjSQdCFpRJNilxlnBVJyruKhHGmCkcw0nc1quybvSP1PjmDO
URoJC0MF/UC+PPXiaAlbtHveNXRZQZ7AtokZJfY4gHR3ozzWEFSbdDzuoVYQdcN9wSbiVMDzGYxF
pyCnubIAu85rGarc82BIsqq8y44Y0RHxwfSjZmeYcs0w0mWy2PxV1IFrvpthBNhTvlSIVnI0B47T
M3j2XCA7c5PtQph7Xey6Cjbygrnx2NpJ9k8NVYExYxjfUYSUAuK7a1tQVaLxb4dI1sWly31rnN6x
V1psU0rE1JQRMv1KbjuNa8svjq+Si0QKiTHO9tnwxPUAoTdEJy/YrR9Dn38mF9t3m37z7RiEiZZr
kppDoqH0RBiizuQ4igQdQDf1mm5+i2v91ceq1h4QAVLjDSWBmlvGpqPSVB+BZCxYnhM3yZtRxiT2
r1k9GwOuxwy5ReiU2EbuXedpLmIadRXwGQ9rpslJ3GxPTuaeV4ja8Cuh2vV0eif3mF6IeeD6S6Dn
HWEny4cpRcvOtiNc5irNeFtcfdtdftdV88RWvlh0rCJb9xkzFLjzhPJE23oKIkobhY2nfmUVRM9f
2LwBG7e9RAuOSqKdVd+ErsIGghAuJZh8sFkwHklL13FpHVds1cVZIE8wo5tH/bjpHDrhSoQn+B7X
lpVdEWaxyfV8t0kKmV5z/tljO9oeD9SR23VAJ9tXNhAUQ9G0KDeWhGqjQ2Fg1vi95LfTI5sp6otv
58oDkIC6ThhMZIaJZNXViwqaX256O+sr4Gebf+G1a3bL7I2sRVLAZNxJ27UKb+XsPPmVbaLNcOwB
DpK6GEtds09/OnPqLPHdpHCjFLQwsY1jTDmQlmsvmkXvXeHL997zH3Fus4L+KDzqtUP8iG4qTjgf
dy8qtJs34wQK73vp750VSKr1spfaVM8JJv/xLZ0DJYwMDPsAQDuwLCYT4guclrMvv8w/noLa2BKp
ldaEWJm28Y4L6nxHx1mlrQtDHuQWKtr9Qw8SXVrRX/QHDfn0tZcG8OMtTOumeZQ3LpKO1p65758Z
S6MdXjJECvhb7OyZ7ZP8kfN9zcftFiIowdXDRlBQtMzuEPhFJPdoxt+wJlyuVTUELSPTtDquzx/r
/V362Xq6p4ofCvVpZmWALTFGYhiDvmtjIHwNA06Hs6wI2owD/bmhknobkCXoz0iKtCjHw/AnlWqu
yxXl+skKH/82Nq/h5cvX5dgO6zV2pjjHra3mFiU6t9tV7wYLCpE7Wn3sp0mNxDXw44QLbL+S61aC
Dkf4eSoOw71WwptYg3AqgxxJwKRZXl3UZPmu75OICmSfL6JU9OUt9oxWZTlFsJbcBehX0smlRgO7
bGgvW+LTBcLPPdit4PIOqZVc0QdmwqbZQoYZu26EiPUTkeEajXCKZ3akHwFMO1bzyPQE6F4+XMPO
B9XoWNb3U5ushrbDixAUGlo40+R+RFU5LGiC+foMuDadW8bS8e//EafCaoQVw/c6am1eAehimPiZ
mURqWeMVPxQ89ZEoMBS5QTLpoUnGTJjiWkj4/QvG8h20uaYyJO8Wm6hwkGEKaZot2Mxp/U25vCdC
Pni7EIt3sOKs1MO3ODbeIN5Kmr1ROiNOZC+lk6cAobViXR/ZRJi35rYwoHQhXwFeJo5+5rwaW5bz
MUGr9aL2XAqFV9omWXl1jmRorpN/HN+A6hZUtvMRt7WiBIbD37PcSju9JJOGxathKDjvWUd25uBo
DjlNtEmT7QEB/KdJJ7vpRFtn4STtu4muF4IDvRgrX6ogO7qNsPock3GPdN76Yuh+ssIcz/OOCPPt
Yhhpnl1nUZnpw3fXSSid8K183f8p4zY7gduNBZJCYvvFItUF6J3EXekMmx3xoHTmHLFgXnu44pLf
vpAGDWHY3SuzB5SpjaBx5Uu41KoGQXji5PKI6G0F/JYxDItXx4YBTVCAL7kY3j4xrIAWGmixei9g
TqScKa5NhhWAAJc7WGFVUgJHfcQDH0o7v3kozPYDN3u9GUdjgoUYYdE1SsXPBRk34FUzBr5KvLI3
Tikr4kXcHNpmAKscRz0Sjc4JSxkW/1J79puCsfEjicE3atGPTsimi4O8rFysxbNX40yukFSl7L92
Pl06ytgRZ41mszegWZBTmPdPBNT3vV1+3yfNv7GDeo1Fav2t8qQ5zU+Qtkf7yCcOGpv1HhhTdHX8
jCmBIG2JVUnREvjr6kv98EQq0hDie748ZXhWMY6T/Y4HWyl7qlYB51qh2y3oH7gSfOU2GXZsibO2
KDAKlpE5KorN4xSOGg3DAOd5mYRGxW6KnE6xm0+IBEAVGt96fMoM8dj7xCSzP6/hIZAk5Dpec5pm
dL3p6h6/QdZBb/Fjef9+tfRaaieEecR9lgR5vGsYq/4WM+Etxr1zEsvAIzBgbXrL8KAKLT4SSfBK
rxeDq4O8i5HKGoVVIDkU5r8V1G3OdHUHzps7mpqSoy61JLxhbOpluID29fkSdt40UENBmJgLAAi8
6v5I7585O4wy8X5Jqrutdefa+R0Vpq6r3BOZ4DlaBjwdiKRoKM+aQlQh52EipYyYFErGVRtTiOpp
2xjl1nAQf3LrhJVt7d/Y/TEz60penC6zkGIZlz/xSBrg+dlW2ygF8DsaLCap/wxnBN7T40qci/nx
r0CHTh9X5ltF/pDPpCgSu63OnSSPrqeHo7xp0CarrrkeKhwhb0ErRqiHsl5Qx7MafO7Qmn6lbqFy
JBZU6JNwJ3WYhkHPY2/vDVdxpTwNnwSP8RiL1mpcLhx9j9s/4kbuYjVbE04p0JcoXZmO/mwPMvga
NrSJJ7EVavW0T7VN9c7MW4cWzGNk2I/8jzqgYRLjxl/UNrjB+vPBwjbNJnZhbW1oQeJlYTY60WBQ
4lS/EnU5pdX2Y2o4dn8YHWNLCK4p1ZnC0ec4acDw8iRb+kUJQ9EYKUQ9OuHseqFyc/FndJW1L+JD
7KuvTaP14CI7Vtg4Ek/K7eNEJWzeL4b2aCVfBmLvGHWx+vN9t2G56EEseDVuJYxrOg+74q8zggYr
vSjiz9VPp6X37DHyEI/AHsOb7DUhq5BwCQEAqtzZROsBzeNuZn0Lquxl3R175xn8IGWL6dKPnn9P
IUu+sRvGR374BZsDT+PMsX6PnPrxQnrSijx4fw8nW5Tg4W9xqG7FaC+MF/FSUFrvq1CfkTvCi9pT
W2KX4kZSXrre3Xt56tQUC+HjLipv/SHNCL4UQ9TPF5laFKtAoFTwW3rgmsZ/W7S3Eyi5OTy+FcQ6
USYczMtyuffFVlWx6zzgtJt6AIr6UJdVy4VK3Wn/E7iNBv6WftFfj2pGI6SOuCVGtaWBZu4MJ/qB
f3lEIzJsO//Xl3tZrPUe2tXTubHJH22kGnUnIkDWqmdk2ow8wK7cmtwQLXQ8f8EJQG90D614zUFB
3N04zEUyl156aXiq5eH4s9H6dINXoXYx0e8KefDEScCROxd6igXpCVCnT/a5jgQwoRoJ4BfTxTbS
BRvRTlzkdfEY4vGgYprf1ly3CH+pLmOrpvamiucrJFnTTInHifkV5m2/bwk8I8BAD/pdjCB/5Nyy
Q0MZvhweWebMN31Yr7sE9H2eN3m0kT0N9NSFEDxuRBqodX2aTnKFX+4FFXaCROHXCpk4CL/EohrW
8X37/1/Ooh/uxKAAS/GPgRne8BlmmwyMsk6Kl/UQnmsFX2+6WoWoZePovon7lXlpuDiuKhtRo9Ma
7iPOrF2W823b1/2f3KseaEKGpVLci1preqXv9kPqQWrCSoUld1diI5IY2nTnD15/GcmLEQ5CFp8o
kvutz4P73ZBGoAJjO05Ehirme58pqCRWUrHy7126T72SNQbNfVz2XFmLtcR5I39ftnlTbEgHGX9u
qN3QjBbBfKcdXdgKIjCW+5IaOPchR4RVThkkpvW69+inoWl64Fy6vXDlo9HhTVj7S7d4FI13FQ70
71xgTjrycxd/9PTb79XNLK5mXWi3EcIzDCcweNF0Dq8GwhSB1xHq14xSCawtUrKZRyUXRSjZteLN
FEZ/5ovQS2xg5RDmpc9fUU7vTiZMl07VvvZmidn6azSFL6hSZXnjD6nphdsXWOGWG8lpI4D0vjWG
amFwlL5glcc66VrHqlq07ft5b6lxQ+DzaaA0awRhtnr6+efWuzqffVnYUyLrjCccxv9xa6zi5vOx
65/Uy786GJC4pAo2rj9fPJRyF4YrV0lb3iAbzUUi94ISd9U5bAPpnSk/kfpzZ8HHcuHvybEv0iWc
ILb0jtulMJbFZhMowd5N2FggCQV6A3j2sYWhZZ0NpbxE54Z1az9Inc91Tuk3yT1NbgShrqb+Cwcs
moOJhoVpMmipYMU794PJUOKCbbTXEqRjj1DeUaaEbO3k2cvbeJztWzyrlMzvxsGp6Ux+ppbNi0hq
l1L6fOJbpK9vmKJAENtO403oRvYeEQnJbdMygIYx4WDoBRFSWkDKKoJOLe7QZCdmvZVmIfaO7Htl
7x/L/25T4Ld8najLlivMaqbkUkt4ttodN0Wgw4+9DTxkyS2i/l+wytQg7sHjbTLsTE17CHcEcgbO
8wYhUQnA4LNT3Is3aUzC1cHGvW80zkifXj+J4MvFWyNiXvdmxiVUFfeoH9kqp01rFnNbeaCRYY5G
GD77e9V4F/Un35OUBO/xVSDCoexAEKNWtTkpGPByd6oR3GO+u7YqsDSA66T+WBvwtA7YwU5EE8Ml
2Kne565RUBIzba5F4ytH3NF1X5+FcHuqEHwKBFM71xTC0KjiG8CwHjraUGd9CURlpbu3lydF5d8w
i7yQI04R9SaTqLUbCa4XP7IJG+FIfJpBhoOqI4Oca1d1dRTXPHt8wbdN6Kxw970tv1D3lzzjVYrH
U+cR3iKaWH0zuRC2v+ikyzCaSI/5HAeibGpoZCEmGZ8tlG1q3askTaqn02A2PLrQIPCG2MYBKe8P
w0bgEqsHLSExsaLe7lJf2ivBhKgsbdeqsba7adu21N0S5wCXzlwkNolBQN/WDgszE/czf8CDU1gn
scC0XqtnhyfqxqrstMdf5BAga+l2yp2N0WtVx4WNTQJ32jNlHkLL/gMNLJ5nSSI8tb1Bt+uxccyY
1CEwAUdiI+90RRGjz7HmRtmD1XY+JuDGf+rA/+lTD3kA4cWI0PYZRl1YX1wZ4Qi3Q7o0b08q0PFz
BdNWPuGYSTr22YarQFssn9WKqFTZT88V7YzUCmlygJkYHkZ0MSeBvu50LXxmTnXLVRIgzADHUznH
0N3kq7GtBe7azeoAJVgBP7dK7m7xeRoar+R3qwdWleDC5wnwzJy9Aj12PB5r98UBHKvr+7BBV9YY
NMJjfRt15688MDc62TRhoMXJC1ISpdm+bnEk9YaRU8CNJq9AQKxdZHG9DoFCWdd4fS5Xbb4IrZgd
OFU61WCv2WImDv+wKGVvO4EARyqeROWOEZVrVKP+0O056nqUtPq64ZBCoNxJkmeJbQ15vwGEXXDI
bAwFtLUM3n6jDyUcXWCx545Ihzr2FYXmQk3S+Qd1xfoBSIviyVvrn/mEXflwFkKhhLlRKpGSBWgQ
KaFE3k59U+5XXj/PouC29fsqnjEWrgZxQeuDvffcHXBL3oLRPx0z8hzms/3ZVVMdVlZK7O8A3UYg
pB3RcBthm3gsY4qWNUspmhFVFBPnjNkQnKP63tyGRXtcAx5U2Lkt3Qg94A/Jwg13Sq3cDjuQ1grG
M3tBazfTB+Xak+qPUasSMBIYBiLUMeu3YiXs8qTDXJFwLBgxn/NC0qGmsTPO5aUEG81KIP/JQPD5
qoezpR039MY+h5cmBKvb6r+a3HtdWXwollX0esYKWBIBtmiY1kAVQHkqXsIUrMDEZBkuaLARSs5Q
dq593KhYG/TCUzFp/4QOEo/58+JClJqLOmLSq0IdyD9eTGZuvSAMiyD+ENl+/TiZNTcXng5c8PaI
FQ9tRJ8ufnAnkK0WYTEF5ZdHtdMWOaWkP8kyKeYEhrvSv1EgnPI+wRbtSkOVi3G4Y5ejP4kiTtRb
dwzxThKX8IpH2cBbn2vGGQJ3aPFx7GK2UzRQ+pNisSptaro92Q78fOlGDxXor/U/D1rAfMEpzCB7
sdiP1hhNMkQjQKL70bjat/73879wd0b/AK3hQRR/g1QDwTNeaI3rTl2NoL9D7CavWEdsgONCWpiy
HBEi/WXl9HdmO05YDYBbflO6j8Be6Jvg3VpSl9s+BWdMes8SxRdh+9OeVowJbm1lH7xWJ9imuX2d
WqKOVewqS1vMrmNznVrbr5Ks+q4/BRrVI5lbW4CqSzcKLhkYTH2WoJFY4lqi7VVVAVZdO0QE+O6H
ESBOtaxX8VjHdVRpKFy81ydfktdbvkNcRFnZuak3r1FYwSe4i3BwO0xpjLKXP4VWS7MEk8x1rijA
s6qwz6MLuQY6SrJJDaSycLMqz6+r/alqTMHBRRzufPWN/YxEtrrOK/2SK1Z6Bqq5HQ4nw2ZZ6t51
/PLivipN7BFwV7MxBH0JfGVYhwWp30hp3SIE1mRTuS6ya6xzKgXpaqHVyub44q6GtgZI0bGGdzQC
qN40jUzMA8zxgZ0xopVsSejxhUNCyfkc4cz5DjCACVFHqFRHcdQMwqNtTYDUIbR6cFvDBMa1bdf6
mO7JIvV4HPnOwlaW2PIkNWijmZSeav28uN7U0mcuSfsg2GpJAL+6glfx9hDddv5Vt+kYUEWQsuDV
mBZWKKUFHp6nWK3dBoMPPD9sCUo6Mu+wL5pk/Ox7RHXQqSEDFJbYY/gVk3LVB4YxD4xaVOckEmgI
OQSQ95nth2ej5XyKXHpvlz1Ej8Hb2zRug6TUrun7hhjK5afygmbeM4HXSLeOOckabdqIStUD0DK+
2/BbOOBAbk8wSbq46KafgTnFv6f6V7tmkGVwa1uptgR2HJ6OgDrubScmKvvVG9IGykWYb3WNhfME
3i34YL1AWxVWik53DOK95Cr3c4M2awEr3LBYARfByBa242EM/U7I5NdeWpVgD8mLPPt/mE7GdaKY
uSgc6VkmWNliX8OBpH9SK1TzTkQSGR24PjQpWrO6xouOl88XieC6dCmic65uAQqeaLAWh8KRAqj6
diI+Px4NfaOuePuCMP4rO9OW5nZvrg7TSo8rDQhMKGooAt0zwFvFUe8esecebx6qA6Ce1Ygz6fDP
U/T2W283FzoQylJw2xzxFJfHUm70HmNbKnXhF/lSP/LLc9iCs1oFryEFm9BGS8O5Sio1nEEueMGq
fgIZPuq/R+Mk9eEKiMBt0BKEeP0vAi/02InErT0LPa2cxKJ/YKxd+sYDZoHYLHZD8qrkspzBcmLu
D228qub1X3G/HngQKF7IEOB4oq3MP/q98jIcAjQIOeLVSSIbOtBDR80TZ4yoi4tHOsRs9nC8wL9p
Fp6oix9xd96YKMQECLrZ0mzyYt1yUBHrSs9H0/nYNaJRMMZlbMl/kHp0aBz40VWDdudrUMtzDv3e
Z4K5Yg9j9D1pZktXXmFfjOw/hHsTCIndPlT78PJHfk+MyXDeJydX/NKS5UthgnDdn0sZgh3q9R4b
iMh1AJ7bruKUepCiRE/z5BbXIxirXoJuRlsZGZCoLzDgYfEOgXhkFOcuOT+DehvIjh0BhsHjH8Ix
y0MsjYWIOBDrpYw2iwsEuUeHpvhKFTY/+5LC0q8d8dYzVYrlbYnPdZMCwhm94S+JplI1kM54PHzj
pFgsmRh8KJKBu8GlMuRXux9931sTiEa1MtAbNxWiNruPX5ciUIMvIU1qvb/XITZQ8RXCF8c6yrHT
/j+6cXFZVJhDxsmcG0zWQwf3qRvS3A8gE4F7fKcNPjmpgheGtof+lPYdb9KLGcmH4sq3/+s4DBsL
TcUOg1NwLtfr+iBKrN3/LFXCK2iNJ93iCsT+RWG0ohkFilLOEiYu7Cf0LHO2VzYBlNK0omKX9ytD
xNWNJhbdFaHX5RpdktDyQJQssfaMsIwqBHyi0E3OAwkMsBOP+07+5K8P6tudEyVZC7genoPHKXqg
OkbYkZ/0I3Z1RfuervrbIuAJrfBIDIJzJo+wxnSEu24pdsl+DeuJH6iJMptskyRcPCpAxdvmgU75
lznPBnuOFLSLTL3gkdzOfZeDIMSpBt7SmwbL//mju38c2w8owtfr+qNwpMeMchF4IYwhZH0NAbky
JFMGIDtIywtJ3OOS52z8eQuUpm9I/5YAVvdFoQ6gtt55GVDulOk26r1NU2ra1t/in/8RtRTmW5FC
DAO/Gr9aBlolHDatqr3Z6kb+Qogyb48PF7I3bWZ1Rmi1/a4w7JziFCkF8AXcx7ahIlfhO2HJUXTy
V/eSErdU15Ts2WWOXJedOVT2DtF/iM4N5LRSmuNBjlr1leOcMHz66BTNktH+JO1mnpUkdKJa74fq
XNBIJlk+Vq76R+t3AtGm5Z0NbS3NUoRGJ49r3WRkdqf2FsMWir4kDZgU9H2a1lLdCLn/GQiRrCYF
syfCekHoe1+dlNJB+91docxxzwSK+oQnu0FGznWSdxvtHCiXELoa4lL4JsOv3OI2aGSVLkv4O34p
qhUo0mD8T2spZ6BGXzAUN7wGendywy+QM+E2w+0XWUh7GPaRWMoHvhRjuzvUoy/5lDVyKyQCaGH1
Jc0FK3TsiCgDKTcTS9C0mAb6Nz/ge8GeNbIl0vTPfVbRo88SNdw3SKlNZqEK377Zpu+znR+CxPH5
Re4xEcRSOy9RP/kRD5vfaHDkkH7hG6PU0vntBCNjGn78J69H/8Sg/cjLxwA05vappBsBSzzq2FF7
p002JGSto33hVb3WOQe79s9ESLXVVk99zVcPuWpUgutqTQT1qoYFPoVYZk4tXySXskfTC/rFjdrQ
SwFpmOT+UZqoXi4HuB4Qc9wEO9NS134w9zfFFoIWs0VMlCErrhZMtInk7NUjg3siaXam32Qv8tcP
KhoHPIPlzvmgmiAkY7SSB2KeRXJ/JtWTZ9hlNazXNqC6uBbhCcpU3bltiad5BUo4ng9Y7Z2bY2e/
qKYijEPIlGpNiQaVrb6KsVNR4P87z6c1hgMEeTWwlG/0U8b+7HNaR/ZHvq1rweUV+ncbTWaN5mSh
gCnfGBoRgE720XSDbKY585LqaKnQP9dqANQ70d9fPRJsPW4x/nhnB+MSYvDUx774SHf0fHTiOMXr
zZvz4LgyxQmaJ+0xLsmbEEy9CoO4vG+Aw9hW6iceZkCdsAJwHI566Gp8kU3MKPh+uaboz+oijYMv
wdLG9Y0xEGc+rWqI2XwM2Zx7uUvN1bvpoDeQA1vddxuh4VbHM/6J9GVCl+R1ZNZtewO0U/D+6dgq
NKqJFxYktrHSM+d81BeSp9riRDy7+YCaUGQN5+zNqWj+s1fX6JMbxzS8SGrOQGt/mnRAfw5ts6EX
yRoPI6Cucjj+MBow3Bhs74eWZIg8MTHHEe/SeCNjtIrnqQa0zE6B6Xz5bR7xF+3NEIWmEtBEos2r
XeVHNlzj8y0V6SHXcEVbOC554SQCyhw1kcgNcSZ2YM5iYcvpIYwN4kxUltLrDI1ECXOQWW/BorNA
p/ngq8c65oNFwv/bTPurgoCHI5X23+7z6xvh57V9xaP//4WjuMFhhS1LSx//6n1JeKeqskpTkB7/
yBTyDFIXYB7IFiLXiuHOElhpgJyZaYRvLzuZCGXrd4q0cvHbph3XKoeQbe6MN95rQdfM4T4iVXwh
l/E0rons8P9B+p4wjH7pS5mW6y2bwUFJrfKS5sUJsKT7e+t3AFd6uuYzfjsGu7st6X6VgVNJJWo6
MC7rswS6ORs2mBxzEF/Xf+E1JTbHHyY7f8MA8+iK/O+oUNYIGh95E8XTmA81trtRBX3QgZLiqsaN
ktyG7pZ7qREmdoFu+uIFYops1O00PdkXDPDA0AqPvwrZ+utR7NJy6CKb7DhjRMlEMBM9VxTgyLiP
ivifJ1WBWMBOCuHroP4M6y3br+gpl+WOoZQ70IHAlRrkNViGKU1gzwdv4eGgtdVlaZGaBlLmZU1C
8veTG/XUCkxKV5RRP1PnbunfgEiZRR4AbGBJApmjbKk0YUPUa8LTi2AUNtoLw4grNKZJ0r/8kFB3
qzFOgZB3ZfP8RJrNVMdcAM4xqkWWOGpemL/L7uzOhlx5tjLD85KP1HwEAOSxDF02VO1I5G4Ybbld
tKy+F9bOTAivSrHy1jtmaZbxhYbHd7uNkNshN+/qS9perCsd7eXgEB6pg3008uAnICmus2NvjZ5n
0NiD2bbJKP6hkUQyBxbH5U+UaN435vCWfSC4y7UFx37/sMB3QQ93yjv+XuksdOM/5BAMag+l7xrR
IBIrM3eg0PeIy3vxgBqXAI9JXwyYBuxNixlF6BBmRRduINJYc21oLTODQpIZinOhZHk1Tk9n6z/W
m2ej9rLKFI2h97kFUjdbAi5gMElFsJhCBmc5xa7gtwSVgty3Tk4VcYVhtNCKPSHvWHLI4ECKdP+c
5Yf2c0Nth+LnAb/i2U5Ls2IWN1Agidt6tO96LHdxhm90Ez3uUcg/aUalTEeTKujS1LFe6FCkvfCM
IsSOtohgG3LE/Qk64SXpYippPOE8BSo+9YLR90bizgeVqsNi9cMO3/fLKPuQVzaR2RcwvZBN7maO
6Wfzy2mRAh9GA/ImN0/lGL8aWPjmkjPZRF2W/hxFuSXGzRVFutSouQ0qv5CCCLcEeHnAwIBJNZen
B4NDOVCV7niScwaXBiYHaCQhPmT5K8QpwBkH6i+ROgNzXFuibpHePmCsqy05OS1FS8E6F4S7+rqa
F2tFMPM/ulYwBqjiIKuO4KbMCxL2fYYMYkC8UupPEE4GOv7UAsUXtshVny9cIatQJ1b1lKK7qTdr
jQ4zZNkxCFsnPdc5gNT48Mw/A20OPgEmrYs0ivqslR9vb7NGp+RDdh6FWInWTq3HzJ0/4wBTmBCB
a+Ua+nBFnm1j2VgSo0XQIcNiqm54e0V9QWSD4Pol7W7c/GeeV9XHxrG9iIXS6Cniz0HmiqPT5xvo
sHGi4LBQNvYyWsqvBovs/ngiPW/EO9WkZugtheolYe45S6zvr74YLTDiSoIAXokY0AwEc9nrk6rs
LG3/EO/2IliEBAiclSUQFFeqmv2cTQRbl+XjSlfrzRN1mkmKod7x8PXvjgf62kXmhTVJXxvA7WS6
fcxZZf3ekckhk7LvzYB0nv9JatnyrJ/YMZKxLhS60v1CJXsAFtt9QrMXQU1pRjSTddUpatgFbamj
kVtr4rOSMsGBi2u+krR4J8sKvnMVVhmgo6a3lM94SyGTgndeXbWVfT8JeIlJZzx0A1tzf+DuldHl
y61YXw6Kl3lnB/0mxyrE76J66d332SWBqwworrXPMXg223Yy0p2tLvcpZI2cR6eb1oOjTe87sBRs
BeHOCaHxNFkFJ95rhXcSjsZ9Ou4dtZOsfxOTwOSyC3cjjuS7/stTcSL21HMtv+DgL1vcLrhBN0Hq
4l+Gz1lhBCQHoBEB6fwjujD7AX6lq6GxIoNKOgsQ/ik2ZDd2XuT48uGPlgA8tLFFAb9AnugnW4tC
WX1oOptFeva9GWzit3Mm2FUB9E/y2ie1yhZRI4rVxpbTYtDMMHo06vJk9hy5VPCzu/ImJjQ942rK
kImflhi35WCR98Z9ooDfq/V+mAj9IM3N7U+rf++8xmiZTtkRzLup4VQnZmjGHhuPHkawiTvvcxJv
OH93hmY4F7hMHZmmgyINauV7ZpiWks2cwMFYQXaqrKhxSnzZIm4iXl7dSh+vpV1QwnxNRW+nG6cL
KdB60YVELBQWy/0Kmqy9+jbuFL9biLT8hfsaDuJAIIP2DkqYRXfvxKXviDz9kFP1rHfuWO8Zezya
7tQfapspFlaVdaSTpYyBQ5CTAzyYmDiC1N5Sl0bTnYqEDLvrLgW/i8tYAUMAQ1GYeIwstRHV4kY7
Bynzmp7RICaiOh6+up4fg6ImkWTexW3xEQB1fSRSXrF4xH3ida29lYf26RfXjok+XJaqwJWQzAUR
7ffS1gnUWNGi7HiqlH8jlBGBLhwXKDRUtAUhiGBcZkfvpazEfQBZwS2qu4TeCznvq7YpG0I2dCEs
smhURbG3ajABd/O+w5ZNww4jA3+py1OSLA4qZiDCqSBIYqYpMT7RYPTLEVKReLU7SHHAJikEc6lE
zCLwStVI5TrHIWNHftG1WNTsxY/1AJvqrEdeNx83G6drOVYXDDY1bnk4kB1k8kWD5txBFEaDOHfM
IHqztrnrhNFER5Jsl8mG0eBGCnEA5GrSHXMzcDJQ8yhXpq54Z3Ip0PmSCcEEqgBiENq7mPo5hgG/
WvCoKQSEy6OuWYjkokVOZ6EwvjSusYp7vnmyx2o2OCfjAlsfuxSiXQ0FwcMir2SprYk90SGWZwTn
nht1Z2AAdD34tDzAjztO0HSqn8w080Ce3DxxwfX1G/X0Ab6ZT3QbzZzYIydrjOVVmkDWc06DlqUb
8PHwgh1MAWEOaliBBwqoALoGGdyawPRP89qrP9sU5DjZcsGgxSApVSn9Xp/Sp+P2C2TxvnTPfnYk
cvm6JxLrqJ/29BnHbLmM8mbwDZ0Zj2rcnUxuZANmUTYjwwYkcK4CBPN8FtmILnYYRsWGiora68Kr
AJ3ln1+Zevc8pnNAswrNEhJ94Ax+ymlkzMXVRUmsx7SW3FclkgX/nE8aNC+/09cKC5AtGFoavurw
EO2yVGbCPWmqfy4qPPLM99KZQ38NcGQEvoGTle6qhkzeasRLBXGZDrCuBAzxOFVcf2KaX747PWV0
/QhVFoQ8+wmHqRKRonNBP7wnd0i38TYoEkSGEPoxXl3rFFxBuJH6xVt9wlmYnzY+37hIJOMBuT7w
eBvOVulK8322ijqfJPXH2JhMkQKRiHhrE5WuEUn5V6RuvtS6gzLhlXZArc7CjmS8pqu9Hs2eBzPQ
sbBHJB6ZI1V35FQf5YZOJwfXELTXmmI/JKsyvz4SDjJ9iqWnVXc4aTBvMhAe422duQnXJGcg5Jx4
E+9ZKrbCzXwNHpiDaq6ZVSPAMrc85F8UabSaBoXPU1v39b0NGvQ0sMNGSeVlP1OJ/FXHea9uxRQY
1mqVc5jvEf2oXq34M7xX+Qsk3oyLLiMKcvMGRbsluWihWak+oMrnuHejsNtLbgO74VVaCbWhueTP
h/4f4SlOSOceqkcGekUN4GZRQubWxWxEpZ3TP8cMCYAJOYxj1vwQLmcNVGzHyDq4TT15FvCkAPHe
lKw5Uq7INSxdOsbh5GawuX2/pqU5p5/tu+ixUxxucgiCObJisDDc36JI+cusczpZ/MCmMBYZMOIR
oQCE7UYq3nN9PrB4HSLa0krvzFks4JmAcpE45wmBcZ+rFUaJw/w8pOzA6qClzZmlGcfarv26RnLe
nvVAkcm9TUZ8dsFiXCHfemZxKT3lchL5VMRrOUATAbBx45LQEKUQxnb1at7BCLIVxFF/BQVJjfQZ
l1FGWLA5XpJBkYsnbb+yTK9zC5fwJ0MKLek3yOf44R5ZCK/SCqaIR2eOb541qM/mscfG9cny1b/q
dIEYW44xkSO1VZKf/8uM3UxIihXqw5SzgWwu20pu+TEHEMfsDiCSJTlkZYChO/FLyOQU1NPRvHQg
VznuR/Ib2MI0+HTL32erQmV+eUqkIYiQxCUIDJEUy3a1nP6pM9WZrC/XKJ5K7JyOJzqsFl7DLhGz
69Z4eciD5/+ZW2bxg3GDTa8tccNE61oamrukF2xaGEivTciCV0LXRwJ1m0zSO3eQiBVKJPLVEMKL
fyxYZguRKYtyhRPxRNE82Qjgd+tmOJFnZdWmFwJSriAsL3WtdYt7uVLHtR5X853/LlMHWLlJFPTm
O1e99BJoZTK4kLL3n7jME/NbQnOVnA3/iNMD57pm3ZNs7hb4Wz/cc6rZMe+9wLc/jbk8RYFaTFpz
MrqIgfCpbWkQhSvM/JI5zS+3UXEBS3gCJufnjk1MMtSmLwwVPQsrhX4pXcEQaoISdp0QAXf06H/E
xrUc6Y0ypFjm3KAMNOpTUWrm+a0D4pG2BeSTp7q1W+cwOsXQFuXkyF2eD90hHXlRtTfr2BJVjwPm
S19ajFvBrVmCcNEsgoppvpTAOxmVadjYth8xl1FRa6vZvj1l0mX+ocafNz4BGTqNWnHUlI22bMl1
qbILGfXhvJfupYJTYsDCS5y4Vbh/96vNK7FFwkd4ziPeQQIsSuoSbKRPT97663rgnmt2pBv8p8ns
1mVlLXxhdjXqaDpAWbgshNf2nEWNPcUftWI09VFgGJth1l0BvcrGZW09lWtDbNQRM4PpXA6Lp7YT
e1elNoMrG0eSE/x+Lhc4kKPhOWzLC0utL09j4xCbMB0U/mMVpLTHN1UeIvWfjeL889h+J65bO92O
46Z1h88EehazJzUeT0h9/qlonRR5hzBiqU7OrF8UIzE5/himFzx4ti5rkVP7l455ziQrl83+dH8l
TWpZSJWFE801aAhkdhhC5XU/uNUfrmLtZLOoOj8N+oDEXj6BXHc9gYpBLYYeGkGerLq81asLnd4h
5cn/3ap7PGGDbc+92sLBeo2/Zk4jkdZn50CSgvJ5P7HpVa4svR3d5TJZaeoAUbk1SjYuKTyFVRqd
tPlw4cfzT5+ef4GjhC0D5HwuDi8besOZ1XLiwsH6Gz5uxLRcFF+udKa0MB0UoScZa2cHqgPFke6b
lOtgK504LjWRskJ2yeUlU8ngVk2W9FmozNlxQndd4IUZBtDrKQUgrNzAjiHWTzCO6uLQBPzLA0uY
F4X1UEFmYAPeWi8o8SjET7wauxlNxnKaIXHDlsrYK/0Lq6X95sCkMSN2wZoJ4n/sJ7lFepNsk7Ay
EBgMthgadKZIFWw262mjcFXErvAhkW+R8x2dnrT2c/+MuP3tLkpd6Xdt+USrDVNQrhLEsDSJ0aKU
Izv9wo36FGT2q0EwJzWtKUe+a8HezZNl9ECGdE7Ua39FJ2MxGiDlh9uxFvMzmR9tELOQI41Uu5NX
nRaPieSrKixzR/iY37OELPpLvFLIJBK5LHCYCTZmUWVYvGvMmaqUnVfD8vLrZL87FxQcQgawjaRX
22ZS+C0p+SnudifBUJHDlN8X6AeKPWgQgFwDoWB/A1z9NcKjCa1X5HBnmUN+IiOWenu1RUY9YV2q
BlRFK7jHYsC6UD5Z9IIOOjoYaxIHOcOHswMo/GK2qX8uPbNqKraQEz9T4EwPdtznq6slM3LkSqo0
Zov64nMa15GW+HVIpX8khOwCcOSUQyVFV7vFoTEde5p4BiS5HQ/0lgSl1ZIUdWs1WJVfu8rHZZQY
V/EjjuJ4NmPmJEyqyyHMnaH1HUGWEbUdcYmSPiGfcwGCSwnDQ8CJ4KqYhDVTJ7+AtJif0JK4hKd5
k0M9W/hz57RGpVU06FgZ6MOpmxHAOKKNX8uSQmjOxnuiUZGhilqmXTcqVIdRQ0Ew2i2MZ5670GDy
iwrn6dlSokCBMBG564cNEp/fXVuVjlMbDLeb/1wK9SAQGNHvGJD4dXPmkE2438Q+EK6QDkdtvL5P
dlVMHqTaHPeXKmgja9jVheRUyH04T18VkjQEFqjqutYnEUIC2AjT06ravtX0XJNa/fymwzj2EMwE
t67/bhQMN3wc8tM97hReEnfkQf4qnCVIMf3x8XtvOmqPS3NsL1b9ZhYbDsVDIL8dqtK/x5kyW1pa
s3xsoRj05iqWsiZX98ltfWB98SjDe6RSujBYphPyBiOfoOrCrNyVaXuYBzU0R4FcqJdFhzkM/XPn
zUK2q4HVvjrglEB9la61WpnoTYckRT5zyiR5hBjggtGqwJeLtpuOc7O2rnzIMXW5uEoNm7RZLRjp
BDY+CJpsKbmefyaJSkwm+1qPwAJur0+MaFztJSCrQZKDdevW/cgedzqHGP+KiZ0bQZL2DJojfwNm
NR5hBlGB6wsOA25vsVzVKNRQPfrgyc0sefw0YvgoMAXBQhvVuZVMRhCNyqg91SDB69CjSwrXafoE
dSNQ85P8b0s23CkMa7+cYQetQ9eWxRuyX9a/Mkl++OD/beuI9djwIH8MNG0KThq69uf1EQttjx4A
m9cnZw8BH8kBLc8HtO9se4hKkIpoj49DcCDdQkv7fijRB3lL9kBt+TP1lHzAtGL+5uwqScyOuIRi
DF4BSocdL3MNq9+RGjHxxE/O1fMvoKDgQb8hah1smPkLvcVXZlV3Azh6B/GaSs1fkyiiU2Mh4Rn1
QLUR5MrGfk3aL7HAuWN3yXUuMo5QS5SiKSeAFqGU/2ZVy1L4qJle+gchckIgl0rYUep2Uv5H2CRR
Wvo8r/cxmsnuVEH5fQXeAmzWesZqIJHfVFlBOuh4nFPvDGkanEjGyNmpTDeQEajy38EUQvngoq6k
YnXkjgkjnFrJ1t7ekALBLT3gBE0bqbcpaeQURV8FkTtjlMUmJwQgCsPv8PG6ZlVBYxCE+memoZI+
yhSME4xtkDUjsxnktpH2Z6evYQR+qJ3hcp2zcVZgFTVlFeDpdHDe/uF9LIei5ObhrJnDyhTjOPQl
ueX2mEFuRZHV7z41tLijLNGjZB0nQV0p7TJdWok2e10rLOmQBiKpl4qcEjwLRiHigywLc80+zz6r
erok0qeU23a4jI2ViadoR6pkqzCY3ruOyESGcBR4y1UWQOdqL0I8vKtKSHJ7OisJSXMNdbDR9OJs
0YHr3DHSphXYp5ALIjDSeCVWzSM2fT0diG4mnEa65jUXO/UmiY5U5BL02lko9/VywDkL6BaHu4gb
W5NTlcX8MJST6t9MrE3H2OSQ7a+3dkf/gTrmbjRA48evFDvEtgSjtC8+hWJ15SOtxIEuSvC1+xI0
s/ny43vMwybtWBIu1Oo8SmjvvwojEf4D/Uv8ZmIJMEIHaBCPdek0mXG9LWbN9KQqYzgrg3h8XjOS
MzizD4zmSwGRItzoGLv8pOG+leDiBDSTEPofLZO2WTqmPBdKnWZgy2X/aIrGIfoHCd9NofJDXCZ5
kLj33LXfQu9PIBpzFfIzu4989i8Iik1EZ7/dTrMUS+4wZj+U1orVokp0gbWnspNa10aMzxpcqBfS
X7c08vGX5w5hkk4DqOT7fBZf2FIcX6dIPp94il/UXl1gwQxurS/QqV2+GxYwpAiTghVeli323xcQ
tOmcNg9mgiZ5HyJGWnx3RsIkAZuALCaTcPdhP9M7Uzkpmd9Pwb8OvKQIzgx2xxCSLPmXmIo0l4Vb
qQVFPS8jT7VU7IIQVLg21kqPrpgkJjxgLq8hWLQn6+p5fifpPJDn61mQW+v/9A+Xtx9eysvhuf4W
u+YbYl3INOLaar5f5Dts9VnQry0/UKuXZBduOxz5mpAdVGwoOFtqw2IiIS7+IT6lKZDjbJgdJyJ8
DeCkAekeNHmONsBgasR/4+2a6CxZk+PPFac8djRUnU725ig8j/y/nM3comPT749n7f+h298QcSdC
fH8AGeP4TPJkkvPdGueTA3mYkD6ogm8vpHNfSn33/iObS4ZHV4ax1R9YAS8kXeZU8/zKK3PgGg0x
92hDUT0PTsHjgf7HDRKRF+9BzgnTQTC4idtjsyr84eDg1SisXfhRj3gZceSqoitWhGACnoS0gOUq
iYnEVRJC/KNaufiDAyKoMTufK3WDS8wHaLPK7gqJLHHfae0BQ3ZxRD40KuLEOBkFlAPrDaFlmBjZ
ZZcGEDR9jMEy3TmKyiILfZCqUegDYI8DBs7WTkRkkn0J1KZx6Oqu4iLEDuPNnT96g/8XNOwEJpDx
B4rhQFfWqXj8IB6MkhDrdk27qMfd6r5tFyrDEawmOa07lx0dDDG/NbPFJc+CvB0gYkVP+zw/9o78
iKYiihEw0Vu4Vairxor7RsjrDRoNW72/4u8bns4AsAYRCTP4uCBrLufVDpBUeNp7Mko1fECo6+2N
g1wmX8itdZXBgt9mBlp0xn8QYtSCOZxC+5Ve4c4kvD6Ab32z6dqTNl6Tuh6dBNe2Sq/7VNvHEA2L
kr6hjr1ChqkeLFtG7+EYFJCamh52xc5L3C4cMsx0SwWk7+bU+r6muR6OYXpHJCRKeVgFUDERgtBW
5A+Am7pW3LmtnLWU1wid16jIKp39NXE6gzQ8zKUDqCjctfe91dgnmY386lNuttTptwssr9kuZedU
XihYDtYtsKrThpe/IOn6L4uaJReKPED7sxtB/7a2pEK8htqoahvxHKeu8imznyFCskpFjKG5uouG
RtZu/DWxAGzQM3CD3pK+WaH9E5Df1rBS8azkNTXNVfv2FhziHRK3MkzaljzXcC09CkazpL8z/hBg
5w4Judcy/BGeJa3ZibjGUc1XgJGojxmN6AEAiCIHJ6Z9G52X+Cy6+dyotME90DKHLMTl+CCPHKwu
vxpoMzTvdeKcwh1KXrzoOkT3MejTmBCJeGVKtLd1uUBeOSGRgyuqnUkmCJNRjyWDeDPkIbNrnYKo
jFQj3rp7d6/665ghgl6/CqKS8wUYox7m97pVwC1SHipwT/wV7KdfqytCjCsl/VaQhRtn14I7PFYT
E5+e3r9E3J2n6oDcPm5Ef0gEBNh/vbU4mlvAYA261hOiLCx/xUUtI+f6xsV5kxlN74AeuRtOZpga
Uv+B7c45w1E0exQAQIlNn5YptgHBhgmR2RJpIaeVLaOIOpIUASrpil9nqodVMKN3Pv1/AyECNvGS
E/vtyh1EX/ACXMVJamCl+KJIh434BGJYoBjpoQJYaYUOTEKQl5l0PEA3ufKuA1jdZ94jEf/zym9J
ZGMvBt9EC4hVkqOVNOKGb40y9Tm55muVnub9zgLNtiQ/g+FDolSgOyhmEJc/A2NzYvQFEEOicQGD
Ia9UnCePxZ7lNQBNR/y5BiXKSl6CaGY5xxS3sbnjCHflu+Idc5iQHWEOAs8oY/KqCZ+OILKUB7hC
9rIKVG32DbGN1OyF6kPAU52662arJaQFiuaeRn0Q8L4ufijnLGusRH8+UK/uPremTH7Mfb2SRLf0
qdGuUKZtznJF5UCG2ysTAMyG2m2cay3jztonZLqw11v+/+pAyM2NtUgAK0mVoKKzHy2b/4gkZDay
TVgsYzpeh0q9d5r0z0sRi7G1Jigifn7Onwwebn7vz2SSDJJrQY82RIwhpEHwTcl9791IHAWpHjLA
14WlyhbkB3qbZYcfFxHw+InzTPlzWSEdcmkV0mKe1ZanT0qTQc/+hwBNdi+3+DgWOGcnvRL0UyEN
OHw4kgeCqqA2Er8HuSrWZCTkzP3qTh45qRwr+qpACwX2zSZwd2aC7JtVEWqQV4/KW+UxotHZggPo
ghDF/lWg2FhJP172/wnPqhAH3OZs55LyKJOZywngUX61mZ/zsfhWnCTbNiGAYDYNUwPiqMnCH/m4
WGyWUCBSxFFLYAtTwkGLbZ3z1NayKUER0Ab7L1uMuOIlD80ffP62M9mzCC+8zDu0a+NnyvjFkJQd
qVGVzsUJa9KB+UZmx5jT1+zBggLD9g5q5nVUhEUCAvV0bG10VJ5u8Or8PbBjFJkP0NIIMFxyD4TS
zcffSOAkY9K+Ok9L0CFeTgwqafU2ZvxPbmybQDCs85DdStTarj7W27tGyf74m9f/v1ApRZkmR5+G
pSAPpaIDzeGxg/ofokP4yp2gXbvnb8PULNvDxkOGiTJrwFDi2Vbem+MGWMzbGXVFoYdrL72NLCVt
5uCPV63j2A9MfOBI3EE8Vme/oFqr6O37eQUYlKp4PWSDVK7pwwTGRrbX2rUqZ4qVnxBbRI8FYe3e
5YngTnFFPIgeP9aqoXYf507gpV2A9W3nuzkcqDmBnyqp/o8ZbaMVAOg/2WaudWcHzBJsFl2oX7tV
aNf5A/UTheKKfRNMlFO0XsWbro6ISO+YPGfBDO+lZNOzpb1gRO1cCe72PcpzTyxldYtlPhJr9zST
WARTnOJgzhcTJwJuV9XitWX2uQqIDXdjCxelphM9EN/tTo2/zqk+Bcze9bagcbDIvPuZhbalaDQq
FYoXCcB75GhNB/65W4HqMqS0Iki0fLtUnAYA+z+Z7cDd6hAz1I61GtCj+s6z1UUHBiZPMQNyAP1F
U0UM24VySfEQZMgd3YyRj4BS3I5gT5PScQnjacyZdsNQgYMo/Wx7iGgQHJj28AGbWWbhBQ04cEFf
QBwMeCleCf+/l+ssfysRG/qf7Jv41kH/Qd6QyuYEOyuDlHt3bD9CZhtJLhXnW/si7GiqNMqS9ne0
yvSAyiPkGCkYIseCcIBuqN3hsiUwO+oFhyFlbDWriiU+k1eqaokwmNEfm/NUovCCgVcX7sNc4IEc
/Ga3AU6SCZDn2cYcXhJOsrvFYezyebHpUz2txca1WpNia/rSac9h9NBFT6V4+kkAoOey3y67Igvo
6OzXdKzAXZGAlfaPQkfcfym9Iwg3BP/p8vpJG52+cjrAJ1v0QSmyawbSkHGLyg2c3qH3fCLByGBO
AZJaqLt026hZcoyTHwi1baUHgjykh1Q5XhPts21PyosiRXv2CcqXOrJZxFn29H4lwESVmr8IyG2K
eVQ85hLO9cP36B5uTfKrUT5njCX7Sa2MFlim6aJXhrK1EOgnuLdqskEqlz4gr2xlo2coJ7bprLzD
HTdUuwgRzoIw6sWrdJcTK6dFUiCLIBpKY76fevJE9mD66s2vfg8g6tyngneROxYHYtpcFQS+hhs6
rJcH6R/mv8fQg188eApvk7EWxn1ck+LyR6f0sba8+xyz1+TzTAsbmPBTxn4lWtYajpj4rH4JSPP3
J/zr0PVj7aW0Qyv87CZNbInjMkoIZ+gGKrMnKUsObZXve0+/UtCJGnti5QZXunTNVQqMQfa8P4Xn
V9TAYMRsXEX9HLLh8nezWh2dR1oyokeIbU1pDrTfsZexk9q4k4s+Mq6CQRxBEw0AGX7I0mUyUyYB
OAE3TgByBSSB1MLA5ZlNEogzKkC+iZEwGjL1w6bzAJjbmQjF0OkFKQrkLIIotYzG3G0I1qCJgqMI
Otc50ej3pvOLsltf0s67XDwCwFJJ/OeP17Ig4hMrNGH/kixAzcMBEUsyCwBVqbR11SpaYhmluaNa
yvAPM7BQex+Jk7cPbVLM5KYVzHtAn01SSjbMj32m1pUs1XTSVEJLAcFwbqhx9k9VWMW9zotuyRk3
xSeXXerB/72Vcln8ReHhXNPIzkQkmfdW/GCfTJiQHukdi+ApokxgaXOb7biUeeN5FnYO19LQdhiZ
JzcF5Bp3MiVSFSefanJCxDhBAn21+h1gY3ISTGNjDOjekkBxohY4zHbjTGA7vOKzaDQevaEKDfOx
VVsCfFnFFvxRk4SP6WuUCvOiSaVajYG+4+Cx5reP/vX6J42NqzGLczFdKI+ao/lVsa3kdZmbiiEB
g/nIvoIqipoAanOIP2jS9wWeL5puY01PQ93nnml72g2SOan7e7IvLOAiHnBIt0Q8TgAeVIqL+BbO
7zC0s+5d10nrW67IGPNvj1PF78Sdm3Go1kl2WjwYIi3YIX5eBDqx2Jw0HZzPUtMymdyr6TR1b440
hv3tzpHiRnWEQmbjFNzk3cDMfMc/iPGLSeo4shes2IjQvyu3qfyEL89yGbn5exjH2L14DPZzynW3
6HQZF/4p6eTkQgUDnCbPQ7WKKVfqJDFoa6L9us6A20yr4AbjPFt6m9VxIlN0FXkSK1Aj8+ZqMOW/
ojtj00q79NW4jBGLjCR0ILmvGYvD0I+Zb4caO3Q9mO7CSrVmdQftBzEksGwLeRSjI3nPveprgOX3
u8Lis2mTjBnFyozjnMc5kwVuKNR/ZOeNGYJL5mDjhUKCVqvSbBurd/Rr8JiTGX9ai+I9tBHPSo+I
ELl0WuOdDc1FCHXmFZ696rMX+k8DZvOqUB6qXSbiaObxwGN4X1GJauCMXpRLQtCECtLaVMVFRonf
vgTfaW4NHihYe4hnEIcK8qqpYEukxF8OawzL2EU2ymHOReuvy21UsIq1tS3Uv9JgFQO7IrXUgfZX
Z0S1nP2Ep6thallqiX1D5zbww22Na8/W+EOhY5q44dg3yOE5+KAnmFqOHA7SNikdHiwrvYlFTMnf
R4Eybc5x2C0+/gbziwOahc+71RvQEdhWj4CKY7uwHAzf3GzBk4ONH8irJQg7WkKFWidYND1NyNAX
DvPQl3p1Z3KFiLDNPG69/CfxaUYSsZSziMuxHAC7a6A5oRuQ0wzPR3kUYttUzlCcKekbMKd8Jpfg
/tXHC2jm0wy36EEhbk+U1ZuGqp80cdRK0BuoTkxsSW2+78uiVbFSf6iMwxn3dIa6IIFK4Gu2W9e0
k9uJAYQbV8wJ4m6/gpws0QQgvbCPw7nGD51jjJpjA82nnAs6HnETH7C8o+96a01RRFuHsJGxaxD7
XhTdGU+yODDVF9DsqAeuSMcpMBdsnfMP7ch0dlaLRBAQg1Wn31QMnHX0nRtruuStLwLW7OL+Jska
wKmAnYYSXFxqaDMwmFOIhPuTXCKDU0MsCyqSS7LgtQpD2MKAlDl4/xTdCLw/Jil24HnJavVcSjRN
YZfz6lqgHzU/33Qz+WEzOMmeakf9Dxa/uuXv1ibzwNnrRsCpY0oSjLo355fYmwn2pEP6FhPCUTid
2woqqhiOteMvChxAy+FSM5KjaZjiI75kPX1T8FQSo5u5dJOkngNncR1bmd8uG9guxuQ20D3F/8TU
c1fIbVAEUaJxCTfeS7Xps4LIIvoKnrV0VGoY3AqH74Wu5v4aCGy7hzR78bJ9msvhq9NAau7tnAK9
j3axIT1GeEQec++k+GTJMQGsYj0GCXywSVcwI2Sd0P0CWIz3yb0N1H5YOq4DHq7Fs9WlPGyojyZn
pvC3jc7CoilhuRRuAsDD4NA+LUyRaXxlIHC5OdRC54UDmQChGT6d8ChDSC5hYbP1/Vd/MDT0qysW
dunCWK34BvyQf4gBuAQmJlXQVo2g7pKViJB8yprn72gqLwUQ0HS5ZlbM127SyvLIVDcfNIKKZUj5
mpf2jw/Dc1KvyupzqyM24Glp/3UNnEoSCgi6+Xb4fbIV0yA2Zi39f6sbwQQJkDtK1cOps7x0iD8x
J75+N9eCXF2oFNlbyHDsISSBCpxl68rGHQ3EvipTnXmUtKZJewTygzU7gdQ4ZoJnUpNGBTOyHdal
NmbSufgUbFlwuvbgJyxxwyu3Ex6Zn7hU5OfRcNUiKnt/tmrTiLhHImWYk+UGNDPfKiRN2nif09wF
72lCLOQzyivgAkOTQETqpYrPrZeS0dIHqJpG783v4zUB+vFpcpm61YNPle5nuQ5cMJeNVCDidhHx
f6kbjNrUC8+d4ZXwUzihajrwipOkuMsBZdUugA5/gcZh7c4ILNHjiqXncBuhM4R/2aoKIAYfRf/e
QGb2K2woK1S03QyxCZqkYWcwnYViMbMAne4TsnYTEi1BRU1LDD8ttUD/BACRCnH1HzdNyQcSOGLc
LIn1GZJWDl2Y+OU0VCWg89lQRlJaQJIpIy8LMmNiuQ7dvsuSPSKw29v8+bzyPgAycBhdeS+WWRW0
i1he6eWrr73Wr1V9lss6KHJBfY00xhgZXGZ0yFPzUd/7VYGHS1aCK2nxP2tGdM4wx949HP+pfzk0
+Azfo/vKScA0CZJ7Tc/AEea4SqjUZIcYh0lVifTML+nOJUIKuPbnq4MzmuoilhsOt6dWc+2uOCHj
HaGofbKshVFYL5cG21JyI6XfwpySMC29QoPVPxxlC7SL8UL5dvrWqCB3mqtEWqHKgHz9y8K0UsmB
ZLaSNdg2WQzVx/KcA/KFyThxzv0f7zn70wckMTdJP8sa28atl9ShVpOZ495LGp+8rl5B1vAMSmjs
iWchIULVlfDoQSQot95roIZ4aFIqbc++C4vP1aUiNdD7w6v33x6PPzT6cn0cFxp6AcjuyGuZicf9
cKW/1tK7X9YdZYODj0o/A4/uXkfO+aA2pJw1pbGowPDI3UvG8w/ZelyhRkG5BLRRHTpjVOZbjiBb
fZBgMXH1PM1IC3JCIUiYi1wbTfW1aYTJJFgtR8BnLd+ijKtSDwDxF4IFeX0J+W/iUarkPSYMcxyU
Sv/a1NizWekGVlpbnhpFJXhAl2b0W3MBXemF6ksxgKVZeL+Z19TqjcSeNetmiCjQkaIldITycj3v
QluAh5jULhVBWfIGeQZ6y/dJvso2eHaq/wE5VLkjE+PotPpvzenM5/4OlkfAlMW1Quqp8xzn+R50
U3btpFV5zOuH5F+wAT/yeCndW7NzKNEqI1IHqRp+k9HwlZpIgypgPvP4KV2o25MDrHpvraWk4dXb
q6QHrriCHaagg6Py83PyHI56X6GjRLoQUnk7nXTUIVsPV374DYQGPDMCJ3+lChUzMcdPlNEgeegi
oXIGmFXj+xiJNIIw3BPLNCFENH1X5eBvv3Hit8ENT4Cs3gpSg7/5svYRrIe9X/GGMXsWdQ3hMh3v
1o90poFuQd6I74JanIQiBJZfa1mOcdnOSnZ8U6yvyKTCFIKaD/fhRLifvgOw713+vU/WLC9ZFesQ
0h1NHGXd0+disC903BxL3UYEBWYbd3y2icXWDTpi+mmsfFIrnLrLwOQ/kwas9FYIRWJ/dnFAkObu
pq7opKgiw5lxt1BvOePFuSPMkA9JjCPH2MLeLCcvhdWYnvXE5C0khRZBPYB5ES3dNR9umafgxTn4
rV9WFbjfKL3OhS0EJI1XPA6CvUG01Gxwxjz5hfhTRMPMuaU2+ObduUzPohUoSVRQqC8quaoio9NV
2oH2NUVVdwJLDFrPGWK8/M8XIncGOvuxCWpkeiD0TJfG1/9goOoy+99bt0BHN5JO4Q/a+8Vr3uTS
b2tfPCL/1DnuXg/tut4963SBfV9hLzgFj0T9dOB/RPgdjVdoUhBm1vora+Gub+8LSJROT7N9XD4C
WcvsNph4XEqBgt9mX/MHv4DlcL+oCiCEvIjRnakpGtxGkqQGYM9OAbW2dKCGbwE4krIbpJvokke9
S8kTCbmc0hn4Q2J2ErrTESByN/abf6JAz95Ur9tksE37zNmrJ4P/pzoTwGm7XHHafc0//19osPPc
BiI6ADj+DmQbNCsfbe6X4eV+gAOUXAx54jUTaEBYh7IezoOWQGK93dFa86eOKquWTBX/Lm1U46BW
iwqqXpZ8qBObYaYEWI7yatlA1EyqQATxcz5j4twiS+yM9GHhO5YCHAZwAcl1iCKph/hdYqjq3Zvc
/nHNdNGf6rT55onugar9K+tZEMnoikq4tSaymLEmE3Goimp2MXK9FZLXSZyO9eNialJ2TzSgVzdc
PXJRVHfzC+Sg8awS3x7C6HTbAp53zMth3mso04vkdLxR4OGtCSgpTP2yjSrTeoQsUtDm8pu+mCUX
ecAdvtMpDaXrHaMO9/dc0t1v6/A0wO3cjTxeBxVEIaCfdOq5ZR9nHpkNn8jQN0yQwJoZa8UahgXr
qQLYph9qSQ341EMD55BN0nLxnvmR+skLZyogYeLOw/xEEFSWaBngGq7WRV1AsAxDcU2CS8qhujwk
3dyKvFtlE268B4CUsl0S89AgqTTbWKlDx40FrhErzp2ffZXYKVNzZzF06JNKkqvgQ7lXKuLQydvv
8M/CNnryEs1lv7bTMuO8gzTzxS8saHI8lb2KGK81x0VB5kwbBZxSytk+DPrukX3FmsoMD4XzLVmR
EUJH1iMjbhQ+xtES1G8mJ0RmkQeoPhN3+UcN8Xgkec0EeJoYGtpHLGCBwY1f0Y6cISWcEEqmlll3
4S2scKAARfPQjC0KAyoQClbEtiG35S10nUgS6Lxq+l1QMTIg+y/uAnMpElgWe7NiRtIKmddcivkN
Aflf92VDiRwjYdOcSRAzrG9p3DUaAb7Vyfw2NHoc0h6tu75xfcro7rh98HFZmEhMyMeATs5Yr0/5
H5qVGqfQvM/fTdY84qdVrqSoWJzF+aU5BkBNENBSS4WG3U92jhxfCl0MEh5aJzeJZY7JVoV9ja/5
JbSCEWCJGeUvIDyfgR3WYaombOGu5tixSz3upCxbxuKGvi7rr9MAjkeKMQt7vhpnrMqFjlAshHxw
XgTe8CSm6VwKdut5wM0MnoqVK0lcpmQJzN1hV6o2hPsqhbmmWDzUF49SR/HfDsnM0Sc3ZE8tLjrE
vHPqzIieamqXE93zCcP7Iehlhve4w182oF3iarpNJvl/4qdx2tggkk2CRkrRCKDUmHPlZmXxgjFT
hWJx6/JbTlNzhGlGskpQnK4qUR7I6gdyGgArA5dTkx1AkxDtNTs6DvZVLi6aFGZ3KwSSjbudXd2Z
Vb7kxmuKr9Dfv6VL/iIF5u06LzEty//a8yaI/3FArnvO0lCHj6D7ozZK0ZgVXvPx7Q31gGWlgkOk
Ul0nLMLcnV4LsGo/8P0EwfjCpxIJa7d+u6OmNRYu3dMcIMq5kDdIzdekVYJlwjblygo+VWWGPjfa
ljvYqi8GmkTE7HSdl6QMT1hfsLwu6ZNwyJZcs5HNQXod7WVmWnBgi3X/zOY64do1gy3+5zFBezdv
K/4T420/rX8FQSJWxkrRyzekCS+G4/bsmEQDpEEJHOCcE5n2sCs6xd3moejXBe6WBcs0AmWrFc7I
zCQ8pfhgsVhgiQ9v9fKDbNNoaiXio8p3moJVP5kAqo9qEAMwuXJkEpShitiy5s2LYK9lEdDp+FeC
NA0cqcHADDJjJKdgb24LbhOix3UllIpQJnxFkAbjK026xiBRnVMKCby7g9/25jSyytfU9uTGABBN
rCXkKRtshOSHzTVvLUEIOyZeFFX67+W5Y512Ov6yPNH0HHgwK9EhTiZa8bVqJpTLAsv3Z2ZnyJ2k
JCmo6jQp/BbD/IFVhiwieI+N/mcu5D58NbkQy6YdvSyTafUs2e6oGdlbUSqPPoZilPxmgPl3RKbc
i7GU1e3+RJtxAB7K3+KuyuKHfZ6CMA6+fwmvc/36hgu9mRZ7W+X9tB3Y7Flw/64X7NT3dU6AeahP
xe/Gfcj/KiPZi9v/xmW6efhyE+sktokTVSGZM0/96jGnoAhp+q4SVyHIRwAqfqi4GG52gb0KqD9h
XAbdeF4MHPuFNgbAZ403LhF89kcH2YaNATEFCVhH5S7RBOQggV+EMojY6H4Is3omAInCFDG0dm1r
bX4dYdb6pDM9zIz2ljBN1FIW6FZfpChJywpg4nARJYhmUFlnF12bBOSLNuzrxhVm6eJT1eNngqdk
wryZYskBzGcFiWR3K84KFcQk6lSFdr2+vwnGLuMzWLedPr4YEYVszArQt0dbA7df/NKOvLILALBt
ezrgwe/mUuDYmZJEFZU3HAov3z7dUBCRqbONHHzjuX1rr0Be5Lp+g1sAvZ6tw2iLJfA82LzD806V
hNE1JNAldErt+n3x7O9B9+fQwf9UbNjbjMVkQl+ENhd+CowXfhzQtHbYn6EEDiGbqanaDbX49gMN
m2n8kBwZ5TcgRP95+cqxP+BpOQHXzzG4/POGkIcnrTfrAPNbSChyG0H6hccPYC2lNeZNVXU4HLEB
Djnul/dFuIKaacrh+Gb+QXVtoibtqsyf8xRY/VfA/5iWZsFzSeEN2eWHcitdPc3zDu9wnUShQFt/
Jgz6IG5fh0EOMx7tS0Dzqw9sbfx4G4+4jOzkzQ2VmzqQ9/r6vfDv2ZMWoS353yEz/YsYPLn6iTc1
ytbPZrNeMLLKJ5TqSg+cFE0k+5oHPR5GecSinx3e8jDOr7NGb7RjV1PevQTiIqVmqXgqWkY/qlg2
ZZ8AyPbeygschk/+dschrKiCGCunCmFXwXRwzucvoohO9Fgv3I2FpqCBXKZF20rezNty4tWFy3at
rO09mfvVRacQJZt8k+w1sdvZeG+KcMjvarwImgOj1mAGCC4ZTtywq4aEb/ta48OIQ8Xvkek4Nmrg
Bp1/+y21FtYPGqqhApXFkoiNiVEIeJGHREaEKaZid+LQCuhZtsnckkH0Wvc+3RU6s511z657GqKm
39h/d9hTekwMq5Kp9orzgW6ghMw2IDvEVIX2WyMmxpfG4reYeE9SApSx+UDfH7y1P2i4ujHoWD4Y
an97YCuF1r8j62fZkUnmJX6ZvpIMEjtVKNEBJVxA+rJeYUlzaiTzPR62FwRBoa1NfNAJsJoV/RMN
ejTMEwmUHm3705xI4BClqTwqyqjOc9bkZGnzaG2DD+UnvQUzbiC9l4DN91sCwSL3iZw70DyyJy3C
VefvXpmGFBbs2Y2wqM2IyV80JpZK1EWe5WN6GK6AF7o5s3D8QrdLvG0ptaG/WYoSBozeWu4Q6OIv
8MDkp0umzESsLAuLG5GbjCSJ7rfs6uUZ66a7lFxnzGJRizQSKw/EK/ba/9qMrJ/2nIeFmaePynPL
DiJppW/+vt3AIJlDdcJ/3dC4Q8CAaU/jKmhA5+fkvtneRwbhOR2jGJve+Wgpyn+CGTEXL7Zy/KbT
wHwvY/vvoJRyWm0vECTDBxKvTJFljMJc5aHR3DgKGlZxlqc2wPSwBdtJwuA/YRPeTbMye4AczaBO
0JR7wuDFSpulPML80oZGOKLqvgnVKdrNIyS8CZCNjtJNbbChal2Tzfqmga7AsR+SDRK0/YuPAm6Q
HeZpUXFZQYsWLRXVmtOri4QqaD46s7zcorVPUp9d/q0MAnOd5+YGLH1Ac5dsA+AysFJNeq4TD7Gk
5WxkltchP3WR+jLOznQHO+HzbeplxBHCd2nLPtW/dsxYArEEUkfzVknkqNlEoNeBNShPj1vMmMA1
OMPtuYaQBT/Mf5xtHBHgNgtHHa2k2FKawltMJt2gCsOdxJWQgex3Vwk0sUDz4zpX9FEuqjPXr0Q1
x2dO1U5lKqaVhqi7WzEb9n57g0F6VVgs4duEBQzjeHcAaaMAtuz5jMBs6l+Gdl4+kFbcYtr1RQf2
kO9kidAWIwnqoU9gdSO7EDqKAGmePU6ZPLYVIcfRdcefgCshlWbSNpzphknoLIJcGx9HW2xOJJfV
tpr0y/++7R1EN1xgzooIQp+juql162ufmj3nN/Jw1ot11dDgxkyuw3AQ+WQOg8wlD0DlTjJrbzgI
glj/yBQ0p/fzUvY9wKHq0QcCG8wwf/i5VF8znUJxeZ2XgoCrCPFSqMjBgir2BmqJmt2tf4EUbdBF
cVu40fvRIQ70ObApt/48BQY4wigMSV24YvRNYOBvUcIBUHvbcaeUeDUbx/7mHSjlzdBjj75FoGC2
feryflXVmCH3puDHGX8m/Ds7H4ae1RM3DsyceDjh+dac5zNGyMfiS6EYhecNkiJIDhWgRGFdRMOX
bWSVZn4EfJBjJzZUOxZRX1fqlhlC0KpObzkkf8cqJ6mulrAdiq24QpctL+qqTVCG82eK/MEbe5+n
JEHesPtVaiRhEmT3QUntpG7fvNmXrntm8q3Du6vkS/czzDg5aGn7FiOgiSkCCc0vheEJiczsA2O2
pXgZ5hRZwfVykcYLJJjQUmbnT1SwAFZj2qXB7/H8Fcg6jZTBiVij8UlAJv2PWlHvPl8HCSg8Xjyk
yUUYw45mm6NUbaarrWilvpBZQM+4t4X8+4SCnL/TBPCUKYArr3mCuPWZjRYqfdgryqz1o+fx+TLv
FFvBbPNYMahPjic2F5cewfal+5Crx1rJWBLuka3dbAkCE7gnV/qP23ZINTuGTxZjVeKMFBQK0uem
aOhaxP+SYWzZ9Sdfr46BQ7bVwc71yliEp0630OnSYX8kkHVQCAJV4oAShs0JCA3/MTQzYTj39o4/
JwbAMw97hPh1C2NQ83Axd2EsZBsaHGkszbhP2q9Fhh6aNQKsSRle/0m7OemGI9IgKV1X5dw8r8YH
OB9QfZVsXjTMKISObwwnyNkyLPhAtk2u0qmpFeicCrwcG3qHxqqkLGIBP+N20cKkzlJWzPzH8YrG
lC21cxVUef5OpR9I1Rr8f4dS+UK0pVxJaxnfnC+z0W1t9aqHRB67EiQqd54iv2a/kY+q+51D4LXn
7Y70yUWNN6EBLUVJcAuEj10w4182/Ee1IbaXAx2IuDPllnnGGKz92sQaAWvtrZEHSJqgubqHqa7y
j0LW2OKAQLA5xg1qb8BiKWGBOPUev5nlpk5esBoxawc1aB86tHcIAhTFQaEBRcL4tiLjioeraMzq
2jdtieEcj8exSKzJI5U+TiDMzpbv8FstHh2pFqBTMyqf8BcBZpcCVH80/s1xOEQ3paYYbcf6Z3ed
jCnSGhRSE6jIa0rv0x+zD5CH84ObEmwTbLpMnQeAhRYbRYWwcupPA4nTh00s5Y+LIlXjQhoQuubr
qDLNYOLtJ0Xputx6c1G8ohCIU1j9KH1999hDvclqM+OQa6QcEhpPqMQtyOfM0UoZXYTn8oVJevq7
IABzv+FwmepvdmkIxJE+MzJdXf+4EjVvSVTNwHbww/i3aeoI4T7xaoF3kzMTu4N7IkZimujp3YNz
DQScgpmgtFVetF8DQMb5J6F3ab/1tKEQpp683F9kvf4G/XkDkXv3SeCOpHM1gcyLAF3ML7GFnXyQ
eoDXGYLLZvSkOAHxh5Sdy4elo/ceRgCONmCCDATPHTsfP0J/dxMBStokLysyOG3jopgBWuPsXokA
Y3Rx4Koto+2umtCx8COg6sf/8yYxEyI5TrSRv5htGyZw/X9RvcNiYixqEbG8EfaXs3gBh9vHpsCf
MRaCj/W+2OTSlDInyxyYb5aUDeq/NV7jAVBc1TQ0Yo2KjjJBtmQnJZ6w0orXp0JsSqFd/LJZi1vw
ct4fydQSe/nOuSAMIFfaTlFJg6NlXgG2N0+UCi1el06S5Z1F9bQ6atGfBduvDa0JRXhZGg2oWflX
obfrHM+9/Ysnxh5cDRY7BaNzDBdxKS1JK+W8vvNmvBwzdVQRHFkXJIba/u8CSEpBy7quOqEW9wJ8
jpKI5anp4Sv5tMFNmU2xTTaZslS3b6UeEfKfv/XWe/qIVRDDSzdzDOIP2cNUKJGdfKFN/cNTPow5
y4kY/nYKvPIpXBC9YJuNP8gu1Sx5AhImtbfa/KAcBNHOsPMT5XAQ5w6wQ3BCkEl3CzVUNh48m22g
5P9l8wVjdNaMgyzsoJQJ9FCWZQrPNscb6BcaFVF5RcVXIFc3IPc86GD4iBFGGj4EW8FOdTzRYlzu
+VrrF1uV0L7c9JFaTNPK67WTuv2YSbuUxMUjcJhTV/MOjZZrV+hTIr4+dV/KPzIlN25/32yPC0b6
zGKFj2H0SehfwD+lTGohIgMl/xK47ou/CluRmN4TlE+QuIDcQMDlb5BpH5RTVrzSiKfHY2Pl3Zq/
7bxbuOViiZRpsCF7QQZ2PITGIq9rM23TjssnyXK/XS7LrPO+Q/vPRF97haiJ4gFmG5QXzjuQh2RM
YTLaGWlUVya2Q5vSha2Y/CX4QG/0buEc0XI+cMAXo/U3rFDL7ib87l8vtEd/UnIb4M/N+CM3onAS
YCJJabFVtm63JNJZ7f4j/kHMZyN7sx7t3kHik6LzUOf+E5FFPZFDQtb7yWrMrE/yR4RqIEz9TySa
8m1dM6d3AlmpouVVGRnNBIm5DCJVyzKoEZpn0Yp/bLwls9kVahueoQs+YqVCh4t2/2z43nCxOAqM
KDNnZveYunnBeZTBcFC69r1RRRRb5f9L2gBouyBTbechkbU7N0D3Nu0/L1QEH3Bv3w2v0qrQN34D
nL3ToWhMqoiPTp3ebw8+KEJHUOrjNhW0Bpu4tFXNrwQraUHpwhaE48ENNjd8tnxaEbO336yD7oBp
B3hdk2vUlS6wYqcHqenWwMwm8Eb6Oe7k03hNA/Om17Sexk6Dld+dgK2dP34bHt1Bok2IAMSeJtCP
+76M78ZHni48tds/zyVhhGjGIy7fnZ46rk+KdjNPvgvCViDiNjZD3coCdKKGalxBi2H6eL6p5By5
ogOJpbCwPRkY0L9kZ/Kh8HY6yKB+QVNY1EIUPdMNRwVQW8993cpZGt9kyv1k//x723Hz8N4rE3l9
UTkghAUKKjrLZkgGanNr7PSb7Y2tH/nmrnConBJ6FvYs2/IfOVVmPcDkeqPtHN0w/x0ZvlyZBwv7
oqg61PvbnG02jxi7L5O2MMvlZijtH2SVHnrgeaxseOB2jUr4HEanxGogGcam7WX96YhbbOXRoMcj
nbZ9aFRGOOBQV69g8NduMx38pjemWLSb5YnT/5JH/crN1BiO050M2Elg9kQE5SZWIvl9w7CsHUer
MsvoBJNkDzZpiJ5kkNAeO8llVg78qGnUSlE1Z1YT/5RLK7o9Z6P4sKpqKqnFSOA8TWmA+tTEieLN
xIfHmJLBlw5U7YKN1rs/IOrxiISVldL7J5l49tGDJuglOdJ91c3XSRZ390vZ7dhhMht+tH6bhh57
rg+k6HX5+rhcpeegbvIhUwzireVotjBt4UG51EIaehCWw+jBai1jK5xgD1a+CgqyPpK4FjOGDYGv
raMeKm/Z0JjwBgoG7nqJC/mKGJXaRfmJgD/LlCr8AACKKwZ6K0gynUKYEr4zopn9X1nuIT1uVvue
q3cOZ39u0mixNFXjSpcx6Y/xgPPnAoxXUkYCR2CMF/1lJq9r03Trl4TKSOaSYJOH1Sw8p8I1OGFH
9U0cPLKUmY21nup9IrGZwqCuJJa3ZVbH7rR62/cAVPiTXv+9bSc/XsHqAt1xkBKWCDev2nNr1Xoa
4YRji5Qe2V4NotpbU57l7iTeusROladVCSnQr+rP7TkvXtLwcA9UYN65+1ob9t1ZjH2KnPfTxf7Z
VdMxNmZgQ19/DQuC5Qb0E6DvCiGA8DWz+iDEsibUOJ8bqw8JAAnQ3DGU1nXwDERsrU/8ALEKE6B/
N+oQI/eUQrbr1Cik7ZVgJ8HCnFx/bSXE1i1MFnHQ+0m195iphrvqmvBWTd4c2zujgwkTf04x5ij2
5XBGyKR1qj2Ikkrh3V75WKKGxaARwSXYqTjByTptq2UfH44YNsXZp/rbf6FBrJdTO/5fjasCc9p8
M9DF1QO4ozn8GDleeVz0LYHsRD9vboUKYCrVmrNcrG4Zt3/DhIyN1da3xujJ8cQRpcOfiR+eCvA9
oxxOebdX4HXmiDttzr/q+zKFtWxOxD+K9yv3914gGLW5dfJgRzaZ3oiY02+U4+K8TMs5uQRokxcC
y7DG28nU9DFXUx/jYvIRSLfzkR0aI/IQFpg3PhsqyBxpCSf5gxJ0pvR+lfVxZMpFy/8PEOnBLd5/
U22d/fUvrZI1yi9RPDKq78hQlT5Zvx4VCULZrl/SQatyIGcoXU5P2wIcTj81ki6gm5EPxrJzXjTQ
BsTSw903jNEasb7pzYbngbSM9qfHKemPy4E4C+8EZgimmrr4ajDtf0t16glctYnkkjGXu3QcrNO4
ZnLZkBUUAvhNJO92Y6eXl0QWqZi8W7lgdBverencBXxst7mMsXQpEarzt5tHNg/3nt+a12FgnEip
U13RFKOqUlI6bruXIelkrotrjJg+76DqJ6ZakZzZDmryxxU7drvzJZKK9U5Zg/BpjY27QGzMDQDI
44hijkAowAY5HkjnCpixTwdW/Kju/2nRaIJieLOhmci/IiGA3XIeoGA5nlRDVh2XlmWatu10iK+e
AAdu/qgXnht1d3VEryzeWCl190BEZ9IsrInm7RbJ+q7h2VDaqOz67QMYZ6PXMrkgBgVJn56GXTsG
+WXamAfby3k1Iz3RCS3CIV+hxffBqhR4k7PZkh20dPaHoS72ert9dceNEre1q5CZZCWlkKvrAneD
9OMP6i3C9hAt/pY5cdYeqYUIv1OuYMTKg69FL04dtvDsAkdRY9+yesy75BGwddDnpwon2rk8J7+C
AUQ32y7bAJxY3snif+78Ju84BjRh9emjMPsLLR7x8wLVL5t18Dlj9JWL7uONV8qM+mLmdL4LPAFK
Qq+SHunqRvw+iISrwH6Shy+j9t1upUk6dUZ+F60R99soV1oa7ReHbu8rlMs3uFpUD9LbbgFejKga
yK3K4gCCkn43RRd1XmIwXl3+jIwYD+N+g3O5XtD2pHywHQ5ptQ2c4+EhkYgSr794pRG41K9LbYOh
O1VU9uJiXFs3RRwT3wbrIFbmgTtbWJ3z+usFWem5rBrahYfdXHaEEf5XWS16ntn+W4oUcx5WsmBG
tmVHAs5K/PgMe4QcTO+BZ+WJgtJP8iU7Mzeb12KHQRVe3EBjJoU3YRk6Mf1zY+tTU2g7nSfzKDIb
Ud6KHpDkN1EUUHEsKZ8AjEBuDq+Ie7HNKR9I0/3Ny/OnqSA5yW8jyxcD3o+TzGsZHuZ44Vtnl3Je
LngBw7Nc83a9ORnCtgc2uyv5rmmz6eow4AsgZ5d/mUMSUejWGGrqEkkMEBQT56PrOhPRaNxEwKHu
8n/DGA8s3MZWxL45tmqoj/EzyOxbm3JMpPCpRF53vity1yvxtKGXSQ43q5gVQd4x7KU83FymL2Dk
+TmJMB37WziY527Pa3+ZELdkkpXW2Dt3BSuhFwE4X3/ytV9FonVYqW0cdzH65EUP0LJOt5mk7cla
UYfOdw96nWUFkNKds2DxK0UoHENz/QkKbBfGyR955heA1B5xA/mRNajLUdliuzjRTUhNUQHJQ3U3
XAJWGBtrjltRaNCGOVtBHxwFvH2wNsPD3NK3io9NuaPfqn7I30zJEI7phHQ8XAUMf2/CXUbJ40tX
I2PfnixyWK6EB/eMu3BEoeCMA5thr/Bl/jMP16Tu1bOxN3EeZBltwZetn4uPju2/G1BZvBuZKt3W
WTVPLjuL0Ai9MYwGfoxxE4sXN4Ny/vICmZSZTq7zjO2GVTKx+2ApD2OwJJUuvqM+4nO3lyyNhpxx
soMRWaCjBCSlu7qRr2c7jtDSl2Q3BYkt+fYxqNXEAdT4FYa3oj04Gso3DlWYCOLZwfGudlcv4K9o
EQ6JH3mS8oYRQuCWNHFMSOH1NB6MlTt8qRoB5O4zUzZHeknGZFdh7YkrCjYldLvCULRL17n8btp0
cAJHyqYij24ni/9DtLL5TAj1K7G4MqqzBmGaago0LjIELw3VdiTRz3riMIC2uyQN041M0smCGr0h
KeU1vZF9gWGTc/vGaUfjVt1CoOACVosAL4X5KXoW1Fvdjw9dgGE3eLZqG0yul+akRnj/TK9+Ebb6
qSvG5mDaW3n+AE7fmu2/Cp/D09TuME66Bv0wsAYlmJkWSprpn9BF2udQtEKmorhdo4RbldJbCeLG
gE1kDlFHXqNjRI79bwvcNKvNx+usIalfEdXDJDCP9lj9jUTlbEz1oTB+vCzloYVM2UT9AcjL0TfY
1vtJ2TiEiYDFkjdD7kc0hlD5Xv+Ety5WUf6F1lxt0KPuKgri/gu30bRAcgp2xiiuw4goXpQl+wuS
19Xqc5V7kLpivsM2sGZhYRL6L/gbAADMq3LYj70xqW4Fjn6HuqOVnBbYZyWyVhr8YK0z+Lqh5IVb
Czh7NGMefgX9fMtGv/xjPoeotR0DECnD12vQ6yKh5jKEbic0Ikw2j6wtUTRiBfPznI5hihEJR+DW
5gs694Yh3K5nC0b9DzWVp29yMJSSlm1AxXMb9V+pbErD9eZMkUt0jSaU6Ov7CGVPn9gne+8nlxN0
foNPAMz5lzShEO/ZwmPGo2XDl+2uNd+2xbTDUjQVYGEWFMEmGq/4dPhMn5pKQUFWDJZkfL3uVQyc
iFjCTAL9ALNH8Kz/JdweK+rESy2FU6Myn/r/kWaRCJBucNKNfUY5QwSHCXqor82t9g2A26OgXkjs
68Ks2OueBcewjc4HONdwL9YNiF+l/WT461lWVqcxZ6+LWtMf5pcT2fwrNw50iPCqesIim2kNlvWT
2lMQBPX1sjdrI4uFpKsG/RRLWE2yxReR1/5JDF+kPcYifk62zIg/2/SI5NVgRTi+ohR3988GBnCW
eT6DpzMf/+kUEJFJwgRU0hzjNXV3/MteIr8ukjvBmxUOFkcr7vRYmMR6ydkZkPmx5XxNzKRQuOPc
P6OgOsq/ouyoV86Ke3+fS+Tp0mYbuU2JOu3sUib17e3zJc9pqiUGdUG3Jk6L9qckZqE3abLXGASs
jEBxFUQbNWg7ENTT9kWEsBP46IDIYc8g2a0ibGAUJbKxnFeycbabRFewNx/6myodbgj2ILQQp1Ln
9zk1vgFIjF84fCcvxhd9TP4XnOTUOrqTWxLRvqu3YCSMBCt06rZcIk9cUnWn7wBsxz3l4vNNSOrR
LK4/gXZPQFz2sbVCttfMorhr1YdcFVoySVjlwPNKk+0fHU3RpgRfyOOgnP/4YwWroTbhrSuO3NqQ
nG3IGRWQvJ0Jhkh8LXp3Af0WYudOYkSGhaYq/K2fhQNmnIiObsLtlYRex7/LkG3fUu5wjZrFaeRq
z47TisqJCkfaIlq5y2odWUld6BtsONVrCIqGKeUr5riw/QyQmGjGilyeAveXaeVEgclvbBWyqXlf
Ubz6/JgaWSo4QOkVcRZ6s2QUrKSR2Ct6kAFiEX0adA5Eo6+AkZgTQFTApFsaCLIboUJVwoCF6XUF
u4ctXSV4fsPNxOY/U5fsc7IM0QxKjxG+LqEhBOVgGcdLZ9spwulg9lpZAxXBOdYDs7qr9g+Y/Pb6
V6+aZ214l3hc8LqZj/QIgPyLAm0t24QvV8hpPh3Q0LQmacdX1B/7aPyMZUAhENph1IWIQpUB2bAS
ur7FhJwZB9WP9NFmm7BJxSotywsNFbpqi55jCoQgkRoHku8jsjdGXRP/m8DFC5JmkhyRKigSyhP0
3qmp3SN+UIzrrUadFwMmeRqk4O18MAXpxnZe42NsR92UoQF/S7cPMv1wkVlfhpyNkrir4lhdqnq5
b4TRHZvwHhJNbqy9pQ/cBRLBZVjfY5A+Y2rrh2GUVhM7dlNhrOudOJtvHnBs27Dq/FKge8Wsa/As
0flgaEuwDliIebPrPBmb4brd13HKrmYipQ8egMnOI08QuqrR8pIaP8hnhVdtKlshR8WMFAMAhyT8
g8lQWlDLgHDp11vYE2RTXVtxuhE0/vPljm2Gleab6Q8F8wpt0FTATFdZVVOruCOdIooHmR3LfhUZ
qlW/HsX5ODzV6kw4m6BzvV36HcBV+N9RvSrCpK6eGxtJT/H2PRItHvqvF+aF+wZrXo/2ByAFhWfl
sIC94RmH6eGTTVjrL6Kwcr3dTJE2CBJKg7QgflHgVZHXAA3g7h8sudBqctPBxwDtIAfyv6ko0Cei
wl0RRT/k2o9QpXuSmhRhyCPNT3/gLzzqGpXSpeZ2WYn+U2EnEslIIMhTVg23hsCUQDXD/+o6wFxa
F8YdUYGejOebxio5pMtQNkUGp1WEcRCV6ADC8C4F+hDqePW0Wid1skBcUd83+yHnSrCDhpqlirda
WqDeV9MZB3k3xEznt6oe7sgL9DTzK7iJ0t8mZ5P438LqL0u0UJOVbWh3Vgu/6GT4ndcOQuXaZTMa
aYjoWIsOJ6J56ff8G2VQY4a88sBKT3kdTT9A/gb2I1x73a851N0bVIPIGdOrLnqS9OSMV4pw/QAT
bQiEgO6jy60Gj8bPVLSWA8ZpyFy291CuK4XIhaSPJctFLNtxbE1miFiAgKbudJMb/avT1fslpUOM
gj2sLwapoNwyV5tPg1YOqhxzPK4m9U5m+nNQKPCGikZQTmL4vkE/OJznBe9a+FE0tkcaXWzAiQri
A0Gat0bfStQ8nkSpoD6ge5kavrg1wQwziO1ci3bbefAPB8Br2rA+MOkhvkb04Zbn/ewJx3GLlZXW
EDlZHDkjH8U4yz2Qb4dOyOakOj/1hLak/0AmRLYpHcz7F4DgGkoOPrzwtS/vvwQHnAEyvbOtpiQH
5y/WVT8AJuIUMlPHKqUvS88Bwqysr2fRMNKMIN3Pm05C5YyvPXjNwGbtKsfnEXNTM6Mrtm00NVJ8
nDQolEOuIPq1fsyeoWgs3IHS2e6eQ5CRY8uo+b0uHCbau07FU2tOk96g7+TZevyJO7DavPVPz2gl
qode/28aDTFurQvJhJMO3VfkuXAireve9O/nBJLeh7TV9Jz3A5cEm4GjqI+OOw+kvdQyG7XhRzE8
bzGwF96xSzfJYp8id9MYzBTRNCzsQfyZRzda8TJ0S/pyIcbgR2WPyyW7BaPpyxmMjnPdBAZssHk6
aA5dJrdRt2NcbFA/fHTNMoqHMW25hJZuUJH89aicwkQwW5tsBpxRix2tisge1uWucUEKFif39guj
HuDgrxfqZrd1+hguJM/NTfa2h/mIP7v2GOWGD2LPvSSxVadzBj/B3ksUpAfZ9I7cOVJstF3cnx76
fwpKrd1lpl2zmC04e6b5fSTsohctSDf/l1h3j2fm1XUySD4mVRuSwBq4lNU0KekqHQBb8XtGb4ZK
Tmkg2WNT6sPQS96/ogtEEGQo8oTUQAWvhnUc0x+FaCVACbykbQlHHaC1GjQzoC/q6M6aqBGeciD5
Uo/FsdTGLFe0K+nDt46EFIx0yHmrh0bd+dahSq6ycV5IzPbP56cM7O/E30lPZfZY3iWbYDgtyyg5
tjgrDq3oGT2sKWvkLsnKkSh7qpeMlsegvMxZwE1MG/dDhJbMpiC7Ie0M9seH+BqCyQpHo3YIDv4x
DLXDP/GrFm7Z8edcJfejUK4YhhAWpWEOXkNBpUqdMbtSuovx9Cwuz0B6ZTKKumQf/kQ+On9NLELJ
liMzYqwSpOljK0e+meiXDDsw9iGD5eQM0rFl2/qwvIaU1+Iyg17j15BlSLhkPAot4ByKBIzA6D1B
6C9+xAeP9zUx7juli5iLhOYddY0+UsHjXCM0Grqk6az3VYvE58aD41FA688Qo6stVWx4GnLVNuJp
aMf8aeQZ4CKJxGYYb28FQM+hCNrqM7xCTv9IMd/mCgl+S+yxM6o51dKEXO1D+KZdPDq5SwMygYkL
7X5SYWHtX4GpnLTPRizfzo5TSaQORFv+MkEWzzisZRLfpp9vc6JplqjxhmWNHLNrVvvtyBT810m3
boBCW+D4NwT/z5w0aieJiAEkBpXbdJ+nRapj9af2xRusl6L77HQ3SwP3GytvBvCltMsPdKliQKXK
ygEq8ZwI/SILzqUXwrAcTIXqdLCUHZZ0mkqFJVclgU9lvZwMAvDWlFs2YsXCemGBB1cRobH56WqL
j+nJd5zhVMaWIxK2V0up5iEmn8Unl/LqsWTXPRwu6UH+RIAZcHg/+tYdxztFjC+H/Q5F42YGzk7c
DtT9v9sIHsmH/USiMc3oYjoX0Hww+Kf6yBa8a4VnZl4GPZ9rPSB8GOfUptQDCbaHyFgT/gWrLrXB
sRrZIKD/H40Togs3JNITTwNQShLjZM7kvx6FEjnPuD9KbYB8CSKSiYVGv2YL7CWoCXqNn12zqcI6
VF+I3pcUHxFvXqLc4wqjlmssJzsQGd3CdKe4xfEySXoeQ9AA2+cRjCnNUtJCghLLrcUAoYMsE41Q
4Faac6+EyD2uPqsXwyXF5j38dmAk3e0K2/HJi+33U39Mk/pHhlmvSQf/qFnsMC9C+MTJPxmxjlk1
WAPwWDhJiel8dopGQ7Gs00HeJL2IJzO+BpnJFYpC0HHZvdWbsR8P0nwceI4UP7wbIDxPa+hYAM+2
8iwYq4cFxaDytxOzykY1WiBYPPXqmwfAknVD5ovp39Jl7uBOYEO74IeoObKjEK0m0/4x9QXHvWnp
miym0oB9ZeYLUoWCusCu15XpG3L8uhEsC4BN5Q+4EMpj8snvCTpTBtPMBKWLLZb+5hSaEEqKj9HF
Jkh74Jd1ds8JnWGZQYzPP4q9h5jtZO2EAttcikGzJW1vax/OcfcN/O52TXLNKwX72wIHqqFCRKEJ
JiKJhRQc+Dw9yFSksmENJRBqfKGJD10CIfckE6Hl6VqxIY4Tki+/rTsNfTHOqWPjwE79ouGVW0Wk
BKBiA8vKZ3vtaUcNEx19nK8G7joFF9bQE45+Gsg6MnZDQUFVTMdUN5DNKSpHF0gzJxJgNN6Fe1la
6DZLyo9yu/11Yohz1ZqTl+pVScUL3dx/iHoRljyL5BqrTckEbgLfp+EFHJh3DvPXjw1OjGNtRUAC
BXEqzjetnVAzqhhG2oglkM+1U786NLiM2/jL4jsmRfPKllKesttTu/4lIwKLmhHAWKoHTmny7dZf
PgK0oLuh567t1sRGVzZN5Iy4uMPpj+iSG2adZO++hcfE43GVO56PvkZ6GzubdevivSiDf3+Yff+g
nqigF2wxZV/2Z/G7QZmakgyN8p4j72cbAbcyXFWndM+LcjS0Q3Hc/QZk6PTlwWyJKxEqjuFNNS+W
UT0y5EQdZArGUvuk5jDIj+LLAYBlrPyURYzRxBrz8g/wl/sJqtJ21nqqojCuV6J/PWTu2s6nylHu
8yijAruWinesjpidSAh44ebidQH+6Aehhs2DAIyVrSbo0jJOwl9VttnfoiOYgHQ37AB3GXbPxbFj
JATSqNFOBhCqGNZWkfHA+n2QwWA4hm07vWfXRRR0BfXng0AfBP2Q2uJuwv3Ha/Ye2k5DE9u9D1yN
O1bxhhqf79tBTJunN48QigyCy9+orzgZCgf9Xgn9VHNheFaob5BTNbRgFBCBkhopGOIVTXeEh8zk
HGW6T4KNEL5XV/08n5mH043t7X42dTIzFbF9TC4vBnzeECnnN4S8DMb0Q6552QpXR7RQo494zCuG
q++XRAJD59ciS2OKJKqMwBsTTeRdCzpiO7hXVd/vsr2f5533Xv0E5ubZzNsYpavHOCzU9pWOJqmD
0RVXOMGHBxipQSpqAsG1kq++4T4EOoqohCmbu+9P7j3yEkJNeftv9wfgTe8D4ynfDI8fGCre65bK
xiPkJXJ5lA+Gq6GCcynZXdXQVoYURs8kI7LbzYU3tH+BYD3U2vzUyRdCFuZ/uYlTYAzvLoa+eqni
uxKbS7H8KZYb3qYWLsz518SfgJtWskUEkM5Kxh7rntpTKMXaXtiykdxxopM3uVGOgC4ssOG70hR7
Y60Rp4cmdHxInvY3qVERsuzaTs0gor1Nei000srLMUeSw4ztIzBVZ+MXY5mWDI0782xOqypm5bJO
PoqiUKcyrfgzkuJGolpTtkW89LHrvOs91soVrgJ2YzZM0ps1bQI0nCvC+Q0BTcrJ4+NffLG/h/S1
xkhxaZc/phOq4ysCAw8jcB8WHy6ofIINML7V6S3/q3bv17hmA1Xc8jemxVprMglGZzn8cjXEVGCZ
Y37i9zDQioxbmPoKOCxyOEddAPQOiNXilPNV55kPlRor1XUgeRNNk/dcJB1+zA24syLQnpHQAVUq
zHvy6GK971UVg89BMActMg2KqLt78F/ErYOubVG4d6WxWIj3UNg+QiL54B4giV8BEmWlxsoGRDyH
A5C3RiwsQm/fdssjFUVjSpsWc4r28Nc3LfrGY2QHUvj1tCdgM4VZySZZQD/r7l9lB1bXbnRIxiL/
j6llm9naFw8++m7D95Z3zyzXKOYaeINSzWCnVjeRgjymVEKCAdzCzbUCd8BsLaTKtTk5bHU6bIw8
42MfOODP5AuL8hamY0Pol6sHr50rAwsc+/WRDMZc394yFH+DxPSeJ8oVoaXeqZFw5TJLg1tqcX3j
aG91aFt8Pi9ur7kLd0ecb6BipNiBYTyOAn1fQakDeXZZwoGtWHRDC6NB2Ein5RXDrtJD0ZkAJwY+
i8TrY28yx9SKYZb9WPOXNpzDCGHuNP/cAZHIKS5lvWhunO8wrn2AwX4C2luwgznsmicDxor1bK9S
y4DWTVw7tOL+iik9vyAdlxrE0WX8q49ZiA0T3rsj29aTaG40f4MpS8ZAHcfAlvWSxiP5YKgIJd1j
FWdNIAwrAJ70CI/0dae6n23dHynnSJjHJSaVDnn24VQS3J4WfT61lEng+ujXnWWXv7N6GNjzs8rf
2FWmzGA3LOpdmGuQzQr84KFeextU2BHfLzo5l0VpC0caD98eQy7B8Ud9UUBrLrbfoZfD8rrbHXEb
uiyrqx24OxJMGn1IwZbIRItvtwFSImZ5YXQ8+/GPib5cYshZW9djUyjlZlBGG6cAAwm1qc9cVtYM
YUAr9j0LwICK/Kw8v9hNjDfoDJHIjEtIe1TprcxKPUwxgmctCbwDBp0ca8vlfvZddi08IG4hcae0
f3oL0Ppuw5VNZ2xGdiA6bpYLrHddnfoFdxN6vPXGgbiFbP+wTOgrfFql/qYOUKzMqwJRQFaAT0Lm
7DPPmyAr9n+1qH3rLOmw6vTijNWunQY730bv7QnG3IV6BbSF5dcrCuNVTJR1TzRhC6t4k0kK0qbJ
TzAMsoUbFsXcME/v4mLZYqMqPDeg1xw50LbkamOTkM3JGkHx0gP7fj7ial1y7IA2Kv8aDl5tjzoE
/mH9nyUmR3RimOIvjZSjttlv4jDwEjzavfZYVvFClVBL2I6oA2Lje0f65vbimOPUydr/lvuKuaKZ
pX2Gyt4dCIV4oB9R+7BR2yLOcaMiSFfKC6HNi3LUfSsaYd9YCiJ84c3MtY9If0ZTkZY8YcPfyIk5
wUHH/QyeHh8NCBzUiv8EHOlwK5lAhdu7Kp57NzExqZgQ3YMbVPjuV8SWxlCFmvY/c5LY6b3GX7k3
YmLvYCV9g3JBQU/W0YPN/dfR5UWKeDxEHRFbaKD5DGnWjGk5kCltOW6+ENdFWOrJ+sjo6lvesBce
t0Lto4tSm04yHVbCgr1azXvV6Itm/VRpMh/S1tR3Sur3uo7vcsFNCImPZlOwqIPxkDGNiCX/eaoC
2rKMrby6Nh13Bx3kFdZqeEn/rUmx0IyYRjw5W20SgQJkz0bGpEdRXzH+1d3t96BVhS1Q8YbfHB0Q
sMoK0Pj8Nzt8NN+IRecApt6OtDJyhZGuUc4dn3rhN/zDQMo2YmhGgx7alhtLXcKuGFVuro9VpFoX
eP7AZr2L6h0Jhpny7qfuACAuq2IIvfrx4rSVP7IhC4ERS/qX6LA8wAPcbGgjHGODVGsOrQrXyzNT
Bl+SIgexlOH76slp7jQayreMNEPTUibAZ66R1xQJZ6m/17VTBsp5Tkho0LmFYjO1oZzbvoEMbZzV
NofRU0PSKaulP8ZdURKWB9K+0IHjweDcN3iKYC7Zo1cE8EdJ3gLhiutWVSgki/OvuM/jjj4ERU4f
npM/G73zswJb/SVOf6zoMOMyyTXf4Lmozf/Pxn4CJS3sIEBRdsZMQv8jBPZpxpE/8rVdr9CXmHVm
r+cReYsJZkJxUYLBDuec20ZsUXigpx1Q5p6j8y/2OrYbdELaacbQQnnl9KC9rgD5LC/RL6OPIDWM
4o7am5Q9WdF/HAadVMS68h04YAzDCW6Lfy8IL+PvYRmEyM1rMrkgwkoEPmZIvQNoTOtLeaYk0x1q
6yHTDD0T+F+EcyXCURH5nUs0M1cjEymq8HA1EQpvDGB66yp2PbLGjDQTgJu5sQNfSUNgXngeHxKm
nH2POiyu0V+XvFJCRZWehvmpzRo6UJR+frwHBCsBP+jNBrNXBjUV9uKX2VSK4P0li9IXRAjdhO1t
E9/1Ony1uh0VuwO1zb3ocIyraBn1q6Pvb6ZEkGuMvgW54uBQVPpilibtxBMIrN6FDRl8km3Z3JVb
5wHAsKD+/3HHxQtiywWO+ad9hOSceqU3HleHO3vA62DzAnsd9DTJ+LYozyg8YDpXMsHaDHp9A+cf
5crLxefe3Mdje9c40PFiiACPS8XN5b+XceXIvk6EB3Z/pUT93ObKYJOzJBDKs6Bvfm2oHBA2XlhI
6Xz3naF+5Dnsx5PXKCA+AGGQS4Ehfeap3qlVN/Za7xg3bR4qvNgvYQ/sI55xRf/kpx7fg17XQMZU
hGVNLJFP4uxEBy8ebqAZVFYx2Qw3P+Ko47QLel3dbIhTjNktmmhvOfEkM/udPUq1lPC0svT5pEVv
hYWGFLF2iWKAAq53qHnwSt6a6BVLXhUkhh+P/qom4MXarE3l4wFsXIph/sl+DbQ5hZfomQo/ysEi
26sWTqotAZLcgw8oY+2MC8KkRaHDN+j3G5HihEW/j0rHKOLtkt+WHVh54gf3RACYqQtkic6skqUf
TmWATLNnpQDji12bQbiQ+VUfswTDS78i9B54l+e3SCx4lUhjPEueh9VZPsPtMsrhgiCKb9KEuyfM
EckdAlFpEldNaSgOI2scNGQov7w133uRE2BmA/Mud/aD5kkWlnDvl2aQERENu0Zdj5RM+XYh/6U6
ZfmNOIl5Ou2WIHEMM+nSHmEQ9LtumQffLiArziQZfo2/d5o1vxCsowNwLkIsyp118IGJgxF0L74T
AuuKMps1QncdFt+zHZ93MsLmCzAUMJ2zI+tJA3cVyJjAsbWEt7ucNFBwfTNRsX9kCG802ti/6Y6b
Fg3EAsry+JET3eZ4pKwAJStCnds3GPXi9xYSzoLSwPzCkdl5KghiiI3cHQKo3RQt43UsHrShVWax
6qVKJkUXNY0W0tto1Pt2boIXmWA2LeQgEuy/SJsalFaf5zJUbuqy0DaOideZhMXOiFnl6B/Dar7X
f2ZpAIrrLQfq4Ee3EPCJswvJNc7OkdQNu3FQash0de9L52LWT3WOKepQQMHl23QD7a22figPz785
mTX4CHlUfrw4IwtCDTkAsK4inWT7YKDhY82W3AR0vvC9cwB4+VYRrI7ZofYNx3vXAp25tqnxN7Pl
pYId2M02Bj6fyiq2GE0UvGSrFlwBbkZXR8qLDzEODbkL1CSWMb/7nBhLjShsk7WJOmC29ajSWx49
EZRjZptsRcawXQE7yR1/ctYE0VpzmvO5O4xPYK9MgG+NtQQtwwgaE2zYhp0ZmWW0mYbcrws+ZBIz
FXf+o3t2qEjjpzn2O7vutDdHsFXbKQm7bhgB9xHYa1RnaZ1kwljfOdk3LJlABHj9GytyOUHQJgrf
9GNypPJnOP3UMi1TM6oBDDwdpT9XqqVYYveEPJeoVgz+pWJ2hv7bbKwH1WoL69UiIzcFFotgt3Yd
WgUeB044CJryJFp/CgqXkORQOIPTy7CMvQ0naFo1Xn3R7jUaRVYGa4eeVkEim9hHvqY4AbTUBj2z
6OcRN+KBe3mZ5g64Hkg9nuLz/ddQwZNP+zlWDcwH9a3NSOd42jELxbh6HZAAfpLLXIBcFELCSbM5
biI04xRPhhWN/RIW1xsNjvp+oESg7VU3vNc+JX+ytEuTCD5b8qIAR4AfVfmeB8KWGTDmKJLJHC16
4V4D/2uQOfLe/i6gyQ8o1LsZ9cPGBwYW674hcXWcJzLRljM6If48WtfpP16545+89TByga4susa2
Cjk1SAlrJWfaVKm8g68GRH4WZoBIPwpeNyZUYvK5ZG+DjBfrGQZ12JWyp0HMaNBXVmr+fu3YxsOo
Y7DEvtnMk1Q9PFO9UE6tEc1hWhKaBJOsyCIYWh4qYZEH3KZ8f0wRAhYIVLW/iIpG48sk1Xw2q9Vz
qA8zomiAs5Zi+Z0DgeQevr+MRgan3ewX7+7CHxBGZPVHBK9cAMUyLlM8W6857VmhdV41oZuRL1Gn
ezeJlHzYzKlYQv6nRF12352IKVe8K4DoOnm39MmWFEc8h4kfmn3pTyRJ4goW8bGPy0jVoHBiDsj1
uvb2+v37SmoyIJJuJNEbuft7PvyowRLxinHl2IY8xTYC3ewreRXaJdXXFldvKUYK0TT50EfAHk2M
Yp3FCc85zTkEi4+/mmD+u5sBebqPDVNe0OPncIgJ9OHa2gu61Qic0XOhvVjOIBkodBbNr8wpSAPp
YDJpnJizKU0WHL5Lh/qYbt6/HcbpJnpMm4ohT/mko6Q3DGgUGKQYzxgS/QFG6mSNLZcPyWBjKL7z
BOy0Qv2hPckVwH66NaGtH2UGbkHpg7MNbWtaFA9V0GzlGEJ5oULdnp+r4cvgPGUcCeTFGLsKUygA
G4ocFk1A/Wv7AHpyv9yO7Qf1c2YTYw/vR2VPsPi1KhvDc3tXNl76WQt0mXhvEkZjXVPlU0FntnyF
mhsVqtsyd+rBYh9RkuymUJJRNAN7jOGp2piG2RhH/Py6hVrt0tpSrLDnm8FeLkRMACxs+8koao4W
ED6PzVsBQzODSqVtdjXvFX4kq2bJmuCvp7xRtcg9EVkDYezak+m/kKwo6P99a2HMUu4HidnpX5za
TYeNQDw58Qbdv+RPHDyfkFtUsu5qFSYTZ6tuUhpumzJqL2QjRE3Kjuwjyz1fQG+4eNhDvv1Eedbc
N3PgBqf6FbDK9/L1XAris/c8kKbhYVmsVDtM7DD9pjMIHyaN5xDTjeYB/DrJCmXJ/vY/8vHIDB2p
oNjQVUNoEWCVUMuNVY71NjvpHB+2VfGA1TMDO260KTTt5alnMwyeOve3VCcOdOL7qXgqEl/Tki1V
SUTn/NKYSE4dvlBlxywHk0PaXqx2aSgJvTg93FpqpIkiTjXKnQrJsorVxGipFqkT2ulMj23nZKFj
9MP7+BJdVWuIJRoibpR88eSyTfkuqGKlTaMYeXg0aDifcKkRn7GRopKGT7FD1GnY1zuwaQOji2X9
aZLEpkrTvGRKUk9R0fYaCzcHuoJDUJMvfX/zPRYyTVWSRj2NQA/8/Q8V7mZZgcgmVPZqHu1gFjlK
qnRQ1/n1LycM3kjrRl9PYnv8H657bN7yOZUmlJ4pOiEHR4BtWAVKDkhAhm9sfaXhE5U75PC6AdMs
1d3G2QJiOBQldkqAqeypXGIZyq/moxWi9ePlwN41ijODxRIbICHqpkLdihT3svMuN4wiifdv0TGj
jzCAeL1NHHIFS9NwtNMZweVtmA45vDeC75SK1Yag5891EJusTyz2cU0RNkQHPUJdUj97Qf3a593W
m5gsGl5nxDKk1XztqHJRq21l5P3A1iLLfhOiTylawD4lgEmc3+waP+hW76H4A+ZkKycbyHL57vPd
uV80CyQj6DCqF7Cty4f2RuGo65qbq7xLdHVTRVe9wkDT3L9CEfhZUOiJTJ4BECO3IVB1gHJcUS3A
BQgPVBbpxu8R/5YuZG4HGEjNdK720PjxIKIfRpseoL/6FrWHu+1Ow2XsgtGG9ZfDxdmF6byhnBR6
arUIOrC7jXclhc3cZX4VTJOaUpEADAdcdEZUXZA9WyDkWs/oat0w9tzETFJtNw8vNVtPd1xRHEcs
IkT7fnOl3Th0bBit+aWMgUr9rc6+E2bLXXuC8qJwIbh+ZTNCzVc4YdGv0HpL+w5WGh30FsU6FiDm
PRIgCMmWNzFyQLedwmIP7JvPfZq/FUrApeLs1aa8rnyfrK0yldoqRYHvB+nxK8QuyeZN3uIv7hyx
uNskB4agD5yhyDvTgGs+wsMr4dKl6X3cfkKfOjGbO25VoiTUUocwO56nr5ZGNsu/xsgS8Ihzrx4p
ADmzC70ybIrSPXcQa88KWgkR0EdfnqPPjSw3E/dSPt0dsJYS9/o8GxvhzVrwZSJNo7PC0u4u2l0K
mGrk5v1diJNpWia160UhZrSTK+xJkitbLXx3K4fjk7gTganz2bO/8Y8e1VB18p1szRA+IK2zZ0MA
aUasHr63XsvpuQrOMh0ycGYJ6eN2Uc6vo0JdgbmIn9UZ2WB+yt1OO4DPbM2x1l6OzY6+Ftcwq5CA
IiOfCFtuOOkHqQqmVJPbBpeJRSzt2QsCJoIsJr+eZgtPybQl2dkhvP+4BtAesUGx6fw3C5I2ox9f
orWBPihyt8OLCV6ih1T7D7PIm0U3GeRROPRXdORXph6S2DWyjoMT0MSiPkdNgk8IRV5eN2ZVgVdO
fi0D2JB0IhaGZ/3vf5wqs1ZPQiD5iA2vYsvyvwGAmdeC5YGcBdOpE0+8qKYGvEq+OcQIRfQ6KzW0
EakwBf4CYCA3iPSAdWSMlB1u2bRMMR3pivjW8SYWUrBq2sjgmdTn1KXrZ8nuAjkpVLFRQ4eOsYZw
Y1h+bKgpNgcJFbsey6nMZ32XOLWsKkd1/Ku+qtdcaWlmPhxoLYEuPD5gXIbcaay7Kl0Awub7OL5L
939HcTgfb5F7C0aYqNijykElt6hLS0fKAN+PIcB0cvbrV66Ep1UfAQVqNXrO14dyWML+WCvfxbk1
R3HK6MdkGTOQJv1zS/B6T9aArzSE9N2gIDKq4qi6ui7ozerh/eUcEEiqd6CJvNmtzbo3uV7uWiKc
LvfJs88CXyeV+qoPHG5bJXNDCeAAvyslxfoO2OO//r4dUa21M2qR0ClBE601+Wc784Z6jDF6f2OO
cjH9+Hb2dH7CFmQ6qrjTrK9F+bua0/cs2zMkDK2owUs6kCzQUZWc73NfaGJ8TpIQFtJzyCP4ZI3U
g6UZ5aaBM/JTLyywd7sMcVNG5PH1rlNrWjosB4lnte34DouOsIKTLkQboI2OkGGhkjXd8MC78qpp
fCcM4RHiNYYwlY1BB/2MqUlSM+qY44EI0N7u0ATXrVbYgOUCjzW/qvkxOFoSXDUMXflQ332dYzca
ybesGSIbDM35tdbSigT65IIYzep500S98oQxJCMS4Ej85lYb/EStSb0qj7sLHZcfm0fnwOwR5fQ/
0pvMW+3QrGxpaO+OKWb2S4qk7USng9sP+XE+CgthQKuFPrAY4z7I8BcHIyf7Jf4H2MJV50GeUpuQ
8rNk0N4XG8KJ32adoncshkwgt0Kp0sch5fZ23ZvvXwOF7CJfqiNK4oXkNq0fLgBikC7ikV9VYvvC
FGkkz6plGpdSjr4JqI8tpnLg8/8ptTwz865gu9XB8ZmIvYRe6Ki68mnW6mboMk9LkrKctMndQcy4
xxfVxXS96TMyiKroFUdz0SQQexRwkEN6sDpVmf2PlC4u6V8c5DI2DwPyX+J1njRP3vZbOSq+84u2
hLghkx2pMBlYwCQVg+tT1zwvqVUShE+3Za8qJxPpccnLk7uzINrwd8lZeG+/KoTSPC/XXam4OcrB
pBdvlKYW0/Mb3g6lO1VFDYmiOUtZjKQF3lEYiX6g8M/ZTIETPhDDA63GcggNxyQ5xlC7bYzWcdqC
SHApBMGqIUUJRICzWCEaFhD7sBcm0gmoj1jmWSP3BYRqriyAKBo14DtkhvsfcXpst+PBjSuOO6ZI
ITChhGXUpIGry48UdIYi5AVGJ7mqBqz8/IXuC81UuLz9qftw8qh7uJ1XQxB1mRZvyhEFrPvcE2Tl
xb/9gLTAf8i+L45rQ4QqtM9z74OWCnb5BBHn/MZ2v0oc1ZafUvVVnkTMu5eddeF/IJn7I7nN0edw
lrNxhAjSRdzefZihRcDztBPvriy9jDDugu8tZhBvsd4u2tleROtT2I6cUDlcUliwgR5Iz1BcRMZW
qCm68f9IS/24jJ1F3Yu+xwfMLOOMw1j2GosgtrKg/IMexwvQBAQscHuU0kw/leAtXLkJjRAZu+Od
/J8RPyDz0FWvrcU1QMY9hRNuEaRemXx7KbH2iC1eSEwXCTN82IXb9i8rc9Yok7liNXg5WMZHdX8V
vKYDik/+HuXWXUErKSfJHDwjyfT7p/pG8zbwigJcafyn8kuFYxt/bEgRtubEG/udscOO+xkHTo39
cQ1w/0HzvAhV+BocwFq1w1f06RLOqwxznvoE9HnMzOdMrMyGXIelBvOj0J2eVNFtHrQq6P6UIFA0
NqKMQQilHs7B5p64UxeHRGuxCeeG62nf+USRFt45AaWO9g9rmOn98AAe4dBaRvMvfHjs3hTyJqPH
4cRFzUN7bOXus2Gn5lRjyFtuzBKkRJ2fUJkGhhMZXpCjnVyCXtri9KtCowhIvcT45OYicL+ifYiC
35lXCJ8+jWVYcDh4reENKnaDDY07LZLDYAbsQZ9GpN/8agI7i39apwWJ8A72OsDx9J6G+zdx0DZN
sJMmd/6hVkXx/2bFfMXK6DU6jKC9xAPOGZd+sPTiNMaOZh49/MajDdz0h9NsP8rWzqv6l3XP4sVA
rTMhUbaGTc60JCG0QVAeqn9pBhVyrmtqlGqb2vrEDU6V40edUe9rAmYMYbM2VizrcTklAZ5Jsg+H
opGJQsRjXJ9+eVcJIN95AlViJByYIzkD70TPvq8ZB0qUWwiuJqToCqy5fpBLg6y7GP/nRKKFYiBr
QHEGdN4xv64qn7v6FxbueD2wGNtTlHzA+sOlqq8qCan6x41rJaMQ0GFxFZdz7z5umHxvkFnzi713
btKHgnuV3oHdqHJMiEyl3/TC7PU+EDXE6sDsLtAHxZ4XwqS82+w9WOxVr2bL5G0V4x3kwIUcnDoo
UnEGTtv/16GXROePKudYX7V6qBN8TK4s6JXCEzmWo0XP1Wf7y/vIIeFHNpo2C9BYvbAQk4Ki1Qcj
Ziu1eRO/cfRTVH+K8XUDZiWUER8Km4L0wl1xQfjkLzaRNspYr1NXYDdbZ6wpBHFCYYsYbL3LUQ4I
apVuYz0sh53kb3eaWGHAvCzRyXdsXdgZeFkCDEMDgk1SurxNq4eT0W4/K4NF3EVG2m7KkJsxhMpi
NxhkR/5N0GIaeGGnuItfGV8o+mXxN1zRM9JZ4btbC4FuK7q5CBpS54ZztOgIqA6ha5YM9NoN93B8
nKDDWZSxDRm8H89EESdLofSdr1zE+k0F9piUx4QFWmX77YOu/Ve5irR+5vjBMs0fVDG3d7unCu+B
/1Ep5iVUXfXiaHvwMB+lCN0d5prRMsdoPKTB3E9DEwds511G65ESAQuSFdsKkN+tFofI27Yaa02O
Dxk1mrhIzJc/PAuXIOAZF+VyOr7VtCOLF6XfDh3MhgCst2AWF+PVd2KdQTel5r0Dp8dOhV79+PQ2
WSMvDP+dJjgb8sdW935v91tel54OuA4Y7zdMLmZgakI0rlQn9XWrRTE/BETPZWQoAi6CIwHGkWwf
R2AO8TTJnvxx+HmBsAZBhxlZETDt9KVerqOSZjXEAMimjswHKMauCYSoEst6BbJklxn8/5P5d9SK
KssVnnyI+w1wD9v22alc8F/+P3AljNcJCb4bQwf9w88pmjL/N5pEYJMB7wb95cb8K9+KATVSQ1+l
I/pIqFwBhBCpC5Gv3XSUBEr1RPMOv7ZA92KL7ZA+gOPYb67UHN5ul6Od5IL9KwlwUo/8x25GYSjl
CStisn2icxJ6qVJFFOkqD/d7E0M8JKPzCRxMhYfqN/VdoMgfSXJ71QZCjSbm8xGP9th13vjo/LVK
9Ya+k48RQP6bFRoAGWJcuwpxDIpv7CndmJ8KX8rNYQye/+0D9qTbY+gepGGfVFVsi2EwvkFdY/ns
INrOLD2G617sDYNnfsYr3aMgrIIO277MvOjQ4nb1di5xncm6CyQZY+s0X+VyndMq6io9xMI786tu
bChGujlWaR1ZfuGrhIuEWG/gseI/AgsykT2qt7P6BExFPVQOLoSnWP+Dw+nMChnd1mO+9qH2H3U2
pg/bmRUjX0k+ZAenz79DzoKvFMN8f7hYd5/nbmcPV1YQXX6uBcEej8rTuimjLaybbrzWp0VitMze
SbOoAnbzPUByNzB8bH/m4nEQgDqX1F0t8KKg0ycQFoGa0Q+H6z1DZonCOFDVMvSrOo8KhgzKNnem
MgZBjyNdEFrUrfoBx+0oRilCGJKUWcLymNK8XV1kCeyzMthO6yPrBh4YWHvNm1mWiI3A13CYeGTT
8aKE8dB50SoOIRfTmN9RZeC0KKZeoLqmwQJjRah1tBJkbb2+Y1VzokY6Q8jZ/AzEVgsqdtYYaz4b
7cPvcKRgggYUy6A79K2dMmGDi4g1O8FaJDyT8JcFzlt+aE1nFeELNZmY7TO/f++AEZ2dqiynETe9
LZKtHdI20CR8wiDcLXDFo2DRO/WDST2wEUFHUFViMppuFZ3TRSnutBiTjvHhkbBZHahn96TeAsAg
JvV0wnXNzECFTe1ljDye4Ela+rwngSv5eUrpTlm/Y/O75EeU9Mc5oxDAtRzXooKBby6piYL+AO7Z
nDseYz/t4rbq4RTAbSe0Rn6QA7voAehi6CPUzITa5FJG82VnF0TVpEJQnTb1RyYtiC5OyjOyak6s
FOcLeNKX3uJceEhrwl7ZywIicn/6EW3LHs7I1w33FiQHfcLWerRlL7wAW52Gldzr/ZuY/awV1RSN
imM6kDNWtJPUuXo8lv9C3M/JXsnpHKdn4DuMHwYoutqXg/01fBeBTA/lz5ytXg5hIGcDeoLA7aTT
ktGql/caSuew5ZnqOUgyJmiSMdLKO3tAxw4u1mn0O8IcDuWFqtmsWNZ7Vgb73YVhUPcOtW43qyTp
yghzugWhCUucVP98JLkDR2xDOVPuj5yYW+D8v2cEPx+nE9SRYetC8JC4doyxoqICLlqtM7yRrsmB
ttj+j+/cbIzKz7KUTieF4JxbsudFM9PI5I1RIIcL/KKAEneSHPRthClp6avRbSGuKE5NPztRAuG8
SaN7/IZISTVunusA7t7w8WKj4rUaKQf+KXczMptHNkTGGxoasdxkyxBoIyoAAX0H9CN3R4rRrbL5
XUVYX60GZmlINdbu1gIzlsIHlg6B5307ZKkd6OsX8lbkyRrhNtHIY754tfv3Yg5x32hLAr85HS5g
yFpPqPVJ/EP+4dQgsX6N2KyUAaYU6IkV7NH7e5T92UiiI8q/TkMbJgV521XvdJoUbhjiCF4lHq7W
9l50rzfn2KvKtpsXQpBliZ5fs/Ce4D5KUVHz5q1UA8RdoIRXYeYtrSbySwjiELR4heVtyin6L8um
e2fCZ8PBA88wi6bXdRuMy8jqA0iK2Rs5wAWRv1uBNL6VfwXfBr7ZtOxxeFIvqIp6iW87vWgB/R3z
1l99aue67KgEg+E/plX1cAsvtf2O+HxxeAxroyOojU+B0N3/jHW9pwPqM+ZlKT/GkG70TQlRfDct
6SfvYD3g4DUbmzyVhpmA9N4RKpApmNeC+nU4LD/YWQuPcVxa90LPBnibOUS2QKYmituFAgbBGgkT
dz5W6qMNGulaRZTF3ikdjilv0bCarDzA8XU9GRcRU074zWQTDO8L/84JDD3pDA9OvHD494fgd0B8
pYvTDTDhmXx6mgqk6mEoTIJ3vr5svMmVZ9xsYw43yjNuOXRj83jjqNRxxqfupgOXuu6Q4hvXvork
CxFhZzggNzfPV2wlHN5Sw6LcKe+N/0BD4tSHHpIXNegXk9X3O+iMs9hIa9yaBFIgy9dp+W/bDj+p
wgJq4rpAIMhmj8F0v2S6iGkMWPkijy+6z5DdsWy9D/hPvxmywnl3N7Xo3DfbZE2363mdNOYPLwod
IOEQuJV5180SzjxLyWy5lVef0iGDBj0rFlvHqnYoU51ZK/OLs40mqrhn0dQIX+feoShty8mDC+En
J+YAjutwbfdB+nMgueyo49x6gWNqtNZwRnTYcUwmAKhzWwb7ay7QmSuo1Sevs34Uao5KpsCs9wL+
t9ZCaTbxus+fXHS3QIHT8xlW7KfH2KiAIqno/I1+Pv+C+elO6OfbFwLgqAHfZ01k732I5/wCm+So
DeSUqvkNeAr9mqIngG5u/XW7//zBkrykukhz3/3dQmMaIr439V9HWRSe/S5WC8IwUNjBTmoWw3ja
MbZ+jXV3jaKFCMNlPuyZQ0T0NmJ5pblXoFmQ3JGMgWA97xNqdE7eIfCvFEthkJEexL3Y/bXqZQaz
xPMXJJ3BVu3Dm9KpsmRkxDG35nEV1oaV9o3uuYvfE/Dei+W5H+SY4JD8Swn4qznlE4pO3qb7aKXK
pzbHwwazre8OH17xlkI2X9KY9mdj5sJRPnIf0pyK/SDwghuO2o8epFpEBOrx3cvOLszwYsCgWxxV
eUdW5lUI67sI6/Xuf5ZCOTB5y8/eesXp5CgpfwwvFuGb4VuXlqdCufegd5Ww8Ps04uUlOxmQhuC6
VSypUFhMV59VEk60NLz7hjhJzEEeqDwZXInh/+WpgDd0+u/5Vs2C20VuUnVjKmBxJNJEfKatOZ8D
pTgiTNrggDGsA95Dqgl8NSkfi2cTVJcb4EbBMXcCUvJSG/Dfg37HN+SCtGWRnxe+ubWXtZbJFQ8E
+vVYaTljCvfKhuSoJykFEpxOkPz544/2XiFgdcU9QQiMeAObdCrTUm1PS+MiaY0C7jKyu9VBac8x
3E3tRtjrKqEs+Wf3AWka5txCHoKUQKocFWbz2+Tc3l+ximorrAyLj7CCUqf/pWOvUlR3meF+0s8g
Oc10G7EaSQTHKSuUc7nS/I4yt+EHO4fWydxPD+b3xMACF2BWdEJaMsNDN0k4ONDxxZr4+WuofdSi
uWpmcPxIKLcG/j7zN7m7prOnrfhaGJr23H1AoZHm+YR47A5ycOrpx+cC9mZ+gyonekOFOw7/hXRL
r424CDkCMUCfIb1xsigWbzBQjEvQd+GphaNcZt3shiMaQniF2DXirnkwx9EKBEjZyGpUyKTuiZkw
rM23HXiIbkKzlFLN1WPeT/Bl3R2jP+mspC0qWYxHAdRprQPja6y/mFYmJywXjqlCWWxbnI86MjKh
BUUYL6jlgBTTYjsJSvW/h6EWU7FJG8w+g9oRfAIzfabdu706lOoZPI+pcxG1Z5cqnKT5oS4Ru5+V
hGrRE0MVrhqhgL2KUkKkPYe2yzGBH6CQFKGFV/X6wFjH5VcP6y6BIHNfUmAQUXB7iQWtus5LNmGW
Ms6w1Wi6txrs06QM4xeg7XdU74qW5HGyOCgQkFRGY3vFKe+y++7nfGwjBH1iiWnwHpqtqucXiKz5
at0IgY7RlZjCbXa2dB8k1gfMAJk4ko4Kflz7mDuhrdL2c27QevjWGe2F1e5LflfqpCIASZSkPpEM
8lRU6W6X8ztYHvID3Tn8lrY9NDtRyr8euqQ2FQQen7oZzXhswVAUkQneUoX2ts81Mar+BgjKGU1Q
iWbNMt9+j7ostcC8m1Sb/HtnUE/tjDbwRImuXku9QSHd822YXOAXO+I6YIhtpKrew2/QGfRRN+NO
Ff72U5JRcNQrSsUsM71LtHVjQ6iire9Lq9rX+XZvMpHB9PX0DwrCSO1gKXI/3lYaXuqHqrHb/dMJ
7eStdkMBxWuiEO/TWrRAwng+9oEYGmk8u6c39XueBovIvrQSB2IoC5DxJP8Y5Jm9IUKFSilEVvah
vOaVGYXrGo0BmjO/W947QQBilfPw3rXeJA80LOkIunVOBi4OGtiSn3P+20aDfSX5DIGjTWKscjv1
Vv2UVggS7/cfxftHu0EeA0nY67RZCR0ch2yonOY/KDGBmnYpSTZ0QK+7XhI+huRwYzfSNalp9GrJ
vphnOhLWL5kMc1ZZuQ2YvHjeF/Bk+jHdfoCkjUgrG6zgO29gEYeEbcAVovswnVjoqUC6hsmeOPCW
fKdDO3/KJcWkZcxzqDM3/O+L1PvAInWBuXLxJn53LlQakrnldfURKOeO9Jxu7p2XAs7g8M3nO+3D
Dcqtg24vpwGnR3lcBYOa2q9YoWe/fFAqsLSEd78jrWT/ypPegH5+pfRznT5kaa+TpDdsB13MuUv5
vYuMhYTWiAKMfWnvz3dNL3HgJIG09stjHkWL9G5ugxVSNQUhzzty4BFRvNlzyMHNh0QblZz/OGlB
Gp8JQ1JB3pvdg5jDzU3ZHibbkhTyzl6yDT8gQf1lbpXNpvay7TpLjOkv2d3JzHuTymzdDAXs4hIX
Jbjlc4Y5996axLur4pVSKRR5tRZTq5y7aPOrxBp8kHf4iDETsA67/0Z80fRe76rUudUluh/YqkVP
krnLz0IdodzZUcrXQ3ZA+xsHxJmM6HW4umrzN3VyryMOVogl7KVK7DAdATfEoNgbfS2iXdSXzBXw
0nV+DxjRBHz8wb9CTVspFiXqM93EtQ==
`pragma protect end_protected

// 
