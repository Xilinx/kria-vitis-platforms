/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
bc4WnAkqx6dlMsl5fn3cAprcqqxHUHgVY/ImIQQum+cRAB7ouhGGGf7iFZf77q22uZ5IUqV83Quw
Hyk2hoLyHV1tsHXgJxRTk+FG0z8kNO9UiseME5aOM/+f1fcoxpdwoF5Nb9O6O9ouJZW/9wU+cOBn
deDxs8Fe2cl/gc7w+7aUoFn4WojygKnIaeby9NCvgShnH90A/5GxWomjUdPAdBRy04fmF471qpG3
rcDSX8G6arFIKQEh5UwVCLxQIuBK6e0cztUh2ocE1tgu0ybaWCTYOjp5wNkYHxW0TxCBiXthO/Y0
21pIqRWTmcspQgDYTjUBBMfo4xnplJBqhrkXZQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="ASJKkguRF7cNZtn0GfYOwaRh6RbIlcvsA1oAuucVfb8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3296)
`pragma protect data_block
Xy3DKr6jQ6T4G9Vc1bujRnKDb1axZ1tuwRcXu2EmmVax02TvV2I6fGFfcdOJF5FWxpvs9CskbPvn
DfZAZ4TMOJ70wI65PXKD5D1rI2pgMr9jjXDB4XdU3AccSNLsEGAngi++0SARYRv/NhACdFU3yMGj
+cJHcfzXM3lej16yje8R5hfzHJcTFEQQiwnGT/iY+Y1WyBlyLCH4LAGq0VvOHhSEkZpw+aLJwDro
hLMUCUhpTUUvVvakyL/vU7oIq6kWnvzjEDETvDqj3lKIYtRb07ZGRf5vagxPgP6IaEtRfWp/GK8f
bmbctDCj6YBzlsX2sNLDbTOXbqfMxb1rt5N2oA4aK5pEyfJq/UZzdRCGw+8h/rO8R67zUs+CD07m
3xDzS/Wl2vH9YFp5MDWcq0MDbcrkfrnzo08zaWaKA878tVyIP1/I2maFpafhdn0utrte8f+hg1CF
iCkTBeRkelDXNDFKfJTk/YV2rcCcWmM4t6UjkitEoElPQ1FWQYGWpPVHbv4Sw27WFtUYlStVeV2v
teR0t9Z6195d6JiiYKxSUrm1k87OqpDqjC8S2lXmfRXRRvktVtlzUqh5DHJ03nPAW+Kwvqzow0fn
djqhz/MzcdE6Do848eCVYX7l0wXgN8xoE/hXbL2PFTzfTARjTnsEemHEwrExXCEPbLh3RoLqOqzG
QZVISYKeJVGBG9kqcH3laxv3KzsvtxEDM7liWD95oDjHccKM3+jCa+EOo5B4WVycM8ytGD54OZnL
gOp7ovVw7XL6B7GQve62H86iykcZZnsIDUWShP/Bbyu/9EmmyfXwzCqELLyq4+CJ2MQtqYmo+3SO
ePMkp4jN8i1TqBBXaJQWIRiXg6mFgR40O/MBdVMO5pWelaBcRvxMf5h/zK+qWJtNbhVMs0tZVXtU
oj/0tkyW8+1zakrYBTHWsErL2YS3NyRMxujzK0eueBfBk8kbEjSUjT0Nfc8j8dEmVQXq/g6ruObg
hKpJ54B7g+PfvGnMWvTyG9tVX6jZ5mjWsYkevA2KXf5LftyW4jnuqxbjSYZw94RcTBu6U2V1eR3B
CjirCIzH9e8BL5qvIJeawtzPfbGUAOcWADFPv1u8gttY5jzWedqNCrccSV60SzgqN7yMv7D0PBxY
QU4lvvoTGZGe6WwcnRirvZABqjaG7+QxqBDgMpG0XDwFAhw2teCkQUj4uN6VhJeLt4gGGDn8w16+
v2iItLoR8fjt8z0B9lAsrVqgO4aHBpe5PKrUh9lYcUpvg7nOvGQ/EF3mMGdsZCnEH0B8fy0WeRNy
BakOGQN2m6AyLrJrOSdWOaIkMD4Ad+FOLZI3FLLi5ZYMDeL+AOjISUVqgSWiEXpb/a+UyNUoU5wA
mbkDPoY2TIxz3GeiDqFDpOZMRPnTjDCFDuv1njJtThbn7UW44aozeLHzRsjyTNTlpK1a012uHTeB
R3RMMS6CT1FueQF22RQE9TAExw8Rtp25rdVRUjNpxu1nNZfksQYN5aiP7bPhqIxND9bahjD8zaCL
38H3vUGwXD8CEuzEdbOrKKQkpfa7Z0d+6GisGZhzs85oMt+ItKAySTAe2jWxdGSFWCf3NwxRsPoI
SJUJXmZYtbTVmourdkJHh7bQfqDAkSt4ncHJcLCfrElkohzJT+YNpz9i4SnV9zYLxtp9RnHYNE+f
qHC8VM5icPgI9HAxb2cDO7K6X9TJUc2rO//nLnDHGe2XdfbShqe4haO9vbgVQCeQbv6ZB1m7fFmD
8dMgPkac02kZrBTAGFyCbdguVP5yiq6yr71xDKm9mSOPXNSQGufwQNAUrkSl6JBA3a/gh7i+FTXh
FA/gNIa0yUPymKGXRmB+mSeLrk+db5uD6EV1ecvvk3gPSWAeHN8SB7nEVrIvGM22MYmhFUhtQjn2
IC371I7S9vtObrIhs0jqhY9upRQ0R4PnKN5b3nyUlKULhOemyFbaQK2GI+rBHUkASKRDLVLuhd3G
Axm6LyFSQDFmEoCchkVjntwhuz5aLcBtFM6t2cfaWk39L91dwdD/VkQPbGwv5xcWjiKRTb+or9Tt
fRQpbLd+H5vR9IK8E8c+FeVo+l+fLPP4Gw1pGgz9KcfJT54NFwzzFO5vLfWU19LmQhBYpcdD2ELo
BckDVPZ8FpHw/zQnQLU168Lhh0R9icbTfDZLzGfiZUFYu/NO/r9oL/nhCdHtXe9D9myRETi8+HKb
c3zDtFMdoDu34AgD1AyGUfSpzBduagSBEHHKkHHW93L2yTJKZt35ucwL1Habw135Zcfco1EsK/YA
xS/6id6ZYRZPiB3hoqATo8fJPhAWcmHj2Gjz8PtW1Lw5nFrOj8vbKOxkxmfndG/hdHAu2s1xFPaM
f9T46n0OTqRpbFVDeOZVlqYAjk9yVezFLleb2zHJTwrown5SMy9GrJVfHDZDmDzOe70HOg4QpZqs
e/pbHUKeSzqjBTKmK86pPanJ3bCGikTNRpP7d8EvYOEicA9I2TUknIov42O2jsECw5NsDU5OaQjs
j56MM1HBpdf4+fafYFbKueF7G4dcXfwRKsPCXsJpAAlXA/hq3rCo7FTuc6VJZrxfUQHrbN79x20O
d5u6SVSwlOYyrey2NbrmRSbA2FJ+ZPbZm1zGU7wGmdTICDncVsuxDUzNC5VBrAqjGZRBxNBF3f7z
KKxTOyY3iteYsfvsg5F0XydVshoaXM7VAsJE/Vkeh2fGx40CnuQN0KsRPCfPRWD/qhk361svZIsI
lGv0c57LLcQdZ1YS6IsWCLjc8UEzeqDrpB5WNH9uNR0dVVC1xrpslsnbErvbiUJk+NrCJBdl0lf7
EQMClVNZom3jcHElZoT+Y8WHncyHHmjsf/L5C/JhXP5g2LkbaPv+0aEeqXYFPHDIFKXQo/Q9KPeA
er9rptrvzZ46cf1JpzwBppPQWX1ISM7LXbiDjZUx9EnYUyiobvk7iMaZEDtnoBXX6++eYMUfJ4Q5
YptcJvu0mfS2XPw0O8MNZ1TyEg8eNwKC+O4N5UUCG1pf8iSQEPMcvBWpWStZpuTUy49kr6VC9cLZ
8n59IEXwp7kufzlgLulXaG27kVeSQ39MEDSjZsHou0ZXvSl6tQdC2yQaMwfuorNW3WFkxN7/ugq/
gC+7JsBckgmuHtOOU/i8v2f70iza8AjOYGdA1fX/55+lEClyBK4u/sJYCfHJd2Tqh/cjAw5gI6tD
MMm4Xv8o9YyLWPB8jb8Zqpq2sse/kNBavDmz3Ok5Vs1ouVKg6O00077CjMxxRB/VkBNvfzF/u2yB
251wz9ujgnGf3mS9xKEbh1S9tw299CRQDqJ8F+2MWvzUKyZjb4Rju3usYpOlekXPEOxCsNC23o/v
XKrSKlhYoysjFDYZzFL/FzTru6htISIo3L87onYzRi2OQNfYif8hGZpwP8nkXHY7AkDth1/LPN8A
xQ47zBv40h62sjd7SaibwJzw905cX72FwECSwJQBLr/wB6Z2LsJ9/YSLwHfs2KoQPjjJsSQVNS1h
O2REepZdIZfr95QAi20HqyjP8J9GuEI0vjCd34WlmwHkUgLrFf95vHgyC+7PJz9V1Bkei2i4j6s6
PJpFtHTtnUgEl2ydEYb8Z2vlEFhwiPJGNMdPQ6XjQtjZmoFbi33QQE3mGA6lnj6T9kzItQb3o/dL
M4TdBHafRmbL3uYRxViSInKte9zgxZQpxEu4pWpprIYg9Ec1ey6+lR/EM6oN4ydqs6PY5SI5Q/+7
4CIIsp3tDJ0kWbnJ4CwYvAZGDPNbWaTS7LkjEQKEuo8yev+zY6bMOEPHZWTDL6ArxxDkDU7ld3GO
AGJPTfSbvIoGlrsr8ri5Gaqjk+pI3MT4sP1GAO4HPBdjA/yhYH4RWIf7K22yglJRtsqpGqWNlNLI
WC7Mi782bYkgH45TQbmgL+79R7zSR3mOtcy5jIseDhCmXc7enYyNda1pi+YMsOR2OUe5scLNJ1co
TAU2qj3IdRjqUR0yEqa87cK86qdyqlxK8N7LeKujb1IxaGUc/g9Ow/Rh66bPdBf8nf5efbGejkho
nL4ZCO3GsKCd/SWwiMloigcp6IbuiYO194XDA82qcxdh20ytzIWv5OWF2aC6sC1zEgPDpvkDWLZX
LaMdsD4jteYFj3wXwxpEPTMIGajE8UOHXrPLoqm8J9ULgpRQTUPOYl9UjNhJGnHbSepVWqMPBP7H
xyoyfU18jcyPubIOa05AFEHVb9TGg6FOTsDYlBkBSXHcmLOGUyr1TETZGD0WTb1egWCqFY1hUzmO
eEdn3O1kdGgu+g7cV1HaJwT5un/PoxBYD122L3s3EUYBz5crYbxiIhcOu9PKV0NbHDrLRJ/gL4d0
UGGtp7O4zFZjLl8ToxasBjPM9BKx5fd57ln4nlnxuDIrPDnSR5zmE8uoX82R8Eo=
`pragma protect end_protected

// 
