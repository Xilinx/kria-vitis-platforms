/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
CaihNQWwu+qKJWjcmdIgzgKIXQ8l3vMImmWHnChjYqoa51yMcErBScyiE64YZSDih9WCUqsVfjEZ
HfdPZ9ljuyASaDAJWOBnJBbhrePBDPO5jKkFmPbv80QoBXSWaNMFc5sW0Ulg3lCiE5qq9SVr7IMd
vkFVewJkI9IJKPXIqEiYLMio527A7EkzJrjUXC11BQnTYghbA5n7/6q2WIDOwjQ+BdLZXxGdIUKi
ihIieqBZEgdd6vwETSGv3sSorIwnUPSueC94L800xEEoFQmghwgPGvLA3IEIqt1YNZfrY4rcuvTH
rxE5ve/ar6tMYP0QdSitAf/UOVre3EWtsP+Jcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="IxINXwVvXQ/n7KwTaYrPoEaEACBK27oPy3cRIdl/LOI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3008)
`pragma protect data_block
EiGu1ShDtOnFp1/lwt6VhdLFiQGwTUsYQTz5DZx11TvMud99m2FdMW+PHUhMkLGt3KE5Y11rAunE
YznnnGpyww9YbDLxxYxQpjrzZFquVryKG7pQ6GK2V6U9Qkn3gU1aD+G90rGYuFLdIExqa8huwsLZ
xxEGBZw13zObAEbURCNmeqF1OfOlyP+vtLotqYGaXVLusVH4bXe1XqRiHTC7UBJSwNN9IQATm2xq
XEPmNkd9H+jUaJ+LI/1fViJ4BPt7bOVrIr2PlEgsKTbDGh63Wo/IeY6GLCnDTXblXaFUqOlP1bZn
h1FOXqquqVokOrllusUnN7HspaThkYTh/DdcXMB9NxFJTk+BbpJe7pTFsAcrAoz2qJde5XZFGvbn
9v5Fl7qHjnItYUFFb2ASWMxlx/8Pz2PMgyBGK8dmu85I0iyWOPXIo/47lW9aJ5by3wHtgMgWQJu+
h3VcjPhculUU4ZO4F8jU/aJgLw+rLbd/W/w38oitZa9cQpaPhJijXsiMx48tG+kK0jRGLypHXJGB
SIloVrxpi0/2yjNCXPjzDVLgOheDVUgKIQaW/hnvGi9jwzRJ73kNMFvmd+lcH2RDHQoZN8asEUyQ
DCxUwg78Vj/oh8H1wug1XB5xamcXhBueAHc6CUD6tlbMU9Szyg6lbcYW3ceruGxlc640NQlprlp/
WNbNH8HRyJ2oI3G8+P4S/SW1gj5Du806lNURWdXZKcFx8kNHQAmuayiTVm9uAmHYmgOooCoZ+4n3
tvu7tHfQUBMH6LvB+7GEqWynox8YhUQ5yEF7xv1+o0Bbw9uNDEMBpvMf1QipTO76hElTCgsu5GaZ
uhh20YWZ3ik8vX9Kfuehtc3qEq9fYUoIZlbug01xvqWdfFXojqWHE6c3yot/3ebGMkPPvTHRGYok
pW03XZfw9VJkNZ7Q53S1UwCthQ3EY2q2IrCo4JYH2jnI07jQwdk3DvxJDG1CXiBlEmJCCTC+qEV4
9Dxo6t6yBuUKZWtvzFdyXosUKFs3LooQF5D78fIDyTscRcptTUYQWm9yaMSEgv1DB8NynST0C6NP
MQhBcW8q5RDa8ltUqzsLQ0EG4TYrNi5vEF23WRmSHP9x97bLNFL7XPalQV9qdDExEfQaklo25lHu
ErunzGUyj3NXQwd8LmYMBlRv4qkOYI9SSrd8O3WImZyD0yCzVV5okDigC0fiNaI99nzYQxAyl57E
YuQynjz5diN0CBBxgWlCkr/UMdSjZIiyodB7YoiLjfOvgDGipx2y22vxKINv32mn0iycSVBRX2nT
/DVMR+gy12m+ee4DugsUk+sblAMEkJe1CqeNsHbd48YU2iJHkqKRhYPaK2+cs5wrZFOP0ivgrVTc
4BoVlSGyqCHaLQDXUZ9pwDKPyf+1ex66fuit1Dt6rcebYnvu2/mYItUT+fAtV8PL3GUqOIhK8V6w
hkalwR8L1vm0qwIX01zL9h7HxFbAjcuI/Lx5ishyFGvqJWjZlV9uyxHuT1WL+i6vKLBRsz1xd/bW
KeXnVy80Q04hkD7YwP0k3w2t6rty9c5ft11n9DZKSs7Z2HeOTNu61VW3/34vL4Yum6Li4kGXMzfW
s85mvo23iVHHPIwbydpp/yOIw1BepBZdZM7UvxMxvZeLQBStdJdUmL0tR2x6nDrbTSC80jV3dtpj
VLO+oRZuLxzVUu5SfLaL83GW/1pZrRySH966q3GO1uNMXN4wO9wsOxXc2jcyZP0+mypNqHu7LwNv
Yxu94K/MuS/g+H+9TGGIUUbJpMaUAcxq+RKpy1kVIRvagSsJiaIItjh5MgNE/INtVW1JqftYjssM
k2/o9t2jnLyr/fPNSTERHEedefpLGGulpY3e47DEoZqBaPNRQhmaF6f43C4RlxJixDtQ8IQQ0txj
PqIHvgOJb3LpvN7XMb0DTyWijKtb/VbMjCk2PyFgsgeIQUkC6EF6yRq+rdE7+PRTKYsT7sSVANgi
YRf2gGwh6SqXO7976EGLsfwsA/nThJglm+LLeuqwJOJ59jCFf4LOpZgKan77c6bygMGe2L5lq1pP
TpT32J++DMP49ynBu7mybd5vfyaeU1m4dK55v5kPv/3pKv1alogu48dwJ92hjlUzXxYrhQZUsU59
a7t0xlMMOB16xstg9DmlS09I/iEqlZ50fjD7Uvtby52FFbcbOafnRGkstLo4oghDkQhNfaiIJ+In
kQUDxEZDL/CCpOxA2Zd/TxDJE3B9mikZwXeRZtO2IzoLairvnb+BOWgt8TadZsovWpmDuGAvPWhu
S1BKqH5II9b1lp6vcph6c/rUYIUKCEVzPf8RPkY0pHcR3uS4q54Pr88R4z87ffDAOjKVZN4JeVf5
9geqT+gjXTmc5ys7Oth0hWQyGx1QKyRWSDakcESABn+kfYoqPCU4N+b1Qt0C7kGfwQ23xJw1xQoX
wwgALXsgjgqsUON7/iYRnwMm4k5LiJYEkyjyQwYG06FUbi+tHceKLVlePA45YQls8MUoEHt71LtV
LSYm99pDBbIvRHRnxFYY3dEwGJs72BGj8WEpe0l+Vp47x3AMxp70hDfmnE4RZ5DyOrmHDd1nTjE4
YXoW67MoKPYAKJeCjYhpnMzKElyc7W3lqYS+aHRNfFJMjRcK0BLsYTb5QzIotv45+7OGnXEwCl33
jWhHLumgST7D/jqBrX9qqdrf3jeg0IuqkcwL2o2r6aylDe5dAKsbySz4Brj402+ars2TdTB03BaP
TGCUrAlAwo4AzZQgMIkrAN/5ZDqRVqYVEn1dl5DjeCNtMPJA0dMKlKbAcK00QATOkJXwTB0FjABG
DpwnpC22Le0uWJzSn01fDHzrFmJgw/kevVDLAfKWMur5CRmni3xc6HThSqZPsMUlIuNMw6FctwO+
kPpvkoPxVy8rTatPBXs0qrI1i+6MLjs6OhE6TfZ2NnSji0XqI6dgWBQ1m7L3B2edA20aKciULH9X
xQf+OKf33vtRvRGpLxWDINKB289F/E9QThzo3mb2IFT8XWHCXkNq+inPfVvz7Asit5MQ/HVk4DOh
TqDH9iJx0cJkmleR5FIzPiomap6KGNuwxSowAwFvoGiTxColxi8Q+3yerQyhHVNP7BsZVpuJ9gLO
4h36kyN7qBtUBcUG6+KLxfjAaXmIhLA73zZT2sTi4fw2n1zpbOSwsA22VtTpi/daogkASQGAre5M
XNDSOCnafi6Bsdz7ReUsMhIkZ9+/loQZdFCnMGpPzX0ABitqWG3mftol7vUxAwy6waGjQfY5Xgq/
t7oCvD55lzNtdsMAlToDMQ9yshSlidAPSt/QUhCA0cdTz65EuVJFLz6TtkJf7QHQ/+SXKxS0RZiP
xJADGLY6GTTlK5JzwVgs5ToD0TixvAZ3bfhFjRDgn6zsw3Zvkok1ye52WnJ9cevJPiHfzljz2+yi
QUEf2sClCDSaiAniAiksPbOXbC9Qqwv68A1RH/0EICVhF6blkrYvboVbK/bX8mSnG9HR1xz+GoGN
twD6nbtmxnDcYt/OVRU1AWM/nuwyDmcFAbO1WxE5i9O5zZCQbUyS2Ykxf4+DX5A9reNCDpMs0jpU
RP+9nAYA+amxHYwiDi4UIouYRpdbEitGWIdocpFTRZibJSGURPXZL1QVREjaMvjOr82BA2dHB/Kb
TjHsCxd0jLYbB5WQhO5EuAfkZY4mnUQIMfpQWK6XL/jHTjv5rib64xvNu/EbJklWS2cw4co2CThl
cRpcud+DmCEDbVN/mB8/dCTwc+uPPWJl87hMZneIt5DITu0D7hlO28e+kZSQIG7r1UsBs+YVkxAx
alHykU4rnngmRJJekOO09nZRBP3lmULyI/cOcIhNP/la299wElNOFG5nj/rn+oxHecaXLIGPN/Oh
DpyCLek/W9lXo/tF7wzqWSUBNHmIZiXcBdVc5lb+5dcR83wnpvvpYlU5VDL+/Q4dnD+uP6+NpGps
SQIi/Lyjl7UL4B8YM5p09zOuL2jX/PyeYbqe4IhngsHfQ+UDsWMYlq3NgTU=
`pragma protect end_protected

// 
