/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
bc4WnAkqx6dlMsl5fn3cAprcqqxHUHgVY/ImIQQum+cRAB7ouhGGGf7iFZf77q22uZ5IUqV83Quw
Hyk2hoLyHV1tsHXgJxRTk+FG0z8kNO9UiseME5aOM/+f1fcoxpdwoF5Nb9O6O9ouJZW/9wU+cOBn
deDxs8Fe2cl/gc7w+7aUoFn4WojygKnIaeby9NCvgShnH90A/5GxWomjUdPAdBRy04fmF471qpG3
rcDSX8G6arFIKQEh5UwVCLxQIuBK6e0cztUh2ocE1tgu0ybaWCTYOjp5wNkYHxW0TxCBiXthO/Y0
21pIqRWTmcspQgDYTjUBBMfo4xnplJBqhrkXZQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="ASJKkguRF7cNZtn0GfYOwaRh6RbIlcvsA1oAuucVfb8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 992)
`pragma protect data_block
Xy3DKr6jQ6T4G9Vc1bujRmksSbyKrAHqxljLVpr2AqnA48rS5l64C2d5VTvu/WqjYINVcCbrEZMB
YvUaPSPWMNz8kJT/2pPyGcEs/pSLilb6PWYxTxCDh8baHuHG8IQ0+zeObSjkmJr89Uc9XpHXZXRt
Shwt8BPcYLfTZ700qAFVZq+c1s6sPflc+XTgATiid8A4qTMqoo0NT/NhSgGeNXJGjlsmkJZtSyq4
SYsXq/jGp6bZ7agshXCzRuclRv5D8SljJU/f+QTTGm7P5HvamKd8XzzofLqcJpuBGc8PWefKVAP0
MZQWancPwM20q2aHmJqlX75rsbI1uScd9QdXUlz3265S92+W3cfl9YaXmjYsb+XcbxfXeYxfRO+3
wP/yOq66FlpggKxBTP+yjSBrv4c8biJgV533uc4MWhU6e8ZqR3jRNL1Vy5PUrielGGUvv+69IJzK
w2EJJsP60qhHdTVOiwpnjgT2oEML/Ba9B6Ohsfl5dyfWgCvWeI9IZgZzQVQtWGEfQFy1ySU1JhXZ
CzM0X1god5tv7GSR2MkihMNvqxPZA30i4/rycG+5LYJNjGAlFF/Hiupgdv/TJ9RfigrxLEoahQAH
gYpR19r2PtMHynDqYV/7OZM5IvNMkSnwOoqAw5kPcwRMqnF9lt4swGFw2k8LNVmUYgyaJXexcclc
A3TEt5WbXlwj7TgrupOFBsKsEJ2H4xub2QBo/rAyn7ScbELQplFc8OtOmF5ZPF/MoLyaNaN2P6E+
8WGh+vT1CtG2fgEON2Zo/xAaOXrVqbAjahip932F77okYZGS8Pq4U7h9gbe3m1Gq73ATH7iNYL0G
DZAQ3fhtRa3piVlumQW5SLCOGv5AoF5eTZO5ATEJgY12tNe4EODwjgqRsIieTXdwDtkuE8lkSJtM
iapB4qnVU8B/RrgT9qRmPPGGP/wM6m0oz4fWkoOqN+SZaI0/8+WLpfPgq3nrD6X1SxlatKqhA7CU
K6emEI+0AyaezvpFp8lFmeFKRbgQMznplFQx4Rnrv3+PWgyC/8gKUFktXddrJvFj5w0d8mD1wptX
cOpFE9nsf3aCbSZArQZ3p8p7L2nsUJqTrG/uM1ZwhyVjwQWoFHF7Pv+1kqKon51Rgr8mcva/+yi4
DPxGLssC4GJo7gKycPNjwuQjESFryyj7topxnT7nvSCQzuTEhXBDP9WEF7uxJzpzXbzAiumEkkHs
5nsoCn7a4EaQNZCf48LoPuYPgzoL5QgaXCzXpIJv8DdgqJ/9XYBpFzli+pl9QU1uiBwipl+6bBFC
be1lkWebYvLrN9JDa1iwr/ZOZQ28eLs=
`pragma protect end_protected

// 
