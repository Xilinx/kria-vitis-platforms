/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dD6sJjMckNM/hk590wWgo7QyLBP7qvuv1GnV/mfQB0w/i/pvS4BJcnppdBuizaQbHZTE85H6pboO
mTjEC8kS1yUyaRKX4KpOmRsaXVL7/iV6Mc+EyHoad/3cx2lAwTCRu6nptqi96Q/dtiPbQirlE0cr
bj2VslWvQXYp7agPImHpkldpbIx4OKKY49/lmZgzjQmz1uAl0Vpqn03TZsorFhKrWNa1NL2PWEvy
H6r6Q2NnxwJibsxIu7/DaDQZ9tx7P3Ox5rT/+t7OV/sWKJMNsqkendhSkyxMCR6Z1Ip9YxyEItGS
Bld1ucslP9zp60t9CzMGZcj/WZZ+ve1NzjV/uw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="NlHs8opBWv2KH1hFnLsdY2EH/Cy8LVzvJ0P9w8zUaYI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57840)
`pragma protect data_block
jOrE4515xgbASXSOIDgmJoLAtk/g59085Q1NX+alZrvKwESdWd/HvQY+Goe1eZkKJPrxZnkXYVeG
kqPdbXo62CMZ4JWPXZvuN0Kl3xE0GUTeexuiKf3FoZ+dcCaI3wL137czbjknojzYqKLS0WvSV1+5
6J2EHnpWjrfmxVYhiqqMhou4lzyOOp9xXA/RXa344TddkqrpDP/Y+MgffXNuyr8eCgGXl+u2L3qy
Azsoo5AoNaP0nf0Aa8r7uPpX2cq3sFrs+M5K4GUSrD0VGltfjcMJChMQcOUx5nySreE+PLeDyCDt
Rm6XC6UqyFL3tE56LklPgvIgGkB9zQRZfBFHCULzHFmXAskmVoynINJr5bsvtsMN0B2s7yjnEmb2
vwToEkv4rkiJfC3+G+Z2JaxAukK1VF8817TIjBlsvz9vSFGktLpk7bz8PBqDEcZhy57++dcMqJIN
26Dv/UhGoG6De9Z78GTrKt/DyyhlZlfyaggADm95r/hREJFuP94Xj2kECVLx62lJmg5RrurbVfNV
9q+eclgXbKdnDDrFFQH6XJ78J+v+LRo+23ytc93xP3PtWhlin5+Uk1DyWO3hFTPXGoIPemgyv2KL
CtvAAC1rqRL4iDbW4deZPywb+WT51+wPMjzjgxKJiENTw5D1D4s+qXN1MgsKqZ4gvnp+XhsuhffV
qPZcrPcUp7FuXB+Wl5vUArglOvLCFl1auPtGlwPALQ1hDYFjJ4k8k0nO7MFxccD8ajW5hSbkSSex
4Of2sM9wM4AJxjh3zCB42nlNhaygwvOdWZ/c+waIahkiJBCtABxn1Vgwnrr/9xz0IG7xWbeze8a5
RUpeMVTzMFrSh/qJq2QCPjsUBY/YrYUsIiAXWedEUHMsJdF5bzc2yZo+4NjLcv8cACeOr1k8UcKn
THv7TX2HRDXUUNr4qZ5dEttbc0iwJMqSNSDaFNzwY9xAG5ketFA8gOeiZ/w1EufdvNhPWwX4lcGF
Z6w4fGj2KGwYfxX3m9R89LkbmA3NsE9BR+cTQg+DVZbvgcjpj09UO6bqlfsVU0ERKz8jVW+PkcnJ
nou3f0qQHQYv89P8ZMCm5jxeJK0TtSJq0S5FAYiW2jcEFAz/0ErtN8OuT4SjD1/eIDzzWYKxItJo
sqq/DK88mZtrdirAmNe5WWIoc0yS5byHajGVC+2rmaC2uNYaY2xnK01wR+UvSPMgmUAdhmd6D6X+
iB+cUL5p5m3r1+ysZW7cjPNYV1GBnl6ArKvIjfUtUUVrwxQzKi5f+L9IY+Da+lXoYcCfTs32o1fB
X6BoUq1j2tc2lyvzf08sAn5LbNvoIT5bkD82lfQVxTUBKyDRa/1WmxWaZ1OIrgHIdDdCq+n8e/4e
MbiYfSg+ANSnp+3d4ZAtRrLRRF5PFj1B5r8OtW/Gs7+2TzfOthRqB6sOEYhGiZP/HHuFpAcOQ6kr
YqTId9nQJ+4M7urg9ugTS9B5hwB8M2elYXNzwMU5sPqFFcCFYroK9OfgHKtIMyVHWX2VRQikFwDi
nQg9BfD+74jTJDfahqD4kzA2bKr/uXaaObT+ppKpimWyMmYm9qnA9aTkh07cYp5InxqhhPFG/63d
SP3w1NybGDmlnYl8py37lrR+NAv/8yiyRXcShY0zgCWpkzk/X5RlsW/0dIs3jpBnaTlJK7YGu4XU
Rx+2xSxykJaJqy8e5Lops/PKUvTyyxnjGQTEyRqoNlufVQHoGa/4x/381zTX4tDuEWcaq+AqUiRN
C5/9ZN95U4WpxTSRuv3zvRrtYjR/orK0/ZjbKmqX27uwfcSo5UrDjKCer2NNFhpvvjZWulQ/nFme
9T+r72DUoVGNMj9w0Z8GhUOrOGdOqrX3GFfRubNEqtJIL1++VVcFafgidfBXspCFUhXOPOAhufC2
VBac+xRVK3ZvQiBUvKDMdv297ryWeEm4UDCnugrp8YiwyjWTPMvivBTGKzl9FN1W1owaKxpBFmJY
VnWeZIRHAOF3nB7bAAOXMm8Y982Ux79O+GywSMxAOlZu0AsGdo7KIMqw4Uk3fiIribW+W9+PCSlL
d/pgchAwJU5sPx35yLhuNXHfvf64G/U6r7lgmZ9nYDa8HSL9s0IiWezDV0V2FnspqwBJE6F783AH
WLfVhDcbxAMymsjakrjykR0h/5FUaGqzsU4SkFPo/0Lzr0ltWdmL1cZfvt8aaG7CLWCfbvRexW1U
mLW9ypUGnOZ+lvigCT1L8MDgXZXxuC3lDb5nIzkJB3CQZmUNg4sV70pGf7NKox4zpRbwbNfCNqh/
5W8URKpmzjeT/lrMwN60Se2D5LPTtvx4QYyus6pzi9XJY217eD2BQCZQDFxgQq6UaQcVfOzECVon
YptziPzn8q2phaql/dcnUqUMCOJHoyK07N2Nm3O/+h44a+wapykpPeD0YfG/o5m8D4aEWhhpF2bn
Uj0xhIWv4p/dZBeVcbTBGlWgO8ur/6zBygh5+5X9atmlkL0ATr5W6Aw6W6D3drLPDxN+0NVeAT4T
f0eDV/WP2fw2bzq+uKqAGa9zhH5t4MG9hlqJb5OyqmJRRbcBAh0ilLyNCcRwPiwAs21V8KjpXn6O
R7nvZ633HTIHZKHniAG3+H/2R6dZP2W1U1lt4bFGaiotx9SffdmQ35XDFrNKmiPu3H6hr5xXSqYq
2VFSR011OT6M2y/szRzA36ow1+k6XwKiu+CGb2OEAAy2t8xvwyIJ4PvFoSPlhUSDHux4MM92NY2e
guMXKQq1LtMu/vzVme24cAK+STIfKBF4iQiRKjjSxVxEuPkSXPTa0UMOh9YkYeF0G0r1mA5MEGnt
vb/GB1J8bXcseFI3hRmx+3hhG3qmw9ST41mBcEYQMlqvgQND48DF9LAZTDOPP2JWdTS/SAFxsKdY
YUQgFRahqrT+uwS1Kp2QlRbNRoJ6llzclexz2ibV8toHIB0SVvCc5Ml27dH6bEc75sklQltagvwS
XOAr1+iZAuTRGoOwuA5mHT7Rk+dRlFDIOdYAMuggB8u+bfyhKiKnXgPLmom2OQ4PhN2e0q/5T2XU
w8KuE2oUlHpe5JiNZdDsgE0JjPsDSeEsQ10i6JRPGX8o+fJXuWKjHLBIhHNgx3r1hnkz/X6TG9hO
IViJSrYya7cRdLSxmAgsoJzmRGcjuEnNzgIQzivtZUJSEUn+fGzDpcduexR7glwcntiwCNDSHq8U
HVXJxrdFU+zk0yTdx8/9X3jf4VqvSxaJA6OwXKTh+sA9p4NWvzkcQt2BW0E7vOjpGGYDT/rELvB8
eKzLV09u7YDJsytO9wqn4dra4AAW7Edc/K7009c2r3FNYHj/sXrWqOCUOKF/NTQa+ybwjK7vVeLq
7DqzC1BhH3z8uZ5VNYHc4kn9icQjaoYS/lOdJAABR5/76ZbElfA2uWIidb78+FiUFMLBPtbk4Rti
mBfrtfCjsBNssSyTE+7XNANwnm278D4lTDHgqzBBa9I+ujS8KG6f0KMgqRe5kqs15u4mQa0t0/Fy
lCdYzPjeX/I5x0S44QyjYUnSo2liBYg7m8CayaXUeo5thCFvCbXK88ati7ZY/BY1cgykedfRblmD
hvH7kk3ZnpgJpbPyZ7Ap9a8XAl7/X0nPnsBTeaWv5W3Q4mTvbmFi/qpFJINhNB5ugzTFEQWsRxk9
U2OIN1RGPTor1SekK34cIQMV5QmY0YZ/3WbJx+IH0t2d3KJnjkCTDwFkAMutgbEp3CVUEGnA6K8w
cKPGDh7vHVnOhy7Pc+3pMsLHWSI0gddgxJMuS7OEaUm1FHo9VBOM1u7/+edZ54E8cwORkCrMy8MU
zERLDpCPc5QpgiR/nSKEOO0ii6o9NOVlw9UKCFBnSuihibQzbjnN6/2GNqmDdUDXMYQGqJxjGHpN
uj0xfJm7M9ZnFlxPFwbBeyljzbNuAycBShAQu53YzEuVbFztQZJqXRAx5DlA9p0TJ2HCjN16HM2W
wOIa80pvhucy9QL6+EQLpdTVzLQv51PHu2sy71LlpoZe6odXKm5l0pdDcF83CSkyRtUjkp1+CX3U
zURmaK8X4WZhwZyo0osya1tgCuGtj+XYNmHVuYpcg90Nvm9j+wLN+xKJJNw+Xn35C5pKQ8xj5lzF
7XY351q6VIUdcqe06m/PM42cDuVJAH0StN6bWShuGS12cgnzPuDcXaAnQ21bggtZs1yLQtNVvsOt
9X6Fl/fl2LKJVeOOStYNsHwy/PAiqM6Gc0KtfvqNGF3zep7KBEd7+44linKiA3IMR12TxmHTGJm/
QfZMlfI80bL1PkJHHKLX0tBq6qnaKGw6wG/AW8b3Z9stIwF3LiwKfpXYS/ucEVRlbvb7sbcPWVPT
4yHZ1VqvWI6Yh3TIRuQ+NxM70K3ihff8l1+mQ7v/B9zN5odRp5uPWeVu55y+aF60kKyB2D81DtiA
XS+a/48zbT7Hr39Bfa9mh9PgPlalLocdzRM+ZjctkVpmVeSWoGyvKxruyqjFbT3i4b/8JSdv0iwy
lz6JP19mJFQmO+2WOOHL6t7dHeEKRXB434kETpG+S101oQObuiqCgVZt7z46TGicHd/kkmvyYKQA
CZ0bfM1gDbWiIDhl5VU90xUvs2ZhMnPPHb3aPLudXOGKouLaRrg5ke48fiU57Pluc6KTadUIjAFA
Npnw/JNB2KbeVjCCk7WrsLU1+iCSmi65J2yWmlk9hb88vnxFNCNN86+lfCidTrEOvIN1Fi5PmFTI
mjDb+sqAuZcQrnQlT66R3W/hRXwbibRGbOQK1MA7l6s6UoS16tI6+k/cuEqDqsWKH2jD6JVAbJEV
16ukQSLD2HRPgIN+vAuZptkYApdQHxkbfjeNqH2haCFYmPNRCbO5peg8UwolJBXvtIudg/jiynAY
Sk3wUsPfg8E26ZOB/+IysLuyUR9AS0xqSW3QZXGti3zftB+Ffx8MoZAqU92vOgCXlQhvl6eRbh9O
Tg9T6IEllX3+b5I6v1acOoI3doNDK6OXJ1v2sVY1rLnQ0qpMntxIvHJ0X9JmOgCJindxVfiqXNT0
NOmhQYnrcA2xth4jLQwkxV0hujHAFa3Yizd4Zz72QMktOmXETQCwXdVBSy90mvPmqTU1H/ZhsJS7
/qxQHjPDPZgvcebGjO67PeEBMXqHLhJaLq9isNyZ5SXSrnM1bE8W1dq8x1x1wMkilsR5vkulZCXl
OFm5s9Kk8N61w8u9pwERJKy+Gbxohs0dv1he7KF3TIreEuEXH467NeweA0xFUXcUrYdKlkcspfEb
RJ33+1jmj1ePHLScp2ZQmxxj2JKydmZFaxngQ053l4Gslxnd/ORI7RSSglRz/gtw+3stX6OK14th
F2vK0LKAqULDjjN5obXDZqtsNCEZsnDT+tCbK3w4ZeRyhHUqBNsI5kXaBnmFNP7SO5KzaIb3YGvq
JO7wlVMBn+Qo57xFf9MN5cwHyho85iVg2obKSfV7ZynRaZHiH69QxSsSAlCNk3Ze+8u53fQGci0l
z/PIS8sjoPMVN38EkLeBJYPrQrSN8APCOVcR2NDSo3Q8bgzBYYWApfeEQq7lVhKXnAeZcg+cOKs/
VJw49BMNyYik5skgejYtmKDCeHWGO6APqN9FaTMJN6c8mjVdJh8s331oIUqkbIG6rX5UoZjhceMJ
zn9jf6Ji7/ZOdBDcSG5wFsOTb/YgH71i1X9J16QPUsNj2cOP8DTcX/ovBdl0njLg7KRZCYflo8Dv
/Be1wT8DSu8fjP5OT/UFanJ4oZ6pUR8gf5WzD5SIo4LzGWE5//nOucSTbyYEgQzkQe+GkJ9F+7H6
ba1bVHt+YYBfRmc2vwH8C1TCKnc7FPOapENv0GzXfhiPgX/xrG5+QmvoooXh9Ki3KTlwT6H00UWm
jJB1mYYSzy/zZbZScU4tex2qAotk58JCQC1B3sJZHohv65lyskMdFKx5KWVwojdXFx5ev3q7FbRU
pXbFAp2IbrY2RiMj9GM7nMY9AS2ceyp+Yey6yRrKslzA6V/2R2A1O9/VqHfOPTZtc5EHUu5E+R0+
z49WmRVgpogkYj4PVqNtdNdhZjQz/8Y0hhggoMCseEA89u+yyyq5YNHB9pBOBxKF/bmD7/Pw+Ld2
bhf5kyZnPJshJXeN11rnPJpQat5dzWIn1FmhLLqhbczAZDA3CngJQA0Spgk233owGfq2eOA0oVbl
ccnkViKZm9I+i/t6p3YZ80GHSk2dwic76NeqQfMqh5hLdW2K32KC/Y0QlY/BRUz6drzg0mu8hMOc
RyZ4Fe7cmLIHUEdswCbFwsut7MOyIm8GATjoCui6Ai00uUhPszVVstlM+nV01k5JPQS8nfCG2lRL
qy3Q0jZLt5HbyCriOU0Rbfwm4dYdkDbABBMvZit/5QsNoZHX53zhZzOwMlrf89sdL+T4+HWU9IOp
I4udxC/fuFWTwlIEOzId+vN0in3lBlzcExwGNABulLNx7iFSgnQihAQy/7Abd+2RpCsUrr/PvlXj
Xkb+ZIGlKSr7hoH1dElk4ia8i+5fuSdsiuSBIV7kjaK5uB5p1VvaeOBgBuGwBSqe+lVx0GwOBF9u
UPcVnbl138KqOK/1Whg3iwdB7Bx+9f8zSTLd0UQazlJ11Zmx0dLMWQj97X8yumGF8GrCNEEJ1LKX
IFRu+eVi3K4zwBFu9ELTJLJE7fvankwO0VOIBcdou4ZK8rAAOSUbfIXUHYD5cYRVpbY4tbpdT9Ou
hH/J1xWjVuE90siwdAhfkGWuBAhHDKXACOhgAViaOhcZ2TEh3A64R8GOeFDPGdjRb2gByUMvQrES
EwgBrk04VHscRHK6FvpeSukZfITdOnduL86Ib+rDeCuN6Mp/RjCTEsDwpeki1pOVDqbl8pXWOjbt
UH/OxFgWISdvM+S3n/JTqsQycDbM5bosPIvRDwwekiw7za0dsotS1OQi4kTI+W2MTJJLWjCeJqs0
Qrk6ZK7R+iz9Et+Y3CiTi86zhfYlTTWCAPiSB2TuU3WJrYqES1NZaxtI3tNGs4u/RuPDFOe2SoIQ
mZvUshMqae8SnRdhIlc8R2Xp7XAH/zh3ejTdTVLtHjaRSC1pwSn5SQAl1MKs9ECalPaMWOT0XxtN
05StmYwJvnRS+GzZWS6kAcCoMgVZ1KhpxxRiodD94jjkCvH5tEjS/ubtRwhyDZSGjgsdyP935eR4
v3eWsdPF/ufumzkSq9sYyHvNccb3168G/Wls9l1nxt7rTi+6FUNfK3A0aSFlzTS4VWuKfsBUoweb
4o3GT1FQVml0RkOUCKpmWxJlAQsyunkiMQFKb4jzFlmXMRHyJysdB0l6TxYfADzVn5GXFZfMOBfD
/BEQGy6iC4QgNo5ufOkUTj+26r5dNe5wGi+XSD1LGxr3gCijc52eW/zeRJffEUIiSD2zUR5uC1Dn
+8SAxgXsA32XqWSvbveH+G80XOONBD6iB1HLPbRgys5kOpU42a4o7jFFU7j5OmMl/npBdOk8SN1/
9c819HdE+BfJrPKQ60p2AWeWg6l2UMWkimsfg6EQfdG+RzAojOyFe+8q8TMzWkJRjEFsQfg0OB2t
BEl0Z8GP2EKmoquxV5hFN/67/j1Np7BA7v248MSoDjgLp1Ju+MssnnlPAo0IJhoXdzgBmxbt3aXZ
5ey5ONZZY8fVqEZF1s0deSElappMo2eGADmGE8nHSMFYMV6WURconuyKp8WAGJmOunvsqbLJ5GKu
BPZfUEuiB5dtzDtlkDCedV0WvjLYGgSb6Q4/LHaU2zOYteFpp9hE4x8KL/Qzfoc2Clv749djcbVe
Mj8oesmYX3MeIf7a0tTLmDRExNGI0xPIjClHBFVhrVF8qwb+xrLPNcblGrBMOhhiQD11tSODpaVT
RsxdpGa0fnuhJcXf59gn2bWuUqQ6NvHTE/mDvCon2q0Kp1Nd4CU8s1BJNFyIqotshYN6Fv5qURQs
bISOuZWkOM9B6KLOmXl5n0xkVdFZXRWh/VveGDKiWFoxqOO//sNwaOUbtNmw1nS+IuvobsY/7M9g
T4+QK3VuE2PySZkgXLBPwKQgwTaD7PmzC3tiJtx7HIwIRmM+HrQUCP5tpvqIJv32vULpX/xrmeDL
grilNUCxuf8srJa9Bkxt2tqRnOeESd7J5WEvX9A0IfytkJZthdLov8cKGEd/Nv1rFzh1VG5WyBwG
t3kfo3RxTw8RHCAPWISXAzag6w9n8zSFbySbkxlGva3BDnjzP6bVOXx1c9DdpRdknV1N89F+Enu8
j4wvzhoRr6Kz7VI0RfGucysNgdbHV58me089Zw54Pp568uXSH93bQa57LRPm/hL9nj2nCBn8u1J7
vstyLi9lvBiml7qBNtTUk5KU6bGh00/AFOpF+Su6qkUY3Vs9KJybYBgADipNjE8r3F1PJ5tRJdRh
GFNRzLgZlQwVn8aiOWeguEoIxrhp0F3ExZE8NE2qC68ewYiWdy95vff4vQdGJseLm7FsjxvMwnrs
7NftAgB/mcVIlZBAHCcCAU6OIzqQyerKD6g9IG1Yxi3/yP6UPodWu52ja7J6u33YEf2niLvq15Ky
Zu4nXhtwmrXgQtsAo8EgCib928K1eFCPdqVc8SRAS/3T2xBUpZaB73LcvSoVKLwBztfsXrE3HLnx
khr3IeojhLzMRYDnCBmR7Dq6Hw+ZWAr5PM4jXUCoa+Kl5eMRBr6TFC33PZtrM4GiPs35Qms7YRDW
XggrrE2z9XfJv44KJGu/t5dNG6+sFE3/pOcQLSPl3keMqTZnW5z5Z2dCDv0gZwZoQIEXYxnSRC8/
AzUIWJz1AGsMFvucIU907poJeNB03+/VRFTk853dhI3mz1uxjaMRLtSkNYUbCJBJeRgvrFbrRfJH
p6kwIoPkB4k3tA4Xr+kvVlOh3899zCcbuHY4zoceMUauuhuJtQd26oGH4miyT82TDAwRxcoh/x58
YJozTXAFFlnGOM+oj0uTfsKRWaIjpl8uayMxV5KZhfGMbpAgTChUlnswzsZHRGphF7XyRlO0MjBG
sQVQ4IZC6RGBKVFfxiVfSxhgWh7wILWId8wm1DZfIOefD574d+PLFuFwOG1y+Wav5SZLqj/lPoX+
/MvMiXnHyYTLUHF4/66l3+L2Ouc7N7t7wtJTDTyORT8OVTy9H0UVmVT0MtgD8f80OGm4bysEnQ1E
+aNOeCTqLTdTwR4/8l7uY6oS8gCCPedxxH/EL+/T6ga9/ka4CRpmF0b8fVfzMo4Zovl24fQki4q4
LGVFK9A+nvvFLpJvzpzJ4FEYv6tDU9qgS2boVKzEzSGhbHh/OLnNdkPOJf+eDKUJtbztbbYQa60m
ejFflH7itYDMggMrx1vnOjBQ2xPPHCDw7TpwYCDpjmJ8CWR3JpmqdpzqQuZNaglbW6O/6sSlwLMK
vKbnui0fAMX3uzgPMUzWZQBlysirpNtOARVJo2ee00X1m9gzobMb83pGETH5hWaqgUFa+vq1siVt
KskYr6g4jFsA+vPvMT+zdlgLbRQvrAPPbiWxlVKfr1mlcJWV/Hs3jG/gK06zWhzzWWSBz07uFI2o
aQER2LrOfvRI0a9BGebRR2iSU3FFf1UdFvc/93GLZiZa95mwqs39lk0hE+EfFimp6zaI9J+E0e5g
G251TXsNrQuxCddq2RcBlg5W2nPxdZNxeq3JffkwrAyiX9FSQGj4QH1DrJ/K2VEmO+AW3O8SFcjo
Zk3E1XZpnMNrWMhlzh2ioMFM9ZoG0SPdoIOayb7lB+aOcwZwpTPnRXgcJli5MhnAJ9xtxchvgn0M
h5W2aHEwduQdOMTQTPXVKjT5tAGT1E4wBTRgilUnCVIzmxg1T/BmlzScIhL1C5CLNnrnqH2S097E
Nx+N2RQABqkYUNznFYcKP8DxezT7eW7h2gpr8GLYS5HJ28tWn6UtYurm+Cqb42qQWECQk7bdPq9V
1aTby6UFlp0WsWmIzey9u6n9jw2/1lpgxm/fjEjoWWTrfeM1dH7qBsAgUMOkeMc5q6jGL3/cYibn
QiLUpLtPxwwjlzpZGv3eENQvrXMrNj21JSaLOXde02yrZlxo87at5WNNSTFu7kFuKwsSR6ifzF/I
73QoLfawYtuyYL7SlC+IXU15UjECnhHhuq1yHJn6xkIMrCssaO8dQeCPkFMT4naCo+5cJ2KRFcPU
ultXPBijQkTVQHboqLZ+2R6y+iADiV3qqsGhchyVGjw1jS5dPhkebTytGziqIhBX6pGGY3JdW1qz
SppIl+kFDy3Ow4ElTrmzAB/BJKSNDO9TbF4YeZd7DVjf9kf8cG8gwYpm1fgjVj0h19CnPZsYaDih
Qos3/CTv4Ye0PDufnsMgg1YVs5IYBzMnZK505/0jRogsBbhsy//8viFZBtw7lJxsaJpscyYp0Nrr
9wb4U2tmHguM5sFz3IU53qEIRZ+BrdR/j14NH8ISq0vlQzteYnm+t1vMS7fGn96ywjgiBLbyCL0o
jUZhd6bGLmug/SMR5qO2EaOdCL6zyu4Sm2t5C30Kkwwwbf3MkdnoVx9ZNU/rQV0YG9pBqUdEQH7T
+pN/ilhddweCoNRVWuSrIXUdv8rpawWJeNjO5RmCb3gkZfLSSE/bsV/GHOGHlMgADwVkfPmEsiC1
7JFONZ0g0XUof8s1zblsS7UYoQ6jQZiiaUyoNLEZKXkkqXHAo87OIsQp2JGjVHplcyT3edZkPtDK
/lCWXl6CNXbgz766IDbx/uDI4kX8NhO7eP2JT2Cy3e81L/ZvX2WGxXi+9c2DsAL2ytzomHaygsKl
BH6sHbsyFibxq6Bzax2a8gq2Ytp55DCyipOfkMHUz+cxNxnpqDW99OV3nBS8ZPDTt/B+AWN5EbOC
CCeX2JtQ75wApZNZ+FosgOYkcv/KQD+ECU5P1T8uLqVsCk+pcmIK00HRnWRaXS/dgKmBkyqkOWkA
/hxBbxuAD6/FzvlA/1QKFH3UunmOfSpW6LRQmUFbBl78jWngu7DdOG+HL2F74CI4gyw+lYfh1l8k
1OS1BDxQdYEsz7Idu8uCEcWtTp81gPmV4f6+TivLi95Gc0s2Ro30QhvWIoIjtMUwPFrC40j3SQEh
k2IhHWTlbffWSQf+5mEIAiWsuxFLYmOMmzR4vfKt2btyExfiCt/1fUNhozwZqsf34RPTx4xW16ku
6qjLn939AJy9rZ0LV8tUi8zjy2GpqaPJWfKhXq0SptS8pGeBswhYwQYM/q3htbvwZbBCY4k38wtD
3yGlCGO/4KPZQ+0a976xIJt7q3Wo5eK42aIfzVrRpTzFNYLtduXg/TB/bJA/UZud04nC162l520V
I45qlWgwCt8477LsMgS5Uxz718Hn/mEUrv2q3yM4X1s3GLlKOWevINaZc5GxDbzXDjf9+icVyYhg
U54BAL5bEEC759mSKfQaqR2flKEpKsapKZfW6yfRWGOEZEZeW0W4+nJfCX/PGIfKhxGPphJ1h4Q/
eKy8H7fDoqHKazPNCxNS3S3LQ0rltAevZTsy9CyHw/Uch7z324n6aZWRcyYu6QhXK5YMlik6MbfC
8Uxx8P9k58vPMSUP77RbeTKlSswc4TA62GRQlXSO5TF178d2/RwcPIURLhOMEBS/xM+ahlh2RXUY
L8ucMiX28Hdf7FNZClr73u7aVJ2vWPdFhfBku4JuiT1TmVrzF1oDnOCX07UPaeZPZB6NBqrwnCTj
lAc78HUVI8HUOvcFwpJdQ8fFhnZeKo1lzlcFu4nHvvpjZVeOuzd21fSoZXypxXvGQVoTf7uWvCqJ
TLnjsVV2NcE1vfoMgPovWIXEPx0jzBVdXhZqAnjuu8c2hM2/A1/4AZEuvSOs5C9mPfmdOLnbepIY
7lZMn7pvNqjgdISHslPo6OGiMbNaI3U6OsomuCNEmcTpOdo3lZtQLQp5S5G1HBlcL4gO7HWn2P0H
rvGGDiVPt0jfSLZTSd0XQJasZA/wcAa5GTlDkWf8Ret9DtR8zGZIY5Y6QH6yqBJIyYxfDsL3RTIR
REh5N6G2RBVkUSycjhkTwWlVpiP7cWpkdZIA62FfnYOnEVGV1X+1sKpM0fonR91u/BIfHUk2Rk4B
FxgfsG1zfBPBah80Gx3WPQWCZk2p4y5Ji+7UEIhPlZP69/6bX2SH4HOw1J3WtqJhjLWXLaAP2VMi
Ox2KFDAc4pFPaspWLVRtCH6wP4QexQSg66ClpoMCf08iuBZRk6YNOa26roFLu5kYefNwbS0jGyFD
+DywjJR6W9+OFT7DccPzIPNpf5qZOcMDILtX3E1ZKTbz3yqEukIwt3s2YvtDQKq/hJ7M9ggR3IVI
jB3kebiX0TI8VjlBmTyIqoUOWgQcIFdy1W7Saa+zNoym7uA8nVaZB4EOM5q+s89oOxjPxhioTAIa
sWBanWg7RKWN20eoqKpmc0Ys1szyZ/+W2NBmWtcv/qtfkTtUc0fsh7M8f/0l8j64WJ0Ue/t2bD2R
zAQAbq+lb1JD9H2gobDlRbhkTm24LMHxDjvtK2xtXn1OxfpPfgN06g/QxAfg+jMFOjgo2DjVmR5G
BId+ORLpX2OWlBFfP8A+hko9BupBpT0yqIQEu1sWFo6SobIk4kmGYQa7WXTP6iCTkW8ZEZnXeh6h
OtycQlhM4F6IinZrbcBwHOM/Cm2Fb+Hk/qN/HJx83qpLXXQHzV6KRG+TAiEHHbQ/OJzzIY2M7uBh
FLnCmAcl/s1AFJnGnL1kKFzdbfitrsb8H+1I+XivBdMYae7XMRoDjIdnpw0ENnuUp9Jk/+ugr+lG
Rn/R5ClR0+gNPVPLRUV5C839DNg/N8i31L8g9UPRZO8OVo6MMS2cRBFQgdMOvQyZthJ2jCyqIFg4
x7EoXj8mjWuc59EhbkTX4CFHBC99UB3Akj1VqXcBGJuYu1g1eYyNxGA+bL2xDuSwRNbrC/L50meL
gECj4vx47UY28oLE9qyrTa0e6Wr3imiszckbxA5S/voziSlzYpemDp2fjcpP4rzi60PCYPhn7ud0
kIxXNMxqqxWEFmq9PKmsCcqRAc+ynUwx30hkfe6zrc0AftEnjBB2jXDusbE94OjNLc1FGqZYUzMo
FilP+6+0g4WjHNEjGMKzeTzg4vwAAoqesiDaskaXFCtcUELN/CFLfeVdqpsOmFZ/jSIOxjcMHRU7
ExrXvVdeog+gOMkA+EwaT4YM8Ee09dGk+N3jycEwhTcivMMrbxtS9Sav4NbYIER1sFZ3++oVSgIV
8G8Fjh3NEgMGMWknV7pV2dg6aXAIVq8i71wb0oTUypCyh4k1+uxC9xUV8/M9DW8C1sKKZEm09CXN
ClCHQChxNc022MIlgiEvgzvvmd88KZZg7tR4KseoegYSj3TcT9o6oHrT3BrSdgQxDB8BGMvw7lyP
y9rNLzSaj/tLHRstHHPtxSdgtfTwz1gqIb4LhyU/fpOomih3rO9i0ukfWN8SHcMRXDMS8XBkHEC9
42g8T+J0sxcwoaCpvIodIUGvNJSMuERSxJ7bqSNAheOZCdxYjSv7pZ9FEQ0bPBhSU7EHIGm+6iP2
aDNT9Wz7B0P61bzAUxRhy9j6cOiLz+b5Zu4vNkExGwGl3pNVjy5DpasjgviQh20TCqefD7pTUtyX
ZMS7kzPIbMoYM3Jba08SSFTcKL/jLJiIIGA8qWdc3xkGJzxIXFqAOrZx38zdc5+CSJfPu1xCj3mi
0/iHdRTE5qiPW1TIdWSQWCMyt5RNcZVaORuEhwfHnvWxil0vPw3MvuhzAjUBB19ocGIJ9m1xLWdl
xyewfZL090bLd8Ux6iMtgn+La9TRK0eISz128tDXujyKkjj3A0XWavPvIk2lK1YemHGcsmwtVa9U
YUr3fT1xs3adyPuEx4+c+lpmEWT9ZpzTi/LKcFNpM8insq+PYpCc1pkCt3qFEem5u9lKvzAlIkLj
ulCd4jjua+haDk2LF01ESe5677/Qd/B+jNkUvuGa+UfDLK0jHvO828zcHTD3xtpsFajJ9VusAexH
I1iv12yqvIPBV3j3IOXX1xgt9HiN/qle0N5GhIxl6BPf9FA3pvrHNpRLhauIj0gXGHz64PGG8XkV
tFwb0gAa7FlFDHYFXJn/TMh5ss7bhvvARcG4ErQYM9Hz6jIPyNZH1C2vta4KZyIgxsxGQas9mqY4
5KFtDKEsiD8fyoSY/UDb5gV55g5Rx06OnIsG2oUzOToDJ7r0SopdTHV56wbV4zQbXhBwIr5Q+lz0
Hcji4tb5pcUH9nCIMF+wEC0pmP2gI5OB0iUkxHT+Fek6BjaJ+qt8K73QcKw8GmtSytJINlEXz8cu
uRTZOBKr3wAXR+GWA9pfbgyeKqMZYOs7Fz6QNOiuFZqEjSf6Y8kFq9V4JMnMmPWfQbKq21m5qkFK
R90pI91dk36nfJyWGfrnvw+OP3y0kxMc52pKOXPGplxMeApOTtEQz4ERSpoHWFDo3UddVWPVyNS8
m3txjkBRkogCjlPymGR2B5r7Da6r0LhzJ3uQXEPUqjQLb8I3EaYYslXPprhIDgFTLSpyqJvyoSOn
2BJOGPw0xMZ6DS+gWmy9B4kJR7wQYhQ9T1J1ms3XsT30jzzD1OZB4rYrvx/iFH4cWZRshbl9zzFH
4zVXH6yItLQ07AyQp4V/npQRMPV+PKrNNywR/NyilWPxBvj14UnxvxSedfD7gEEUXS4eep7QRx01
XXgBcBjUHyYvnJgr31h3oQmuZBAi0ISS9U1iXHmFxuDmEoLU8l3UcIMlLaLhMC9wvM3mBX+TBGy9
u8fREOqKpLQjDholN8EJgeV8fzS56r0XQk21B776atKETGGjRsenxcTN89dBm/gGPl0UKrkGU26s
/pGantO6vMHdSiIUBI/+1EefsLp0vipxduRxTCWgD/nr+IXGEE25VPe1MPYJsVK9OnGnNl7d6nZG
OwkC9UXv6laDty6nz+laX2Sz2ymv2FCBNp+So5Ea5CGq0PS5+/koiUrfFL/uiyy0r43knqnw0Uz6
C6A/POGO/vFeDREKr81CvMz2zClVE0kjV7c35mffrGyutug+tz7aVHz5OlIdhASyGIYl/6J736o4
uywMebe3okdb/II5hCUJ1QI9IqCferU+d+aM9XekHHMhpHBWQJZqLPiHLTlfq4hkgs/boF/AmHv2
e/fjcu7DTcdly9d2fhg6229EDBQhCOpCsNIRyHhtpfUyKXNAlmSr3Da/LS2LNZ7NFAB71LBgLeXW
Dyr6Hbxyw8o0KQkNTFQcqz8O1QPkfDoiYVIJSHyKsUXessUeO6KSRlIrSyVoMTxbsANqSyiyCjkZ
ot79sxuKAJcUdvfftF7wMInPGfQfPJrmEKtwdyPsjmTWRoDyU+kj6+D/izMhsAOXq6d7u1ywOQVO
/XW3SiUKCT9YnZhX7HMu4Gy6axPZ5fURJsVt/5e1f4GPm6RYSbZP0gwvH9U/3H7z2rqS4LF2G4Ti
rp7uH3IOZWz8FY/22wd6Umw+wQJ+2svDHqstKPECYN9tjTdH1NVLclESl44US1Lp4sB5KY7a4XM0
qWq+/PMnh1QIyrb7xKP0t0m3/6w77UmG51fnh4wXKfAl2Ln0Op84kxx5pPMWNs+5qY4djk0Q4ivb
TkL+0H+QVWLYriuWYKoUsy+Tn+w9aMG/rv92bNjE6paew2Qr0pPYjyfnAFo9uS+AX2ISXYcweux2
ym/EB0zUJcFJkT35AG9DeFWgMefDl8NKIWAoTKidPJjxU3irVGNDZFZwDL+c+tY8evVslz1wTceg
lVaQTjLQsIbknNGbTT2brt2jN4QLhgJxR9NA80jDs7yqPli7Ebn+SemeoN1V3NjrMTat/2uSyT4x
KUt/HFowrvP+FQiqMDXwaGYTXAcrnH+An6f4lTeazXBDkoUKPzkn70+EeLfw6MDn7TwThYpeKBwB
VKHDGj5ufNWZ2P8AwwafZ0H7aAcD+DvUOlnMp+hOdAJTMGiJ9chBTvYtBsRbpK8z/1IjM73lQDY3
XhZE8RIEUZhQb4tCsfDQj2DsVvUWqglwa2WEpt/UUEPX4xxFQ0tZqN0pgYZDDDFJrNvwMSCxPwf/
iqy3+1F2pems+ZiBRCtErtvw2KCAFGZEZDpT+YIINLsGtZbZOfc65g8no4uuZwzSq/OJuyTAtcRh
7e7czgzL4CLPhrh5sIjAAaoQsJkCCt8FRKKlo1eKqKY9GPMdXGUVDEW3h/1I46vA6T7B613hp29C
JLrrD1UD+HsZJjWyeOlunPldXpC+IkOdOwgqtkfsLnYkWTvXFTaVEtSOZu8CRauyb3KVPOxeEsaO
9UPQOXC/J0fITnUSFnooFq5sDIdh2xY9T3iZEtfSFQo5hnmXVz++z4uZfGZeaoF6P2ir+vmoVnLO
4FKNsfH/EE6rKdzqv4qi8vjRGR2+uAd+Rejd1cjtNrbIWG/0ZbRgldhmKDUfymJhbEEfy2pIhwYu
S/kE3SdvT/oZjah3Qg0REEHYkGxhhYQpHhfgKMjrw+Sb/y5lsGm95LvwfCfrmf8as9Bm5ElHnG0K
62u+mtuKQ8AcW87N5A1cNfoGEjdMb8bBQhVS/QHB4xfXuoODSVDG46RkYTYpoMNsPzlpN0/ufTYy
fLmMnHSpZSBlrOXd6vDuQgcHK30tgFDFvSh1rU1oFR7hB2sx/4Wxa90HOkot5pvNAW2Co1chErtM
gyN/iWOTvl+SsSpbiTbW5MTfQhnYiyV5r6aVzkVYOJ+0yRTP5P9keDiJU1UANRbq7iAyb3GaTx5f
Pj1CYvnDizOUhK8+PxbhpFy8rmqqVNWW3Pi3YPVQJ/KcmVSFe3XUaaELFKQ8f9vnhZk/rIO9MFRW
gfSD6TYlDa/LOtrSKcnvVW/YScKguC3/fVNQ+RFFKC9SIgN+HGK5jnyRwHV7MwlMYkRsHNBjyk/p
2aoE2AIAqAE/4v9itWIvyxg6oXYluvRrBnUTpxa6T+AVcgMv5i2CPubsjhdggMl5adIm7z/drRa3
s+pf3o8Uf7u4bHWZxPoMoh7mw7PyRB9W3/4YSj/4h/LSlnzy8A2zUnB4NfHNf24DEcyapAgHkZJY
m/6IjOwHpwD0XosXWwL24xZmBqhA7LwXIDsLTVV0pAIMeYAMMUHyC5iObhMjJ3xG9C2h+FG6cVWS
s43rGwkYejHrZj51/rilNTOlMmdbNNKTUNtpuJvfGTIPEpviq58r4FyYHPyaaNsBLIe5px2VC5DR
4KZYC7p7iC5SzXQOYRgohKWLg0Ol3VHstW+QukO51yLPxzGR2irnVSuAb7RK7/pSYMLJjT6Pgsz/
/1cIEVR2ob9+ktRxyKM+dZKmJBHI0g6U5LGwEuTe/a/ruRbh2itXW0bNWUPkX4BbiBjUqvnMBPON
8CekBEccrdEGz0Ix9yRtSW+xedkj28wqhkamZnHGnClquzO6I75IdE0uk+7jY/GVJK2ZZuB6ZeU6
JRPtDg9gZVQqmvAufnaVoAJWmZbCXD59q9/Nn9GAmAVCNMmitZ9kOHGn/LniQ0osNrP5OTqVwz6l
eiGb+wLRWinm4kS6mt7qfdTxxFaWw/osh3/jRKKDFIySTPbjnSAg2BildDz+h2WO/BJbquw9Ld7l
lhJMgjQocwj6w8h2U/RvM2Kj03g0V4f5BgSUzy24jfJRsZC0CxhNpULlPFx/eIfOc3gTOH+PrORC
RomtkoI2soKI9sVg/BOfwXMkgJGktBk0PG8De98JxBVdBMD+G2Vq/KtwZWVaypVnsaHc4v/cZppY
SM4McwVBUdXWRtO5eEqMVPSpGlKyvB/rhtB7SUkCLycs0KHOb+O51Olqu2ylh2zPNWoI/hV4tceE
99A3i3neNSAgWnw8mjbm7JTGATYJ94oeuNlPo3II1l4DA/FtRw550ZG65napNvKb+5p6GDRLBooW
5/ABvNf6OCXqczJiYEjFsL4YhNZNK7Bvx961wKjH9qma11U8yVNp8sCBxcxbXUk0SwBTBsZYkdDK
Na6gG994Wdn0rZE9g09h6lxAnVGmpFhieqFXUBIlSJy9LIFq2N699XIpzXjKPyAKh4kT8NLUoP0l
GwRpMmO5lQBcE9plWVVgJ5QYzRVi9amnj1ZjFX9eAWP6PEOfIgTkBlaIjrszNKvgCiDQaHkp/4Ug
kAig+pmhEQr1haj8IITedI9UrXj32ZX9tfK2SKeBkJn5vsdXrFPYMBBt06KcdIRMPAzBh0aquzuH
QSENHU+YRxMvT4UNl8w9COQVJrJmXw6XFpbrdeOM/7mzGLuVzo1A88K9xTX4yEevndvvtikEFGBV
qy1GZQus9zMPiVDzNIkpgVSGRjMx9M/FPqzTiag5T1VEGvqxx38wnKziPQOwyF97Vlvi58vIRuRz
BHAmz1Zu0AuiG+24fGfhXQOOAMdIqE0xyOuflM7BFEAcdH3gGZRl9KVH6o6iFW/toyJlhUTDjjKk
YsfmPZmCTzkSX/rLiYU/NoSo/MLi5nG5lJHylGo40qhEMtWATgwOcKiG7fAS9GvnwW0P9SP5pA65
BPBdR5Xi7DZyscA4umFDe9BVxKE+S3rcKFR4X23PKqwFgufY30l+50eyU1KBdMqH4XpqG/u/pLtG
H1FTX+iyUp5uHgpiSifsQv/f+3j3731326iVR826EIZm50kRKhO/pKrbhgTT7n6cQqE9axExnlVy
o+WDAV67/sr7hIzB/UEUwwipzPTcYYr13zaueR1JGEppv2T0cA0zxmjEy9uvDyPOcb3Ar5imI3cB
pPHuO1pgfVsDdNwEOeZpgqW4a0VBqp+hxLhxzlUV0rKOhCzmlHpaB/hG84JOxnaxvVjVgJVgl3TW
hgXAPaIPVQDnY3SSoZIaNYXkKkVEaN5WibaLSg6j3QbeQFRZq3WE34ahfkX0DUV8WM5xrzIpB9p+
txm0RDnNZSjFGsB+K00J2ZTcL/brtfzLNPxWddoZW4aWdf0Q3qx7u9tttVOal1A4WbGsajKO1TxO
7GtZCbDwWbXmYeNhNrihTA66ClYsvD+R8VgozETcbGlil3Boua8mpcHlWHdleEYP3IC1JVDX1YDZ
XJVxXJGFeWxwV3CkEyvlSDlqHAEF6jA56ccOvsvoHMPx6vUeYYIPFG68vy0Dei9dqv/5zKjdn7FV
XMuUNk8a9ktfxk+stY86W8zR5miDO+m9khJiR8gSuqIcjUttkGTWlwhexYZYjDo2lV8/+JyB3f2T
ZehDYKjQOdwScBVd8dTepmucaEWS8md4xjUJCMXNSLPgNc3Cn7Y7YCUfveOMNGwAe9Lh8FvZPKo1
zg6tboIZTSHZiXfZ9b9bh4NTYDkz0BbZLEp6NvQzQM1mHtDCBsmxc1bQTsUAswISUDlExswuVMIu
QM7vMt7Rx8iz2FSN2eb4JMMsx/5u0E8AzdqFb4duUZAnHEwBb4ODlN+lDTTE6LsRPRq1SO4xM9fQ
MkDPhKI0zW1aQZ9OR8xARIiMhSHBAeqME0z3szi+l8r9yWB70lYgmHK0Fo74O0zCpgLj3OuUojsg
eDAyzNgSML3GbvyCJ/n6Nz1XO5Z4+AMKMJdKahvMZwNId+GIoJsqwg9zpkCKu8jLRzIMOAKbolK8
NnPDJFRfn/ly1NlEbBW3r37uj3AV87fC9pIcybF+WquGXMDB4VC9O5qe06CqbZNjUJY0GpeBVaTU
E1kUIzDx/INX1LZPgNhQBywWrUPdBPszWN5Hk59xdyDX/LJE7P+KQwWxi+lr+hqabmc2YH3DQGMb
shjHnlbDwZhrhBnoXgnG4K2+5cDknmRNtmw8EoWgPTM928PhrIBcI0JbzEGBdDuhieNoY8LPa1/t
JNIrhvaK6BLHfgtey4d5aFT2aIalMrxQAisN/wCbZxkXcf4A1fPufD0iptNm9Yw8ygUllD2T8QHH
lvC8N5bawRAIuPtXXInBgMYKaxVYKnAMlYD2nbaOh4DoGQKvfGg2dSoA2X+ESfb7NQ698vqzeHjD
LFqy+K9L2ImXr7XxVUmFw/1NRJwgvZP/qSTCuWZV9cMnB6aIwokqlI3f9Z1DuUqyTXlI3ceCKHzJ
BduubIcaRZOIjzBmMhkAORbBKao2Zk2XZ9gupN/ycaAMs3UqYCV7yL3pIyVD53ivDIsdVLAC681a
JAt9Q58HwakDzN0w4LSVI4/XUkHbIUfR+spZfGyLkTSMNvVF5Qp7aI9JQpLivWXKApbcsTDoIOB7
m2l2Mnb3uMdUrKPq6GtBgAp433AkB9e4QuDpNb6h09E2HbMlijSt1I+V4rtMeRf80UnvVV9HOBdB
7rcLA+E07F2WOpGU1GQ4aNB6ZPl4DlaUbBiijkiexTppoteIWtl+ohai2ODkXLJv8Zqm9RKKyHx1
nErr0pSPaJnwMg00OaL/w/dvP3zFssLS0l63aL3RgtgPu271LpKLueYtHuShtxlJHXHn4LBu0gbj
mxbi6/7GOu8+1nRjNL/HNP18231DPTdGShq3//dcyikyyFol6saZ2wz5TLiNaWuI4ArAcrHeJOen
MDfi0cpJh8JJHLHdcQL9g1zOTby4MAzt5kI04wz0ZLgQDtvS4gOZAKZ8/iACxhbgok593Ccc+3QO
gdBWByBH6rgbv7i73b0Y1j/MJivy83eVEDiGsmCzZnTkv1hWKCZOIDqHDHUcOqcpq/+Cis0rbUll
xI7pZrvbpnq4s2hieS8Om2WD9cKSqWvvcWGRrVF24Z78wWc6fPJq9Jhl4+MeFWbCOQRLYUhnv9eO
1KBYLrXhqfsip6CxJZbZS1tZ5KA9qEZVPEKPbjxqpfBogTmwctzJxrU2jRzdeViKWGuUFBsIrtjL
AvkCbfMofGwDUqBw7p38AqHKrMvSfqr0ui0T+A5NBETQBElyEMO+doIWlogSfTgZUzh246k+yR5y
W0rW9aNnSS5f6AY7hHbI1exwAfWclhUHrcAlyoYbyWKe1JgRGAk65KMH2OG7QlWvgSsX1lXzfdri
2LBgzg7nP+KhdbKMhhiGzSXqkTz9O+DDlMV5GZdGTbyusbO03ubP3Ms3lJeQ2sj47Qv+d1lUrp6/
cOgCzISilILQHznKPZ0ug22mMZstkbRz8VUqaviZN+q3vSOZf1bcMDJGwwy2LXvKWgL59UT3J1gm
9Ao8hQOSzDhXU+4NDJG329XUnvUtPWi/G3gxsssGFiwRhSQvqEcS6xuvqxeU046UR/jw2iWDusBn
yWcEBfOb4eTdQT2hT+ADSV0L06fFxgQYqr4DMZTTB/96puEIKrKLXlokepIRkOkNEOSXFgUVtj4J
NXwvWL051/PKra1wovUuLg8QyvemD3sQpnLRHNdyXR7CUHxjrs/OdLpq2wXZrE+l5fQKvixppWyn
49blWBe6Xar2yZZ074JTFAlbbdRNS1cX5Ev+iP2vAN5+8FvDe6R6YXB3VTrWnMOxbItHIDLCYNxO
chFPa+imJFW/fY8cOyNDsRI+F3ZBypr3czFR+H2Zh1ObDGengzC7mN5pm1ftB1jgYaF3lsZjzGEP
5ue/FzbXuEbao+/fWEvxc1Hsp1s1biQI+2cFNUXMGjlhu9efvMtfwpYKIsOhajexZH2sXQGe1PVr
RUi3cTGFYTOioCMM9Ur2nnccAwZmcnt3INBnKziAQ4wskDQ6DmmVf5Vuo5KzjAbnRt/4iadognvy
zBj1S7a5QZ9M/Yi8KgklB/gGYqKx0m9+56jGS9tnAfONVx3i6FzZ7uPuE9ZnAwt9paF01+NcGyhB
QDGiHClFAB1D38gZiaFgHfrrlHKcJCk6j91uX4kpfHHoACZMUFdKGT7Z6iMk7fREY4jgBP7e9wHz
vWA4ABcXEKaBl0QcIftaGdYLRJbjSC1H88srB92DUv17iAaCJ9v+8k47W1grFvXGOYPtOI7UaSK/
aDTM3JN42kIru/tFSMsaXxWOdHiWrr3FD2c8MXAd+gQ4JsWe+m+exi9C5PONjgxzP+IxAFvdCqiM
ad3SoRdKhl50WH06dsUUJI4clTpuQN/7zgke70JUR2ZGS1PrHOyinMGfkgYbgyhy6xs+rGybxk9K
erN5xB2b51aD+X+5Risxp1oxDy0BFd6zmkvyxEVgdfKFJAKmh4TddDuR7cHA4X7eS6Gzq+ymkUK3
vemh3Cu/FuCRLb7DrShJtpDhpYeg5vZhEqbkE8oTbUsvhloGGacuSkwK+qzQq2QjPIKSOXUGAHsS
ms3F3u9r+vnnR+ZZzuaerk5Ln9Yl6hS92LIxbR7cfyZB9eJ2tOegvwc1ck+K+kFSFhFqxG+Sd482
6DwLv+uc94tEAo2Ls8E1kbeYLmtLWSPw5gIPVU6NqGZreT6GEWM+dMQ965AQUvuoyF+AnK1ETRDD
sWiGV9xSWTCAd8Ckbw5RfNDl8zT0rE4V/2h6HYmFI/e6uNUlXuinH/tSh/iZ8Q5SHDc1CneCyUIw
hpfTuZgqDPLOK1uKKQ3XYG9T8Ak51q4CgynjS/UWXFtg2esxwNKbau8wSdh+9P8G1AW+RBZLpMnR
OF9LrsNH5JK/tXo+oDrE/NWrHs8Q/tm6Dwvlz/GGG1x585X4zceSoNCVnDhLEOPHZrUkppDk6GZ3
nIax/T10qaWG0V46CFsls2iMmOfCoLckh/0v3DoQsEg6VUEyqpaT1/bBzV2D6SfGU1DRkmmo8hey
c7oKxMQCnuKWI1UMHXCR5pwTOjqKeUx4RbmmER98kmUT12jZc/Rm1d0POpbFOGZ/y8XSRIe0RXDe
Np7vPYuyfKHJsW6GHsbvEkcqzOIDhlFj1i17c3vaMe1sqYQJLrC20UfDkjsfhS2/2btzbKf7a2wV
ypH91aj9YInNS82HyTzoUoXDN2H5LfcqJn9tQdqGfk0uaGXrCOgSMzLKtL2/KFag0MI95gt9Kg3v
87b2Pp/qwd46L0oyy2pGOVYcV9knucFvX+IdbO/8ZGQfP9ezfDdGyJoNsVtrYzxEj0bb7Buj1OjI
TpaNDOxla0K1T0HISS4gNgzhEemJyK59rR8om+diW8gI3tq/32aIjOSn7vNCIO2lzm+0BjXR9ZFp
dIJGl32R3LwMnTijkJvj9KG8GkMrIpGKbCyle7s+kW7EBDXDxUJ7H28eruihiHxFRAY2cVMoArOZ
xeaI6wxJ63i/MvBp5VA7/j03EJwuGzPCFkNaWBrowXyA2bLeg6/z841CAgMNUNSchcOiDMlBEkn3
X5x7ymFkXq5rigHsQP9a3LqSxT6MOeQmKBDCUlWef0RmqG6tIGKBWyH3Rxdf+f0iyAVCQ17+7kJY
MDT69JD/nB0+7J8DaT/AXRVAsSGPwy+y4r680GJssDpBgcWuUwSaROGbkoksb/N17NbriCmmzoKk
e+cP4Do6QZxRnlaYEwEI4gIggkIESmRdldg0iot/PafpoHarCpbiPmBBZHiUd8P4LnP/6xlSGQpU
tPTdidVktiZZu8MW8GprFC1+s+eZCgw9wsXtclShIXXx6vB4lMpefomZxmRdUih3nLaVJLWqU7kv
Eiu7jvuDowRHr4ptXGi8Pt9fNrJroOrIkELuq3n1jtdzg2wXemUI80ywr4sZj09aTWX9obeCrcs7
SMTL0n/0+srh8KhV88gjhdopobX2RSDndUXa28efNrqVKJ043EhaTgDl1EMm2qihhBWYdV5TVXD5
xF385+atzbdBquSMfDyKmJCeKCZkgK03W2HY9OzO2nxgnboZQrHP9ECLwTeTC3gXvHjncr8m4k9z
bHdCUyt9YD5d5wkr9fck/UnbaiHyMpLi/1fO3+pnEt6uUJoDotAhR9CDesRqXGguBiqEDeug/mR/
kfy8qrHG71YerS4iJcCi0SgnlY+Q8nnVqVTDLaC3GcGRRDYUjoBj+FwoAaDTRKv35psOvLLuA7qL
STcUmAYPOVqg1RDonV4D941UX4aBp9srDX13qt6gCW8+ax6iR4W4pLN+Ddiu33at8lwPv4ayL8hw
hk2XboG0INEfCGf0K0v7HzKipWsEj9Lho2v51S4dMydmpBzwaBx810BBhBkLf/8HPuCt6+ctxwXo
VANoYWnATzEnMhKZ95FoTc6gKwLc8l8o14kIp9BPtHVxlKD/Vulp11rESZdcNDcZKPuFyk7wuVsk
3SWmpoa20e7Bi70woK5ISquS1f1RNxMBNgUExwt+rEv63a1J3cpMLPC+2SnrDh7Vad1mjJ6giJAk
O7JEeBtC0oQoo/hOeiCNqP5mV3gZ0ivzSpuvdx+GdkeYVaiMYpvAnJU2Hi0sAuqptAD9elDMzQGh
+Nu0ZZpxZSulH2hDZ+dNLvCM6k0K5mjo39k1rDSt9haHl6joqwDwIFZpIz6rWg0eQANgCW2PX2K9
fwE/5/ZJvcjcLQvJmdO24TcgO6ZavhBeBkUzUhBaz7ptsc2pPqW5/vnDMVaZJmKrfxH0lrcVuU1I
nu/Hu/+sjzxo9HD2MsNQUfVJ12Y4VW/21qzIBMY3QZpTNmWn1XXjVAjlC3xNORyNrSk3q09lG9se
RzEdYkrFe/CNddf46FEmazXtHJC3D4dZ91GKiHVWU2TTGIsNkbfu0va/S66MXW9Q3CPlE3JHDA4G
MQlpu/WgxrmFvMGcjfW3MKyTMZAMjLhDdUQ/cwrhP6rl+31Tktc4mvGsFSdNseoupEBArV/4nHoW
L8yf1+NpP1qSi6XqTwBWfEcHSYTKayDrO4/ZB2/FVXtGlfD2pPiUEm3l9RSlTeB80c/dCatbueIu
Mo+G2ByKiUTZKkcdkSkKhqsdWEFErnraRr5E/L90fvydALu8rZN2YEvYqNbEOk1q5d3DrPZk90tr
i3DAzbBhFbb6/3c5/N6Ro0+z2uZwHhwZMFYaNqD86GJStkhafAwxSl+AwGDi1kmc9lc91gTvjGKb
i0CoVrw7qzFMesnFvuryqmbSHktgduROSHHW7IuNjCgryUKZZRau84Sap3imRCaoXPWF65LPGzzH
IVnVRCHpvBSJU333R2q7Izwb2j6ujiw2580vPXA9hNe6cjpQr3IlGiXXjb90axxl1fZTIuDu3D35
R3myX30vSiCNSv9sYmvAhusRBXN4WqOzQ0xDAujfqiC02PtwwFtV6C9RuBkPhIvdnd/oIlLDwXxx
+nYOg6Igrc0pHxvdlcWSc3PojSFcpWygYuBfQn5uFNre8yysn4MmUyEQszFBYD4W6f8g/BxS3O8q
ntrh8Q9gBsYZQHxYiYGWViD1S1VK/vDldHk3gn7cYdqMr2+mUfzSsUJ/OoAQ386pi9tlDc+I2eJg
ccjyR8WGLeT1bpFiWZY6JHyRVzF1ulgtcnJc7SO9InyIZzzzqE1NRtgda3gverShz9t6PhfLBi0K
hYU19DX5BCjsS3as5SN/+Y5iXHeuIympY3WgRnDF4T2MefKJti2AvNK7IC3WwpAO69rja+oKMt5t
xvwOAnjgrY73jtUQMSQA5APqlaPtxn+TG2wS54QCf40gAhmVTXSEWMEs93YqEevnLyoz5Hi1CuU3
iii5onVzSePtw6n2SLM9m4ANfp+YY5e5qqJ7GjaLUvogGCnOJCyfE1jIXAz0VtjL/7tii72y58K/
Nsf8qQ/u6u+4AezJtI8G0EQJ/Cfsha6vydCPNu5aD/kUOKOpLVUUO7O4/3BdpEO9Ic0fqxy97ZDb
LIvNe0RRaZyi+6IWCaOoTSPDXKqSXh+xVOv6mojmnkaobKYlHeTDzcwwjKLJPVd1SjqVJEA1EiKw
t1sIGi5qDEel45Z8v6CJkiiurpgxJ88hTS+3qWzbRosfUQNAh2dsWd0uBj+5Zhnlm68TYAyIo3FF
2z5gOOv+IVxNaIJQv9VYOWZh+z1kDl2oQE+BE6XH/PpaKZAoXusX4ak2PfDtuPi4HR6fbAfMYG2F
rRKsod6R6dYHexCBDgenXs2bbxiljHv5CpJ2ZSRnYL6qTvJqXBXVPUU941jOWyrVuldLnVY92RdU
W4sfQxv+9mxb30JjTB+jhxX1NmzxgfzZAmcNCzzboW06s5TG/gjTXhAsYi5Vgh8RMmtnTnmaEm56
4BlDe/WtsAbTxf32d5yk5qeHR4nnYH4Mzic3/hemyHCQCR4itGlfJ1BTO0/PwrhWwsDO1lYbxSRm
jt2rDCUmqG8p/tJTQFxQWPyq4hQ11PagtKtFVwCcDhtaOTCxt8R2QFtoxR8K845QcTYhwrTMFRK3
LohYdt4VyfDcbm4cJ4PSheGXyROkzwKYmQvOEXoNMe7M61m7JjIU4ihdgSGN1G6xLnKvxucyaYVD
rj17tadbY0OOYMWYjoTziXWNABgfSa86ePHRirybwIvZ7S2kUVp6gi+dZulVE8jQ18b++KtIrKsp
uCD3vGwYFjPKPvGT4HBcUj+3sF0nVIhlmLARSvoVr3x4cZ0DJZDJoOO2XAw7Mk7EDMMJZ4VdFd/J
LXVIO68RX40OjXpLtTPl1O7mrEeLyvd5u1qsMJw2ncfc32AvFgh/hdeRs5K0cdc4f08QGLkS37ix
1NGK0VCRed4yh5siDIZYLVhPjvL7hUpjN93TBtI2XVldmpgMOyje3V/zxM8K4QexhbIyUcF5r+Q+
oelqoG/CQr0JRPpe8P4aWknWBlvwtl9IMvP0dUmGxXJwAjMkx/x+xhXMfZe49Hh0BStdL/KiYHmZ
6VR1+Nqdv9rt7l6K2zmO2ESubWpOD4DtX/px1Q9/svst6A7KA00ESQn0sRm163jId85xn9Tu/dRo
hM31BuOPlbH+h15HD1anzQOvbZnv5lOtPCCtH4JFYW8CXWosRpy/+Lb/GylUojf1L7l7pWWtVVKy
yEjpJKR6m5VvmGLIFeTXPyM/czO3RCGtU76UdjU0unEUbkmyY3unTUVwNSLqmCNDpU/EZiA50IOK
TKK2+1GcJIcsNcqZqfLRg+ALWz94lsfGDe396lezJem8Q2ey6/17q8if+uL6JrzRnJJwW4ENjWNW
lHmPj+ngsUMeMtjTQ9q8DpD6hUuMPAmWJmNuG3b05WLBZQY09s96lfH4rTmTgZSUqK6jcvvj1oXO
G5593wDXfhwAN0atvXXRPR7Tf5RUNCK3UrQZQTG7UeNLBrXmEA1XuUynFB5un05kzanmXZG8NHCi
Y0k0RxM8Sl2DqlkIsJjC2Sui34aEYcU9pfKkJSvLia9NV5kSpweRB0n2QoYzQrai3wGl79GNcD3A
Kej8t4Eb2D/HvMPO1u8yKnDT2raGhxXBsvIJMgFHX2UHWlt1YiYrhrHACfxQuwOeJUoUyII0oaQb
KWikXrj4leaLkepSSraFjnoVQXpPVL93lqrdDZoBNSPDJf5I2KWL2o1d3VojkGTWyvNhBHsAQ9ub
Os0mCF61dTqzKlQUJEt/JkCMcJXoNusg8JPHq3LE9qMXXIHSh6QXzQq/6WAD9lYreuti+MqRTLzc
v1ToOYMLrXXjYInM6XsL0n2vQ5znOJpOsHIz8Hlz8qnv2bGJiWKmRC399qe4AbY9QNwgjvJ7cbtC
mEot64zBs5DPi/3BKBFmxS2nX+BPLZDX/aCdPSzR4O8YvQ5E93/NQmS2fXkRN91sSeq0baYmEYeG
IkzH2xcIugKz5R+DrkiIrNHNHW8vGvgxw2w5FTmfGrwwJp90pj5NSkmA0eTw6lE0VrE+VkoxEFNu
EVK3z+9ABaoa5YwZqm/bef6bmtl6zWlNlOysAV7YYX09Arwu5er3W89D0tI/FYCsN966WbSJ9Pqg
oON5XmFhlPosb722iXD22xg+U5hA8hc24yhFmFpbEpWc4Oyady15SGXOgk0+sVofZWntmvI0qssv
S9p5kwB31DhbYvUiU9q+92ceXJzP5Y9mw5MTjlhzjBzptoNNxspLnMT83p3X2e10xqAmcicSxIsJ
L7WLrby6XS2zmLNOL0rEVvQLtfH4Se5KBw2vcVDZm+cjy+m/w/0PdkJfAb2x0rctZCy/nnH4Ko1C
kff/4Du4YUYGOUXpmVUie7ADrdo1q5TWttUOU8Bc8ydwxbJciETX2F9KxR27uHRoht/7YxDJjsNi
B38GvWjJdZM06IpI6ZJAXHmhjrl90J7NY6OG+obxQ9LczGR+qbK9WVShFaHbskxy61Xix39397eX
KzfE85g5gxEOjkBY5lIQkwnVplY35JzgC+IbjCOAvczgugPvDXt9mg0LSq8irqMbcbZSbz0mDKal
bY1XYR4A2+2Eb2niIvzsRMVS9QAPEN4nhl9/J/6BdTglzByRbdmLQee4+to+3iYLWzbwQqiQdwWq
2CsD0FRx9t2R/jiRpkYldZSPeN+XA7BUSarSI0uAPXdjW9S5P4kioYJQ4uU8YDmrBEIlyhlwqNBA
ipWov1XUaikC5IV99vfUKSonotPuKVGB739P8BtI1cQG5lACPaUnv4f4+kMtBLiKLT42h77TWpKv
rnjvSPRJfsExyaFqbQb3Loy6U0HKeGIXbCAYY3xhLP/5TolU4dCLgaMHvq6OMDirq2iTK7D2qSzC
asEOK38Bpi+Dq6x3W0iCjdi4DsLACgpI7nhpL5ij5YLPfenqTo3fN7SpVbx8MyoLrPBc8kcJe4c/
ql0weOjGYdyjf8+Bz5cvXrmMp9shuyXEuurVDLLwCOlwvKnWzXpMnUpG83XduJDinuFRKttiaEfp
5PtB8NxFzqxIe5G/mEa1PnO3jSz6TH2NnUUg4o6j8gBS34Dy5II28Dm/fkwk02WlCh7D8grt1Y+Y
DzJKCV9y+TX1jd8NJKo0HkjjfNCZw46P81lqdvOH0kQ8OWpFD1MmDZBW99hHzVZ7OvyQuYYiwkEi
MCKuAPpA5U4RsFm4CLhxyOSL9j2CEDDFgGYwlcpY6bnvIg2Mv5ru0EGlVHve8/dbNfafB8acMbps
d35UqbDER2ed78pm6dEZlmNuc+zGIABblhT5TI0ck5+v/2cBIM0dxbSvkHr8T7QM6p6GeLktxZMk
RVfR0Uesi2s5dCFNt1Cy3N+Z3ICYArO0bO8a9Ab7VZbg5fiw20Qes0bBShG1JdeeHItUxu5tPdym
bioP1Oi5KAIl8cL7dDG65z4evZ5PDgPuYN3SYdF45QAlaMm6JjayWKILevuK0H1sjlk5uNbiAW53
jv4bvMSyfyycLQ5+pRjmkIa0O5vY9bC4NFBX1FysI4clYbC+TTb833fwr2WYnINVDs22EKZN56Fm
jc2Ph25f3aahDsIQDCaC3tUnA8WCShf7iH4oMmzBHGfy72qjqvvEtOL+G5qgavAF9JzKFGstTn6b
ArBgtMCi3VJuXx9jFHiK2r1/YseD1/uJRhXhI9S/1aK02Y19oljIT8xLPAOc0ny1IwAh9nqwIle7
kLj+QV4/1jVbReykaGnXFHnH7FTQzdRdZcgXTUj/ZPrxb4jeqQ2W6uOE7g3+b6L1o5Zsp4U2CNkP
g2IXmncv/bmjTo/CQP5KL2EZIvntR+SHrU2t1QBdc1XnKzhDmNy92jUpLm8pyxZfaJH4y9gK4fP9
stgRvXHXJPQU5qwUGICVb3wrKO++uYLUKkDPCNqzqiQWLb4p21uw9ZBluK5MgIzztIBMNYFkFCZW
Wb+h9axiBYmF5yd1uvOjNYjoYMzsV+5Nc8bHZXb7LtSSSe7pLdaq9BJSlggkaSX9rxUxVBb3ahP0
gnZEr9/KttXWXL+db+NHaYmko088RcHy1I4iZe9IrgHmJU6GKr090EvJ/VDfvJ6mGhSssD9N7IAi
GK1H36Og37hif/Y2noCOOksZzcb/akKIVs8sVW8FJ3POYmlr9TQx+tRsNTGJIxoqV4K9Z82rkWV3
Amyby8jIwtyu2ctFb/VYemlaDCWq6Jvywulgoa00DakWe9xTiBxsx8x0X0dsHVYvkEKyDPJ2wsMk
UlM4kPUdAghipfo5tydbHT907+w/9KJWS+StS4BG0jZ+ScYHZzBFzpUOtP8dk0W3aPG9FKI2UVk2
g0/F2vniu4/gXZ/KlVSNNdr/xFtN3wj9vfffyahOdrbPuwYw/IgMP4gAeuPpHWaGaZew/5UGZ7Os
PYfeooiFxHyc9szGMLoHQp6QSEl5SslSV0hWiobgS5THqbRVdsWW0muD203c3nRUT4wkKCFG1IFk
3bQw5Nlqja4b+SZzel8xCjdiJV9/rv/xZcp+0PlBwKwtcU9MsSFeD2+/7ZZlk9blMCTzHfv5IFOk
rXVpQOAgWH2/4lqqGjBqLGJqYP8Ckz0Q78Y3D+vEsGoonEeBOlJsxSiOW2CKek82RYoBknEevHIX
gZhAOzZB2bB7C36ghBX6lo+cwOv69R68e22WraEmzY6WTvNXjAqDLKfnfpbDBPElygkN3362yFjF
JwAFnsuIQ1xDOFywY/ej9cv1arqYMOiOrH8A93IjOAl3KRzHhlNy67CU5GJGLuLHVd1P8axyWqAk
yCRNv10R1GfYBhwwPCdHFnuLu0mA606mVbhCuxfzJ63Ckkf/CbNrC4bjhc/6e3DDcXKmguPpYF5c
/5KFsYLtRmm699T8PPhJCh2m2XmEGL5gzd9f6sZEHtFpsT5JYJW3FjQ6oF35Xg610QtU2numFmuX
iGECdoSjjF8uesuhCPxBZlrXXKHec7wuzMjziDA6/nhp1oWCU32x6FtsoOr8xqEMQGejyEyuJMm+
6vHc+QDTmPKNg6fOBDgcGYq8Iw5fbiAlhDSavFvbGAL8xfzfgNn5+G0+AGXsd1KqHeQpz7OEwSug
ERqAOV+F1Z0TviVJkIFztP3tbxWO1BskIdoSCrjHWPZ5i1kVC63dfQtsX5JUt2vpM0pqO4vwZaDu
n6VFEsVzMMUF9+r/Wv1Edx40jRVACXJ1PTgHyaMMnZu9uzFlpX1H2t/ISTjooqf6L4/7bzbFZwJd
E6BUAjPFEOhdZ39DZ8IdGA40UA7BErC86fHZrHnFV4qJCF3n9p7LYmDEgg5HruCUhzU2aX1kNpxD
z+nhNi64kLqxST24ifE9YD+EMqA/+WidalFZ6DtNfsvlEe0XTjvEqyFiLHqC5XGBwZP5/IHcvfNf
LRBBiipDG8DYMrX0+N9L+8YcjgC4HfhxfbD4UpGb61vEGHZo1a6dhjUngwme5ZTGNh35PIednIKf
inLmQBfTOvE9g0SzTG8BXOM4f+2FMpTXPKaYYty5/FEPcwPig+tlQE/ke4Tpqgpkuqka6jbsd1oY
AJ8YgVtgLFSxKIiIOHVZ8SZYuw0uctQ+d+rSeYjZxS1fg3FSRXqY1nQLEETnEjZG+KMr+XiPaJ41
6oow1a1dCiLXcTalKs37VYDAjFm78VYnB7/GuZHH1wU+D0Fm9wopubK/Lc4PfpBVbOpy9dk6rRkN
qOOEdaBpZIkd0Dhx1k15p4f1D5rsRVcv+vHv8SwgOJ9ZWSESNFcgq/IAnqoKn/7KrB7ZPjh/VyV3
dvraBgV5Nd+NxZzzALZg1MTmM9PpROTkO4FMNFT57ARGYpqyAvUxIqU5q++2XWevf0TxRs5JkvhR
JtNU4CwabqtFipsKanKtFXaCJmAt+91/APTJzV03MRVroFWzjkcjxXl/Ecms4lqIW1kxhRcDKb1a
MyV9BrXzaljkya1AHslYBXLDlABbZnESKfm84hEY9jYFgoKjQfiZzWN+p/LxXJqAnjXlqF/LOGro
I0BKdUBlX0gkJnGk7tnzQoIeDEYCqrooqBX5TWQSIfSWLe/AEz8P5XNhM7r3qrfcF5W2gilO8z+0
maQAjWFPLcAn5exeVSGyG3lu79Ylz5nRynvpXWU+gk5xHLDLoMKedZZzBU7HI7Oi0ztLQeETTIiz
r8n/j84P57AhFrOAen1DRqSkJFHJ5CkFMPzV1Fbvl0uejlKpZDCbmyez/Pedmx4XAoEjQl+N9imb
15ij/DK1EqxUJ7NPGE7MkouMzanv1PFHiuazXVQsCztTYZpmigEXCbaqZYSezAUlw+x7Eht8euOB
Zw5BLfpTJdnkCW8mPdTnLrl+QgP9/23reYRKBtfxt3m3yTs7gWSIJMN+mNWfV1SFZnNekOjJ/gY9
h+atiH/FJWTWQ7NPVCUsvw1JZpNLjSUQy0LX5V3RftFcMDAGFsyKGcg2MtB0HalEpiwsJPgmDkAm
uMN+rWxUpyDdWb4K2LTMn+eoB0AtyTspUkQPLGZ5fuyiSqqFLvJGGpWPj1rl5uE09s0x54a+HiVS
GEsWOMKuwxcKElFxVzG7nzm+puholSa0Be975ut1wZv173tPTYPa5oJXG3E4J7PKASBnZXizp+Vy
MA4iiiNSHekJvMoKT16PYnEuLXiPFnMeEsdxMVUtgb7j20j1aY+V6gtHcl8iLHeHAokcx6wJ9cU9
2ah1OZJCaDYrMeu4ZWpEdT2gaIUoc+HU448DqhW82sU351C5HERSx19OFFpkRVB2tTAGiGN3JepV
/QnfA4tScghUc/2a+M+JvH1rjwH1WUCzcXwhnAjpQTvK4eg9bI9EdoUbK6y8upzPC23RtCZlh1WD
yq5InyzUVEG/QjT/LoToKIpuVfOE9hbdeVdu/c7ImULjSUpg20OOw6shEMFa/jo/uXmYbj5RGWKZ
wzDAcw3X7/yMS5jgC7nCggZkRlIFkcfbb/O4fr22hh/d8X378e8MolzA/4Rak5au6i+n7OpTFiwH
Qolvy1P4PIzmO8jIoCq1FGKR2cHBfwzo71flhE6M+67YdWaA+V3fsSGKixRyBFOd+LZcG56fLaZq
aRG3YT/sdbB9pyBCi0P2UWmMdp/7zzcIMFDWOUSalNNWWWNsX5JfblMEptu7xqPsmjNo5GbvzstS
N4YZ5SFGouy7UqCRN5y4a9WAp6raZgAcAxN5zcACXT/omxqjFK34BS8ADYgglf1WqnoX2vZFzcJd
AVoVYQ3JFa+fsL0AuSR9pb1U1eKDQPf+vT8qpDYa5wTluWvhd+7PGgCZICo9Rs1zmCOojpHCbRo0
pz26BKqku68Vmc7/B1l5jsgjjU4c+APEYg3AiHCLBKyUXwPplIfI2DOlXl/OymBP4D/gyM9ogpuT
xZHKFvYDi9ZE/MFllNfVcnJaLY+RSAetQBhWEOoEPDRuvPSRhuYkVUebiC9A4iA0aClqTwzYH0L/
zWjcjal4C1WHJavlRq4xdxa5lfn6PkVSiDw0EjZx1WjQeYi155Ic5rogX3VgKBGXq7c0n58+eOuh
Wi361F8PmaaQ8csZxiJs6J3BnQRNwTc6n3FL4OVB6rKv5mQJoH9LGLK9TGpH/zHkFcO1eTZitLll
YijFs8W+NuIKdO5t55YYsCZKkfyDK9+D+oSHLnLLxVUrVMMjz4xgefzovMN1AWf6iOEMflCnnldB
pxPtUm0Wz4qBR41QqW8HL0nRkKdEk1Iobs8wVUFp4Nxm0pAbrHv+A7olDDO0sRoctaVTX5krhP29
m3IKWfUO7KItvTy3ufCoJt2UHe/5G2AV/yD6K13eGKsHDtJF4eSGqioWGndFt7CiVQZjmWWzet5I
h/nayZvovhYYv/ONy7dYia93kAMq6sgrLcPOwxfG66Ojzlq0GEdx1tG4h6icVOLDpB20nmJqZriV
qi7kHv2hGzdJZ+KPSiEqRh99lnG17V9OeD6JgYjMUeSwycZW2KivVDooGieQdwq7qa9u/MAbSmob
h5bg7/lKDDcS5ju23Agel1oXK7gAVkH2o8DJXzIX6b4EZP2YCGStldp8DIBeUkHzXGciEhj8OTo4
pzpEC7vtVdHlOopuDNqTAsyzqg0MNwTFj6BMWb4Ba6RUdtiyyKZmxcOSJAYSF3/l7AEahzveEv8x
F7zWR9RLo/uOu/hLvPBNpKqwheT/blGa8kpjzQ5hTNFc3Kc91zcsWPLfRT0ZyI2jLS8kuM44ocJU
A0WTJDe7iK93VPYKdmCSCmhEkO9PZ+TtifznyhVxIDWktdLbo0zmbtG5oYDAz75WdtnpLGU7Q7Mw
hmhweOBvFON/9tyC7cjzHRIVAftK8X/214nq3Fyt51KWb0O8a2F3f1+jZeO8IFRvkgj3ul2TwBoI
hpQGzCwlmws/DDxs62RLqZokl6FQyK3UY0wRUjO2p74nGwJRYHBRHqlK16WiMbILa3mfBdo2VqMP
Y37bO2H8ZbDdZQbtC7m2ayXcLnbmRyvPhOdnBLtK+8He8xdof9hvRLNA6XeqLGrEQMcy13A6Y4bi
5VQa64PVDLvTaNNNPJdgOO/xbdRA2fTb9OX77YmRAAi8qlYrnGK8RDH3XLK3slQfy4I7y4ohmNKy
LzytTdHfCJSSaw/Me98sEYyDtex8BY6jSDXxPkcy2SNDeETFs0mbQN4pAGTHWsvW3p2As7XXVckn
+iAWDOjbrZa810IMAVxODl2GikTvKx8GfgiZ69syD/yHPvTDciqFiDc65c/TVyWV4MOv0TB2ib8V
9Ohm3jMfShvjlOgMboZ8FzZWIcsI8g2A2CoUYB+PsaBOLzj2Bmrk7hbTeZnzf6WZoQKdYOJ+kUk7
gRbAmFH1LYofKTNKdRB+1YZIHMeP0oKkw7k69E1Ax7UlZaCkKHCOKNYOTbQZ6QmJlawDB34qA4L+
sjng04hb+3oWpE1KBi3ZzSjxjMfZYe3QhtgC7LwhwGw8E7UFGss0nNi+HMbXuo5dhQ3smwb/EMt3
7/5cxWBWbeFqXgnLf07X341gJw+4AR4vOMY6oT4tmuzS99nnHZ8ZkSyp+Dtwi/LGN5ef5FIGd3fU
Emqf/vS8uIUlOpcOyQ8XKXvyxrCe5m/OXZeOCORxExlbEjlPT0uBoO3oN9zHoFHFJx637sU4+x9Z
n2f++qVqeP2nbRJ9FdaiteGNy9ZjMgztyFezxjvdSEytToaV6MrUWrg4xStWoesZkc/uQyRpC2jo
cyWvF0G4VahmM4N2XYjHcxE4XppfkJlVHBtmH0AdEGZ0Tor5n+DhXurY8qv4QGywAV4Js5xcGVPa
wTzj8mCBsWQmBwKQZVGgc/mmVcsvD6+g2m4+FgzRd6x97pfVxlrDZGwcC69RUU6ifG9eKiZCxKWT
ML9oBDYgBtEjjodfT6y05KIHbH2ImWhOMnwJxnyeMOIE1PncqSdw/gmvschoY4Seo+dIAQULylsG
/wW1MMT1b2YGnEaxzUsc+LeMgH0HuBkb2eJTV8VgfSweCrVI5tqohSsM/yKtFPoivMoC7aMQt6Um
PD8ZRKlq+HPr4nd+fJNom+40TVuAj3/2LGwGaPxinW2UF41vE6hoGSHG3uzz709Q5QGRP8v6RfsO
6rZLCvGGZeo+NKewl8lVRoVDEg8htJw94U7X/KqjN1t5ZR8mfzPV5TBV2cDQxwPbeHkBGUR7qE51
L+OFOH5tFR4qmg6nbchQD+gW0kJavtLe0AE3HupATwssiYCItLpHqhmTrB5+wTq9VnxXrTiVUuYc
j8dc35JK/kgUk9c9QcsQiYh76gjpD10u84A7OGFkua/IhR0jCzfx4LzseR3/pufGVliwV8Rq1vQu
hq/pmwgf8Mc/mao98YWZGX90y6QHCT/h4XO5LTYF/ghTlt5nqJYZZYWC13DODZaYhZyiP3bXNe6y
SL+U0/FyUxUoq42Q7sv5n30SHc/eqVex+gxHKBCUpatbANpn4qLXLptid9CtUeBqk7gWS+QWdfdP
UXF+CANfpeJAdYl5shA7XBTtB1gug4rpVVJPmHehTpcGzGSeXLmAYNZc4qc1TwJ1k7GPkC+UyuC/
/YFNxu+C7V7EQlAsweEmO9FEf6jNuluTxcUKhWBTj5jq67j/3LThC1HMosYpezF6+HkfZ+R2dlZv
P4Yu7Fc3avarC21t/jCMH2+tnynDSZSTAtqFzs6/1duWYSdR7ZR+I0sUtm3TVZn7GHxXvUGfXDWv
yFxisEVqD6k9ddC7Kz+oBq5m/24/k/1RHfmz/UBJT3NOqRgsHfnPTuB/kQaFKPU3AEbSAEgA32sU
NFw/o6ODCS49FiMA3ZsjL5UOHYNFFewHjgEr6WTHR872uQfyEUItcj4YVuy5ZeX5YhPcLBTBkbgq
ZLUkqmSMkqC1jETz0pGP2lKtMC+jg2swb8UuDcbhxt+DdAArxXEGcn8Fl00qlUJaqIT2SDvZdiH8
p8hJO0a2qTATz57Ekc1/oL1EhK+dgFN8V2XB1K6KEurxhV8lNHtpafuz90lh/Sb5N9U2A78Ht3uX
1TA6PcCi8ZN6qbaulO8feVkAvaK2zZ5+qH00kiHKDMz0mFs920g1xNlJTXFBU6s0albmATKXsDpU
XVEeOtIR+DVwsmfcwN2gHq9pw9+PdWy65O/jy2K0mnkaSVBo3Fehu9fuTgZMHmFICkWUuK/MOzw6
rRkWvZcsfoR1fkVV/3dOu5GWt0s1NahbfYgryfA0H6rmIkWFeuvp2SQGo65tiMa86R/Zmp1HIkxy
wZ677dMQNZQnLOZPSn3LPMgSSllryMRBdEvuVXzkXWPerGhwyphJ0I/q9w06QWbHhBsZY3ssnASE
VPxbHW0JT8Zqq7oAvzU7DlqxSnDwSbgYYFGbT1IoTFWuim81vqxYvXn5IO7YNzOjjlTVljksFldJ
Ej7UoH4qdBleQ1K75d3gdMSRKFLoUvlZOeRlV8WEGmRYqQb23PTthy1oFjdDG48gswlvC4uPYUNl
+plzrvvYCLHrejcJD3pcApArq4j5cgXCdrGcvvUm8/k4IK+3GFvJ1SjT2d3E6NAwM/KIR+/udosq
WRKH199G3GD/gE7kzczM8Z6QP/6WlHAa7Ezfwy4kHbAxgELp/aedKqTMi/+NR9l1ate4Enwx23gw
7SbfN4eTXhy31/kMe1B/tHndcjrL+e3M+e5MTeTT2yJqL90qSYCQB5bIasRRkajh1Wc3SD6rAc2f
FMH/tERf11OQAazWZZPnEcyFf7ZbsNP4TfoMqZof77fMXLd4iPzPFb9nKIHKjlFc/icWIK5zZGFf
3GCedgzuHeiHcDDKXfciL7zQod2m/HTvbE8bj/VIRh3jXpk0oZxvitH9DOeHF9cZPTZJJKjT7anb
7sh/wgmc84T1IhF6S1kNC3sUg7hdw1pzGhWNSPeTaMGiXiLmuOGRMJhLKyia4zrsCVT9SxgaOSC6
aU5aVnNjewpubR3tTGvhegPtnPgHYKFxwoHuOyvVGJoovIQBCNUOpQ9I1B89gRGexyyJBrHBA9ww
MiUJk3/pWUhkezQpX0ol2lif3F5UTfWDJga/9y/5MIADWRUQ2HhHJqfM+9GLV6R1V7DyNKfjtPZ5
FcvSYJy/jYr5sFWSzHskLAoJdVLpdFRiAyISMjCYGGc/EckAcQgQFiALyQlpksWKQUG2Q0qyTyGF
KrkoABlcLRSFBCd1RrukkdiMdR21oPiX6s69LHYHC1s8SRIWwckTNj76FYlVehNiFbqqnl1fnO3G
tPFoRgPWE1nCmqxYN5GvjhLYUOwiJPOi/+RompD/0HRsReM4UBrwOrTZ6QWJ3UVuXVVaWLFpXRrY
CxI8bO1gBYEmPFipOXkqnMUhxOLMpDdy4fU401LSlR6CO76wJiI8N2Jvctc1ORKxu8N0FI2NpzFK
c9UeKvnoUihKmrcRk3xizbMA87rGiVQCz/aAVOqXoXJzWIIx8ae8iu5A7/BN/tQZXbgQR7j88R6k
9we3upyCBVdmH14NKFQEI3C/LYLFucqKIu6dGBYVPoFi9Mhq/GJmTid/ikinO+txfLpc3sZpVK8X
E8Hnc/oDUhTPY5GrzYPX4fUJcn7V0RuFn5uCtCfk3J3QYimoxuC4HmZEp5OuMBm4jWEtZc36UrWZ
16pB28n0UNohRxf75+XWHEXMuwWtcW1TPoZYlwXzQlcKMwqRx4g7SrWlvxrhH/ubtIzOtmQep0II
nLSUmEnQBpnvjTXiabbq9y6kEprPB4WOM+M5WianzvMIo2L7uC9S81J6WnMG0Yd5t9bgUC5uD245
Xphqmzp2jPUUtdMSTjQsR2ZNpD7QeOtEge6gDKAf+5gpeXV6zBtAc2oyIR0UT4dTxAnpY/SzTwlW
WXdlXBzLLCxaDtEVUxfELEZO6wlB6lQR8km3+UQxBYfiy5aGKrKOXx2GayKeLazyViJtZbitvnxH
+PXCOy0+xo1/GqsxcodvqA6d8zdPtj5Z3rw0TyR5kbrDUvvxgI6ui96yg5RDrTc95K19vttCGRrM
SMSvSArA8sccUOaROThIhZbZS9yzLo/IRdlUO75d59r2Jek8c7/lL608wpptd3mebD8mZN3M5mab
ZTUbN1msbgtUQg1CiS7zEGgyU8447lckGkd5lH0JeqyCkJek3f9ZqqxoaItfx/IpaLpGC5JDCnNX
HCEyEpo/yu8iGFiSKUbQfYxkKZPWqpnRCCl0nrqEdWlzWd/KJD1bNwVj/UuMz9leVqoz1oRivSt8
zVGeEIboDJ9fxv3JHSe/I65C1EKZ92V2xW4fr1cgxRMX/2zUPnpOZdVZlWZ4BMp2afzfE8H09MXu
UqIUqagT8X7MnYDIYw/SdzCJibmj4nsS0m45Ut9xkyyyx6NCh2Orj/8oQzx+P80pzUzXTSPwoTb0
yG/G/pzBBbegweUw+po4pNLv+/L4CFlflYA4J+z3gAEshk1LgiaQzTNhb24xolETT1Ys60ya6XgK
wvJBOY68BJDm7qFtDF0BMcKmKC99wI2m69SnQDIkT0BInB1nfoNRTAeho3tTXPwYZgJlgFR8R442
xT+UpxVaSdGfGi9l95H4nLJAMLzYMMMVNajUmwM5BR4Hn3W7LrBwJbuWFjkqlr4y4bJMAtKkSnZh
F0rbV3DKTpkpf+QuwjCxJPR+QddqCfuOYNgibnSWfmOT5EZQ/7SKc0U4XbdPDSnTVI/OmH7BVWIs
dIyxSxpR+VYtqw3AQ8c2HxpPhFupFDUPMXphOgKwP44WW1EuzGRESkuSJ8Zw8rHyVMymO0HVS/8M
QbobYBeetmzyXJUHORWMEUyljpn14/rofNlQanOpTzmeaqhq/FR4XxkWoRBbM+pvsqpBHz+kAZZG
3bJMGfNguCBxHiCziqxjeQ1KPuP0DROilY4RaPrFZHZ9b6OaPe/aA+K/X22vftPo4fYqfcE54gIU
qkCDCgEYFJFt5GQEMmGTCAUs3RWF0jgNv7dWpPODcnwjhk8mL3Be/muppxaLT7hklaRHZXKFmHkA
H2Nnwc+6NHO7sW2YcJkDz18tT26nu6u0Y3t7kSyRiNF7+AofRZAijyNCtysSHyDfmSxLyvWkqT+W
D3fvp0lobyoJHgBKH3tEbBqO8xydqKiacwca61N/96zE93RyOMpDYT1XcH0wkbMjfn3DbIZ/rX3q
vQ0NRH789MkZjnoxKiWztop9nGlQFiUcZcoR1C9FepvoU4/mCyuxCLNiXgF/r3vCoLkICcz1AGsF
SOjp8TiG22K+LE+mueP3j/7LmG2PnI5/NRJUGcr2w4j7JLeYJ1SgW87BAbICjxog2eTKdn0/JyNS
F3vUwzHL3c6dtt4XhZhPX4Qs7Kg9rSwBp+/LzAjQCVkdfuSRTtdX7h+coMkmc/ZsKEF/jdcikTFs
SxBO4407rw62oSSq1thwsDVaMk3IGM1mmzoOB+HmcGERU9pc8ROSiPxwAXfYGoVA3gzKgiycw+La
GnpHawbXCziM7GZ3ieyuuj2Ith1qnQ4CHq9gc9gz0bEG66BeBwsSbbcDJ+M420jTluE6Gzx5yGJ/
ApVaNz/NhQBWZfDKvyiKDvbkzMpolKu6R4Wo9M4cLBYiN0K+V7q2z+MuRD2IHFmAJxPuTS9J/qWK
MomqY4idUuOQsVQykLDzxF4MpYooJcfdPDcAL5svjEFlF/8Frzzguyv2xQDzIA+pdkqfYuZSgCzB
rQ4dcJN1b2WbQ9nNbm7RZWCt0ZBklnExtoH+B038gawiUo5sfkhE35UXkaAzn1ibMly4JsX6mKg8
KQ36Csuekt1q1t3TfJpyJprA98XFMimA5khR7VyYCTQxBgoOIRlToZslYhtsL/rbvBx41jGs7768
I+qQOGtabjrIwff+UDL0iaipFE9QR0aDj76v13uw+h7rAJ9Qprp77TZiaa9fBlgFcafAYj1NregJ
5XutNdAOOaa5sKc274eNcsQH+OCjUy0qse52egXuUn4zyxYJr03s7+NeYhsJV0OJH3vfOHlVacSa
hQ/7GcI9XGA9XB7rvRulX/KAhC5X3JYkoyqvglGx+u0UzVILixos/6qSLsYSx6IvLsm0U9wV/ERm
Om4e7xRLhWYKj+L7PP7OUM5qLEv5/jvk9BiKppOJ3snkK0iQ5/Fj3W4kVMwZzME2DuaCJFHJg4mz
MGeOqWjyQJHH9WWaNITsHYb7BgcAsekBUwTDNOLROPaKOgv6yAt4chNGcDszIK4O+eprdWFzFBzf
Quoc3sSGuKlTP9vunUdbUUh7UjmvYieh1hjUb4hgJKkgrKkRqytzP/ftAqxAfbNiIBEobjGRiLQj
NJak/nR9mlrdKVmZoxIfTtkMsCkeZSjjl2yCZQIQfqEYWeR+qyk0Tb+RApFwBG04kBQf0Inb0Whb
wYJ6Rrj1JheoOsxAxTzvBDDwzgObJ5lweHiNDAiqDp1SguMQpq/QEWRSqt5/aOHXKOQ12t1hf7T9
t3OpMjszkcX3bSJJuCXQMGM4iE28vvxgOHlQiYA9E9YkeqmB3CncQif5GG1igWwrowGZ5RkSzQRa
YEIk64eKksxHzf//RFebn5DLcUFOaO4eyrS0v3+q9pcTDWuKWlqGEWaxtlu5GtEnLC0pAlt+WXe1
Gj6Zsm1SPuvtj5Sqmc3M0chnZ5/GggUYXnF3SVPodn6o4/zWQY2yFF2ETuD8HPu1oOmevogmcpBy
wWuem3ySCxnKJK/7iInHnSTojv7F+CVcURnRUQuxc2SKxiwQm//BombVM9v9yDPmexw4uEmjX5et
HcTjxyJpegk88gdFJ5CLqqbxqELXpu70uup0Cb7nB4ndxY5lutIex1grJ1jUuEfhMQKTEtO7eFEb
9tTUy5p6XPX5ncjEiIdauARfc7QGXuIRoZd8N6yNyzgm0DpEr1RdbtUgBrLzw1SRrRekoAkkf0R2
do6aif2x2YwvKWuQQIYbKcsMqBAs3BcJEn2+jYCbHudFDUk4sxLdXT/vY/rQTNOmTFvwAKCqpjFn
aSrNuCWs+C13Xxy/ZyGYKp3i7zLc939H5xOR9786tF81sW7O/6bUB78cV64QSPl/P2cDLkNxGJ3C
+41XP0zwxekn2NmWo5116ms2WVUHa7kEjklTGlCYn7iQp7NSXgBwlMqsgmZtcQqaBMyrNKaoblBj
haW+aCUznRHo9uFciFscxsl+qAbX8AL59vG/j1gbhiBgIDlruMvioBbg/IkjUdisL/4fvzW6ALMj
Vt/CuPOMFrH7jOxKdQicI8/Ihq+Xrx0QNLatdcOzF5nQTKQ772qaFYZSaDyr6eIO9GIQKZuZn5h6
bgN/ulsa/kb09mO7GL3+GGvwdGhWZyZuvvptSopGhGav5BLCBjT6uBMiBcKfCm2HUGUgirSg7/gW
oS/DBx6/YqaIaxG7cjNVITrXY2AMV8jXAjb5PPzRcXZuROCP7e2huleRNzD+K13pgnCUmJmEMYgK
5cpfnpNHBHYwxayd09kcwMdhX3fiwzDxwvV1lmWwgKs6CYBP21lsaZHVaB8dqKbbFsGTEHT7NWCV
A7Uke0HcLSjqaCVqSa0MMcpamYNxTKKrJglSL1Uq0wylDmYI7WZ2ZzrsMudExrr+03fCbz1sawoB
PjDRSWTdbmoOc4cDvwwC77uu0LexOv+CzCrht5aEY70EgeK8xc1IOK29Pndb9yPZp/2NVqaSR+x2
tIbElHtrdTeoL4+fr7EBnVgBV16HcumsVv5JNbSAFmvJydj1ArN0pwlktNqiew0WEXxetre1Gkys
Sj1P4FIzdv12ut5B4XO8YvgatuuyDIfMpw7GHh1cO7gc3zD9oTwXNrkAMKR4jPNIV4/OMkGbBFV1
Ajb5S8MpS8iQcKfF8ydUk1Q7sDTv5Bc300Q6c1WZfRV6oTQp4WwJeYJpmYXXIP0DkVnlZdho+4e0
aww+6juro6+MTZIBAL8Bem/pid81uEOEzsePphx3QpibmZYT78PCkTiryCegbcS25gbnWDN4hFag
dUFET1zQU8LVGLcOwgSTcrOTYeLn+sKRAhNrG4JxR5h68NVuF5q1smlcTbq6Gws2fak6oP2oNLsG
wX5Xl1z6HS5wcXfx0iy5sCIuDeWPZ28P+8IVn4CK72F2tkDtJfd9wSToiDJzv8A/k+vdya19N94s
GpFRJ3WNJbcPx/ndVLDgL1cYzmMTHO/WxaOqJ3hQcFVAKvxz3qv9/OHy4urFLUeEYHpL1z0GA+6D
6bGUxdQBXWoP/pz5DHpK/k2Xm542IoHIs+eWiai2CAP7zKBENWin0CFYo3ui8SWRJJ7TMoYpxEHe
DpNHgD+mxZhnf4u2pUWtrTrKTurUyAAPB/JxKlAP1shdXPC9zqIyIv1x1pYuc6JT5H7x0cgPO9r7
PQeKF3EYd8Roz2oSSj121/gVqThnTfVTorldZpjfUGfJ+eHC4Ty9XhfpPIQc1ewxN/+WcyFiP678
g9Gbds/m2uD2C2IgWbGU33FHDVrPxjYyZrqXc6WM2ZUzlPeXd5z/C0XNlithjs19YzOkfGUNIJib
XF/1bypwEMQZtesvv91Mc/YY+3jI4kTc944VEhwgNqZ1zrg2ddmOjfj0Gu0ZC1P5DFL4VvpsW3WE
KJ5J3uOdX5E0LmuZ+1aGCuOtly/YfoLjgTVXI9dQRM1n7iY8c6s++cs24oyGWAQhHnJ2XjMK3bQw
e2a81Bo/nO1KV85tFr/b2ybqaZiq2K27h+tP+rWjHbOcc/lTJsI3KQLXToT/CxH45JGHk72W6aTP
eyeRmfPd06tb02I1ketunZwrfK1U/T+d/4VEqJn2wEbeIVyVl899HG3ZQPKjox/Qwr4SqTzxBy3K
NBA0h9U7tKiNCCt8SU5krDjOcAAU2J3jIHibTHyD7z4UTI4wlNvnakV6Q9SBzKztAlBxaCz5/xbl
3WShgwX5gBPZZPRqca0eIC0hNZ+v+eg0zNDqLS+FDmep2CuIRxc6VW8eH4RQ4JngT81LA8Hf41YN
755Zo6S5BE7KCRFuoaXRu+XJQH0XXvjAwqac+S7RhDNi2bQ8RR/PASqzK7frhUg18EArjEM7f8yg
GdlebOOMz3vO68iqB/WVq6gz89Y3IZov7r5FaJbuZ2npsAQovnSxTxFLnzFjqmNGDtS9//nSm1am
QFpcnER2AN55ZmChW8wWj85qU/c1ONs1cagOt2NXex13vsHGKuaDIXXpI3kYs3Z8Di4BxPTUfwg2
/RRvLJ/NYc3cG9VGfdXynDZHW9uo2grSHejB4RPjeV6V41Y55AMn5gtdSm1kTkvs3yudlPJo6W1p
9M07JNGEUsFGBWCGZHaXingUd6qngOrcw3RZusAW5euabRVEVrV01s+jWWrDHCO0l94L1t0iZ/5+
g7byZOLCHHzeXsMI5AqfJUFqd37acwmL3TjE33SrT4U+le9dQigqMoINQBTvwwhYCi42+XUhz3i7
bgk8YpsGNXdNKHCgCEsflIQWRBl9yyzMk5WpjQKyo4FTOXS2pxCKjzPQLMK0Sl3V3RhqRbjcPyLE
ypVEegN2GKpLJVnY4Oa8i8fekfhKT9EBhZNsm8GJTkCYpQnT33PoiOssvc0w4gBDIAcLKs5eusbi
HjiYghILwTBuvlm7CgTtDVfeah8GDdZb0Vxo8ACK4cH3pAeiN07QaU78Jd9KL4wZqHYmZSeb/suN
Y1coHYIOh2ztlSyIhTIF95TH7BxXtyRTs84A/xWl1uSeJZfdqeyow5cOa/lP2zaDi9Ie21QYk7se
aKfC/e4td+U1Qed+fKXuNhaHDnyIXn5cwg1ZyONMR9lFR/v322Ob34WM+CcEtHeqyG3GEaACGJqv
DvFrhstMzfPO34qAp4m7MOS1SO2fhOFlb18lz92Utjc/Yyq5xtppkpP1wPAUANCIw2pPhlNhy4gg
YAhlRaTSNFyDjdHk8MC7xtkXnoCEk9TZM2Tjp/z/Y4lrfX8vLxE9mMuXbaXtT67lppdj1O2gE1tZ
3W86eMAzMQFmMIvZQZ7vXfi9MtCRhR6dKmNKrfnETCaG5nPs8iC5sdPjP4IueRSM4se1hRKaMVzq
FwJlNgiuo4/kTVR8y0r6XhJxAj4rlJF5ILJNzsGQwNED1cpqVtSGzWp+1Obmi72B28fW9yUt0BvT
vrttAHIM6NqCiUKtaFE/X9VLXhaoDoVLe835GEeu4pVQ1YxO068ys/HMoeycYGPuN0at+e0q9rY+
xJsoUfzv5lubQy1/8nfexp6wJUY3OscZyXIk7Yr6vOuV07BSR8WwxAi9pLDZWKQx6fbANp77NJ+U
T/rPanDgNcV1SYbrx0WiZBjxeCeI1n83r2mLEriu8dKdnoiyZwpNDgFvX6qyH4JdN9GWtaxoPUBv
IeaSWx09g0gXESdxVhCHUy0WQ8wSoCKaFtNGrW4hQYINJCMoCOP1O428qBBIsor7ePX9JpRn2hED
zi/djLHKYLYmbr/+FRHx+jjp5UlcBi/6SGdlR6VU4oM8/bqCeDAktxG/7qGeLDh/YY3FfdiV8bWc
ayb5yt7t9cJMu0FgOfcba2YtqoKYNyqv/mqcKVxdwQWbehb0Uu6e60NLH3l9/WuTmsUopb6Wcppi
E7GTDeaK8m8G21KhGHoiGuSalLfZyaZFxTWiEZllHzgMD5bpw/1B595mglrBhdpINoTY9syI2xpU
hES40vnPhqKd+mJaB8PRnTIniow9iGWvD1uJDy4ZyYXIKSd8JxB7jPYWKdHWwdjQKVDPdWbgpkJ0
pNcwJJw3cFZulYZW3vYP9aQ2RQ/anRueVWg6YE1O+HhiGrLqQtELR8t4lGagUgG8jFMdLnTISDaC
msCjcdCvi1woXjAYUUBdofT9DEmCA2q1CBH9RtYwT3EP1BOWkpzWOtQ95O/SRXBNVwV1hLvuKRfw
Uvoo+ulUiZRawyN6osioRa+255n3DcAA3Hi9L7AGyOiGbe1x6eA5EdBKoLq+9pOK1Szy169ID2Q/
ig1UUr0HOSVj84pXw48x02Z4Ufb0je3ujIAcFRKmtDgUeEnre3hRF61knVOwpwLhnVMr+Wb/X9lv
P520JEYoti1xzdJYVXDBDIl+9mtfC32cxLmKnlG5VyGGJb7dd3jMABOdRyjZojnoj+UoMLY21stE
r6ly18ueFJVHNlm4SxsToKbllhSIpwGi2bjYbMkkZ6qRyac4jRRBCN12UpSKRRGLdO4/A0Z9Jnx5
rE6Jvj30Q5ZdjmewaeZDdKxq/VCbPbvcnD3ExO2bdJtAvxMlv5OoQA9cOdCINHdnd157I/LIUGan
HITGhjQRDAazFUa/gcIK754+1k0v3GeVFn65baelMJ4/BZ2NpUVS03uX5+hOITXH2pElyVO163VU
eV5ag1zJCBMNFSALgfyt3LbxchzWo2jfcdVtOetIEhdEeoUUyGSLEnLnyHcAeUlB7UNiXKR97o+i
2Dqms0uQ06X23cRYM2dfdHTmiCp78nBvOyXd8n/VK3AxYIqIOF04SsHvCAfQn4Dz1t8ZOind1Dfo
/5F9HBcSQaAOjG8bgnSmArwy21pf/sGrD8fztXl7abYj0Nx9JEGqInznikzhJ7y5Ctp5uiN/yPtl
dxQI8uh0Rh9K1zBU4FImJty1U8+is0BNuted9gnRH7yAF70F1beiVL93KdTUEBU3z5/hBXjx6Ae1
6LfqyR1EfAIKalm1VVK/GLmypN1MU8KhwQ1E6VxKBi4dZtzSOALh2Z5yo7gbrFRjcDQib6KZunN/
ZVkkizsfmpObeBAx+P7pyelgAItoQmB4pP8n83EK7JP3mMzf67GGkLmc/Lq+3tQ0Ju7T+yENMnbY
PbfewGHgULa0LVwVFw3uyodDvXDDET1AXQrryj4vMdC0skyxa8/zu1eafJsBxJrnNr8aoVldo0gO
vkmB01EkjNHd3O3iVZENokwWiaHnH07wat1py08zU6Ut5cPftxBZz0/03xfbxUpb3g0Nf9jPXqrN
PFuKSdfbT/VROWtbFYQPEUjp7Z1GqpGf7hN28PKvShQ+VRH5xPq4WUUk3PR93xSPv8qR9YJQxkp8
T5HatxDlFZ3FyoutwfNBlaY3P5xj6Wv3hLSs8boyqWO3a11zHaN+2LWFEgZT/ZmjcOA12RRf38/P
6hCAYH+cVd4GHBqhW6wmJLsFVYCDI6LeXFNbI+7D3UC1xCdudQeaIn+WdYqQcIUbgAl5U6VAQDIa
N5Gsm86a3w1sPg4UaISOD4xh4DxSo1se0VFXph0ZJu89VsIUWzGVDzZy9RjG0Opvjo9bMGWBOpJe
JQAaiUr0jpB+ZZcS3aDxEgE9DCigE0uuWaOyK9RX3A899X1Xv5+HT7nQgZ6rUGWDb1T8Sknqiodg
US1NmcvveklDQNXm/3U7r1zNdXjr1A6RviJATZufPzCcMBZqmQezPHS0l9RLV1e6dvTa6HSIKL/k
ZKaQT4rYOm0GnxA5yMtihEcMC/EByHa78FZyXdhgXv0CjUZWCcpaiPt5fjAjfq7QZ+Bp2R8mbY9N
Qqv0SmxImbHOA6kYMjy/lnHNHBrBr9vUpD6YSyD3ilOHbswso5eQ5YVSQ0t8jx/3SqSHeA98HOwV
74VrS14t8I1gWF+rxalCaT6nAA+4xJWqydQMVfuvtiWiKqllpeZZxNEuaR35o1rFJgWwWfBneEez
m9SJF0R47XrsepeDNY6Yx/Yj0frXIBf2uMUBhDih/XNvrqa2j3TTN+Wia19wl2n6ONCItmakXCP9
PjW6ec+7QyehvR9PxV7aGStlaBtksmvxZnnkK0Egb0y/Wfqjlz6gqhnUqxyMkpO0wLV1ydP9R5Tx
KAsCDkRct1oTnzOVofJ4axlWhQd7eNz1mF0fP8uMbdcxaVitUVPSQtTSL5U1Lqm9G0fD1GUvItjj
O/RjUMS42N/58UipINWOBFdL2KcZLoNCt+e6zpELkoYV0XtLFjRWaHfc5AyKrID4kzawCDMwsszn
VdYiXo78MRVTyxDdPR9OtLloxdv2t4857zcXyA2UBPfaQzMae/0nh93Za7BtcazDiSFV4Dn30WRn
HgB1pR534eVKBbbpTc0gtR5nrnQTql/pB8ktzpPqGG3/jmc3FLNmNHriHlddTx8HNhbSlkUAotAD
e6ThIPi2P7V0sCVUkaXnC4G0AmVOFIa1PGaoe2mRiz/VAnElhuWldl9FB6gcwaOBSOuQsMY0SmOO
L4ZfJRdcQ6PFSdhFAoHgQLcQvsydbnuy3hU6Ys1T8eTcfsjErZNI0aKaZa5683NZI/DuWzi7Mkne
uTvqCdFRAGASKA5/dItAf8BH7LiiU55v9WchUJ/GCAMw115mLHNGQKImaAvWqhOFaxvtf/LpbCIl
P8xptyYjAchjVzNeR2XOPNfWgLBKZyq9rhLGlhc9wji9ej8CgxB+YmXVsbUObOPBvP57m11MWukU
IS8VBOKyze+zV9B6CzcamyZoksS1w837QGdDTuFv2I3GjraaCize23CBuuGE8Asp6eqjFpg0KpMr
hKnVK1fyV6z6/hdnJiC+lEajS9OQ60afa+9jodKBo6j4BudIub1PO65Fn6VI8SIDT1MepBUkjtlE
mQbf60AGJ3wlVBiWERuoOqBSIv48MfKMMGPN6vY8g0+iYHoy5ZiyrBWWT3nrD3CRzVUvbQCkIFsy
y6hz6HMVCeIkrKFHDEB2FSB1/uiYutx/pPCnJonk47BEBz7u80Eiu7mrhh1y9T2L0SQXT9bdRAFu
bsUnOZUxlIzjbtKrgU2JkpVjRnYtHcyxgqA9VehP069Gu6LfC1J6e7TMcuh5OD25pmnr8+iZYlpI
pqjyRa0grdXvtWCCxecKGYHZ7tcKxlJ8g+BTpQsb9IZN1NYgETNIjm2I7j1ccoYcKJIFmS2g60Su
3XYwzzQMkiJI4C6jbgJFAusjMKdnTwohPjeB4tD7XLLyFRLfCEvKqlNCgGkpzE9eNUsqsVrVX3eJ
5LJN7p2wOc2l/oxLw3f9ZrGtQHz+m7JSYSCKzCzzU9+Y7Rd1phL8d1U//EjMJxIVTni0Cu0vD7wC
v0PY99NnykqmkJiYnpGz2Urpz8pzVSiqx0fQEjcQswPLvR3LboPtH+np8/g/KJbeB9U1qpZcFscg
K4TMH0gDTwBnnspsY7uuZbvZ0IsqHdhXAI5DzQcBM/3gd48uV/3v+6Zqy3ASmsYBX7yISCZ0K5J3
guzX89K1kgR0MLF0g1t/XQjJkboDqu2ugQr5t5tIIyUc5Il/T/jNDCURCis18t+eSeD4KAH+DZ49
4Qv932N1yc87xz9OBgm5xaN4v27wLAof/e7n+AxAoZgkptehhHN696UzNEE3wxPUgESs2HYfb2Ah
3OZnkWLeOK2oLbnQLc5HzIRtJROpXgWP22ieTvKbq97jcaBG8smMrPCUvJ0Iu9R2PYV0L3npjZ6b
aDy9DNRc9qUglJtTqn46BJcpEtFu/BfmgJ38fp2is4Rq87HedZauwbrXQajctGbbaHvkQYpnx+46
lholSoHPnZrrSv4x+lBOfFkFj4PJ14yKT7EOc47RNnXoTU7vwSTLt03yXrQuhcIBQpm8tjEmKVLk
5JKjH+ZTci0b+KebcjpHOLSQw3hzok/yirzQ5OERCrcCGzwsSHU5QJrF/9+ESTcaBV0wiA5UagJL
FVzYKdo2UCf6LhHrgvZDPM7yDPST0DRIOCv1s2Qp1UwU10TE4wvTtSeBtrf/ZO6EeW0OmGEJTjU7
LyU5SnUI3vIKLADazP1p6nozb/04dhR15YFNh4ZeAUuFjKzG2dvFNuRgU6lGAWafJo/F8kxJw3MG
KPjvK9S4yIGAvK5WATKj6h399yU4sRv2yukWbNdXVqHgZt8obcB/0ydHG/GcEUt5YyAgSnf+48IV
7DnuNgbn1vWmghhlEdQrzjuf38TSxcLIcIHSdwK0Y2d6UuuS9/KHXXZlSxt4QwYiMuUYMyN5Bub8
6sy0XPUR+tSzMbWlOSpshmg0WYt+QJ0qpzoLVcuTQ+1+YWGejRinhnTQNq+ozQZH7YG6KOe8XL1G
GPzXpco9bvcIv3bpkAFkl8Ba1F6th6/B8sPi9wvidqbOfOfgzNg9+6smOqErCj+7o/3CozVz4HQ3
hyxwJTrEdaOp+krXg/l6oGAx1RT/IOHwCYbVA1+LfeSpEypUEu69tQURrZiZHKlz33CTbyDTAykp
jZTTlnMhvoAuhIguEj2i9QFyQhhrgAaCm/KdcQ2oiKqbZRQ5EqbMyBqWaYNVFnyGXlOeuajFy4Sg
P4FLRach83d7DLnv04dpoh5XMntrgRXBjZiAbPQJtRP6uEsPamnrM1RCKqu8PO40v6rgnO+dzn9k
mb5y9iu2RQDm9T6o6EWPyz17Z1GsJkfDRrHVyQ7px4ZlkwoFHmbGQU3hG55hI621bx7Jv/H9dV9p
aWez1UvyXE1JPZqon3awAU/L+rsQQc/nQAWeR1yxJrctIo0db22HDBCNXjYVOzOoSG8WwLBha4SP
dsgJ4tq+dm+YtKuIfSc68KlvoRpS3AviuOXXsGlQyTzMzYeyP2tFK4kLjaJysYb/Hb9Nu+R32QiW
yb/wt4kdVeRrLQt1eSXOt8B7J6avJXeJpKAn/lCRIK75U9AepfaY+IfQXZnK6fjeVu5/KCEaxp1o
HmE95sy5hLHQ02GVT8Z1MY92vXGPE0qCWv4Bc7L57eb1XmjfOCcQ6IQ1kAy3SjE2fiYLcloYlYIG
T49dl1JS/H+zhLKla68pdE4NaNusE6tBmttcirya/VxBhDmCzQXYAFV+gsv1rWMtMIcr1KCl1y/C
dYo2H0EJZ2MEuF086VaI0JhfsQMVm5+NXyqQOA5v9dxLUYU55dnGumi8DFDBEA/Gn3m3JxxwZJd0
MsboRoyD9HlwUs10spD4y71XN6ikE/Jmp04fiG59xvos7W3NzM/MQTvuYwkAE/SyQGrlaQPawd/f
j3oQjoKBgfnBX1vy8OH7kOHCGWf2dFla7TAJHFsd1FderpYC4bw3EpyTLWowFoHnjRIe6xy4rafj
mnJVK8fUrtRPEeko10U80sdQ02uxIjH4TOo2IiTOXZ+4YdJVKhxWNHp/mWP6cdszMvoYt0kYMlSt
R+x6HJX7cl2l6pnhPHvc3bh50FQGjBaXbYqHQtSr5GiUyK6Un7Mumi1OfYnaMdj0m05OGneXOCmi
hcg7Y/tXVXMEN9CH2Jd5BYe/eV7kRZJ2jOfXvz3ccZ330dNBD9g6nyznbqx0KTD9Yh8GLdniebhZ
sS9iovOh3UQmgWBW265Wv+VZCiqGVFq++8HbJUA6hAyCA6JfQLFb582QyJO+xHsaDLiWUlIzBIfm
rwZSEwwar8T6GGDEPRI3XSnC1gLpXzBZShAUgEbofV1+2muDF9LihlsxgKPWN6xHPfAJgY5yMuEJ
AtLIF0hL/2mVkvTDzCcZWrvDANI73Ucz0i5t5WxrQdvJ4YovYFBa8PWyjcbRNkpCqhA+Jd40xWdZ
TfsBm10asvw3DfZups/Ryru0IpNwnMJmvbPhQqtrxWKrSVelsYA6oAfHIUghvwMr1IoyYDh6qqrk
im+lrWsEyA/8/AfKkZsE/H2QjMdRnsGTTX3PvInOS9/TKNKzVKJpREqnErw6hY44Xx0kIzw7xj6B
SXeOlJUzH4d4lrk2ynct+U2juCdznN+N/pVRDrZxuqaprkrY7PNmK+iRV8uOX+3k1XfX+ja5KP1M
1AoVpK2jRi/7wVBVHR9xXwB3+lxT/h3Ivbw15I6mueKyuZSsn0szKD0cK/BDUqkoHzScmDKrgXPI
zxKSOUbUVO81YLgT/WVhOroFDfxg7qCa/axkd5CxuOcQSvZvl08XCNsIinIrug+wsHpvQyecNvDL
yldHtvaL8no9fQw5Iz+5upNTFUJsY0gnZ8DFflOO3YYjLKLADB3qhbNz+xXXyrsLEQ4ud9XGCddC
uhENtwfsRkvFMGSySREGpLDj4xfE5Ib4k+bOBWAVMevLVZ+a6M4csAqOXRJLftKN6AHDlYQO5w9i
kVptBHeNOpelIN1t0+ML8urqozzd9Q8jdzL2zo7ay2tECiaipW/FhwXxXbVzy7Ug1UZRWlCZI3Zu
VV+PDtN/3Driwzfh/hovwxBHVosWbzs9kZ1DezEO2d7HHXihhuxGOvt3o+NPayWNq9atdRTflFIk
9I26kmvUxSLO8mP9ROaUEOnI1ezpMySfBRB5liyMKE4Yijmq0oFlAPIXLOcQ/D49uftPQgfGSg3Z
h6OH3k+3BuBwFZbKKw5swJmxUaaJU2hxlK1E2sfNbmnqw1Va1sio5z3WrM+cJWG32JmP/ohegWBJ
eAB0LJGu3CwjG6Ct8uV5oiDsI7VfKsieQkgMpdERo+MwpxszNp8TBZlBTeter34eByX+gghwuo8M
lv7KTPySxZqZm2TacHaKpBa0S4xIPx1Khwp8wrXxMIONw5IdA3rWz5sASjzVTKMLnQq4rtB6jVIi
VD3hBYi7jXjlnUd8pGJfHXDqGKNJr30sWy7IGrX6BMpAIO0GrH0mJiq33x4TVoeg82Wq5Ziaofa4
68Ea6IBGdo08cwXDAfUKSAZB3VI5vPcLYNXzKAmnaKk1dDnyhFsrC1cd2TG26ENM2xvmtTCjAsuf
mp3sNkCRFRzkHefOVEy0MkHKp4JvLc6h+uzhOXxagFliNxO02nP3L7nJwiMgtNQG5UFTmDhSJDD9
VB/z4zpLQgQbHTQb6AOSMe0uQZY/v390Os48FTcY6412aG0AcqSXZhdQ6pgSYtQUt/YlSuiX2Qqj
o1mPxVVDjgY4ZYm04ra13V2RvixCMIi+ld+34kRDPnDZB6jMDGPLRXDbsdV/q5duqT6zuUhQkMae
o5BqelaDwbNZYKDta5CGuua6unUbeC8Qg3ZJHmYKsjwbrDXZ/DFCzdswxaYMIZweIpSDtluxdi7+
GXvEUzOt73ATKEXEct9JY/Na4Q1pFZTqPpM0ksoZJaESYfieuI6VU54IrHodWPHqbhA/zUXoIN9Z
HjV5hiygrXddytUmefMTCer8kaY4OkfskscWBxislGIbTkvYEpebrIG9FEA70SGTfyNnXtnJT5JB
/7dIgr30LduHO/wYq8V03ZKLyuv57RLQpEEQu24EqXgJ5p8XKOYXJAvxsK5WzxEJeCGIBJQKm6Lx
Y4cZRBOJZyQWP/vpfLV+/gWh5FhS6DbXSPna82zYRLzHaRZNoV5SAzB+PRZAHoehkf9l/M0XeCqd
3V5imIQIMBHRwvVJ6rTBZV5AojekyEEnqsV2yM57OUxLv1Z1ijjy9wzzxMQtZQ9xbQmh/LO3RJm+
dTHOv6OQzgadu719UKjUn/6P4n3kZkBE2orWCm85E+Tl2ExZqza5yYqmlGszlcEpdznNxZQZRtl1
SnRLOqaJRzLqR0zcpjq/xwSGNF0aQNOFDAiWSL2znCnEwoIk3aMSKRBwuO7bg5De5UlSBVR2Plhs
AW1GKYtUs4SFwY9G7/Us+4bLinQSGMWqstSK7w0DI8loVVm0TTBSUxq7jeqgKxwQHqO+llV6vPYi
emH629bvjBFX/xGXGX0pr+Z4QOwsNupb7RXGRHrC3mcbJIzEi7JW+JKNvQ0WUqOZodh7Nsy5SLQ0
czJy5ezx6h5tEGAZ0mGZcCNj7Tp0WVub9kvJ5b/9qm1gBiPC+aR+3+qBuHFT/2dsOtKit6LNOmgG
mnPG4hXCwkaGgEPNmwnPn24XFUWqB4zixj0OAEjMra5lNJfuzsH2wLezDMv4Gfqnufa7qTIa24PU
yMKMr5Ne92/U/DQJ+fVb8GcMGeNsWfDeKwG474ROxnmDAPlJUSRYm9nLy+rugIYq/vL+2v47O/So
Lw24RYbghwgEWTZ590dMUxh5/STayml0CE807R8nGyV1lQ5oRf921nzMYbzC04FNn+MkAWVULV6I
wdDDrWWt1yjTXO3CJLfYMGyS5s7lO4Word81GVRwtg6m32mrpRO0kOAfoBT+2m9Lz/bOkJQUwoqc
Kv/okc+09V9vbEUmtqVqy/M86wnwNNhu0Vv740dW3C39BHUjOJxtRO3kLxfoFHLKzAix5JLU4TL7
NjIu1xsYF4XnFw55uilkk4dcoCu3SfiPDTVk525bsh5j9ALpYkayYSYi/huVG/4lTQFa+8rlJpUY
AMh9GhRWVkadAR6gUJ98nTgtIgfoodO2P1Gd+OOzwuZ/ohJvODdKRqnjE6GawOXkvyXrakE+sAc9
V/aL4RN9KpS/9v7Yfq93myE11UkA6b72CE/tinwpUjxqV3gD38J17DRQWha8+Xn4Dey++kkxon8J
ixIt0NpUIGGS1iEvnC+U+huWobnS/X0EHmaRvvoWiQG7tbeQusgPz7yaywy/jLIFBZxJEZ13byFF
lcSWMgDJ4iDhqCx4Nu1Afw7dZS2tzjYB4M6h3vk3zH/7+iEYP1XmY/dcX2BT7cKA7SQxmtu18Rzf
5zUsuC8M4NToKENCeaei7JnNyYWMcW6P83HeI2bVbJa3fidfQ74yJYawsTvM3XgsLBjoNBQw6QWi
7knjJAmNzX0fYxOeKojjhEKxpoTC43qiFBqrlh5nQQmBa9uvLs6WPKsDDApEq35YM8VSjWOOKQjH
CDStB6DI5bIUHazQlLPEOEV7W16hPAcrRRndOKTsxtscQYuY+JBDRg6q59rpo8ULw8z51zBVYloO
Ydl+ySBuI1jtq+ZHZWf5awBaemrvRMbVuOlS7+zpNmCB5fMFlr55+kt8SAZgkvmZjNhqsjL7g+7f
oy1ZwzCfPXN31EfCfcMhtM8VA/4CdEqthjWaOPUNK/sQhRxl/lUFFPE8Id5l9BaXsupuHvKIGgGb
ULLY7LMlrHVhIOXGCmmJHtlx56XEmu67HmZZ5KzC6VLoS+NyCaFbRUFv45VfUdIsQvSUVl4MERHu
avEDx5xZOMMVutUlUWjX9/AdBABYzaWUXQYdpH9qBhpOHZgGLHLkCX8Ekk74CrnUE/XWtNXlxB9q
kyqdfWq3Ey5YIZEmlTi2NBSEqQdiCOayA2c4+e//jqeD3vMgXVbDMVW7u1bc6aiNQuRtG927bnZf
5cmMO60MAI85mKo9PCEmetdv/aLFsyjZ3/DFsPi+9LWTPnsfftcAPJ55/YsAVDaL1ywHvlQ37veA
TOIIEDCv7bDN/CADzoxcbrtWyuVL7i8zNNCeVB/8HDL8JQa/TgTDsETYO15nSXxwXFllvYVmtAlw
SiY7+l/+1Zqyi2t0m06/9QUfXiNpbMjgx0rx6g0KtmIZE/9nliIMSo1IANkpEmFS9xojzxkl0yNg
yW9Mb+7q6c5h//sQGTZvIi8atJ9jO+v1haoBhl++ZESKUyjXmp3cMQaf+Xtd1awWq3BGbdW7RzU6
c2t0vknxG0ssgu1U17FmB8aK6xV3SjqwM+V3OJI9hX/i40Q4qfC+D14uhGngvZyiJbam0qaK7xGU
rCXcG+PS61n8/fLJhXFeudsAdfRwdJXsydLjYc25Zlk7p4/u8JTvupdgtYSPeYkgImcyIagLVg/S
cQQkEGPdQuYoXbTT47JsIswSJGBvfmsiOkrGBraFs9l2yycdwJNNRWAOX8IfGLoVE+hJg6ANDciG
dUjkb1jV63ydBEqFL+u12y5tUthi/wdumn41fYFRZS+bC6XPVre+NeZQPdxQdp04f6KDraHJ6yPk
iwAStfanRjrsgTw6IIqatWmvnsJ9XjiboMHZJvfVj1rDEQ53K8Z4z67sa+i7FsOzAv0PWLAS/HNX
A4aA+0EpaF8D0rXpcuzsIxSKN1h8TjcCm9oDXJ1dsUTK6/B3iaq1TrZolIYYP9htkkjZw+QpO5PS
czzQkXbZnz1SVOrpqI1cgFXPornQzPUW482WMvdJHN7gUsf6Jvy6mQuI+ql1w8WXJ3CCFJY2XhgP
GJ1BTe7o88/rouMEMXSDNzbaeW8XafAkZsi/Dz2f+shp6OIpH65cqXHmQDFY+6uRKSrwPti34vkj
T1SX1NvnXuHpcEdA8gBbYEr6oUWGu/paJKhU8r8MdmN+RK/bZk6iIVdYzMxQAUuvCTsurykbk7cJ
PvmVffzo8pbhbQaySlmZBFd4XsAMlLsYqbu/s7ZnJV6uPUEPVD8hZSxB5mNHsac29Ke7HMJZZlBM
I7UKUBrdW2dVOtCfbMiXOvx081gsJ0E9ft9i3GM4xQwAZn3P5M99Yua7xoXjhxrf64V119f3AxMk
aqyI/1zD3bYO51+y7CMO4QW0u3HLlIp2iZpP482m2xiNe/ngudsz1qEIXqskQOTzVftCPfc86YCC
Y2VA3caQXUMFcw98A/HwZ99V3r8UItwCrOtVA2st12Kmbnz+E3KscsgJtFXSSjMxoQcHzTJI8TV6
uf6STCLt2ldXd1FNeEYn8LGDwUftRUt0uDsYZwyJ4tX2ZZfKIvFHSLMd/3HOLH2HObRunRvReT99
9Pw3d2dCgdOlDgYLLFyD64SaaPA+LUBw0/MBYZ+ArsUcSUIe6Psbg33Lml3NrsG7JVf1zFK9qsHJ
PUK55QGAuYkPtzxP2zcvKyU1ieqxUXmAn1OtJc+Jvp5ZiGKHIl+r1TSDwomF1YnT2AY5nZDzuM1N
6+kUcoRBkWL50iEoDcjxlienPUMGbdzk6HlTvsKLv5P8v8yhWOaODtUaTBa9Y+a65zxncWTrk5d0
YqeK7opO5+H/9t1l7vplH9ZPgbC+fBMopP7I01+HoMdHXnN5AjpWtLoAf+VxEIsB8PvxUjzkAu6v
90JH8yhCtWWilwXXNIAiU20aZDZ3M4jbVi0ML00D/0BzDtNT7CN0Ii6W4eVGLObBYwhfaygahpvA
yTaTQtaTDPmJ4PIdlJTOYM3BCZiaQ+JhmK7+pNgMKwTDPGlcTnK7yaMaU3+u5TszuFmOiEiRvwpe
YyttZfFPo/mq03UHRdgwLzT2X1XYsnEHZVkXylVeRkQmXxRqKaasLJIxJGHey+sfV6pnxHJyHW7S
M3XhIFl5Z8xy0BmiSbIdUEyphpFHnbOgdSOalihPQOcRcN/1EfdrXplADd9Lf5KZtHIlDLDKDc3w
h8ixqjGQ7zCTPetC9L7MMfHms4QhFqIz3d3sUTZER+pMfIm0oMlpXDrWRzDSBYz0Wi/arp25kqUk
4C/8GsyFrKJi/ahErqUb2aTuJG95D6YfyzoW6ACik79KwmCX9xNfEeZZbw2/ZtVVOX7JgY4qL6QA
80HIgp1i4Ukx0tTXIXiCaxCLH0YwICjbb1xX8v4ogbZ2P/2KXtGxrp4mBLO/VJUeR7efFQQQvat/
F6wwDY6SU9Tz8sm5D8YgqXtdD0xWNxd5sKr5VWZ0S8SKYRbSMo1XBX3YyO039+npxLD4n3W3jNMS
nj2c8HRzRwuPGtZ5Ed6u2ZeL0F3kv5KM+Ht5QqUhJqcQNtzDKRRGkVNor4pYlgeX8ixYwrXkfryk
Ug4wDbe0CZexnkH8+U5omVKRfB55OxQ/dKLsMROkGtJXqFhsViGg+NDEyn4kosz2jySrt0+8ZnZz
QynIy34TBkAFy88ldkmyJXBP4fRFArfc4DKioL7n4Pnrqj2zHphjmlouevrsAZgjioaojm1yMkWs
N9+/+lHYXFh3NuFO1S4dNfGs1kmfUNop8ppXz+KrFn/ii2OuSRt60MbiH5qaFBbPX6sHbqjEjqqM
exyuXVttHT9EyGyBd1cmyx/Uup7ZeEeLs89WkG/jmIgHvlbfw6v1/z81wk/x8IEPM5a2vTLo2/j4
YAau4sDxjicCme9oaJeKTrYKqUsAZSp5Mb8znxoN+uEOre4AoWvJoJBpW65As2ASnu7LrkkpaG/I
Vq5SZdZkuE2zTKeEJuERgR7Mh2z82cOrbg+F1fUpbL/4zdJXTh1cKRGvo3T/bgwisZXuETj0iE5k
Mv77ly2jEDwsUZtL0Dg7OS4ElQHqeWOX3JlvLcj6QVfIBRV3z8dxz9EQfUGRwi8AC8liR5zkWRcf
iPw69m/SxfIXVFp6yZHWApn6QTgInoDqBnHdi3/d3dEjJ0xz1bhb6DdK7Dvl0eurJrwopCHzsXkV
CDuDkE/GukdrLkdnYeWfGQ2GcXe4XQVYuuhEj1oDQmu5SZyJjSG0z5ln5cs6WTE0nfaq2ARbhGrp
WpJkUUVEOGhavoE4VsRx2isiEUU0UyUpIUVB89+yyDiAhx8Zl5aQdYRREwRQCLqem2t0RMbllkVs
BqrtHmRa9Dcv0RK+rMmkgR22h6N9TX2HTQ2kKvgQeC/ed1jBRqgsDVXEm38uBSkOjWBOb6SS0Xak
qB5tNqb2oop2Ru3y4RoW80D2JSCJgiNdI0wesdewwEI1QYqdf/oOYXJHa1hGJrdCJbxYt84ZItpZ
0rtuzfAYOHwsIq3tVBAxHtksePTQpJocGTik0Q/mROL9ALBCMHOt5qv3izYHCzjuEjFTrKu5vixX
Sl4onKHq84TNmNktO/PZpqTR3NcSwP0rvykusxqnItfqWGJrbTDdpbv1N2s+NRMqIImA0Bdh6d77
KNWvUdD1ez2cTc63bcpfdqW19gc/P84mHDEZR7CPeeIJqSXHotqMJdYKABRJTuIKkiZMDRGRqtyl
L69r6ui/kQ7/t7VH7n6qP2a/ttSl4LSpzviLeum14VKWAMFD7fS1G37hT6YlmTs5a1pvAyLS1+ii
3Y6DgPR8YghRWzy+xoIw87StSHJTM7t2lGB/FAzIHmQoBbq3VOG2qfEfVdydf96O9N2mvqzCpxOn
4vGrioRQuro4aIvDKtB8EYC8XsiVipYAgSgGEksd+x/SppSaR1+p4Lpmc8kRoHiELmB1JqeKD7li
Fnbf1K2R8Kw+WerbZStbGtKvchKLhhHXByXJCMVgxip0K7bVQYbPHYaDro0yZDW/HNlpeK46XZwd
+1uP7e49Z/x0DLaXB5YcbGGQLQTLmrXlZe4Nl/Rrccc0LsepZnrxuMek5jnOpy4w+tBH9eWPZQVI
2JuvT6L2K750FOpW7vVRceMh21g6MQABPHCHSM5uvUN/b5fhJK61/oZQZhDttREKi4mVPVTe9vEQ
RY+W/CWQtjf67mr07Sb2fcDwVXLSYxHpuMJbChPo/tgnmWnT5NQEkDHi6qhf6ujLDgDC+edYue9A
cY+UR52UjcQkxNSYg9MG5tzhYsRNTZ8iehzD05zdpEvt1yQ7K7QiPMREWGzViaJCyc3QVK1DhQZf
bxcnzASjd2PXn421LG60YwFFxS/Hv0xOX6XralFcV+9WkDzAml0duhY6QDI3FLh2jg/bbb9tYltg
ugVfc1pFMicm3mCesXSVXiSk4lpPDPuY0g1OCLhNvHfNHjvP1uWz/DqZDle4uPkblgmA8GhK2k5J
V9KfnIpYQxfzWuN48zv9zBrQXu4poCaO8S/lnbYYQhxvaWIlobJlIqPn/87NtQB+5RFvBesa5nqO
yA9AWgsK/J1j4NuU1Qo/mbYopY7btNqQdC6qdaWnTUAYA6ekOLxi+TZJI6Yf7aGqvENWoPEQGYX9
y51CKV6LHo3WYaW8m8jNDQ3PW9/qy1IykmMIc6VJYz1zDTgA8IybDDUj6/IhEu+d1hLNmyxvN6By
kGO6MXegVW3jkT2d9748f0DoF7/gTEFkbl8G8GWgJ8c/ya8yAZgNNxzh5cohkfLQ6c/VzrZM87WX
9MsFrLPou4M47Lg3/BAzo37hfMduZOA0nQp9NWo9pwz1W5xQntWUyHum6MCNUFLqiQNfajXGkeML
s/4BT3uelkPNK4GEVb+9lTHKeEJXqkK7Vfw98YBGMPln4oInsPsT6G8JLJlFCvC6nMLgm/VNf021
Pp3WyyXy+T5WCBgBDJF2XYpxQ/UJRoL7nEmH9YhacAmT2oUbZiYcEq4WIHnha3J2pSCfcLlz4P6X
sU5z2dCmXE5XbXLGI7rSLsUjWG+c9HrufsCMKnZMW0ju1hUi0tOqphH92Lg/sUYx/9hNYkgXXb7r
JnwZ1umVrw+nI4+66vg4XwcWk5EmbPPKN4cyfdHHTC6sJj/SsQmaZ2CabtUJtqhuVndi/ROUKUyK
jMCrh8UYq8xGEtbQgABQ2u4/IBDPNhkkcU4zrI+5o4rlMa0dl3nBEAOx8TiD9IFgD9eDenFJhoiq
UiAAiQi7CJ/md3Uc2SuzmQmQ7PCVc9u7qqRwcH0B+v9rZRRKqlhTas6D63S5GmedpKr7ATF+pJ+d
F9+GyZBICoJg3XdW0iXby3bXqYIV0nGbV6/tz66voo5BWWIALsXNzbRqy0cSV+/b2nSPkAm49Eul
pTAtqbTeoXUom2LgTlflyskBEhRxvu+VVrAUbdQCApEaSUjiTSRlk4R60m/Ddesh96tXtRufdTRq
ytSHW3sL5r9DTaMAUAsqbhbtH0UK/8vWh4tuVwOdLLVyVCVGotJmaJx/AuP4kYxIUPHcN4K0qTzn
ysx2Oss0kzb85DQpeoOkKnY2iU/lkIfscGN5WyPyPA/ToPdNkNTNTyfO8MjRr7bKJXiPWY+7PUTf
eC1BAWRQClDU3lSMxg21107XtIv5BGVVJZplZTmJ2s9sEgz+XJBIhc6WUZ4YdU/V0cKQLpdIUBhJ
BMyYwwB6XZ2lfspDlePmitdn3Wny3KNhzghKZ9Z4Ndu7bznkanhgVdIIxK+gmg2KyPD9um/U1H59
rzpx1H67uIcIjt2bWmPD2Cp4FB5iRk3/rU7yPSWs0NuAdeVn6GIrZ2wXsiMTxMdFY/2eR1pyVJzH
uiTYFx89vcYZybPmb5/3siRUACcjQtg0+bIY5pYGG8sH3tqgNIV0rYSgVcCRxdOMUb8IAEigPzsP
T8XVqcl/XVsLi1CKXxDaf0RlXyzgNIboio2Duo7/aC3dIsEZ31SE0AiG8Q456JBelPiyj7KQPEnI
/tjWULtEZLma06KpyeLz4D/CrG5TnEpZkOw7r3EGCgHVE01XX2XLE7meULzYoSQ7liTCqA/Gv6x4
DynhmWZzee+jClqY5YRs++95idrCsIcy3ecISpEOofzc5l0GcG/n9qDXTNyCDU5V2+tSJouAwM6C
Ldx1yCAq2JSHqZsYNYveyQ4af0NxUGPfGZsxttOHg+1Pj0ZjHR8LD8wBljTNm7R5cZy61UImn5+3
t8FgLoSLDY/rTD+HSS5S46cnCVKPy7tdGBk/QRKe7rWCBn5nhYDcAJOZv9A2P/DXIolEwY1tXY7z
cvNGNSdjwpGWZWWX+bWkyK/cPmTWQ3ruuUFKPR1wcPlW75ERAlgBAl73xZw3nhwLpLJLBbPXIzEV
KSQf05mxWcxjY9M4tOWxY6zJ4gtPFSaAT4lpLByajpDFiRGlrBZUUFz53Z2xGn4IGhJlCyU6Lh7n
+eN0OKRlNuENKieDVjtU9w88AS2hbu+TcCH9naeZ1aQKkcvEV+eE855M8X9t9sW1jFplz8+zyaGI
PoTNr1R/b7WtRdD5U4yiiGaTKZSSFHHARBC6tK5ZKPt6cqL/wbfXQ1a5tkRjdraBhEhugeVWGm95
Hz7Xwdsq9S4oV8WA5Ya+Y06Yu/XwN4Pvz9qMmPEQik7LBGVYpsxiaBBSh3bFI+b9Vb1vBj7xZZ2w
adPteEwmjo1FJ759ejA1I6L95SRy+4aX1HbK7YGbOuqSxxms4z6aOr/z0+xtpvgfDjpRViYSYAa9
h2HtUJ+HYsUkqBoHwjdcHeVAySbeqcW2uaYgvMpx0TiZNe3nwnX+O5aFdStfiZQLqWxI5MSWJq6j
ot0T742a/LlTzBGZm8ocz6T6RaPw+ixcAL2ujqYzlaJuzo970uPFyTHNQkG4GQIxjwr/FIBLkLVL
AcKJ0M1a7BPzure0+F+61TzSKcxojDhTVyzKi5Jh2DrFj72Ctc9BQPG6SNsR7ZdlkPkrGRVpljyn
5Aq/OIHBtZdwKbnSvtHTAa7Mulh0/TPUmFKXnY1SOY+Jq1GPzNtY+1OlEt2j/JOboh1CIfGZasIe
YH8+SfUG2+HP+F+hBhx+O5vJk9cD6jzHei4+zQw57odNnE+wGpkFuTT+yDQyW9pOiyR5FnCAzpaK
I7Kt1H637id4jenXNRnpdFai63LHt58WVFGv9HiGUHLoVE6DXASD6UWoS8k38vRocUEO/Mj+JDBr
Q2i3+/Z5meF+NtZY5C31Hwv9TWKgrWlXSbn6po+lS/x8B05ezppIC7Xdu1oqelZemFxCECW3Ns/y
ciiXdd89RFhwXDOqzG5JSs9LNRC75sOyubYiPaJUae4h5w2VRm0EAai2qzIFi5XwM6PmN+r/48bq
TxymJ8ijlriA3VG1NrNB8hSThVwGDjpzlPetDQb3WkEX9bWYCdNaIvrcTtmiZot05TEDqjOQ559i
92as+g+uq/Um3OTsS3YVhGrR305+pYy1TshGYpoayw8uTUFIzTZBVGa6+mYvwwGslrpIUeTqVp1H
M0h18k8mdM3348PsLUH7mINEfjwZ6zY8pQM2rtIRCOWXDXBgoimPlCX3iswYW+I6LAe0S1294xeJ
/l4n5rChmEQ9/74bospnRjq//Hl9grrlZTamnqsPc3MkpwLKrCgkejlrJLUeFttRmBKm1R5ZsNm5
XpJYaRGWxvnRaiYqvGNPh9tf8Gk09vrlz6yPbZTszIwufkr/W7v94a8bwnYg7FkEN5tvH5n0YLLz
XiqV+zlmqe0ezlKQiGgWiJg4rSnDP2VLBFhywMPwTFtqwONa0d96Dhk0yHU70WiAG4Je7IMoRiJZ
ShizpvWbknooGaaHXvOuyQUEX7+aH8xBlaWoJGgCDuuBZFt7x4K9fUO5x0keyQC1XVxV4SydyDEy
bPUSYTa7xX+5DrUk1ji1bsV6s57Se74Lk2jHEPiBkczGQpFfT2cv+acF+CvN3foTI6/u8/XwUJSM
wfYVAfoyEkLK8zTJhNxk5tyHBw1L7vCDygh1GTKKvWGQUQ48xQnz4Y2LbMZSmhwcgDMd5rEGPwdL
6g4XJtejltfCwggt0ZkJL4XUypstTpz1AsbEJZ0I5yFKo7WcaepgGiW5xUgu49Ujd/trLLGSIbQA
ZKaih/GCJo+Tk6RJUqWMKLUDW5FK3KiUaYZqdKbBjEab5/6wAPVX8p5JmnY2Z0tmPlAKzz0cR6su
+1kV9fxJPwSq89LwxNQGFie2XVfBuGj3qm1k6zPMmvGmtCtby4Zwwk+Y/jFoX9E4VDPQ14iiUquz
5T+zs18eCkpwhYzNwZxjVAYpo4hiCueXPRbDnurI7BfOUuWl2P3Hp/GqPskUirJ9pxwNFARIGOx9
Uetz/GsZ6+Oa0IO3rfjHVQbLhz9Si9Y9mdKW+SdQCJvJg5zbl5ZYgAwdFuAPf0nwHq3RVSITP2ba
TndVGQL1HGruvsUMvuNoS0Kpr+6FE31DnZ7CpEbKTyxEEhQo1F6Gu/kyhzB731TqnU5YhBZNgxHy
XZls80XQDzPJfPYkJD9rTv4QF3m3GjBC3LftbkCfFCfcIC0srI6Dshi7d+a3fpKb1NCbXv1H2PKZ
soJmds4Y1vKWjjZ3IeRthhM1odsnSjZMwF+Ff3bljYbT3EYrxGlV2BC99l3II495UCGeDjcFkS8D
9EzvdSUP6tifeM1A+wfHu7FHYFFB34bZePstk01bvdeBC4v1yf1K/c1cqCitRMKlzccTYsGhvVey
LAJk01bpkjAc3NQU7WrvNnGKbgeG+3D6lNJqXYa6iuqw2NNM+HhrI3kUKW0RZyjs+FIFDbhzcILc
4XMRUSADXsFvDOHXlQTR8DKq5yGAT+Abl8WJvMPiXSSLV9AzdV9rDfL4sb0L4FpeTDCa41VLk83r
rwaLUCJdYlbgxyHc7R6xJnVDZ/UFfNbOTyDCrwBjGfgtE46hS8kQJK5b/s9F3vcL5FFIyHkk2K9Z
/aHBdnwzSWBDw6lXWfnsxIbxGRu9n326R4JOld5fgs71LXjVDFmAVxzXUMDCN+v1PAWapX+w4KoR
owGq5573FpIdL5qgJsbZ1SaEO0gRLFO2J83Kc5Lml6LkbRTb8ssYp43QvAJ4NRdYh4jLKvIE3fXX
WTn2JFyz/+YxDn0j/DXZXb3VQ8C8ffFR3mcmJrw9l47Y2rpA1be6V6bb1kyK8WptSpbbZqmgVtVS
CppeMOvwQ5zisJ0ikWWdfs44RJoQfzvT6nMBnBS/KR0CUlWDZilZ0I4eX1SyBBy241Ko+rwSsAAC
WA1xI/SuVaBCGqNkPh4qTqx9+XLkfWxDT9ijul5FyblTm4SKFqlCyRski9H924/F52uofIP6vPnU
mPO170asxecMZjGAcc65s5fo0fSlEa5m33ZIiPiUWp+eu7jp+PdQBSm80Lu0RsxLWyFuK6ydMkKZ
Z/3Zb41J2u1e5swLEkail/Ysc4IBs6fMMOYnZbtzZu+Ly4A8rKJQ35jLStut572HGIa4mlD4vJWI
nzasagfT2+mIfjtWqpcw5UgIXUQVpRx36ApjAmoceAIhJpq2S0ns7WpmKpyNRRUF612MsWY33lAS
sPt+e9CQobvEigMBQuqZG3dZOer22fusl46AVHUc3K9UiKbPtGdcRmhxcesW78LHNlQMJHleMBmJ
qmcJubcumHYTxisY+LusBKBBpLQFSrzzmkxduG/MCDhm5eSJp+6xfVGkTSI5Gv7xuDztXNajgYbd
hnN2OSSpwQtIXW8whzseW53HXgirfGfWjgQD6e6kOZ4ugwdwwW7ZKgbct7lRcV/F5PWyjlyhC+4k
XkKhDRJxo4ObAYB4tcy66XziWpYWHVgwRmyNhYS4gDp/11FEopW9uCQMCFMYqOKN/LrmkXIQ4R6t
a+SA1uagzZvv757kIBiMzVU184odXpRmHDIrEEVNNAV5j6PTR7nd1EKEQUui8ub+x7YSvXFoerX/
wEQgdyZTsYrHn20r/kMc/P1KQPcQh8KOrwdL4kR+/FRFU6So5BtWHEdFwEO0tfjfm6nhsJB8dumH
TNNZttt4RUSkPr3uZr5g5ADbRZQBS4pKfPawf6Ocmk7V7lE8ani6wM2oq2ZwAyEYXdHPF7KgKIv/
8daitv2GdizSNyqlG5ulo0FuyGNTpjFil0WYDiUFjJxp835MjO4/PE8ZZhbm1lsg4YT0FPSeefFP
LEvBF7VHflPx0YtNmNSp2HWP/UADZ26zgmXvo0rIMCz62+NSvK8gvy/ax8winEnjMdJBp/rwJgsS
u+RNG2XnLms74/HPjGuU5uu518UkNcw1U+18z4NkC2JPi+hL+Do8J9SZYw91gxKaLASfsMgaIGwD
2hczAU2esjnRmmxTsQf22r/ww/42SYPPa0+H8WBCfA0xfRXP2Aav5nRUahuKxDPB7iv69InTsMle
Bs9rZH62gJmza6QdLPw0/eDEwa1KtNFWlvD+gZAwOpBlbzEPbE9QSj3FpjTBAu5L4g0P47jBn9Br
qOYZWD4V+bQEI/YpNOTQmxz6P7tTwEw3s3DsSVsv8uJgES6/m83kYNrW+YrkgVrK3Dic1Z/TaV//
StB6jw6ZTT4UdHL3H3i8lOhSwLG3nUH3gj+l+ZjpW3jcou8q2+SW20xucvmeaggfjP2F0lgWe/na
PdHsC+sMRb6gz9AAmKHw7JTCiePNdJRaumFMqCi9LYzgBgCGt8gGEaJfkAapzgyc4ZiIukYJYKg4
ZwMR80ZslW55ImY6773ReCgoHNZDTGwYVSTYtOoOShiu5J6opRRc2+JqGZ4WksTRHvq7Uaxqi8Mq
lHp1jVCjUQOwXXonJGVXpumbXLKQJ/v+pDNDfYdno8o2Ewe0KIItV0SWF89cNwN5IHXo1uIvNDxa
6SMuV8YbPkWDCqqAHbgn1HpZGf3fM8E2A3YCbhIDbJ3UGUDdmncypuQ/nAtK1+B4Hyna9Vu7AOsz
2aZC29ym8jNdDLrbnUdC4rRdfJndqNY19AfYQNqEuuay/tT3JCuQKcS5oUUz6x+V6iLG405cseBU
QrF4dZY+ZkMEOf7Ep4z7BCK4WJeU9xkQ7ZYXkwbozjLdE6xR4p5J2qrCyUvq8RetpqcasDNVOML+
/t3WTcF6G/zA1U10U5n9su+BtBsb5CtkvaPWSPZH2RjKx9rOb+P3CKAJMRtg9KsKUSCtI20wd52c
D3e8JTRlDK4tGnrWkgorrF24aWfqWivZXHUM88nPfvEUoaO4kq+XkjuITfcei2JODmMJpT5AGSlp
j0Pu6CJxwUOpopvSVwsaxI3k6N6R9n59CUCi8aTzx5p25qBV1Pn7zKIHLGpOM2wiVqz06hsBie7M
KzjtX/tM5cIXYytJvSBcIVLeExN43nnFs42PqKFHeAh9z6Z8OLb27HGPDjNYwAdijkAc4gzSHFNh
o0vSUW5j1OOVy/8EctmeSypd3QcB0zSYlZE7iDNKmexImxcQlewI71a8KpuTtzks//O3mtAYUuYi
Rt3nPWckcG41uZczixF0aXYQYw2Sa1iT5p+HM/YOVgQCmr92faXvVhdy8fJkdS9VPMO0aLG5wSr/
/u1rpEGJeHovUtPkKkgUbA3LJ+S1AOz3xO1S8uN/eb9CSHtX3eJhXG2M1BgGyzXsYD1yUImxGIGN
ZJ2kxrDY3dj1OxujyuIT++tNDDT7ySQL4dFlkUDx6lvdILbAX/8h3xgOmGhpQISUJ5ynOZro7Fjj
ehaToH/vWgslwgY/1m8fBMvAdA1aWbyxa+K8T2Vim6VHMc9XwLpAV4702iEKAFzcHJJwtWuojEi6
L2EaPVkEyqK4HiW5JwGxxGHYBs3ztYEck8HZ9O9xXKV9BIeCZjVUKQrdsihfuI7HAYRi3yOiNt+u
aucMzOMQ3GGygDi3yZYenBXW9ClrNvMj5ZqWvO1+aB1tllXMjJ0iASgAbSEpl2TkUVBBccHtlm3g
ezGTJt1D7Dvs6QOXmk3HZkUCMD3lu6Yg0uBSwbyWQ4TMOsCCJqne9cstPuoO7HtJ9DUOkbqEk8zg
uYgntARXiSjgdzoxaRFxb324iGY/hPgavD/86y0xHQyCA7cwaB/nhRqx+FyxrxhsPLRKoON8Bq7E
kyvPgwYJ7xpwsHDCvftL6hQxVNIDpvwbx0G/yMujSpJto5nAHv05kijW0CJieNi+Zbpn1Q7Z6URa
N8IkQFnlYTeyHvCWn12YhXcclXREQ6QKTz8xil5tMqjGYcZxN4xE2XGYSBCwH5C8UBXrhem/rZm2
4963yZn9xWqNcnSMXIY5HiuIhAqCFTmqi8lb8VOd98HFXBVKrhNj6uMDy7OT1jV6U00sMlyaw+8M
aahuygc5KQZhHR1DxCFlEHPMCIOadWDdUtk0iT8kFC9XR0QARNhAIWdXsm+mFE4449GDx5LYpOTu
ZG9wp2Q9onvpzraDVeEWyJ/8cMQmP/pikj9j6yathjwkr/V723CcnNH0gcLWd55FTG3To+n9231t
RNKNKKLmwTT/tkTAtlWhnixsFSvI3McdJlvjzQnuG96HvaPXHjIFHo/L1wpOiR5Xzsg+0Hwsv/ae
GoZtKSBUznqZX8amhM6rsLWWGOl8Jd9KxXWX0xcxTUO9jAWPs0BqoOZd3KMOz1B46PUXOOfGUeYK
XmY8CjUcXrB9Tkt58AIA1O4v1kcyKIuth/Ak0wR/8/xWLXPtFxcjadK94JFBOOz6LuwInycHk7NZ
MN33PBwymLTi+y1uK/DXXdT3WhvxsIKx1N7+mgxzT5MofEdYt9dn9GG4KpwyLc46G6HPMCLyJcPL
8ohxdRa5ecAoUrPrsJcQz71kX83OrrjrZaPoYMgIkHBWGc705i00Kb+N6iU1upUYpzWVtIqQ8W8q
xWEcVfpZ6sxNAewM/7M5mXsg1B1I3z2DZzy6/2+hHUXRQDVHbzn/gAOBvuoTn43ol76ysL4vbbn+
myhn6sQNZ7Y3I1cBLjm9FR2atcpyr3EBCg0V6WcY6WNxX1AA76mfAYWl/Q2NP4F6L9hyA8Z05Pz6
tpyKkWqVPa2TTdR5XgUZNWn6yOgPmOh8AvAwKOg2ltjZ6QCQ4cDZ34ZvuPsNKzwiY806wA36B7XT
mvvMfL5CoHSg4+kUwBu5SxELtNwzxfmPYpsVZE7v/bV2T0I0+xhqdJho4PwLvYQ+gL7/5RbcKRXu
iG2lrQqvL0T6jcenuZCCqN+d0BEiF+6IkyuQfJBdrIuyXui/+tHzYZEo+PyoS/t8fqK8aC4ox+Cj
vn3MlkLNPAtOVJStDBIEmg+1mghRKvUys/FEYMwWKxyyC53vwmlK5csu6E3QBO0zvxlir+SRJ1rm
ygqKD2dfneicrewUtbE3bCV7Ipl7KtCW1xu2kcpikIzOq76gywHk0aSTlkNVsqT+e96izFj96b/c
m5KFxLTJMCnRgAH5CLfKjWvf2H3jYTIChnV5dwANsixemtNtAzcfmU6w7A8aS8SE+JLFR7KCH7B/
gSVq+Vg8w1JHKbp7Hq5d8d0Q9xo0Res1ixHy7TSpUbq0zzxax7etYy2mvve8aCT5xDumxuCr2hic
H6diZeC55qsNV3+fELTtOxeaQ9MWb33vr54BiOhVQrDaa++2GRgUi0gC1EPB3HHmhGi34tmkqQ8I
chRRx9SvNoMoGtQRm9Jdkx6Z5R/IepgKMIe0NxuVgYYo4Bi0cSP8cQ9gK5UfJND7eBq5S6A014A0
0oEzsQuerI016be3Od3ZXBK8806SD/MRjYNf5C/gHD6LKZIwPYP8G586rHAoFRF6reAzNTdED1ZK
q5FoWHX1dNjD6l7ij8T88FdAFsnGrP8bWzNOtrk1ufDM/HYpqOxb8+KzDICFXMV6W52xsHYSKTs5
T8MJSW7jo8E5neo/w5QqJ9chc8eHaLYSB/YrE/oOpuSFM7h/b2DBduB1yIPnSwauJ482EYAt0ywi
z1ex+iTU/b9g2Lx/OGG/v9he86y92xI10duqLl3WRAOvuEP+Rn2YG8Ok5U2256LaUrwyS9HPltGF
l+8+TPtd7sfLwhdLmxHN9+3w5eW7+tBjdiwL9VNZUo8tO+Lf2UNKchB1zH/fhpQw1fNagsSwFnB3
x87SkfyHX0dWFZGzp63Rw+p257iU5ZYwk8auHdJqFqWiFhAz4omLsTF5I/eEcRULZm4Mm1q5bvG9
YuRmw6LG8xg1orHN/QmZNoqZoPgHtQMFvGbX428E8mpt6CqC0uJWNHIBtuL/hK6VoyurMEkuOFa+
lotclRGnbTC2j4HQBGUdS/6nOJWyzrM+FbcjI1u9eYfWPNs7i1BsDJiplnTxJ/nTf3Eg6KwQ7wsy
ZDJDdYCFMxMYS5x+rmrFR0wCTLXGltCFOSJuau3+7/pEFZzmE4WlAUYTrqzRy8QF24LYNCRuGFZa
Xfu5Vf9AJfKYQ2bdWMddzsIVho457ex7y9b5wllnBqWk69XCTyyq5egJLdUoh/FthmAmlmaN75ty
PxAu8YvIZCxik2IKMJNlK501YlflUsmBAUPxyk9NqdyRbjDk1qlB2vN/ubw777aLgkjaopsT/YJ4
eyIW5XZNkaH8XVrAnc5bGS0L3BsHzHVFVncMMBy/fK4+238dmuZu+hUVtRScYzorYt23Qpaa7bO1
ZRwiwVq+Y3oc2rmU9rQz09FNM9SuotXcItwETb1Xzz48+tXjz3UMYyWpyfj3iju7T5SOvgDRuye7
P1kk1gM2zLROTdD9BfvUwPSEpw+PNVpUJ84uj09SPFMtMm/sWZ5ssMXFCk+Y+P2R5+ibUnDSuVV7
BleRqBbttcvYT3rwUe4R0qesy7RlCgD0lkHZNCvIZHeqq+ZqTuUz3Piz2HOAefzyxkK7X/iQw+wG
L6S0w9Fyfg78YCmz/XrYbmjRIHoz02apr5tIIJhHYG35yKnMmouJxI9x8P3fkKQeNy0xo2MRi2ts
vik8Ndj5m5Dftr2IQKpBCI5p4ihenPLSJPkPyf0XwFmJLw7p7MmC9MKe9lt3ZFCe9/BsIGa72oI7
Rija5P7q6sL/WVUDZ26S5/tyh3cXUH8f3kHB/vwMvtwo06FcjOEKf8Ee6E94uw1K7uR8/0OsV0JP
fBlvVuzN6ZQTP1pyH1N0vUmwraRtuNGjCpm5MXm9bgOEB/pp2Cxsa7OcMIgVNxZVc5zyOr1KqSGY
HYxz6zhV+KvpIbjPiobvLcRqX8tFtYuflTdIGMjue1k0NNFGk00uLNsGhJKY0v2ZUh6vvNgKNRSB
u+BnEYy9DOm4MIbNY/LO+TjsRVIMsztTIo5+aXTbkpxS5++TMTAr49//9DBmjfhVG4YbgHbf6TLG
5RDU8WcxZI+40Bcui0iG68lHcpGrwNMtGoP179tYDXGimDNvmo5fGcjEg26ghA2CSe0mQxpzW/5t
p6J7VzZ54b5lgm2KreEOARiXRiuwBI3HRyHOl+S0lT/hoQ7HmUusbjNOoC/3Ei5OMegf+ENEvj3A
JwgPGIzqb0jNf/zq41Nn31cc4qFE/FbmVf7l2CQZu14OE0jAdvA5BRy+YKvVdQuf2w1NvHuCEAI+
FoXFuWFaoxTmZySdtNQIhUkRNEdMCzr+I2vhOhnlyxmChyYwlWFcxJgep4Q1wBg7eHt9YC63qx0n
fw5PRGkrHRnFLciwGbbhUrYcLN0iLxghrXN/C7Ux0gEStJoFxNMy2neWt7zQ37L6ei3ZWblQJled
QoJ3h5X0f4U/3FOdr1IBhu3gcYlst+dRX5KydalyTIiFUtvZ8Sh/mbzUTMsUj7/UcSj1SeKY33dU
mXZPQ5kEAnpf25kQ3RVDIvtxR/qk0/sWxbW2dsf9ClVaMc7+qqlndT7DLn6jMgZrW5vpCFNk4I1h
PUKIDVxN8jCP55hR6JHL01ppBE5zKYuqGtCYSTPDbnaq+iI1mtqxifRoLdAEK+kWvNbX+RrVhqT7
TElZIkMT7KydvXb/KxiuQEW1xyJftZ8WHVp0DSv6AP01wc9zc9l9mQbHtylrzjq+ko+uOAZU1Y4M
vi2JRuZHWSfXvVoYNXvtlV6TwX91GIRBV8rRcCHZDFAk2m5vXiJ70b6D//UxxEUFoyrTOhoXlJ0m
lmZ6T2z3qHPiHFV4BUqc7uRWHf9emY5xH0oDdvRioQMNC1MMJuo9JLvP7F7Z+gng48aWtg6Gw8J6
TNgbC8Zl7FEBNIf5g+LnPIue52amLeOd0gF/3qCrSUp7cPzcss2GYefXOEOQOpXN+qtfgbx3KdvY
0AwVUO6FTMnVx3Cx0tJRtH73rIB8ealu1WX+5X4vByI7PcvpVUr/uXsGOoZls/4RU0rhCpQrtqm5
3aB7TOFNU6yIkjbcyg7jStddOlR/Y0I2ZDxn/62+jJOaBfMJ05MXUWGIkhbA6aUrm/gRfhefRSaU
DpCxkqZpx5xbfXdigxySIJZOON2aiqzzKk7EjqwTLd/QtykDb8yI6QL/hnojAJYbJ93zK4ctqWOg
S3DBxpwUZ25LA3qslCWqI/gQwKcEw8QSoumvAi5CUx7ZP1CpccZD36TQfuHpb8kSv3cHXLxnT+Rw
qzsiKIQcvZMvyjPGD/jI1Wu5BQt/exAJx7GAbGdnD1swE9e41F9Rs+KQu5b6nIi99Y9bvW+9Y7VH
a6ORlHgvS/skaYpKYq4zw1I/2y4u4SzIj974gotkkMtVbGY5aFzX7OEaT5b8Gu5II5DhUjqkmxfE
id8Cjh4noabALAJkLzEfKshUp9okmnd9TK1vW5QqS8qzwYRlTWh6bCLj8CsLomyJ2YNz4eAJeOAB
fkqodFxVKxWAMa7uhAMMKbqa4r+OhEBbMCHWgvyGQwxDBbrP63RpJjwL7vAolbsZTeIRjuRMrxSq
HjiU4lVcu23X1mLqgW5lX3Y5s2jOKbjHj/sdD0nOPtfc6tbXv4shzvlxAiTGNFlWzRFfOd0Z0ngW
FIoDUXq5k+5Dh+OIpbROK4DWodkUo1aUEPmFIUJolg2WqBGK0y78cew98muFIkSW/l0o/hgnRCAx
X4JTZzwosho4mCOCAyzfcstkijVYLgUJI1spkx7wcmxYNTCgquc0aRnJDOPx041x9HEvV2giWBnt
rzysMZie9yulJzpG7WUm0xMZJpZWmRL8jkUdizfQKrCFZtpVyr2BQHV3+8Q3Ybusr9FolEXK9+mO
nFb30oi4UlEZVq/kBh1sGt9UMsEuPHvq4iEUVgpIJyXtTkg65xGZPs0rw6kZG++6uSPN8Bia+ypy
oNgSf1UexsQzlqhno46r4EMnRM2FgzGnx0Besd8efUAx2iWJJ1KHij9Vg+ZRB/TTxBShk8ypaf2T
v7OxDSqWyhc9eOzfwECA/ve+p+36irOQaTTXSAhuaiLhX2CebpEQvkg7umVGovS5wgT93uf3+Euu
zMYNOFS+fMYpK5DH1HuDxfro1HodsGp6WqGnpVNAB7u9zfzMDYDedo0oiEOBUYnW+DQPTosEfMiR
gklKU7bTUdGIXeK6HnXkcbC3P9avxYs2RQ7dSMPqr+P4SxKaQsPf/QZLj+3RvZ24ZO5oEf1cNXbb
nUAywNx+mYEBVm2aX4MqM5u+nMWp5H46ROjBUexLA9GiQzVXidtvfxwAiMZ3KmlSdsYEsZ9BrekK
C8pAoIbGteG7QGXoo77u0vrTSU8lOJfbif2HPs6EhwzmAdbo6oGb/F9UHhI/6wKL8MwAv/6GcWoB
h/SY3Cbm/Jy8aGPdayjcs+3MJeZIuijKktPdDZ8rOw3jtuqj0uy86Lwr3/4bC5hBheywUInmYoNl
QfbCdj5KIAVNg86MYlK3dcuai+rl5wmKhuu2ZA1wcGa/tjVNPq8ZnxacUx4kBtobmy/7eXoENav2
Olm6Wd3imuYvdYEKonQYWAr/zn9ndtPGJLT92wyl4V9nut0zUfFAHbAGu0okFxww4F38g7q3/Sj/
l1rF1JH3Y9ktj2fsFt3yCiSgEEFfFbQtDu0Tb+XK2eoUyCWIXs+x4/qgF9O9F+L+rn1phgBcZEVI
9qsDRkzVuo97kuRz/FYh0zM1bba8Sft2Dj6PWpJdEXyE7YNIw9j6/wkzYO2vjp1jP2Pe509COVhb
KBFbqSp5z3boBwUXyS9B1wLMs0pQgcRlSnnc86PtqG1dsC8Q03UKPL9TEmYND8mPu9YHovGn3YVC
v/4aH0pEslhID7gsSvQUGP8NIZSyqN5ijD3u2miNFnYu9hrg5u/h8GAsljBLGBMkc0ZsODjSsTNI
XK7UFxuQQrkbcMlNrGx9SxVY2Of5WAavz9bta7gcbDp21bWIoyoePxhu8mH6JzqAU/RpoYO6PeoA
vWjyk3y10nlqhIHJdOC+yliwk9CTmzSxeGpfICzPXe8RN3vSfydzvf0/VHiy25tmaBdGcnsYc+At
3DcqKc1rMZOLHJJe3k3qo32oMYYmZi1PnWLir8FjnMfsm6jbdCvFWpSqJekqa1DJHOhWVrf2ZB7u
E+YSsrKVLb4uBCBA9/zXK7AindgaXNq6f4odoe/fjnkKl2iYDrtBe5KgzTAWyVORo97ADRZj7c0L
1VjCP3b6NufGwTwt+Or/6I/nQECYCtEE6+wViqiDiFxqsOKdR5adPeqID3GqTBzS0V9kiBHBJGZ7
s7OldnZqSetLEij6P8OMAJlE65HHUKbTb9toD9g4yemYQpzhjzCQqTDEe0hXoOKw5q4yHP9oItZc
H4h2g1c6dU7xA/DgXZgkCQvTVXIRZxWjIOuH8N3HI0c9eT+N70lQNikB8D0CmU4DQM9PlNXyYss7
GD+kUVlkZ2PDM0Z158AREY2HCLXf8e2R/QeOYhbu55yhpl2SnQJBGVI3FTAFNH0hhNk3njrSr9p3
I+9RZPQDK0f/qR0oWPrZKqdF8zL8I0zrkDv+wOriF2FWtAuLcW0ZJvZIopnAmGu3XYYZWPGPm+z7
toL0lvfjagfOCSyELyxGnGh1dhSfPK48zntFl8oqQ6vShwlU5jk9ap2Bl2avVVOfDyZtQy7XH+9a
wxtCCVoBRRNXpwytiCJHtgddCghc7r4dVqKghKYtxbaQ/S9Ait43CfC1v2Gmb9620evA49NqgvkL
LRISXnkihoc9CR19l/5p8hU16YMUyWzwk4E2h2DA2CShzL3h5fCvkurrXQ8pZaWDdonDBJ/jjzdS
xakYYTMPWlk7mKEj5xjmJeaB65IWMjEVd4HYC/ol8cXcspffo8lCkOP2mYoPd33FXMUAijR/6FK/
bbt7ueG+148/mtnvSQD3kZ8eJt7j0q1mYvtigbpDCvSF2Pihzek+LAzBJPMZOnVvjq+s8Qm5kN/I
xDqtR2MSYK2YGrz03K0uIbaO8qgNsTb7/IKGhBXxW0+6z/OvRz7CpIPcVd+9TR5T+WpApr5ObkVZ
6tWz8ITG12qlKmmWslYqXEfyxiTe7ZDRz1IVSQ0dMgfgkHpFODdVk/Gz4qN7w9Pwm17IoTNOT5NB
SWHPz7kJJjHB/lUuLQ4ALFyHdj4Ey5SztjWSGYv9YX4LCsVoW2rjNp8Q5iMXN4uVTbZ0VOnkwQu1
WyHTYB97IpXtdZkNp5TNx0mj6Ixw/VO2ttk8aZiLD/dl6eWvXSg/MT/gIPcE/H1VyfiiMCAuyzME
DQptZS8BK8QTG3pLQPvhkWtBpi710GZNGPjjV+XGYEOu31IhfBEVzDEIAdG88Yx0J0/jl1DFBJD3
BV7sF7wcOZV+4J7KYXpT1M+zIuMwFzeGomRRFhcadkH0TcSC5zWHXlF9WpO3BHRsLI7zF7PDdSgt
e/BLptza7T2Qbnm70OPeF9ZE+vI4B5UxWE5UU3ruAcBWBmTBbLweOqab3soJ0gAwSyl8BdYM3ZEr
mhyK3dppoGpR9jMLHttZH4m370a1dcv4hLtwJADmiCKj1jHlShPARzp73l6LrF50O5FDVue/gd5r
hpSMeGiuZ9oBhxH3I3CW3g2xWVXXdSUlgsJHpXKAiNmuJoWu87h3nwaOE9SHv+VqWFdM2joBR1qN
zHi3uTXuGRAYr1xA3H3Mpv7siHlQh8UZk7t5jC1anxlpIXrw+5jQtDMWRFghcMm95Vw7Ca4MP/yt
gbkxPOSZG92tz+WVl+9i5FuyOFUSht9Ni4YmQbQWBHJnrmwfqXIpYV4sQoWQIjtrKnZY81i715Uq
Emr9ZjQ6RoQ9UNtyxinqdKgCVwzlFNxNCBCdIVw7XHjihX1AEvudL/kTTV7BFWyvqa8uDa+uji7o
gQlJcQE27qGxWha5dDLjTaC3zY2EDU4rEip/nZiYe/6pIfMe/vkbS9eOacGlXb9kR26mUbKbHH5s
ETj0jmv0wrDAtbpRFmCt0NuelXohEeDIabdBaw7Za2RioGUz+PcUxtLuTPRRzUdeDFyeFwmlNIFT
VPDVi214FNoggTuVtzU9ne5w9x+STT21NQhfulbW1dMAOkGDYMY9Gy2dLXQknMtmzqRfOqQlJfm/
VSruNaG1UP0ZFdkqVleo2fHO2tpmUGQoPJzX9bCUvV/hr8bqPTJJhXGPUyqR5Afu917x23c2mRBN
lbB4WZFzUW7G+Rr6F8VvTcLCuF5rEtzlRgEjoNgsIJqaxY2Hj3MkOEOf+joanXFPIFa0yNhBXg80
Q2/mwlaj2WTocV3NYgZ/awndLhiPsXnc2OAFKk/TcSBL/gZx6SfGvBJliVnhfyKCfoR+E54gjBXo
/BN5eX2dtAjjOrsjL8X4yaI+x9lBiSJiSh+c3ZMd/ndwDOoGezJxIjzHTh6rBrskKwp3zxkjL4h2
m9oMHNfdxqYcxRcsDha+q8vVIFI0Ogf+b64p+0er+gNeuPu9aykDJL8Irke7Mr9bbMUWLoHr06iZ
5Q+vOjkFiYila0Tz5COepygBIodFA3FerDInkKnSSWS3C7S6SUx8v1QH9BkvmLfnZzR0fROpB0Ug
ebUQNt3N8lB4jB4qS4F2gHxj4yMzjtIsEVsWcEdLsHZGCiZw1mfL0qkN9+Hen7K1xGPAHrDNUs8j
wYb9we9tBNfqUE2yZg1FZkQeAOnf8oSVOv0kva4+tSw00wi5/fe0h3VgaV9vL73A9aaXgM3BOkJW
mplNVISk/Z6I5/kB9txtVDZ4Iz90F/YlB0LJ8mZ/rZhdqgSJL2qlOrmrtm7Cucn4bBe0JUNtXopH
J4ewk9689AJU2j3mGl64omWgEQXb41YF5S0He+bbxhyzw8U4DLbRIDOH70wPkCuBhifGmIxAqAaC
WdRm3j0bZgu7N+bR/H94XmkeSFEgxcEvIuMzSYDcGby2jbku8sk9Ohck09D/i7OtsdGrXi2iyjV2
tqOMnABmT0uazgbvpBbeGgDoJE/PSGp8CR+Djfn6IF8ncf3J8oNkuZV4yy4wB/9HrspnoCvEdDsZ
alXV/HVYRMcoDswhUK1ok3obGM9uhuyUfKcIyCLv2eB6aIzbLInaEmJoU46qsqIrtO0upFY/CTEP
KtZ/XekJ2exfxAblp00hgh8w4RTWTp6NXfpEMf3X+51cWbR7HEGo4AJNJGKOXJ6uzupt7nkKNFmd
k+Y/xUFO9oeWtuPr1lMxJVAVdGWh5WwQ6eUwJNCu4M7xtmc7JeJ3Evbnmqv9ce/15ZoK1qrs3W0Z
rPKNb12GDccS4pRP/bJmk6lpA1x+DMgzMaI8fhgbjlpKd0nbBJVtBIsBH2Vg9NSk4AEw5jEZNvq0
31MpDtvFBxcIchhdKefTbPSH/5MoMSkZS3iktQwayG/tMos2ROixMaX5kir9sSObzTs2u+/E5Uan
QcuUg+BSPn4BSUzOk8ZnHe0+o4rDQTHtmIGaW9CS10k8Ap8HS2PpGSfdsu7i9KFkcKsQjyEYowym
i9B4Oq5mipx3mr2UyPWkzeH/hhcCdLQQczASdhMJUiahcmOuR8UQ8AqgtprKXHbppcIGR/rIcLDj
cuZ+TFZjLlRd2WaeK0Y/CQNonbXW3ia6xBqZM99opZnx3MPdeRW8hWVT/IKXSnBmt2lLI+iRm+fN
ruLp3IulOD0IsQw4gn1YnJwehYDjwkl9lR+qY6GOjtvpnEOu1VQud8xnKEntqejvTO+hJk56uNDk
4qlqDTvhuOoXVe0KY63USgydKnBKhyLJk/HqXHEJdSvV9KRh+FIyfsGfRvPx0IXjDunD6hz2Cv0D
TxZVTJBH1PUF6m1UlfcQwjlGYsCIBYr7p268kEt/7SgHBY2xeC8m2v3I2n7gbtZaTzM/DJ2kq/vO
B+1sE05S2oFb/iEgdrozPyUtRcNtOTf8m/W+lflVSzfFwtMC3Wwr/QnN7Cd8zkI+2OpwguRvkGy7
bTdMjokY7DkI4Vla1dzpJANKM7ak3G+JP6btp/llhFDX8F+UJeEt2L246UXqPh2YExQD/G/9aIzK
I4t2KLo7eEojpYftBksxkAtNKrvRnee1lPOCslqJUahdBIWH5J+r32Nf7i8vvrbN4QJvt4o60ZP0
7VyD5damLbq1qHTiHR2v4Pm2Ycs40M415L6/OziuRxKxde7fROC1zBYZHNx2MTkwaYv2K+MI94bW
pVb9dGc1RDWRa7IIZg0YZlC+Eu1ftW5D+KoCuT85SzpWlTUIbPtCjaWlEdS/kfY7B5Y7LJ1YH/ah
M7/Iykf8CkDE+EqQ/B5/ylgPph9d20dlzcgd0224ZZ1XjwNJWzTmAUZEC3OctP/u1AjDT4LBOTsh
Me15xfTA6p2Emy2+1B6aAEMJgydMSaslm69uQL4J37gKSioMMGQOAUHW/vpuERF6GXrBkbE0gvM0
ZTXF9ii3IXsehN3mHPgobxQNiYTtvlDHdwv+4TUksD48674tzVML5O3NdiyiAdy5mVRIJvPYdHut
oHt4Thpwj8A71pVna6IXRGccogCVkl0hMYzQh5zsu4B3/iVj6hp79Zbo/MtINRj/0XBgtS4BoEx5
C14+hKdk1a6XItiRq6YBkls8LiMA8oUnNxDziVLvV3sSpdxwaZe2cwSZ2ExzBLM9awSPvG+epm2/
btOGk5fF5S1LF6wNuJ4OgRR0NxYaKneLttNjyoBqjRoZMbf/SUIJTeCjeD3bKUxpMVV5nU2vuVlW
A7fW+TwdfUG7lFwM95aYAJFnkE7pXviX+OQySn/n2WvFnM23fyY2mi89NK4uhgDVHHYz0MLYl3Fn
Y6TKCdHP7+zEDjXBQuqgh3kloXWJCCxRr73RxYjAHidMDVaZnMw88CoRBYxte6WP70+55uimwrRO
tk/ir6ObbA7Jzs0hNx9M6AwY0CZeZLxJgrLy84QtmdvtEKs9zOuCKBxJwraKt97RT6RtX/FksPS4
xzmpcYwm1sCgS70fO6HYdCbjgLxwGUMVMHSrh8eQHGYtdyghrzPNfYV64RbAMpyaSIhKjvDFHggA
kAOxzr/8kAQlGoyxiTukZamuL2GcB1YtUffrelh63k0HjvpkeMKduwCspdqQcTgUpTABVSkZTNYZ
uYAI4yyLsGxS7q3dJAB/t7Oz30IzwpJ52OBPptWUp1JoIiJ1hRYneF2WInUUp6RFA8z8SSHE0btG
4BamH8ux4OY0b7e0WjQHogCZtp5hDSyYCCy0GtpY32Mu7UntWla5Wy9T23h0JLVAk1OSkW02j5So
B+50FcwbRUO4jcwMmYsDyV3maRjl3NxmubgqZKm/qFy0FXqO5eM+F4nz
`pragma protect end_protected

// 
