/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dD6sJjMckNM/hk590wWgo7QyLBP7qvuv1GnV/mfQB0w/i/pvS4BJcnppdBuizaQbHZTE85H6pboO
mTjEC8kS1yUyaRKX4KpOmRsaXVL7/iV6Mc+EyHoad/3cx2lAwTCRu6nptqi96Q/dtiPbQirlE0cr
bj2VslWvQXYp7agPImHpkldpbIx4OKKY49/lmZgzjQmz1uAl0Vpqn03TZsorFhKrWNa1NL2PWEvy
H6r6Q2NnxwJibsxIu7/DaDQZ9tx7P3Ox5rT/+t7OV/sWKJMNsqkendhSkyxMCR6Z1Ip9YxyEItGS
Bld1ucslP9zp60t9CzMGZcj/WZZ+ve1NzjV/uw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="NlHs8opBWv2KH1hFnLsdY2EH/Cy8LVzvJ0P9w8zUaYI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3200)
`pragma protect data_block
jOrE4515xgbASXSOIDgmJvUoma82NC6svbmrewllZ04yfBzxUt1KmsOZ3BD1By57vyN/CbRjrB5D
pG5ehbTjRdtLML5HHtj34GAKA1O0KqcXGXWm64FRNj2ugg/OOlrGdhkSCoacmHSHDWR8ajBWQ6o2
ZxydEO0m9ZPiPzskGFexOuxLCvdozySrIZzONOrGvqgpfDkSGuLCz2aGAH+jwx25enCQ4qKjYPLS
YQ3ci2atWhyDvVzYO382v3ax/P6r9Nf7E2G+3QyVvOsiFTIDSQga9nehcULTN5N78p5kw3DjhWGP
rXr/wCJ3scaQmQ01q+h+UxgOOnNCDIbFuq5hFgNA2SLvi5wuXuv4rvHD5IARMEBdljTZgyrneHw0
PhG3wY5Oi2jiNW1dphI9UIaNZhjddY4MDq2wttLKOKUE/5YTSoc5zdxUg0lAPn5daHvNIsz4seCU
PZq2C/rYb7GVpfuMrj8wBdjvmdbOO62PRbzP+Gb97ohu5MDjVNIn35KsnG7J1kg9Vip6M8DkiZrh
z+rKZVOO13wtDvj9YzaG7lrxxjMKT9j7p9lc+sbGIYN0hOj2KmLUk4wzDPTJiMzmHwOBRAgmT27X
CBMCWtwdjWxkeqZXpk4lmOWWxtos3X08TjRHdphPHsDpEB1bAtHB+b5rCfzH5UjtiLG+lhCNV/nG
WHTwmapu5gZUC0SxChSRuwksUtuSIRUWeN+swWg4tpvau3IjVkzHmmGKoGMhGhFYjI/xVmri9+iZ
8NrfZwgJPFCsCP2R3axFZMCaAkCk51atthEJAoGlfy+qQHf5cOC6m14qTaRDJqsDUYWPMQ2V8487
myztSn+w1k0TmVhDK9xgqH1ITTDEW7wvFoJL6FC99c7ftrMQ4LAzH0A0q2bob4iuC8Zu3rvYPAca
N+/eUOt5Lm+Z0M/HiTSFLHDq9ZZSDMkGrXO4TO7Z7YnT/PtLbFrs6ALyoq7D72myzWKPVuUmt9nL
YkS/8R7ngbBYBTTHfi883cTMiS5cO8SHXr0l4PVZHuANVDXeY8TvxY+Td/LXajDzTnow/QCvswH6
CmH0i96U+TGHozXQ1IQ3Dhfuk/MojzqUSXGVLvZgN3IiAAf3s0uJYkqBVADB0caJmf+pGJNiOYRE
OjLb0QG2ZZe3AxBvugPVytb3DPn7aWeW3cusPUX4GUizHve67z29Si+Sn98AyvmacznWm3S4hvRQ
q/zK0Gq0M3JKah7EnbPuD0doSIHp8kmIcTPlrB4MjqbKmMm3a1ot12yjm6ukQkgUiEu0LybBoIhV
5LcNyaOIxtqqeYrYzr0iP7bTGeCKekJMsxi0lCzCnTX6bQN14khzfHNZCZagcDqJOKOaUPt8fkNy
3GJOIohYqQ/T+I20/WqnJ49rzYcpCvqmxH4dTeAlqStSZ8JXYsGgSE6t8yJ4cnyDzynTQJ7bQ2nP
t7lcfFZtRbt0Qm0J7ANCusNHfHPU71q9wHvUCPGuA3oQg79vGW1D+7kc9vY8ZJxpoZwmeTNa8KEb
zVrBhmxcAUpk6RhiD3Om0uwt4G5LNXO81ULPyoZc2p8n2tezdURtGMjRzWexXHvrfIYqMCFFmBNo
efKifSsPgB0FFH9bCgRPrYsM7ZDm3S14oHidmLr043NuhXm809vELOrA1Jjge9Jvkq+vgus9hTpL
n716WltCLHgWP5HxN1gTuEk6BtVuJ/X3fXhcX2YYI6hm5jZBIgaWJXgVFJaswN6rK+U2FVQrW51i
r4Pcy8H/37EeLZNNrbJWFtvjN1xFzqG8mA5jE2INS5ncJTpbs24cK/ep/9/eVkTgR99o95tezBQq
ooo5N2S2aah56bu0o4cDYHfiWI5eoakBK99pudmcYhtLi0uxngp/YiVfx0fz9hyyJy4hlwHZgFEV
gV3P1wwV2t6/8vXBiWnU+9ukHNtWHycKLV2nHi2M5piYNhYt9NvfGSoSXA7rQSToE9mZCr5teGCR
OLZ1xHCaMM+Kj1ptn64Nepb0pXqNekFhLp49yauPToyDmPa/FaJtdl0+CVgJrOX1O/RLWAcQv6cT
tWWbZSDGVVDQs13GyMccZLs2cLTlGxHEsBVo+GFJUSiyEmaPFdlrj9dlZnZxr9rP0ZOGsC2xTTHm
yJFepYUIwcHb9OaH/9EqTAPaCFMvY6qvfIrUqvwyucrjHq2sTkQyqIY5vBXAOcmqe0OBik/Xuibz
baa6XaRyL+mUhuzCUJK5n9477g16TKensEqXT7xzETd0kS9Ze7Upbn7xpvdIijkzQT2IyQj1GHfX
qUgD0DHfgAa7pUyAgrOc1q9PV3dAfUEe99PN9uw06v6YMpgcfE8mSsZeWW9lgp+gJi8lHUAeUx81
RkWlOf53tfq64lI0sjryYFvAb36qbSe31nWWw2qaIMaYPyzKh47VibLusSPTeVL83kS7iprOAxKk
3NDa4dxnH0QJiXyIGSK5SMqr9JUT8OCb4DwDInakwKqMnB0taGal7oWhiwSs9rGIWi1JFz/W4rZs
CtPXWiIPfNs6qGj67rwktviQQh60cGxDk+RIZD2sOOKxDHBedfr9N30VFS9srlNlggsNN33h2Ad0
IZaPY+bNTEXClE9PN71oR/yAf0LXVO7ofop65EAE2aN9D+5v5bHSRGXLZv4lTtiuTRkZlMjgGz+l
2nSrVJvHh3Yrini4RqvH/4UK69KpzQ2J2bJBBy5y7hNk0YF4V8fYyVZwNh4FeIsk05cPBveXmz5i
Q7iFwHSEt8L2wrist99O1wmSZV3EfWRSKEj9o4INwoGVG60t8CxklYRUcve5Zpus8PkyRCjP8Pmf
zDMI41DPiE1VE9ILaTcyK0/Ld7eNW6o+QwK0fk52oGksHAKnGEnhwTB8kH9x7sA76JPQaYT2J4ej
B7cbG8KY90epoUiv7A8uQ2B4KrqrJTI8qmvp/89NVpVJwG42+ckYvQx9gM5EVPhI+C/K8s6bbw0J
hrziIUTCkN85YlF/sb5zhxwQmwwKCtWh82DL+caQ1frRi4bfSCekSHIqXzpKAft9fQbRs0F+atAL
faCInRRUxzr3XbllbURLSyaGD2O7ELY8rN+0VIUlu87BRyrL+2QrIVQL521yiUVapFTfK+vsrmMo
YeG/YHRTHDxMLQbEiim0b6AOKzdux9G5JxCSpu7v79kVVHZvSR6MSzDCxkz7+eVlkkHUBk5WU7Ly
9tXXEHHbTrxCr9tnE36Kfquu2fQQb5i52pP+y5OrNWZEh/rbDw0xduya2Bt7oH3+uWRHA6jvCT0k
Q5MWkn+fxxN7ybVf5xrqNHAPYfI/fyaiZWxzucsggXeh9gpMumNEjtT/XiD+OHxTSHrsLkxlxlMn
iInDNlENWu3CL1/jntGBe4jgPioUWWdf6zx/5Fh5k0IyZ17ggeYGX3NIk1Bz7Mb5l9SvZ1RJZwa1
0FQEiS7WWIA2WiBM0qfyTXhqOnoUo4kitvPc7ODFDaLXzxlrqPvBdbsDB0Lca5A+HtQUxHZgexou
+cS43wfOc8grFEboTCzRIB5I3nThgnSalxYnZ3Q7jZelNPtHo1LvkGTQWedhY1wDGJ4etpk6cFnf
rmpY07vXxZ80+2xhLXTBvdcQV2/0OKKNMq9eicwbyjDmGIz0z+vBM3qsz5g29OKZLquu02wMnn3U
BR4yseWgaaVOLMCnYLWpgfd+8boVm3/UuDKnNdQOZqpuhvODfzWoeFBBsAW09i/DGc+2ak1bM+mk
sHR2rCr2gtA51C9FcSM4V2fsPxh58+JppTwA2k78t2LqDTm2XcbxzNbyC300C6VwCUyi2kG0E6VZ
JLsvt7eZjhYxDqcbzWJcVSjXg11pFvdaOFSTw6Qii+6SruzubAZKx8C5MVP9oT4LAQxxXidwnBCB
uXonz3ozXjsuM1/6BH+VJJyO0tR14ip5hQVN2U97czbo4lfo8artwtaQJuj3FThXcZdUKwlR+i4T
xiR1+5lRdVxTo+L1/EdpgpkiLiMDhY2xG7DjrVBTq0+XdhV/xmRNA/ny+BNhXiNtXXmmnaTkSyQ9
avN4CIABH76WFOxtt1XrSM+efNIesDW9s9MA7GL9RxgbLEVlzjufSJHSBSVuXZmoTbmPDJq5bwp3
AH12uTmlZK5wm31pMi2TwLplJCPbnqICZyjwQpcGJ+tgyNdvxt5tINLd1Sx6kag+ucqRkFn7YtzH
y668aSAHC+BieatSP/hgU1Qk8c0jnTAH4msh6/zST9+1vagzWI/wHO6pQXL7/o7hMphIDSokVuGJ
TleoCpMOWi8=
`pragma protect end_protected

// 
