/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
bc4WnAkqx6dlMsl5fn3cAprcqqxHUHgVY/ImIQQum+cRAB7ouhGGGf7iFZf77q22uZ5IUqV83Quw
Hyk2hoLyHV1tsHXgJxRTk+FG0z8kNO9UiseME5aOM/+f1fcoxpdwoF5Nb9O6O9ouJZW/9wU+cOBn
deDxs8Fe2cl/gc7w+7aUoFn4WojygKnIaeby9NCvgShnH90A/5GxWomjUdPAdBRy04fmF471qpG3
rcDSX8G6arFIKQEh5UwVCLxQIuBK6e0cztUh2ocE1tgu0ybaWCTYOjp5wNkYHxW0TxCBiXthO/Y0
21pIqRWTmcspQgDYTjUBBMfo4xnplJBqhrkXZQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="ASJKkguRF7cNZtn0GfYOwaRh6RbIlcvsA1oAuucVfb8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1040)
`pragma protect data_block
Xy3DKr6jQ6T4G9Vc1bujRvk/IOEpZZrd1qMcI9hmvvRzDk/psCHTMZY/3+4tr6y0P6GeqO3aZhLn
Czh+nd79YmJNM5VcLh+Q6toWNP4HuJ1oOU3y+0wF4fQGdPmd/kP+jEvtOC3xaU3cRJBScICt9zmx
OYXm2Gj8tCn8hwuYUfxgrZhJiji0UTPu8kKpV0CK3Wr2R1FqGkfIAt0yddTBGZe8AyS6/WUT2Sdb
PratrImyvSTUaSRoMUGUDprWg/8nOMhHG5vNnFxmZ1UTP8/rqlpwgGsnbhbFjlSFPL5osx23TxQY
RhQdI+UxBdQRUs5fpAqULD3+ZgI0vxYVTcBWgjxljONnQW3pJT7xvFzVsuXUEhTBqBUDqWXV0VM+
8DLi/TLeNuRX0RzZynAXxTZaYnRhS8modUwifaUJEdAwv/+5ymodl2pPeaHFVn7J53UwGKsbWsaN
Kp50FEqUSXeusWkkvImHPZ/ZtaOq9ZtTsFjHzIw67qwWelN6b4taC9J4jhvwdKigiBEye5v2oZ/y
OXxvjJEV2N3lDqUK8wZEeVivdPAWb9pTrBcWpVZfj6McTLNuEFKb1bexFvzsw2AfH4Jf2vrqOpxN
KjsOWtDuT3oCpy0xA1dAsKnPCeXEw+aLCSwc7aL7iGhwkj5LGE5Tu88KeZMn28fCzAju2KFgGYU1
jP4zwekVnDjnVv7trow2M3bllgUE7glH9AQOR+jhXLrhpplWaCj4AYSOJmW6Ba729bAd7WQLZuXz
LGkr+OClTAQ5G2l1FVeee3lNhIb/3n1z3/a3H43wDOpmjX9808fhMicvuJv+H1p+h9+L6N6EWFqF
lhLrIPyGqLqxoZw8Gq4qloBDXsNaPCLHxHRaJ1p60+0w6dTnTmZHfxmJFGwFtZQSI1sRldkiCVin
WRqro92Qxtxzzs7Af56mmHBFZLFzSIj+k9gh+lYuPPPSHhIrZEH57GEWkZf/t3kTba2mJ8usYVA8
ju1ORbMMQsx1JeZ1gw60jNv73jEY44VkXTvG1czfzNvz7ofypJyxYUENxG1BYOsX8q9DEC4lAgSU
s2c5kHrzoBKBx4JJT+ztFY4b43aQg9Ib2VwIH7CsFMICBXQHidj77jVejB6yl8b8QmJh9mP1HxKQ
EoiV8d7LEwmQL2Vu4Gs2ZcjwO9ITDh6iGMw0IaUYv206vO9ZhWH6v4vANA6UucIMwJINuUFDxb24
ekdm69wHN7TBZrS7pa1dpyxSpI2HZ6zEy2Liu5EdHnzJ1BbvDFlGSFiuxm50DvG65M0SySdXPkZO
gDxk03YXMhPLzyzDrfjsijyMDKuyvEjkgtgJDwluZOa/oU5+kJumX/IFyMAq2Sijhs0LNcjoCf6f
wZKf8KpoJbNaXtN0LAU=
`pragma protect end_protected

// 
