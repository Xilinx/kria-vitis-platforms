/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
CaihNQWwu+qKJWjcmdIgzgKIXQ8l3vMImmWHnChjYqoa51yMcErBScyiE64YZSDih9WCUqsVfjEZ
HfdPZ9ljuyASaDAJWOBnJBbhrePBDPO5jKkFmPbv80QoBXSWaNMFc5sW0Ulg3lCiE5qq9SVr7IMd
vkFVewJkI9IJKPXIqEiYLMio527A7EkzJrjUXC11BQnTYghbA5n7/6q2WIDOwjQ+BdLZXxGdIUKi
ihIieqBZEgdd6vwETSGv3sSorIwnUPSueC94L800xEEoFQmghwgPGvLA3IEIqt1YNZfrY4rcuvTH
rxE5ve/ar6tMYP0QdSitAf/UOVre3EWtsP+Jcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="IxINXwVvXQ/n7KwTaYrPoEaEACBK27oPy3cRIdl/LOI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57840)
`pragma protect data_block
EiGu1ShDtOnFp1/lwt6VhQRGkioQr4+9yyNmO1imSLcQGxdvupVNu0aFmTXbLJdJnmM27hEBzpod
nXpAoxy/J1hxX0sKJiIsZtN2p2ySstRmqfRRsbfHqln0i/y8hw6IFrUrq8ShlMp6kxmh49aJlJlO
XpnsIWrJz4l+aQ76nTEPTaNW/Pyuf17qkjWAoXvuQSCwsu0Ma4RMD1G5H+UwEQbBQ9XEp0aqimc7
MNQacymOSmcQtft8whs1hmE+YsjNbGKHDtC8cnO3uYtpSoG1HvJfrQDIR3OAP55qHqcfw55ymffF
QbZUkkL6r7HFrLw9vOh+26xzVzx2cCYW8sz93yIYXhUBwxpxCgiaz5xZzOfHK7YahLvgaT82sACB
YbSalrksc86m8e9Rs6rpBSxhJM8IRDwf7dYsKyknnP7b95bcnXZPd8JatMLrHWAsB3i6Ai2BXSWD
ry4DuwXpb8iPBuE/IEruI+/hX5z9u0/xnR4WJcF5FkUwHgKa/Atjffsd9tlok0oF/NRH6QWpf6ay
iDyEG6tp1XSnpFkgdO0LM4m0DzQ6W3B9lxLSiowSxZHkVLpcmDtlwZ/mJERPIYLsLwYhSP1ifzuI
JU7cvtiThedddsGTEzsNfCfyQ0CmQcVzMHsacCeFvI4d12ZP21IzlfQquoyE6s1xg8U8sndmD1ku
J8MzzQ/Y3yQ5POxEX4HriEMc3ufoV385rTKLNc9i7T0MNn0oOWMCCPuHtL8sDrVjV4o4TXT1X1aF
2BQOYfykwBCmeToLN8ITv1iGq+ctSTRWJHynldyWy3qYNmM5/z0fkjRMjhKPXOiSJBekQJ7X6uEN
zd8GSroNZfkHUYkQdXsfDe1uWLlaxAodH6BtlPcuRB2qaa0FesD/RtZ6NU1hSUxDfhVBTYtm6vMH
FQmbDItjy+4HtM8eUJSLb4SAz9hKpaXqkGufBZ+R2YkVOxJ3o5kD5Rqeh1waxvAhCZRloTgWI9Ih
1lQ9n+65+yzoG4DxrupVyv54OzZyWlINsN+qNVT1OrW659OmKzDm74flb+bRWtCkxPnjd1vu5LTQ
As9+aFuG2QnP3mcALR/beFOX9aTVex1O3Qo6DjS0/Ol3YQJSLG+DgGeWkzKjajEEyjlxhq5a3OuJ
DmsHzbXBMo+Uj8zsRRrkeFps8N0oH1floZarvufd83IGXi77so3ySvks2s7zPLlAqcwQ3CjL3PeX
zI0Q1jPHsiwbpOTM5IcK5z6Mr1QJGioG99qpGIvHO/ukjKbSnhheutcYnGOnrLCBqgGbYMkGV1Un
cr5hFQhvkaYRObFd/6EWjCI7dHXwtP55ETii1Syj2jwCwnVspk8urX1Hb+4yNmmJg+ImWDo6i6dB
/EOMiQ11frSPMaW1NhQFcuepYikgVz5ntaE06j9nmA28WDJh8Syz2+uCe1Vt0mD7XektuPPkKQf3
nQaVIrBIQWgm09i/WMr998cxkoJQpyXKpaGdFTgw63FyfFb6nsg9Fekzl3Z4PVJEYMD65fto9geW
RIInyQkVFkNMrCCDPAo7CFDkPGHCzCGSmocEiDAIYBp009AMctBmX/Jjryk2R1Ga1Owpfypshhpq
pH+Haf2Hk6ZC8EXmVfIY9t3aqFfeFHqO4rHz/OzaQqElB3M5/wPNxlMmhxh46tPKqtgLPpp3wBf1
nqsDzOV5ADaVMPh3nM98pamDC4bpYUxYVT/GobWH4m1ZA7Cuej9z78dJ3QiYS5/XOY42QMYk5WQh
57fvgVNkbFmWcbtlIi00li+l0oKjxBQMNeuVpQudpFHYNzzVAhDpgOV/URl+wiCT9oxakKXRtI+n
cKX7Yv8kJOjgRifv7NXSpKowHZLa6/wNwyQrcW9HGEI1q0JK91q06f5eO37Ac/7iOnqXx84xZBW3
TujjGKr+GoTwzBTPjjvB6nDlX3ttBupJH98rnQtyxJXO5yqwyvChnCFfMadXmWsFbhxRdlvv6pKr
H6MWnmFwQ4McC7t2vals3AGGJ+tndvrT9QzZtaxNmRBtrDbTkURtBQtKoGD6eT9FTCpDD2Wr0pPL
GpbL1ly6RSHzEZ0l50MCgcv5y8tf6J+6gjr0T7IBEx3uifonzv2sJagteYrpxytUAxe/ujfKiDDh
5rsHnHvKbhkVDRCb4SbsR/xFA9FM7cSmcWPqxxnHKS9zR/5ZnN7FTH/amwbaNIw51Kwydk3RdNyN
nFreteSNiy2aQHgVmz3/oK9asuSm7UgAKN9uPN1Jf9HGdeBnt8ncjlnIDOb8VvqpI9ckw//zJ62w
7I82t9RiGxaEotUOVZ0Jjx6y7Jidz+2T5uUg+CnLGYi4tJvAjND5gFHoNZeHX+E16lUIqmiwPZVq
4+7OXalezPMI6adoErFFC7h68GkOEPitZtaUxsEEqygwVqNcyBGHhKBLQT03Ip03pU0knxWZaHJ4
lZEbmRzUNmsHj3YOaQLKYCjOeKbpUQknLKvRmH2AA8BnTZ9LDFabBcsD+nQia9mvaEy9zG0ajIjM
GYP0k7EkZEjcIxCL3pctXqEYvbzV6WqW2zzKf79t8mocFSx1E709jYsi5kwZAuDkCDFDV/H8VwbX
NRLE3Y+UMo1yf4iifFwMELxNRbdR+kUsHaRCfeksIvc6VE9xO21iOyVPgP5xvnW61KuL25yv6pik
1YX4F/TLzKn/G7EBHpwEeML8rlc7i1zBW0811Vu1NXYqtMZf/U2uUEJqvu/VHBvkO+JZUYyAiowm
xjiwto4Jnohk6eDQse3ee6rX/3E3DzLRVlzUO20EWjQtAIfkEVA7mYrsquPwUFyDE4OHc4iunTDV
U5G89tw0YJKOqWrZtshwdT7KMskGZGMn1ke9mcnHZVjsqZd+EzSyfdBPCowFLPLTqb7gPBZKj+RS
+ecRMmnNfhkrTmXbDqMWCb8nTjalUL0koosUOhC2xL1l0MVR9ASPKQCGjjagL8XGgs2PXy7Om8sK
87Q5Rijz20oT03f5yweWixxE28EZuqR8150/JOoByhtYa09gSWHiVMJ5RQjQgUkW5rbYL03yGNp3
txBoZEC0S4F15ctgym1pxZV4OnL0E5gQLiHeoDU/WGQxC0nKOsztcFjHHx6P6YAg7S5MH4cKuSTp
AGr8K0w/uRqUUy9aafH/zSVz2L2AjuDOsoNQcUb13a8seJbLcX17Zc0AHFOFrZLRvON9KO64Vjbl
33/j18GXYzAaiw0/Q5BorM/iEIau5S6bLJIkVn7Exc2qCrQwzWYWZiLEZNNa43FYSXBqrBOn1YUs
wDoQfHFAmxgGGargUEb4MFNsM2CxQh54N7yu0KrFN8gwfmbo+TjpUYvS8GzeIS6+slB62zuoMY4J
934Py282jxG+FTnyH4Uo0EggSRgmAxmjCeUS49YiDq0EVKaXoPyInr8z3FVwBBFJR0bsO+kBP/fz
QVr6baqEVKPZmSZRUcvLQ58Vyd9qeLE2qY1yJ5wk0L4AoYfbLYn0vFwswL3epinyzQinOsxYzGRs
qoc7N9b7UxAFSTBN8MTj/IWq60aXfTQGMpDKLCZGtBif2/YfCiHMRpAK2ug3r+0aC3juSKUal4YL
/lASCW3Zasf5jDuCd5hr8mV70KXTuAOlRRMFKBSzDnUOrwxJbu7EjK+Fm8FP1CjYHwZTvoDxE7iY
xBRM8zl/arc3BzY6WG3k6F/R36eaIu9UqtfpicKxqv54wjuYERCIF96/dDp9SZl4wR3uufDwk86L
j56n4pMlrw30G0FCNLollG8IOFEMB5cJgjiZnsJKzKS8eEbmwpBSzG7Cup6SAenvgHkL+f6oPiwK
cmhCmWyhhqeXATvV5vqkOgtsL7kahr9wwL+J69irkskbk+ZZpqJPTkL1zKBUoxkHWFoMXsgEGV6U
RwBBFOkQ2z4Nk7cLSaqrVTNpEkOxgWDcfn4plinTjc5Soy4Y/aIPTUb0ojPlrxYLMAg7QxAUk3lc
QGDgPF/Rsm8vqKzrqeDVSguRN3fasM4T3NNC/YDsqzfpuDAiO6HHiqEYDzucsPUyC88+cSD1la02
1rvtKKsspT2LqRjMTBwuncSRxwozwpLH+QZdv/OlHlyfKvZQyoFQ+k420eZ+tba6oUYF8rz1KSfj
ycBkrttgPee6d0XS2dFRscfj56R+BEjX7lAZ7f9DSSa+0Ppse4H5FmuUiQfya53EhEpSCqW7y2fy
cq4I4WoRpgMrvDzLWYbdsxEfHQONbTmvPaDoWH5bK4ZGor0a1RfCTPbD8+DUv9oqgXHNU6rrhi68
Vqfuqhl5ciNgBmloLb7FPCcwQJHSJKSOWzq5YYRG/0B8dnTQTmhSBa0/NEVxVs5a6TL/sm3JOKcA
gkrpoyo2Srn4Wfc72VyEh5mhZM0+0Qrli1QgRARrhgZmvAvW33qxv2vGr8XexSvTaxbSyUYXXQP8
koG+ookg04yzv74AFE3RmtdFhiQM50Ek8Z3uYIOj8hREHY/G2AqHIpsnqjs3tPtxI8lEScJHlek6
lkdDpeb0uvfzNbUsU5+PrDyjIEZcsVq1MQcf9jYwGzUqXLaG788Q0i7i0tnX7EF/TvJB3OqWqPsK
NHmE+J9ojmdbGGtuzdnBx/sGeXsdOWnybmiSB0Nn5j8p+KjJjw3Ym07eU+zSKzxRwB2L69ksiAMn
Y9BxaxVWC7DUe0/3xCdkU0LMpdk96eus17EKPov9vqAIm6c7TD2chMVF1KhnxBDu9t0sIRQ0Wg0S
4i7HgTHV7wcNu6oF6r+tiVpqZz06S74Q/ftRxS6Ph32C0Lug7A/pUB6KnaMK5UNMWAzSLP97Kejy
Rd9ngyNSD/eUYL1aUstLMiP8JR72/DgZz/YBuYW1lCve8f3lO0PxJsEYL580O0fLdk6cgMwi/2gs
ByTbAyEKwTtuJO3fAXDtI17fg8+vvcTmTZVD9Qg4x6bmZH5XL2SLwSH0Dw1i5WZ8pUYJLh0KDFXK
tBuiDFQVrElZuxLUB+Ey4o10g/xtczgwZO44Yb5RLIOEyE/Rry1V3UDPAJ8YehbmSRM1/bTByfxI
aAVwQWdIOE9Fuj4mAdZ4QLD2jd62PmLzi4nA/Rx4OvWyMHZWMq9aWamgSNOS11yXvvi4l82Hu4l0
uToH5oZmCVm7ZrWHE0QKrexaGY3+aJUONPxenn6WU3iJ32wgzm/Bs4LTrHk69Cyiz8UkZO8I9jXf
j9APmcSh/tth7adMoXONOBp02kwdKzmS7P1QXvE2+7B1XqmvJbnmATiOTsIkYIP6fkC/PX0Yu2qc
SZ+dLfUZfAiPsDtsJPbqlBzeI+pM1w6n2GFrk0YVcG2zccFyyS8Hsi+hOtJBk1F5jxtATRB1jrez
/iTE58mcn6NfjKadTu4DuXUUziZ5EPk55BdyR1Uqcoa9wpAACS9TmjBMbpn0jR5bhn0S6FodM8Ly
/73KCSja8OazKEt+ux4mLwjr5Uyz1lkq9p0E2G1j4VY3qTD5TDy/FLk6jfJE3mPiuj3vT3SIQmW6
WqD+sj+Kmy6NUB0xwyld6chv0lXM71CU22SNDnEKw0bUWcXY7wr+b/r0Zz7RsqlhvUYHwTss6vss
3rY6N605jdS+cr32fHzStuIz2uLXRyF0cZ7aMs1qephFgrCerVu31rZ9Pul6hC3NsBQvexYqNofo
wIM9OOzgavuhfh00tlHQhyVuZrJcU3cMS9Q5yZFzNeeRxJGsucFW7vNaO13qb90tS2JVqd8yVanl
KXR+lLEXUU2ubaAAdGwDcoljHG0ZW6AQVhpDUkOxX0hCpLI3qzZ3W5Fjo7i8HDe4QXiPfej20ArI
GVGG6yF7Vx2+lfEyuy9nyp27p1BC9eabF9WOkTFHg1jRM2KbcZweWjGAUZ41G+5lmJBljgFa5lsr
eB7CPICHkj/RDm2D2xsBNpcOXRW9IeRv9SWqibwZrwW2+R96UCBznrHjaf4Zws3QBm3hyGrZulVQ
sNjRfPbmMKl7MtvMhisF7Bfg66zaNSOUWEoeR4fKJdRju1wxJTo1Uq7TZBWyIMdfeB480DakAyVl
QiinZcKhFaNzQC+2z02trqM9unxUZDDayaExzxh2HGS3IGf+umNCd+o2zhVKx0VDdMGsm1Dii+wA
WcLuDsL7n7t4DZ1JoTrrBN0VBQs1SuwXV0bcnyOyvIqaSdR2jsRHu8pI6Hq//34VjUXuD3YgN3o5
pQwTE4NQmp41m/8G9durxqseQIBdiVrUDeLvdWGZiJMGRLEFO5CFNiooPmshk9awgvFxudmH2Aab
CN5LllvCfDz+dit+r8PawODN/gkYpApjoWVM7hJ88joYwlvgOK2jRjyQdXZG16jmEeanntt0Q1fb
QqDyyoowNrSBMvqPkHDtQiG9yqFs/1IP/dRNYj5UnPV4AAPJ/VwqtwSNxEThIZlRznStFaoi/HT6
GDZhkPeg3YFBMgQr/8aGO/4M10hPUpace0+5AY84SBPZovWaVFnJ3OA+hcwBT9LOdx0VzkJyYCUD
AbBnVJMZNog9dhHpQkAnOUvHUjbS46yvOm23S+z70tCMCcDwwLTNFXUHKQG0v5HH17m2Smg/y6jI
m+a+3UEs0vt+DPpbj6aokF9aYLTrdtTg+f9tRLFYEoxhK8u+C9ZOPBItS+a+Zg2z6QYcHZs7trnT
45wHUBzuBYVqw6e5LYqfPoHr/MYY4fFB2qiy/o6PTRBHcHfB4cmiU5wIXOmo5Bk3oi+PiLjcA/sS
xSxpvceprrxU+V0l282bKiOEIExDqEYWrwJmcmFizMno8fyG//hjnE+pBzPBzPyuBF69uwFSQm2c
jl6ntCgHyR2EwC0Vzsg6Jl7sIacpMZxIBZf4+bxQngtRvcl8nBibVv2ZOuMTf5iA6YRpP3WO63XD
gnnMSQVyZGL5MrnpYHsbEmaLavOIbqkTtm0e10j9kS3cL96+AwJ7H7UsTVGvbz/rx2rg4R4UDR8d
J4861Wy2DYs5fjVec93eyWZ8Lia9StknGVligSWrQ/+5KElGMcL0/PxdDRXZskSD08V7MG5ZhYKy
Xe7IaxaVbDvVKswQB+2QC69ijiNOXjeoUWdU6SUlbMaE3K5jYKD6DhSoLU8aeXtkVym/ADW2nwt9
jeUYYCjoAer43oJYAFNJgBE4kip7SLCvp1J0qUgIXu0vgNqEmT+aMcnedwp3pH/a2SGlgCmumIGG
jOuZVd21aOcewDUIdT+0qP01viZB0h1rIxXwpwup4uvQhuk07wGi+7eCL1UNbd9NjbQNWvuL6QQZ
E2FSzXgAU7sZoTz8wYW/FqymSOVaZHsITAmTGchOeYKBw8FR+ttdU8Yw12z38MbkGU7XNTBjzMzu
cQS1M3Yo/EjpmenQ6k2xirL3HMV0urDoeUiNAFBykE3pFEvWXkdLPggcmT18RuYvDab32p4MP1N+
MtA8B3V3KjuzE2nJs+9IwtuzEcQGeeJj5d1D2t4FSohuWc/uBTLSVYxb6wJ4quIBhW+24dcozhiF
3OQuZXCyjN+AeLsnPTZn5XBh6wKSIJz+5mzq9qnY3tsmmmyefHYB8FPu6wdAwx0gdjvlHq8SrPJJ
LOkkPo6VjT0sJFhWTawQZVI0Fjv0bN1mVvPNV5ytWpBWlSlwMMLsabMUftMKn873Ug/UjmvlIAhb
zJGFTVwwx2A9vlMZIVIwC8FumavNrH1Na0atsD1kDylyzNL+jTnXe/uJSzID5C8ZvvPYaT9a2BQA
Y1SoaClze6SqxDcwr56kq7HmgBCxMDBN0NOXISeTqw+V3UOIGZ+k/FvRAeJ4RCGplKW5/nxiTtif
vMkv82XvA40CUtByHJNCkBN3c5LWk3ObytgcjSaKg7GVVX1wMXTp63CzvShcrF3VutFncnRyXCRo
rQfyNMD61SK2HjaZX94XWU0/NLyuvP9jGqndo6VcR0LAnoxTphn82rF6MjLp6fyLrAYCODKIYDno
SMWBAGeRcEY7oX5bGpqV7/ivBfQMEeupc+cblaDuRmTWcIbXdE8tdwUj7NDtqrPt9FAU01yVoktH
zLUZA/6riJCGmxVPhBWFSeIT6ibUcz8D6PtDBq/3KSYAbWZXLGH55QEeQd2aVIW42d8KrsLM/Q2g
R5bLdh8mmQNv15a0/C/cmAP7xsNlaM6h6Wc8L7MHMXpTsknbUEhC7fowd4DZvW8iHJNJMIMxbFJF
BhdRBimT4lFzx/JKNqNw2xgmzi3C16Gp5qkueqNgG2iR3Y8SAWlDpVwL6qZPCbG6IcSk94RrYrUV
u6fBPM6K7mO0exCseLDQUiyFwtRvlMhZs1L3dFvqEu1Hibs5ncfmIWk67ks0HTcCz8kdDjePqi7A
FKymTTQMJEU1uO+67waxw9iQ0mD7TXjOgG1+hkVavnS53k15bh1FciDvklfBG4i8q48fkOpolMNb
edEaFYors7EQSRbzLZIrOJnINDPd2OmLZ5kY/8Hd90gCz8wlQwc+pfE9ShQ68IuSil+hqQCgpq8s
RRCmv8vVuXR8mALFjxpH9j4PfRQxIqtrwnklI+STkBcAwa4cOT2L432fjvE9wES2eOJ3b6acde4i
9w08DJD9XAprnPPZWQaXy2RvvA390f/rpnh1MycziRcW3aZi3z8iwuRqBs+8X5jGZ5WM3Y9aPuq9
WNW8vCcthoq/q7oDiExLxkPVsLJe2YQ8l/amqjRdysH19e312mYb2vMyn8nHLAywVmjWq2USAcQ5
9dQSXm5PEJsPo4Ee2DjBjiSM9M1XvXcG5X1YWqjxcHM5XuGI5B9C//zxpXk6e1ldVzacKF7mckaZ
rl4FTIO6k5LFk4uKLPjbwXV0OPrE5GTnk78hP9VMmGmSFxX249cGaKc4bi2PWgMkqOmAyvOtBRUc
izyyh20yKgDWlBce1ebqxc+bTA5gXdbW0KcTwOg953nPwNvByvrMyGwF3qy25fUVLC/P1pSzOUDt
JWdpi4q0BcpjcruWsCYoSr0RnXT0hybr8oSzrtGXTQvR7qVizogbuJHPOBRvDve8EvTMTdbLpVSm
MXz3mYV83LM8iWPhxFl8mXwR4YVsPlEFQjA4XrjAPE0Jm+LzcZyrdIQWICjXkGuV31TvXC/MJRNy
PJXFqPoMohrkjvvHcrtQ4JwRm3WVOFUVbs5DJOfbifUcWj/Nlwv4bkCKtWVOTQ7wnFNpByxQ08IS
ryVI//0IdYahFk9KZoVeGooVxguypLelaFUUGyhf27+hyHwFwiAViNcp/LID1Z6mWSciS7iUsCSv
QthrYSRR+O2TUH1e3ATo4ztwAsDE1QYOQuxJMZf0AW69JrQ6pjT6xf16yKeswyOAcRytyTMBnvHm
2AbBm1pGLwAijfrZi+kKEWP4mKiQ8j6xbRvhAYVAoMHZqSyD0PTrTd84LJzBfa3Ih+AyBduZ3zym
56eF/uDRMoUyGGRlpqrxlsD9KZOwnj6Yxp0xa00N/3KdFPn3tZRai1KQKHOVPyEaXuEfzmFsOnVb
peBA6IDjvA4po6JEpUlAUyc++sVd6A9TIyEc2RN9vvpLL0RadfX9YIQI81kXx5xrHHIrHUXppEMh
uUHizDdDR5IhTJ5fujdggAiJucgAJkCN+E5dfyJXkCoOTUghzg3lt5QWjZj10RxzY7YQfhtzF+bu
3+6+0eZ4aexh8KL6+Uy2eAvcE/ZqYxG8chsSDqAEGfDVzhxCEScNm0piw+7hRplrtNP6H26RFWtJ
ikXyyKmMo4WHNW91Jcydu9+EonevjYGg9i8EkfanLA26bzy4Do9I9RhQniO8qYm2fmn2uSK3dLaN
8+vpp8YfKgz132j08pQYdapZrvAmnSArzXMOqdT9Cig+4HENAMmlqo48yTGlH9J0uzJDOTD38erc
Jw19rAEjk43A6/cLk9cBX2GCoE+bwLCyXaT6cnRypBFuLVOq6jQQrbtP99HxtwyITb3oePxVy5tx
2/k+RHqHegJuEa4rMLheAHZWTi1Z7zYrGFCTcEoCjhyoTj7/Ua5ZSJu8/TFcjkz04M4EoNNCmu6H
YBUTECrQP/TPfOyBt+4uWk4hrLvNxUragFkEU3DoDbHm0qBDKc2DkH40fIl+d8FbKLuN2Ghh1KN2
dYP0RJTGyCOCowbTbrGiVlnGgzRSGxfpZtfnyR8MwPb4VaIjBa/1VBxPHhHJe57ZTMYiUwL/NI0A
rGk/d6OdFF2IYaZhNSBwEYR9dkR48eWiqRYOtTmW8ISRle+FqUwH7Yu90spHFe8m83zWH9HVFyvH
F0vjWfqMTFp6ZA1/BVpGsE2zAT0e0kVbJwvvbO1SZ4p4uGtq6S2RJOEtqdTXQmW2QLyCWcjrowmv
JoRHOzzRnJupQIIo7BbXelTbm23xXptRxwti/SE3oJf26p4r+H3cicwKkt/GIPN3n8ItFxEC5VqY
jezCIKdLoHKxOq9lucQfKc3aNbn+Sx6t6meZT7CNjtCcMjdjIVUHHiQsEpbdLGMDj6AzaEGZftm1
ISRlkSl6f+Db+UzctqPgj0rbsk7PiRZjQSL8rT3xKjnKMPPPfLUwhjHj82c3uIZr0WbFLuddE/al
0GM2sFOpFG3IDVeZUsYujD0HgN7J8ybpisKy4aYRhFxsTRmRwJetED2W81pKAP69ss/XGbu2kK/U
pmhukE0VDi94gpCp4cdtkD3DKquhZpaRZQC44r/Vwu/Kyt3Nq6FS/y+oKOwwwSXnT/85Kl7MR/9A
Y/WSOS1zKiRQHmEXkss/p5zg4SDHANo1WV2TifRnFYGtDs+DeLcBVKxsc0SDY743Zh6rc93mvFwc
FeGtzUZvlcCjT4BRVlxYQAPkM9JVlfoCOE230QvPSP8uygPrOrGPbBCY0q25AIyTlIZvvEm1fqY9
WPjnnPyJWKnkjJ+GtVZOpby9zz3jpy+7HLtT0XOIaBxiPxKOYTzvCKRfUr7A10u+Z/3xUcIrzMnH
us9QjqJeyGkhDd69awpzdAtATk29lK8aZ8YH0S1VflGnzresLgSl9/0ZxX8Nifjmo8nwcGYmu9Sk
3CPBq3RGAgU6KMQofOKNuJW9HcPP9ICXKh4i/DP6GZz9iroAGI+CiVXZtGJq4s2ktAjuvK1K4/5I
2Ur87ywlZL9VD4yKU/BN9wBoLUVAC1DSqnI/rjTOFhwQ/UCtzhtUG0BKKOZhsQ/kIfmbi6zdgmfX
xKtY+9SpdtLwPP98i3U1SKVFoX0ekKT/iMpaOJARflkWmDHP8S7k5DLV5PAOzeasqgdk5pFJr2yz
6YS9hFxK6cT7eXDTJ+nNi4jcj27g7Hg+vxWBiPg8oXb6SH9DxCZCLS+42VKy5Hn/4+VwTWOrBZZb
wbnj3Mmx72kwRSsDB+kdKvqkvclIH1RxLKJMQJbWfq3zEa2++dFh6k7WdycOjEAsMjyLEBeRYu3S
JD0P9Njt/7WYlLIJqFCfxti/ULahcxa7ywq5yA5tpM9YZ5WvrBEYy5+7gNNy5XNVOyfLO3E4Ilo0
0vML7LGBmIg3ubwQ+fxgH+4Djy46NVarDvyftDsRPP4bWX5z8hG0fw8aBcgjGaw7snmgwcmFMmCf
KbDPneGP6Ux0WohyeFZR7+LpTpU0hFzlyFHaUXziYH1CYjvHuCaIuCnlrBSgxUkcoD05ghNQgWUm
6enEvw7l9ONqWbDpS+o5t1lWrKl4f+Huj6fKeBT9xc92wMGzItGFFZggjwRFYvVANz+/xVcxkvdc
lGV5X6wq1sQkYIVwJG+h8sdwJBm7QUkRqg2V4fgoO+atRO1p96UKkcB2MalRyqCkprT96q8Ra561
r//y8dQ8CrI06AfBDzl5bvAX1rgrmJuge9N7KSZag50v+Pr0KKBionJdQVagc/O+itYsENsSOS/6
FaZywZC05OqdD1JmA3hHlozJQ5zJ39pIq6H74x+M2zcFXdTTfDbmBK03AVNmCGDKapQ7/nP5a2At
2Bi++oqap5qUiWUYzZmwH0lTtlLsEeWY8qSceMWTVU0pJhKSKyJv6gOi/aLY7UpWABnr7ubVz6xP
+6TG86KUdwVYaZF7k1PMJrQ53m1dQ+Jlv9CrzLp2ci1JYNf5k8oRUZFar0NHxKfn4JVfVkJnnBa+
oqgRnTw+NlngHhfcbCPc/mwr9izUVKMzvT35N+lo/OJpNvA7C8w2o7/I90i26FUmlp74MD9Bq52I
+Vvuf5VKvxAe0mYBaxmpY/FndZ4v4ADAqH20Exo9WqkdObo+MFbCbdiJ0YLc+Au3QKVqB1sE161M
/g9kIMe72Xz3qKDRxoym5Jjh/Fq9prTztdP3VgcnPwyleyRF3f6wIXApJhs2FUzRWtt8XoyZ195w
lh/gOZ50cIuhKCHQ2EqsFCoQJcitetnL54OLJUW+l/zX4xkv3Nu5VfECzehD6up6bTcdWLq/oxZl
XiTdtxmycZtFnHhq8JnmXGH1xIIxMMAaF1rMTZYc3NW3+PKhub9DFle+RBeEAgfXniVEtYFoeGQ+
QC7LDfRGNVV/Ft6ieSIFHBuGRQwm4d6Vp9AfQEGQVfhoIN82nvYdP3zuj3dGcVOpR2GYXN90jOzo
eGfKoEFWL7vFy+DJSg5uFftviwRVwjH8suCFLR/l9f94+QLjo9ubc4cjWQi86PMxeSLTL8Rs2coF
LWg5YbKltHdFyNShZVXLFGD4TCovlzSA3HeFipSHvDXjcU0BkzYmVX/BWsH2fbjQQd4G1YHjyJz7
XotuEH+aatLmpvBN4aqVUtR1b3f8/14lsnOxl/9gyhtUk7gy2P44Uu3w/mM+15LLlnMqCnn6HVJR
Xd6QPwi2aLL+X0TMYBijI2MCVNnYXzfQAXGDHsLg3CRVovHaGoYkrKOul20f9wt8OeH3FSOis2MI
0zuxip7MiDJrKgkaZSfXOdYdGhs/qLo/c0S8VJApyQbx7HlL/sHfo0/GKfFjG99Nti2iarEZ7par
2qChg5DSxsW2JhjjEW27KdtxzvvPTS9LudRHm5bycijiW2CDIEfKyJCkLgExExH1HLhoUcPZJPhS
EfVy09jtcjtILCQXQ1k91JfWvZ8umS/wJq2BkcOY6F4VKql0GCtg8TMcP5Wu26goqORHTvz2RcbS
kRQsG9vipVrPy66qoIeOpHJPgH7ZyuYo+54cM2sfKVvKq0K8C3qg4l/ew9TA12hRqgpGNgd2xbAL
YPH3igK/EA4tGe7K+4ZvOUpkl5Eh/VEZQu/U7myBKvXZst3dcBHEKfcza+2AACNaaCrqO+xoR2NJ
+ATvPJJnzsAVO0sUQKeydJlwXgBIsofK6+vj2UvxSlM0JiX45DoDGtNFiSxn0we6KqUg9sjXClYD
xePBORkh1hl/Eg/n6BY81KdbcRKZLx60IHQNlRx51DvpLCuF4ibe2orfuAo3y/dZUkZuGqTLhae+
OvLbAwk59bvClhrorQ2x81Oh9y7TNMob5/0qSjuTp9NjTTC0rIeShp+nzatiH5z8xe+RkFtLmYaG
u2jzpp0QVoZF5F5LqR/EW9uBHAxI2JraXLnLHAtUqqRxrnuHznp6xL9OTFau9Tm+SKQFqrTJJgmo
bT3VToFdQSO3vLvUWPRE3F31GWBT+CebfScgjCaU9XpWojodOYJ1Ln2BgDhQgWJiKAk6yjAQ3Zaa
TeczVGhEmUrl5GGShLi6s74vRotr+phyF45R7SzOt5udAOGAewK7lmun/CGqW/ADQiHTGwV+ncg/
WP1ACBKiWBQSq+2FJ5mT0QYUotX2glNgtmPkjfmEoBhkeMDaNeCKtV/wZKdNlFbBu2HT2PwAkZU7
6h1PUiL2p8MRjlI9zBbdA4KRk7wrJXM16MC9DH9FYtN42q+GmBVKn+YyeSRR9Uvt9027QIb8SkWG
4FcYoxCHRa+xXCMbwe1qPnAyibqKuDfhE+6WcyTrqXLTq1M9FeV414lujSOcagx3pnnLjxmkFAHz
bOU+kh+lS1KNp0pfEMz5uB0HbzUALo4Ci2gLc8e8Zp9DCr0NwcmuKPHvp++aFDNO5hNT/RaM9EgE
KSbN5qcSHwPYilDN4WrUBoVDPwOM2ZY2Jsz5x6PaXc7ypaxtdbt6zHO5O5axQTM+TOmJ1KXCGWlH
+t5XAxLmjPd9FhfcjDngecMcDJSxnV3sTNJmADPBaxqWCFdWt25f/oQbQneyZw2mc8xWQYYOykZK
Py9L8QR0UTtLt/MmUOEjqFNR188m9y7PDR6P6K/IyDZotBVSnoxJEkL/Ncuh5dRpw7tvwUPJTfq7
tecsRf/T5omxmdFMQUEqeP+Z5TdD+nLFFK90OEp4UfWAup7cZkgTdqXZMrGEguqtcUnnrMjvom6F
yvzqoHVXxaSQWTWuumQ4NVsrq+/vtBaz2Zw+eT10xOmc4e/2viZuGaKBBs1ntY+2TnXfPzFWR8hW
a4wSOWk3mKte8ZTyiZl6glQ3xrwTaYUzt56+kDJ/FXmfbEgnVmXY0faVTcHi3zCJyfKum2Xg2fH9
8Vc6fQXkRWsGNkQ7fHN7Z8FBf1uv57+fKCJaYJ698ZADQl2tJZmqDtKL+2U+IPJ53lD8IoSJBcSM
63iLhts51lbbDcg6hEHaFRQA4qGEOkXeNOyD9WBplbpH/15mff2m7342Reg0P4bnGl5f/oI6qfAQ
mOI9veYXn9z9/xzAxRc40sNpwySdqCuWBfr0LJhimAjspL6nH3ed2wVKRjdpEluRCX9BorwjHfBL
4fcArympkHgwWFATvn8xsC+rnBKbtLwkyEccveJd+bkfNIh8W0yYEjpudJAuzBv5aT/M37+y6p5I
DKWfGmPG/930Y0n+1KA0BcQtdFERXv5kk6jv74T5dkFw+vPGgl7I/R6GN0RJZFWGTLnkM7X+d3X4
eOP/b3J6NTjQKNW5davYP4GhIQexxEDcDB1zmtyYbwzR7wqa3ffHl45LiA6ez3U1hICDE7/U/yYi
xih1j5eX3LwloNDYWFotw+D8yD/5wpIwn8gynUN/ilVf0xtC/p0d0Ti47KL7i2u8LwsAwYRp88QX
MHo2OjE7FvJ8LxB3VdMYqOBaktHYp8Ox0EiFbzSC5TahD42/d/uRLmFa3JOEldPtkBOAgztUpglM
ooM5RZR8Xg/UpmuR58h+Gmi8DpSeLKK5WLq8GQ77k4wat1IO9RtBz39a1XRsxb4Ia9lu7gmBQNyI
QA2Ed3mxwfDfOI8NblyHfIZqyS7YA8WQHUoRUagOIxALaxRAbvtYzs4tkQcBv0pi8K3XmR3VqM6E
QUhIv3VrHsNMhpyqIfnVjX8XJhzLned3TcdnAgbxq/nz+NCm2ppUptWIgr99cJ/xQ7fbY2DTUKFP
ZWWAr5VPrRtIALGO2s1MiKbnSxa+48LKLJmljj4X8n0kOcYjmVu3vVKrH8ViXd8z7yqJu0E1nz4w
on16maGfJA2XQi1AjEWdyaSmqGmCfDS2cOk3LTgBC0yfz8VfqJl+EMOS0++EYQu5+JPxBl662zKp
WoReoh+E79BcsmVGd58HWbv4vLiaZUZcwcKlxy54kgSEqdDcpgDd130STyKA5rPKqbPK6PET729t
zWjtXNpcRtXtjIUvjH1gZ8NSDstI+CRom0S1QFsIft1D0JIqZ3nthWcFGc5zFSa8tgUz4AxlQFP6
ybW3DXB4RLLzv1tEVbd68IUrIw9pyUWZSKAld48C4w35hghU39c6j3psOwo1d/CYrlbdAYrZFr28
OwatAY7m+E205fDxQ5pD6YjXWmQGznY3CGkkDPWxvuhgVFeICNM6jh9CbKbuVUdVx3M27vT25pDV
okPlj+4NcC5yNnRnKv0dkTAdman062+Jm/FPkr81XxP67rsShDeigFQEG0grPEk7M7EvumjiotRu
qCksuNT1bq46xoN+okwKq9UhzmuolR5xxVkIVUGYiorfMhf0iLMuJ6n5NPO4UZtYVF2mdLn9llPa
GGFwsSCkz8/KQgCCYGm8Vx/NlXDQ0/ZUQlDM8bEHoXuTHd8nMfpAU2H27XgaFlpKlMPoUE1NH1bn
Aw/SKRakfTfjE2dyfLlUifup5Xnngf6wbNOgao9g+ApsgPXeUUd0Mg9CTGvG29EJNPMIpdsKocVW
w6y72Wm2MBfF+//O1RYy5S4nu1QNkanWouw4wupoy2wF0v2cBoQuIfHqQKo4dcCyGnNRFrPzg8O9
bSfPt5jI2+eLOihIVKLD0oP16N0BLSkbsU4m8R710WNfEgMV/OdkCA2wu9+oufnhMFiwstyC316r
vRjBN9eCIiaA/oqt7yh1GDspy2uULFp6vZTGdN/q3surh8FqxNOAy79sKMAd0uT06vw1dJy9dGAt
RCoGabWsEU7+psrst+w4cAuWXlBWISccO0yF1bW+uVRZ6gDTaBBJXqfCfHzG4G6rHSqFHPXJpNW5
JKejHMeyyK8FFIMBaZ7vtHUd9gSStDZHdnQcalz8ypmJ5YvOco3qx4ix3BawLCe/yQMLYVKl+aP1
r29OYL6RsMHnZKOyb5T5U4GqRE3p/Ou4Ug5Zx70KoX/QDj5mnSvvim0Kt6fsf9qVO1VEhGtxlKaj
4QT2z2UC6uLxkts3sQZOo5SMDIc1xAAY3Ku8OspYUVVsTj79IZscwagIU0i3Z0KU+OGtJMWq4R/W
XoxS84cpj8bh5RYgAwKVhH3iqe184DFip/MhfwKwgYBmD6i7Hp5AhjcSc2fdRGUXf4Hpi/zVMGzK
bpUAh4F8aLRm/L5TRpMbEMefNFF9xEmW4JdWxwqXRlrsGe7CVlTwNhYQClNcEelzicJrQADgnamR
ZkPJRPqhVkQbUVgve9WfaNRpc7AVVLROyc039WzbPQA3gOKMFpQAxhfP1MirqqqDahjsZM5feQUH
H1yRIrTUKW1ruYppMDxUGntJOL/0y2ZKMRnSBMdQGhDJI0SDUk/jpfKIC9a4TxWznAXPDfIm3lDN
Tn9ZjhUPdj2YUaTbR+TQmXNXrhWQjR5lnswoAkPSU94QvZj3vnW0Vb87qPfSCK2PyHrhu0Qe8LcU
ebpTff3tlA/9uISsKfJZ5tJ8sEsLFMA2OF9M57eXwSzz/+Q9FwgKYGES3OoIiwNi4a8jAsvP/8kQ
mEF0InisrvLw/cuzcnZTe0zS5dZ9BfTBnMHMJSz+F4mEWcX6Bb/IB3Y13DERw8P+7Nveqw2jHm1b
g+rbof6QG/AOuwAEPF3MEglCD8JA+EG2YhxLhG1V0ee37TFqJUn6sS6OgT83YPkLFtSpV9uOYd+i
AkP+pcqt3G7F6oW6GnsUfxQB+Uy+L5aQlUiyLrvOwy5vHYE+hGhwk5RAqmh2yzV+YbImSUNUa8Of
w9WO3JNnLs5cgIDDXRvlfNkKOuHynNtFC5FUopud5ksnA6imARzPCVeDZcl3/9+vIgx0pj2rQhQD
ERYduhoztr75u+HI6IFvNvPf5O4SpsfYrzV9Yagdg72caB0aa9a9opda3v/U6uvl8Xyq0ttY68oM
GtVv7kbYRv94BTZrRpOvaMCs9H4F4kQ9kdRMzQS3/U6LheiVTAnH8iO59xVOsDMxzyxdc0W5dkma
MyLG7TbTIv7U2VxwOl+Bd5gEJfYtV+QOpshKG3+c3GLVYUrk7jZ0Co9RCau6NFwZW3tYk4fwqz/Y
QrJevh0ng4rZ9q1p++UwuM+lFSU0lcX3WETUdLe7dQd+P79WHkvvT+zPqDtuz61PKd53nI1igGDe
f0YHKLswY3jbiaFQXBBl78Jn3+rHGDU3TlxpT6Wd420cc42CVhMkNOe0mfPZthxFi4omv/bjSfw5
1IiXmPVHdpevRH18gWb70LXFQX2pvBEyjjHbQIRTSfx1UBPRQB2SbgEyzF0Fn162q3OaG6Jw0Afx
Wd5X7y3DeLWBsac3PnlaDNwL6WE7VIqCPTae+cEMUwbLn0GvY5l4wfGdHpLvJ0A0l8VHs8ui0BMO
NauwiiRUVfznnqVf2PtG/uXPsjun6bzD+VOuztrqFQ/UhUZsUKo/T/1IdwEsUlYZ0RtJvX03UNCn
YQT+Y3Fdg1bml1UMCd2+Qx0ZrgowRU1qaw2DqcolSURiM+ueJGcMmW5l2kRa3oOODsrd9nvqHrX1
RbxLdt7xVjdyOoNa+OOnsn7J5TLJBTwoqD/24lBpcomnPbRmhU591rjZhi/qum6gJdnh5szswqLX
MgF98lcRQkRIrpykM2TGETz91DY7KLDEnzOSnnjxfGzaEunyCA9nH/zVGg2qeLSI1DqtJw+6Ur4w
ktPCq731PyVpQi5xZLipotx2koH/hbUsBGxqha7BS32S28jvEQ/XiyLRozZwtmfi0RREwQ/1iWhQ
X9LzQs9dLHxCnDjFTDprSDXmVgAJ2/TJreOkTAeFUO2MXcD4KX2eAP9bHib4XLMLP9CfzXedQgHI
u5b1TFf3IfmHUuh4ABq33E+NSgh0menPjKtHK1/Y7SJgXz9YpR5cdzHF8zpqVKaiqxGMIWURO2uU
ekFbCJsVqYdZWw3B+8a05bcKwXMxdCWbUnxWM0wxANyDKquVKRqyXNB2UbU/eYOGMmWia+7qW8CG
ghdJ4LoSslIzewU5b6NhOd3118lvWk8HC7FLNLD1QQvCDR9rfb0TeI2FwtzOMFLrWqd6KkuLdXZX
9OKWLPAp+5Bt1LmDMMvI3rLtKJEv34wSnNSe6flrmdBB3l3KY7XddsBHXRkRwBryi4a05CtwCue+
Rd//3D2GQ45XvNfK4ULdjcj8bQSNSTf1zn0n28Zny/Nk3EtkosNLSlNLhqB0Vdi3wGzAE0UrgDdp
zzGN60qGvJSerm4JrCwHeGDvQQUv6x+ZVVj3oh/gMdttp3C7KUD96pU5LcvP7jLi0CHroou6ZwuK
9oCPIKEN9irW0qf8bnZttcoZ67pwt4WQkM1hWqBi6/n30Gx4pbaPZXYoE1pKsQMf5cWNkH2ZPkbg
C0hNhG5ytX+Uihl9HP+UO7Tjcnw6CR6RFPmhzOofv1WbP9W+7CHgOn+KFd3vgVjlpMs2GNN74y8M
pIl6kedeOarcm+YjjBl2yax8F1dHLA4DGO4qkAPTxu3GUxtVXSU5vnMG0+9585KYQhIc8MceclzU
avGEikDIsE/o+W7qILU2wnhM3Uw7JIVdqzSFFh/zrr9MmRLB7aq/7TaSoNbfekhM/fTCQVaFegRH
obLd5pcgng7/Lbt6foHs7SPmstCjHUocAQyQtNpAUUo3e4Tqc6FYdE2D3qUCy8+D0yw0KvsfIsLS
WqLDxf/c9UFUpGrHfvv3b3iqvLT9EdEP2PKsK1hHecwapRi+fi2QIt0Hn+W/ZrEMbrSpI1a83iUL
GYoNX8iOS7eSmrwNv/Zj+/Rs4v8SRFT9GkqUALWHK8+4w4Atr4gPYcBfZyQEl/Kd0ZJ1IyX3QSVq
jlmuwqdFbfpPgVwYfioYRPBKAzbTizgQ/GevRHhssUU1veNnHm0GH4rAhSZSMEMPUjQmwQyBbSYy
gqjeZQDPtYXds+o6QO/EMLDB1EEnIvs5afiPTFS3Y1c7XcCqysLrMdX5gMXpThdPgleAz6CVA5Na
wowTsDwrWuf8wVkXLRK1U5HvA6CjXTCHVtZQq3kh4lQw1U5TgTxp+dj2ODEzPh0BvLw1iitLaUyG
w8RcPSRX9+Vp+e4LO9jiAUatrd29dBXwKdzcAEF+TaJ8wc1dMx7RcwNI4HsRPnqqKrc002OcxpCs
gl1eBN/osO3/lUOtjgesPIZen0l7zae4LQcg2jSQo6yCnPP5PPtfn0YuCtD/6u4Mrxsl5N1EN0ce
Fz7lJ5x12mLc+Gxv9ACJwNCsuM78rXVCC9W3+XGN1lyiudDzFARigRVDZk8GO09pmBv/F2jXadGZ
fkS9NV/lJeO3ZCnJh9/I4JPMcgohO8Si1tU0LtvR1A5VOhhK4tuFBqEOwDdVC36ZRwqZCGOud3V8
EBo89FO3DQuga4MHHOQKe58waJFYyjALNpEie+WE2RE80jS5IaVFHE4ZW6159NMMmBS2nLi0a2Yk
xON0lHPwTDMiKg6az9BI6CDyFJ2AcEM4cGoAkrbsJ6BbYIZEmy31SR2hSZ6SA6SblpcOfVxiBzxU
5R6DzC0H3LtLcqm03kjI/x7uy3S2eiLky9rNta9gz4hQigEP/Ymusa5T6SxJQAJ+wzqmzCRGpQ0Y
3aEcF63FkklHz8iKMM310JWpdlA3KuMaDXt9/m/9KnQAdqD780Jge1O5atXepnDdP2cpZYiX4aS1
3gd9MzoR1VKLH4bK8CWz9d7FH5/KEUkNreI8hRqyOyeb98wM4M4ai1h7XQZUK86gusH2mKT5aIiQ
+Ifyae2CxKJQQcZ6dETA5jM6rL8+VGAshrGHhNCViA+2Wmi97f1maDZyiFgCCnWQMzjaaEuvo0j9
B9eKSeDn7AgP3BTgvAs/Zu1VOE0wF1txed4JSoDGden4mmwiQGixh9oFJPIkKZw8wwXkOdjl16pi
JYcN5syJ+CFKzoIQO67O3Jlmy0C2Fwuqoei6MQz9YDUWYzrDTi/DWpipT3mW7XEEk5Yur4jUE2Hi
4uwmKbEGFtDJIOnRlQSK2Xv79GOJphyNFGQuAa316L7YrS8zwm9MOjPwGoEGc6plzcm12Mt1drYw
eSoxi470j9TLYiEBj0+8C7nqfmnillBIK9r/Ii8BTiTw1tLHQ9ghC0x1KQCDtz9184LYszsqd7fw
gQfDEb7ejDfMdqbp8V8IVcVvunypmvK47WPaE+PEJGwoevXzXR0sGT7D5q0QesHi7dFC/i8LKkrp
+iHRq00PUkz4VZVA3M2UTAyer+MgKJSiZbQxD5I5kRj8CMwQnoEMB9w+13YoAR+jghHDj6D3XVeY
WxE7KvSYljgrpkH4gZoYbSZgSyE1PNxHCLBLHzvIywoTA8v0yb5xdARDwY4FG4uKgMOuF+lQv1vT
j1By2pugD4lzZnptKM9hcaFncg71JE7boVLjrnlJr3oEkbLTrz40tzlu914VQakK2KrbyYz38hPe
5Fg+OnWxjJ1tQEW90E9QdHXV4W8fwzBl4n13P/9xoEcx4bwBrTXB/9nu/W5jivv9DjTBq5VVkLHz
ENUuPNOtTatOF202B9xCAo/uoweefEkZFhi0StvrMR75du/nCSiAEwrA0hbME2GGhQXAFeLNKJsi
2bhIO6Bm+D6JQHi/92n+o/HSJftB5RO/9ArwxO62yiJGpGxZ2d3pRBatz2MISOlspXMrOsTECGgE
ZIUVTf6q1Ed2Vl/8pDATPPR1d6yfYzuGAm/Qr92RT6f7W38OhT2Hy+Aa/q6IaDoKDwGPsEuyP5VZ
KLi57SYrTAaYwISJR3n7MvD+hKaJzSm1dToHhBY/AT7mimNWuZX/Oy+2MAlZMKMPLDEbb8zjySsV
E4+UqoKFS4QJSXsHe+Ir/wHJlBanVIv1hazEPNHwM1uGwOCHOUvnDJ5vYSsdq7TVScE381UTxms3
XFt/A0Wc3yhTWREQHB11OVVED9pdI45ZVhGB6ohgxh6g6DIymBFNSxLdBr2N5xWnfaeyQ7q+uoUb
6fi6v25EZEbXViCHvb8pU4i+xkL/xQPng46XOgXRl27vbHiampD8KuGQ68f/AYwime3yFM9PiCXy
wSGuaf0NHrllpn5TdKXDbr3+Q+VjE8c6sMGlfibiXPKniPCOqhzjJIkfidGADvDcJ4uwTyB8A7nK
yMyb/ifRMAmQXbcbZRYOHedl1tAaZLWyxjGnfizFr5zChTw0iwQeURBzBePo1A1ITrc3IQnr0Kd5
cTa6vQH2DDsP1oVgz8wUXnaa+CysymFUR+vGI+wAxFR6ALo8fzzekLvLLW8+9RnrrdnKRWSvo7qP
bSmBNYTedImNVTEmI3XiJT5ua5mJGVE7tqS21QMTsomFiyRvmlB7dlEd1GN9omb4ov2/wWH97xQK
hUydrUAXXkYsCtx7WR713k6qeq7QatDX2DagAsMhLvFjaEqroP9/iiNOSjXC7By2ZgxwPBp4VS37
en2ZDP9UUilkLTtAK7fEt88Wad2EL0QOXedJRUbifGtgDSOspG5idrdQYHlwJJkc6YdpcOfK+0wK
bJ6D6iu2WDoxzzTgMjui5tREVgf1eI4/pv7zv5CRXcszUTcXcEQsu7JttfJSllSbVkHK/SJkvcTs
6Ur2avnltyB+1XZ+SUSXjAd8b7wHzdU1mWjzA7AVgvfmP3TBm3hK9xXXjFzEhn6mBeH1V5gG953f
XX8pGVoxlV0c4MW4qb2t/WymN18T4WVSZJ0Om/f0TpNOWIAqTMLzNYnYcF5bwJOsprtq3QbubGwN
ZTQqYpw3yE0u8DUGjAnaMKUbPuoBq2rWOIEA5uozun4IAqOlIOrz1h9vfEVvfvBwSdqbFnLHmpjR
M94A5oTuxYnRpIX2mjwJ3H9gRSyswj68lJsAnpz2tHB1Yp9lbixHW2rWc8d6qccDfyvZduA3YXli
B5S0f2FXHu8sb3xcUkO7qrBYxpIwXqLQs5363k4uO3uTD5KwIowyxLPobDRVIGV/t8REKdqr3kl+
dyRmGCxVJbP4nHLEJOsCdqfoLHxSpBjEiimNQAlRje3ZBtDg0S5XW4FftlDiHd/obeBK7q7fGBUZ
twbAVPtcPuuyJMcxP/A1BhG3LtkSIHqD4axp0sTyZXiMhZ93SBTxbexuDa7w6G9HnAW2bA/qsfHu
gkItnmkVt9XEz1pGsCJ5QNV/hLx1tZmmTeJ8YABkGK+wN8U1bB5TQPDA/rmunmZuO2VePqMKYvTJ
oMicgmCxT9u6/pxE1kXlBLjAfncLrhJ8Io2q5EV0VtHQi77EqYexrUoEtVEp4c8io+cKlLNW0Rsf
D0YbyVuCNDzyuMmdrD5D0Zhj5DqWG0/SynASIW0r7lr9IEmFxx3h0XNPZIyi1ypDP7Q3wTMgxBDB
0hvQuAbZfT7RpCsJFMwcWw1zQPWOU4ZNuVwr7mbS39f3IDfXtv0Dpa2M3Pf436uY4AvcuLjGTb2/
D/WDfJkJKEmBnZzkdov4HB3pRHxTNLMr/ohlip5KI6gQESTq55KTLalLXyYe/esd+7Xx4S6sahrg
YahPr2blZZJbjvTpjXTfopV+O8PJtTx3Ekq3EKWm5RP3P5LgRueu9h61JoGYJAF7d4/dFy88B9ul
Isg/40tzXFGWDvK7Ky1CAUXoljyHASnHB/saXumLnZdMCNTgugEwGQ5eD0tYUzUqDfaFmv5f4lQ/
Js4J4fLtFgjj7coru0v/2avsfeYoKVjrJllQEuOEMjJjGBGdZDu24tHEmZ1UeF1qdbrWV1fRgCGa
L/dks9QaQNfdbELw2KcxhQwmjAz4YAKyDUsCWT4xX8qVa4c+8QOV68bvgJZooEIUir90ATV1KHck
4DWH6+JhjQjKMzB1AB/6sVLAlcLOJ79uLhvyPuZAYT/yrso96P0zUT+zelBEqDTMoQX21nhnCSsh
mdTlxkISNcKCVgUVdP/RsLymgNI+ukrlY6CCtjN1Mh6hfh8iI42pUKN9jBR2SznZkCJs7LJ5ZUk8
PYz7hWza2cIKRrozSCyfaq430eHF9OzHYhCdovQegczoMkWTgx8nyvuP9EbhR+4E+xqmm/OKAGPM
OE2GKVmNA4NNESKOEWboaBJDsNaPg+7rckdYwe+tGincEKpiLPRWYtpfjqbinC/kcbgwsrmdGhPY
IOqYl28gfo6e0Uq2VuSwjIUjqm+SITRlfSik0f3MzeqAhvX8ADywt5f9HZySEuplOMArq+nZNiod
rlMY7QbC84fy4j4ev2ybmKKS5kTJ5aUGMWIHRFRXJlf0YyX65NTtdsXKX/b0EX6MP7kaBssJx8H3
VT8lG6XFPB9eRIqGYiqIIhpbEuVik10K+bnX6TdgfzTVT9sJz9eZ2MuID2fji6I+M8r5QoTGRGzo
53Z5eBQg5u1zUzDef+3TexFYHT8xo1LON+JDfG0hBIPUtSmPDNCqM8qL2BhqvMzDam1EYJIuZRlT
hm7ojEPi80XCRCFstyRZVNbFmY2hH6F6COti8MqjHHuynb0CdYexaM0YWrMAtQ+xj2yN3Z4tS8Na
a2IjbLZIssFkLDuIj+BWxsQgfKVDMV90/w/JWIC32xSynoagtqO4TGWYcuzC6BQiyyMB/yq/aq7s
Ph9kW7wuf7JutAEBCcBpL9MkQwfBDKmjpxhF4i1wve94cdswJISu5hR6hVRvtAkf0Fdal+54oIpt
dGwaV/4XMnN02Ly6TYFbyDtsCE669glGCvn6QumdjFwAe6qiA/9dOIifj+AzFB6VsxgLnXiub6AD
VpVh0WnyS3Uoc01/fBwN2g0/nostOYOLjoLIXs3/b7sJXGHhxlBrIOyTjPV9+HzWmRQZzhIRDca0
1dhstr8rCwIqA+EJGaai3o+aSUXzE1Jq4JGgseWUTg8Gk6sLFfTt/oh3HLO/qL7ULM99Sz16GGIz
cPZ6tT5k4aPQ+EtRlvZCrE/IaxgMyImv29WPJLpLfZDyVwJxaRSXCWdm7fHnfvv7K6F9qpWqqPKi
cLz8yRjPhNbY5nYZb0Y0p7DgscIGcdy43U9rAKEyPqVPhvjxHb1fWdctIk2/LCQtVgGieVE1BpAi
UZmjOW7eTGos2wJV/9AqZIA8ML2nQMBzpw0fGlQz3Nu8oJxexfDw4kInl1mcqcon4/5G35szsOZm
pzG/o2UXR6zKz1C8DztWEVawZ7Gd2Dp+Kso8wSnJK8qhAPKudW4RA2k+ApRkMLmahmI/0yWhQboS
b47Fko6elXY5rcjkLKb3lHwMAxyHv65hPp17/JhC1rqrXpal9Qp5C+8fLZXAINQhhb+DYVjxs0++
Q7Sgnt8hFWgTfIofYaBIKRb0AelQp5IFpHexCvgnqki1m8C/XiJ8PaUwT9pK8tK+ONy9yFVJKcDg
XzCZ5rwzINX4Rd79D1Xc0eRt1qTMtbOmEFMSfLtEgcKVLViVMq19s5LWYUhWSbJWWOA86BgbzXrw
mYPTuNydXdwjEYkfj7kvhbEmpQ5nW0SZiidlUGBLLOfjsVv8UmShxySwhS6vH6gpjA3LCmkOugTO
LqTUgJJOv+Ofim1EFXLQPdw23wUZU5CllJ+vhKlRCNFpYMsG5MkzHfTK8Vh5ykkdwy0w/Z+dQJpS
2FEqfhnKlsPF4PU2bGTsX+LOCKQcpZkrCpavWlnIqKplcXwFsxan9xpHbvkkbOXtSgJFStasjESn
Bk9yItZI9lFwTvhJ0C27d8Wzk/S1n3bEhVZAyMld0qjPx8Ttv2xyXC4ewQRja51VCAAMa5uNUU/n
cBPYqPKWWpU180y8redKkJm9JuvJhmeZjhmUhP2+H5BJiFwWHpwQM92o/MFxR8B0eiPrOR3SDTqE
7rnTCfQQjMcINzI05pxQx0b4JFEZTBmlh1CvszJsfCfbUOZlro60BT4hpYXY3h/cL5cG+ohw04/8
N1dmpCUOHWZRYDMMsn9pHpVHLxldoPluRLT4Jqlwbq/XiuZMAxcy59QQTn+8rHGQMI3ijtRH6vDE
3X02YQPUxCd31/AB7v1Eb8uV8X4EyOURL9Bq62He0gKC/U8HmAS6o3d15RsXpmxexN6OBoggP6IE
Yw0bZbuFAtdMuc5Fs1pMe6ZzcTaihGdrFY4/X6q7oRrBy8xSElPMmlligHLbsrq147A819TDFljT
2qyjgJhkcq3LzIj8zgjvAVtyAQtOpdJf4vtzW43qu/vgN1kRc2hKUIvX0lWetJ8LKRgKRjWAZGln
pXJrM53CA/XfSfdYs8FBQIj/c/mqoIXJZfAP/tnVkQWuEZz7Lh4KlrYx76aq2pBYto1eRccHgVYS
dIReauvofnKAHMpV+lzlbpZ4QrdWCxxlBiSZ68nl2Cp0Hf0UDhgC3RFwDFHPXDjoFxE8tXs5GFBV
u+0bhPXeaerYGK8hTkZIKnhTL9UODEUFCGTwmy4rOJOQB/1iwsc7hqKJWG8f0WO07f4Sm8xEUP5U
ciCWaONaMXzk5Z5vsryyFlHq0hi/+CEKnJHaEvXD1SXd/wvps7BfaCWxpiqr99wZ81HZ34CKuKYr
wh5sk3KhIjGoZkU5j1b0X6WE71PAFtejx7FI6FsVF5io8C/qZpQBARb6LnO5xNfYMmvd+o6AE+ph
WK2fv/gjghnIUsQRXyw+jihhOSTrZbZg25V08e8UmOXwpdZ7QEXwA3NyAS6dnQ8pJeDHUUxGDp3u
z4X4U/JKP5GOhU1pkCeQWQufByDM123nWQLf+WoSh7lQegyCpfPGsZU8cKEhuwCLAt2r6Ma8rlUK
Pf0B4saIvO8v7SUcKak7oFeQz4XGe2Mkd5hNlFb42NAQ/xjlML7VdZb9ZKIL5fim4U+J+vmai+/V
PxegTpE0F0UoiZRKNERXHoXg3bh0LiCuPiu8wf/g2nYHzVNty9zqnaMZcDo/hKDydTiL7Kb3/tXb
bd5TD/jqivaiFg0GR/VSR8yZ1R5gjqaxQ1b291UHBe8y4aubhWWPmxAiv3bpvHKXvALbnM45CVvz
fNZ8xrRcajROkpQ7fm4hYQCPMghipgYYL3P6DDKkBTAJQbO2OaBdv4wQ+iQuEQihrHaATyVr8Dk0
RvgV3qE+SFBawrMv3dBE4sRi7RN9Ffbw4THJjRSVQ2gAIVQHg3bRTwPQ6UdD9WjVxT3QjUFQot6i
rkQ6WCx3SiVcTjJliWraWhaw6E9QhO+WYLAvoqMwZl+isE9WuqS19InLYcJp1IAK/lzw9/6LWA+S
GFfpMifUsRU0HhZZR9rw5XA8paixvXj+Wy1iiPgNDSdJOJeCAALC2vH+tWZNFy5X8dmea7K5ldyh
McWM+7AYYl9gZmxX6gU6/DRqcn9yq3rwDgP+wEEs/jrFd3LDzAlJwMp3/58hsxaSerD551wR4FVn
aPtnYC95uzv0Xjr4DXCqsHuf+LRYNnQNb+olk3iCriRM6yKfHKkTj/FBH71UEbIPnJe348Wqja/e
nM5GWqaF5GgH8qQ5jB/JsyJyILxmch8W954bwijmWaetuENkN5gjtv4lEtSddWxnCZ7/PqpY6uB3
p+kaw4SfkZXIYK5YBhNCVQSzCw6Vv1HyXklwlABWMXVch9zbctKmuu7XyNjgt+pxpk5nUR7GSEZ1
DJxo1SZSGMT1B7kdR918qNoSBsyeAl9aOnavHGpun4eIvGt63uZNZR6ttDzUTYvbwmSfwbxkgzrr
RTg4iix/l8dq8DVY2ffwk3SSO8urg5wE7yRftMLjGJdZA9a/NB4SMciBgBzadGp85IHUDeYnBcTq
CNEDqtTpFSlnBxTqDUnnif89zvAWKAbD2DIL2BP4+/HwUIEpagCjM+LTr/PEY41aGbND4k16M9Ib
odBZRQ4gmxOiXv7+QXHVwExj6xOM5GEjvSGLkCIwYgEWR/5+aGJwfjI33UQnJbYfaWEsr8F4bV3t
Y+EK8nyFlSHz5ckw/+b9iLcdrcCJu9rRlCY0+3pEVkjN9Ga2sjvPvwgq/lkwlsUk9gfa1z9Rr9fH
0M+W4RF4XbV0xa/+0UqzZ7sUqn7uOU/nSYafmb4lOW1j9vryXawrLFGWkOoO9l8NffZAZmY7hQyk
GNUMdhdp0jNIcPGMYCy8AP97bNzrwpi3TPSTJ/q6j1DUgQ8L1OBzZCpICXJXvruRmbeFNrxUqrMh
6gjfuX7ZYGI/a/x4lFxrQ1lRa+0ixGz2xzdwcsh9I/fxqNOuoJ4g4H9uMWlR2Zqs2K8PI7thZbtY
sBy3O93d6he1CUZEjLAgjayvZ81ANmIIGjxAihDIlymQiPjZ3f+hAsjHpaf8rOvqqq3NFjc1EWVq
cJ5Wq3m5pBRrVbb23SmogRK5bnFQdjlc73aToSbi5KoMBP5BtNHDxtSbgqsXOpODod0vEKHzE3uq
TnKkjuJ2Ibi9hwXf/5mraBEfYSD2lfoD62MXJ0TE06pTgy2qcy34iclXRofUI/58BXT2NAzegcLI
J0EVNgIc5E+cflbh1oBXwRHpL/3aEKaVph1FCgl0y4yfJRWVTL2eKwUI7VmZWE4sArCOJk50llhl
kmMbNzmX/QvjZmQxziw8MremFnmes+nxuWc7y4oK/o+K3A6xpuRZFH9aPH6JUWJpKDvfr7/SNPM2
ymVA5kZiTQa0s235cDbcW7IzmHWh3KdqlotGG2mUQ5eLAMNmKr/mujGZcjkr26YnZahVnKsROx/h
c77IV+0bIV3D7c3Mo41GSxVLCt45Z+TdMobwZjlDrIpcV6ibgCpjfEvUnsQUzNpoQZO3KuAkdM0m
XF4asYt07nzjsZsbOv5Wjtk5PN+DFjwJqmxuFlWw9pGzpAao1A7vYN7HHduAsfb3xdLckWZ+m32p
SwErtaDaSp70kNkSo/kMA+ZsF5KG0+sMdMsbb4B5vIF8I/mY8bCSq+yahuVGXcQFIEsVwvYTJJRS
ucTeJKoDx+NrhpHH8QiENYTUGcJOLERLmr7HbjxhXcQTV9SzUATbVwOFBvuwVY3osmBTx1EDbCh9
q4Y8UhTOSeQ6SqLpxFZ6LD/T3Z6a+IN+eUjYCkthfa2kQ82y67V2Ih98OlhBL3IQsqBL2BidGyj3
dmbp2aPLqbj7ccUhix3Q+j1v1hbvV7gSjMO+57YCuKjpARa7iQ3zgEyYFSwU82S+Cb+jdxickqSC
Nbw1me/5hVKnTNMCecLjbkkDnJKgaYxlszIy/tyL3UEzDurv7AVs1REK0406XNIKBdYIrcRpeP9E
Be7fY1ut6jsPXtESwLPxAKZk8PCsOFOA7U9+kG4a/8S4Vn86bk5lPUs+ydT9zQ7kkaAYB2dz5fCT
p5vQGhwRoa+DW6BtiRbiu4XP2CAR/UXO8dCjrl9WjHaO5RE9ud0/Ns8W8sJlpkvei6xaA0HMvtzS
+Re/PnqnPL93xdvd1m5IWh91IUm/humVxgJbJCZkD59aIAA75wwFR9yCbHtXUBJGbXbdTDXDnCPR
AEcVyZ3vYmcs5+Zlk9OnteytK11YTYPwBXA3ocbP25DdD9TevB70RK2TDP7QYoFM5vac7QysJKp/
6wvKvqho8P9vxW2SuC4Xp6OiMbEn/MvKYoxOFayCEDaWOMVPpHihbBAKfAV6WVswuqEeOZ0hoK5V
GvUqp+syhzqY6iK8uFLosN6sj7hWtCZRxYP+tWgh/IaS2Wljg3+ARqMsVKcqknAcCGkCaBN8CzUt
y4we5xm0IicLTUD7UlmTtwGaPXXHj9b2SHk8lHJqWusIDq3AJrAaVkyQ+K3Dm7/a7/1+nTuWcwwT
6UUine9TPfs+92BfqO+2ty8jHxLqo876Go/hMyix7zMTrlXnbsDb5MeEKPAGssiXDzlFYZ1nTI4t
mXow7M4Xe6XQY9w+cyuPq44KyR7/Se6ZNMYjGhkbI1fDyCYd4Df7q1TpBLh1GuL49w/H8uo+6YoC
GbtO8wwQPqWagl4JbZmuaFlDLZQtRjz4SDNwsjLLp776C63+v5pwQrNC/AQ+jj5wrarbqR0Pbe1e
drhLCk/H5fzp8XbnvbfZ5p9Lk0u7gFWhnM4sVaQxOtAAwNl2lPCUgB2Xkj9ICr5g3JdKEpl6HE+/
oTojAAkxx40FIQKt7BePNa8eU0gQ0fLOROyuFiW/ScwbgoL+9jndgRwSdpBQVOnonIl6IuhraQQK
gF6KSq2RGZo7d0owYJcODGHeU7WfISO7yANQb1230Wa7zt6DXvDNeKWuKeU4GRfInYfGv+M1ve24
OoMlt1e0JfOLTYMIqcS7pa96ONuj8Cx2o9xUykESZ/loh8r+TBpoaoQ323B3GQQyyOMa1zU2BNHF
aCpdLVX4v7NjOtP/pv4rai3XFcCTtXLP195XrCjsYbSwpdpTHShD1WXglR8iXcrXScOCxLqaFwMf
Fm43CIcad3lRpCg2Xb7nFcNsyIDVtJik82mbLaCroXqmYL/p3PEatoYdgotmwBw95YTj8ZQfbkoA
me5J6M12vuNeUD2MNSu2uDDIXrWbqenKoVYMx9buH2zhxE0gliOtTGSfj3C98vmhN3iwqaG0B00m
V+fyjxpjhMwQW1gz457uUqG8ks7hHA/xgvkyq/73sVMqFsPE4AAL/tAy5pbbvqsGc2Prdmnj92Cu
gnAkUebXih2W6zo6mwvYMobVDRG56BFFPYCfnl9peuDTTRTOKYhFpSG/A40kijTUFuGovPxIpU+i
O605h1ZXcc1p05WkORkKWEjDLoIEOvQLbdcILvTb3oTlFnQC0/8pqTm7dJiBbcLjldU24Pe4CW1g
XzF0NqIsJHEjIwLjB7M6qPj+BUxxxclJbVJqmO/H8vC5hxJwT86c3JAxl5sjvTNgZvKp4Li6SqwC
RBehmOKJdHsR7CA3HHXc2g6xbbeTDmMRgKzydRHM6D5SvkoAUX3q4nkCYX1Gm9Q1qMz9iN/cx6dx
TYzr6D88rRZU4P4SirrgvFvOvPC20o6yzw5sXBkwxRNhxuMFmnKcE55ZKGQVNMUBOSMoaA8AnEiC
YkrFoWyu+iXX90WuSPsugUFV54GKmsH1TbAP6QJWN4gudYw+zQhmOMZdxerLYLb4s98dbOaSK0w0
zDQK7UIiSZjzJyCwNWsfFmtI/V/dCLiZmHqqvmG5ViOrSdBISbrqtTDgKZf9tK04pFLmU0KHZ3Gu
PE0t1loMvnpEKmSi+5n7wPXjYpxJPnNJwDeOmMlwKvkpmUbt9qNHaWHa3O4ofaz6+2cNFuhCpOOU
1iTC4SIfy1M8A/I0TiIbS8OFtjsgM1Jd/kk8os6CYCRMUF50ADLdn+bF/JUFlsYqCF0WaKk32flu
O/g3Y8aE713hRFlX2dvZC0xYyp20C+938O2MkExnNjXX8R/h4qZtE7xfmAN/bGJUfBNsSY1KR5mg
q9Uskoz3VkA+1kNQm7inIE1x3bM6U5vnz1gMfvJ7pB02YaJLkl/F/WVkjezAryEKWrsJmPVNY+5B
Cot2X0yOGZtjiqMkaY1iNhlqeOAVCMhO1fpqyDTqQDh8u+iFT7tPhsCUmqO/+UfWboqfS8YoCaC4
OxKmgK7k17IM93t+10QZVK6TRF2RLlaHURtmglimTFD1Kx0Wx79o83agR9ACxUcw81FVCH+4CP6y
Gmxm8ah/d+lDWcN92nLxQXR/sb8v2aWGm8qcSp6Qda1XZp8yZ31WOcjCarSM3UZaAlglygG7xhkc
QMB2RQ7CltSaxXf+DiGX0BoCZoE0WFpKbn1+COrOhPl6hfxgWtnBU74TnewV9GQN7Lu7uiqbumED
BoFwv6kRqpaqdltDp2573wOrV+cfp2jfFPkgRbc9Iz0MQvZHRG0Zy4G/FfACAukIKHYq3hGlQ3Jl
2wbhYkqrAirp4Ujrw0/EBimH8yaiyDZmiRWVm+lHCrl4OrHxN7WtWlw3ZbbrD0eTmVUPkZBzBaEl
S+xOkbxQ0//Fjc9sgAtT1zXjWcQIdhmn15SKODLzAxaWa+TYFONaO9iZudR9KL8Yrd1rGzRrz4lC
LeHmOEnZ98gITritYx5znOpyJQa2GzUQ6uGAAgMQid9cSgkMvsPliLGWwVcv0hbjFyONoiYyuyC2
qmbrbsdA1Im1eQO2Gc9l3JTMwleLc6REtaoGNR47O50ZRHl5ISXXPdVTToifKSQxyl0ZjOD9DATF
IWhOtrAESxrtcqUJ4I/XRGz3vuGHswlaurbvaq+wTYshkb0nrLUgUjLHB5Z3BGF8KZfUKd22Hj+m
coY+kbXCF7t4eiu74TGLglfYW5FpkKHE0xZ8AxJJdj7LBeC6cgjwP+/CapqxQCJX52+1i82WwCs7
+hvHVlt1ZrIg8WP/E5JalsZ7/vPXyCgpmLhPoGmZrTPkz0Ofii53XPp/SQfMw0ipKfhzhLKNldge
NERsAnM7zy/+J/lVOI50dDshQT5Ts5mqoi9I8/kgZ/vgssqn/M4s20Uyy4LFgenY+Dn6uT0gCy8z
5HfX9+XxYFUzBEwFSfbMD5lwoLdfIzKK4DGH4pYX0a8sbcmYauaZ/cZ4ZwbQflsgHmOqDOhLgR4+
Nhm0+W4M2Ub/crDk97KJ3SidGaGE+xQyy0FZL2kKyq1v5glSE8cDKIKJN/a7Ck+M/Y6gcNf0/6LQ
7vK7OwTd65p0m+j7Mo02fDsxSbM2+iLL1j0AeoXwqe+Sje3+HMFKvC25/dzGwpWc3vh95rjNiRTi
+8lKrnIth0DWOmdOBrkh7O/WlwmqGnZxDQV3K7l33u2KSqmhQNEvJGrH+Z2787KkTmPd6GhueBny
F0emEqOEJgWdW1J24Mf7FEi6dHFF/azIUaAoc4S+ZoVfoweFsR9HXcaq/0l1E0A60uUBug3bHxP6
D4CaTLTJEAi16dnrZGpPhfyhPpjQNf5xLxK9oR3oUOyydL1PK3V4SlAyJ5IGkA8O2BOUa4hjRXgJ
ip4VUyVeKij1GlSX/fY3gRNWe9VCXQvOQTP0yxqpRapqKU9zZYu0uZMq7tVK5c9+yymmkTaHgJAB
TT+LZ52joHlFifTbwTTLFljgd1Z2kTmDooTAxFJey7/8EoTgi/k15IqfI6LmIbkxJanWGVFX+lDO
HIhnCUJLm2KhtufUm9cr2DFgs7we9sjwgyHq5hD1xvznLqFYIOA5EQsfqsANB5Pcc9ppH/JjVcs8
QCu3OwbFvy93ZVpTqG0W1tpEfnsE1zjD0f7kcGIHWnChmL4wtccjJFJ39nmG7V3rhJJCj2GlrhhY
n8eMunYP3xik494QZKgkrHV2ySpSUvPayDwA/qySXFtUYVePR/j5UYfQ31UVMlD/4HczUnaUZcXi
OZw3zTPlv3wosdmE7Hn94BgwzAiPJur8jh+RBv1k9v4utsemAnCsNfFRjDKFPvWkdVN9InQZlo42
Vm2eOf6SLxKgL7uDB71keoWXzSXbeJ8lMgQluYzpkoLDy22HiF/AEzdpnyQrf4NzluSaUaL3dGDb
K9faZaFVnK5onqBTS0AEBAX5cdP5q7hSDY51dwtALagcC6hr14G5a+MY1Nc9jQHPPDznmAcOD5mV
fHSyzz63d/bvgwQPfqOw4Zd0uU18AQNK4emGpKaEDD3NlZ6H3WlS9461c8wLSiGZj+MvkQChIKMA
f3O/kxcdlCf9qFGScbOy6ki7jqJAEzkTHoLXfYjfzJ6ewcEcVEGMz/7zv1WT2rNARwuRMVnrEmyr
3c8IGlg0qdf8+u0M33C/z8BQAWOdGbKpQh/lkxGJ0digJ1bMokgqzL1BIy1W4MQVjmfoSSAHaZfW
CC6o3k0tVCmB+IzRSkmtGXDS3DOHv7sySnjS0cphkTgg6UplSiqsrdqJR5T+VqR4R34Zp0wEqzP5
U2K5QNlHMVtmdcR4yWvyLM4v1/jHd1mtvoizdC2VdK2c1U9Fe6cKzatqPKUdWKOTc/RUFkHg3n3x
rZJ0kzkCPL21B4dgyK8Kw948H7OHir6RgqHs8SI8lYEC9HSpVN9owY+52e02jjgNJRK45mVOUr5V
MAW0poftTlLlxYT79Ym2+tMZHqqQMIV65JqBNN8qEI8w9OGc3Ug7Kil2fXTjDY/wLqMu+SbWpHmI
O0g+HvuWFK80lQkFu6Qomc+ZXIXj3Vp9+1B4M8C+ZadyyCpYzrDmQSOzbEtDzPSFt0BkzC605a+K
0kRaPrJRakK3FXM030ZCXa1JRtAxDWpVXbOw8JDtWShlnN44AS4jNqhO06troldMlGqudrtbD0y4
RWAruBHLEEgU/wDgXf43hJfdVlRV2oPEHYWXKHwG6c+I8XcpxtZUc57P/dUmji5X9hODbmmNmTy+
xUQ15yAANKpXHGxM5LO8fTXTax0Y+a96P79nYY4Ubi8oq3VOk9v+l1Ks21+gtavpzXC9ry1PkRVV
mVZL1SrIM0rIU0OfngdC4LZRuiO626hq7KSWBgjgY3TEDCcbKpH3tcjYmX3P7mg8juok6eaG2IMg
xcB57V8tBolesphXEE92WccOl8kHDWsL8msmlNG4zgQgNIW3eTfLutjCF947jXCCVAksko0tE+Zd
bNtDGmzuFKaiJg1wWSDPOL+8G7gqTEYncPKu2Ng+PKL7iMu+IFDsP/p2uWoKB+COlJrUAuFshsJJ
gxyh/mvzxHuBDQa/SCcPwJdxD1dAuOBRWqB9CfO4F7GhiJi1GwHGLp6g+amlOmvcRX4OUVga0xsP
43XLeBn0HP1N302gay3xeFPeINIZIWVH8bdyDTChWv73MrY2yjcdQI3XoogtIQg7do6LUXJ0t22S
Q9+4ihCIoCDmJT4hPsGbDvWOSJGMIzMMkJzl9RjRB3Jl6XMxWiCcpoORY3nGU7ImlwO8qFz1DGE6
vclpVI5xOM5El+4Q5thdtFRSf03yqQJkGNZPLSx/WWg8xiTTAR6Vgx3vuNtdoNbr/XG9FXn/kp/Y
x1ZgcDh7vbtg5bWzSeHhjOhdBmRywD7Ou3gqX+duHCfNYWMtQ8izTunk00ELiN5AkSlINalviQF1
LS8Tu60j7eBkn52ClVQWuG++Lxa9BTGhtHW8SyVrLbPY+955r/jHVZZv8nkOW2AmtsJA5nVF7my6
XRxEjjJ8l7DK6c6doIqxbDg+D9MvYZ7BzBOEeTTKT6qi0wt7ewHTICITtIqYTip7C3Z4elDNCwT2
7gySNy/joQoMNR0dyJxZeDPCacCzqbVO2IbfXAQ3qMa8znKVYVQJVmlh35PTV9z0HQKxs9tjOYno
90Ak/RJH9zm+2k5DaquY9SYLt9gCy2PeQDrs9tRvAkepD0lTpwUZ9Vek3k6Wjt2rel9KVtQYg3Pa
fHB2KGP9ihUj4dLQ8OqoubVeJmKVLm1oCguplIPH6FL4KUGGW9LAyEc/+VKK1g7DyDncrQhMrBZW
QlsvUn1wzoB8Czv5oEMV/co/Jq/YPxLzl/EONedyYOlwzHw47w1BJP+0mAPQ9GFnxKWGr6G3ez8S
YvQhUeYPPx9HHyghqRkzBWZDzjAAHyyYHDy6YMk5r6WY2CtUNqApQIQ5IqoweTAdcEbHvOwPDaNO
/5YRAqhe0e2byLIdhcWUw7JmDYb8Wm4CqkZQeeiQf7HJmwbWWdUN5ZoSISUvbpEwLEdhsVMeH5Yp
Uk9MMBOHWQNLnrv6MU/ddSWzZ9cvnDdJY9fGu7QBKb3QCU/thW5Zc0EWrEZCjw5b40Yq4/oSC1RE
ggRC37hLdS67joQF5DjxpJUm8siQlSCW2DwT/E5NgqT4384RXom8oRaMzdbP7VGCDVCMCqMni+br
sRVbXgVPV7ktbAz/8e5qliCze2lmdJ3XDbYPKhNzhoDVSqIcJvjYJp1SxFZg7+GTNlZgpbSxTFTQ
HYhQFYrmQnwVT6bcswm/T8jOslZ3jGW39XbVxAfOxN7bN/ZJE6/awH+2jUCgRymCLO6Ejp3ynmWp
DwPIPeEyJ0d6qkWXF1k+j2Ld7KrC6cpirFo/OCisSdLRuibmyUhsnUtOn3mmhnry850q6PAVWB6n
1DzpH/+jakS6yb7NZvucens4co/x4QgA4kIZub2TceyHVj5evl1qC/OhjFTsoDAb40a1sZmgd/Hl
ysZ9jj47b3fQXNVNoPAFgYgUZ34pCMyVeT5R/3kq/QQp7PziymMTKq8xu003bxCf+yNJE5HlwwZG
CCxTHixrp6Qyjay9TuHLEXJNRuiOoMpG+JBT4IopoNc4R+pwCTPzpZfUTJ42p9IurnrXLeeeoUXz
HmpWKP4NDmwPOur4BaU85A73qNQp4jVQEXttLIkLoRqwsUSrwqnncH1EKnjeWw8Beg0Dr/97P6Bt
aKeB6GYq3J0Wds7rUaL2H7i8v+oUqeg8Xs1XQb2CV6dP+frvNEGqP+cCImDGuqeaRjmyXOuJfeGg
rToDl891VMG6aYXP8WDFNlTe7NQztpGrNV5y3yD+9Byfs3JA4pQV2fAgbgeEviOQAb4+3JXd5KO1
TU1F+yy3URm8BK6bm5v1cGQvoObb89k1xgIKOSdGe/DCifzJ3Ahf2Bfe4V47epBSDj1HHyB8GG/n
yXPjrIsfglIlTu02IKFHRnm1gNNAKfgfYj7nav1W8WZlyurUfv7z09FPDcuvYrKoBjMa2u3ctYBQ
ReQXaepAHkFPDz252pPpRCeXPSEm8jJv4uu/4ygVrId88ECFJ0xie6dWRLTT18RDSXrZZZ0zUvLt
BJ5bQTTld+mt7FhMvJbVrOpBAFAEHl8Llh4gEZApaYPfah012q34JHs/RVd2rcyOnu+xLkRXOqHh
6EuQeM6sLqRAlNeZAjTeY2VUc+PbfXo16VnQthTbvLBmBnie8Rk2D8Ao16WrodlfZSUfg8oHWNMq
ygK5NGKkRqzHIZwcmPSKVOI8s6OXfp5wPFrAd5fPKoY1yLe4BwtuYvNFw9RSoO7jDo9DwBC/RlX8
oZ0TylzAjsx9YxDTKXeoQcgsGbf5w5pY9hlFlbALoOWVeJ3hsrlldxAquyUMBqDnBYDgowmHGGHt
00cg3neZ5f/Y6kMClm+W+rE09TmW4iKAiaZeEHtnKxUEBZI6o7ABDo+AT4/j40hpG179d+Nvdd1v
kFQx6Tw29Vty6N1H3iBEgR9F4ZblZrSp+xhbJyQ8qzFujxbqJT2iP/M3Ku71mHskdmiXUzX2aVl+
4bUDznwRfjOy6hJE0sDSGcUzYJcP4vPiGrUS6d41x6vbDM9yfKlkVW3z2MDYgCEbGA3RP3Zs6IBA
qK869zWvtUETZ6f9McmetZAvx3ZodEUYFF8k8/BXqEVN0lBbVHXsKsNTmoR/UJs4odrwd4sFDih1
nqb101uky+eW1OiQMjCik+PQU8MDOwibDIg0Mn9bGsMfOEvjAkfwJNyOoB7QCBDpuolXpsXfgrML
z0SghOJFVbXC5Uf9DHJvbEGKtup5Gbotoe7yxgecEANpF4VY0p9IrBi0639/IVmG3eySD+x8aLRG
jTjoEjn/sVuier2vcZr6KbeBHDyY+Rc5z+wPzyZRNwQ6+Tp7vwAWq4jaCqGfz0K0OsZGS3YX8xj/
UvIoAaczq/kIo9FznrpUAqsnwJJ2ZNtQnk6bhq3AiIxA2cmoNbFEJnY/g2o6XTWUmDyNEI82su5z
9p9n2ol8AOWOv7Bt8oQfGBCkl5FsxeVig+KyVRyG7hflzHq/HCo17TI0YU0Q2Q1ZogppyaeM3ZZh
kM+Hsx8sxbgR6b4UPmlqV9zknZ2eZ9qdbXK/TNsA0A92Fp+jfmbP5M8zBl6U41+yUEA6Q7t23f3u
pgMw46ab/9weDQ/xHqSmLb5amq6U3aNccLyMr+RSU05AdCv8sU463NlosXT/aposn0atA4N1/iI2
A08WMDiU9q8nFc035iqOddfwpxNv90M08LUOsJz1EQM+NjW7XezMQVe+9v/YoC6CCLzYnWca3zCz
PqPlG2bqoKGfgtbNzIF0e79wiX7eO0upZywHu09XClgMgM1XK4mOVIwkzcsWmtMJKEVrHvSHU31+
LujrwQ/EkjidNiDeNOEjSwvkC5kcMAlgvkWsifmp9xZs3mMSZ4NVxVo9h1LRjwF/3fvt+MeM+O+B
2eV5hR0f4NU3Jf0tvfTrENNh3qZHdtIjHmzuOcYlQ1mbVwn8TZ1R7NSrtISIedL/xvZ1cL1mIR79
Aa/MSQk7AFOsu3E7NpvllE3MoG+SF5p7UsorJOoumhGIgSKrj9xN8JmSGgSwTCJcRQfBz8fuKbR2
y9LiC+ytdOFe7sQ+OGUUwJ6X8SG6TEC+YB0d1LgfEKubaORZFKzSpI31AI+TbcGMYA8G+8MmSCJm
SKYMNyTZZvYDZLeyc/kGlHKL7GXuj0KHXzu23llZb1AZiORgPbmX+jBrjnP5JMuXQajgraWzLnpA
1KW4A+P23VHc7e8NBfTlAY9SWRt8HGAmiRSaZz+sH7u3kDYSGjPh6D5+FlEVoTluyk6ValbxVVG+
gAhBmmzCDDtmOalWjqOamex2BRwBQAMaT1TOO6GBr29CvxOYDWC3EJ8L5jSU7pWdDz44tv0rr6Ak
yc+qiqAQ/EmonzqSz+Y5jHAnRhiaRMPgS91Shji35FigCo3DeLSkFXygjeA8dTXNUzstPItVyked
dK9S0sJbHcJIUriyJtKL3VgmkmH5or7S1Ncji4eXuyiIcMbKejMqWO06F/EFkoQvlAsF8hTl52VZ
BKrLlUyLXhU2tfhgms68dhKxOCG8xzWhHCbf8u88dDBqdzLbizixwWCxO16GgClzk/pZAWqqOhbg
UXRnPcMfuMFh0MQtivqoQ6vDgBoogib32ZJrAW2rFCkzFUisXCtcBFKkuNAc6XUmZeNEJSJQa9OB
aDmajiWPFcOGIQIkoCTXzAz583eCgkK1AFDwCKlGVMhEoKVA+/qBKU2JPCJ9etscVJr6Jwgl9rY/
rqB1y9u+C+Y5omC3f4dYZh6v/bAta1h7rOi4bGuYcxjc69g2o7W4k+vbTVj24dQhLHq9GyZXmx+u
06oyKN4icAQrpu3GNpdTwqddrhfpkiVqniimFjGI6HXY7c/17drEMr/9U8xOdG3OjCXS2Aay78D4
TIMowTy0QBPz3sQqT76KEN0BVTvOXS+HjeLqqIQp6eY5c3vyV/YZDNQ5E9jAD7EHEQMfXuniVunp
GGjQKaMtIsi/AU5R1molVGLpvwpm6hZw9tAaa1dDwHBUM6qcPaPzE/hr+7RZ3Q1hiiCiOwjYy2yU
SMUzw9PMyKzdWRVdOfJ4kTGXiSMfd7WBW8UeEj32PejTYgQZ7WMkAcf02D+S67TG5kQRHQkRa+9C
9S7hzSblLUFf2kKigaM4dds6PvpMYeLwGIkhBd/fHv8YADuD7s+rxrjUYEv3Y313mPoE/TrLzq0a
KaB+r/PTU0Y6ElR+dlDjsg49bHbV/QgeERUqoSlcpZBR7LXe/6tlgNX9tA+pOkrHDA+20Kdk+aOL
udvUgX3Uc/KhS2p0Ml/BaFfbmSLRJtW9RThM163iqeRNuONIJ+5NKIXE46IimiqYkHMM+y9pFsWG
qPN51rfZG/drEe5VBmXegbyiSu37LjrRc30GAJhWIqVUTxX82vuxtumFoZqxculX+kInwJ/YrgYC
YLEbhw4ANpGywkuwYc9agNKVsr7+OGnx5qHui015+N5G3KMcrNwIa+oN1wVYbwKqZt6VB8oCyX+m
SbewNmypdheqGhFAxhMlhOeiS9L7Zi4AUS465RyqEgfgbztFDvLQvuliFvcMyyfmzqwz8rzu69zg
0RD5tZd6DzxbQCx6ruc3EivCJk6tnBHlxXO8LGouNUrQfBz/oCEvEF1mbuK0ZWWhbgOb35FJy6S9
ihjiNY7sd88CHEoN3/mx1ixRPU4+qDez3wGOxPx31udS/ylSKU7UVN9lRCatn90SVXWUXi066HrA
3AIwQZY0Qm7z6R0nexxRgBpSKjO2nf1w/6/9dkR0kz4KhYSusk84yNgn97Lte8sulrKv2bL96yng
vUK6PFAXZW5gwcG++CSKl9wAsnxISHZhF9p/QgR3dPt48hpeowxiIOEgasxwvdF1iFCSQq6R90ZS
1vLP0NKVLS6tnBFoemt1PTGo6Rvo8+T/3hviuji+NAAuNlkZwMASNbiHNb2m4YLSCpnQhp2+Etzj
s3OPXRRtPUbaKZgSfskwbLDQXRodpn/G/moVqKql7uBnB4qmO03p1tnyxLyyacA/bh4uFD7MJyjd
R5HMqF/7+fPT8BZhlXaEnk3Q+TWy3Lblsu0n52/KrZgSu9kArA4uAb39PkVz5XsrS4ohpENwUNkR
h9nIfX2CWe/1o776DKG05yGWRSbwcGBF0Kzz8xZO0hmMwdVLK9QRG2mWbF2XyUgYnuSsTYe11Ynv
fm7x5OVg52HzqZ2YYopq/WS3os1s5zuNexhXq8AkU1f3HIZywo8k/oxnXSzSrkEtbPcAqwuDcsBV
DsNwbc1JrkYJKd3pJgFQoJ7qm17R5rVhvOs41VIqPP6LOcvp+y3ueyS2sig2iJ4NQDR3bWq1GXj8
z1LRK15sn2kW0BZnvABcShRnXED1JZPBLwl4IIf8LY+krZ9OieSFVA8oJJPM/9nEI9EpMp175/Xk
rbtwyktxR0H8dAusDBOis8rMpy7VlJk4bbBJHgZ6zJl3wL5KgPoHdnF7n3214AT0n8rGujRsUiGT
OZINFhYh1JfDjRUWZphzgu5xuze10rkQNpncMYIZ7zpCqdpE8rRzDQJaJif+7tW5IKv1jQEKIsXe
V2rrhBAZcgwUP7c/0j6WtsKnmLcHV6E/KidJ3RoqasNc/1i00WUqMj/b+9VKJuHlsZZwmPHhFcyL
wqb7p4Bu+aCP39OJCCjOeTVfHVFN8BG/GGoEB8cyPxSUQobfqjjKlmFMw2qiMtU+0OmdT3j4JN6w
x+SI+90fqBf0f9C4gQzSq5U8clKS9l9aS07z3hYm3OjCn2Xv8Zd+16Q8NZUslpXa35FFui85nmxT
AFqkOVwP3vspUsMrG4N21B6QRHc/FMt7xog6X/OgX43Qkesc+Drw+UD31Ja4PVUy4ZETpz4/a2s6
/OmJpAqVyIkN9WaSgmausMinDL8QQJAWpCAUFfwWgGzumluSHf2VLoKw5yksA1zaxN+q3LIrsBL4
5HSfB/dQV82n0bZ52ONb/L3mNJg1xsbsHne0iT5hh4NEkWrGqaNKDg7DpUUZ60b4lj4hiosBC6h2
1jzH4JIbXF7hgl5T/TlS61VqOUuOdiCD3A+9iUtZqh10blc/2Ytxfrfnndckm93MiAmthxjhGmbe
IsUBGv210Uaq5peKfOVmkO4RiNVvqYRa5vbJk54GWK+TliVtx/KOWZmSLPVv0RO9xh31l99WlznB
aifkjVKiDFhASFAr7Y9mzio2WXoRO/IFwdJEDgi3CztsoSHtZCNnSkAulDXYlTPdJGj1nHItzX4D
stiWhoKKuIRm1phVks5Y0F5BOE/vWiiwEHwq7B2sH+cU0WHAdhvuP5bdn8YjMbHnu9Yj0DPPzQ4x
WoxSHURplrHeZEjcuVyQk3BO2I2ZB2siaLDY/WrZD6Xzx96oYrBaKH1HraBX8JACLERrDtawS4BQ
/0Uq3w+rgCpwWSNd66pmjCuW+cCfDrBHy0bvZqOQ/EQel5OvTO4fy9N8nVsTWFE1o4qmeXDFz3xZ
LyRrRsW1YbsqqNXxjCZAIb6PLUaGZUneZ96b+o7QtQMjMiawklWXtfIpC6Ew0mkhMPYRA9BWwuIA
0ZQP/qs/d2qrDuRhDHJR1E8sX/7bc35afU4Gdz9XIUdRXl2srxiJphQ3WvQYNwM9sjrKRB+ehLoH
MMviq1Ssdd5GYu5+FIPbUkGKya//plc46545q0dIlSm54U8gn87ZOfyd/tlqwyfWH6+AAQPt8/wu
bj4vzKY5o5RoMIxIQgVlnqthIVvPbILk5tlMmnfCRMeYS6OaF6TkOC/tWdX73D+uq2YH5DBubs+2
kPzaQM/Of6+hfld9IW5iN6e0EIbFfNouZ6w17aYOyqg6kuHk09CEQisfZ3f/nlMp7UFObrk3g1Fq
RPyNbjV+pP3iBK2XoVaIeJsevC1dZlcJp8xYqrBwWVXsFXcqwLVfm147mwrJvpxu1nD6mK/ny+k4
dvoBw9cCSKXab5Xqp0Ps2t/if59v9anygiADMl7uIwHAwcybeb3jZN67h5HjuB7OctdCN1uNnWgE
t5g0Zm9xwXH1Gct2cx8F7ldTVzSmsWuC04Ju1dNgl64O9UHSQm0lA5XMG0Th0yeHPfb8s87xAXQ+
7NK/8yN6RyLNZDQVs7wvg2hTkoe03WW+wbAg6Wi9luaN1RPdIpKTRNzVtYhoEGEa3579NjcwLPpC
TT+xlOVTSgcHWMZEZ/9H6faapG70zVTkM1976DRpfx5D5d4blfPEnMb1HrhKCRuSKzeNpivN3ygs
PxjSqi8AxfUeTtz6D1rWinSy8592nfsKcDPZLHp1ePYlb5qy9yfpYd1VHNK3ITB0yVkvmFIK5M0H
0ub74z0CGgmCLRbZTWccddccDHA/EAklcK4nNXBvs/R37M0+d9fctcaknImE1Ekbz1AF6QhhSubO
N6nJ4N/r3zbJEm04UgnoQ6u2P6x60B3z5RRKkvoO1mwA1m3MSufy1Rpt63Wr9e78WaW4Rgco+y/r
R6Dqr0FUu/llKg6yqSlx4VqBPlX/szLTwMw7U8bIOqldopjYXYWZ/mwJ7pH7VSRW367qOmU8uuK1
OanEjdxo163vIfrHpIo7K1myo0GsKu23Jwyr9bgPnZVrv/btEQWerKKO8Jcew18JFXKz82YJiaq8
snUIyFY7MQqIJzfHz72MTkIOuk/fMze3RNVE7VLfazLilnGBGUesYVO7t5W8EQDF0smlGtiE35b9
PhQId4k/3m9Yyp/vhA3ElQHSOz8GYHRmGS8d3GBZ7kti+kbwOfyXTk2WTfYL9ch7VINIMFCQB43J
trsLzA+EbgmIZZrcFNyloL6srQayrhpjSkwzabicQeG1sK56F4uz1exCLFn58jbvbW2acC8+DYyg
0jAhzbwun2DyCddx1B6jIr10VwIFNAGPoPyToivBi7ymjy3XkPjUMtQ49aanCs4xPJcbeqwzrkhM
Qf2PX84g+2HUEs7Rw6bDEnMK8Usx+uO6whPBySUHpbRfuPp9Ul0Wu1yBo3Lr2Dq8oRF8Xi/eu/HO
zBRbE60Hn2QUMJJZUnIwkw6M1UdYSSAZy8QzEroG89L+rnTII/rxOr66rHpeDHNpDJ6XzpU6F2jY
Nf4mzjGQsI/ktx6crispiQfKWbvz+t9Re4tMtIVN/sJTtPyx26v05IhgMUXL+Q6Az6X77lQHUkI8
onkSxWN2azuw8t4MiemBMnAQIDaqpJ80RI0xqbkAUpOREuEDtqca41XfOuHkJWHoJ9XWLuR7mjN1
3K+CVsdtgKm2iq0KxewkV7Do+ov+Jj0TaZxd8cnkl/PZ4D28NMBgvfaAkVfpbAY2DvB8lqWoAgOG
p+DGV3pEYrONBl85ejZmjKL00IGHzCWOB9GM5w4cynJyxu5wvfs8IURi76EPVml3FKOBQOCyun6Q
BqS77/TOqxXpv44ED1Nxmwee65MMs9FIS/MesCazqSq/JzCyw3rs4P5HYs+VPyIKsmjvEvynmBh9
eoDezx4a+oaSNrbrRpLRJ4Rdl6T5WY3ElyRkeUDe4x6N2qpwKim+My4zUY9ZysDAxZnNZp9EdMSG
NKLavGFOg+TUXlkrp4opYXMbmybDTW8/tIFvUEtfLVbwYR5zUyL0jr2wnaVgE9/sQ4cClUD/Cqk6
/Xl9EQLtPJPwbBN4QgVPwyVSNNeD4o7sCVqHEYgfKPHeNq6N/j9Gzbwl3Z//nHaC2k3buYUHOqGX
X+UA7NIviy9sPWlDZKKGvBH20NElkZ+HGWAOBaKdNlNKC/S5JHTAyZ4qVCgPfAlEpooZWj3DWxDH
bcZ8Ctv3bH/Mm3tybDav3UARB3iV3ynqlhC1KY9mFZckzg4Fdj0iCbB0Wua3iwtC7QijoKcJPptP
1x3rM/QgES90P6IZpaWZRRlmdQhz6tESjXLakabPKS+ZlaJaaAvf2CzNhu+RpVsPXOkMeG3USRVn
Js2gPNXuayKMX5y50Srx3CK/TIBQJrW+rBmz2UOPFLU+flvcVXeVqeDgvLJGpr39Ud+80mvxkAlj
2SOLlzSVRLk95spcdpStzyM9AeOCFbkQG1KKy3NCX0F0JZcmWeo25TC5yJow6KkT+Ll5mIkfE+Ch
YDVIDCfVr0kUx21tq2BSgYpNgHJ/j4TBlqYvzVtNVJ4t2PpFCM9PnRMzAnp7c+tseLZnH18RHOrB
BMvx1h5Nl/4bDkq8krhfPKuOpLRwg8k58PYAqgcqrA/hKSYAkQXDIFnH+9VBiWDRmWWDvDAPV6Ma
00ofECfFxPHv3bb9R/pM/InJ5QCbs368yF4jYpwN3czPv2GYHJbvuGugT0ze+GqW5ZOSO0re3p6S
xGyJEcwEYK2nUQ/mr7B+qtZmx0A8QeyET6wMoleR/Oi2Cc9+or6d4QqIaS0sMspYJFJMYH+A9THa
PPw8rFTxXtuDYWjZiypJbDkhJSHiDhydp0Xsbvsb41vimqS5PG651hhQ24j3dW+/CBn/9BTCCE3h
K1ilZnMiSx+b7b2W/DNLxpSBUlGzr1i1sSCzAhNK99VV8zabGU+YO2WohysQJ7pUhi7d7dPSVr4J
wYc09BcijjzwTifm0n4/1sLi9KyiqvHcO4hBSw2pqXCasg3unqipDLD0V/v5mlmo5u2lf2uqhGs1
rNLhMIx+r0rf9JHurX1qt5INGEmlZawqLBlBIFKKzabUEVa7q5J8MtYWOstZNCsP1rvH9Y1OG87e
HSOgplWUoM7g0euDGY9j1lM4jFBAZexFIiReLJ53WX5jaozvRpK33askPY/OmfwwoeUkrcIumfaS
kBxYXPqCtrrQNwQgipQqn06ixdFpktNszNq8DaWcrg0cgmyNZyDCxgsjZc/KHcU8//A+lCFsD+W9
fiXdut98Vn36w7alqDWtSUGk0S4roLbHGB0IqTwEFGrChJRCG+0FNKYBiFjzYDRzFTyeJ/sYAboK
2l0PCjYGMpwbLLEHlGqCWChO0+QDXpJDh5u4EnDJVROQoW5CM6wXMnelIEvTpcCQ8LjLVMG0zduw
aK+5hUYlUkkHGPJLa8lHFBfiupz2fVuzW1ZIJy3/Oruz7zBEoG+mijIx8lVsQjKSB8tvKpS3XKnk
OOir97pTLhUZgdfOXa06HisrUAgpPfEEkpZi+ov2XP7Ntj6gETxUYoqkPAZntsivXuzVnVWymd1y
LRNpnpbqmCsJvNt/tF1SrTxBaUK34EYepxhJmS6oG9loKzhNzNpt9LKrajf2ZObCFAEeGpf2To7Y
fKZqAH4qVO7KRctastTwL6KbW2hbXVKqoRdvC94qvs8b9PdPZNYsVUKiW2hKxld1pSnLVzlDvIC5
6dihGGnl7DWfomBQwSQCYWkw1KJPZbH6aVDD4B+y+1kpWJV267EHg4GqGpITsxSyyNezPnNqroeb
uQwnfvJLaAqTIl+eyd4aLxkBbjItrpB61jjXvAcXCSa4G/paiXxnm09NwHeA/eA1mp29GBLeNqKD
hevM+ZIqUXys3K0p3tu+NtxxYjf9CuliDpfzSmem4R042iTC2GNjJyGHLwM4FF9hN2YDFHztyuWc
tiEBIS3Kw+58FJhR8vRyS6BCiq/aH1A9shLvwgs40BuCIckOA434d78ZvCetXTJwZxWMsCxRTCEB
5854uCutV+4bMdptfpb4zxqwUN2mF9VxMxK5V7wipsUXU8XYVtbZUDwBbdTBNb57sKSu3OFPupya
FId7Lx3WC9ryi6TgCFcZV6M4FkFMc+0uuMTrOk1jYfahLNCSxcwyKPvOztaueKqE7Dn2oVfnI74U
iCZwW2LC3cZNHH0aF+Bwn+v2dKIz7RLRJtjPgpOpVz1zl9qw07Mbs6713scdftPWsXsSZKfucJvf
0+jzXJXC7hKPZOhWpdXP0KbeW+tarAgLgC49P4LEx1wWZvLvAMp4/OEY/aVauDAQmRZzPdapsdWu
XVQy3PTOGbHCQqcw4ddPsZCVHah6UdaO7rTcZ0Zd40FaVbkVX5KjgCm6RcQpt/fw3FjgFHxkTPve
ciDjsDUDeJ4Ki1iwu1gai40tqe+/pfy7kdYoQWYnlsx09LWH5EDbuRMp5S7QL7ElMj7eLGBsHnk8
v/gWWzBZM+WuUjWLrnxHUeG2S7Lbb6YUeEn0o/geuVUvT+mgubAM77Xzf947f7JmEir9hNzWgHk3
aV25scLCm/gXd4nRmeiOfU3MKRiUZw4duHWZVZrF6GegQHbYMp1uKLlaE3AVjs8tRtZThhqXdR29
61Hw1Cw0xiZzWgoQnV3V+IWQFLrvOhteuZsgCm6tVe1D7jfj6i4bg3imMlLKnlvAcOHvAGzda/Bf
mEXxr45RQz887n0ZYXK65gyO7oMR3Cn4GdbOAqSJGyAkKrfFZQkLOyh/FtURbNb97suIsp4WaQaZ
8rgW5kO1XZd6u7hygDDLoOit+g09aDI0kUK2nofbHdYP1DDUhN2bUCUlxhiFwjzgkLpvmeg2G1Sp
vtF8KUmrzreU4VCua8N3qu8CSZ3p000gGHAKTVK+n4HnaT6pRx4VwqgmTuZT9u9GYcyTtbmNxygc
1iOYq5qUHP1rEifHSO9lc6n9iXj8wBsiLf7BPt7POywGj0C/EyVwUXdj7gU08IWb0vYAmus9DAn+
z3H+zza/D294SuVru3olSBOXJ+ModIiI0uqcKd3y71z+aEgO8Ru7TeWWlCFlODtEFWpMcDAK9Z+H
c1uAfSAakWQn8Pe9Y9qWKxbISjNs3PS2dpedQpH6ML+Zm0nGhjjNbGz0CjQUB2avEb6LoUtMBtLw
NOd0r+eQm0RlG0PBb8lnHaGxBzHR1uTavYEMz+OzO4AGfBZ7Pi1HQUGemKe5VBEQFRtYflBV/zGp
wEJeQvnL8uj+3Nm8NAnZYvxy+8hY/TCSpqy1TLRvFRdc/WwafgtqFBCeE0zweAyLmHGZlh5jDMUY
MWFbDCVztSp6LsZgOxg0WPaoWmPODrhfjJ1jWtssGpU1iJw/P6sIGwFsZp/2M5mynF/otegoI/pS
y7Is5mtYEG6C9jePuJ7mTSoZYOPQwhaUfx0ZkNQuQ8+E1627r4f0atITdAmd/1tknrqvRIcf77fP
bx6lyPpLxtP96ET5/cOOx2HKww0G1ziIgf/ZNA6VFJI6Uv2IYLO+/HxvzAldbVQB4DiniP4GiSQ4
LO1T6UCHmIWkyM6vfS5d6a3hRGC4ylvzyx998NAwa5TTt+tRe6byOn9j0Vh+pUAW6VRefPNfcFHL
e+4ZCrQEnE6h9EKsGhVKA+86wz55pZzybi37WRr/wIYJmyMfet2Mkqj+qawzcGKsWTK5h3zbqQC7
CRDumJrgxEM/YBIUHfOLX2XQT+cL7mkGmVFgmI1bduO5Wuj2xzD8LY7RVwpfYbc1vyn3iE3IfUIY
VNhr6OcFQ88OjIO7d+77kZD9zs5Lm5h3TxzAp9gY3X9h4yoPK0myVnnw11ZuVhTa84O4ARlJAnLB
PjUER65l8LFdePomADzOj5qg9xIguogcULCHUHd8ye2bFKIYS5yLySNlG2uI36SZB0n4BF2om8Ih
dZF8J9V7lhExn9TM2Kw4e1sZR0ltwX0hnssTQm9QUn1C3mL8edmckMg1tODyHaEO1GlspN28sf/X
tZriev5cTL+cnDrV6PJ7OWO38kjr+JCnx1tvYUy0J1k+W9UeLnZyXmk443zt16FGfyydV83j3I9b
ua+7vsngoiAY+BWdorHBmEbLWe3S/WDJk2lGMf00oFXtFpkZZelWSywWDbEUtHGt1L056fqK005Y
7o1Lt25AXXYJWvnxUyeeJyamX2ghZ+7EZxBFlkYKXVarZryucCRU3TUKbutHEpRuWzg3mq6q5gGf
Oe+R9QV1JB2rl/l8noedoMv5tREgRl4yJcAcF8Q98q39+u1zuGzeEBS+9XwI7tCux/ncfdd6aeyZ
+YK6bgCMvaWadi2GvIRXOJ2lYG1re+Q8ESjrNlxzR93zwmfTQl9DPoJMZ8aqQl2lxq1iQ/5LWK5s
mN25IWyCKXNRDkdJT9ff4SfphOTkou/nr+pmws+PheKC5R8twYE18CAcOiiMD/NbPjQ9EPFBo4Jz
aib3e8V/XBy7F8xmCd2OJfKxyqNse5t0gyC5vKfs/Qy/UM8ZbFiX8uOSTj7j9WocFb7v1Stnn3ys
6GGfG9NMnukLG+b7D4Q5sejb1VYbCntvpQdLxJptSIOhzk9ZeP9YyCRwDgkRrLt6N+SAxHZXuT0z
nyJ82ZcKTCDIQ1hTWADQbDXgbrEGu61W1dLMHbpKFpAlAyCt0b/UVj3Hql2/2Nv6AlBE84GJbLn2
MkxGHtbhTR8S2iwlqYIye/O/h+RYms1hB6vxOn2G1zTof/ajTB6LksrwbF14hIojP0wwg6AhPMvY
Soa6gDB7Z7O2COh7b9BmGt8/UI6/e2W9tD+p/WrIE+Q+QFt//gN/KYInp49Vik2R+apJJGCaVOfv
jR/zSqZ6d6lhoDjWODXpsQjGSeYU5ine4fv7utFBnITCWQL7uzonuGpbJ+nP5MrewjL29I7aWgvy
qJJN0ywijKwRlI/sfuaUiy7KFtfvL1I2XHRIiqBAaCzSKtpnZiSQQDL2hqz47WTPAZKxBHfbcrMX
EXzhqG7nHNZHW/oCk3NlvvT2wHiEkDxBkk06uwGLLD+me8JOhKdOeyQbEztGp7U0gPH8Fw3vkLYv
/SPRbxv3Do4vB/kz5LGojVa/aYKn6Qrb8qFmd1PPEYyqrmoPoX1qMJQEjTtR1HQQwwOfnUciVhdG
QBseteRSI0WWVUfZbn1gbe3Z4BKjBTXRcSOALlE2Rn9y4V4Dvoe9K/xJPYDtd1dO9OCKygOPcYh6
AbQ+fyeKJNoSYMBboPvXsg4j8ZFTAmJr6I7cHobfLm1SwOXNgiaEcLp5rJt6IHpNCS9aYNzxn+zS
olI05t4DHuVchAFP8Yu91e8LbNZDmz5bBy8gszkkOP+nUCzdIkuQ8a5eRUgZB5RuH38baaniDvHN
S3OKdLihgM4TSiJutKeksxYMBg/j504Exd64VBksv+hghpTO4bi/Umd7vEgyaQ/LKnmwDMvsgubl
0J0+Qk97w+5vweZlunxaKGucCCQHsLBSYkhv5bnjN0Po2OTKn0Zsh19Pk1uOvQiq9zgat53LE/Hj
26y+WUxJhuhfUuN6Pr4qbi/s9xa8UONi4gscWDVCPxIANMlAUh5X4Fp/8tsp1B88dClOy6ooPD1C
4w4XLuwizZIsvJp4ed5ERPMzlOJszRgtKGPohQTHE/AUR4rEigroOMgQcPxWHR7bC2ZYz4xg4kUm
pKqb2RIgONLWhtXaR76VmkDhIdQSjvBuQvo2xTSt4Yti9dmibet5r6jxGrib34ztYMfc6v7kDrva
UMNta5USa/fUhG7mfwM+er6LmGuwGDs7U/AlRAI5J/0ZNGzy1yp2b44FcMbTjL/9LjNiIFU/mYCz
NQCp7a2ip/9DnZqBPDbGNhoCBPb7qH8TluOIMmdH61hp6c7+HV844fnfWZNh8wiy+lPZFhg1P0fk
y415OJtOyU4DyIm1ep4E3BEm+jAf59vWlWMKuVO4IDqvDKAHpHBsWmUU2M4IVgMhSKkF2rY/56HD
+mi9mwuksleu9G8VdP/64z4YDjnj+3/DpVDgYQbKO+vwbk0nyuycgodGlix3yDBT5Dz4vOo/K85Y
Ly/JjwbLCPQVv81iMsmXiaS2ZHO0IgpVBPFbZklGjgyTnRUwqvhdaX9aaJkIW4FvvuVT0TV5K+K8
y6TwwZGTMGbfwoE0jzckrTtnwZsadkyIFIVgRQ6+ohEvCoj4nvQRmgOrIBXsHTJFd0qmHBT/bQva
zrDtRLbZmuKam7krHHGTrNJopn9GQQgx+aONus53p5b2RIYw68eHoNi0eC5Tub330NwgLQIVIJXX
WN1ov4VuCqxFwqRaWJ/jpqMHxREBRsMN/NogU3V73Yxt/I6J/kNo6BdXCbo1lZwPUln4PTlWCm20
umDUiAdW0407j4mBUfNcEEeqjd2b2zPQ6PAOPPhiPW5JDxRZ/2VDUrU1LDOzyCgdktFp6dDya3xS
XMX7ACoI4cS02MYhmr7blxkl8+G/bSyTe8+YibsVFJLapJghZd6+0cew3N8zm3oe2rCP1LAXT3G1
6r2s8j/7j4U90JktLxeCIZs2yKBgKigFlLwYtZl8pqvJGGqJQxr4ONfPpLXevG2/OUHs2PVmfy0W
zI97gSgQI7dO1SnFzTa5a40e6AcCMBkKlTXsLRP8l6pjKVfonhNtsDJc4eSyGXCT91Ah/CU78iz4
oyzaudDjpBaQNQtTVDMh/smwKla0BQzhb1rAtOuF5DlVmZmw6H3V32zSnVSgGrH7HUc/Pjsticwb
t8z8w5CFa9dZoMUlkmXwIoRDLzLNTGhj/PSsbABj6kW8nkE/E8pvW4Fjs0yCYDEd3Of8UZuXlJ9Y
TsaMNTZHD+RgwX5APi8rj0BXADG6/NWSiQimzwl0P2vH4Jxe5BCKPaEy1UQ4N5sui3V2dD4xA2Fe
VCazlkTTmmY0JVcq4+moIuNSGpVY6orovnKGYTvdH6QGJczWicRtiHV06y1684pTc3Yh9u91kdpj
krcwB7bDjIW6ZpdZDaNyfDMn8DPZIwE9lYw9mgYhmGsZzeODr71AUFVpanpCkSze3p64YGPiln52
y0gtWfU1AU1p8BFXzvLZ0IUa8oDqnp2X3YfnjSVgP4sxSqiIH4+y04YM3aoEPXYgdZOt0cKSp7Ha
cyXTiSIIb/Rf842S4F4E0PsEsEsuBoAUTTC6Mnyiw5RBDKFOzsBPllAkhNdKCU485LjS9sVobdMl
cbee76KNp0aN2tooVmgltv2ygKssEgVQm9trsLq+cUvABMRtrX4wZatd1UAA9pAgmlc7hsXPYWGg
Gb2/UR5f7mYXQR0dVC6d85RYIhVGUMLsBD/RzDqsN6LLX5/XZP3b8gHkZa3PG3gsKLKGz49N4yVb
mM3w/1tQpVKDJXvy5x70HZlU2nQjrL53rqbklqU77OYKhSBabA73M1SHKs0Ecclrl2eSW8u8VUaX
9EFkCriTDBOGF5CHfv9QU6IgV53chRbgbunlUWsriTyHPJ99PZESBiG2DFk+3JTndisA3Hp90MzD
VKfRPygp1B0fZI7gy9EuSfA1RtWpfhGu0ezPsHwlZbSNpJk2KT+DZK/xFb151mYk7bk3kOzMqWfp
n25WYUBTmJDU4ZPAWAldjLi5+w5iNq7CamF/rKCT5zjX1TUa4hs3+9BdeeAS1ooiMV0ZHwyx/74P
lOV4FBNQX9kB1IQgwLqvEU7LD8jE73rXu7xt+EqlQ1sKP6Z+4Iqn0WEXp3esDNyWspwZgKgz9N4I
aOeNeUcQ+4/dnGTTlOJ1vArXscw03cRhQ6+ArhtLGuMTTLhUnFSmIx9NrMHi1cWjI+NpxeNl2hWF
LDXFAhQ2JDg/osap7duEa2zECzD/p9a6u5xWkhJm2jLxI3HRg0n+Db/mv1mLSlSu+42hXTYALKvn
CYPK6YDZ6LeIVfmrMHiuLHZAPMkYmxYmun+fdcT4JKW8C8aGegrLwGuwNpirh9SzSpKsB+AN0FB8
HEWgpDVAYf8+j3HlqXq2gHDqGQ2qHE1G3KPmO2uxocwH63tFL8wJMJGOcFFmG7vThuLfgbtT+MKt
2dU22qhXedbMR/EEzrn4E94FlQpGTkdm68X3zj3XlB7DTdH4uzrZtC5s0cb+byqTnUZniQ8T5sde
5hos32Jc+f2YPxMrWgGdTi4f8NdwlqUeu26eW911vpi2fTSM2AOce6My3j0vzQDyeHm26w3BqKpy
RXaMV1WssvHo3q4V7irHbU7U3ozZ2iAlOgOzoQZGBek0/g/Ptf/s0deQJ16K+rur4Q6/nH9HK713
lgpeWjxj0M1HaCxwieriO4oX09PvcQoMnx6Ifx2XRu/23hlh+EASty+tcMXofARmuW5h4DJjiwKB
SiQXnS9VqbaVmJ8Ak9Q+/dpOlliOrtP4CayS9Hj0EZv6zfyO7GC1POx46QWqgPtCA7L26Z0rqJ6f
a2M8ofg2my0kb+LqTaGjRA4vaBEpkgYhfma2JqmTrxZsSyhYPxccitvmbeFoMt0SAT7jzpENDk5W
0vcIBi+iQvwHPAiegoLR+zToqUDjafSNM2h0ZGo5YyaLuMUCelWEM31c60SskXlZZCeo/0badLFc
78vf3E/DDQOP/iz8kcE2bNW3Ku7SsxaDF1lMAf4XqOXZbweH64bC6us1yGd3iaTt+Shdu6PGAsVs
Nns92nbgrvfKKJQ0K2mBe4YBBYbOrLzrLi7rnKNt2ufEXDxrOmHxS0Mt/VwJSE75x6AC1X5X0w2g
tADbuaVClNbPGI+QnT6XbtVYuN/6hMLg3mXBiHTjyOc/neL19s2ZZMQu8gPsvanc93/VBR9etMoS
Xhxs3QLMeKl66ozBENI1QcYhGbMCL8sHLB+7cm475Wu+KMvR3gP8SqqeUmWf5J4/jUAjY9F/ozVV
FHPYz0+KDnjFpE3t4xSAtVOHYTxk09qxjVOU2wC2uY6lJxWFoXpX2Wsi76dEE0v2+52yNtJU4OGL
yS7jOVmf5CE3p+zD5UoZy3obe//NGIhT+dpi4fQTqHjBUEUbAeDWzxkPpOv1S2L6jGTW1y8jZANx
Z6IFWAermzQ4RiNC+FThui8Ex9BFuzh1NPufWpNg0vfH1tIaNLXys85wuUkpkbpQmSfiHYKdW6uX
KprStWbBZuo+cT7bz0uZb4+K9kyYou+LzX5Mg+/HHLwA1ah9M0oL3iTa4XqlFf86DHrlHcqkaH6P
sE1QTbZkue/m+K8YCVbVysBKiJUvFKeUYmhDUMeouVjdXurMR3X/u501ifWtuDp0PpRvdO9b9Fww
h16BOK8zVt34az14aaiam2iTMmXjyIiMgRNjEK6u0CmmA6jjqIhwarCkMTzlFLUjweIslvmi2reN
DyYZKXfjFolaARxU5WoV+ijvCLGkpE1sOiLqDF4TX24dAFgI3LCHSdZUUASsbL/1E4MZ5YMyP7p5
ARDMnU8VvdbYTL40cw5PZrYKq/gE61UO27l23G+m2sMD9XaWl7E4GOMdIgtn782MYmoY88FYNZOW
2FX3puP+TLr6s6umPwAbBuMcndlwzaPBuMSj41u+prd8Cew20PgO0bpYSZxeBQiko2juA5/B512k
neh4cKPasouEF+qpFOSGmcgZRr5QU1Wnr1ku7mopFsn1gzVCiwnQQ/L5m6XMStuedPVQK2Mwreqy
EdbucHksbiTADsKw7NQN4b4MYfmJw67V2XuC7QBqaRzTXApcSvCHZNhfRccmnxMcrrblZZBwHtMw
cnAPjZvVk3ECkId3u2hz1OhTdwMX/cTn+ZDaix8CrBQKIMVlQXnOLcOfa90N2bz9bWDvD7UI5/Fq
4uq30Le8vKTxxQQmNRAms/Fm/9u5HK5Tx8wkjEamApD1WK4HKr0o4WECuyRvzkgZeeXhTKVBTtTa
FXpbCn/DWynHgGzgnG/8q9nDpAnempdSBljg0Pa2B5E1PQvuDRjWlJ7FhYAFy7xhSy2fWQoXdSwS
rsRA1Rj/WsSfOOr4sisj03DbyZ9AdRTV+KZs++R1P+3YXV0U5EDQzye/GkF95Jo/F6oXQwA0RpK0
97xEXutd85+GcJebBe9dr/cyr80juIyhtHyY1fUSGXfOgHZyJswsWiHbOWaOMPK/q/dZnVkbIuW3
8vZQ9SjkmPK4fQ1SD9Wt9SyNekr6WYSKTmuYEE5seKOlR3Q4MtKHVR/j9EihyIVn1Zs9er34dw3c
O8hzF8us7p6P6/qnKXX05ivhDlMX9yWRTmaDTJS7CmHJAQx/BwBSXdNyjVquYCTPsXuu1YUHSPkP
dmd1CkwQpK1lMAvlGFq1foutxrXPwVkRJqktbutgiUZANjeil3W4bw4moeum8vyIFciVDsgRaJk4
TUgLsw3o4IZq2zPJFZLJ8zbiYXwWsgdlxbxCvbYJXZ4b2SmH3V3eAqC6VJ2+iTLF+ZMnNakfzuCW
+fQx8N4dG4/kLK05BRaQ/RYp2abVR4YqQMxGmPTpUgiVDPKp6LWdZJn8zEzcVUUUBePFzRI1YQo8
4XjJ0MqlBcjI7TL4XTBQVKVNs+SM22FIHSrgVK04y0dX1UUh9NkIyRmc45H5K48fkiV8xntmdm/u
KIZgZU491pOr7Sp1YORWicA25Ez90N7ovL62LBWqxwmJeBt8i3XybARD8y3bVxsnCzItXaZuIg9w
jUZgx9g+FzFiZNDPiBmP+QariUbuGNT9I0n0zmrZpeHUBVrpz1seuAg/e0W4deqa5DL16/nyiFct
pWKJkXmV/F5r2at4J0/mT0h9IwZzmaMDKetTFa0Z8CRu6QR+0eK/dhDObMnMDc4VG8XRmxPw/gzi
IGhVh3dWNjFtB3FcMixhlthjbxEpDJe3kxlF1V6vp+UqmZXbT8D7uOYxw9GZPwOq7hF+Axquw9FC
Et5dAv7/xTqKxXYn3660/pFmtC/9KgZ3SVE+PHkpwzDCRPYkh3KKimxHK9qFJ/SuaNMObxnbEoBU
cGfuWCtMCIa5CGmpTTNvWKLzjBUKziFpc6gSSEQdrmvpQ0/3wVicIlmRJgA8umxOm289kRgaJqsM
xbj9LIU5xPY5h1Dpzp7NvNPeXHdDCR+xoTujUwrNloyfBjAjdb83ZewJM8VL+KgOefy2WHuomTPU
HdhAz+qHUdvgk3pQw96FP306T6PAEOolXxfPIe4j4N2bmd3HzTG/7+Bq23OHOL5KsTCb4R5QMEwW
wz5iuWrihxWOAE+B6ZzRmT3LeFw/fqxs6TpMpR0YAH9+/572Rp70Su2l8p4WHWADsdiXYCJVJlHe
xXCBngBPdVzsDJA8rqVgor/GPIWeyqLHHqYyzmw0WCS+pPdr7NwS16m0NyIRr3RCoGmgPNCJfjSo
EJMdQSdA7C3BGVJ/kqI2H4KiN1cBRQvlQmww/Ztm4okp2fuhUlK4dBkFNmwCLK0tE8sK7PKRI7Xh
6FiDWoJKjJJVGuD/RGfx527+foNiYcKyAG0JEZIXZmPGbCRDAAmeV5Lmf21+sEnYFncUb4t+4RCA
1J2wzitCzLP9ODAt0Chg62niWysVL6aiEQz2kVKeYsaRY/jFTEBe07oty5jb/ep2iBt+kMw6QZmT
E9QJVNO/XjTUbiNGcDzLlXUOguWkO2K8dZleOQ8s68PYTd/U+nzyhJ5MQt1l8ipHT0FlGMUFgpWH
80a642CLG94I4MewA0xsdxBNwoLx0efbDZfnxk3/eDYBnG37lMLzOxgviPT5Tz1ab+2BM4UGgLRB
toh6SuCKJnTim19o4UPbrvWDzPpZubVYCaSQUq8aGFjLcaSmwXolCV3H+lEIWUzBgFhzJyFzeK8u
TyXWL3kw0Sks5/a4SaC5TGlKVCBtd3D0BbeF/zzE0iegCipk4FwMOy8r1q6mdaqx5l7yo325LqYi
HVbUbmnsyRCRegZBpvahtnsBy2r4eHxWNIbUDGtCNUpBZFhtwmzPPFu4jAcHXhpaErL0Z0p7aVKJ
9hx35D7ws8WRivPcV1/m8MN/savcYCN55T782mXB9dbcp7eUn9/ljpS8ka+H6EFes5qzXaXP6Z9y
/crl1crIbZlc2vhXunMJ4GNDdaXzq9FbMA9gu3eyQAkuRy4qxj/8J5+j3pbm58NWBZhZHSQ0sgSU
qGHG3Y1+WG6NIeNZGXPV4+VfEHpOojvh3eCdy9OdnbWkxg4Gm2MmR00g1pwWT6pinAcH2a7DsHcr
uJgWw5A+SJpNhLsoCgswrAL48kG9F9E+N9RjnBdbmE5ZOzKf7Noi0NSRPf2UXDF8pyldwt2O7UU2
TW9fphMrzz6PsKVhQjw0f7Cp1LW9MFys9tacWPl0YFaey3abaTYgNy3p2adzwlSDoLMGtcoNnRsk
JLEjL/BlwNfCViKVTKd2p8nNOvXvfArM8jVsGgZdNLkCL39JGkZ2UNn2No5P1QL409zkxxBJCBKB
jzQPGEiof2R+yWoWVi02EdLcKKVirvc5O0HFmD6vwsjLplBSfL7jzOzhl9ZiCEVwz1wIpu9bFB1v
b17f+IKr8vbuRRQ1tZOzMLu+UuoGrsVCxS2pRhVN4Zo5KiONwMGLUZNHAf6L3ihky6ud9bw+xFua
QNH1Y2pn/Imz7Z1s3V2gDMjn4lZ4Kvge7Th3f7Mq82wt7/C614n6KJk7LyUxcOoMN/BuBLT/n650
Q/7N+iO/QSXlIIctBS0ge8OpE5DQh0BFbDsN0H2yXAH6zbV3pSpArVou/pGWHX0NQGCaMVHOAS+a
MoEe9eQyC/VwzSI/5Ucvp//Ww4aCitKu+PuToN823RDGq+lnmzgQh7Rn3uk5kvraRay5jeKWjj62
sl4YsFxBahhdbrjtefsB/WxxqG4YRWwKDyxX34rOSJ37NcYqzaXeFTi2iKNClMzscSs/hJEV0Uhi
UbIrFsAajaCKnYuORx3jw/9rgYo8dy6u1TsGWopPWvBpYn906cBx+vw/zts9Hb8ijq7qMGrPF/Y9
87yvZBqCc5KucLKreDRSwVut+LzOgCGoqGw5GBz/th5nCMPgdlVndWYqcuEJAahX/tSJA+6mAdk2
LCcdkJRba9xl6VrHZwsxR/tBn1EsYmEKzGkrHQpTQsiVN707f7oIITVwp65Kga4uPNeW7ekn1vQx
6EUI4tpY4YAIT3Ueg7KgHoyslPqtbWUIhiEHJGGwhW6N1XjAGXOcTM1EN48yv5FHLvWGe4MSadDv
HhTKFv3ZcU3qlWRFbz3Ya18tknuh/awcDffecPyunteZzAhSgqNwEAiR+jMnCvV1btAdcEap8vTZ
r+aB9fhGrV6ann5CvgbcoLlVDTjTa3AmKKTWqGUuGGjLulyVRNeVZXLmpmD3vKPdCxse8bOlqctn
qAgYC0ebTQVn430XZ8eO/BLdxl7sfL0e11jvrqdFQvq36foX6xTm0dkMiS6yqQop5Ibr2y2Y98H0
1o2yZzcjjRc5Ss5kq10ae4uQv/SddLw+Um98i+PzOyMS1CDpzIvydhquWb5cA0BbnBhJoINbuwXj
Va9B+2aBIBt7E6G3jcNx4jBOsxQycCmUt4j3t/tcTSgJraqEycYayZBjQFcBCpH4IHzCYEZvc2si
oHfW+kBTprXYMKmEBx0Y1RXdGsAfuaP4elTKB8JYfzN8uEPe2CP095Dw24YYylOs8rubo7ZroHBF
Cm1D9FdOn/pS9XlsNtfWUivL1rYi9FNeOum4mJAvV17xNrv3vb1wmKM+0dPqDjFSMSOvDtVhbl0o
KyKPk3OnUV8AuF1GOGSILlupw+qYoKyXdL0qLEwMpzoTPlW3J/HuIyuL554JYylttvWIvNO8Zpks
4rB3fokU6g6Bu00LuiVWyl0ilmHysR/EwpVCzsQIeVCRQxR/cnhcDn/kzBMkvdUnr+hj2OPjSlhH
VF7ok8Dgwb96fF/wahZEr2d+N6BPZ1+EKF6htdXD7SrOaYtcTSgp8hHgOHySQ7CB6rSHiap0Yngg
hcFS0dHWGAkvznUDubw2xA8Trxria100R0TiKBVlomjVYXCXnrwWwGcH6PuymuZhYdceSfhEZupe
gLd2mnZ0+H9kJKMJ7CvmJOLr9ddVri4z1MBvaWLzqRVXrj7wgy4dp39ZD8id6B5SMXlbeeXx7C/S
QdXocryJv81TLNGBqPVXK6duvGnAfHpDETkCcIYK0l7cgoKnaHwLyQkqtvRlKl+W+3yQWlAg5JIZ
7VAxVRI3sLIJAsENu13uzcOvMTXxv01fkNAdu9gpzBLozsrjYWL5Fhln2lzwI617aaKGuF1jmoTx
6o5JgSa9OUUmyRY8OdjA+hDWa3aWET6MtDO+F4sC2zJTxr3aJ1mJtrY0DVBjYAH/2GZn/zy5+LGC
TvaLQsIUq4jtbgP8CTD6Dek0wIICbzBp96d+HvR6a9hL6BYLq4mLxduiYpezOaJMZxJJy4PaKQHs
V3TIbsLucEx4vGaZYDM4lY9VIXiU3cE6hTGiibkxFR/u9/7pBF98C6i2oN2rUIF89IxQnQnJE0Bb
llECCKE07rN6pxoOD8ibzXdUn3yhwnDMKOBADvsdws9LQsidTbUR7lu7/OnSu7jmd0yV360bJqLn
ad2MK7lbE1Fe39x4syzr9K/JdL7CGQpI+mSFg3xq+lY8hhT7Vy875vNpBcQeNsT2sMWpjM+1K0ff
k3XE/GAi9DEpMphpb4Tej0EKDDYTQ8A2UalmaVsZVGkfzktK5zH7164CesXQFgtGcQHhv974zM0p
gTjJpGtR4SZlqYM0Dxb9RrbcA97uw42SJYlzphJ4tIL+5j9ZOYteAXPTiYWaV+rSAS5nhkNc28ne
uPy4NE2f6BwQJ1hxas+ZRkccF5e8Ole+OhsaiLYLIaPn6khzCzjHJ8fWXYEO++MUmS+QYd+YCsRS
/8APsXmyjRHiXc1LxBBlho+TlGrv77Srwc1/7tZmsb3tqYX2w4sawshEib7HKqsHqlOv8gJ0Xi1i
AVenwuzQ/ZI9DnjdwVaQI47Z7Argp2sob9c8H+Jcj0NsS9cGoP/z61g2l8Rn/Ylp7hPoKEvk8A1f
T4yQ5XB+sm+KhhL4gpYmDK5a+NuLtsWB03RNVMHpbWfjZw/qPBQ66Qms6M0VF7MeQ53hSUBYLeFr
OHmM253IXNYmmfLo074QvGHCR9Rnt8Pv/40hB6yUPLB/q1dCQj+PihpVCsey3gFtMmj2CMDqCgEt
PYt2Y1xSyx+A3QdhbmNoA6A/fHSInqf6SqTw/65L9AaO3arstiYMX/+Icg05rcf/jS6PAW7WqeZn
OehQrYgSdVVfqpnKJlTjAQ4MR24972YrM1rKkqpxnMRBHwX3wk+MEtk/QiJlrCE8SVT2KZWPUB7c
pde4tMfN1RbMMJSiXCt2sVnej4de+1noROVYxeSKvrk5GVIHzEg/K5xVJA2NagUTDJ66edd25B3z
VfDX2nbs6gwAPEPJOKVOKl2O/7SI7KzcDR7a1ikxERPpldL/bQYRUsD9TVOXtzM57HIgVwqwXvb6
mWLoX9YzknQKglHOP+snL6WvVukkGZt0NtCjd0ZzzE5qrxmVuIbI372PUBX+kKlL3dMOS98xiM/O
42KLehO8JvQGFuHsCvJWe6+2o0130lhKDxlOdN/9SoyCDiMfVbRUeEhD3inoW2l58Dl34TX60E5m
oT2/iqgTWmTH+DlS7Zf9x1zcMjfxD2zw71dlt3wPvvoWza+iYtygyWeRIuGpI6BU0hr7UnTq82cf
Xpqr0KvY9JMR6oivHsITo0aUMY52dILNoreHomzjgj97z+dNnSQuQm+uypytvt98Ypwv2fBhLpmi
aoMUmOFWnMM7d9u0ShK4O7JAo85XkBxhjJUbzsGh/Ml1UZzg2uiPTJi+Zlk6mZb8rXTY+xtJFR6o
8qfsI3KjsXe3V2D1SgAKN6Zb/TfhprYPCOqlPzrDhdWiKXx8E/e4xpkAmzRk8aGbRlQD507Rkf5i
LgQ336a+65TaXkC1VQbUbGeoDRX4fUA8dqKuB9PFZ/L8fID2rh33SVVbFTHHWl5SDS0lkDK3GzNw
1BFdKcGrjlw8PcCULcbou33tCA5tSWYWqiv47P7ViENV0LCh4V2uw7Vqf1bCwa3SVaBMjXeGcqua
uLiwawIQ7F76kBXjMC89XZaG3c/uaGhzk+f5nRPlqZQ53XP3dPONegq92NAgYvKR2snOQqvPDVnd
MPTv9TLOGRw580XywVgZnoqi9w0hjtRiX5VllVmkNt3Z62Sw1lZdrZM6lCC6ODeXDlDJ9h0bnSJC
IXvqxLdSRNwPxILlMyZXFDl9iSzHW3ZeDUE/TKHpNT/Si4wzauJkzQdcqg/byCNkuz9gCa87EXlc
9+SgpVIq8owTcBEzdr+3ce9AXxpX8p+7c2HPR6NH7As5wRsvFT5KpdFX9OHlwJNYzi8SEtJjknOl
UkRof6fuoBPDpTUcg1Imgt06ZbDl4Jvw2/Saett0uimpHUVIfx0pB9QPJ6ERdKi5Jk2ERulfiIPh
mr4gKWyenSwnWugYLa+/UFoo7yoE1AtzGPdntksdvW8HrLJv5lp7MC5s0fseTKTiRClCfUQV7DDG
78ODFG50SVzy1FvoU4jyzLRoo9hKqXkEzwU1lzqznfJGkM2DjLOzfQbBKym/8F7V4UtRlBLCo/r/
npfmi5JKPvBaykB78scV0s3JMk1Qv6nSNH7ws+eGyvTLmLUKYatyIXqFrE3R8L1pGDbQ2IdbESr/
vKV0sgzDO4a2TZBKQn+uF+O/vjyuloF3uNOqmTJubgpGlhqoor2xHWiAQlMNDWY0l9SXmax5hFt9
l+vn6FaWJPxlXCoFD0lDeQ6t2l9yQ8OR0DO4SVYCabkAEnlTExCGgFyvvih4mI7fDBmy9cDWlAP2
93/DiqGA8Te7MOjsIsbwYeuFLYPsqnhdkZFkERpMVLftYdPIx9bWzFvHdDVYdmCOSyrjNDTZbdqV
JrjyR85r2AvjPHYglaydHGeLj4RvXLxF/y7CA8Uk4+k+InLsKyl83FqNki02c+rAENBHMFuV48P3
oNrWS1OyowE2l2f1QyAVlwWqndB6ymI9Q60TnvSfeQviinARjKnnPq7KGkufh1occlpdnmLJaH6p
NHSsYQvb6kIIUHQ0ELOqGrh42tH+RdZlSGkjhZ8PckjHNMpVcv1IZiari3j8WlUqdGoA9bikOeFh
WyKeZ7T+p5RZoGW4+8RF4MtpupXnIbHjNF4IuYI5Z0iN9DG4havwxbQMeH3LwI6W5Hq3eIx9OxAj
9ow4AbSk841zWEd8ckBzRoF5n3FwFQbkEoM6KjPphkMuW6JvQ9uuZ42B+2h1u/O4fHcAXGsvbL5C
S2CFz5MKDzlc7+SwO+mfmhCsOLs8WEUWvH2zywpTYHlExDfHwpc6gMuOi3NzyedLgGcGgP3Zu454
pAUDFfhQQcIlLsv3aplpYpX6NGxy17mw3thS2MTcMxCAP7VPehSdoov4eYme1kTqiCFBsuqU9qx+
2wLg+uz8IJdfamhZ0CERB594xnfXXm/RRlxGZnMBKzlb08BfZudUQa7QWhAXPhYy5klQlJbneAa0
AYlANBsa9UrD/b8qNgh3Sljo9yUUU27If0mTNvDb1eWGwES+XouJXf9XAhcndNu2AD57gjcoCHzk
EnTMnGV4GhLtEWvvZyHe4azbhUGhCnWkqHlwds0uzo+vNIJ3bej3zAjPDCU7jaDEZCgCZzCdLdTR
UGmMa6kaT/F5V8iQFySF4U8ofpXU6+njLbBvtZCDHDxooL6aV5jnPdSwJ285ohJ4EEwnWurillfI
5FZ7puc6zfhNSTDRwOXhFt67dxqo3SyQKbMbh+edfhqKyYq3+btoRsVS7NpoTC5uoRXyN74lDAz+
xR2WpIUS2qFOIO2LiEg7ntGz1AVzLxRl91fsgjI7RwHBLMcH4iofKTNBw4tIcxJxyL5eZR7146a7
WoQNAoyJ7cyRRjjvu2ijydN7ifou6iteDmiGnITL3BMuDnhf3hiJ7lrVQQ7BBMbSAJjs52g00HF3
tDrFxs7+P6krFwB85CSqcXjlu9l8/OYYSzuomRS3/rmV39V7c7BDBBOUS93f8eNVrCAB9pJ3kQPm
HGtcb66TpalUoO3YfL08PvXNHGusklXO9Ylmn93A0+T9v23w5z8tsBJyCJJPprIbXa7o4NAmtUZY
AE46PlG/P2dML2IJ14ZYmOsKkoAzrQUi4SjLU3N5n5qMS4o3pbjSURPwV6eSvgYieJjoBb3HonBl
QqMxgEJvyJ0q08lqLjUDli14CdCNZSDVrFkUI49WAQmStj1xo7RxeFr9pxHuFYILNdoMBsk7o0Vu
SkDeBSPaJTdsmeT73zMOhK58vCGiw6KrhLE1VzcE6mhhWFz5TiGw+RG31F99eSLyrPtHA0aiuX2C
5+aEIWKUHh6IlUPtk/IkGQG76h7388lqfroghwSOhg7IcNkfTzX6inuELnO7lxMY7ysa0kYpJpxs
dz13C8D/HScfSEC8CC58LWO82KWP6rOe1l3VfUstPhhTzSPKGp2vEDIUQTjokOjAJ9gdZT9FKMlb
gZjuW3xdCnoHRQwABW4r2rwznHrAp0VHPVd6VLc9V9O9ZHAbb8r77JbTTR/9gAhEUcXSvmoyI+VD
UTEiw85wG1Z4khnUKsjOGDCQaWVizBIfTNMIKKcznl6VV8hqPG5TzrLAcuafSt+4zcEZD/EmFkkv
7Y/A+IQsmn1TFSAGjOO+9WFkSeoMcWP2zI6YeeyK9z5X9uBcp5q9wwoYKLw0VPLOHzP6iT/X/udM
hnXnLzVUD94ZZJp5qgjVNOmWCr58dUxjKVFcMkAOhTJ6U2rIfi2583eQId9hC/3Pu6v1OMahTuPz
7s2KhQLZH01Eumg/i28z/EIoIpm3l0kFPvh1ZHyGQkLMwAvYpY9fOcyESCqumZIsp29mPCy4ai2P
UChxSOIpq0KSCoF4+U6RZgyPyZKWm2j28LuBZHyHnGa9awJhA0I/5VM3sf+SXk/rCXqItK1Emwhy
6w/z9HYPV1U1A4vgUc7tPPRF55gK6kvvOW0WABPzT0PCnNm+WSpnGd+q1P42Cz0x1jNO9BxrG1O1
JJgedLAjiP/X9WlqWUu7AFhgRUlK8kylFefYbjIG8QC/G8c38InBr7xYdG6MO6iFRb54UWe+vhjY
XH/0IgIQsUz8s2sIL1ME7BiTaqQ7vtJ7f80qU1VWCPnA+Mpwok/Wibu6p3VzGiB1jrz9xbATRaOO
SCggrlVSnIx81v+5ydSqf0KZGBpErS27cEiNkO0KDthkFiCn8yPf6SAf41KWOUzpHLth9e9HAXlL
1qbaj9viRr/c1UbpaRc9b4KVe5sXD/y7I4eKqVPC3O9cy3yVM3VeUkzK/HFrMXmws10xoJ6uoKOs
G/tsfkq/k1vW7WbKzLrPRqY+/tBMUMS0ofeSAi3M4ysdSo2TD8oW300wBj/jB+7h1ONF1T7MXzQ7
Jf/dQpWNGmgPMb8B1PjQaemB3HIyWJvC1h1O1twBgp6WDj0gqIQGuahr7ODzzVEgbDh7eTv4lZ/p
p6Yq+qQu6oGr2+0tDAXjUan9Z+kdffurgZARxGfM8suiHypjbwXJ/K/bqsbEixMUVxchuYlSM9lM
1jqUoe/sKlW2mk/g3xeEdYFoMgqj/zMWZaSBqxjvAqgB3NDbNwIvOx88eWRByJNW/rvcAqzIr2cw
5j/d7ztePxuy8YUI9OdXYTEzog/CP1iRyqSqcEBQ/y+bbBS4CGXfwydbXFtuS4KU9AHHqPHEVgdn
969y0eoVXeaoXrfT1b7v/PRk/EsZ+MgxQW/9XL0b/c+lGw1mCmqLt12IUqiTfr+ODeIWYYYFXFah
NYKeocvuZR5K0ASp2B3aZE++ShDYlSWfHSaLNwMZ9PurNneUC0iR/zMZw8T5fzoYGXLyUtt5C8Jo
pWZKEzBhNUtyetXJ6bvNypeM1f46Msz9WAeXo92ApC3g6LQ1pGnopkE8tEBvRnSoZLBqHytg5FfX
7ZUSYreARhyYiqbuTPyAMUHhlZESGIAq/2nVcka8BLWT6OYviHXWRn1sqaU7c062oMKcPP5pJ+sm
wBkC5MW6ZpKQazPy2sadLD5+wa2effCFs3jagYSlEc0E5jaAtbwIaakYTbfrlwqx3w0743tCsOqx
H++SDnyJmH2S0sNdCFLKknohOaQ89c4pudxckGaZKZBXHCcFIevPwBMduZLb2T6byrVFnfgKK91Y
pMw1mtYECQV9S2yqaSAerNbuS9hAFJILkYKfYhIQuEziS/cHs+fZ/t7zOfKVQNo8YaP2rWrK7gl3
8FRTRqi16VW17W/tF9zCNRzSairNWw8YtyLL7vABuwovq0uSUEE09hkmJ+BPEgJhNuT6dVg0f8Gg
5HyBqcv1LRKYlwdFanl2iSntaIMt6tieehcaifd3yibfrhBbfEaJUMV1Wvg6FVEeWynRU1yNI33Q
dN68VYd3eg4N0124dFOfF4fRU7AjbRr/BTJxc2f1U/GKFT5ljKudqsz9fRbKCi6zADYMew1nSn+D
Xzfvfqxl32gy0k3y/kzKMGwCCL5Aq625TUsdYFcdfkV0d+3067UJX7wTIxJclTiQcxFBJM0YdkhD
aAjv5v78IYj6Dec7DmFGjjdjLew+5/8Eu/71S156ZGnTGZViVAbyG4nsPEtNx5mu6n4MB+srages
gDysuXUwQF1hfTHHkSECgM/NlETsn7az+ozb0l+RFl9cM8Y7Yz/j2zPqxeEQHeawTJ6rc/7iWEki
dyaklGqrKHtzcl6iS0a4TQeArZv4GVn4gA/G+SIfwG+N2MTLn1qQE4Ig/gubKxrsXO51T541T7aH
1fRlL2TPoEeVwfDELs/aFAhdKjHlwIxrn/IlC1JdYGGrkUPjkdo+Re8nE+FWxyUW+/UohNuuUku/
e25edIm1oCRXqZ6a96mhimoJlHYgNXgGfh14/YN32cjXe1kCw7UBnZkFSf+ckSaBh/xzFE2Hry0z
sDgsfrryJQUEUecE9vU7ui8L17kIikguYsd7l1dECKIcl5sYcZG30WQn4+zd99kRgZLSkA+EbsfU
fxqfC9OcifHxGZTiyX4v87LjOZ1s7JI0J/ulFNfwZ2T1unk7sQDUIi4URoxgAHGg3tgtXYgMNWEQ
Dqkt3492uOQLngH4nkjm1Evnr3z5htYC/oyKBwx4+L2rpZNQ3fNgARVd+ouX0d6z+Z8vLX7IZQMm
GFq7oLLpTkK37Q+HKAkSHN3958wjB8URbFWu8iG50bCHJI1deLNDsV0PaWm7LWlXsloEH11u6dbJ
7nSdbASQqB4MBvPLp227lFE3RozvDW0G4qWYFBkoZTvK/p5HB4trjo1OcFOuwB1ZKmpvmAxRiN5s
Uq9hTsFJ2rjpL/V2mcotdtK0elNwKbja+lsA2O2NrrDcWHtvV/UetATY+EDR8YaZUTgrpeMqJLzo
ocN6UkYaKbYEAB9yM21QI9a29cgJeMlbTX9RASEoIN2SeA2e19IfaFOwypRkqh0clcpllMM2QuY/
BtjwQcmzWCukEPD4z+jLmt15pwf+hDgDOsNHD5FSNe5nptrmVGbp5OQ39E+B8IwE5UN0R5redtd2
+seKSuXvQkfuaeyKSt3u/+SrtCTGbxIAJBPgmd04B82utirFS6pxoE0LiM5e+2NNWKJobdGbvlGr
s9F5mUi4r7t05FoaKPsRLXW6rdPFiq7DPi/lpyOM3UIEfuDyHZM3DOd5hzWHFdVIBF1WmWGlQoIl
If/fJDJC4yjqvYYZwf7VBJTAxO4/JwW0D/b61VVcW6Fhbb6lEFchEnCJg29VJP8OOoafLE/yp1z9
UOr2K9zfSDQCO4hb2s44aGE74v5WqEV+D1nQIIhPpudTzrUErUEuKNh83cAiAIdh7TUVWVZR9EEf
ot5IijDRoiWornsWKsorJ3klsHLKR2pshCtc3QKehoA7Fd5wRQTFr0T+Xq7d+FtIQaIjwImFS5t+
Fhei3nyQtLIzoAPUfIOsLNylsjjrJSfrPutHCppl7MBHM9rDVHT1w13zLmF9TwdSxMCdM7PJ0FBB
8K/ZqGCBtCChlqHWjnolmIx4+2mnWeKlnB0xLItCBQDIhgbpj2yRkmPcOnibbRvnt5+0hOc3Od9b
vGwO2S70x5tJvTpwnov6y27iBrKjaXIOI4L4YotjKsc7Jg9wNv/6wvooT9MdT5JfYzWKN2FYzvEh
Wnlz7r+RDwHHnQrKoehZf5qpSVQqcS0Sqhkbz+2ZHiw3kHF923/jT7Kp1h5q27v6oP2s4MB1tkbo
YYvrFwyTT4MDZC0bfQ/Fy4WNLQOBC+RTIWBKkWr4yCwn0XEDNJYCxlkxZUwrjFfhA/Bv8kARjlRQ
NdJ5TD5t1vzgG3MnXEdsxRQPFDuZphPkwePBePEf9rxIqX7Un6u9biqof+MMFlbpmdFOd2ysxpMD
u/wm0aHkToCCOdwy1IqLu22A4LNrk9uppCZR9bDEu4R4XYmyFYUlHSg9cg4me90pAVusJTceuTIu
6TyUt5/UxhzRUIcU8mduTlxekAHqRvM5OPtzO0HgjC5zTfErV161hr9em1ijwAiwykqbBFKOtrSm
SkVwg2cKNEgn0+mP7eMBXJ5L2CmClk54BIXlrGmafq1Pa440EV+RZ+UYsfPgH0BFu5wipDM/s/0U
Kwf2DLG+ot29ZwNuSzhl1OJTgZpb6hkPwC/AkHnG/7+5L9Udkzj2QH/+8zuzn5sx996v6c5WoOvW
TlC8ytAb8tzK2c1cVNac5pYygqmAWoMrBxrgpTkwfdtBsoGzopaYvvOwTpTcBALJ8m7BANUjpu+w
8TBi48XK4W4DQAP86k4dAEW8WvdPomADT12jWAKlNRBlJnDOe1Gt/liHF53CP+kqlWv/3BDKAF+z
YhE5bT1+Zwn/ezN1yweOAuvSWkzdReUk5IpRF2Cs3iIggr04BCWVx4i2/crTk0T3Jj4LmC7X6kz/
nbyzHa+CCbsW4x9eYnkTST7mtQJNB1Dxc4h7lzjKWKrAJnky/HxDxusTbK2GChE6khh2rqOofQK7
FU0eXiu9ITbLf7Piv8UuNMLcFtNz90teVLJ1BWEqZKO5i6r1bcdk5Ilp3a3Pnw4kaJWrJBLk7psR
EQWbA6H1bGrcTztdqDWaOaav/f7ymeBmX/p/mU+S6tILuBqPcByG3h2nmXD7mGvgdyeKk06PcZtO
sqph0i2yyHVEQAA6LI0M6eZVEp46/vsXZrW9eTUgSfEvmaJuwCdHHWxboIUW9Y9so9bvEXHSAqGb
/YqE2et9gqSlmaKMrJtsv4BCqvWhPh9nEQZOg/OIRQEwT8hsh6Zb3aXiyvboPFUMKViCkUJzuaf5
xL8LPNaP/eh4g6P+3DXKuTJQyqd0uzfrlBlZsIxBYza4W5ZYf1R51mcnrkKzenTkjTszRSdFvVkO
D5mqf9VYNukuebZr9DHwr5NNaPmvnR3hwJW39C1c80/77PfXyKunqAF1G8lu9adZgDX1Gzjeti3I
nIfYhGofoOoyfby0fSaggsafbcCOSOA7IyFYQWp2nmwlBvV4UlCAce0Rh40njX1lFcJIHSElBzQz
fS6Q3ZHeWfh3L6W9FPimsfW3DsrdmvgNRP1Bs+dPhzfmpVPPMywCicvOPZSPbJXotWySxbyroJzb
a4xbQ68m+WtM0f6DH4dsOJ1QSO6ZwtfvsMW5Qaq+2HeVp6/2pxcksBhVFjW/ueZzEs7z2SSvmtx4
xJ/dGdQGmXhwWwZqyB9x0q2HW1saF0YDB9hfBm74ti0m3YhQMpdNTXhCZIcmrvVGRnhL0U+OPiPW
yGyNL3/NmIRP9XfYuo9RwO5jW7wqlST9UX5b01ueQDPSfGUde4zM3WUx8d2f0/cq/SlaxgBkbcdM
PlO+QgeddnyygU3Tq6efNuwnNfz3zsLq/mCJHdAVMvuIBG6FW5+yBvp/gTz2Bu1n3OsmXS96h/tx
bf6JxPLGZuSCQjA7xDgcfgrnvWemZnGo7rYQmAktf4xivnQDTn2eQpKZFp3ygFTc1KCuAEspC1Aj
Y9fg9i64uupd7076fxqRB+pAdznFJ8h3VJ7S1V867skuJDx1fSmaOmaXbK65SfLQqMWRcCT9W7ny
NsZUHildBTPH+rU3ZfGZ/Goy2UL/l5EiuzAc1ekUbwv4LVc65tZlqZwaClPBk8O+EoBGtbm0kfdt
3VvB9LnZlPOmodTLevQpQUXxgtWR1+h70lSXt9gU8Jq+76tUj7iwO9J1QEHZaj/FN6mBZhMqchic
d+ITFvj7HaJ5PpRYfZoiea83lpp52bBvYIWTJ0jB5p8RuhjaeOKmAVT+KDRg742nZonMZNkBZ8CF
P9ygRQKk+zXN6HKuVphu/pPrYAx5PCboAkRXQ3vUbysI6RgB/jW7rUtyxwVKWXAyHN7sNpffR7cf
I70jo5aSgRnBAgtq9BjvZmk9/dBoie33ghXXEFOnGBDqXdB7bAWhEPxFK8PzHUTGWuj5bkcUwhIN
z5qxbmH9QQ2AAI/JTBlYPEZuERv+jTY6eza7zzIHFbPYabj6HTkjfFYi+2rCWp7MH+kvU8OucqnT
Khlw1QkM+semD1SrR1/Yoant410iLcult85FjH4JaXUtrRS0psc5TPibcdlxyisSwv5RdQmd/nYd
3zpgoazzTFJT8oSlUIAk/ujrRwjpc+HTF1HHbWQVuBww/86dR5HlVv4XDlftvcMiPgRKsvtVnV3N
nJwyjEcTc4++pvJn+H1+r1RfTmu+Bl70Rv9mQ/gu+4Xt/SNEYh0vHq/38GCQG4RDxydIKwbH3b3h
VJgNbR83Ah/mrINtGoT2yez4kk3zuFbrXyWmF9+duUy4kfAT7awZBnALa9pe5va2pB55n7XAjrcK
nNVMspvp1b4jMtMwBj4unj5YO7/TBQYDJUorbkJkbtENmy3E2SYsjYEJwOk+P9N1aTlpnK5ov4Rj
1SClnjGHnSXi0br4z9RE4dT+yAYM8743AfmA8GQZkIhSMo6RpUslFWa1MBwi6Kii5F0yMgsT6mlR
QiEDHDyZn+iwfSa+frQx51oWMAsQP/GX19JZGNs5WLekGHJB2d9DRzyHrzEnEn6YmbU2xxIp+ew1
pcRLqArldT7F3VOfXOAwxTZE2bSU4DhR+y74RWASCgBpF66NzbIzq1MZseWpN4qjfnOi18YTBt/b
uhqx/UpTW789DHluqRh5QrOLxiCrqIs+qrHou0W1X/Epd3Zi/7/5gAJmLU98fKJXKqul5/QwqW+C
Ua2TQALFKyPez8zlCu1nBc9VvHLqavl6RJ3D5Ijo1ddH9GmjmYAwrHh3rYXAG2co7FK08PGmKaH+
0VUA4umgdRYqz0cqrNdpnzd/SJyqUBLJQmsXjMudEWokDRr2wGk3uassGxKSFUWx0BnEYmfDH3aD
eQsNk2h2SlRLI/+oxCIILiQ4X24n011kjzlqIX866dqskE8IH7HDkJ/MX0x8RB7X1H/octhcDhiK
Thz7sj0COp6stLCgvtOhsXjdc9s0nBDj3XXPCuwAyPACG24UXZKbwXL1/z4lYWdS/k848monXfcf
M2/htU8O+vrs/OvHLM4DBZL7kszEjwR0p7G79jsVuo2PHCNtbwiaX7zyue+QP3nk6AN3Y0LrocwA
jCxneQYFsRvUwAljXVlOLu/HySyr9cGjyAnRTcRpGkoyezx0pI9F8dTVTXQAJoFSZr0GOVtZQAbq
aA3rpGePQkerVTjYldarC9KVXDBIS7aQy4V21JPw5xR7h9aSmh8htVFXWi39dLvsjVTrn8wbTRiR
esV1K5Kghz51f3oko16V2hcMEpIORfj00S8CP1OxI+AtEprMDkZLsGXnQddoX+P5A1hHfWwgDsT9
f46bPhN6rDF5OR3iY8Plp9rapZ+K0UxPMHqWA5RuPaXS+5PXELpONVaIHDk2kersmpm9WfwLeC/z
DnUHwgFvgm6gNZ2meyIEdgteLJ+ET961MWYkFNHin0HsKtO0WYyUL3SoLe1q0xkzJ27Hcl2qMkYK
lQrGrhV4V5TPzT6lRJRAbStrHNphLKkSk6KkcYS3ybwdVs9DzVMoCmmuoR2O+kfEj8zBCISBlub+
8bAFiX6cUARFFz2RUnaU6eCYQi7zpZd4G2+dRYT7cHjQLy31tSqAz0qcw23HBRqjR/KahpxTuMKm
S+BX3c96cL/YlPx8OiJuzsaHO84jcfzeh7VCnB/uMdSYLeXwULXjo8rJHfMsGw9GzrruOhBGGYn/
TAQmhvrMLjP9wszi6u09gqyOkQAN2u3yp9CJ44SNHvO8blxsu1Sc0Ae+KggeLxEErDNyJ+JiZOd6
NJuCnt9bK7C6djWpRWkd/kTqrYaGGkg0BjQwKXN1lHZX1v4JcU2ch72mE74Es1KT3KR0v5zgnWmP
8A44/xjMcdOS97KqIEsxbYWZJ4MYe40jHZKNp1+qOVtuUwAWyLH+EeQ3tXzpXXnt6NP8Da0jmA58
WXVibCuP1vtqn8U1ccmN6IZQ/OGzS+ylqlYHxkky1kRVodeZqZ4T72OdXh7S7lXvhEkeh6akCfsj
1fu4F7kfOBiHH5iQTw5D0LgFjlmc64ZUBFSrcNLNlAqHFqBk0QW8pG2RUwjKIb3wLMD/J3UfTpK8
eQZv8jr8rkacjyS4EsFEZ+Lk+IfDB9JhGcUGP87iKYn51WuAIrtoH7R84f32FwIjCNOmgcIPIPdd
ipfJolzXcST3vwB8dqjcNhh/FD1FCY821sVMMcqFlP9shrpA65HUB1DigySMWd+VCJPdC5N7ig/P
djNog0nucUN9EyI4/8EhOVeZmDR1U4pg+Zl6Olg33tGmphpY2ZiSoKtWN5oyflPxq9pSyyCdyH5L
HaBFkzK724j0Gc4Z1g6ysPzCTJLHmu9SMVfukhqkee8O4m6v9VXJggD+htn34HkOvkpjYXWUnREg
GsbtggJ3QBXnpDWlla5XnhzrIcCgOVfr8QGVlYW4N/K+MvR/1EmEHRdKzNMxNsLwpydSyKfLJDur
+Hu4Mk1GHsNef9NTUrRHSAt7gv1GxXhnFFHyl/3KhLbobPqrDB/rYxLaCT9BPwA2dQeRYgiUfQfW
4QzX4/9rw6enzkvQCUQzSFXOVUMDdog0Y2DfVHybzvlbqeqZ+1bMaTl4JtiGm7IbkthGruMvwDR+
ViUFU/ueBfJ2eTQFVOF5VVMD1bzoqNqhpGhwWd7+zOhVO7BtdJzfL/5zLRVIEKjjiJsKU7jtLbou
tgSYQj9Vhn7f0i2Cs/gJRhyj32h9UXYcvoSEH179dPe3A38i8T27Cj/Zj5NyA3cF7FyU+Bn5mkMt
GALz2j4/0ROVi9V+tr9qr90lVz+xR5ulWSWJ7l6cutAYCoM87RwAlJpsQQvllNUUZhsq/Ijeh+/q
2xiBFekoI5NLxbD1kv3slfOh2DBTArdp3trHHvTvfUa0LmXXjlsFTZcpq321B+9PBvPuUJCgsr5N
w+mB1mqXjzmnFkfWpGdO0KQe+d/2D3Wk9YYSIhk7K4HYETxwuSGo9Yc5pFTxHwmSEEIMNZGV6rGe
nc4ih11Zj1O5El2MxWgaNt7RgpEUCMFh9wqUyYJA3ZjOtt+PlhUybU/N3zjD/SFstxxD46rmKcgR
we3fwL3t16RefqLDrokNZ6OnxRapSOjTQkG1x3HMgJsXODraK9ZM22cxvTYObbggiaQBbUQHEBFB
r/i3KMzdYLfPeqMV1TwHlDOsyicmG0e2ir6YmjWZKbg0nPqBo55fdf0K8wXJ2Vu+cvsxen3BFFHV
kI2nu7kgVFbk7UzyTCa8do6SrOn8+psUrNTwf9fSZlOhej9SR8eCFqBnkc+xcSzjXQ/cqb0Q8xwd
d8SBMWnXONNUfcnFJWdY2TSjZWitNCl5VywQDEah+u69JNm4evj9iaSjkGuHdK++qWj9/GqqvXRB
GloYbgPNVpdxCJ+6DI3yoNgGpw5WuB4H22eDk1aZrA3ILyTOGSCirFGdaIbSV5S5tp13FiIRst5r
/ozUNQpHn+mN7SLdqby1LgdbGWf2WKBUkw2mj/80GsXTFLLrmpae/+MFws15fa0yH3AKmgPI7mCw
+zK1PxVq7XbiKkg4tWOMawAYz/SJXAX8IKz7n9tFia0JfNTpE1YGf6m16+zUYtBI9xiyY0UeKhio
9sPQUY3GPNQ+8Z9FeZAAH9BtWFlcsVyBE9d1J/e5oHplR4risInYyqvJ+G2Dw29g+hIb9jMXWytp
ULIBQD3jefM4miuInhXtNssQGpiDtob5ZjhXVw4Ino76ItQI6wAOJ2xSDYDSxPWk07GCtJYFBKC9
gSvBviaMVFphiwI9+pcXw5bZW2drI+7hQiz9TOeBwpKjNie3phyBos8i6JdwbRmqoEfvFSOLU6Hc
v20g5eesU6F20JLEx300k3qBVc7yBkGID6PbtR749O4ZQSP+WJMe4kgiu9LY3dOqGhB872+xMggk
X1R1y07+/yIZ+pdby+Umhet70rj4bJzx7KXRD2yw/x+ZmTz+VkNdyAm5eetdNrEJu74MuhEsXmED
Fq8d4f01NgZOwaCL9ohH1pBCJQm5ttRdSCSnqYaPA8N/7m3sQS4Da3VXZn+jM20rWHihH5vJZgJ+
gJC5AQ46ZNZVEErrvIQElBAi9/UAJT/u9c7le12gqEPD6Sr5q4tYgBfN+B2g5l9tHTAEXTmg+SZG
FdKluvvC1jJuEeBAENESA/IR83IVg8LuSADbNLOShvx3ESZrJnFnTsaHi20zJ0OCOPj3dzO3LS3J
K8tJHtQtVDnxmq1JA2tvD5UZMYGtWcLHns6eo5F/s/6zih1vHEFGuNYfQRMHUWi7am/U1u16G3ap
fw0mXbglvOyT8kXMWKQaNxeJmcNjveDZx5zB+wbEpIwgb2PvKUIG2OibAGL21qGf3kFNImj4qv4p
eKfOYE68iF3SrHNFABm+oPa+9M7+teNjqNtNYBDnv8eQu7gT4MDs8Hl+1wPcXT0orySSBbAUcLYJ
bBL//Pe4IJnwGUWdTu/9KQuZP9NFU+Zl+5Sls5Z0t8/NrHz9e/5CTj6gqR7/7GBCR3/bMM4SzmMy
62K4R0oLKL9nKVtkyiLQmTlekLq/PIJk7eSdijevvzxUzEOWdKWloapGmZ12vfPMR7VC05x43q+J
0GmgY+tW5QkvgdS7FvEA4n+VTrJAVSKHmi+8fNI9sHTpxHdliLpQ3NrRW3b4N0VO8chUvfrSNdx6
nQXgAd8vhSCFTq7Yb0+Y5ZPPKqGoVaw0UjuE/LuKUxOjRiZiMRoqaVRWXHQvvEWo8H06Pz7I4pGc
WW2Heo5W+iOAWy3wNcoG5DZm2cHFsKDYpF3UksFdjesxedhYbjXcBPy1g+vjAywas6KwHcOVMkU/
5B97I79aRAXf6RCCKH/uCoMZ+m1LjAkEm6MwTU4jk53hhK3VSo3LufHrYxBACJIBbS7rJFDWBAeo
8Q6eJX078C+h7wM0gxybCvwozsBpWxz+cHqUC0Di92ti7GhvDGS+YbAZCe3vshltJUjm+pFAWoO1
YKcAc2jHs1oAUWEemMztNyl5P9Ab6YqIV1oj/6CVZLpci7+uCJeuv7GZp7KoyUxuhIGYetmcstOT
ulhdhZUqecrliCw2Nnq0jKr5Awj3vOMZCU0eH19k56Er+nyZWXjpQzRPRGTR75tbZx9+plR4vaju
H0hfxxl9SM6cj79YxkNwTdWO6FSIUybeOKxaqbyP5BnCzUvgasvA4ybV0xEga6MiDhENe+xxNLDL
Y42K/26/li+G4n5m2QhRAe19j6rUOJSeLMPHhHbPYmQnAspsFxPSuqGTNH58xI6QTt6KspTViC5X
4YbXIAA/+INOQ65TkGU6uTQDpcOvdl6GbAhwm69VPQctnKpD4eeoME0fk9axPyu3ipRj1Be7agcQ
NU5uMDfNt09n0wNWXDkhUKtzEyB0w4TZQvCMTHkYpIL/Mu2Bd30WpGns0xdaP0Hrb56EClXhrCIK
siMnjb6O8INfreAvTVwoO3AKc+PPHySyfx0RJXvHb0vlEREGUD4odEWt0FEe6v4zemYSBDTZxp63
Q5BqbCylaAhq6lJmE/ZRTV0aqLb5V+bI+X8LyA8jRKlUmokUuZz+cY4TuNUNC81k0egZX3mnGOwR
CKyUQmgcWwVunhVGgfKBiVUtARSdQFAzMmKwd3mXmc24uHKk9sHITCXfWj5RK5HZe9mpe6XGZXTo
UQOS8atmWghdTOGSoc2kqFRnItsm9Tc4c7c41X5uf9hvAcohp9sYR3aakzqJh5MpAEmtJ5X0fnRm
W/j1W9YIbZlmvhkbSK0PmxXUL7PxTQhrENvSpq/JmztXCwKUemsSr/qm2ZL6n5lZHtwoISUsc0cc
oRlZnTk01K4cFMhK8Orgh9onCXrTzQjlBzNRdszjcfPricnQMs9Fu5BoyzaxfTkFrxhjtRNnBeWy
l0x7zXl2K4apxykSB63WlHWKgwNo+iBmt0Rs7gmRZYSz1rI9RNuwMrUlfZANGpczdIwCK3bETorf
bCpMthcpLhY2+QwY5goXxG/2NS+2E2HtRrkZ+Qfw/dIRWfQ4VwkS3OtZugKXCEe5viLHiDUwE4d4
PqYMbXCI6rbx5bVwmx/zihYrY7nmvEhb+a9LpjT6e6nIvmAqayJi2VkZPV4vLxEF3bFL1bVgj+zl
dV6jf9/SS5E46dnre3dTnUsQt4V0Ggy7/cGuqEdLOtAZpSDEYJemO0A8VU0u6K1g7iHWpFKqIxH+
LFAvRzwTv503K0USmXqrPC/s8QqJoJbHG56MqMCcPpVkv+qazeUIOZby6XJe8sssScezNEKomI09
R8uIWmeQ1boHn1MTtROvIjstlGf58pkKiSDJd73vmfxRB+S06Gm7gDLZRzF9/LpM+YfkhNCvpj1y
sdtsjxW9V8OoKKPu9+VF3Gps2InWz+bGCQg82EMG3j0icLYlfmno3ntvjnqvaUAyw4rpgWfCXLgM
eYiP7njxlSXUcORgVuJPEApnEgDJiFavh+3G9BmlBNEugrTmJtQYV0KNQbYGNxqdR5Lik1Stg++r
e3gU3zOjFdKUUUZ2jOGcO3HF2yg4vPKZHB2aiI714ur/OZIgrPpwDPJbjshwB6xoP7ycDTGaRhLH
+WA6tiZUYb1NC4N3G0bVt6RWW94Fi1/J7FXCcmhhT92o4aqVl0ULB+cqW/URRjBJpredNEeSLrW5
ug15qFYlCdtkRFJspFi1fstpT+LMV7TUFDm7+HtDIHJfoNBRwVoYIqcAwdDaFpMjoWU7qBMDbccL
i62PbNjoo8fdeUo0V/w6WCC/ktn28jhF5jLFQzfWdKKMvT2EgKRIAxwo0a9ExOAY1fHd/eYTYITt
0S50vww6GR87eZBXVw43ahuQkVpWMKb1T5GEZRh8EsElehDJ0EC5eoFEFrnx480VcM/dnjKnW5nd
rBb7LtNPcbC4Ld5sFmvgRotnRWPtrT5MbfRjNNuc5od86V6L3J7JP51lplsWHx0KRn22ZVKOQSjl
sgj7gPh0a+JW+FX/WfDwJP/O+HKKhol092aSgYofWwsDMNMmxsC33WFpI0nLja3bysNL3d9NuGis
+MEhHRHunpztU9+o+Yx+ttK8lPQcQTl72OmQEKUQxBSJhNoX6ava0Mgm41SxVXtdzvDwH5XrHdSt
ubgYEUFrHh6dzKi1oB2nW/SGTYD7BE8/hL2l205hEeWI+bxzfB2ZtNm7diCuSObC+R6+MD2Wez7P
6MJTFMYwKHO9tmyK0cQ8AgBkwq1C9B05fJCMUAuSA8kxDotCLp2mDVpxqtkfYNl1f+G/GHcd7OWH
ltjcv4m1aNBwtnuAMBbDHu8tWqmbfrfLavmaFP1lu1uHnGOouYF5tdaLQDYmFVGEr5xJLFL3T0gL
2NoWFXi/nPqaCunT4t8eDDwUxZlhEMwqpcghHIcMdddHzJVuf/fbw2oa1NDDjGv11BY+S40GSqr7
S09VXMQ0b0M5KcDYcsjegwFzx2APhVBE/g+r5pwio1vvZcI4uG5rYumOb1U3ly6I57dx9KflVrre
CpsBYZfAV6S5vg3mxGJexNA9fmFPVN8kNgHd3Kz4Aw1/qeRQpp2b9txMSGVzQfMRWysSh1uKsoNe
aRwjgh6ECX2g8EPFbwEyFH5RINLv99+7Rl6HivVWipQVIhueBgoVOXpnP/+Cic6OJToR4LlfJ1oW
oNB1yDOXic04Qj911szRDnq6hmD1VgawzaWbwcK/+VTX8VD+1r+fh9PPq+kYSZpAqImhiisvNoR2
HQvX7FKKgdeiRBHNqu9H5EnpicGhzvrpltmapGK51VVmGgbp29qJGJ3jXzyRNEYsiKwCyU/44HGJ
82jZ95jS/G/WT8v3JELLrJCdfhUzssA7qseVmsxwdIMWSSY6YFlssV9UTVReuvgHOz45ho3jMRc5
Jxe4zY7z6wp9yYDs/p6/vFPaBP/fcy6KHMbSVDNIwzZpXCYtNh8UOXkb62cg+ZI8QRMo7Ta2C9ts
knRb1ivdgI2JaVc5qU+eE4vz2r4wOXzgTdnyKlXR6oGcuALU/LuQ9DbJYFh0+oFt4+GX6qoX7ee0
r+wEAx0nTti9R9oBRC8dQtms94y4XKT/TRqyQr+6HUljrylemr+bIby88qLo9QvFbEO02P4kpUzz
hchLh6eMN5mpSmuDoy+JVdLVi9pZRo3mvb9zeieYuqYCleBKaUESIAr7COc7k56n6tf67kD7d42a
gLjuMGApoEkJ8THINIy4jTsB5vDbtdlGQXxfu+Y7JVCD+jNb57gsJ9xovzwSt/Ym/aysUFox/nI8
zN/xl8RbR4XLAZbc0sWdvsXbMbtSCrvQuItL8iFi6Fsbw9F1ClTlLsW32UcS5/n4vEFaTlHeRkgX
QS1oKEdFOlpuPDoA8/FzwM3tGPuYYQm0f4c4bF8E/MF+okZnJfkISXUbJZBD7Lc04yUvwa5y9ADO
1NMEXwKe67go9Tn9IW/UKb/LFC5zt4s+tUaKmiBabgvlZkI9JFaEy4DIUjTnZ9FSff3SeTY8JTNu
edWnEE7Vc3pMIA3by73PgWOXMAyb9HAu8EYtSWoE6UhusmJ7soFcNwwD3T7MaQpFEWmP0xZgcAF9
ZAOYJ6DFaRs7Op6PlYHsNNmMu47lg23uHwvBhUUB1zjijxMIrxWk96E8lCDEkMiPPR7gySJl05VN
SyxFLJfaZMEgozegaWqTiEjbhKRRTONb2Vn+0J5HOGNuzdODkdGw2bFbjQPgGFHmhRHftLhGAwpT
hR5Lj/MzSOZ7NYnMgp5ga/9tZOSObOitT6RjJ+oxdlVPHfBmd+XoK21YGmKTw3nk1yRb+HX/734H
eQ+4ntLSJVqWD6uAhtwd7zoZgNXk10ktgjXP4kv76Cf+H9fo+5VVUtJ15GUr3fSihnCg5+X3EPDO
MEi0k+ST6T2dxhVPDruJeY7xZTTlD9+goEF0G+R8geeIihqTcyPfkygw4D7Lb3B0D3juP8D3sXu9
KXve91LHC9ZZ69PQjqLKDKhV8vo4b6brOJpwOMN0WwwUS6mLnhEcOhMTRvnroW+3komSFGvnZkpy
w5+mjBQ+/AHouXIR2X50yUfJolyYgaDZqQCLj7w402BvhKbQp+3gou9lJEBy/Juhqj282bHzGvTY
ZgOLbtWLAPQZc0BBFPVOA93tPJ6eTssuGoNalYW1j4r48Oa4SZOrJxh/n8AKgNqnLXwCfjgQty85
gqEnxiKMNbJQa2Q48LBgR9caq19uB6dZgH+TnSFhLkHzxH6stTN+A7p4OlF1EuALiYKtaZmOm4IX
i/A0h+M8fpAsv8c0zZkRmocWaLQyA4ZhqArgLqIVXkcFiHC3DNG2o5tM5cyKCEETzb1MSC6ylNLE
/+y9JuWL5A07LVHmdGbPEmm6VwQhJmESPqVz1A0LKGb3H+BOwzZkby2ERo97GzxpaqKhGeEKUbfP
g5nTmMahs+14BqyImb/9eZrPSl+2W5hMNFxD1sWmtQuhy46aQDbIEcqfCjov5FEEMisLu8Fa9Hdn
i2ZNH0XOKJW4o44Sr8CRGmIvwMtPw0Rb0hpx4vFLlAeCpPOyqDdqytRHYzLSnF64GvYTa/dpr99S
5F6axbkk6orfyhGOv2192gCNCjExShWWGQ/bmgBvcd6q7XaAhdwAUzHWCBa7iWaLGE2Na5oyvrCh
VIaLju4+O/b16pft4PVkFsQAaQju0zJBst0+9TM5bJatXo0oFAo6Q783b646Lj5+quM+/Jt8Bzue
Pgm+q0AZvqKbJT31NaKPSm3ZkvXZgFBsXyu3R3jEIjj8IUgpieaybTYLK+/KRd4axAvnZQfCmKtg
C6NCiWbV768NvGE5CNJYC3j1FjjeeIqx1wfkQAQliR6hr6ilbuXo/VFI
`pragma protect end_protected

// 
