/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
CaihNQWwu+qKJWjcmdIgzgKIXQ8l3vMImmWHnChjYqoa51yMcErBScyiE64YZSDih9WCUqsVfjEZ
HfdPZ9ljuyASaDAJWOBnJBbhrePBDPO5jKkFmPbv80QoBXSWaNMFc5sW0Ulg3lCiE5qq9SVr7IMd
vkFVewJkI9IJKPXIqEiYLMio527A7EkzJrjUXC11BQnTYghbA5n7/6q2WIDOwjQ+BdLZXxGdIUKi
ihIieqBZEgdd6vwETSGv3sSorIwnUPSueC94L800xEEoFQmghwgPGvLA3IEIqt1YNZfrY4rcuvTH
rxE5ve/ar6tMYP0QdSitAf/UOVre3EWtsP+Jcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="IxINXwVvXQ/n7KwTaYrPoEaEACBK27oPy3cRIdl/LOI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 880)
`pragma protect data_block
EiGu1ShDtOnFp1/lwt6VhcUR8yhnAB8O5e1xLbmtU8hFkeRUrpaBl1HAfyRFT7nbtX9ANec6bT/6
M5F1wZGG5qSvkCUW8yVN2ibhwe39b3gqpxlAM0Rk2b5g0GPQS0EovauYN9XAQquN58ggK/O+KDM0
63s7X7It+p/RSFzWWRGZS+v0XTm+D2a1XMT2uisqh8PefOCoBySO44oktKTY504wlCSc5omNSe+u
zOKrUyvkLauqfVr0IymzexsmShoC8a5rxCwtiHWtuZd3ISZeseAH4yuuIE22EaResPkSs0AOtuxW
LUa+5ziMFj1jUrwyX7edUaYFWubmHAbAkkw9Hm+C6bamM5RNvdj0nJ6+9kR3k9JEEwFcMnpU/+T7
AyStZ42jqyndQBD+fvcXAhE7unT9l7MeF6FPz+f4fj9QLQ9uKKfDT4Z/nUyAujR54s7JMJPusI/1
6kmMjc0VDkHnbDi2wkCweAVtI13pMf21kgykit61e5wC9yuUa3wMmmwN0K5j3CFUalZcs5zyaUEU
RFQ6sxbZKoizpkyYAVpfJ5ooRM+2IwCcC/xaZGuC28xR1sA7FuTz8gJHfj+31ej4SmCB90pf8a1j
v5GMWH/IC2k1qDCu3Nv9vlIh9ddPqzd8V2kbzHKQIixQUYVEYd6XzNzpOSAo7YP0yS1vkaxpM13/
tmu8VZm2h2JkrlzFuDwth9ORNpQM+dxpUbIiNRz188RAIvel6yq9G8g7YjGY6Jq1qeGPfgm2uqIE
OYHDHJww2kjAzMfBu4zQRXixjhSL5YOVbevDsp++Yot323jrunN6b3HYs5T3zX64N23723OKUorb
BzfFPVvrOEw7oa31ZqgZSsWbWZMOkcIa955Zi5oSnEOq4KNx1IMlwiRrRVmeW2nzDZyOT/6kkiV5
Ay+TkZF19zF0PKmiNq0809vsxErEHL/7oYdQDYLNmot/tAe+f381qkRVEbZrjA0uWw8e7xnBZXdh
276B2htPR1ezVeOX25aKI5B2G/pH+lUnzW5CqMGEcgS1yReFHycsSdJkPGQDl0uTLiAZLicoj2v3
CAT2TDbLr2Obrdb1Xpom03ZaOT0ImqBumdzSoPD+eRvc0qT6AoCHxmNojpf4C2WADh3N57ctHcPk
V7HEOkM7H6joRSQhUNMkeuqXc/t6IH5R7g==
`pragma protect end_protected

// 
