/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dD6sJjMckNM/hk590wWgo7QyLBP7qvuv1GnV/mfQB0w/i/pvS4BJcnppdBuizaQbHZTE85H6pboO
mTjEC8kS1yUyaRKX4KpOmRsaXVL7/iV6Mc+EyHoad/3cx2lAwTCRu6nptqi96Q/dtiPbQirlE0cr
bj2VslWvQXYp7agPImHpkldpbIx4OKKY49/lmZgzjQmz1uAl0Vpqn03TZsorFhKrWNa1NL2PWEvy
H6r6Q2NnxwJibsxIu7/DaDQZ9tx7P3Ox5rT/+t7OV/sWKJMNsqkendhSkyxMCR6Z1Ip9YxyEItGS
Bld1ucslP9zp60t9CzMGZcj/WZZ+ve1NzjV/uw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="NlHs8opBWv2KH1hFnLsdY2EH/Cy8LVzvJ0P9w8zUaYI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 321232)
`pragma protect data_block
jOrE4515xgbASXSOIDgmJjtzDbqqaLfnwtvi6R+i6tx1cVsVCss3SP37f6NOzSsHGetITG+Iu4KN
NfmraTrbAgzjBZhgpQ+BTQFERtCc+AuVe+KaGsNV3juGSbjcSsj3oEzTYbG3rBHCjYW1kq133NWZ
iihXznZcrva0Bw2+1VcNs0I9tZhOVQclOHk6XqA+ds4NC0jHd7n4HBdyo0RCtgcT3SeYog2CRhKn
CiuJCrDH8vQaF3b5n/1/QSWQHMyXiBJALmHGytabtedFP7NtoFxpuEmxIheDEpifJvG7w91hXF3t
XeFSbZLK6eLwd2sOEI0hDM28Ysd0o6eLIUwqBVsBgrn6+S64cpUs3F252irEXWw9x1F/bHOd6y4v
bCdS7OTHCySlWUB5kFqEY+GlXB/mplertyqTpHVUJ/JKZarnyCLxzPDX6r4zN9y+P2xFYQ+T6WlF
Y7fa1usKMX7FRAOqvYxVqRUHz2EkaKHeWoHs0OKxH+ZUtz4lPB/DJwt7WJ7eM/C+AI7YGO/aEG7m
bEk/sd78zkz6ryDgHjX2v2FjP+L/HtX9bzIpoqXFMK7+YjE0+i0RLb0dS1OjfXJuKMDZrz/2Pfj9
PBYkC1RLvgoJiiW8qkrQk/CCX3932cL/gLkFDjoOVuG4cRJ4t6AqNmd2S8fSrG2mJYfM6ADXDf+y
leg6dF22OjI+9H+eWP70rXwrdUQ0sg0iFS4Bzf0TxS+FZl8bLb81S9YSpqg06E6RjQU6KzInYLHs
Trchqewhil2rrpr0E8oER5/sx5l4k2Etn7nuWTFsRDs132v6S6D5CVdPAhe76KJDdM/+UGkLzceH
XA1a8lb47KwdVNIHDqiZE2reahVnsej70lzBs8fnjafQtmkkrrpgPa7jTOYuU0YqpAxc1NeLPabh
Q5EJHMTvkgbN5WUdHRBV7SSOveTdxIMFpVors3QBwhYE0ay8YUjBXTVrEbjD4E193wEYJxomPJY+
zER+3U7FYSfvxo2apPUAADfrvxU0apOgb1DJb0837rEVZVFhGr8V/eV7SVQTfnT/Li4EbYIzI8xD
jnJUJoI2tTRsjiAIwJXgrYZiI2ChOeQUo08apYnZcvPVTxpU6lv8AzRWyuvR00Ab68uZYccaPBzc
v/6PgOF+uhSKqiOiuYWHtOkQxbnOeyYSQOv7oFdRJHYFN1zLanXOY21zqQmqdLuao7FF+bGFF4ev
dWXlbu9DfCRkCcgqiiwFhL1EL42z1jgS0JoHm6zNCcqVdINZ3MjAHNclVwOV+v7mZkYLkptFrxIS
8KWP8YKQMGtCUCla3d1ccoWUxv+tY14EbnCaE/IGMFFp2vdQN4NJbbHTjKGHxKD+xyEjSSpPJ2D4
yIJMtFtdaM+3j/LUFDSHgi3trq150C6adXcyiSaopbf3SZsF9z1xAMj7OC+BAEkivHqBoqRKDD0u
yYG0/hLdgBO6jUvSMbVEXUkW3A8lB12U4gxdjqmjCHTBjqptoV8UjPeN/vSyidV5askqdQfm8P/g
/reny/22SNOjhDtyEpV+5Bo/t5GmEDfvOq0XXfxWphhZ6Hgs9umPa6ZR5371KkykF5Ej1oEqHHDJ
VyzXo1yFkKgIoy3IR7lEPBHzXe3z4/wlhaVNjPYS+u2aNKOWevLSznXv5/TRaKiHx3Xyn5cX3QB1
V2XROzzRr74TYW93gczju/vlmtc4k1E8Ko6GL4v5J3LgqOxCD8BMQtc8cSSnLVzXtMj2gbRmTsHF
fOiiHI3D0c3DLNxYomlcainOF8t4SAlCOe7n3aw+IZ68U9bBthfhROfqfLk3rZykIncuSF63jLLE
D5sPT/btkiBfGvnaXYpOyvU/L6tUwhNvd7Z5d5X4Hq+31O1GU6aRGVxLZjz8kadMo24buL382ITw
lSNIVbdDbPpUbpDX5hOjkD3UxUMLcJI8ppIS9FH3zRlKKEABiWDq28oooA8Oct7nRDZxQgqdj7UQ
AJ3ecq+EcYlHFQFxDXfVnMh2ULhA3b430kBYmM3Rkd2X3U37rro6znVQhCEe1X+qlZNlYPuXHyr9
TAAsjV2LXz8sf3bZvLnG1y+ntCY9pqHDPBOk3Cvey2A/C6/kIBEhuxhe93wTnX+e/HtQHEblHPLV
M0vvzuDkmHpMXFSmDzD56rvaDne4CLW6ygVIJYU6zZU9eK771Y9KL8YAcz0lCGjZjfwfKIRExAxw
Q6lsdLh4pphqq9hzGinV+S1R5JK7XM8RkqLCVA9Nl9wfpv0AxcnFYBwWdVveAxo45N6UWt1LCk3M
d7qSKaD4jCaKP3FS54UcbdJdzR/U/eRNsmaqsuv4pcPpnDEJ/PcliKeKVPVhqAbc3P+Jm4SgVzUz
S4DnVZMfxbWJXZvwzKvlcED5kwLVDtEkJD9izwntMNCVce/Tl0odbqn7iwYAl9MIjhiFF/BZ6Kg/
0Ryp1vqd0hOorOCUu32YnyF4H83eQ/AEXqvLVrDjdMO8y47Gqt7tBcTXm9QulhX42ewuhVUNfnWj
/pYpVTLbJTJesbKhKC84bMwhTzbnUAnn5UqDwd34NDMbcZ163xwp+/lFTt/Ylsai/1JfUCw6kN75
Ot2oTkRFdSQsm/2B8E/doS46BZ4mHI6KZ+utSbVWt0A0TWJofi38d8Jzf09W+lnIpSQ5VuSLtcBh
oC9seD3U9yzGxBkDA3hRxdxQgNd6yVW+vuKJP5xUzTX7hbP/5WAHUVgdhU7+3nZ4aOWjTzgH7+Pi
2/skHcvSouhwFcUV0cB+uGXSLRP3PwwhD7/ayTCGSN1O6SmU6oPPoqKDExl0EL7az4bE+Fg+6+JK
W4hYmlYQFtIXCgq9Hc8mj7EJDNnJcby2dUIQk67nW+gAqL1PY5JW1h75qpeWoKRqm0QET1PRjgr9
z7ktx+lRZbmFXIyoaYDeZrAvRe6Iuq5EQmV0lej0qeAY2xs3KpVM3FDR9fcCaEURc+JQrhsgLzK0
QevpPS+cLrxSNH1NOCakdTT9LTUcd5nANKi8kjqOzKZVr2oXjmlxzwMMtWfUfLFlb8OeboyXjcqU
89q0CNz2Fn7YIU4eqIp9w9CrK/x+yF/l0KVfCyzoNcjBXSq2Pfl+oWFqYJBhvVVpY7VuA8NZ+RIp
E4JGJqT8/l2DCEnbslL7EnjYpWdyMS0QS2VfkfMC3cGdLsDCh0u2oqQ2A5klLeQWf6L5vD/fBujS
J955RbgeO6osCCt8eauExWlQDr9W/KBtoqQ/XFT+qRETQuJe/EcKfahOJgzzCqGyIo/M/uupKC7P
8ysQ/Y9dVEqoYWiyD+IYDYmEhX5JiiCWbsK3Ul8mYoMpm4sCeZqoZ/nhYiFUQ7TXdXa23UpBrzHd
kG18lF2I+UD6x7baC2uVWl4y3yeeDC7XX/RTmuH4wP9hJ+2Ls+KstvIYdPAyqjHRx518NRr4oDqW
6fcFmipF9QEZuSqyulnj1KaZv0vLDsD6A5K8ADOjPF7+/NLrhhf31qXp5+3GcIdyfUfvAgqQg5wK
NvtB+9oid89SMarjZmzQ23lDiDR8EGuomTPVHH8LCB4odne55FTtxIaDpGRoIiPTv08s7QA1MKov
YpUqj2mNARakcXaNkgg7v1oXl9oD7Q2lCPYfcnjgjiEhnvP6oO+i3SxQ95BVQSLGPTa54J9iIBJr
GaADI7qXBGtUXTujnTnorEIzz22TOHWg3hgR+tAlJ1Gc3GulJt0On/oEPnHM5Wvczj5w/khccY7D
9BhE31tcT75LqwkQgvKgzg6WosI0DRaeOP3ISzt48OJd/K//XDtPLUIi5l0XKfaXPE8NA9ZKrRAE
j/KJkUD1zDi3hq5mKFDmNe9Jis7l/ue71F9iFmE38gcd8KuUy2NNXXcSBnY6XIqzOg382cyyCtb6
273/RrA7mls0H41xdOspVsKtMjUiAZ94/uPKM+vpJxeMb7BBu//hSb1kL8CmH2AMKCe4N6oPHvXe
9Bqkbx00bT7frCMNt607AppIN3oO6wfv7k9LWkvvb/B34AN8o7qiufGQnqV1fZLrYTHmpNdImH5j
Ub8O8ibINKdmZh54fbSdQTuYBe9LlmXXaIx84Zr/G5FmHSsVLvMERTvzDz4USqcn5AnNekhjX0UG
XiqNpKAfWj4amhaS8bu5OsiA1XUjD0ah/NZ3zgbKX10Ma5kIryv8FjKYib3u+M7+aItoI5bTqw7v
6/z/7rraQIX5PLHGvcAOg3EKpMuDhnIkgNFQZHRJx4+fQ1+X2UZHMDvgvaMD6Dj00Mv1eGri1WEc
tgmay4wt4hcWw7xMcOJQ/0La5Qq8gZo9BjO5qkGxb5jUcOf8CRNakRz0Z3UNlSLTgOrZnysRm1KA
NhZX4HWoaiZ03KMvoenOwDN2GVewwV8j27kQnEewygGb0cNOfgar0ySKaEokBoQ2LLLWbavbsgXb
+cNjXmlDDmT6FKGZiuS21nE0mUF3urRtwDLCS8goB+GmJF0Hr1P/fEJWptylHFuipXCKmRrUACf+
Orqvnx9G1gikmjT7TPxOnFkAx2dt0n5jVIvOAiKxuRkAo0Z0AdPTzNK5ApqdVku3TGgjB5k04vXx
jl2D247tX0etEcvmKPPBYuQTpbM03fH3GP+6BI5tbUvESvnCGg7trGwCPNxzKkVfdhdiTr2eNtOx
CConKXuODIzldy5yun3QS7xpbsEya8Vqe7VY9m5Nz4Flybp9uFcHfHZ5XiR3Gx35qQTOahffSvYk
T6jaIGj8E0wIwN2+x4Vq1tJ7psDdlDY+pvqDrR05AbmId7tWVO/lupZxuq2P369XQaXfZvm75lYk
oo8tYdlcLFvIcD+bYXMd+aFNhKLk2no3HWlNHsY3P3m4m+LEIdJlX/7z7+YbHDkzYdS75s+t0rE8
ukOpuxJgOAfuwc1nIIjO9Q0265U8gaqZhc1d9NNXx4Z/pr8whw8Pu1fd7GzChWnZB2BlcK/jSoo4
FBwe9JnLMtrnBW5DvyxlD70iQ7aZHhbEvgGz9o5LAMXUFolbENKMpvVgCzqQ1hhoCml3tqQwdBIb
IMKzF5MjQfB1Oz2VWe3qqNN25Zi7qTTTnC0LWeSjTs5zJFYYanw+kMDYECJb6UHmPIiMwOLWXWgG
fAep0Nx0GGYgQ2Ao/7a2QhkqRcvnz2kxBI1IrQEAHkAtRY9XmSZJz3D2hOrOVY/Hmc0cAcAzVuNz
Kf855/wsZWBt1eb8jRnAVZlgTrnqUZEyX8XxWKATiMv8ebW7B11eaE+cMIIpsgMHlsdpELN5DCjH
TnsksJBFRVWj1NBLSIXgvLZIUMpgrqQs42gOpzE9i5qRe12NebpSAzez+PgNlEpNnxlbSsBD7iP0
1TT1Wya4I4i5Y1ZMHxleMas3fi5YTdDv1DGMe5H/uM5BAihP0eP+HlYObDjEtmPvQhgmsaagZbwY
ESK2b7qBOyNq0cPcsrsjaNZldqqfvFQdMH479XO9e0c6DGiSEAIV0a5s+kHKR0Jfq2HKAEub5E3A
0ouzL+ndiN7kfXoBQGnAEi95LO7XjS0OloctqEJAzTMkgZz3tmTEJxUxtkFI6f9OGBYFxTFSKzU9
sttBirV7WusM80/cOFw5Jyesfx8GYXbYwEVZcTiH4lwSKB/CWj04ll8iBFDAVvzTLm1tTeDvA5dC
upcpH8wC19UuqWG3wlNgivu+V3vkd/k3Z5N/N45W5xdWzvyDxVo3qhGVdkPujcPApsfhEjEHmr1S
kqpedbir6ueIyllqPsYZZQoulwGML+InyKJ673/n2kuIvtbLo0PdBM4lPShog6P69jJCuHKgJC7A
HNxi9xVkYNsD4f1GOQGybuQu/BWgMkDCPw1nEZ6+eszxGPwdVnLC54VluRVbcMSXejy0E5Nwl16K
gXSaOjVIXwrBp2rGDwQzNIgrb5pvfff3fKOx0HZIZewN994asrIAypYN0xh4BnoruARuMBHuhSbP
dlDWGtyXbQvWjY69Fe8G7JWpCe1OaEBgNWM1Rb1Xa2feMB9payVApgfaagrMlNnpFUXoYUFQmdjv
4WI3JETSIXGDAA4dQQkBd/0yEoGwHNo6ks6bMOVShRqFqFh5BA6kGV24QYdznnFwg7Z113oROv50
YaeiXIJCvsue3EvhcnhXspoeUmBxuJkDCTjj8ZyE9qpL4yygsJCulroAuCDC1eTzAB7bXg8wDvkr
we6uKZnKbCk20WMsQishcfkXUqraZ/Ss4xGcSzHnoEFG6TckvKbSY9D5bdw/juQOSbi08MMX/r4C
GUeH9Y9E3UmEyESCuWxiF6LyovBnB4MI/n+J208ScYYBpyjxCayKrFTNIMoLurIktYGN+1l1wUXv
SNQX1/9r26yq9wDnnhz2lwPl1gOoJDLXD7/N7dCXUvUMW+JGnGuY35VI+DtYKRiKZS6IA7ILUgNP
lvMXWtmYuYoEcBa7SSoGjJxjancZBhZEXY43Mv4da29DKmQ5YGay0d5l9JyDiqSg1O/yHRwYZyNL
Z+9bk5kX1WiltaUdtcmyrdoxU7NB7vUrv9rUNUiCjwfhY5COgHQMLDJ5d0FRjNU2/Dt/WoemHO+v
BhIvwqQVWTzNJVZPTWaTsI7kx0IupCcdEDS/wdWHfFnIR2veTX4POIo8JAofbYHUb1+P6Mh2aGXL
OYkzBB/fMUeP7iir2wTlB7ncDqgGaI3QiEfhEedDJuWjBEd8ix5SWlmp8fP59JK4UhZcBMF8vCNk
i2Rx+VgPDAmAVS19Hzb/zuEDVwYLx1A/APCJD4IVnrOEKz2oA6Uk/8nq1VVRWaPTdqqxs29TLC4M
hU8v9XwVASVQHr7gdSp8ToPOm6Iz4jKPR1DXP/JAfNOqPItJZMYPK1JwlAGvSQTDM0tLUusyTJHR
398TeBCvoNVvMuiOG1jHa3OtjrXk7esCpm37ZxWCJdB+m04o9blb05FD4g/zd3zUkDkzjhA/kdSj
td0oVvNqgxyr9OH44Ds+r03r+FCFvTlchAissm3EBxl/8jdZX77f0txVQPiXtTJQ3/eM8cfNO7la
UvPEski9STdx2oROooyCapaayHar2N/zYsCr09de9GOwIq3aARfcG7VKJrXJIdtJkRZogpQY5AWF
C8RRcOd4lly4+jxhwLiKpPDfV5kB25Gk5C6NRNBspCj5O9HBMcVFp4WRTO9MlD8no1ZqGA+8D+YH
oqKe2Jiwlbse+day56EPIWupGM96JODUvbN+2/IKKVUo4xv3e54b0FuFU8ITxnukmKTaaqxG4smp
/tPLJeelhkiUbeq0TJkP4VYqZiq1SSRPWQo4jLvbl0xyqbfhBDzPlQTXflqRvNo9omn9w3HelRgS
gRlRrV+49crRELK+1858bbL+FXVjySacH/oyHiWkWRu9dfzYmTHetN10XaePQBHldXf5xNnzCopZ
Yf45Tj/01E64E8VfdlRy1eJdZE5bIIyz6tiV199C1ZJQBlVQiFheQk/pjgZMZsjlN0TmgFa1k+Ix
ymn9GaHco3T9AnWlWflC0Uwf8kCJSZuJfn1GrT17O83xBmg+qI2V3rWazcQrXX0hfpQ0XSMjwfJL
aP2jC62pWIC9tO9Zp2h3zdk6sf0d9F+Xjv2Mki61ma/sPiluO6t9nFTZo3MVlK7umXSiPvGD0OPW
9iKjYH1p1oxim/o6Tx0N/G0xoTU/ZHP6dvD+WpCwlKioAuCeZlCoT5tuj2F63oiMVUAy64gXLNnP
W/CAFhGQvkfxkbjVgIp4fEQ5OviZM48RSy9QeExD2cSJ9jhMOZbQMHgHPZlo4VswkQ+/5G+rqMhW
kLYUyOCbaoqgvF+HHWaXMVkMg/zf6+5MiUSyfrIuQ/cvaPNTHzVanlRPIY6RgwP3NETF2I6CB8eS
ErO0JBuOlYY9XTcB96IRz5jFq+gQM17W1BpvR73AgjN1TAtOPJdns5XyteHN3bLhAadBoiTO+mxY
Pd7b9V2rLZ4o83BxT/eSMP/whNrNO9PTlYlwEdUm8fSUVNXPsQgGgbyxPlsw0jiyH+IOmDut8Uv0
p+rAJKmw3BP1h4kdyXANPO7iC9T7t6AjEY1l/C5KxPT0aNA5SaA3Na9UchdPco5exNa4Cg6cO3MA
aoUIBDu8Xpd8FjEFsq01MmkrGs8JiMPHgWSKs80dZW0f/NdDfkLMhGbAYCIRNC8ArXyUz56k5RWG
4XeYAjR8TNQDhJNycMFeSRdXBiZYp9IE9P2RjPClMeOaQERWX/Mkg67B+T9meriJUMXYC/AwrVQw
l+9lr6cAJQyQHsswRjCYBeox7ftEHNXp0Y6oarHp9+lZjQdmbaRO0xpweXOWG/w+RhWpdtktjF0j
sG3mssANKKSdsnEW1MCnBUZpULib7LPl8nc9HJFov8Vmi6FtXvVf8xiU10wl0LmfGxghZWP9DO3+
AfH0gt+qesooXebfCI1f237bYxSrdzKPbQd5RMbD4QqWcZdqLS/FP1qyXTP0bG5ZfmZQwf1ykgR0
UOH+J/VmyVEAVOTAuXpJEABPlnMIEnSnsn7hHTfuguiEC34Rm9ErvpswYSwo+312bFeVThgE6xaW
aHeo77vPdqnIthXXkIDtD0IzP/wEvzxXmakRNzzpA8Yvfjpd2OmlzQbUc0isT6CnvWJxhvYI/pwF
GpAByR42pC4NK6Ah43qUZeFEaZjDyyEsznw1ZEBAW9vGCdfH2Zi9hk48RO39EChVOQZjmRVziis6
dguPtZoJ06kO/YiQqfQZgAy4+/4R7rEeYh+xGw55GRLlLemc4NPNAuPc0NsagkJEFWnUq6pI16m5
2rN8Y+PFZuj/UQ1ghQOfqFmc6NKRvtFHP+qokNHhqAZ14S5CObUK/krtqGY+qGVT3EU2Mi1IuyeI
Brxiawj5zbUttI3Yof58qY3jESZ4zlZEe6djOswuBmUGC3gViMuIzv12YGKi3OQ9xySdlQ5RZSM/
7iyHK6CI07MEQn1DkwLswxApV9foVd+cGoUkRmZgT8/a/8MoJ0Z0QpiD5PFXNESumAWPv0chvvD1
pe8ofgiOVHmmg4GeOfoPUVBWyWJffRlfEJPYbel/5r72lzfF/LWgBo3zErtj7pDcdNCePyXnhQHc
Z7r9Zx82OqtKxw9UWD8Ti8zGOg8MyIMe5gV0pnk6rdZYoEiyPUsTKIPkbL8igyaDhqud452JXcuu
xONyfb59t5531YMqQsheSDTTC9NNDPz6YVyoPlchGbkBtON7Pxc3wyOFXKxMIqfQ3r9Ma9bd5gjT
AuRjUg1gjwADWKpn7vN7M1YTbO62AVk+cZPbcO+VMZ7wYrzo9rBZyx6idCyp1k5gqv8ee7h2pTq3
NJFT2dNEFQC2DbdlIt29NmN1/h+Ob7FDY348ZNDznqRLCxEU1oJq5asR5c3TSWVltp2QXZx1jDEZ
PM8z6U5MHyQ6CQ8X534A9A50dleRRbyCEihWHOJJ0wD98DN0PB/S4O3BEUGXwQRWNJR/3IfkCMDq
gCS6FrptTgyUVbNqU0TN2T9gbG45pysYLQbB62VvpPKTCkpH3PoxkTo9rNj1uDfMfczh0+km1NrL
qQTpt+Vhrpm4pvGqPa/96g1K99ybaMclw010nVZ+DqlKt3ovzfCBxYYV1G0d0gXT3VD2SfLJDzxH
Zdg043wVpuaP2daQYiYQECpmilMYPhvm+Xeh4KZBSue1TQil/i8OK+55w9PG0CyUFNaWHDOvJvtY
esxDFP27rZsp6ZuyFJkL6pxp3ogDuUdPMWPe6dIC8ksb03ScSQuuj3CPTcTIM+RC+k+qJNgbriLj
F7RRSK/AMaj+fow/Mcs4VYO5fVotpnhD/AYffRGOPg3xOUICkj3IlaPwAWD9ssj/bv/itJoo58Z1
NgHVWBZPBI8DH4wTAh8O1JyqZE4mmaG3xXD/4XFfqSU4C+8Rz2DZ1VMGC5wPDG1d4X+eIRPADCYw
+YH/L1DU135R33KEtHRvfl2U0y7wJdlVonOgVtWR+n3WI30/MUgb8s15YjcXA7rz/0JzKQETbvBE
ZQAaMLr595BqsCB/aMF0EWwnd/VBCpE3VQ9IPCdsuRDiJnUH11e8dAtxINZ9WnWVM8XX660QcFYw
57bZiw9ee0apaj6TZHUhehv5QPOZHR5UIqpWeomnkAvb/hqG1uN5WmEkI89RJwPavxDLSG+lCEex
ZdOVSfUveveSqLC1BJRP57+YbVysD8JLCOFMTl8CBwdj4bSXM8HwzMslQw4QPNaKVD+X5J+onQ82
kpe0eoQrxdrhJ7dXDWnx1hm+jr8oNn8Db++DEG8CROLhKShVKINNtK2GpO5VPzE5OWs4M8PgpnZ1
aRRHKH+XXpvP65/y5MmBFuwFfQKV5yWJ7BwXLhWotmsIkeKnO5//Mg0zjko7JHGjWLAkRk2DAjnJ
n6fhrw8BD+R/Q0IxF0+Ks+kkMJX9JY6mQtF8/llkhNlcqg3kvzK0H8pmAPtvlvaFv0JHM7LioWqq
dNWXz+2R2ucOEYDu5UT6fyo9tgtxHAyTT4m5T1KwJNqYP4hkugPxsBB142vgSatioKD7MvM0RaTU
h+JgYGeFCPA7Gi0dibdaE1kbFYeYakZsyKUdvl47CoU+DvFZnvvurZURI0jWf54AbB7QlZVGTSH8
zu+aJ7fuTBUQrBpb17Fbato/75g88UdPpn1YijNscxSEAmcae0t9Pl9zZHU+g7/95jhK5gXbct4D
CO67LL9tmxYIgkt1x7cZK7D9//ZVYvlWE9ut3VXg1Y7OJx0Gigg9py+uTng7qN55JiyFSDA6aqMj
X7Tj9uNAj3RZCECbOW4MdYuSlFFr/n7by5BvGKoZcOuB4GjZCUXM40VizSRJDeTq0kLygtZGTJSG
cJCY2MVirAOxFvP+ZYIX91Xr0ysnhTZIomqcHd0gepFNl1yCsQR/BC7+OuuFNzBBwDAP9QqOv3Xu
X/CNfOJhpulhp/RlQAXIIrUfDdB4gTAu+N/XAJjpb6YVFidkIsNXkWlBkcU4bLXpfn14Uoa+/LFK
MuX5nGhw538MmuCzcP897iQ32bvjV6hpMvxCPVFxImJ92JYLcFgWmCAUv8d5TW4MLZRMJzESR4QG
xKxWizbGrCQzEWXLtbhz95lquSUaCQmz3g4UiFnRtPWiotGopRttIi7U1frFW9siAUxKvgIdrg4e
QXCZge5eIh2ziyzSPOjXK6RrXbo4rkj2ZkjnSfpdfv9ylEaempv9OR7Klb0sG5dHXKsgdzC3Mf79
H50AtLZV09AQxJRxXsE1RE/ma1tU/eCEMzBwhc3K8k+usEAchguLVF+GOapUZ72S2XNEx1ZQ1Ug9
wsse/olm5wiEgXcak9UOYVH0QvKkvTnvWcX4sxsp0xJO8eF7xZ0KTPTiJpiy+R4rgzZFe5/DSurI
W/Z7umRmdXMaoOQvT76T2gsq8v/hgTGbqZwkWGgUxHSuIK3Biv7Zkp/RiStD7KsZ7hAo35p8pphu
18xi86HtNFsgrQu87dcZ0BUZUfmK5dGq8XdhCdCNRPE+9zckIGL08dRdWqarFNNH3sAwrthn80oK
R53c6pj7dFeFafT+la1/OmWlIjVqu/k9uo3idPIfbw4aAxtPdTYbd3hjX0Iob4KnPW/7OqgetPbX
BlcSusy+VTY9P2lDtzpMCy8/YbwD/SnBg9rkpSc6Q9opZGub1+D8ahrdK9kKQvVXG3rjipFxlOCx
fGcu3fCFsZJRv/dRnm5YyWtEQQShM47TJyyUTof4OsLgS/6DG9ONA0hLx94HtwSOZLy/yLtiLgHo
tRg/692Tagg7LOLHFT5tdwB6bGiiiG9j/Fk8KbCtN/K+qpJhfdtmLJ1HOy3SxZRtHqdJAY1oQWi4
pS754AZzGQUVenQhOl330sV/RWDHh1Uy8OyTBP3VBATu77BM+L3kBk+KLxFdAfr2dw/cOF04DOoS
zzVvEzLyIvdEZOp42hAYZZtwHK8M2WIf2Fia2FHfmR6Is7owVFzUq56hBB4MwZicicB1iWOxMCrd
Q96r1cSnUEkpV23RszxLbcZbZg7pAUf3Gym7nEoHmkk1/tsuwyeLC416Z002Csc7jlZ7s6ESzi8i
ebyN4rPz2LIkKFrG+rWkL4xbpL5OwAbC/b2y5cwy3PoWoWfUoBHJA3srXcl9LmeTdijNFbyJ21RM
LHD/t/PIXmOhms1g3A1wQ916VhuYqOmESPgH9I5nDDN9emdfrVXMgVSwhz6nWktyHI2aNUiMtqiR
OjNDiNU2qGxRPyoRl69oLaWfxgdC44xB0vMQJTizvCn9BfTkatmJ5LlZTNFTbk3MYAv2H5MXAru5
hqE5AJ6XQg+esuHIVztLKXczigYFgi6/1dwjQNv2J/13OoQxQWw4oyM0BTjbUYSUrHKzPrbDUlIF
a7LHSGxk1sqWIOufTvR/gixyylHcF+cwXFcc8BKasOetW5Dkn3o4Xwgq8mCZ1PO/7iO3BpAXYbZQ
X2bI3y0Fa9iwx4E0l4S6zkeSwALH9Oj5jXyd6MCLl2sXpt65UMMSonVC8PmB4UF/jBX1eKPmDzep
6kiXQXmbzbJkvhBAjs4ifyEAWSAliY4ADIyn/adK29NL8bK200NBtyR8tqPZsK4h2pJYKpccnxYO
qYIKcOxSpxGmr7iN7jQnDRRNcQh6xtNtCOPbBt5N7CNVpI0Gwzc4PFpvHpIf/+w9uBN5D13x0ynd
YuuiO81UmEfuLE9h0Ou6SNO9sgnDCc8tfKkgvfyQGyjf34FKeKJQq0a0rE5iVbu+Yaq5DfSfCjx6
Ht6ionarw6g9JbfSLfbKHsLZ/nOjThhWTMEPZTCHeVZAm27sL+h1lbQszdlp33qS8uyBXEn5Ik4Z
cN034wSnwfmNW3XpE/sZlIIPPvbT8NL19vcpwhBN06atCSXW/vyX/N+sC8VNlZxikGWgwO+iOcO7
Hcvit6Ua+gK+JSUTnmfabjjNUWD6fmImjenxVnMAe5YRniGP+3TA0TWbEQHXMjKePFWvZOR3fr+K
eX9vC/AkUwUzbJrsSvR/KiCQFA8D69npnx7PR6hdGGZhFfO60wWfXcTMyQdHzkSEbxEP3BVj9TvR
YEMFEZa6xsZesqpbjpxdWoYZRuPS2LnbnBY9ittuXbaKYLPO/zeFe5z34pKtOf4IyL9Q5p6pc9/d
Two4eCDiWy6HfkrPyLP4Bk8ODRRdBrwjlPXe1TNCH3sLkkmW69xM9g6ZPEIncLW4rkOorN9x+xr3
V7kmOOPULY6aOWoBeATjYDfVJyr1c+gOS8qUlBPnYwQn+sQ4VIU/H7bfKIptS3FFIxCeoy6lcPq4
MO6gDNWqUsTBocCFqArf+HfmR18dvcbqk3blj97UQq+2v5DHod8K32TkejkgPshqXDonf42zUtcV
OElwRJCYJWyVda3nMgBfP2t7K/p8TFmvYFooQJCCEcaqvB21yfBqymOzgODQ9X+3yR7cDO3R0Fnc
nce9enA1HFj+6FvfRsvQ/xv1cyTSpE4MRLMMIAuXgJuxJ2/mADs9zGVLdQWBUOIv87hCzpHMnuK5
Tm9jBWCWzh/4gVym8V+j6IUupSRycnoEnlA0dNpZbT0KEpvU8K0OlRQlqqj526MholbuXzEhZ2Sd
cP1ERmwGyJ1Pwdgar02UD2HNtecllg5NL89X3FL69YGZMj3/5TDHco5p8Eych58bHsoXtSSCizti
xGNYYPSgzAi9NoqbXeJqnGM1a/GvjHpMSqTClDdx7PCIYr2Mr1Bv2G7Ql7nhF8/FBEIN5jZggLGQ
/qLpVLVRkFLsp64V1GdgpHfeLXSPRYMdkTvILm8BKUdaUMxwuEYIegFNRrj5vddtEfyXpNsNJITm
/LeEWDDEPt6oPIwcCAy9IdQxVMu1fwxcoJ9RPBl++v+Fwwi3zDrXOwF5yZWrE8qQEp7H1XNKINgG
LBeARplhl6JdVJJkQrPpXIMEOyhQKsDJ35xpIQx5K61FaHj5ZuKVqLpYjINIQ4ygzhbkOuyBSZOw
nYCebITfVISHGpkfVmY4WlzwvGCAiw6D9kxlWt7/CZovb8dPbxP+bToAWXrcKVD1C00vLMkLkywr
dDYkAABayO+azPuqriRFzX/6L+RqGXU6hUlw9RWKvnf3l/yZsop1pK9QZtJnZnWPJPgmushRiXeH
ttoDaQAfR9sakIdrsoQOmkPS9pie9HOpvw0uYbgmSZ+z0+DUDUaEAeBZM2vBgjh5FMyY/DCgaht6
UHlP+GQKVMeR3dvkHpN1I8q8zkd9Y4rxe3BVtrkNBZfiZtfYgldjOSDxDchyG8CzQWgZDZDEhGSl
RwXpekKNo+KND+igsJ8kKIIbJ9OD2uMKAUUod6kgefytiDvKW/mN9queju1cI/NXdcJSdErtLbkL
zb59GgmCumkistvuoP8to2F6YVjdB0uOrIqDTkEAUo7BdKF85NVBu8kh+154A7Njje9/gTwvVfEJ
YgPJd1kPVLKcnokDyw8xP7OU6fAci+sDA39PBB6T9oPVBW7uKdf/xK09jF7OsAyGiyGINXyPv9bl
FBReKxxH9oXxCxwFYWBKeemlHeSfBUdosqLrVkxhLWYx6UZ3CVgXtQevtDKUCDDPVGB3LcBOro6/
c5Iq2M0/UmI8dBf8+WOlWgO3lpO2Oa9NXEwk8ZVn1lAVoOi2RYezJGr+ygtsHU5DyprW3VBp6kqx
9+w4exS7hLJb31aGRprDco9sJGmjQdDvHkgoSIMihXA0XDIavyh9iFFo3umEADigYDQODB2PEOq9
7bFOuj5otbmRFd57SL6jLUqmsyU+zwZ7YjhYVuBU/5puEeKBWVvLnw+GzrbzgFn3mvyCOH2DeDYi
6602AGRosYSpV8x9U88Sig0qAXnkg1km4rOdZWhdP+PUTSIQOPd0T3R5jVkVX/DbVkRq1CheE1MY
9WFcmJpI5yR5IAi6ssFu2ZjVSJTke7vbmNKW0JPnzo99XidVILvjdKo2FoSMhxTQgWxNYQxpg8t+
kfffVNV8N5JVJ9tKt5wiFEz9+hKOSUr6aLW7gMlHijpUYuTL7HkVRRKArajBu7zkNdRIVgnsXDrc
rvhb+inZjTJr3R/wEa8cdoyF41W9znkSpYLPRKAiIloI4iRzPWe+mREke6+lcyG0kuVil0zi1mvX
ORpj6nTF9rpo1TpzYzTI8QZj5g18LmUIKeciYiw3EgOC8TvWDqQleYxD+wn1FkS/qMdMkfBY2aXG
noaOTT7olvtKXSf3PyrNmzu9gxZc+oxq6mDn6Iz7sNWYGflELnQBoMyXJz7nH50PC8f2VXdw1lNH
oYMTapRIFzMYjlDEvwxEwtmAST2Yj8dpb7F1x+MfOqQY0AL1ZnwXdolL/7O+lWVm9oZ6JnpCirPz
5t+oSunJh+ATxCdAup8QfTZIPA3Dt+bj3oeFXpIzwAh14Oluk7NuzoxjJFT6aWvR68e4xBX9NXaE
5SocRA3h75BNvAr2+qOA6dmdCw3FRAe+I+/A8iKjfE2iSbvhile6ylC6/PRcchN5iOSDv2M4Uknt
KGXv6fhV4EpzIAZrFqshSSKvbYQCjnFATt7X4GnKKbwHZ6OTvRyeh9YKh2Wbd+lGM6GFyFrbidCK
/z2a7OUIIYH+8QFTJ3HHGo6/r84pp4x0Nbox7TyjX9kAT8CT2NkvZy3V3DXNkrC8l5Bn8tG/GIbU
4EG97H3IK6MZvEd/db3ZfSWzYkP+Fl/yNTO38iW5odGxcaMkECQzJYz9tj19aVh6uD+IKsbyVkMu
JhdxuDu51wGw2SV8IAdVSI6dmyDzcdDqfWEYjnklBGKVkbPBiJB/rkLIqmSOfrPJz/kE5jiEnuFw
tLaoR2rq+tpyBJ3FtijtF4vd3CfTFNnPOrOVboIjI+VINQ8LNmgL22c7MXMlo98wayX84UYS0ZVI
uRgtybFAI/qdG5V4adxSEJUh4dekC6Rsz7M0efP1hDQL3KmPqRsqRmt/jSIb0nmmYl84n1IOuQVm
S6g2JzyipEH+gG1MMqXbBNUT11WM+sYGeQwxoSB8Wnrwo5HHQ91lYt8osiA+r1jExvuBHSTAfI0T
CxdQeJbR/FTpLWDV+fU81+AEGK8bAjgLzyS8gDvwuT2dA+7ALh+V0scYJKucRm/IwGMVIvwup7kQ
EdUFQcesgNGGEd2z8y3NPbs4Y8z+UpmSz8th5HEQ5ncGGdoJccZ6IJAD9v1zYmsEc+6U5eGobiC1
NDvJ4QSsCFqHbee07emP1bDElAJvjLZDbq+z+A62o89ZGEoGaIsgkS6ibqW4eZVhb24ETIon7Da4
b2B1AUoDsagUhfbHQ19Dfji03UCXSf3VOmGf75Ixkb1ZYhgqbmR0TEo/O/VQ6xSzgd9Uvs7hHf4c
5tH4rKbPn0/YRjslxBpQ2OPspnWMBKbSn3Wa9UW655niPN4WZyTN2i9lClao1W3KxxtXF2wU0vyf
SSk3s0G/Ue5I0cFztTcFXqgsFKXe8t8CDJLfKYPXw/QzhGgyNRgURWCdCV+73HRLE47fxDROjCl7
5Lm64pYC+e4H2GUlF6/KwKZ/SqgtSpk1obm/wTdTAPvb514Lqf00LL/JKpHlBMyTbOpLxvyfmaw3
HkLIVV702X8H91AixXKtVcfxmw6N1K9GI18sk9fmn249XFwkcLQ9SPDbmkwU8TbM8csN08wqagVi
m7bhCIJejbR9y2KqxkEjz4PfXC8+VvWxWM99L3QbR/SAzIsKDDvndlRxqBsQ5VpPetfkBnu0xDUi
mXqBtXgIibgtm9QGrevTti5AMYe+OFS2o/Siu7C20bnlhpRoukeHNXaP8HX/DLiixZwjua0QZ67J
Aa5f7sh4biFA54+tVzOge6hW1WgCTCIQPkmN9Q8O+/agGy7brxfg6vMc0hZLEwXiUbdEkegtbLDP
LixQsc9GJd/GzcP38pbLw2jRFNH8vXIjEaf/7Yn37DM9y+XSVQmSpdasasamoMidQajfHb5fXX3m
U7qIooBC7iZAaL6odLbTrDs8hH5uL68MCq3X1LDSMfIutiXG62RVkbbq3YR/zwKmgUix7avKBu+0
I+tvZIoQZQ2VEGPatEwHbzz0KGICm2ar7yqvzJeyo9DLU5qK63ZXIPirxLvrs3ZJrGgdd7P+5k4w
l468+6+BY4yH4sBOQ05P7lg63VS+ornakFTjfpzz5+VbryOiVQ2DBV2RUHx86vQFtKYIWYIG60CO
sM51ui3eIoMFYppRu6yvh+w+sQCmOns2OwbZcPOMLg/uugFTD5VWHcYdzMhrTWAUV9LcI7C2+0R5
xURDERvoYS2O805CMMY8piHuhkRVw3xZkpqT/RL97MQp9K6Rl1p6kRk9x7QtERvpcDCFaW1wcmX8
TUATUPViIlttZeSMh7Af0Ql8aiACLAtKA3yM+vW34e3ckfXLtU26ThFvtkSZfiCDUF9u8Hhv13dV
gL0+q6VhCsh9T8S3WGp+92iXLX/2hTjxqshT89Bti54fTETKavf+sGFG/1JA8Rs9ooQpqLY+aj3L
YndHi76oFQrNvrcSmdxEcbmNk+I52B11C5qdcKBrtCU3cpxBBnWehQQ4MMJEwALoZqB4sq6KEZYE
kIkj5qlklR65RDPh/IEbv8JAYp49kbqeGTU1kFNlTeJwQi7U6I5vDikGilo7AHPHFIKPkM0L7Xwe
ttHHItRRX6emAeZ5OOtLKHvZ2+wyHALb0rrNLW9HAVJ/ryvsi02wfZSJs0v559CRJvCk09NNFxPJ
WvZ54SSVwAtawRc9dbjD1XibrjBJ05vdW/tAaVL4C3zifHdj1ILr0NFfCPpOsU3NQjVegELXqopM
FfX2AIm6aBUjlAJQrQcViXYmkRYyDeLT9J0t6qfvi8xtjpsmyTIwOloW8wF80bx54PdqHwv/nNdo
J9JQwigR3LPZqVv4WsvRX4zPiuOyWpNBHiOOzpRWOSRa1AziuW+syzmrkDArhsGRObFZR4dV01Qg
4W4yuK8nnSOL0pPTdoyODljvHOq9u8SYbOPhIiD2yG1uHWpgKTfb2hwJBCk+G3rN8jAyQuV586g2
99xCe1Lx4aqKAfLx4nhkrC9ym8CqQ28PYZVX4wrkBISPPyHV/YamIjbrL4lzPveyAHRKlldNed3K
Tbrim/5h7YGWqIEGAhlRSQTveMBYf1I5H3gRgGKkdkMFKmOmQkTsQ7CjiZBe22/Se5wwvaUxzY8S
wt9YyHQB0rZGI0vYpvrsTrImleVli5LROnkJ6KJMs+Z1CeS2+tZLsV1xuB+eXo/VThDuhO1ZEUBP
TT69o8ai5pgYQuis25Wg2Tlpz1IYtlqjRytJ9LMfPsJXtwEZB/quHiG4Zk+gM2FuVT5JIZfiy/u8
JUeh/xaLS327NLINeN90UZsxFXQY69mW4qGx5fQRPsT32n8n7H7I22Rij/kDpiRS1rnfng0hEFEN
08MCWa6ea1qYIOI30qCIl0g93Nd2x1MdnjOq0xNPXG9SsKZVHoAx5mO//d0emJbfyNGMZ+eMXFQ+
lsu0o/z71EBSAYr5sY4psQ3/7RSMedLF0QLi4lAkTMSMw64zlHpcEIFWOLtQrjB9UkG8JwwMO64I
Z9jMfzKpmR+8P4UHeDcvq5rPtkR9zQJx2fo19a5ZRrIoiq2Cqb5k530MLrL+4PDoAwyXSSJ6FY0Q
d9bOyoBsyE7WP41ZIDnVPOu9s4LVlA40vkaXeGAxFeg8zHQlFFgLBzKVSuo0+fOZMxN9RUqOZzuG
RVWt3BC0jpvj4NmprNoLwvOQDYr4eJrNgx3lPmn5/GEmZV2u8KLvdB0ZteCOgnKchpvJhT6vkoSw
GtXFj92jhWgBMYlo5sBjppALC71ZRT+ZG/4PzJYQyI05VgAQxCfYSkpT4XcazPAt8BMdk/2gykUF
DjrYhHgEYbWTBloSvO/0h7Dx6MazDjA2XVZubEoEQGnjddK10/1rlGXxW4bFshqeXameCsY2IbYD
OOeNUzYI50BX+yo0ecyppFhCHKd0fjawSRiWQCwaIgOxoij6MR9UcmonuHDhhHer2E4GKo/3djcI
M7CbVoFyNBnu9Z8njGl7AMVi1dUthXbiB3lOMtEs7pDIE39VsGYV/bNZMtKIOhD72wibcjsWeCAR
IxMxE6I8lbOwMN2/gnFt4IW+kW3DE+sFtzxfdBKIC+kxq1k81hv5HGyXObJ6pBMyUBok9K6+jhhL
MX6+RSf0LSLOEnPyJdDOqbzpLt1YHpEtyVtz/D4oIJH0PLUmkgFjNM8yF4s7E/9CjvJUERz1+EQp
VGalQ0yIdb/lUzYJaLCalkKDjzu05bxTP5LTcxTn1ZUGx1rGMrfZtwCb7zBkmLQCD1uz87Vl8z3o
XrnsDSORLkvAgkFplvZwzL7Fo0xAwCxP7SwCB/ZK0p8FUR9Zsp49B6eBsE4M4qzRVtXodzSw2hNb
OrnfnfD2wMQwRnfRZ8Yvq9HzoIBzJJZ1aXl+CfVeG7yuj/zx1+3upmaKoIRw6ErEZu34exnykMV7
J4uhROlaXuFzVC2JLaJpf5k17XEe9sndIiREM2WMww0Tj5a1ovDQ/HPRiulflwJY3Ps5WxjIRvsg
R00+vgfK3cfkT2cVNXvBZzUUhq9Mm4NEsTQohf+qHY47O1zqom8WTD2dXKZslnQUVLrvNsBfk9ZQ
6fT5ONMcyhFIMP5u6AODtdEB6nZIxZIt9IJxBtRlcPFbjU3gf6dkQM8GP6+ZS58EpIk0styOWDbA
ng0kxEyqifsYJz3nCzPcWYREOTYtkl/IdHi1KNtk8+BeMhcm3CEyYD0fV4obdqI389sDLH4Fcp8I
ZmrzvJYPnPLnIz75KkEOV8mP/IrHVqTT1T5jJkXd4FE3qU9ysc+xO089vKHHQO1VRVl5ia31B9B6
m/I07sygXQAGa2uvGbvU+2aHcMO8/p04G1h6EdMaNOzyH40EEdS67h2EixNpoRLz5RXBVgGMXLVI
PR1f6Vx5+ItWX+TPv43reLYr3CIJcey//LTxvT42wC4TaZnD5fo/qsCHOEyAJKV3AHbs3RrTG71I
6k34ZNv4cRAM8xauhvfrwqJ46pPVrhDQ6rlTOjynRtgI3KAf/F6O1kTQhzBp457/JYrrgwX381d2
IsVMo9uQVY/DwjaDtiXlrSfWvf2I6v1coIPVCJTNQhjSE/2TOm6ILJm+78YovHUtewm+D1A/ELQ8
Q7EZxyRUcfuKn4gH+tJezmSGGJDZMkWCKOJ36s99XrFIYkdJz5JkTRC6WeZ+dg7aMfSgz7xS3vBW
yGSvbrMJgeaJFUPMaw3ClhGN+U8fFZJSOfJSEDBSWZZprUgkkXiBduJJ+LAeIMNM7vqmQ+KQ+bkj
6lKbm9ISkjFP8u1NqhWgHGeYWGCEF/j83ZedccCIWVDjzDj7qBVBYnbaU363iCmViu3Kt9HM+qDq
nFMFtU4aKfn1ORYiMEZxnLG7fg/zCjdivbjGj7R6Q6Z9ICSAa2www8m3epGp7PW3qibqaQRr8bhv
XD2L+1fiuoW+BRE366R3DczRuGGEHGjcXY9S5bcUu7NrrdfPAp7EL9wCxPs/PjwQe+eQblmMjUhs
p/8nESbvJbSJSQwWaPbjDByJNs7B6QragISB94ktxKifvfh8NN/eb33Tq8QrkBsVwMe7K94M6hqT
5qSWWIH+HNZc18pBXm/Glfd/rkKtP4jxAJEQ89NLVaIXbEyqoEQzzmc7AsIxGYwwf6hCqv2sGE6z
UaKATfdGNk6o4TRaNmyP+xE6IkF4bkqwcHKj8HQWcy6QZFBJILPDUR5i5YQt5/+xm9be8J39lD2z
nLYqB8XtiwUaIG2XhACiIAQ7Dh+31Mg4CSaNGaHZneq9J4L4ZdBFOQnyp/AAxp5R32gbSg6cQ3q+
ST+yHPkk7oVMhH6PPvmbw02TTwoNFwwhLYANb1VUjyzPIRTyS7swo88e7hWRgEL1kVPANuP98wEA
E74uNSLAy7gToEFqvA33kySEm+wJ5xsdCz3a5YvxbG+F5/aYLG+/QU0KgeF2kzYaEoeYDgIA+VCK
ZO59s3i0Li6xkffAvl7w8wVvXEgXWoC2jbFLn/WDezDAlbknphofH3BqNSszRDdLdf3Vdp9tK4Uk
+7MxSb4nruxlAjv19SgpB+3wrSyDi+ESX7gyUEEL5Kju2bSYQownoCmTHtiKnc7XbIiDz1NMqEcw
MK89ii8+FH9Bb1qMOU+gSwmvnKWTESDsAz+T4T+JbyOFU1AhJiCxPfYBK1ztEMqWNxkJpuWrVFOC
cdK/ezZDR7nbw6DP+oZWOkViEkEU1MYXoSoIjDGMeAuTd8RniQGo7/Vf86XRVvlMTYdeXchdJJJk
Cw04SlqweL+5gGdl1ZCHTFdY1eQ5sADT320mCtJPr+fsos0epeQF6C7uZg+zqEbJKMK0WXgGzGv4
HBNnfqgIN8EhKhgq2xBaKn11qp3C0OyzJ2sLKQQVAUmilMckOoZGV9365wcWLv2pK7X2UhbJheA8
pIOqMcXFBn8lByQU+KaqQJWg1AfSg/QS/TH9gpy6Hevm8LYnklBY4H7FYLvztwA2ltsUllUbagfH
up5sB0qEnj5xkTtm8kKB20MmbRcM00dVad6SZ2XkI73MGRak33ME+k+5cG/kUlFi+ADz8GSIzrI/
K14JDsGFCXePWrV/v2hO4cx6KQ3hEaudfRKFutgeIUOoWfSV31erMYOyCa+YfYESo+xLOKRllyrp
E5ZUjEJrsNkNapwohK3EVl/sVW+ynoAZgIqfQBTNGvzrCr1N7OTFWLp95kH8nU1tYvCFIj7DAiId
8wbi0dSglj6zDBFWViKl18Sw8myADH29Xc/XJUDgOMDOwC7paTNqWrkSacJeZwwklbJ/muPMp8Hv
VwNBWCqQHsNX1jObYt4p4iSdphEp8G/zLWuJK9lTKA7LAOVOzZaPo+3euQWKoC6vSNuOPTe1eHj7
ND4Hpjib0o4gvrRZFQTzdeOtKcUeR0u1SizEvor0n5PZ1i+o5GHyU4jiMbD4T5vlQWsH2W7LHZ+Q
606Ha4dK6nNgxq819YBvmTUnbrW7RRgzYMj45f0imhL7SF9q+JArcAMBPn8NY99YqX4RQ3xcLsob
4vWAYk1dGWixrjIyJhCRgN5DiRjL10r8XiYMoH93a7T0Yar39j5D2pLGdNx3qxGcGdmujv3em8Zv
lfNTQZVGxhlXhEciKuA1bycpWSv5Ibi7N3QxXc/atwqvXT6O7dwnA9e75jplSHnEPDaxZwDQ5utF
uz237Oixksi1q0E0nTxZZAUnnxX5PXug+Vx5kNX8esLEtoyysKslnjNcNZRu/Im9gx/O3GbfZ4dk
zZXbUf2YNqogP+yKrlMlP+UeeLho5Rqrt9loMdHly7mcKlSc0R4Ow2XKyLHatNmZXMmFDiSxJReL
cckD22dN/WjxUizK4m+ym6jd6/UwWSsgv9Tmjps7L8RmXiigwD8jYGfK1/DLZ6YpGGEN4ud63B8n
tBRP1PPJw3kY1XFRbWtKA2YS428kRWJGFYWoRYutEnICBSDEIdvV1dnnFBLimyWoeEcLpgbOlzeE
F2mkvk4RpgYiibTlVZsSjkLXWE4MX/OeVuehq+sIqLNM6252xHZB846dXIN1gQKBzbYeaMNCWH5r
D92PVGKtscsRJxDUeTb0FE0nCah0ThWp+tPO0STw1YTRKXvlwajY/eY7FxB5YNPD/b5yhr6ovZYW
TG6sdjb4lZ1R1QIo4GQyq5b+Hs2xy/9MTXtNibce18eI9rMSDV/eB87dW46kbdlnljXFzos67hMh
YC/AM90Kwf+mWV1TelqcebGcVKCvTaQ0FWk63LKY02B1HSkUdJWLvNZXW1QJtK13SFBqNFVo3xUz
cqA6lPLFGkvmcf0qp8tKAO0gMNY8mgngims+/CDQMHuwWBpYbgcGQcfNI3OR7j9q15WViMDqB1Xv
qLyCf0vvbnnnlnJ7edIoovirLySkaWJzMeMNQz05iSA/XX3toAwW4akmD+RjSXrubp2nl+B334jR
TJG95p/75OQiCRQh2QP7y7+rMEL2SXSnhquV+btLoSIGNS5zeqY8U3WBbNEWhXDHED5A+8hQca6P
X2b5Qhh425zqw5SNgIhWH41fckJalzDVy0T9Eh0hhYXW6vKdLMxfLmcjiniItBmrznUbKJLMZi+5
FAFft/bos/XSG/lu6T0bxUc+FW8N/RzRn7d9Nmb6YmdrrIyEmqtlpgW//oPSeLyX84OQK7y3fF4k
LOGOWXon8FhIBWx2gvrGbuZ5YtICRU92WdTGyFjq6DoWs45TyeE14CKR+7gyuOTXfe1kVJe0rEOT
X6q4OxQF0kkJlLZLjryfea6yT7re7dHc/OrNspoDohjq3HaBV29/lJ4zrLIf/b45fFt0Lsh+24RX
3aNBaqaqjR3onKqniUZDXV7kiqP9kzbs3YGyMKWrGbP71/RlyEYav8YK+oineuHBCu81K8EDXvjG
u9o1N8CEuqicBLbIZ2G+V8va5TB8O4LaEtgcn8oBeOS8z8/O6/iNadhOm3KXNkik68mYkfEne+qM
GT+5EV8hYCEZc59JCevUlig2qRjvA1mMHSsBXaL0YP7JL/cJejHYa9f3Ne3S8mB4rORCzq+L/eSy
8yxE5sckkcZmEkYFX3nBaWnY+Bs1iQsYOPA2W+o1su7ube4oEWVZuuQBmS2s+JE0WIA/ujMeQgXR
ianE/zv4cegOhXKLge7vU94shQordjQJ0QCwusjQV9SZew5sw5T+RfhqbVU6mzjOozpGUUqdwJSV
QkHgCG3B36UDJtoZYbBjWLKCQ76iBddfMfPkN8b+mYwWjko76l7V5HN1TRNMwUyCBipgVzFRm5Lj
H6E+4ZPzskaFT+wZ++K1CbCkpQosL49aykCHUT+cgz/Ns+Ue92TEPm4dnR0x8vC3CYJ/9UHrpN8m
E/NRlXtjiRYHE664iTze/hPsZpFHZwskXRx1w/iqIigOlThUxX9KWJQ70pLZVc79cp11LTdFGQe3
sxwtM6MBZZn/0YS2xeHDBOjzQK688rITK1JOC8UeyjoZUSLcSLau6y286c8WuOYZNiIRI833nfKz
p+HX5hxjJWjkHR2L6XJh3U78oYR+7uVUJsp7Hk2O/LWoCqUf8GpUdOCAhvjwjBiUoQdaEZ8O2VpL
40pbCtObdIRlP3Ag1HzE5knghPpLM0lgsiBfOxhdOg087FeRfvE/MbfpZAET5mV4CHjwXHwaYTdE
Wnen6ElYyihum8dDUb5GxND1dHmqFl7DQ7+NbqKS0VdYFovbcyFzKu/8SyPwVJPnbDb42r5m0yWH
HItb2gEQiNzSQZ0wct1G8+7jRTEQ0gmgvLTwwne6yvEVi5dz9SImuy40NqWsAtfXC6ZJ1DWyLHCu
i3JgRiDHTlAtS2KI0CqzCJ1h3UuEfGPoxla6tCxbUZ9+8x8TmafcaHmQyAu/5+6uaaGd5JyvX8IP
bqACDiYDp/1GUI+o/VaxbgXIf+JWbWoYqpke2rE3GMqhZkxy4j/uP7eL4tmGIsvFVMuFXMNqPcMs
3NyDlFWPXDMMBXA3iT7fV/eBHesdKn5pwImKuHMFNV7yd0lt+DFbCGkrrDr1huLn+k1bLG98j7Oi
xpW3ufwC1huzknxlnVDg1bpmEptB5G8pcvCXkfldAomNbVo9ZNU29ZYG34tNX2BZ9kJ7uKvSD5GR
wGD4zu3BLarYAoiy6HkaIvtRq7m4Li0cv7R7Mko+Q7kV53TT8J//owNytLFSPANA4TMgB+jDRzrT
EHwruzWn3cTCHMJ8TA357HFVWCIhY1AArHHqsuKMsBRX2lCpr+0mnZbzMam1j+3ZZSyqXwPzgYar
WcBebz4YpI2msOOdGrnqH0PW5l3GB+7AqDKu5eq+JcTsVjMh13yx8ZhEJKfdQLrqdUIjOGmdipi+
MZwDENCJj4Ng9wprfLKniHSdFLV8ZVh2YWPa2SxzUBAD342DUJGWJ3g0LXdUTwpv8wCyXDV59DDN
zzFrtYRsEUpzmr4jFNpmgwnblOcpmiNBy/uRcnSz4iw4h6gAYXJoyuooFskSGSMdz8JHRiEG/GJI
k6ucryPU2cYQt829Z3w8vroNBIrIlDEWXvVWEXfn9QtweVfDfCbs9ZbdCaPm6idjpaI5tJmIttdI
TEvUJn8Q8vo/uejDYCP8vN52SrInIa42nLta2/0fMu34MKQB3j4yIPamZOgaIO2e2k6VhaILFoMa
9ZdJbjMvwT/VlSel3HytVeK415Bdb85eIlcpcXMpAVtAmRoruGUiw7EwjM+bZkyO8vNLrmXgNglH
bKih1VXBC9FXO2mHFv4cZ02Qru6RnEsD8nChDta8WiZZJ3qD7GTQufQfDChelsQKAGlAVmGMp2vN
EoFjnVIop5NNlP9cVUFrk5RBSsGI6H4dPVAT2EudDfmNE5FRcarn0rOsa8czGFWr0MB6RFv0nrQj
A5tPCQnyfIZXoJ4E1xa7QaOa15zsDUluipWLzXJ49bSJ+59EphdoFP2TLX6rd0jnl1hnqHhS7owt
0a4Fh2Sdsj22xXvCZlSLvps1/XRu0uhxB3hxvE5Wf8Svw48SKSk27b/4v5z1pcCmnR4CS4CAbI+S
umxiAK3eNSrwt9H7tZtE4S5pbdxQln6tEArukgLgVbDegW7LLOAEJb3LYGo/GFjXLDAc7e5O1Al3
T72z02uCWEK5vHFikvCrEYKtSv7wdMMqzb8y+ChcLykO2uPuCizdALeWGUfeNoK+9Kj0rFFmJAtH
2icPSOpaWy7ZbZhHtfYytNBWXffOdwBgyTgDSNzgqt76Q9uNVQ+sCHFk1joPuluJZH1aaoj9rwBV
IPvMK01aDuZGNEu7NbjGi/EnUtouKHe3olGFJUolj8AxgJj3I+x9E+IxuScPNNsXdvqiBLBo/Lfm
OY/OK7Y12y81hsDlg45eaaQRl8p7cxB8pXe2wIQd9SPk5uttD57cayjUTFybB+I2VL+v1y0dIFfK
lQXjQ0IumeMFr4RcG52DD9QFQLwcgqvwviPUUNvllTBgUhKos2hN6s1DnzK3Dh2cIbKMNwVPRDQM
WOP4Q1uEh/13m+mUwbJBPF2svAqjH+4LgufdtnEraUJWKkzKbNa+bil3sqbd7IQA2+I7om4eQJ9n
aYOlL7GI/jDUALWf1OuC5bMpWRJ8MtEnSOD4e+MjFItbtGXv1jq7PLK/avThlPrWW46BzeB6sU/M
pfNMtfMI6cDm/9ueZcJHZIFrol5TcMdWnYj3xIdfXeUQvyJ2u41Z/mi2rL8YpiraMP85aHzJ7Atd
DNYjSE08unvxYmiRzbMAqL1buiVMQgeTivDRsq5qklXaOabeABjnObJbJyMSoWW+MB+roQCaGD36
tG8AwsPvfrQwPdOVLJV4PB8d/yDbvfrx4JujHhm6VDB+DRSdwWx4ayVRucbPJKJRWCQ39Rd4Huef
ypPTlznYmlPThVxVm+rJxxLsIXnv1cicQ7GlaHY9SxhwiVw940bsLqax0SXXxUcFbbqVS1F3v9G9
sUfFSJZL7coaGo9TzESwNg7QW9XSnSvuyfMhyUVvmpO2/f7sdhV84ozB2EzwoviH++XuVluFHUwx
lEBBVA4Prr4DSsLeNvHblfjXLyZFqsbWjHXmJPAodjTML09QS2jUa064aPOyZY1erZIOr4SiZF9T
k1MMaKsAA3qgUZvR2SmZzEs2LSsPtRQrTaGWxAQBF17Ci9eMPNrQSyts0OwONGNYngmImNWfz6Ex
5Sp18eXo2B7LvhdQK3eoP48YzbBW2D+Kk2KgYzMUETiNYd7j1/IeH6jHD4rWmZK73EXVNuXQTmA8
pthPYNf47UvCZNjUqvLcd3vTJrIwDRYlx3mb3QtYWrMar3auchP/Rr5bV9vfLWQ/b5Hhl0RcdqRT
Q/QZEqjZEo/nIBEAUGTUcd+Uij4Uf90BuFNtnlWKzmcjvSJrvJl2HKOdJ+fvKW3l7YqbHsY/DWHu
lRs0Ke+ipd1dlknyBWxCbT0MIC0fYfiB5FpKZx1MSKbpV9MbX0+1vwASxO2U8NIrbNnRukr90ZjJ
KQvSu38gDSb575in1h1npf86TeeW7mZZ5cOWRRHhx3yqTilHyvOEHoUxJiaT3LOhkAxrHPv/lFwE
lQAkIWeBqLu3darlgQgPiZxQ5ZFKOVf33KktW6wxYN9t1CJQyuO0z3/gYKOlxQv8fZFRcLW+2VMc
10BOloa2fsXYf8D8xCJlj+t7FBvTRkABva8rS9pbTV4+UOHcK8KnN2lhSz2Mzv7KNYaajBm1qpEu
Hk+CpxFwHKW+2aJHJpbsJBh8w5JjUVj9yXaoqaU+LJEZEwiHGMfSVjn4JW0KVUSJJ/+EaFGMPzUA
AvOf1WAcCaimwKe/dNpfKndGzV+/DxTmh+aAw41yEj4MAIPsTTTyLJLZM/wEpgDSQfUnktU1FHWA
bM4TH5bkXxzWGRC6jMklPakj5fTxSwCik9ECYC/kjCPqY5/GnzHOUujvdB/COxJnawPM83gxfNwb
uk4Z592GsWfBLTEQ8Lg3jI8+g61dyOng9wlpIjqvVl/KKQ9ZtTz87E3acDcy+iW66E6k6kjxyZae
nWj5ns7N1Cp6kIjtsat2AHiy5TAOFPFccZnYjKgehYAXjAkIIPT508TFAllIfiFIgsOMNb2oscYO
JmIieg9VE0F2SgmMX4FaTSsxmyYwHgi2P4NhFaSvYOWgglJJHZUAzFb1AkIA5HFu7WuCOGunZVyW
nx8EWVduG2pkNTQ1X/FkirrASGGcuMGA2NuVp5WgYzk+3Hde13FUhXRMaeRlTyXMdvsQXzlzHG2f
y/NVPIZ/hDMxHu4SsRPRVD85RJ3QTGo4PBswRga+IXxGzHNFaLl70lP7kO3UtjbgpzEw21bcYlzy
/GqPRRtTS9nEN0SUwP0GlUmlIJ4JvG3fhS0DSdvzi8cLDAjlLZL1gztxlURiOxWoBTQ9c9RV44iw
pRWnDOzpHdYJCd+JFHWLxalaQzhI51vzjTYqn/QpPgEQLasCPdKYS/mo11fFzekk7vRf+2Vby6kk
UAoyrYtFB+F2h+BZ7JDUFqG6ZUbFcSmGJKsyUNsef0BqYUu/IjlIGW+z9U2sKdpRZOnYQ0OZVIEu
UBP1MMeQQ6K/VV6VJJw1Tv0ZdFsfIOg3Xzr0REnSdU/gppUrFfXR61Xad2b+Psz8CexVK4Z7Qh1c
DgqNxUpYIPCsPSVMYyP3QpaJN5mKXhphhinkE3aPo7nDjSJxIvlklv0AoEfa3+aNAj0ohJh1H+iM
93BWoaD0Pjs+xei3o56ZGASIPuyIOst+OD4BgLxWcMULipt+Mn7TNkNtGpWcAIbhMSjjWoFvNU9q
yLdSI2C1DEW24FQcLWRY4J0UyanjWPxIXJEtZJUJeK7G0WzhyLwzdA3/7TaImIaBcCXBBTXMaZqc
3M+AWe9tS6cwCtaUVKEzB+2M6ji0YguBFWlVp2inVEqiCtTUD50XWHfZmj3UYWvQ6hgI5hTVwzRp
GlbmwFdxUqAV12sUCR0et8YdSevvSk+SBX5qFEiFC3hqzSIoNM5TRZBhg7PBYHdLqyBfkLAr9Tx/
7zqkFfOc8wtoc0yDSQ+cI2KwmzmoTgfNvobQkCo+ImbjHMkmENjZGb48cpSsWB7lzwULpbyyZkr6
eYzBXveeW3MsWgEyFuOjgsSi0kvG2XvpKpL9wjETxeJbJu2QI7WYzWzsyEQGjylZZOjpxxsKfDy+
K3GHF5B4o9zN5pCg0jqUusSMAezmHiCg/8Udip9KXlng5HusIf0Huc03rrFi2XGcJO118nWrQSZU
z4YuPqxl3Ycc4i0OcKF30ThtK/WMyIo9qhhXA47HcYM6mh7Oy/gv2bhbgR6S5HVZqpbv4caz4GY3
8AjxVBLl8NEYFt3i+xpBhalO8V3cdZvlooyvj0Z/lBU7hs+vzHKplX2BInUPbhrdzg6D58Din7/H
OUzDKp3hkh/u+j/6aI8SsUs0T3CwMq5mRWDQEFkVJscVvkDuUCYFyqilEchw74++ekmav1LsueS7
SXWg7xlpyXihQ115NnlWTYKbVeJJpZ4gh/CHClD8OA012cP696TtqkLBziG9VZci+poABcxXMMeW
GSp7TnzzWkHWNudYSHHSaVcwa3lCTA3RxdTVBsqdMARhBx6yIQuskydaRXY2PC73jZo3o3AVNMzh
foiXwstixz1rlI7nSHLHZ3ge8rFr0kYou0OET7tjPb9SIxm6MjJ2mw5TLhsbZK2h8hanb0NxCShl
Fx4i/H3shtbWE9zZ2JUE656LK2Yb1zOqLz1ey2/wRXoXV4Zgu8kFShbFYcM4UkYjxAaZ82MViQC8
pvxTebVu3LpeGaszJAmXLxZElfgGu5QkhBpK4Ox2ssGgAMvorertQ4rX+41Bkedmeumv4zSsvhh9
zvAHU5W24/etgPmwyR780rQMZSGV0Vbzzs7pPJp/99KV92sYnvIGtsjmuPR6JXKpIBWf6hHLmESj
9gpQUe4WjKY/OkCdmblim5u/EJbMhk25bqRpsgPByLu1Kknm6K3CnPHkv2NYYTSPnULHNG8w2MeY
ej5ICPXhbP5ShvuxMbKcbOSDWbQuEWaduAHb8krVTXQ/dcW8X1OoCH0XFnCbcU1dKyz2cuGGIiA0
VIASult6MK8irUwatrNeUIrpFDcyTI8EKzUrJwpvqGFjk7cyhtWHyZJtcRe+i4bln/f/iIfeJk2A
VPvArXk8po5z8/ltxU0pgHHbLz4tAq6i7MDAEKhggr9R5pB1gK9XKLSTLZjdR1qJ9o7uejpupD2K
LXZyy63Xsh/k5qOfDVRAfN3ARm7lGWK9Ryu4ErVWW6t4Ivnhhw3uktN1dJFiINtR4+hRL7wO2QVd
eI9rbbGW/9rshFQsKb7QHLiGO+3ljsB7KoD6gpNvzB9F5Hmp8Q9eOsfaif8Z3PbMiDJZMQBvajdn
gxqylNwz5JFFemyqI8BviimheG5m0K1Wh3GaPMEper8Ov7KR9zhfwRkZF5KHhfsURAyqedAcE9c0
9OXkpBpMmf2rtiOh+nZJvBptNFs6gVxOKWJjYWOUIFFZIDGG1zKweJBNjyDw+wmYnoT96PDhbVmL
EMr3JJljdwgvCHsKtp3YjItWzCbS9HgRxNF8X9MFbJGxm2MwOLLUvALFwppzj/BmlJz9gdX6JKmA
yqIy7+GvAwdWBPecLsap41kywpUdDYvUZgLrETEBOAxOuMR1dJVIU9LTJ1rutAXwnIpDY6+ezn8T
LTsyX181nDIx2pvJzhfTtrqo7TAEP1wAyxOVtTRUN5LqK5cH7VIDqvhI3+y6BSfHT7HAvvJ6AJUp
LF6V68reGrPJX7JklywMxQe1cjQtgoTuaZJgJThU8q/QQ0VEbw0MdPHbinhr03/lCkqrto/tlcuS
CGpnigybUSn+4Ww5v6e+4ASIUaJIHb/EtqAJliCIZX+E5lIVIE3YrMfq1GkrJsJ6Iwhfly3ZlIWw
A+biFQL6RLV4lrG36Qq6cBJyLdHrRrsaiY0obx4t8F4fLwqFq7vggXsdF7+grEOJRsoX2ZAPqrQE
pfRVb+15MogeaFEVlPSFo2j1lBWzgMv+lSNraw/wHHwgClpeeBTB/8TrhZ8yswKrF7XwNug+1Qh0
4S/mt8bUqED7lINYT39DHQZ5d4e3udEOx8MRxqkdJbga4ZQrqkfeHWZB7regoOAHfPszlXTKz+U+
RLJDuN42rpMo1/TTjrC4rtKVFW5KVUfPf0LXjhT+MPAYdTyhheu3VKOzTFW+9wO5dmRuK0dOXtYv
Lg67z44pUxgpCdkWFsFdyFLuIXp6ptc6ApMKQqQeO+WI7nhCIHpsmnAa/mPAV3srpKdhFRx1lKIB
fWPDNhnNufMjbV4bmondgOAFxc5+cNIj7KcrjVWnT+yChaexo3CIbFfrsqqJt5uGp+nB1yFVFzB/
JLgH7ZLLEWMJb1C8q/siuNylzchyN4qQcqxwqtyogCNPMZw7KVF+OCAgnmwjrO72Otn3yhRKFjy0
w/RtDlpngLjx5TQ9rqp4Y8UYHHUYJlQwBV1DI86EGgWJoAfQfHOLqkIAbT8Q7x+0099x56Oonp7q
eeclYDal9kVqfHoC5Yyl/7t1SnZLJGVRT368V+/StNodQq87lIkWNiHpdVDQRIQ8hy5aj3pkbOfR
7btslffituLrxbQnmmsPknbViWC/Qx+ADWc6p3keua2Os+s3L1ypK6UkNnieBpi1dQZPv5yuEf5s
OfUlrCQStpVLaxkl61kUreNimmLXpwbyaUoqXevb4h9zho5E3SFgtiu1RFk01COw+2CAz0XR7SZy
7TI0T3BRVfpMmiRQ/t+dFD2iwF+fNvg3rN+/1Yiy9Pnbd1b1iGwANREAYqfBKdTrv50ECmIcB4Mz
X8PCNJHYSwer6Ba6z8H9gfESQXJQwscl0fgokUPfllSDMYJSSAM+BFHTzmD3Gq0LINvpSQZO2Rij
YdxC2Qbq0M37hXpBdRgbya7P/cNDr3e2X3hEakc70z0DC/vH6zzi31SkwZNLtWDEMhOOln7JlInr
x2Z9B1xZLoxxOZPQh7kP2Tsvcg8BBgZEUk8WQzVI3l5S+0C0A77ngsF8BBDLMVC+5uLKtTOXu31g
eSoIk6COApZueT/f0t0F2s9biSsfQfCeTFCJZEsh+6PdZdi8cfbbwdR3lAZOgDtGrNXTPjXYjWqF
1lfeIHsgQ+h/cjGtFsZMCQzfMP+i0asFEwZNfTRgXsbR4QAQ7WtsyRbODRxeJR2i2RdOYoObCFEG
D+lEQvGmQVLOINrJ/+Df8Ao6Ly2zNh94njRWOpJMCnhpH7QWOHrrVwJz7mwCrlkNcTX6DOX9ykNy
TXL/LNY3KQYp2ehrMjtBUgQdB00PeMqns5XgmRop/h84902EB/qbDhNinzNtKTBDPpT+wbYzn7Wf
UAqncwOycrSgfiUQ2SlgxMEChn9KgHz6u7ZLUQB1dhD348MFpuV0sOX77fsb+aLFOND8m9oQom0A
PaA70aGi87VyhhS541gwcXrb1kOTAgYe2oIcMbV/lf0wiX7V/JKccS4k93/q0RSzOfobzs81jfj3
rcOSMly4ghSsQKRHwPorUIu/5zzHuEWPO+BX186Er0HzdulsnD/FVLMMjoU5fB4DFWr2XMS5WWN6
5Cjhj/U4eeT5x9O2ADTWOaTTtNW3605tVFeyt1xuyQ5P+sq7+9W11pJc1nrYuxQdmte39Uwu1Z1Y
J0kTfAkU3IoF13huj0MGSx3//zopHu3Hzczp0GSp1XYHZHh7j7blQgbd9HLhrYxUHwwEr+7s8JQQ
TsM/gcUOOMlVBtuxO+okvQSlPdz45Z6IqBjyHagvsBYMl8fB6j/GAH/+rGTX9aItl4ykTCGzLvV7
L5AdqxgiwuMU5ymGvCW2wpYPCQRxjQijfv8P0JAr/vJjg4jtjw6LjsvXeP33iwjx3x+nduV2Iwz5
pGFVgNxklSylEQstlttpLIXChJDcxl7ItM9mtgPNBVDzj4ZYbxP2a8H/A9sNPVTYXuVWWYWo3e1J
fnByfuC67Gp76MpfSiktY0ovQj+IyWfoEQ5OCcFaccKMMa7EHCgLlzocAbNA3nOf3LuSSMYicgRl
adC9CAg/eFTDoirIGWRHhfjJhbNKt5GIfFl8rpBUVWtjnMk3ZUMlA/SDv/dc3k753AtK23IX+n2Z
4arD9WOQJXqkJ8FJOJtqbGeZiNKpa4LE9sgJn+PTFBJ1OvlyWt4EFPkfuP/auu8Jv8IuTKSl8iTa
/ZgDEJrA2XCeLM4Zl9jG3gvcBltMRKgJAdtEczdjYFdABMl8hAFIf0Jm0AuurWV91lf3HXoshTyK
NYwdBcpZTR5aIHPRsqVSseZHXba9iWfYUhpWEX5UDpx9/Lk5qo0MrSMm16UfEJb6yTISiE0434Rb
fu5ByEFfHjUV3o0Fo5qnQESLJl7Uv1Me/JQxS2NVCEjELuI/piBFFLFN4gHPvvQWSXEEkihGiJdQ
x/b1n4nOiDftk1NHorR36Xg2zsEkzJyFJX4f6JHOydArGsXiOr/ZLopwwQCb7CqZNPC4hBhp8e7Y
9oUVe7Rz+RGRYMyUffn+e4396GhW8c89vKFAzsf+tWeLkiBzZQK5WMJPtr6ZfohItzjFizwPotJX
slPMt7PHcVAK02LB3Z93Ksy0OoVyB9xxrEmeb9mzoEztZAVG85fLMqsWGUWF2tv3hn8+rAwyuDu5
453Ov4DpSFIQ/fDbKwvJaAJntN1HmAfxNzeBLTqNKZ7EjMDnzqzD+R93eWGQTYZQiGKOk63nakyR
4VL78hrtJTxIs6qGK8j+OAB1dvwgYEL3qn80Wug6sx451I6ISvUQ8EKJEKnvhrlLuvLzI91cqg3m
w3+n0tUiHNTfzRS71PCre1ySLvD7XtVbb1ntG830TDz8IRA9dFXC5M3MtT+ezfCcHuyNfAMz+5AN
sUb5Un+CfnbQtk9hCeOHfr3AjKFQXqD+6i1ECXp3uFudVmcQyv9rdAGVL0v8r89Hx0R3CFEOhyFN
BeFygCY3OMVaUC8I5XhDePkMQfZ864BMTvv6gnTTkXQvgKsmleJfTOUeG0tPBdmq7sW31LJEw3wz
QvFvYk1P7ttcLawp6CHwm8VTW14mQHGTL6MLf788Sh5sXDBUSNKks1ycUq0QwBggY1mQ97n2KXD4
s00BG2XJPylmjQSLkQy4lBClPma0f6zBbpphZHGaQWWfpwbrWmQBNmOnhiOpnlLDNeN0Dnah/bia
tb/xRcG9iNVZgS2+BY5bbI5vDdCQ0eVWTyTeaXe++D9Uk6+hjFQ4VlZXG2PQ/kMsGKGhgUAk9Tjx
K0/GNk7Qi5FyBeyR/TlptPr+/hYF/zhsGiwklYhf07ZovhpW0+rWjXCl/KzQ5LpW1Q4jHN5eLvRQ
nFiuRTYwf1Wthyf3l+y8gpqn4T7uunsSEyQmkgL0o3YdF/bgHBRxiUiV9c/ZbI3atg4bh1jjbH2b
2UUFbdXDVWiQmoi0T3n4PTdlFuAUQh9MYsXYSmTw8pcvO2BTxvy1Bjah+qLJdN20Xh9REeY3MJ4f
I+sdxOG0ak/756xsAwSf43EjBoaaGQC1GeZQ3JQktffH9Rk+er0ghpYM1f6esGf5DkEWl0B/GTQ5
qxmD302vm5zEoZyPTnUTLy7+PpDJgL3wbPfFlw9qh6kp3l3GtO8pOWgrz7o+9zqnD5tkqPDxftHK
YXX23PRV5Auiyv4H5iXGJan4ysr4zfMEIyg7Lt20aV6eGsY8lMjzhKFuDQbZUeyXi/USIXvXHYDV
wi1gS77tgKvnMmrQNJjMA8GL8j6fBMr8+Hzs6vpGxNE/O65RIwoyLcfVkK6FkgFmqzPw+wf8NPMk
Wo5TI6dspFZCzWoso49S9KqkTgPdTo5i2dQKFmtxpcG+mz3i50wHlqrZmiozud4Seff9SbZyvpDX
3v4iu8sn7IKunHJVasjTrJEbEWPPIKN3+4KWuxLA5V9HbGS4umjOjAYCi78/j94fGBSdJrN9VYxX
S+XR8WwQirilZDHfhBZVrDhPQxpIdovSvwyr/x0oUbI16Vi5cWOcgJ3RPwYLr1fkeGt4yjts0n5R
n8Vlu/lUq2sOQWDVc9/zRm8P8/d7jjhotd3UgZji4yoK7bndwdf9Dn38jiNKDA/iFs0IRbM7fAgk
yBdXp6a0gP0/5e4EpSDaEo0P6GYf/ByuNaYKx132C88hd1QUG5cAvY1wW8Hau+Gn4W8fTwAJwfqH
tSbUmDIWK6nUAGQ3YpKn86uzajBXUcg30nnr3Yk6fCtW+jUflaOhyc7YtCvAA+c35CCTKy0yUdiH
sa+wHGGba76Lezff55Gh5Qhth4kusQLqNhUhdrkQgpymOP6+G2V17lmfyUDfH82LuTzB58Wd58GF
VMbMi4lQlowtpC6VTx3X32UwbKGwHsY3RQVNCtdz/h1c6ix3oySjnWAn7QMN+MTmQp/rpNi9AtDR
ackUGXzmoBh6RgGdno6oN1Go5+5QHpMw9MMAFvVGlDl1o8fDdjuoHQPcFBceGovPwZP8n+Q8e5Py
MbccplslK8D0bsSFG9EP+GTPERaeUVuSuQT0KqgvD9i9vY9UNve+iabTTZ53rD3Jk5Cf8QzMHvLl
5xTow9rr1zfEdAE4kPF4UJZaPH0IW2a0BcJX5WrUBuiX/Xh3q5sixoPjXXHLiqxs+atkpp5JpgYb
iiNKj62W4Z67GovGzwt7lqrHH7FZInIephuhhYBqU4lV5jC9N4RoMlFA9LCDx8fXY6DHwbNFzkxc
a3/viFx52fk5JA05j2nqEfIhUDXZLGAwCFWoEuOXOBWwMjRDRSLuDlsbuZu4CUridwFdDb5ozGUd
RoaLalupB8fszmgrF59OMmfWP7WJIiE3tW14s/drOpy8Z2flcKn4PwNh0Kb9cwjCPVknsEn7Svmz
jGMQ/7GUPGr/vGbVtgPKsSQZMhlEE17wD+pGXreLrcoFrTZo4Q3nxRnSKKOps5Z5DoqSEZl0u0lf
Yz7aMKm6sdOdTkOnuz9sV+7FgaKcM6iGmR7+CdNU4/E6HWxhS0t7fWw4inePEe9i/j/M8sm9M1oB
UwgIBKPyyVusJs4By36Q6SXvm+zdE6nGpDOKQ4/dncTByWp/cwQW4WFnXjFK/h7mnCarLvf/o+Q9
HsMmHvZiQaVMmiRgkVg6pv/6Z7HtOW8p4Ic88GOyv4W2c5VT4HV6HiD3C2eBmjlEKbzJwGRaeFG4
4S/ndhiONJqRDK00B27jSGgCTVOP5eDujj+xAlW8+eI0vpVLfh2pOwtnY/NUZcQrky7DHEhfYnDu
O55Tgm2eFH+bcA9a0VJFKXGRm+HlrbFRj9Ylr5uZHfYmVznjVidFioSWe9NtiFzcFrO6S+xrFjYn
ac+FvpCY8lPiiVQv7UsrWPttMbbqLETRUzB7qzS3OgkIgFdUmy5JQ/9EUsbzm7NJOUuZX/Z2BkX2
QfAgmsuxT8IXZgDQaOppgyuKCtTIZjB/FCeVw/UTArCLAEFdCoQlam8VhVTnnMb/KbALJKwdrWJ1
9XmHtd2CpGk3R0Ul8w9T+d9UrFyy5pNEdx1n4GKFatID8tjbGjobX+MekgrdtIQ0Syb8UfSWdITH
NxYAuvgzFbKDdUPuEsmMnB4r9HlsJUUUOSOOcI/R0yWWofxKn3lcgsODSRO1Ft112ZxFygfLluNf
XGZgwPY8c/aTiwcR1+aaA2URGa53pWG4wiaPAuELaNCfZRwr0+eTRfobZcOzKnJOqgy5aMYVFhw2
y55krUNYAUSw+bbTLeQcBvwpgFvrjYHgdI+U8KREYRocQPt5Sy7IE5WASt6TUpkdgtZRyAGnynUQ
t5awSxZxv7Y2YhNP4Em1vvIz9QxGVBco9qvYwjf7yZYkFEYb1MhJ1o/wKEXaV4H0ressdQk9Skgj
6m1lJjmZDbV17NrxSAPUegUr70W4KMPQh0KuT5bB3kw2s22FW3XsE2YMi/xtPR/XVhoT56gx2Nc9
0IxzYU9RtYNMD33t5gxAhiaZec5g1jB5AZv1Warudlh05f3wFm0RMRSxiAfzx0RwyNbeedadWhQE
TwSgtsJNFatph33V80OVJ0HopqLvY/X8B/uSQm1eH9tDYiRGL9Y3211SUQMNi1LuJqEMW0aTwnW/
9OV7YMUph4R4gkSAGHu53OYW3JnYewqOSME/aOAiREnvp67t/cnsYSaJqStlkeeTFNQ5wOhmtr5K
3YdlOljVBdry8vbaJ8I3bAxGOR+UmYUcbkByOVEKnIyVYh9aFYhIoXUTP1fo+sXkvF+RYgYdHkWe
XevsJNGXe4/AGNm14XYtj2sJKFfj8D3K9nJcp18s5flh4aZvS2+TXVFqeMHo6jmxzh7aaGCgafv7
PYe5iSFztA9VD+PsAnrCdfFz9hnqZZNo7XxgCmgYGNjW0iNInhZLXeppjgYjTBkudADarfwutsyW
wpdF0ElUAqzEDiUWdhis70MBm8tnYJEJP9znyHVDwMeeMQH5iAkgnWOJgtWdnLOI55Lcpl6ibv2h
0K1Z5pnK32o8vG7XDRoIOmi0EM3O0fecJJyKw5qj1CTOmGlrKIWeS6X54YcbMwf6N6RsSrx02zrP
Cz/x8y9z8HfvHOi5AffX5g4a1CCKmx3CFBeteTmQLWI9nQirMGW/+OljKQAjYoUPPfnD/GIdY+dO
JvILw7lHU6JgbarW1H/eE8cyS3hKsT2Uxs33BrgMyiLcdyY2VXwF9MGJE9I8I22RV+kJZY8Whxqt
2LgnLeEmKx0mQo+j/ooAr4Gi0Qdxs44oNZuRcGnIlZfPqDwDLGpGtWJ23++bYzrLJerYWDkXh4dB
Gbsi9qRYg4GfScFL+kxUVxFHFSNTfOoQF0wSb33YQjATiH1GTkDkCqT8RNjZ9R4wK0s9pMcF33qH
WvjKy8SFD1xNSvEBqcGE1v96BiP03oJoxhvHXFUsf4MO/dYqeZDH3W2wMs7QvpH+YOS/Q0dQ6V96
6rKa55CtwFcJANikDDo4XNyvus+PWo/BfA4K4XoUQtkXB+YO8rIlICMaEj0ad5OPfPzmLQ9UXhDt
IZ0ENeR3aBb40NfA9M9SNYM22hHN1mLgZxHnOW5QqzMwmil9Pr7zSuLj2b4x37rFWQHYnEsW0lUE
8dqG2YXhyttXAyJPqBARrLvOMCclkMkNNsjI0hXs/crmMxo/+F6u0lN0kKcMW2rV3glKnqWf0rLB
smiyR5V63ZbLGMBDoBI7yMin/lYSVPa7wsdajvDzxKpMSpgqEALWIaktgW+VmBVfnAPClGfaAyi9
rRKh0FOr8iA+5SdNYqyaOFyLv3MWyuautU/Ctnko1nKJ9hXj0WJwndppRBn10IZ0PW3jeIyv33Zh
9CMILkRpln0S+oX7FcqOPXKouncCKPfDnIRBJQyrX6kNLRt/FdtBt0QCdJAaO5B4oK92ejmCahOu
xWKnysCHLfUBytrDR8n3Ms2q694M1RjOtYUlCvcOZZEkeevtjpUP7IrxAk5xDPpjvDhzZIgWeTJm
Zdt9wqqJaTFn6YJ2DBn3PnfebB5DS3MOscyKB6N8JypejZjhRl+j2GFJwQodBxsY2M5CrUGXFutR
jboJJDcCy54JiOG+xaJUVA2ERVoDTGkbMFxaLz9cyFldfVqdjiNiiTsWtMG18Mqcbm6eOHdPrW1+
PF+4GhHEndhtL5LOdQBshIp+6wEvDejzNmKUCaanxXphv3ggw9MeOsfrbudsAzWwPznOEOpeDsg8
/yCK9TLOkhBXVfiy2PORjTfth1vkjKDQMiL6XrnE0qQp+M4eT2Fe/H2YJKSz9KiRyHQVk38lpmt0
k2NJ9XEqdkLqr0zNVbZac35uedryNN6/pp7/UErswE51RQL64Ff52rQyj0DutGGlEvuWZ9HDGUoE
HJVsARg4GufR+mt/9SaWfCkOAnYAx9BOUvDdi56Np8RKba8dfCAD8IhefkdcusPQa5PfJVysydcY
VSDWw9gqvLIohQPYs8Owv19Dvkv5QZwDqm7c/cTmOuWbHHVx0tTDciKPVUJXmsJTIYrfCeUu533+
jJGMygzQz0m3hg2KMjmMfNUNQBWvWMA3UdsLZxJ1rFSzfYqQuwjEVb99CD6U8RSiu0PP2Kf7i0xo
ov5Hqp1/opfdRrsM3By08MIwtjbGZPDK1rsFRTdbp1X7LOnJ1wtf5axuYXDWyIyELRhWhd9ZPAGG
JFyh56AnjTPHsaUlsJII5YqFb9f+27cJ6He9lwu2rcB/i9sWR37AxKxcMUoSn/kdA2Gl8QuKLVYe
t9TWRglp5/+SJcwQYa3melW1j5VuHnwpGtBRQ0trmypgZD7pfTWJdt0YbggzGNLzmy3M51Ha3lTY
1A1NknBHZgYUaRSbXMU61/JgWER4hbi93KyM/d6ZeEeJYHedfYM7yt641RlPEtxwd05mI+HyHSnf
F2GCny8qg7vv+ZxCyQWrXSW13VtYjdTghXnbDFFWWc9Ya7CSFrztHZaeKtcS604QXrsnC4C7uWCu
iasUdoIFEoz7Z2fWR1E4vYoCVZXhzVvesg7aLOmBvU9+I1IzrLBbA/KzJZrX9ObcWePHzskZJmZR
1otz9KStC9EaoMTDG/EliIiFReli1Wk6f6L0VXxfwk3XefSihbrvK9JmNtPrmrexxo4wBZPqnI/C
vMHztkXG3G9RSWUepaBDoF8rZTbMh3mKq+wLLW1v+nGQsMFCR5Qb1MMVTki6c3HPdcaYsOjbkrIR
jzxBxpJHEFie3WNDT2u7IL7B9pvdYgtTdmnaMyYAE7YT4b0iTpsNKYy9CyHyjs0RYrabNtggyWTB
s9oYP8snY7zNP0za57dmiMpeRFRqC6mPU/Wz14kupbkUrlYNSRY20P04MCxmM0EL5ooCS7iy90AZ
fxN3pgy7ToEEtTM7Vsmf6c0+gn4upop6XQuyv6X/Qy+ARvfVUyrGHsTiLp8Ux8XebreSBNxzoPyk
fU5QYDz5cUqUDj04p1RTn8ER8/PRe3hOIte+X2EczCXJOaWbFg3Rs/zLXt498W9Qjt50kmKizDfu
bvx76dMxyCILnb7g93Wj8OrYrxpyePLypzB4i3IEwK3j2p42a9KJMhiyHLFXluR4Ybvbxmh0v4hY
nuxOhSfFx9RmIOPZxvBVbp/lGx6+JqROfR1ujkBk0F7nV+Qy45AD4iCwI/uwZnHIofBXw1A0cTRM
wXg+aCPvKiFSCvrSq1XPmd7GPCNIm/1zliq+NjTwwo041h9PMM3I5yvS7D4eIJuiA43W2JjvR3MJ
FKJJMFW/8MK2MnjBLnSMtX8Tt7l2M53cc3K+ol4+4kdl5RTrU4/dkqtFmibpkQR1MC0b1oW0wQPm
4U6Q2qfIoriqntj7Lne0tOEgBrlqbXJwtHY0pOHVjjmTTc087ImsU4MbHZlgU0lLp/d2QAEQF/o2
H4mCDI7Lt1oVmVbmYlHjIwYgfDdfrc7qmTHczk13kAaMrCL0IUfxK1GhiKpgQrAj21lvxj9EfdKC
Qr96zPpvW0w9F4jkUbL/gN6cQA9/bD92T3/Eysa+aQSzNfzpIDclID4AAeM4cygntKcKQNRLdCyi
ccCwx8uLN74IFvnlRiaZgz5BlL+hynfvlq5wX90tDp5pGhkghBgy0HOcrIKwuqjBQKp4K4mj4luE
vwGy0DsXo+nsc77onyrHwVItQrCreaURnLY48cI1+N6NQ3nmZUOKxBJCDHL96KFGqLTrgrRrvmJH
av6HhO7QgGx1S9RgLG3M1vVAfU2bDc1RdJOfJq/HLqaXl2z7mqe2m4KjQKdDm+c8f4jf17R49SdY
Be8Bq7rUAB0+o6+607HwJcbX52iO19J2CCZSEU9IhxY/TvNnINi+oft8ul9h0kcicvhmd218jJp+
cMAmj2+ITw0AU4UWoevA+p7K3PmTGWT/DhLK/te/jVNy50McW3GS20/HKdDmB2RT5+rnULozR1G/
syicUsVJ9MWj8Uaaj+ZnJAEQSgK2qCh1vEFk0HahPDAXyahH2yxkosIU+xldDNhBj8aw4gFDimLY
sMxREnKrXqZFdrTD58ta6wb/JON4ZSSsUNZ7c91B8H81CNpQ5gP0IX6yWvuis4DnTNDViE1Mj4UQ
XEX3D5Jl7EUnTSfO/NGatz6OF3rcZrjhRAYkud4SpDtTvua3/ODtrUMmAyEobwmTikEkE3SEIuqO
B2/1gY50dW9VLGq49u+w+7tI2dlnBd5eMO91ynvwwKwEn8P6WDd67AJEDmn/YT+m8pXs9oXxsdIF
IYXBH3ubG9NkCWn6eFfnWcPAAYlEphrSqQCX91rkimt+e74BLK9sZorhb39DvG64HsSMQ+8h8d/a
V/YatDf8kfQ59+fU9tQvsGbQ+EttPwLkZ4UfWCicQ2t82pjsCSrEAFQKi0nsSb53arlfPQrvftwQ
lyp69BHCv8FpKnN8JQ2Vcj8cBLFmHihZi5nrbV1tt4Jr+7UKegLQLqZYwWzGOT6fvD4zGrWsNMa9
dZ6qrs6ScbpQhRKsDKEu9MWcu+KeC6VMLRxiKU3nIosQDMQ7GkXEh/OsHsv1+JzELBu8IaYVJSnT
7Lf4kxK62B/4hVVSq2QRm4m/oXPEhDhRvsHsAybGLfjjXqDvKhvrtpzSjgD+LI40mmVgI+8WOuK0
R8iaZUmkqzsaBlf836wEYUqKv7hmoge3GdxS8OVan7pR3oHiWgYAxvAHwJwwvgJOweidkHPYrZvJ
Oh35xK2gtfJzeWjyTHo63aARPXwshP9hOO7+ngJWbdv1TzY75HrbLDme/OPUnW55bDgNo/75ftt0
dcLVGOGe1P6wyv8hiWoTJx8wn7ftUuWBRD11aIlBgNAhpcUS0uQmbtnI8EIHqSvM2y1pVAyjr6q/
4CPVV/yTKw7hcS8BSxa/wOV+DKgXcFz/Akt+zkMw9aYD5GezE9Hd5KrUStygq8/jNGyuCiRZQE3d
3XBulLHzvkSWLpZakN7AmbTeTi1IKtkSGiFyk0UAFaiwtbz8twGt7ys/XZTCL3G6oMvQypdYpSgm
QhQ8USE+6c66Hw8hZMnUW3SbfFAyN467boGAxAs8s8dLhGwKPUXHbDVmSiqztUjLP+j2VifjWqcG
P/UvjEvhn4rOZ5/cYTcxHp7zJn/m8RrZmbPy6c2c9Pafi6uGWD+KIQ+v5vW1CvXPuewtCZr1PxZ4
Ske+0xH1V4p1QeMmCJZF4fEkQE/12YCJkPSRw9ziX+FPADaYpkx+/TmUvf4seBDQHH0PWwKCGSu4
yrcK8dV475jBIB8MWk/3+eANiNs3sPWcfvttABEQfO5VrR3BpBFL2obraYv20pMWNZ/qeJy2dp7O
WWDoU/oX7Pqvq5fYsoBPK8qmNUM2XaNtNRIv+BMO9ZuOFKar1dzEJ6GkYWNNQCYyv9Dp/dX0qHOe
p5upmAZxkEv+qHxwFNEyzYD16fmIco+Dmio+UMFOKrLLpnZA93YjdF2ZXhEh487w8r+9djnvmGG8
M9TiEoULEUF0qKTI02cTCjKjCVv9oA6GDwz9Zhk9a9/WH+lcKPQV4VQsdbByMr8fWHaJmqRb2ejZ
gnCPQWXU+PuJ5gyHfCKVCNWcw8ufTwgrlFKCDq5vy8XSVZ5j9v+g1weXggYz0tJY8SaNp2W1gpLi
LsP41ONxYVH/orz3wpDiprFsYGvjkRH1y6aJpUgxSxj3cpXAsus6IW7+mhV0kW7CZ+QcSVcda59s
I5+6rn25pPjEuD6Ph2Jw3pck+302BwbsfVgGskbRPHPZiJaiBc7U25oMFA6lLPjcu6R+vWE3ccfE
nXsUcpBVfziQDRVDh+MGX6WqnhAhL+Kab/ZDgKBKipGvt1VCfMdq77JTa+ppoaxx/A+bV6wjfWLq
SeSArhiU4Jb5HUchJH2fanqZUs4idC2ml3ZlmXwYR+mdKXFIofYe+Ix05riPigseuGHAAe5lUqAO
+zm5QcR011KDduXq0gA6W2FuRtzJyxEQ2sLoXt3n5l+zPz3E/sMloSg0QMZ2em3t4Y8AjxdVu7fM
e6NuWv2cz62ZsRj39oj0ORz3iFs1sloJ3CJvbJ18kKBOfCcOAvhHVOQQtiM0bosKRjRTzgQMlS7f
LSsGgKSKd8zLcvTA9r3owX4Et4iWzWIegf3g13wPeyB2ZDvwzKeu31mXMstRn0tNhSjK06mbXVmQ
1/HJFKp0xTEathhyWAlLCwT8W4D1Va90aqqg9qR8VWi5dBh94k2Vp1Tz9YrwVbwdjVTrju785dCb
VeRJgRov27fKqbCrg9G5uYgT7XKVSAx99M4ZwSDJWA9UOsDw+dc9OiDxJ+2rvmyeNVukVEFodeCG
0oOCZnHjz9k3uAfnwQNQjbK3AXxPCqfxMSVg8id5BM0+6AyH0OmRcY2qbRhLdZ3dK8yT4FitrfU9
ejKDnRwQX5DIny23ZfvranSPHb25Q7MA2M8B6CZHZRt/hOYdWTZwoLDzBwsPf1G69v8jbrNAAJme
ifZ1x4oQ5TWX2olsOeZOyB1TGb7cd5G+8S4ukfb2ltbwILczD73M47/FzEiN8W9WLmKZe5HJWqsJ
UWemsl1r1uCkClc0kiEgk4HvZekimk/bG4hsUucgzN+Cx17eXoFnaJSlqKmczOEqxhe7qECKGb8P
eCxiW78zOQxMz2lla+Bg4I9XiAKfcMBNvRVdd8ZEN4bxpAYaCAtyYTmCIKBmMeqM+yzeFd1nm+sG
Xpzis0FmoAIAyLpM4k2xhKm0hl9nh1vIQAwaH6ZhrXtXf5oCep/qXW0x1noeCrHKdxl4plBkScsz
4qEF0RlyNm+jUvCZha7RijsdyxldXI0vBsQ5LSvp1LqQaMJ86YIhRalsmu8V9IU40EvlEUsDybHx
EIiMDoAgD+/diYbOB7gUkzaDDrxpc04KHeQpTiviCxo7Q9cuLgD5ZvQP4M8luy6zi0/fBTQgo8iM
qSMmObRNB4NkyWnTqAiiQfe/BVcK3OY6H8onr9IOsZ40g6OfKTWSbCCBeRPGFvkZGaBK/DFBPZfX
+fIbd+u0DyNnVViFAfVKfEyTi4fCumuXTNFIbOJWXmm8Aq34niKb5cQMIqnyb7tKXeh1hahAj/sN
y3gAmBuWPMrQv6Zuvc+YirYK5gpA/OUCaITHb/0wM961FB7rBBoVcDLl74ALN86apZH7xew1KwFu
F5CRkqD3Yqk3erG9d6mE9w+BvBtU3EXtb9VzNdw1JWvoUtrqs2WbKCXgWHeCp6lrplQbTEVRIKDB
neMfq3LkTG5DY4aX4VMKnjnjRLABkwcu8kiM6/419sTMCeKspnEGeAv/T+QpZTIO2kxdvnfEPe/T
alSuigGrPpR74t5iZZwU8aBWhWONm7sasbicd9hv70h7ghijtqRRKM0KEgXxIpTeKp3PApgg7b19
Cni2hzMNbuDAPlYCN4y8+P/TXEva4tIk3ceqqhq8KyrsPzThTl7WY9WfunH01HjeUsqzXc/JyW7B
lk8r9TgYBSEgR6ksZwTmkRmLf+CVmCqvQ8bQbMESVx4jOOBq30Cp+JDoUOr0XBtHEFZRNDqGNG4w
uiICu2UTwOt4Iac4S6j5dWzywRu2Ih42ZkEcJ9Mu4MQVa5H0QJ1uAf65+lnAFLnfuxfR7CvnKmTg
Jpq32x3MQgD5NIrkNluGPC/AP3a8QMBWlkmTRJZ9m1GtLSBsmbmLr0aeHt8qNhow27UVj5gJXF/V
mVSlEM9oWspShpiO0d8X5KuyTpbi9AGoBEHf6T0eVqO1Ihfr2QUvFUlu+6do8kf0wJVAR2owAU7+
p6E8Dt1vHeZ3KUejMg562r2CC3VxRchtAKuKQiJ57l365a2am5+f6c8c1Lg5nmCwZzCAdhS2AZO/
+CgZInGRkaAdU3yg5m+7Cxh0IiB7pt+KFQglZQgDTQvMywigJrY2xNsEWjcdw5RwFYTmLtG7TvAv
/hHs71vtutYYYF3zBQHsOgsfmcsOIUBT03xeZAod0Ljnigr3rXxHxTuRVkVfcuoxrPu9Tfdg/bjA
kCf6Al86LwmlNWxT+W9FJHz1B7xrcN2jwOt9Fp8SLKL7kyjHwhAho4gT2OpgaJDUD14K8Gi5MHnh
6sUOmw3gbrbFzF1U11MDyPyd7JpSkGSFEyHPSZDliEKbpPVt6r5bwi32BIwz6XAvuugWHbGMrWdN
ERn+/iFXKrJ42sQXS9WtRZh6Z9cTLY1zuGkCmCNOB9G645q7ebX1ajMGeSA43VQIn94CjM1qy9vl
7o3gySYC4NKpho47RP0WUye9Gh17FVZf84xEXG38SukCABPd58hN8knhph4SNm2gyDm/tQhOCvY8
jni2ef1L9c/j7lUmiXZAu6Oy9+W23RiI4a079R28pD+CUUzA9wtXlQflb/5McDsek5Un2DDsegV2
tnbrhePt8cmmCwrCqIbe6U+tGuBfPTufMeg2fU49ZDr8VM1UXjGtBhsUslHrlE14fONXJRQF91FN
NKYfzMZ/ihhIK6culqh7mRvus1fRYMixf+98f+9YT/pXdbC2Ti0vJ+bMxokSHJdrC9FOajHupTqz
ZSM7z5RVom1YKFExviyPg0XXXRlCEaqIcIV6W2M55akJpotJo97uQEisrz7wLaM4SsaSHfsfUjGE
ohGRCUThbVZpuLOA0eKsleujm3T7PQzylfgsDeboZisk3bxx5IuBGHZcCZabnswro4vwfR9dqRYe
XHonXd1SX4eowl98SpElq1eBM9kyv5fxL38M8HHbC73bjSVgrq4qg1vfe6EzGQeXoDtbysYSKmEn
qy8tsvLHZJ9wFiGRFRJaEntMhaBbeW7DSeaUfA4awzRDS+xMKVjZ4fzlH/B4xtIj9IIpVIbLYJhG
5xGr5bL5F9HMgSJOnal0+wp1KeWcgSzdwUgG1/JVD61AIMJC+Bk7483C3x3Hrqh58X02ZCGIxZFn
6hDqCwsthkOuRuKoHPjv64WoCPIcby/btNOeVLXMH/fZPkFRsIlODnHfiY7hgYJM2sxkdNJ5rnPq
mrfDqxON0dPsjhroiOYjelzvfwa/yhL3sxqlzY3CZOtgG7eDK2M41JYBhoEZjgp4ArRyi1TZpNqi
eP6yCgxu/c140+UlefaU8hZvTnylxX0GP8IoRPXDB9LXVKiiTgV6ssQ1yL5L+ksKfN3Y+gdJqzb8
NqHia/fPm8DZ843O/2IURGw3pF4utIBxUV01SInU7i2+b6Em2YhHg/xHICrMRMivEukJWvU81uhG
88g6Ywxx96P/xAgYjGMMYEKJ6vPY2l+Ax6JhyYkneySkzzRyxe4xXKpQ36T+KpCQQ5R/namNNCaa
5opKK5wxoArpd7IOFwzIhXj3uqcDSG4i4jl7s6oS6PUtmI8kE1GS4kUmrgGQZJnP2X7hfODccpUe
VFHVjT7nnPCdDkdDF3Rbnk4vUx8twJWjbmf9VFeZ2AVnQT7nVuSoc20oSWzCEFwD+epP5IWKPe4a
6g8TrSw7tNWyrWvLTgzC3FAgH4V5q6vCT2csvFAaUQ27niBpK3z1eR90zXHNzZVnH2pbcQdewolr
zvctU/922eoWP8r7jX06cBVDirIAGJPUUhYgor2FSM3LzdCWruyyStQcvn+ngVpb++4Lp2wZx9Kd
BAcN6JCmG9afZ70udzgMndIcZ5Ub/AjaAK8+a5mCv/Z9RizV/X6IXM9lXQQeyqs1fmoAVUnYrY2C
sJkFUIW+vTK+DX820ndCc1eWU15kWryckevuJj4XWxXFc7FPJ1iNmXiqBcPFPJtUQKTi1Og+bSnf
vkI9Btk35TJufsmxFziy6LDYpkOfMHtxXN5Jif7qosOndjMjN1cwbJNxX9655LNKM4vM/B2D/sUl
JWJ3J8h2r/OMylIYoKBMPgLmerA/JFuu9hnXAXtddfrPwANwxd0+2ETRyanYGFIbQbH0J/sz8Onf
7F49RRrg7Elo4ejVR3b2NnuLLXZ/rgPSP5HnYetZgGXwzyekl+iMTfRG5EvsZPUqwMZcbzH09BTO
KtCA+om7ccz3hv4P4+HkFkGyq+Lc5pB7WAdsgYiVy+1Pdzn404C+HrJFFHtgJgVZiXX94JTj3mQF
dGAtURenwSgh3RJ3Mp+A/A4oZ3WIebBC7l0G02Z1/YNLaQVjVPivEgRGHz8Mnisq5ouYV9cC1vPF
QTZ0bZBICcE8XCuSqpOjcwIjXoGpPT1cKbYjzUtHR0mS8BfZqwQbtHdmoidRv0xC3whmXf7Wp/vp
VsZ6JNNGJlpYHRzN/Qbusw0w5/k4ZTpIvM3bgZhcUEUKItxhlcdE5rlwDhSAvpCwmA6KGM1W6Z/G
1tWYHpQoz6oIyDQ6W24FwaG1YE7b7Vi27lNFgMTWjrA4syOefdN/r+zY+xuBQ1qkMLJHOnqk8WVf
CVIrjZBkK4nho2Q3iChjz6RJWdgVSP88tHvmLrcG/J6ssX/TQT+rTWpixgCAdq9N/y4ZfJWAGhNp
KsEfObkZxAq6tNBZ6iNzjl83fUBR1c5EPmuqnQwGxkxnwrmAtkcBX2IljMazNUDQeCiQeb0Q/05U
OixPBLYTpJSIbOPopheIgqno5IWIAY8soqFYDEqsFzGfBo8X4MmfYcaUNnMFPqebe2j9VWQeRb+k
tCeSGOcVk0wUrLtWcVX4PATT2aWgCYL9oA9LxMdLuRaLVHRpSfx0PALby2CeJs4s3HnPOmolytG1
ndXpdcX9cmRYFAypYBTSwQhJdvf3zQcuHvveGkL/FFALYUKfCHRB0pmCrC7o2xY3tQMO6Y0YaB8d
SMAtRr2RIvd97sZfyyehUJc2VAFXnZ2aV7mP/qObZGuoS/vbyJeeq+iSVqlA0Btv2StDAbxLgEvV
z61BxJrEoiKcbYAW8zZEAaTWTC3RZgX+ByMU55O6KSM+bALlG+PQX+gQHKoFd/abVF9kUpq1lgL9
bjd/3bj57KYscW+zWank1xDWoe2WutgKsUew4MsTLkIm2pVEICJbVAAlqOTtXmrOoKT2hF0DFdwa
bO1q0ePHKP23HwlJiNAkvVh/rQ7+7FXyei6f8sVqBuVQsAKlrof4RoZfx7Gi7usg08p3rKr+kaKz
RcjkpKUvq7JiGpAOfzwbHb/h/lTI2EqRI3rUrVMxe4R39kW4zg/UVIv+84V+iedDunCoweIVLXl9
/hnbDR1mS7fc7ELB4mJyYdR3cp1/SH+lJ3qqEOTG/0cbpwY2/wzGkgFIER/4chAV60ZaA3iSNdIy
KKQo3VKOAi92jQhpDVPP+0N7N0dTeOdNsYV48Z/oefqPVLbIhrHRJnmyyPJRlGibMWl5youIj8BZ
u9mUKYR7QHesg9YTQN3xnrNuHWMa9B/r0Nw1QllsZ/1H9ahaxskqGM+/3RX7RblengEYcFIzhRAa
X0FauR3I0aLyJ5aZuxILHjw31Gi5UiZn+agEyJTYr/iJok2cR7dN27BhEQCr35fCHpkCH1XOWY60
YltMxJ5MS81XdrSEzbHD4MBHGuKiF70ytWRXKZ4W3D723NqbWiocyvyP/QPaXwtm/m0G6wWeQVLo
gH536c86wlxqnaKETQbahGTK++RrIwd6UwthP8WSBfBsdl8Cx4OtAYZq5K+ACzOky5NhLMOOComg
LIWKzDsaI9ae2+yNL6uFAqSC1gOd6wRT3rEBkxI94Hec/tKVzG4VvmOl4DWD89q6oJLgVoL4/6Y7
GMmasn2U9+cNTIosHSEqWnQ9sfX3yxOdLvGK2a0Ojmmn5CPzg+eG992Un1hwm2uucGfSnlirovfw
MwPIGhBS1mT3LFP9R65e719OoUkEFgS7bCR7BWRJJo5DdOE/C/zymkrCj0faoroyLRmmIhSOA4CY
pZ0wAGE/ov4+igxNeMAfAhkqfVhX9Gvrn+1Q/zfStwP/dodhp//PSabTyExGWIwbQnx6l474UAcs
DYW9Wj9zIB3D2Q0fB6+DyZWOsNIjr0MryxNEjV6DRHq0Dnb5Y+PwUIAJThuyUw/cKGU1Zqjj+Pn2
/zldr8FE7G3g5vVE/EX3d2sFmsDn2+XfNcljsRUtBY8/ltdyaj+2puIv5OZX8qLFhDsFrQ1AdBXn
UEmPbPtlLxDjYHM+SFpF+jVx3kv1uS9F1lEuWvPpKsyCWJlkfkjYZIIW2DmI06Bb8wz7I1U7UBwQ
xhFfD2gSZ5Y5vgautnegc9Atd2tpPgKAqKX200h2GhQcirM13Zdc/ri8hqJ0V+k0pUuiD5DL8+y0
zv/mfJkpJmCG7ngUHqqaDvmUuT6gM7d7zUEA40lci4jLKOHxjZrpc1wmNNN9W13Qe/dxh3sJXu1c
8ymXcAkGB7LLtTe/WdWIYTEspqGq3FtCzXqUqJ2d4c+c4IJymFSKHQD9ls7DV40Fvfcx2Dn4UjeK
2+4N2YefneFB4CbkRmUXiArQE88Lt9Gi1HBOwmk0Tl0xjfnz7Ai2n6hMyt+gmsa1m/VnPniNh+80
bqAtKTf1lzNXrcaCWihCwSpiYigKHwqNqKmqq/KzUXUgZAj+OeRmD4+U1qnpdyyylw2xwBYO8vSH
MtrKwKTJGN5sayJyVryx7TY+DnZd97cU0rxD75BuG0iFFW0AgHIi1qkie/8ovBie5/+hqRUcV7ok
AXFKzzcTX0IRGcTbIxFwVY1LZ2LaRzt0HyqUl11/n2DAcAkDgwnACWExiaUIf6AcrBOgVYYfLIMV
JcnF872vddb/qq7LPXyRZbs+9c+DanXMbw2P04Cs2sKqW5abl9Gb8TfmUWYEMxJ4uxm2mcBGmGCc
AbiQ+4FAEBjcA3XRIR36jw8edmeTdj9A0miOt6lSX+PZ2bmjrEBNVO3bKCvDnIZztSlgitQJF6MG
qEFO6y5Lfmrj4USv8tcSk+v3JQZZX5nyO9cB1ww0TyhfHoSmLmbAYtxcmii3d5WVcxsAi5bfBeM8
2cOV42D+etmnmPrKOD96erT+BJjKMxjcLd8BdL+D2NG9YocXfwJVVqVz2EQjxoRaLBu12xVXzxCx
ipOeTSG1aHNprUY85D6vV1+F4f1OpyTLhQuVtQpH6PeiOHfNfL0l0jlbWi6EryyACjpyANP4yS+t
3NDZZ48Oh6sWnEakzry7mTQRVWx/bPzPTf2iAe7XaUuEfBGYLjB8hXbELyeImtJdox60N0oZFuAx
Hdx85QZjcvNwWK7VzmKVvTmCC9dL7Oi+vDOhejxioZRoR+DsgyNMwhXxnr99miRrs+MVbYVtJxYH
Xj4Z5f0MmzyAwxN39zWkQIDrUFc4K9JFg85aIGMf5Clw4GXHCdNcwWv2g0alTOmDA7XKdq8CdJ0M
ycTIFCEuAt9WAg5eTljCO5KvRPg88np5Lipn+GFIb4+rTytN9p6JzrSb6bLhY8+dGP/D4HKw8+ed
PTbeh3adKt57GkUY6zULsSh11Zcb8quyGODK7iXOvOYGnryOmzxrh36kQ9nehYdhzegPhEdzqUq8
CpbJH5neOR66eQzG8oGKUSiLFQg9QhmPfskEEt3zXxizinMjO7hhVygZ6+OL9X+TjWxHwqGUtYxI
7x5HY7rxX7A2obDn3hI2/j90zqy38X3Yu7vtLGwvrJfMwIgoXez5BR1DoxsRr1PP1SEuNyLY+5oB
X7Y8c/29EdDw/vPlTjPsFkdl0Z917EU8uS5vtJGfE3BP6IFDf78SED7tinIKAGEENvzodqXHt5wV
P/Uv7DWsrVVquC8NGx01HSlLWt1k0KFo+Ru6Ifp49E+xzxieoqV/hDeOAxQicTT+iRhUn2dynau3
pIQfZTOpCcE2NTMaZyPZj1HO1mPLUrzedwJy68vwkGeQg6fYyZYbYa02bQPcYv5zWLoK7KLE0zqU
hDiMNDJanL5/eSQqDKoq+pJKdlPPzBbHw13ysxdoJ6kzXo1C6qjkG9AA3tz18ziav264FlHl0ZVc
xV5kxzfCzwXYCv8C0HWRugWoHBpYUoyGBwtShwGnv0YGkgG1oA+zIuRs3rM7XZAYLFpq7xtDYMiJ
xmziMPYsDqWNCFhXPlKmPajvOswGMnHig9M77czLsLd+lYNQYJW/eSsHejFmPB7KSVX6kvwJdZ41
pneIDyLRZx26kv3EBWWoM1cksLZUUDCLAKMd8msQcpx1B6l+D0XOtBQeTHLhE3vNb78pBXzCGy2D
vkmS/ln5rmZTOgJW8F0MLQEkHzWdn2/dMh0kthnttb9T+E+yixw1LildrQ97puHtB1bejH05nusC
ofAAp5sATVYJnrMwRlpeVpGhk1SVLH3veSZpX2qliwOv+8APMf8gPPv/2EmZBvzVEQI4db5guMmb
scvC0oznPbgO95ZxWpUoi3hO7AZ7yMfqRLdVrcnK8EgOclj8yqNkVUv0nY4ZW9fWycj9jehY8Uyg
hYOSGWol7T0sqmsynKzB5acEVAnlXLyI4n1NWnNBNgq8MD8yGGerGduq+LRkepJxiyhwWr1CFQYS
hCrCd2m60bOxOkHJu6eVHL0eTvX4oXXi7AkqQ02fURZE9V2t8e4H8G3t9vADnZOahrpOjmRz/Mzq
u3nVheobqmmoA1+4MZJiFe1mIRCG2cfh8F6yPGeezxnGU7I4wRVw3qqQl6NvIW3qPU0Z9G2Nifel
uv2RFMdfKBrYivuIuAaWjPJ0fjYB1tmMZuERwoTEhjI1tKL5L+QTRYFB16ndKnfC3N9UxPDsvEYR
tv0LVOjrokzNTwQ52MT8+681VcT+qkys7EEfi6cTBjE9qH490TQaz/nrOvvopQ2R1cowOujC36JQ
QhR0eaZig0A0hKIw0MP9FzjW4g2khqAQG4u0eR7OGY+KmRr4qon/mU6yHMupuwqWwagqWIb1D8d/
Gaz8rFMNt9NkmtSnQQCpkCpPrhRczKQ5kyL3BWuYdXJMxFWCCFbQGObO8sDPKKm1ALYgnqjdrFyU
+LxAVB/5gphv3wQDyn6kbbFreimgEEY1T6/NacWZMgn/o6S6UIRSgsJg1lNwTJ+5TyX/FzCRvDIX
3ATl5VowxS1Et34C8nZ3r+54oH6loA3o/wifbLQRvxQyPxwzf1HDNjJYWLaz/mL3UnfnrWQJs0o6
HcB7mqU0pdReRiAU+2fBqOpYV56UoofefdQIjtIHywf5pnXvK4jy98e/C/PUVbo5NGIAEdTycVMo
xs2xnWxUA1EZDdT/Taoz3UJKgO16wWNs+B++D6FPZHxosX5Uzeqyvurp+xjaKyN83y0R5TWTqCd8
ZSZUxIqiamu0sypEBcEYfotFKhjpVWdbRjJndNqoUPq7sgLUItBYxdAt6nuJGyRoS8HnHSVNcFHc
8JkK07k6MN6KodzU4iRsoZ5ANXru0WbbwsvpzVJfmW4aS387m5DNE7X2SEtkpCTbKiOEzDjZw/F1
m1co7K7pOQxvMsio5yPASJuQfeOS6Whf6hs1gTcP8Aiw2GaSJz0Q7gC5yo+OcEsTx/n6Wep1SuDc
2mJ23BZN6luG0q7SZ2HLS1zGcY64cbcZmoqov50+KLdamO327/NepIxzSoeT+3aQoCpNvRhZlbTH
Smrdh86CL/4lGq8XifbeOMx4e+1/GYpksDBU72XW2FbS4cuJwWx6AuGg0PIQFNcUOfVqZzo6ykgV
tACLOW2N+/t/BNabWC+yxWEhwYWliiN/tDnYPMOmDF2uQTBPk5+JSE/XqgVX05cfIM68bLd0tunV
DV/i/qQxzRTAwzkf3uNhTMSZwPDzzDTfc2ix8JqtIK9ihnHIbjHQFRvrHUldeUK0WB9o5yjxZzlK
QASiINj6TLvUVjp4A5rPls2sO812bZBb1ytCB343gL6WVCrTcux8Z0Tz+0656V/iya9mjx80jpRe
uzpNKTRcwk7/MV4ZLN1huPc8QnMUk34Sgdmyyz9O+5udQIIWww0rdcetSpHDNMVQ2pTmmrULy2Fj
LTEKkSojXnQoX/CDZYfFGasf+FyHggoKqjaVozTtkjbDlai3FZLavM9rSQ1Sg18P1+VIIPkykTPn
oiMiQAOqomOIkpADJ2SSBY9XaGyzdI5MSiJiSxCru85wG1TXfg1x3cri8O07XEwGclcGiyQRx7Dr
d0QOeLrWKU7R3tzAu1Dg7qZuFbZblFGRzwaGObKPQCmmkAZ0DdLZX4ynstub86LTEsgmxglFZ/LF
K0SKa31AykBYdZWEZS5i3Yrr0Lb1sBOzA29dIAd5oQXgFj1ztYCcrVdgYvXrPJ5SKQsb0cqjcbZt
IsYK9M+T0ggVuRI8oQBKdVVo4PeSoLm5AG3z7wP5S6KdJ4vbBxi3erKkA9BsUhM42LQlidnDo+ab
DpsjF68BRSDsdjJ0lSEu+jvAZ4kDo2hnD7iLv5NtCb7Z8NcPjrDMOaNNUQ17yIg8I2AxMyIvEDGx
O25sY25w8L05ar/IGyDs6iEIypQNYVaH98Vw3FeVKyqFk01CzIqst+dgcgjEYrb19rxgATjfxgwl
P8e8+kIAqq+8xsQcuIJQkaiclJy+Pbq5yYWWIPby/p+z1Y7nZIlYrmK9RbEP4fSArV4yYobYXxZW
weV8MrPafOsuU0o/FVgnqKMA3Smh/Zx28BTA9UFn+n8ao9o0ByN1aiVTBM41fhqzgh/bQ4FQkT06
8WKLP0AvKsUgn9J97ZUfGmtLyuJ2iX1Ee8lwDS/AQXJECfUhq+Vb7tUoBJ3pltRs6wXYMPksHK4E
FyGkU+v77gdg7Wv5Aux94qT8KylME5X6ZjGWRVjArX+PZHIQfNJD1NR+eu1ysEJAax9wshm30/a3
cpF/KCuaPEkaitM2MygfgNTXnLxTvcvSDSvXzF8r1Jow58tgg3Hgq0z9/1UhyuNHVpEPOo/siM3H
RS1gtSWJQ/TsqsurCmkroZI7ydtlELl5c1Qg8quVgfsX298qDhfZOwZHZLlkYwh0kymmH4cn5KE7
uUDsI23SOAIVyD2ZRZU3WX9Hyl4PAhnWxBBK3syb4I19iKX3JAr92F/FTo6o7j9yYcNhRC5aWBq8
+7hJCVqnu6ar8W5ajZOTcwdEeu4UiD9IxtQknJ6rcAxQstBAcKiLStc4H57VgVekduiOCOOrlUlC
LrrfxUG2XzaRCtjNRu/bJrbx5SQANFWpSvNv1sNh1U+HNwtchULa6UeL0OR7Z+Fdoduj021lue0Q
3ydxeFijNCPza2sL/MwP6X4hlX2A9nsgC/mlmV3OTJqRL1FbrWohtHezPsvDiuE280A6mg8MYrP2
9ivpPtkVTbZWp5EG4PztNy0mFz1lyxlUgAIuPM72QoKp2SXr4mIM0oswMIXPUoTJqvEjfMCoriby
McDbVwiiOUYmy08AnQiTzskNg/+o9ALl5yS5BirUz11etU8yXfIXneFu8kys4zLIEY58Ci/DvZ1v
3gvQHzhhBVSQM2FTppHjuuX3VRLq4ifQK0hSel3eR7jR0aEZloiHJRkiQnBrhayYeaPNLueUN0h5
asqtpvdncf15hHKA3PZt66Tg0Zco5I0GEebKliegnnbkAqE2SyQ62LE4NPCGsBcNEQNLg9KF4jG1
yfDSQoeVBqp5oszJ04N9sP51LOlh135zhLhY4IpG0E82tkctPYNPBOd519Oa9lltf7C7Aw5AWqSI
oodNaRvTTt669OE4w1r+Zje0mQFbDBKFJ6QCMxmGShkuGHKuUYOP6MFoZwJibBTdqcDzHegFC/Bj
hvxU8dcr3MUbtbg5sB6oQE/MrJgJ1RYmfYTmJQSuVXH+Oh8lLZfYefgaO4CX1IFMQUOKWBi5DwBE
uOU10l490W5HtDecwNh+jNXeld3K48VKbOzWlM3dmrUQPBfPDpkscClJofuWSBu9xYBjuphxA/XB
17y60r2TU3VqdX66qLz1CymPjD3cL2Ngp5wfnOVPqlLv0EMqTNbG40+fSbyV/qBaxyqgiYrqtHfb
a+D0JS1SZCOn+ItGqdV0gtGspTsV0jxgD+WiNINGP4C15N1tHLTRdIxmKNPyMueIIJ1mtp1GS6HH
wAdnhi66GwXckeazWvBoIsrYmEQpJgyOwcnNVRXQmWLlvJ5LPDrzXnBZZmpxQnJGG3pZrJeF0mMY
EKt5lZpEUmFVlwnTQjerh9efL0V6w8RPRpmlRnP1s8hJRjWNoG9UF40UR9a6uQ0qpLQDfTinBT4Y
69mk/VBec9CdiaRm4VU1n5xUMDTfjrETpKef6LjmBlwUsLTQ2EWP/jAg8SMzHq/JPjn9m6IGszCI
2slCwxKAEN904kND1VEjBLYxeji6LUfh2oaYedCeSY2QpBUniZKz3N6TywV/lgUFosVW8T03d8v0
2zCX3/78aVWjItyjQklsHSBjZpxSl6cuF+tP/EekPYusZ3YPIqooSa7xgLI10+UVkJSeuIx3490n
q4wUjXXRcxRVPg0adRKcBeKM217+cQd78QxY2KNdpmWUrfoJD+vMzA3uMTNdHNKgReL8gs6REO11
9IluQnIz7vVaBr7yaLVDKxqfQc1RhX761AiS5vT84N1bSO7KFSM4MdOgLJhPtuX6o/RqarKluDSx
QwtXoI7RPntnj+B2HCYDEMfzhExR9KSx8x4CC7KvH479XFXjfEV5V0xy+euOIsnwIdyN1QXdGnXK
6PXn32y1c9Sy2mlrHdmvyttDetHXzJ3e37tb0br7qlnb8JDUFbLyPRm0MAip6Jd8DxZ5hgI5Skpr
zxBO04LvYP01rdYtwPRSciygwKyDhcZjP9O9+ornas1vYG8SMsdOVpxttw/vHnz5aoziWOnzwUsP
5xHznsukQXOPGFkOp8UmwK8faGcOInliwRG3H6ywrrjdNDOnb9V9Y1AKQIqys05EPWCMtKCFRW/D
P1N7DycXmp2lph96t2lmRfDxuV7zNIJ1tBIh866C36ni7AFaJRDEFEFvr91qHMRQn9ZLXTlaahiC
hTuyGDzDIAn2sXXckNQ4Eqx/fhZtzoToZhcjXMwa30EF+RjOZeWleHn35pEOP6Xi0B3E1iWPYL7M
2z1DlnyjbpLCZJSCowN7u4bHpL9zHl5VxYSsJkXj7tmglxUzC+n5wGyhFo8e2JdU1a5KIHzh1t1b
FkW91CX5CqMXx37xY+hSu4NLrSXLu9gJiFUhUgzNvkRb5s+LnULvE3U4H5s7Eq23uCaS+HfiiVCL
geDeasMnb0oVOkICQHQRaBT/+9m4ncXmUBnSsIcJBfBN686bEvKFvf3yVHqxtaQ3WX0LgpKwvgmS
CL18xJys08Zp7/20yqF7LAE7kU3RBY9b+oaobO5LhNKwY+db6P5W600/Tsx6oMM3ReuXqVvyQjBV
5+2Y74n05HY9TQHFX8HUd8zoUDB1OBCl4iIhSBJl6adK9lsOJb1vDMaBJL93camHIqUXmLy6f3GA
fU/WgJFdoy7uTdICQ5dCw3eKbX5cbVvJJz45ab4QRRJP32b9QYUuGl+xJ73bdzpz0lJuGikIYY7c
3NVKpFxmF3uWwqS3iRi4J4e8y0ctPa0Dr7Ram72FrTKNms+iaio+4QUDqyrBRJT0XTJ/Di0VCOQP
Vkt7KA9vNCrC9vRkPX0LIcR4jmWQFdt0jx8R49Vv11v+Vm48fu5WPjYF3EowDj/KzTbGWUGK4K8x
7BWq2VL+SOAGMAWtb3r1nRb6diXYc9a9c+nYCkL7gj2jZa7GeX65FqgcJ/YCP2JmRF4AIYi7gRso
bP2XWj086UseLdWupL+fgTk5VzQiyAp9XPPpLq/7ebz/tjq+Gc9oP3zYngv8BcbL4TpgsX6zJASm
all/Fz4ZNJyd2VhYOUfJi5LVVGQSARYU/+FOQBg92cERVZJyvh8NG2uYIWX1EnF38FB/T3/RHcZn
/GRfcOmFCFTCUMjuBIE7KpuVHnvJ5ecl15LotOv9UEWgapqcUDQRYFO+4stBGhlTg06kfxbVvazP
WhXh0CVzddLbw9A1/JVJYjn8kMJm6bYA3R6Ej3Wii+MZkol81ecdsFFUv/3GyTLTiNEYFPfeuyqh
mC0LObPPK0YCPRTG2SE9iUQVLYzy9OzVO/6cxPdETTexObadNAKiIhB1bMejY6SPQsOa237qnu/1
KNr23cr4zjUcwLfBYIdNG3iR/MJZj0xEkQWp8r8vfg+obDnsevDLdMa7nGC2JayLgul22uY64cCR
Kg+WA/91FXX/l2JE1nHxYhUL/ENfU8Wan4Dl1Oqzpa3c8Xt1dYc1cdEWZuc7P0i+lTwnKt/O8wwC
QSmSSqWFhLFQsNddngRMKATOqN3NfxmeXAQ4NovRXg/pmR8DNssUEHDp+wZPCF/PTdmDiG7qSuWf
s7uPDGRJa++bBOnLe+mboZpm4eGTQ40C2F1EDZClwrkAtS7mkRgnTJy23omgWOLy/LMUFQ322Azz
uhv+4Yz7Dx975OezcpBRye23mc7+tf+hVbWq40Ki3DeO4yJYVTDKdrnVFnY3K/x0UZ5TCEIz6lwo
gEO98phyKJZR+mc4aVj2/qkUEt4Zr+1es0kGzN6MyBNGpB4ppNuG6VmK6aev/OuK1+fS5ew89kue
bHr5IUNTHexCQj2INU2M0LPFpivGFlnuBmtIEhswWnqhN9lKGxdNZRiYCfHAJyrODthh0FxNtoYP
J00wiRo/erZ/pJPtkDA+K3VmwW1SJUOhs6kaaVAgOha100AV+or8kbNT3+sIEKMlh1/KUFlk/25T
YNgeYiBO9aV0L/pVfvMYW/+I2TPdC+ed92esXU7HS1TxNdHpvVf1dnNCR1m6bck3+qahGYW/05jF
W7hjwu5vXDlwd0GUZj/FrUDFxUFy4pf/nL9B+GR3iuqALi21lpSh9mwXt0xjVAJbNjqDVJ9KFNTy
Bqy648TgZzyKPgxNqL+OX1WRuVJ5tRiHjvINq4H+7ICeXAOeZQ23GB1f/2Epgz0D8wgAY6hzV1Up
eCmomeoP5l+8GHMRmYCWPI6NrebWrX5NUAlExq+qbxOIcLNT2K+Jka2nQxHZiDtb9HE179h+I+EG
YG56CymXDzg8+gTyazktI1AFBW7P2VT6QSJK4m/igjkBDWOl65Ee01wPnYu8SwTzmHqioCkJ6tb4
b6iRWA8DXeBPWqso1THZf2OcHZONNEq4MX2d9aiHSGAQMog+eyE1mu8COy77EVkMvCcGS6ZrR0s0
ja/r0gM/uCDdEF2vmz+xkDpaMcWB6VqG5hoA0YsSyBYdeK1XKCC4PDjDl6i4dAk4yBSTmeIiwaWe
8ayEhe4RFEXAoWbwyW4IYHoLnvQZVNwOK8WY7Hr64HHJye/13fDqE5f5EvNJI7WrOrBIiCzTNbDD
WfGbcjmTf5poij+aIS2xJy5jq1mZs/rE7rtdrn6JNkQhDkAHpBdi4xpkNS+K9VWih/7j9J96q0nL
SJV9theggtic8lT1qby2ddAimjgpqkNdQHJ8ELPgZGJVkkiVXtXI9N6hE5J8a7VQ0QReK2qnF+bP
J8jCp2R1DtMtscLedKXVrTW3Ls+rQx67Yn04Cz9dfUSvA8Ax6Z4El5djT6/eelf3Cvyj5s2a41Bx
z201dhHK633XneP34FZ3B91eEKhccUCqZF3KoQnmtd0x4LsMfHKVFMLdX/+YkYxt9Yfj1WFqr8Du
IajS/RJ3z87fB1FESsnavT1IdvgbxW7uhqZac+S0sLAYhYgXRhuH7bBI8M/ayLdd42eIqIKMolBf
CJoyizzcekVVRmJ/FmzJNPQ8f41wjktuP4VDIAw76FH+/0oEHACbhpoOWnpvwzMGLGFgLFvcQ+VU
ytZHTeosmOeN42rpiITCRs+wqqwdaYLb0eRGEqejcHVrIYuiGxveCoFq9rsWCrCDHeZ8ndvjStLu
v2USEiEno7xpGINMlT81mI507Z4YCyGYz+p9lppGUNbGr4Gm4jWDsXxorrp5msI4K5wG2OngLXjy
uQVeWWcW9s7LBNYM78OljgGtvAXvIybIo2Nx2idBowbBWLYPkj8JMhsP1VTfTWilPqCevQAyzEyD
JZya6kmFKFHIcaBwMuawKsCWgqEXhTkvxLYJ+XxaFIlAAOcbmtmd6Bleg5NZLkJBywoa5T0VAC2z
IISodLVcfTItZoOb3IzS3oRHp0msxhr4CJ/pKmEIxD02f7BwOk6eXBWkXR7po6UnSy1VZYF4lUhF
8z12iBfF1hG9zW4ae/XCkZr6flliIVj8tWbHanHCYnTlfES6Sqp4Aj5Q2tmUu1Vj7sfp++yONF3S
SupxYSYynyAGfz7ezDT3uL1xQUK5HN0rfSXeWwjBOe0iy01SW590PRwpy+U0yAq/oA4CgD3rmfui
oG32sitQ7ILTw3hObS2I6MFiRNEt3ru6+B6zWNf++U3Twrns4ZFXygXkOTB5He3in7jdb2Na6mCh
kzIa2/eCt6hFCqUXrZl9YjBKGqs/PMK+bVq5/a8E0HOcekU3ULzd9RcROBbZaGymLojEsZoTs/Ao
iKtBGjVSdPocdXyGz8JY67uRFFycGYhnxpfzD73tASH2axyAooQ/apiXhXEbgs4f+u2RFldDhkbR
TKlfS7XoEHqe32VHdYUx0tHLX36pJ4p2RsKOA4LTs7+AmpD6p21PLFcPj4DYmhV9paaMUOLZVa/p
yBD0M9V98hhNvopBD8hjuqHniFSzad4KresYriLRH2HIZ92kEZsWZynPN+xNyQ3/Y0M2/GOHc9oc
QnpuuYQq1d2BIsjWjLgFg4/rMtcT1+mLQRRpz9+HnFMnZ7NXT7C7xiLnZw9Nm/3/oEbJeKEUpjjl
riVmGYxiRhEidtcqSzQTz92aReY+PYyFJwaiNUXuEAmKU3Scmmcgd5eioCUhNeFoe6rjdVKgv0fo
m+zTOR1uq81E+8wgsHg1YumE93E4Bx77f+4JvvSxFU30qHXKXurk/xvol0ZHkMipwalT4yQ085Hb
gGoRY4D5W04rwmQKVUSGk8bMA95ph9wvtMLM26Sq0rdYMvlNORbd05ZVAyBI+O7L4/+qVV1eB+H9
sCTWasEsDB6iM/jm4pVhY1dPgbvHFhJbNdgEF4cHAOag8aqVCQE2xucwEUoEqu7rDRGQFF4whIhB
DDngE6NPZ3xRn7rGqDVEHg65P9KbLmkhqJ+viplVhAkk5eNsvc+6JqylDejdBjBySwW1QKhn1Njm
k+e3CcUAT8GDdMH0xqAQl6X71j9bIUAjCjh9/LXnOu9WLF+flVMJWW5cWHgqJ177Y3hXwpudN+Iv
7vI/bNnvdP+n23Gmmw8q4oVzofkiAK51Mm3C2SZPR+SGJtWGVU9+9wDV0emrKpkNdolsJFdBgB47
1WM65B6uqn6mAVQBkICWFXPW0esy+3ZG3P5J6BMV2JPZ+TOCXcMJJoOOJhckKteS3Tv6vqeiYf19
lD7hQSYFkbexp86FiTWn26aFnMpm8/i55Qg1j3GEsLvcEkG9Yf6JUiUMp77fcHylEpMA67mRm+Ye
Ow69bgoRRXnzu3WOvYb5/uEuzbwkGQKH+Vp2sOs91w3J9SvzZyGd5SRTiTIg8Lx1vLCDzD9eefnn
vJjd4HQqJX3EBdTnZJs0OlaRmHyXLbFf2gEwk2h4r/aLPX3eqQWCXjhsT8o9xfNcpQUjSuKfXBRG
sJHmSK8efq2h8xBpEIGR0kUBq9INN0gP++cF0n1s7VStldbj3Co576dIeDdSExU7I/A5P4bk9Hdy
iiv1rujF7YBmN2fjp/vhDRntG/UACRLvNCoYbTtRhGLzZ9Km6kZ9LWe0mmsZapkICOS6H8RZ4Xcr
qk3RfIRg7/6TIXIxcSz3FYd89xmZhaZNQgh3O+tPP++RSwIWV+jnGfLVi+qrJj28z2XDcP+lE1+H
WiO9tBiLFn9nQTIsgXrKOkJLx4s5Fvcn8AIH2/devoV74gaD588WuMGTqGm+r3XTvZ9A+SlqK/IQ
UxEFideqGlSBLGKXd1iz/kS+nYICQLnCOcfxD5t9BOvJkDyggQfBfIpLMx6cFmW1OQw3T1I8vZmw
I7gbMv38wAXxdVKB7YjXdXqnOjdyBtxLlJCtP0PHdeU4EK2r8tUUqFacGTzaExBsnYO6T/ih5fdV
8XPcPXoohpmqOaL+gHGZMD/dO2JiJwA8j9e6YRAbv/A06Dn3Hr44yS/2f9HDdMNjKyPqCEmLaOmj
CjSIMiEuq2+AEVZng15XVYCBboBJWxKsBfSQxeMdQYJ4hxKsEnuqt0lxV3lcQtGPzecy+761xQZR
AmwqUP7QOweE3itMNA242bnSsBR/wF1VhfOZPPyWIkwYKIFcomo19PtCKv0W5L7Kc/vDqQLqFODF
IX+jtESdeePpGsEiAw5nJ48z5siQMmfkRmYJpELBxh4luxZq+HqKpKNL6Ret4OIwEkmYICeAb/n+
+cD9U4MAtVlt2CxqTp2GrQadER8aBm5lMrrtPabIuGVQApvz7nGpoKflnH/IvyLuMwwQNGWXakal
SustO/ZiViZ7ywyOnZODBfiFFiE8FMcBhkoyinvOCyzalM9fehZlTVd5HWyhqdyq4zM1TE0mI1HF
cCEFOrcdzpEPx47BCY7tBUEPNcmVzEpWpOdf9+8IgITh+LfIUjdvVbsjRnqj/Fr7PW0O4sbrvj+M
2u27Uj9zZihxxOSP8St4Z1Oiq+f+vuab5eISJCwX92icCPDjuA11dHBUMJ29FRpkfC6jEoSCtgo/
VJAhJIMM5Ze2HbWBsNyw+9HQNLSR20OBjf25tGJiKDfo88W+alh83PcJCTqRXargnPJIHK5KzYFK
UYM3Vz+yRzUHB7BVAI50hq0RyQwzK/iuPQ/Ymq7m9HWfG6J12Xyi/38CO83T6nWFLG7WdsWHwPBy
dTjGiTEUAhKf+wYb0vo0qdZnDWooHDEsNzbs0mxuSugTRe8Po7EQ920swFTpflOATfuR4jW7rUB2
6s6E57Jkpn5qj3wtfSDlPc/Ef8YkIFH9GwIYs3LYD2q8L1QyHfV4JMBEMd/UWan8imeJPvlBJtuG
QsVBK8N7LwrzsZqAtCrGmbqNvKy1GjnbFzrTIPuRSLPdcWfybXlwtXNUq43FwpAIril93Lios62A
oMNAFodzgC5Y2RLlrv8XkENgRhmIUOYq124RDflFEDJNwMxESwxbm3/Y041OMztpIF75ArxHM0am
B+6ezV25kdowqDoi/lkOwReEwBIy4gHFiA274qQzjQas0OobI76OsSiu1osW8YIn0EocgNMjCHJ8
PmEjj8QPzJCGNjP9Wxt7Sr2sno6Z7roLK1X3D8hcYVLosbq+jyZt75+NxO4aAv6HvQRLv//6VEe+
WFkXg0B06sgnIutwm5ru7N3VyUUA7QISuH5Wz5ws3yNQWnq+wVZEgWaj3g+MBkJOHLAImt2zl3FO
+S5q8yeSiX9zSfoLaGUACjzVvuS9Zk28fhZKFvNoeNo22CZ+zCi3GjEQ3/eHXObApyTERrffk0By
jHSQ8uCs2j3IKUjM5xB94pRImIqlAp4NCDpO8vHUr7aO/7ckXGMUwPuYVw/25kWbhuUHrEAR3oMP
ZWDCmlP9bQ46g5OuKZmz/tLcYNE/fFyrCf+fcYiVxLt3+jufee1OksxbLpxiTn1YNmz/+MiFNRdi
5D3jx7IAyKZnevRmMznKMkErFunn9nHhUgsuj8WquP3xh/MknmxrRKRWqIAtdwrh0YmFOkzGKRF2
bEqCBrPBOA1Ovb5wcWmzafKZ5TGFV3KChXVxG6UdgK1zzRLjP16WuZ/9U8/mE/PcRGkv/luXEo5C
k668Fnz1s8Do5jWL0rgX+a6RwLpVHq9dByZxMSDTVOAiQdvLOc2D5Hy1rM/xBUhyVVRp1XjQZjlu
wMyEcLJ1dSrf2Mf+wVgsIS0dWI4mYQf1LDuZQibn15+1vGBi3yJg0k+cs2P0YjYFG3GNeFTcrFG5
PrE8BfFTnCACJ2sjmTG2rQ5Icw2WVKtciXeO/4x8ZBE1rf+cf4Fg4lRvcXtbr+0Z3o9nlBxO2POe
985O0gQFaGoJdLEvHkF5zouBcR8bKoZ0HKPF/R1vbo3l2XStuWF7bCwds/sqA4jyDOSKdKJN/fGl
0fDSx0/PJN28GL3IhQacJbaCWLQCnGODnzJzYcPFCFvqaT6OGx/qIX8GssMrbR+L6zrzQ+rGDMXf
Xx5frEfnvtd5EQLpEenZz+GLFLn/6gtbHqx4f4EUylnbH+gUPnL4INKjxgN92GTLaVGQXCgURgna
zPZleTF0T9YzIu1gPPjgjrGUVZiLR4c3F5hp2+1FuI0p6JPFGS2zvc8Eb9aQ62lo4Rl1K/HQKrm0
cDKy5hCdCurzAoyoDcq+gornMj6S0YPxtf2WTWTsiaNV8ILbHv+mdmv6VoaMgAZHkNg3K7IOn75x
bh8L9bHts5C3v3vYnNB7DT/3341UvkfI3RyJWz6ZNX7BWGfqdk6FWZH+LA2mj0KFK36yQv3OcPnD
cfa//gEbU5WPMfm8a2+PsiJSpzA+TTWn8iwuvue4KgrgNyeBSZpC56LR+vdjcV7OpTpw4IkHuWVg
fIiv1b2lwH5pxt2a+/y+mmXLI+MBSLikQGIIY7iNvQ4ob81I8l5ecBZgvFOKclsHVK6Wr2AVYk6c
eqzkyUIO1sMK9ycet845WmpHoK6G+QasvTiw0JkmJ+jIpqdCs8iC2uFMrFYujJuBJLvmKsZgabab
oJqDLvTd9Mxot0nDQi0r+KrJtCVpzLkp1/NBXPZPdRy6LybQ9tMi7Ax+tHKU+FyD51NGbwYlHnli
DdLaHZyDPbE/5Frj4gMTefe4guey16MY6sJoc9qMYZ0T2Vq6uiozrDfJTMoYqQIBEnNFumgiG8+z
8Q0wejDbmeMarNxQCCZCnEfT1nYuzaEgSnYN2NXD/AQrJ63o6E9FTC4fvVSc+ZD9qnYYBqS9K6ZN
lA28DMhiSOpJuB5aRq+QJNT/Z9omXb8oWiF6hwoj9/P/Qv+XafhtEL3BKbr5SZoynFU8LhXD72Hx
82LH9Q5m8xYln7/LuOyAnbaA53tbRNF7hUqoPa97zX1iEIjLqsrz0pwRgsQzQ78H6QIFYKMZ17tx
U400/SZKu43aj/6G1B+OTPm2Gwkd9JV1yfipyicPspJzYASWo2k2OhCJx5S7wl+jZM4a+9UFbSCq
gCbbXCJ/3kg2jvieW2+gNHX9tBrfJzhEEwDxvu30py69x7hTHrKPKOdnmyvTfKGYa3uN1ud7iOW4
dyO8eJHT+bqooYXW83Stjfp8yuH6TKFsKjZRcaIqDTvtL4gtkMgyoF3+BNZSmetaLMXRW3eGkbDo
lkO3sZkYSIbjUFFlt2ZLUHUALwnLFTJ0CBRKr2I1f9uruVgENrTXGjNUb4PvxHbcKbPZoR89niZi
34U/THLXtwtjUFsxwlpljE1UiKK2M5Bw8ZQOh6F7keOD18APuCtvi4bcGNO5JAWga+aJvWSDg2Qj
5S6aVJZMc2uqQWItpgFdVZq1MnTW9K9hLsvQYiKId3apWzM17dQmk8n8UzCzfBGyJYnUX1iY6q75
po8Hj3PpZs4BcXob0okkfcDiQe4EAHVirOV7W1DRGkppjcxmw/D8I1LHCjPzEByLs+Dcxmkxeojp
9WkJy8Nm2PTAfa+cmvdd2SvmY6vU1gFt/ZDymahO8p+TNzYrs/u27rtDaSQSvepD9pcwy3J9XxPz
2PYUC4NiDD8ashQwSjxXrAX5VfiyD6L02WfoR7VM+sdQ0bYRKndU/gmqGszhsTdFa7h6cJzI2RF9
H8UWF7KKdeU5MizT+NamwLNjTfzlfAONLyz/EPR/qrWR76UVCEKmkP8xEfC+LPY8oxhxAqJnv2al
nzlO7CyoicY617As/IAopqd4E8AO/p9DIq4J3kLe7FiuLj67Amy3it2vrUdsdMpEr8k4dX1xJSKs
gQ0czKAiCKQNcLuFCc68vChO1F3xapI4J12qlPIZfqdL7WOueam/6ttN17pssy0UABhmZMJ8O/QQ
eH6vRnsdD4LRSL8IybtEDhIkh+HZONx3yR3i0jSTZ+dap8e41b/WB9UQ9+OA9jgCbwVEDKCIz5fR
Yn2ALtPlvm3Z73mk4jzWKoR+kIEbkJ7DwTP4nF/XcHIqQvI13aEcumnHvRPpLlaLh0PzqwqFmGCE
9c3dJpxCuMAe1mNMIwJbJqZmV/kwR3S5M/W36cyhazRHNUT3rnBlxGw0OWWhXs5Ow9etimT5tsvJ
IDgKCfWVAwokxOpqADuARLAMNks/J+p5TiLxjHFQjKruvdsuF8aGO0DsD+ojwbLgB5E5dxDNF7NA
EfRsZtCNIyEpnRdNDXLAdOS/23U89Tbb/HVbLpNelWPW5zRkEHp3OlSyqfJaw3ivvqylQEgOi92S
q9VjenHByLnTc5YMBuwfIBhkh1grrFyEuaJwieX/mqsXOumYHumgCryjmPwICYe6AvmViKzReit8
RVv/8ZnkHMs+c/7LvqM8i13kyA9jKFga/hRTq3I4MAOSrAGacDzgSd8YJQm24zHKT0BuGw/Ejo3z
kdgjcB9e+4XrKXGg8FKRSPLlReDaAYlHVbjUq9Cej2J7ctUS6R3S9NP3xEZCYHqIha2U4tmI0Ip5
3W5H+sfDyZnGXSMdLWhQ1Nlw8gvWMMwsmAyeSnz+lCiBO9yWS0z0fTA8rnbOhLfTn393R3adk3KD
OZfOgCNf+tCkNjDu4tpQVpmFfRLr1YMSk//nAGOjSzcvX9QsLsOzulexvSMNTXJIAu/oz+rKO0tQ
sYAQuk9VNK7LBt48W+kPGwNiiisttY6DH7DYAlGNQLtBRfVITtfri0pTp1NnxH8kLCi9r/nhJpo3
ofjJ1FVyu+N0lsBCLDJKmINbjkpMS+oVSZvQBER/fz3KEA0QIzAI+VlWEF6rzutbWGBC0UuGbgJT
/9j6VZaUtj17aXLZBKWgfSRSmLU2Vsk7L8Wx4x1U30QO6VJx8OiONfF1hHu20gKZU9KhxSvz3Xd7
cKlGQchp8wiuuITniv/UtsRkm92HZA73lg62O7kAXsZP74k2yLf1DWs5pPAlPJNzu0+4OI9sV3/E
b4JGzJtva5oip1xrmj0Zgeq+Do1swNjkjnGyLKHrWHtqbau+lpxTIa1bmwEsL9SoEUugZ5E8kh1X
u1p0tWdcv3I80gnxJdJ3BTYbNLl2S5HTfSbpDomh8gGJjk9nL6LhWPU3VF0I9YSDZQTcDEyK7mKz
ZajxmK+oJZwiOICxHDdNTBMTzvEvMpG2vktMFzKpr8o95c1AgyFQG3WjhA5nXX3/zTJgzOFS9CDb
S8YcsqSTnrvoDJc8v28hE+ZtRsW4Vp3MF5w94lSjmydu4ZKuT+E46GIxnoWhOqGBsrF1GEPdpVPY
rnC3N8pZbcBOyoW+8hzR0ApxqOJXB/5szE9yARo5n1CKB++RlFtGnMHB+Ruuqh1TOk+HIj6s7RIA
3YaYeVx5L5LNHNfHGS4BMf8ezV3p/iTxFQngBPV0yuLCjy8VY/lo1N+SxYY1mpx0irxvh/2NSXUv
1FZY5xXZH6UgHm6Kz4W5KduAKcZh835mbcL7WlDY0aF4I5jMtulL2rVHliOY5TktO32zV2eumll1
XRa81fMsajirlYoYbVsUFVfXHV/CUhlRKBzfAWnAc63LEGu1ABSceusjY1l4duAmwf76uyU2ol3R
bIS8tkeDSAdLZDBfsFu/gwJCctWAr609J9PthcbKjW9P6b6bx0XEcTUvjoD1jTC3HhydtO+G4ymS
OFz7X9qUwC10LaFJRINaTWIUByLcHgJRVUnTPfn+aD5955tYpT+zlYGx1i4c5hBTOaWtldIyLfjO
OG3RkF3rZG2neE6mZIubKqxLOjCNgNjgMJhGoIv9w8xmZq/qfvasbJKGB5bIN1xKclHgSN6Q3IYC
asj4gQUk1T5pTC1wA/3J0VlHPqJBKfvV9ne/RAmzCugjeRqSN0cT3+qLVns2WPXQAoxyDnt0QbRV
ezpqNB4grFtyezp1nMC7m7SosL2O0TFbqvaOq9CpJ1T7JwBJDFPJrTzSWB5FLYOTP1T9tcGL14Io
BiYMac1JVHMQsEC7abdtC/y6xnGvX2tZsNq7cWgM7LJxvxzQZDsT/zqNuH/PA/KIVmmUHZ4+wSzA
nKrtQcTO52EppISatj/ujLq0IAvlDf6Ilm5u35EzHe0O0jRxB/zoWJT7fQVKkQD6MzUF3tZlDF7e
UiZDUridoU8LakOCwWYQSWdcMnD48h9tXoOo6KAYsLiwiYWJ4gIR2X/e8VB9GPKwK/uc2fZj7M1x
B1Bj3jYnfPk+kWG0RG4ILBiHrw6lvN1kuqlCmFp7sl+BB5ZFQ54UXFFUiDbjbvQUI2nP6OpROaa6
1WQchzhEpXxT5kHn8QT0jmTY52rY55OD0bPOWCbTpvp7Pbn2QGPd6RCBaahgOWV3hVBlPo5FYZbl
dvXq8oOS1FJScY+oI9Fnvv1O/YTJjSkhAYXSd7fCogxZnjT3rNfmqWxuz5Kx+LXaNv0pH+d+0RYk
0HLTX0i1F/nSElF6ruLf65NQmsQas7tPQ4tCdRCxaTPPfJfjBzDsOpvW82R/C0+lznqcXEizzZGT
mIPQgVfJskF4olhu9dGeC5ZSQV2yF8FJpcPQmti8y08howN1915vuGRwe73HEHahLH8+GHtOJOBp
5rEb1/0yYA4Gd/KIjlsRump30HWm6fXRGZXHpYvsi6lhHx3/FBN1gFbzBM2ssGAxFR8Q1AxpPIac
eFPjs2v+OrFoC3KGK75IaWQHeU/5EktzyevJtkclsTZNYR1sGgPn09X4zHTpon4RJIEL/9qDAQbD
hoHWU+jXxRJJ9ZX846KFb2dAeSfe3w2V9zONWEiLLvVLXG1BPgTllHLHEeQVbetiqrfB8PqgQ8iG
7ayXMU6slEET5xUGJAKSy3ZTTeRGMZddz52QN6aMjt6LcrC//rxrRu5coQttgc85+F9xozP4bIYx
HoiyHxU3H7NJX0+9SeQ6wqsc65E/PswJL2pv5PKEuQlRs/0Teny1ol7YOP1Ep+i5R7SOrPeyn1hB
42IquyUUPF059sdvDj3UYL/3RDIiBskXDvymyPkU0UywNyKEPUz4da/sa2tLmlFOfmRuvaC/tHNW
FA4dqHhMp3XbIR3d7a0r7BKUW/UFLrQDrgWR2cgXcpwJyt3GPIk4D+d4hvvHVzRSxdnzj2VvDtfA
+8yqHnD5XeOOb25Zd/FSpEVaj/nflPjRb0cVdlAysNEFu3oCQ/YrzX0ZV8pQbxqLvqrRhQ7yPYep
prb888YVwRZxnwSKtR8ummRi87rjphY2ox+nQG2N/yMRFhE8qiFgUYYeRCJwtqLmQaoizMS1WORv
B+C29wilXw/Qn1qRbKtsnP/SiyLMqrTkDAybERSlHPkjqHRITYx0lO23er5taQsQ/Gc3r2l5sypl
qJfp0nPeDNI1GKBKnyYkFKS/Ztt1h6wkVeLK137FAiIffY3z2eGma5olD3BSc3/XbqiED13BT6WK
CNNRFC/UVKCERM0Px/TEezro4SAN3wM7WnPecpE+gW9L/PC0tUcNHASPA1WI4epZRuffeZ7F4RpK
L77J8tntLMvTnQLnpVq5/o1r1UW33/GOmpu1K2ghQG94VTrfBUOp8SDFxlKFZ5+CmionVfAk0so+
v1BqsW+9yF+Ph4zQ/qs7F1iwhOxnXjZluelJU8Jt01dxRVFYFf7DygNAskjotZvD1HlUjg5cHl2l
phQaoN2f+63UCtrME5+mY64hmfvTRJNTYpV8wD04jO6q0ExSFrMFfwCsiFcfVsb+VFTrwSg/2H5a
yDVZ8hV7zYZT59d9Sd1Kma4tntyUJnMc+zWoGWWreK9HwbQ03CGgj+JTBK3hjIZM/ljsp08u4Sie
tu0m5by3AHo7p0rMNvavuspQAHpN7dRqCcFC797FDgtFVGf8dpwmpn1nmcd1idRy35DRH62RyM/Z
55Ujtg2etrshV5HiiOCzkApNPubMiH+C74yNwQC1+dRcDjJNyColNQXLM731a+Iave/joKSun4/I
97Mpe90YIbMl4zPMMTu8v5PxeUxgCWrcihacdWCH0QJMzFFRTCbs41M/gZpOuDZHGalUItC+VKoT
4hLtC7KxFMf5dBwphaHVIwqfcCRMEoPopBbV7yHhzfp6rB6SlUmUoyz4RY05FE5xOEaJ7XS7HALp
pVt0yL4t+1Hc5Vw4qFyYS/u2EpHKqBx1EV/t9hToWUfEWfxW9Rhho2+B7NuzVD7iWzLa8ee8rGd+
VXj2QMl/JTnPAL+lvaGyVN0Aa25uLdUPiILyWYoFkaFokhsFxZqKsetzh88lt6fBYNZ+DnASgDkM
crO1Z5eHTtyWLRqz7Kwm2kAhv4KL42D+DNnyMoPykr/jH3zKdNDa7SRIlvECL1iQ418omtXYPrw8
4H+HGQsGocV21pBZw+WyRgweRHodTziwq5wbuIYvKkRwIXN4VcUhH4CQjOFBgbnF8+zRfNLtCiiW
ttIhR8a2zHy1iCDAqVug4rSZwLiZjPdjxee3tQvDjRKv/4JPl0baeQPa3Ylca+MvJ792Ve0kEW+7
MIbtClvFV8MSj3+5Vi2YfwdeLbqWktSogTtoiJQOlAaYRtmQnp+r417Lsua7RO7CKEra0C1ictR5
PazAA70E1r1X6QyBn3FiBD/6GPlYA33HUy/3smJlp7km/q59tP1owg26dF5OOz+PRESStq3ztDsk
/5RJLnNhHxX1Zbb23/YSi0cQnHmTHesJa7E87XYzqsUWfjOnIETJbw+gabRumdm7pjIILj9rmNNb
/mQoeN3Qd/fxz48fQBnVxVFQBPVPItrci5vcyjJ9oMJDM43q3X1a9HXQk0umFvVxNeQC4AXEFe8f
5oOw3sq4TLVvZoJ7vqvHlv5RrKg74CT4980vDz87hg/Vm+fcd6lmUbYOeO4YhS4xETgmNg8k85gq
2PGzOvjdqq7eXgDmsw3y/3P9utX94RGxw5997NboCWN4rnnunup9bmO0ua3Gu04K1RZ4s4viX95l
4zt3XZvXNK4yqAUHffWAip5odGljz6rjE0onaj/d4xinchbwVtVkw+3ilyETZWtIxfYeCwD4Z7sa
rJVvqxTolp/16jtLknL5o9cb67DEh6DLpt9HrXnolv44R6U40qGtr09R4elgDedcxsVTeuEV2SOa
Fkytg0isHSFKzDTsNx4wZr59orX6dZzDuiICeNuNJe2DYStv5xt7TYKAOt3R+ssQti8My0ArCYHE
B2krMI2OEnqrsJl/nTLkjVCeWt2K8QoFaA3Fhjbvz4i7tEe8NFGwYu5PX3ymehwaFpXbAQwx/Zwk
vLaPF9qE/ixdNgKaOKSMTzJv1ft4Ve0hH4NAnHQxHB5Gv+yVdyYqbC3ghrSwCUm0eniAq/+/aFrH
QUh8mUWP1ppdHVQri5XIl98HpmJnYzZuSOB1Lj0rxKanuTNd309ST7DPL/0v+dCZ2XEbFu2x/6Y3
T+oUlHVOQ/MNU5oKbqrYQGjmuh0a6OdzTx2l1GmKPHD028oJu0VqsOaB65opQr4WcsW/2wFg9KD1
RhyO1+7d/mi+LxxgcrHT9z3LPTqlNfvdv08dnj6PDh1FDmMOvlfMFU/AxVoIfV0G7BABnZQ2KPGM
WqYihffzYbylLR5U5phmkZHSkrA0kS8BZ2adjSwEbOty1htmKEQBqMYChQI75swUjnk4NYSwRmtW
S8gbdaE1JbHaQpx9VwP5NqBBNJQtnOlhjFx7VgE2AfC3DhbH4PcpqAXkBVJ0nH+e3kOnuR0/jjse
fHNJ1GwOEZwiIFGR68TMGSVdw1jyTPmojlVQHZBSOGnoQd22mwQfK7OTvwWdlPKcoMIJE2gdDx3A
bQ0qkTauN8bOjfxYq9JULXHtLXKkFS5FS3g/JpRl8RzHaLR52ScZJaYOGil2+1877Ao2JPVC96/X
XJBs45g5UVTI3S5s43J8SLQ3YzhAzud2WCL8qZINXSPRLjJq/x2ORDHBZqvySgKP5najbFPouEIC
kEhSyp/TYqWW9FZdFIC/Vs2uBhy553XwsvXGBtPg1PjkXMOsNwiUn8FlVE0T4WE75sfO8Ihiz+9d
s0a1HtcZPVE0tGz7luucSwPb8jb/cVef6T3kNnTRjMp3fFAmOWC1TZoPjZiYT4GNhZiwSRNvVxHH
sjlOyPXIGGhMmBdY+ZNsndZ9JB+FqIhzK6gkKqKvg6Kxp496BfxSnLRXgm1mWyMI9sTscbnaBQWA
uE7K6JPR6SKQglkERGxX5/oB6WUSVJpODGkACQ46BZnD7m64xywK30EsWxeJR0qSoXdfUdXYmnEA
FtMk1ZhaR+gfa8nBRHnksXGN/5GAbjH8mGeUggXfs5Ds2tTiIfxhguul2UkyVloYXmXDx2r8yCYH
y2EvxLG95GzAVsabuFBPX/Q0H1hhS1U15900aepqrE066zQeijhV9XzioiDYs9xo1zswEnRjTG/N
beNhRZIHZVHbLqghaNz1FFRDWraEdcVdXOa7R410ygbxUe2C8B3Tmz7AQDbtHV3U88qEvY61PdJ+
sJm7REw3vP7oiFRFQca6pK/dGNih90waidOErTm0JN8sqXibzBesXUzWq+tfNJxELV755hhe01fq
mrqIbG12dK7K3jtFICLvxKa2DR4cgpFkja4sP+3DZByLbD36yMpdwPz7Fo6Yim2SzyTAMudR3GLj
ma2T8GR0fTGvmOAB+LrIl4+/f2XKWLOGLeQkGwq/W3QEfD2eq6qVG2Cpe9Q945n1TfqbGoTIRZsY
UwG4gQCUhErEXNHGJyq0uJlk6azZWHWWDy7e97ZuloCzEjjDxrdmYMlFQzCoBKwRyqB8PvWg+5IY
smAKMAUV/kQhJOPv/XyWxDnf1+I5iPuaXXkFqq6vMxbKDlrcItTjlEHYO17Bztb9IY6hFW2dQdrH
UOJN2eJ9VTQmmBZJCJS2oFaxFYdiHMdlCOdmVpNOwg9hLYoJF0bA48VcSgzggQdfl1f1Q7xlZl0u
Pw3WVQPTC5bRKP53OsbeSqAXtLPORe+99sNP38o5oSzKKzUi50CP8hCLFvX/M1FjvIotFX2n+CR6
C7zxn4T9sWfELkXF5RbcpuQy/u0Zi5k06GaUMCViY3xWw2JCV5eXuC0u0HUndN2Hk4LJIOy78uoZ
+lQsKt6DiFmC7Cxcz10zp/S220hcHqN7YoHRqf9l/yrzYDS/4zf74RDfuMMbMSYhCTtGSVvjwB+H
nzGSX90ZL+xbrAkmqyRyx3TIufcUaKHn/nAZ/2mRFF0o6BFgMTj2bWwO4QGQNARoBe0NGIfm7JIP
JlSU4UVhOci5P0zaZRl+mUVk+FUlLwZ/utqCC/266yxhlcyz9Qr+KJQAuOdvnsMfqF/oCvWfmoIN
BjQQyZcdA7UbEflK6PeWHswc3yvabj07evw9DUKN9FnhmOqnl0SLJjD3KrmaJz+Qew81IhJHso5W
lSsXRPE4bMFfClmyapvEVwOqSm+nJafhXhwee8AJXpybwYcud4IbhZQVm2yA4xBEei8xdRCSg5sw
jUoP43Wr9iR1V6yK7o7RZoJWXi58SbvvCPE265esKM83sitBJG1tVhy8lR14qm8Q9OAg/7nE3ag8
Ni8IdtiehQEv/yyYndmyqNWjtUn91f5BuQUlkSoO7DlNHeD2ZZttFWnZihXD/7Tk19ziyT++mAUr
eoB4sA6vfNsG0hEaw7yUeHKbaTRohNPThTijyRIlHObHL2XJkLgZc37bzRtxEI+l1CMzpuWbuliW
Flozc6G9gLBNp+A5JE+19zA7+VXvHNcB8tFgBq7+3nisFnTWantIrJUJvUV2v7T2ivU/Z3QA8Tyh
RV4cKQKuWuSr5NsoAji5EFK2QFTAiqXARolSZB297eIXKQJJ59tJd6kz9Wede36A1nt3MIwKlwoD
RPCEJchI5RL5JJvvPpGaqGgR0WEIjmDLb2LIwYl8vlMTe41plENGNFNvR2DNX5IdpIA4Obi0/UPp
naxeVwjjgq4m95LA1sb++3s9ju44fQNV0H1PWpsalc2XJSHz8PUnXwB2jY1CRkBlRZXPg+kQhe9A
BjiGI2jecC1qxvKdqA0dy0x9EHFKlWDKK206aU8YgCx/4tTc4gPEiWMccnsFVVJir0MYYjxXe9t2
zFHVQ9gHub09ac1Dwdv5yrdDmKtcqWV00ZxpVIfMzoaePCG7tZqwZ3S94mIC0Oi5N31YwNU5OiCj
yiU7mp9/vKZpsKr2ONzi8UKnq+wfHLNRMMprtknNkKNSAY85cW8e77BMpiXlbF87tMoF16Tgnm4x
tQfCOSqAwSv85d31IQ+pEanCOz5vOlCogO6IoLkk2UixRLaRDH3iVVOwpUcfiLSysEtz0ylO9wiy
9nYL8mBLJEho7ToU96XTLkp9n4yHjv3baHu4FgMXND2LRwuSbFvvUkRtO/R3vAtwFRIwGiZn9udb
RuQJ7TJh8VDhS1nxyvD4JgFRfnwLO+n6lUbSEvKxC3Cr1PE9Y8eCQwUGIuZK3wKZWFOY6Zg6MSLv
8jnX7LW2K19VHhrFmwRYPG89hUf8ueyzxX0ga+0Y6NvCGmwfE6A3dHSt602TxCyJ5obreIyXWEPZ
C95aFQOFV4Dy6u4XnenUtzURimEyKnSXKO7H0fGhXJrMKwgWSrfIYtoFISkWxYoYe47yWOg3Ej+k
IRQtel4M8DToDza88IHP9c7hQh9un/OCu8z1vnq9iZMAId/Ba80apbPtgEkUzxerBgxLsGpLotk8
4LBC+6/ifJVSAEPWkbb+qBm9M4V+SlWxW7B242vEDmfZ21MgDBeuqMgUYbwHnOwtGa3PyDqKL43B
ztEGBc6w5RNcWnLYrf6W5VZJ5MPjGMxrZYjbrX/IORT6Fwg5XxzE+6oayBt5e/0iQcX/czGoMDOh
s/DOJWIJS6BwleGL9YybkcKx5xCSEr+x2EDayNTmNy6PZfnOGMaF3t5kdKaU9RlZXq+VV+V58S0w
SB37JYz0ZaQSv7GmjXqwySCla8F6hf6/5u3MEnOFE569zVYso6UZh7C9P52dIQ+KX0AyDZShR2dK
Eh0BIhXpuAf8hhjQOcakw2hFjr/vQL7VXCUeKQadtcvKQ5KNAqvK/M2Vz18khUkrGrsTLdzx+ElX
I5L6PANJcGHHG5s90zvy/Yaonac6h64V5tgpMezzqt4kTvUnD67bXx8RofeAk0GJMIpi+9fW9buq
wiFS8FrqZxQbIIsIScfYodh9PR0f+U5UFJsSHcohXrXTg2PAcXNXqe0GFNu3qXm7sqokImEw0IIv
jUIDCQJ5L8krPzMEjPeArP8Iku+o8XZ/zsZhpoHNm3m8ipFAUpbc00FkJ84EUMGsrnUcLV2PHTqH
O/wkGsNBx3tdq4RBAbSoJ4ppwVoAEZdhFk7ollVk0TbGIuwAaNvrzSaeAuER4LGCylGaVPlZICKz
r1Gfz7gfKTEAiJrtUoKh0us3GKHBWL2n634vmKQwtraMTRhHkCYQQppd9xz7pjXLRRtVl+FGoMiT
XyQ1pxXrpjqCZvVDw6h0KQHOcInKb2qr+30d3P57fStg6jk1B7XOh1m9GTtG+aD1VE3TgBju5qjJ
R4PYhNknSdZIwdKetAF5SLsOcwirlk1rUpzYFsoxRq9JAeab45f9xYC5TJ8/RkynLPmxpo40VUP7
WFwJUVdJvZqA7IofaAbOBrmzB6NTFq2Of2SpI5VvQDcY4gQA/RapD+qPZPZ66/hsZW/UbQpoW8Tu
1lJUImKDZ+l/RoQwCJlVJ4307sGYM6Y5ZI/r5HlDQviIpoSG+QO1RP8WUkhnBDwQDNK9bWUUFhfg
IRO86D1CW4BwMoHHbDvc1Nuqpjgz+2MBvRD7K68QoJrofiGBjCAGxwFT7pm3FpDjVhApLgDNwIh0
sCHRkyHbRpU7Gn02T15104V2/1XHwk8GfGdul/ii32LLJqnt9nu19UsjwuPXw0CUvqMVBrZAJLW2
AKfg3/lzx4JYsFemLP5CpKgLWHSrLC2Vfgjr48jg0t5fg5lUSdJ7/U5BdnrZ1GUww3WnUYekSLOC
ycCA94RkAA9woAoBoCh/M8/TE24x/YluuPP/f+XDrI6fx+kxMgG6G7Xaxqw1lnaZNGfhTAms+pMj
IijfHdXKvyvHHTLYg4QMMV7C5YiHYxZyB0p/pkJesyz1dIYtUimsL96Op/YWzkQJFiVR9MK87djD
zN8lSp9UNoWbWx32oYz4itUVpWu+JABiXw8uikJRiv2kYPVQJ/XNcslzSeJ2HOo43b8wOpEGyz5/
tNCacVJLOICSgu67vzF0fs6lbY64o3fb/MYjyJcBwpGcQfCk7/ZbLU40/Omqjf0STx2jRQQ0RQlw
UJEzWNCQ15SsAbQiwgXQTSMD0W55KYiji2nLeZTtcF0466F2lIy+Ew/xTCmtPwJVjL04XtPlM/WW
GkA4mzCcIKGNK7OPQZFFMB/lUc5Oaj75OjfFttVpEEiUVpI7lRzYtC3y2PpoNgs1M6vI43Mbr/6j
0MrEkfmb6ZHbDPxqg3uc95ZVP/eslrbgsfeTPQ5JuN0X4/cpuKsg2hhUt9CiN0qumru2OR0t9nRz
IAefan9THuNFjub346XUjjXJZuKyi0B2anbVoXPnmS39cQGoFLorce4On9mxXwV55M4ZfHaHvEeK
J/16g/rIY4SzXaJZCeR/HYLCclOwDuGkOWGrqzKJa3zQn+heBIJIs9suocv+OgfblZKdfuQuR3bI
Y/u9IwmAXc3XtpcuD935OpW3ysU4cO8eg07vE4gTyy40zDzxuQNYaEQKTSdHS11YlZ3jl6wigHco
n68QLqERsGqyzc3iTxr2rVjrNgms1NBIyk0X0mLC96j5D55ti+28FRTDdpDlST8t0rLmHepnVd6P
jHwZ7S27n/pKS9qUBB65qyA7A7ka0A0WUNu969VGt7wWQxewgTC2znjxlJa5C8oC5MziBuPr4VVy
b6atlXbVXVhPnLMKbrIJIIpIccG7Ma3oQVH5ylWhjzy/oaUEwCfCjatyOZ5aUlEZnuK8f7invO5P
N9uY6Z1iZxzDyLJ/LvNGwLWMjQ9sT+6Xw/L4MYPng64XBFh3FwHLaJG9FkEJefNCYceQKVKb9iD7
1VjO89SotIIyWH9QcPoNO3/E1P/AC6v+pJ+awY1vgz26eLbqlNWzq8dF1CBcIbVh23ENSJTHLxYc
SGiyE9o5otZ6suH+wyKIYZrDNX5kllIfv7lv7B+7sLJ/7n2AZp92y+roTfzVAJEp/eC49IX1GKIL
GFuPsIhW6tA3TM16IPCwyPndWW3cA13oh41upi6YYE3dprg9H2KyOAGIJ0hkV0cHE0FC9PDfCF8e
8rv2T0w2TEPHnx2E1Mpq1Dp2Ylt5CtGLY9hmzuw6siLOxz1tnguH9fv6L895Md+kwiixTlP0Oeah
WtNKusJSI6MQ5c88jgcvZSaA67fkPohKL7+0T+lnOchsNZjiANj43gZ7+VVLlo0UpqbnZdgt+5uL
I6srPsWfn8vK6XRD16KnlNAqfVH0g+CJbTEYEM9oI1+mw0UQywsjD3vRqU0aPN3FNlYlrWHYYQlp
zinglOqCjF4nYARiYyngpgsAG4E0t0zJTVBz9SKqDLPKNxAQymxZArPpJWCeFXy6viKOS6IX8Okh
4Bzq/tOmGoWInIwSBTusttk5a/A3mVa6FcjwRE9OioD6vApBz2eJB7xura0R41/ahyXvd5z6fEg2
CIePde1JLsrVp5zgDjpJ4CHBFErhBpMdn22hlDdVcjkAyHJzarueq42B+MAA9RXbOWWQUrAivfvE
z1ELreAg9m8gMwh1HFGicHLpdYDW9/3csnWmj3oZw56Lvs3kbLIIYjC1Gzr6vd8PUaHwF446yBnv
td9WNg6BaKilBmMhxrPMC0pp1y7+Yi3znWYjba/tgO0qgPD24AHd7hnGoZPXR+WXcwFPVbzS4A+j
43i6yLvmMxTOjkvgIbgQh9LRmtElDYZExzxDGiNuvADfnsM1daFiwCVGFrfcjQn5lfpqWPJDfUHi
MDzj6ptzn5lN9P5W1cwo9w5v6n6cRqymmntC6Yk0ztnWic3C6wRSfSj5RcdMfCZ1qGX5J59I6pCp
3zA8OR0YEjK9zCh3ChFAqC3hFTQ9YthXXMuzZT5UbsqJAVK0WE73635Fam6BqxVwMr6F6ptbQCdO
xmZ9ysb9hFBGDGu4YyUggNgxH2BJWn7Z8qXIoWotvoVRD0hq367bnnjyPSKntSLlMTUUhTzXuDtX
+HWt27oV3kN60VAnr8vtAVBxUdK3zVKo7leNeOo14iHfn0c2wj4KcF76a/44WBAFnWfJ/gHHbFo7
+AXFD5u7XuWSCXvX1dre1CBCU8F3yT71v1gCB7eft1ABgDPSk3lm1pdjkCopjxn4+dgxdKft7D61
zhpBfXdvKzXnH+JZWMk6dL7MZH9q0MLt1qrhqXxnp4vgUuBHtODVG0F7eGVRKTijvAuKOCZ/ntc3
Cp5rLd1anuJshMt7NObTmagCAiMaivQa4CUNWoVVOJFUQhiWNwJ0nEtiQaW7zrkBAggxnKrjCgqN
jy9VvHmobGgNt9msoP+XuRWVJ6gfpZwBneCOiVdqdwocO6PEadRIAvof8js07On3/9prNkJLEAKc
xKxS7M2GfcdfCkBnC+SGJM3WLInnAh7wVkVVkgc+5FBzGHuA03SkYYOs2bk+5clBb6/xL+EkKsBg
jInGYBdtcK7KCyiKL6kMp1Nl1JCivzhvXnVkW0BrMYuynPx1CAy2IINX8vWcZkKpmiv/aKR1i15R
H7e9pMRK1N6WYuyRLXp2spRZSzjgx3TS9YpeTvj47H4Yu8Kq5AT4tbKkCXf5JUbNB8Y5RUVlM+Na
uyk2s9cB8dNoVZwSz500HqjY34/vanD9/TVrcohz++TZwOdwHnji6A9irgWW1Yvg43hP57s6rFd3
EpA/ulGkp4FiDu5o6VDsuNJZMRf1+mo7vxjBlTgvOvaBqFC0rnWgkP9wh43qH/Fq3L0S4J0yad6+
S6LLF4gAF8cwoI3eB+DTMaBqaAOhbDoF09pVa18e+6g32KDMQpAL6nEtu0kPsd+BG+qf53WC34ey
4HavSmVCGCu0Rzy97GUKoeKTPNRtjVKj4hOuDUKd/VCzSMBa646L5SMEDUp+liDNHr0jSd7myHWF
SnfdADbWSOe3fh2UPERYOtvwMFUib5HMidh3FdtA8HkrZxv+9QDmg28VL8sbYWO0Gasn0FLzy+tw
dQ084Ix/z8sfDSK55kocwfcKKqnQyRj2BcJ0m22PyL4QbqcS5L40+bMBzKpB7FTEu42up2Y5B3Fz
MXbqLvui2Xfuc9JOvgzj8CdBQxtl4n3Mjn75YFrzQStQ6HMWAGUYbGLn8XQ2Aph2CPnNzG+7N8E1
xxsIwjl3PUUNE5AGqKhBCqEM0YeT/4cSiBCjHbvSlZz8gm4kGhbgPOp+Y/D7jx6bAaYGHmT1BZIc
gna7ZgVLkU+rEZkuE2E23ZePnCOsDTcnDvgjHq0oRRd+z+7Dff103NxMi3oLztAJiDUF2wSueIVP
/Dp5aiRDPy5RetHLro1nXlbZF8jj4GS6xIXrvOaUVUu9R/I2cVNqlFo5FHK2912HpCHwC+NWaqFX
Imo3emMVR29MePUMnXEGLFmpczwcGj6QGsT0gqoV3F5pJedm0gKhry7hNS2uTWbOzSs4CC3ER61y
XF7heshTUbvoDL5P0mZQEV5Y7YJ1XRkOCBsJHeCQ0AR1WoZE6js/ZItTOqSf8lXXIZbAXjSM4nGI
nr4s6FpTijAciBCXdizALhPoW5ejaniSAGr6pt/8yNdrrBOngGz2yiKtbQUH/qf3F+H2Q1x0tPtP
kuHJvo2CabrWPEz3D9cJyqu5ofIiT1fjreRT1fkAtqAKdvuq0SD1zmgnAyTs1BgfHwtLxci76IZf
9sIb+SOZOjDOKXG3VideAfTB+lhP49tjAJ8vl+KGdYDGpaHLkFZ/sj2iUwGDeAdLuJh+qsapzxK9
OOJwe+9H6y6+/RnPmdOGtEmWR649FsOg5zgDeYTosq1H5CbESxKNWReHA9E+f4IvOFUKtQTNbAji
z0wS5x7N4mlhHWBf4cZFhA/0dgvWTPenFBuBZXduWbd8LpQAMl64YgrJ7Mw9J0on4pa6QM7lr9qp
ZarcZzSznndyPCnlk3xVOg2M0a3UQNrEwBDDu/88bVbr+CJ0zps9sq+dsp5bHFRp/mmb5uZOONnC
SeYfEYG/mavtC02MZOxeHtgUjOiMYBBbB+nfWhQ55Vcl5BLbNYbBWdBi56wq8gRf+mGchdFmK8v8
sAiEvXxvpdNvXOTCRix7GMcFPEQQgssUkvUE6YeMDLCB0B7jH3I8FEM6CuOmMo808VOIN+HryxcA
n5gw2A59KH1cWyQ4NYQdRYQwRSSKG1D+iEXGK5kGN/kRlNkN73GOMdzl1Uj6gG+WdTBR4m3W3uUG
41qzWPs9iaeelKmH1++QqchuhyaYsCRWkHu84XAK5bGdckfjlXYcFvIIaPh4Eu2OMdlqE6zhTE6q
+vBKxXQIkRx8I0AM1OlsQUYXT5wupHGOP0IAZ4+kA/PitXWDRafdx4UtBZSVZCJgl8CFAB0sJBVU
q9bX2WV/YHX+oh+E9sk6eEUVfNRqniflPeMI7T5oWzqFVGe8hai4auBxDXs5ACEXCvAP/MnXyDiq
jazuIYXZDL4h/JWewN5ec/jP84rfhu3OyoKx7Kfl+ohgDdNhbiEisUcJbT9lumPL8k9y8nbbGPk0
Lv5AYSzhHf9VE0tDlPU0OJfQPXfgCBQiOOtnPHZMykeNQ+jGvUAr+j1XbvUnszC4rckgkaY4kqPB
YnVydHiIr8F46HVViAficaXgD7foLAilNoF6eft0JBkpKPPfYdKKX98veB7gQyQihsy7+qtSgdZd
GzEoIlDGzqL1pLly9+m05qL7x3tMP0wS2kfnXxYGPpwp73z4EZe+wMsRajTN6pHDvkDP/TPOnhg1
MqebvlRowTjObgskYBYDODM3sq5/gxXjIscQf6C23NLFQzi8cXBswcHbX+peiehHsFkQUulHMnKz
eoMZSBZ6deISduuHbNJyn/cbwoo1BuxBnAdsUxWLWzDQIjtLO+gq4zUxddy2uPsfo1T+aIarHirn
+SuAgdeJC/YejIbruxRruyDeYwdsoHlbwjDkz3I1bCiqhtRT5LEaw5qGSpv+n8slk1xauaX3bWFB
/40R8Fc9rifNPxLBI9wLwPKuCiQUfS92Bak/g8GHKEFM7nKslPp9zcHXnVdPz8gl3nAIPWpc0kOC
hool1gR0tHRCoaecNVeRTdn27AzIgVoiOPlsd13Xzr9cjHIXh2Gc0L5XfyGaRGscoeYgMOUU3Ufk
3he2DmglTgg6KgQCKtG2Zqpe/gQ0S9LYMwNh2RKR8NzdaeW2tGuQejAxbUrqSmPqxTvU2Vv3+GpU
z7KBibYIglbg9cbyiteKAKKPrkEdjO0bJAMP1aj+Ok+szK4q0ynM9zX/pnrCDGyhlim4ZEq9dxE2
JDw0VKyFdJrqmZPjn8ydjnnFGBaFY8Pmvm0wXeqJvxQhGq2QbfOPkhy8T2+w2cQrul6gU2FTVq8A
B0P2pbMSoHpF34CsBD3icVE41sa1DRkg8b1B0NQZbefm8JcOGMflvrjBemW6e4Z3RIolDScrPFih
eQHSX4mvsDN/JUHI5jcZS701OfakRqlH7Nqd/KHW8HwXQcSnax8hk++m3JAWKL76gWh81ZPT0tTO
nsoGe/vDrJ4/A7kGyOOvOwEw+6+ZKtJBguWhh1SNWO5/ShYFqWGFZtpNO++9arNh/bG4I7EgHEBL
zA+3qzLsPGMZApA4zBOpNeJCzMh+XNTtCedAIXRNeh3ECJXxykMx3Vn2G9uuIxm1tldw+Qmj1fQB
fGB3EFrsokSRwOV/6uXwry/kim2YhO0esElxMIFq+iXtZu7QMts5YHr+CVRKzNYO6JIUJVBjBrNF
gbZ1BTZS0ILjsEJB/UoKfVbMa90Y7bSkZKTVTGM+iYPexHPhJcV7wRNr85hBaLp1Ee5R1G+Iqo/Z
ZuTAQWDkAg/q8t8EeGNolGC53lBM3KOhn+AZSGaftmsn25W2c05LaB0mZOA0UvGL7zlp84kksbbd
UbpjCR/uOBZHUrlagVfye1BTrdccutXuhW76hRReuCmXd3P0Bl9nrKApd+LzDbd6O69LK1HuIIpo
X8nv6AFolwVaGytXTyfNuu0WUkc+jIjeJZBCGp7uh4vIxJBx44vVTD+6Q5o+xLCHK8nNwPZZuqDO
8b1AJ9ub7zbx2PKJX0298LcRtmKCTwpQjn3iH7Ui0Wi/ldLvR37gkr7Ip4qgCy9A1xohWIPt56Q0
1XIymVyBBmKn9wgEeXokO6cVvqRWVvXLOk2T6OFlIzwvKJ2oLtBrl0quNGgymLxfmXEULesptzUl
f5ofl2e/MBbSFB+nziASUJF2vQ1Pjg9dUv+kowCVGrZUAuRVGOLUz4B8+6P9pRI1/bnHDyX/M0bF
5H9jSEwjFrB9tZIhnXPHyzDTfcdSN7XKZl65pnS8WYg9LCalumPS8VX6lJ8mAwkf9Q8bgKa41bPR
f8a6YLqco22gBqn6WhKZekMmzAzlMQTOEnH8/XQKdFtUDglsupuaQQdvTrJteXqRPoAYze20Yew8
ETqymx1S8tY3mUoWJY9ny1p40TBK1KKXqVo55BXpcl3RhwRlkbELsgQ9kCdkC9EwBuFaRAu7ESBU
tI537WD4wGn/RjRJnvh50Zl1ksB9VHM0cfgNaUqFrQMFfu/7Wrkg6ABWgIc5OjDp917D5NDoZWay
AP1X8GVj8ha3YygmI1OVxrPZTmnYqThiouaw6JrJrZCa94ypT1Jg0aKQHA8R/MVFpWC7keRo0BtI
AUvSYgXc5YnqqNWWD7YnuBnZSp1upNHs9y49cYhtW7lDzFSADR8andljiNR5MyL2uYONWCZuxg8O
Y7ag8yF+uPZT+LCOqmiahBz8GCC0miyD1001yetruzI0e0w+nj7BVfO4sbt9aBzAPlzOLbpSfWkv
lVbhuc2r2vpGZ4TwtfO8jUVY2lJRIPb2OnyC1wxfA2NAFuXC33lDQMM+rIy12IAZwOnpMJUHQ6mm
aEe7fjElW2PlSIFV69YQQuC99qtZL4H5+EDlvsYcMls2CTi8SJNxIYmq0n0GXPBL8NO5vcRSUyBr
ir/DPJ8MALaATD4qgXDj6BqZ4eY54G0dI4f9pbb7VPJU0PywV+fGUEO+aBmGNJazFKLa2dVZCUgS
CHT0BiZnBgBOckEyN4CQXGw4tdvvsIhhrfrGQmh3qTltFWf/h+iu1EPBrLMopWQfWHnGhyTYfSXD
+jBqc0irU6mETbtMgA77N7vS+nUc4w0OcCwHQJe77A8yMblAO1vtphRwIll+YJYXO7SX9Xk4Tq8a
aLm0VnzBVFtq0rTnCsQbyNE0yJlTtgFbd/2AlXdz6abkhttxdGmqqwHUjqK+Qly1sHmsZnR4Pjqz
4Ve9HO/ViBIstg8+/yji7Y6iXKCAkbM8wvNpNL5ttC5Cb3hc+mqoK5o9ykkk9Tbsnk7Z3KUCkPzg
J8jQV9+otlOQaQENC94hStYxmGVgrXTuQxzvFi5D4VrnA2OO+oseVKpT/aEtvZJvUAjswEm6veVc
lp9r1eQX/0wJEXjmU5Bk/7QkzB8Mft9CFdjefVXSiJJ9egMYTtyNtxmd1a21pjNpgxv9D+DeoP8y
Wg7yxGlXDzhKHJ0avXFoSOjRW7OWFbjbB5c3p/mv+ERQnH08e3lZak7ugZO2Ic+iKmWj/elShnhH
sGlOfAY6rK4iThu29VGtgSpcTE3sXpXMyiopjAlH4s0L1/DeiCL7KyBrIKnIRgl1ZL0UcD2UGqym
PBObPsG8c6j1xx9qXe3zlnjNc/cNg5TRkv8H1Kyj/PXAh+MBloJOfQnyHTKflvixRB3Aef6p5DRb
mY6MyDqNeLs0hR0jOdMO/VHec6MTSv/VFjZ+9Nr/36HA5sotztM5kmYvTo+WkWb5J0/EhOVHmXt+
2jaIXKZxEojgoMq+7fufaso2kNL/b6ntEWyE090b4h5pfYYfV5LLxqLY7EDQQAkCqVKacIlqbkNr
U/5EAeGsbncSWHI4ZXP720djt1sg7uPjWloWP8ieE+lOtc26sDazlsx41vbCPkKL88ji/ebU8rmp
3y7UJrgKWPIdqH8VtITzeKUJBxpo+9mWvEPgCOCthp6r8+vp17Q5jaEOWDiEB+Miv5bK5wFJBKB0
xAbwDvMPHljfnLhsE8lXv9sCnAgUwA+xdcX6uVOdz/SlHGxTkljM+rsR/92m/wKH7/ep9X6jHlg1
7KV6gk5f6PeCSZ0WCFwcR5CXU6B6ueXF7SqmkhDi1A9GCIAUBMZjJr7qpzMkrYshFa1Y7QgyvBor
h5ZwZMyCzbQPvpmM2/G9k5P+auFKIpIpZyIeIrDdHOE6sxMjVP5YoV1cRkPfJzVU3XRs3iYDSF/c
3VX99SayOVgWmmPEt/e3vyPl3HarubkgtfhZEmluZUK6y1v5NnLtzsS6Qa+a0JcwdiCefae9Rwok
gNw11Ha5ApQmRnodOSYLhYDvEMER5errDc/hldZHxNtibh3ccqNw4bPiI2Yrhml9Uf375Dcwns7p
50wV+AnfB3Hko6OZnHc866vhBYKMmi4yhFER0VSBCOi/77FVdXSV/mCPtTHCeLUX6CGR1cmEedsw
LeGjl+Cx/ZdnWvSbqcDjUVi+ZrSgTd7kqOKvq4zu+wT3aKGEEdZWdq9uD4fyjFj+I5qV/n+G05TB
0fNbM+lnPJKS8+lV54XrQic87gHVFE4iW6O7+ZMU9EFIGOPGmqqe8rT7jW76o68ckDFg/hceK/M8
ruTi9noTMdAMhLTO9NQqUfjYG7jIHVCEQ06BfFE+pwJvDEr6MoGwVX+SkEMEOppBpoMqSKvXMwMD
m4wjy5zHG1BL3rTKDmklIXJmNeI5RonCjGJ5imsPu9pvhgF+lkq+8Yj239dHeBy3hDtrWf6QCnTS
vbAeBci4kyqhDWTVoL7qOM2aQTUehRedFQv9IHtj2ij36XEMDAuHGI7hdHPFJ1to+khuESxlLFMQ
rZ9S1hSXZ+jQL8FmjyZFnbNrNQ+iEXQmX39izodM1tUKruRJGAHiUSAwQ2UjPl1NDLLHtq20wtuz
YQj+WNfCgEPBQik3CEYE7whSpKMrD0cn4fLhIC3vcQaSbe7fX0MmVYyJxRlwW3vy/ylH4jSq90rO
75JCdl8FWW/d7L3htZcgDft0fSZsfNXZiNR3lgiAV1cgFtvoxE8IuVkMi2zd5naeEKvrFupjTzga
C7LfaI/txNEJYlp4J75n8nvIKMlHWyIPV7IoYXUBbDC6qEGqUBwJizu57xrnCxmxTqOFATtiXQRh
E81maebFJeiU+wmAFxdDHrkcYvIG+wE8RDRPM6etEP7SLHJDi+g/2I49yPF3LOhw0baveBCzMyq/
2NZQ8tmcfLI+Jsk6WOQC+1EBTF8+Srsmb+34F6+REZtQbdiq9UDO1ZR4h4yqPBFC0pMEielpAviu
TB329CD8DZtTyzID2iS3JJU7/MQhL8AyLGjs7Ahy2lav9hn2yq9ZNv15j6eTHUdmsrNofbyCnOHo
TKILxaCUofBM92qM4AkJtQw9h/LGk/YE3Qp+VzTZ6KDSno039dOqgvuka8l5utqrhVSY5HYu7tpV
oi1RK3qJFuXg/sPsHYZnUvkYyV7Hbx/8KFaMTFCGc8rtr9OzN41UGhjp+4a14lVnP8nrTPDn+XKa
3n725glHmBz87xaS7g+tEzIONnu9p381kHYPXVWRJV3DZwoMPnPDYV3qjaG1q/fqEyNbkCGpG6wh
XK+UGZS7D7ikQiTXcDAbU2oPOCBYdCdYQd9rgXmAtgILkT5XY+W+aq/y3Oxb7TuphJ13D4aZTLOm
vPYJOcVS3muYwLF7vwFh31ZalwHPIYTDcYHKAICsFRS1/Xau62FifgOtv4NN4ceNqJ+UVDmPWAPE
XEXGemlWdby/u9+EAAJQJjRLZvqC9kzSKLE4vUcF2y8XgnWS4SpfFXTY+mEoS8uEEVGeIWORSRmt
6GiHC6qviV9otRVKxC1NY2DadSO2F0nfSZj8UU/gkh6qXyvSOSP8xIznfShemThcTWK4i5GpKnA4
dQkNtq3THuwPj+qEjTpG1oWsKXUDBIuuW0NaR/bowRHGO3XTjThAJfTImsw7Tz6ni2qARiWfNrV4
6scX+x+XTBkbJn3TMVFD6M/AoZDh5yzPaS+OI/B8Gc10qDIU+vjOvbdwHSmOzmTLaSAgetABKaDV
OihucF2Peud3aqY5SVYLNdIhBUbAoCjnUr0LHK4mhzLThvVWMykr2LbImq/5FxhheS+Al4QAqbDp
AchZNm4Kw34minTbqRoyP3aK5t05q45D9lDXByT0PxRsjaojtShnt2vHVxVlix/LVJhQDJmqZDm9
YzHWaYEGG1pNVYbuR3Ej9KE2lkWBIZ3/RlXQ+T+tPfBgOaFdzDBnG7bPp4ropeiCT1u5HNHR6yXX
/U89Mu68FAnASNF1fE1ccTgik0ahE/7g7FQHBkE2HDhvSi/+pktk8P8yg1SUvGsBXQB3qn5csqfA
YZyPkBWnNpo6fqN6+5Y2Zzc3GP5vyWCdPJ3JCC4zNq8OJ5JF3awtWNznt5NwF60Q5MMa+FRM5drg
uf75BMMO2U+G6WnWu1WGEWNMiFROkDvGuBientR2PzXy/9+P40E+fRTtg9lZ5jjdyohXlMoMjJNy
3uHsHSvRWefuWbjZem6uxUPmX8J9yGmrQwKXHGIm+CUi+uN7EJQTVoHVUKySQEKOkXwO/WWXtDVs
8y++egJxzJgPbTEbXrNz24+SO5qQFfNA1OZZWhXCi/mMo3IhsflZaHcbLnN53C44GsvdQQg6tcOK
8lg9Os0IyBfqN0CGrdIQ62yiEqqN/SMNhqMXw2+YGeBEoT6iG78pDgbYCIR3EU5Hgr77czmsvKCN
Os0IE3SC3Oo1S/NQAJilj04fRIowvNSw13ozuDJqr1r2CU3DbCTQcu6AnJr6fjI/DK7wb+2S9VcM
iDylP5rQDwjBRCNNpw4jBCWkPS9fnjdHJ9krpa/TP0Z8xyMv0EJdUgiGSGmXT4KJqH2IrwbV7HNO
JmTb7VUgquzLsc7wE3qRV86t9nHOSj6+E4jNXk7GzxjkSw7bkBOUNp5eVPTj8X9ZXN3gUyidlfqM
Mzm5Yvf4TW1Wz0Psd1FjbUR1WyWl+qtDLk1o0dpjaUoh2dkJ+nPyLBcWy12UnFUIpNWcKKmQEy8f
S8g8jqvURAHDlV8EHkyb2Nr5Crffryoh92TiGnzo32O7ge/+3e1i3JDwYaFk++8B0Ol63NEDQ8Th
ZcovKgUVTyNFUW+xVa2HbWHWTEB0kLn2LF8GdzCK0WuWrbySt4tavnm3muU9pzv+lMOA1hbIypaO
uG0mxEco4hMSuRUwGORJOrkcKCS2jNdjNwZ1PBn+Wuf9WUCw2dOktT6clpTu0VKlg3TB7H7JtKNm
wPF1FJU+sHKCPUgdrEn3abjw8ygpsnQQUww8eHW/c0ZP52yjv7IrfzLcTa4aEm9i07adN4qzEQcQ
SW8Q1951/bCtAa3JveQsDKUpWMm6pX4pUZPlW9AJQ/NIsNwvkLVgIuMqUBZEYvBM5OQzzApG17nQ
sJ2+uKo9FzHJuKEpvV+sYRO2wxcEM62HNQ6ZMJZH61UkaN3BxXo41iAD7IGwNyQyw8VAUlXuf/b9
19y+Dv7LU4vRAvdsv2CSZ480/wV+fwsWoTjenTEixxbXuIfqhBZGvgkkeUv+nKxE3RvfdIV0/z/E
TS1WybXYCem6bOZx/pQhEoASjfvMaq7knc9+XByC5T0gzVr1FNfezTVjU/vyI9B9F72GZh7mgcoU
4IfqzbmxV8ydWb4+iQ+VvIZSrZGC8KFfEtNhygw8rPu0eYpbKM8ATsFzQ885AnHOU00e4k0JCMcD
IgpT2POyy++/atVPM8My9GSXG19ymKgbtcGH2Gs6wdhnNrqgd6SKnzkT88vUgWNeaZLbc6RNeuX0
pMLyzmUnDVWRGLbG+aGA03pvAf34NMp0Djp4hcJC1GKsr+M2r6HkBOZzL67uVVnQK9y00lsle9e8
ScQrI5AREjJ1cD5K6U6fk+aW4E/hERNJao3fbDyqMCsVqCTYgdNpVCQJKtCicXerUaCn7hwSHskl
WA5kt54lY6KNf/sib2DAL0J0QCKjgUqiBOviNT5POh00Q9ZdsteN96AXR5i7opjLYUhQtAb1I+VY
OiVmz2dzrgzkn2Q7Uf2Dzxuxz7K4WyKSxp4SXdPuWQCB7QGnFIGgYxGx1747i6Rtx2PamA/lpgMT
/62NUCTuTGn62qfA/9Z0vDUTiDdOIByZqP+taV1nueZXK1NcXp7won/ogW9X29lh9avKhfePjcrC
Mpn5Fxuw0nrp/aSgL3ysUAEJVZdwkZwfl+s9vsG4jCnVb3IDcLCCVDDOMBWV5TNWLt7QSCaQIQlo
o7Ty3d6dPs1B9nh3T2y5RCZsaTBUQP1MftKnfAMrrXJs516KuRr/OPIuCdTfRQK68bPUdbxhVfBD
7KR+MNaVTouVurAjLrZedY2JZAbOw6Xql6nwkCqmGCdcKijrrefsP1UPk5mURWzQ1J7wmdAHgNYU
y7pE+tC9DFCyiECufGyS8o4G+E1nEfYeTpIzbXPlwRjEzaDiLZgwA522/yV6vKKmvHGrlzVuUkE0
V38alciga6BHZMwHTGnDvKXBjbath7zL4qJpFErLK5Vsdmea/h/8aU5WQ6OLvetc6oP6XoV8J4Ux
fTJDbhkNIobwe4nu+c85kjl+6O2bM0vYpTJqoDVJr0v5dEP64aPxE+UC2XQj78IUTRsb9MRTE3fx
jB8BBER6+SYjGwv9GZuiCW2My+vNzGX/zqSxr5AiyVGTE6VfJJeXZtY7uMROVjnVuShIiS+ugrpj
QCY3OYGLZUenXLmB0QFh4GMCMRe6cLz8b2lTXX0Nk9WG+CjxQEEwSRyvpRBVz89OBRS1/3NEXMjU
XE/O+6PbmP3RWBCX3+OHFpxjN3XnV6o9v9qqifMKktdQrIQ5//UKXe9Rc3t9ag47UtLWIIg0Stb+
xtYjREZycoDx27OtWK6SzqfI4+DLcqrpCvkqNqwoIzEPW/MNZ0HoGe0jdIqeT39TZbp9i73BuJxv
4lbWwiEmoDOZCRfhVkc2d6P4MZwVmKz/4lJIKWfC2gzGzMEmV56aeKz1R918ak8fLHJTaKRFBL8B
cxTass6NIIVMeX0C0YYBCXX44K2y5XngUN3D5cuVElz94Zhg475oKmNvGTvtgehIRpXO0vAWOvTJ
RaHnfg12n2G3tBasidW+SA+zJ4iLYx6ou5wbmI/hnf/QaPY/eTABlgr55N1B0xb2HyK7+uP+GWC8
m/IHTMIcV48r1885rz7EUkNSY5OLEbDI9qa0Ovpq0sSqY2JnNxFM9RwMQDtSuV+W2uGhI7sbIT72
6xf+ckxFlVYouaBSAAwlEAK9KJb1WzeUJB6YHFdWLoRsLBgjCcvxUVWbBWSeuHdFOE2YOyXZ2k7P
50Oat36zPGfphacFOwBQP5TWT8XwbS5lWtPxyfEn+irH/UouJm5xn7s8H10yb/w5dNKhNhVGiH6H
usIDG+kece3AjpRMworRuMXoped1Wwot1XrjWPNCnN2t2p9sd5xouITr39WxslDC25nwAqcEzh3e
weZpK16FQgNPzMcAf+tv4tYNYmcbYr/sgrnS8nxcZw39GEF0wIlWot8Y47mKuO2ZwWLV5S7qfmWo
UPe9aX+qPAnNLHFxtau5+JRQEV2brBFnskmUuKZlCOd1z7/VKFmwkMV0cezjgem/LPnZAG4Rh8TJ
vCOVPnFBET+a+YpZ+6FeOHzLrhgppbDGyRFtSULUXMrmtOjkYd9Ax20gc37p4OznZN3C374SD2X1
tS7Zk4oPt/FDV96gd9amxW6rO+xQSWvZNEF7BQxTie3Q5uQeukWMrQX7zI0+Kfyg3t0H1kNWzk27
hzYKvFmUT2BSoYD8nGFvlBYuYP+ij4H02R4vryf6tDWF0u02d3WGVWUMZ95zbrYi4AyeoFic8tPc
n9+jPO4FnNbi2a6yBOtWjsAUO4CMnrKkCLrv+rIv4YcY8Wef6j3gqoMe/5E7CIapamREoGZahwYq
aNvP72RfixywpRrX3csHQC5V4wMifwihLo5lv2SWxYZKJbO5DxHp75yXp6Lw9Ty1CvCIKAaci2O5
3Qoc6OxmF/tTyglPW/ttRct0O0F12WNwoq/IfVTzVC03dc6Zyr+jJbMnKEF7DigP27XArkBn4PA3
16LFbDq6DFVbL1ulMDg8vAX/pkJvzLxh1ZOw9I9zVMZ4vPf5U66C9d5COdq995GQqWB/Denkey7o
2HdJvrQjATF0S/ZbfG2MSKyzvRn/Olyyx9orgxt/+mEHXTCT1dGXU5WbSBPAxWiDXiobUuaw1V1h
QHVZ6pOEO+66PvWK7OP5vthcc1RyCLDojRASUpO3vUX9fpDRUOvZWlg2GgU4dZf0WrA3TUZ4lDNz
9vCAy1TRNDd+uZYhDq1keDszMP41JVtuju0j8GFJdtYAOXej6UKvKHGFiqcU6Mf9TyGb6mru76FO
3ShIvpJqiDNQqfwUhpEboH+prW+DKddQobFy9HzkJB16ybxslpW1pU2ZeYIL6bNX/WxS+3En2aZ+
h42AFv9jHI9l8XTgQ216UfTwnFEHfKJsDgL5l85w3apGFgKkrvMm4Ju1j3ZqiiTUZVc7HAH1pivi
hOoFJDMdog7ZeChwat2Z784u9+duNJ1v/tQQTOu4u5jBg+nMvP2dVLBCMi3Iws4vCWy99qkYqhpy
wm4JYlzUrGHqXCNLCz2g3sBySRhvBLfd3adSYIs0ojEG1nwfUD0/SeyL1TD5XCYRqQ6uAo8tDl4k
jrrWmbjhGeh6LlamYIJsrxhGOwsexjBydDBiWBy9qOopfIFrHO2X7Abml/W68eRJnyEYc93JR6zw
BRco+fbr4d6wdI0zH/jICkgLxqVVTixS2QeoLTTt1l6Mhy4Bm4lqMCWMJ1LXtEMT7OMGLfoPIXtd
oVhzvyyptbzQJs5h6lbCxB67REWe2obegFaEtjOEqi8J/R+yFkGYjwz/cc7yxS6wMrlDEQCotmb9
wh7y0ovUNKQxS1wIw4xSKadsPYtaz9ZRKm0r3qodByDsQ+azhh11cakwFzAmNDSaCKmKRSDDgzsG
XsUk+CGgfDTxjxSbLz7hP13OWnl2rFz9hdjln6gAvaN0ujoQxXsWl3haiWkHuBgZXmUoeqGhl4+8
ycchqf2h9KZh2zzgDsz+ps05JdGCqDUnD+e0rrBZzmMxQ3gohAdMRUl7Fw9fAQp6g+Bd6cAj+jfX
CtIIT7tsnCu6mWZdoj+zndN7CsAPDyBFz7ogimIwfuLScNIh+XNi8did1HjFKXDW3nGdSzs8ld5O
xOb+tYrblJIG0KYAElupVhTlCkTNY2Pl85x9jqwC5AlipllWDEnPemZn+WjAnTvZdGdmuDaWwi+E
bPfW5BPqKZsOFnsXP9vk8FQInZbsRnhZvkUpB/dttsZo9O8l4s7wYbkY3us1mPtMPjYOhTrFU1o/
Ok++ms49ZMeVl3mc321XFmbAJqLi7jzTrECcPt/CqKIVU3dzIVs0uGi+OtocrlboL8jku2eh/moe
9NxDHzOZ2D+uCRubnY2Me1sfojrT0AhO8Ks0MLIWo7mNRSmIEwKIyj8P63/yhkBEkB2g1IA6stHa
Vy8nIPtRE74I7HAS/BsEb/xdfHaE87xoORgMxtta3LqIUqcpIqXLfQ08bMHkYDTaA0klaLaGQkV1
h6mUA+3Ht5DzTFC2jsHMrIu4aOZ3yMgsXW0wiohTGuUVm0Ky+DFqEYaszKtEELstEeWnvfmfephJ
EW+oVKwaFpKYfUKCE4sO+1YWt/pI3ctRobl0fEroFuo0f0sUIOfILhVRloEbrdIw9tgeIFB2rRvv
AlLqJ57QjNbtXIbciV0pYI/U3Fy/0qzdURo+sCRSsE83eA5kQfHc/+6A/KhsOC2ZO2CU1H9duE/K
HgONxqykz/k00Ka/zvF0SwqNL+hvkqh2e3ldc3hpUPRl787rL5RaTTdFboZF8xI/ux+UjrHZ2A8m
70gVGX1g3xRHrGW2F7EO41RhxbaLh7bmH2UofK886bXIgtK5ZLoGLvdeFKRmOhbdYqQ1W8aJJgb7
OscGaEZ6siu8fNm2Z07ys6ea7GwwVP0A2jnJEBMGVyBS2l49zBOoHWuA5HztyNqZtjP5b6nHG0GC
9R7tEJjpUN8dq07osw1A1Td5wwG37ITsl8N9snqDy775a0fOCAIcZMiOANhhSMm17nxI0uo5oabh
rnFhmU9NsRjHXdmMw5YprhjY7Zo3PHPulSMjuevI0YKp/oJG6z5I7GUhBEv9aBLO1G44GKLHy0FI
eWAjcpudm0Dt5peKlxHZJJgtaK77ukEAubUuC8qtmFGAUXhMXmvNR+CHVzYvzHn7rGCkPUO6jbcO
8N0l2+hX4M8fFR0zFmyMa3rzYE+EEsq2Vh3parYOTtFuM3y6eE1dVO1KWefAj/OFWGNJW+/GLYmb
ju4FZykrKfjXwzHHZfY2Xu5x1OezZdBHckfDrKQqrGtzSOIxaLOOXZpNIcl0gxRmfTDEDkgKDft/
MsUELclh/lVhGYOofyq3IL5dhbX+OdaTAZgon6stVsdOGYHWwTriYMeHsSvgof6uyfku6+NC6Eg3
rbnTb1xBijusDXOerRcb13MHzpP/8NbJkej/geXVA0mcoKfvQl515H2bslv+lNhU8B/GAk3jHOn0
qCVdQISVzJlR2DFhm+v3KPULJBQUgDMzEPLJ5p8W52hHWNRVwS5mP3daL/oZowhH8Nw+rNjA4B5z
1hBrMz3NKv4N2pS+lsRTlTx6L5b0Hoz4+dBaYMa/1mSL8s3A/lac2J4FYVgNWB0dLxHwhXfox/uJ
YKPtBCayf4wFEeROt1tWbPMV7ecoB2F5I6ZPfyc5LPOto56YbsS9cwHGposGTVUb6MgjBJzUvwrb
PcwT21ozX08hr8j7aNH3eoupnGcywWVBbI3f/xpcdUKE3ibiqi0ZZ3+mORiqQQRdNJsVSz6hLSbx
IEt8cATPdvtmQNxRehFe7Tnnb9hQcD3M6+V1l/pEf+Qnryd5bmmlSjepoOAL03+Q0gfbd4UEALLg
jrJF+z6JD+JKFD29Q2xLpLizb2x74quQFCnmCx0DEDi5Ni55DQjZ/D2rj8jG0pUgZaXQDqvrSU3J
rclmL/A1sO6NtY8ozJu5E7dATHQKgzWwg/1H7ldSbsE5bHnqAkXc+T8lPG+3nrA1n5PgY7rzVP5g
hATyjdXOTIF3GmOA/rkOPLgUIKoYmVDMiOKK1mtN8h+9XavDhFwAQBt7kImM8CR7+TdreX7plk/K
p8UElDLYZhaCo2iFzSpXsNjScZNeXpRk1XhL3x0v6Ph4saIaGkF4G2zGIZ+keGe3jtnJonBQdNgM
ZEGGPO8nYps2RJh1PR6T5y0fsdI9TjMj1UJGspNUeSHgduP8DghAT1y38lKPQue77g/HZqEGam9d
iNRThDGAaTkS1vAw8TvyZv3IjSX03AdhdtdOhLiZCbr9TZ89ZJV4qg1zOD7dKr2Xse5GQmG5kALX
pftKmH24QZo9MH4lDRq3j2UHipk7rQNx63/Bo/VTk05UvitthnCw6avPMY4XGbs/Ot1cTYmGGX8d
d2/IyCk+UvDTI1ThCxKCjMSLkP0rHA98g527H70GeUjLkfoVomM4LQHAnpSOd7H7LZoC+BizJZX8
RwOI7ILqRTuPCjrjZ55EaLr1fmEIrNyve95alMjnqABh2QB6QFcWWsc9BJaat9lryul1vWll+QV+
UBkb4/JoRwsxowxXTvAD1z5ad5ky7glDlD/dSQ/A9zwwYyJO9h29HntpPnfgHVvAKnWWQzp1wqm/
dDRMLQxGYEKcMVfEWmSMH6pn9H8p3c7dml8uu/0WVBehRhTdLphfVSOLQfMpnYHk8jN80a7LS4RJ
20H7ga9nlWnCIH5W1t3o3PlIWsPBhqXemke4SQQzgYklUMe11+biPHKoqihKbBzLnWbEX1PRCxaq
tMQKG7wYF07Mg0ISMBLyrBpeXwCQp/zOqQAljG5wFyVm2hw54/2IRYeTIiad6VIhrNaJ7FIRKdML
7pWr7QlaPdeD8/mSKSKMRFoNcTwixgPlgxB2VxGXJ2OtTWtgjWYcxN6dycEPrCZBxK5m4euBNb7p
tWJd+T477rFGFCII3ToZG8dHMKp91++aYO6V5nNO659LBbqomLcDltRdIayTWqT7s1kASMFjP2jZ
cbXmAZUIzqjuow8ujqjqz4PKLGMGgBBsdVDl4dbaYMcXxh04QiGf0IC+TukHEhl/7iRd9FY4upA3
YwE5rSptQaLmQ3dUVXYpTUXwOz8iDnQylj7Jmnjfg+lD/cxsXD8tI7p4615rOIDUHHcWHRSlQbDK
qNrnGWHMnPfIli4CDiA7E7hYz67bCjxiaBYEpF9xwcGwSIo5+oEduWH1EUyFf/np1z2AVVLi2hA1
51/Ck1ukkt3NyDDMQ/FZE9PwXJ3WNbobe6Q6b9k9q9ajNYTciXHVxWdn5b4tvewmOYDSF2mEPm22
8BrCNcj7v28pF/ctGpT7YvN/5X71CE0YAN2H0mmHRDI0oSoyqrkufZfalqnf/EvN1HIi70gwvnDC
DvbdNPVUoITmyIHOhWs+DDvAUQxjrcqM7v8hFk3ngBAPjTvivLoHdcN7ZAkbRlAZ6GkjnzrJ+G7+
kcYuRFTj8iZkutjvkk6PH2zHLgKzlOs+1wZkcFdbMDVCZIlBqoBDe+XQMEvEkpInzR+LXIeI29hR
vdRWMGnqtimoOJs4h+sGbn7Lkf6D7dCr+drQqeYhype5ws0x+Sykree3mqPX8GYo4r5zmM4CVd9j
5QJ2FPfkZqsh7F1ncIw2bNZJ6E7TMvRm+c2Fk43MuysotFhPoU77xSS8XaQnjKUPaHRzslGzTU/k
z4FYXlo7aj/lCO4DpndVdvf6Ck9HNbY547rrn4CFXiEsi+K0dQajoyc5dH/F4tU9gDi+gwmziesX
Ga35Os2Be+qBLkTQnISQ2Q1RURdhgK2BrAAZOsinIDTpZZViAnNIxtkgeC0IzIU5XrLoRaoVRtcM
Fa9mFdSgQG9LCN3JJm7YxxndWFWMjWLge4AI5x5HP5TfPmGnn14cxJDgwInJIoqXeMSe9rMNBFTO
bZAVYEkfULQ4IRYxJzoK85uklF4FloIbHkngoqLbWpdyVzzsfyqSKfy8pV9y8kxdmXXka8ndDJFt
/13VkE+w4cCMuFO8gaGTg34rRHAlvgDxHQxgot4bueGgdZZrzGR1EvdFq3JT8BUkdaYq4owV+NdV
PBawf+uqz/GQQwXWh4lXdk68mhpadswh4iCuVZID1Fv2ITXUIMn92+HAZOmUlCNvkRC+r7IvvOcY
ge8SY/XkYi9iXaYJuIspopSMbTST+GHE1tQGdbN3KMbQ6NNWeZ1MU/+Jgn0B4fmYPrClp3WI3Tcf
sOYv8qU4NZDyqDU1Nqh6Z5jyZYbpo3oW5ie0ZJ/68d3Uq5BIO5oLc5PWVwsySnhVN76JK1rVIdY/
IKW46/PKTXXoMQAx81elNk6RMUitKhHG3nW5lQ+ZFLdHLgN8TopcHGYURx/tICV5/mC8oES6x+yr
2wOXvMgiLMXbhJ4uBosvgECyEpjf+iyzNRYfrCrwdjQrtmIhD9geo19gQb6wDSJ/UtUePTOi9DuO
COTvNF4AXyU0VeXgPMnpognpFEmyfNWZelIWaKQGwgVDfWGlVpUlAu9tmthVZh50WxOgLaubKphW
pTFpeCwJ5phRNVe+L3tKoTLdmCVaX4NkKOT90Wuc1dwWuBfpTXLYVtrI0gOBLI/18PIS5rA/exWv
ciVAcVNb9SSHpNAEir13MkMqGekniM425Ll3dlYTC18pWSAh558SmF9Ul2ULGnj+xJhkz5WX2tBT
qO8xStuBCW9Tfls/m/cSc4Jw1PYS1NBzpciNqREb8cE8IIZ5WxosQhNHsCelmH92mrNExazcpbDC
2eNyWjW0BJnsSmVYySLSVJ4iATIn82a6YYHksMSZB41j6yho0MfTHxo0yFT3etVGc33vcVggN3TV
xfcy+AnLpfZe6SOC4nt8OQYdr/fZAs06jzgNXflsQc2kaWBmj5x/ZTQMd4PKTiI9SXB7Gsi8jbmG
NXfEiwx/0+fyZkIX+myhQMgIrt73SFj+mob7jM43y7MWlThpl0lzvnsJ9ILXSgWPJ+Jw4f3BqezH
4hYzB++B5Yq4ScPkV6yvdipxM7r3INYYwQMj/KSuKIXVx3adVlxn/05Yxip29vWqK7dC9MZYXM2F
Wku1NAc1uFu2l+DV+AFAf46nYGpfK0Xu8Q+U1SfvSptOtvhI8NnkuOKoa2U/iOxIAfXyCR1ix+VA
ksvWD/89yhK3ZlZqZUM44mn54TqpBCUvwli/1fYLqyYGod3yBEarcwBtwXLfbSy5xYtA4sYIMRp4
TM2WMgewRUBEpI4FuNA3DFmisBZAH+p+9LekAmTJ27mL1gR9HtGGIk9PIlQgbTfwA3JGm0olk+zt
CZodZViwY4/7/jA0jek5PZ9IJIkf8BVUVRS87lLID1cuTObl9L/EKtJaZG/ZKPkCym+KW6tXsV8P
N6vMxfMWGfel7s+z+a0qe+NTr0U4T+gF1+PnKsB9HOFdsEFOmTE8oRmHK9uW2lSOtIXwNmMNlwL9
k8uFAgb2gQDarFC0sek01oKDVwuoQur7i1qlzREPz2pjVGE1PDdDkjFHPeeq4T2kzKMVeeumt/Qu
TaBzUpQuznA8/3/E7DkKW5exNKeLttAdps0S4y/f833iDK7E2UJHBsIfGctnh6jg5615KoOUyJrT
irDzDYeloaBf5wm+CvOtWAhWzHMogBUX+hir0+XGHNeYPOE8ItIPn9Acg9oK9uIb6xjXx5FMXCd9
xVxQFrSfUk1n09mrnIbUCHhdmOkiu4kINZ7ygsJX/VFTvEPDTJp5q6FSJ8h5n5wzG1DU+hRb4gs9
e5JAAEi7N32jy5X8uMknwmskTnkMXytztkBD6e/aYHWcjxmEsEKcJzKxP5IzmHdoorRMmvtNqWeH
KeUj1hMHvH5zX7YMSBOnQFsJ4eaePQREvupKNbuipBw20LtQLIa7pYx9XNvPdJQTuHgQkMdOnzdZ
TJ4ZcF1x5JmAYMA4+RLrN3XofcVVtlAaKFiDNV/t7s+n+9toG8cyzpUv/ofiw6azOUbe0KwcfpTh
qwaPZ6Jk3C67LSh8DNhefYg/CH782siyFq1pUiSNG42QXqHaD8PKSNIS4gEudIFRRDdcSxURn8al
FLa/kcL7bK09ELFPdot/WW+UnLdpISVWfH+unskG/jY3prNxVh2ljMdXL3ONQBkSh1BUlj7+M3Kl
VLUwhrTBgs1Lmyja61+t9mztE/KIR/jinEtnn59XjcSb/H+LCriXrsFc4VN/ggzcAALf+cSWBdtx
R2ZaNfUPFnAUibq0FJfk12vSyNSjj8ryviOI4hCUDh8ft+H41piHkCVv1vUAvR7TduLjchBLk73r
EJSZ1NEypbZSK/3KzDGVLUXGx9pBzcJnGIOsGTy4LaOfSC6K7hBR87iZAwNxzZutZGC/ooqzelhe
gomIu3nRLVPbViNcniAdGX0S5cSs2Md3C2SNLivYZ8LQn2n8MJ2SiNP7IfWMmYIdqpiSZNWkH086
BvfVN2cj3lGDRnHR5fH6MqXA+PPBb7rat7dtWJZGZkeFq2x6uaPRWzUbluGipYrpt3VnHNeijfLw
srvBQ5UcIeYmWL2kSKFTI8YkN5XDHcN/sd0O8SzmbEe0bD/fBuvXEtONfueO8DomYJLM/4vwvIhx
gRNPtS4BdnrRyqm68VJ8kFUCnSrSavV+7SbUWonxq1HN+9QH4RYe/771QSo2dSiOTm3o07wi6jdk
IBl5R6sRk3z70VCEFglHMuJrCYZsbou35H/bmgXVMZqYGSpazcFBZNJeYRAn0nrRcEmNIhGTCgdK
5nz5Q3RdNYGf7RMCyeHSpeblh1ertjO5ASeQkQQyqiUkHeB4e7F8ASsVBkae9bHvXqo0IHOE8O/x
U5ph+dMJpGL8PZKPGhge14sg6KLWgWuJa6maAEwiZKrgjNVr6xJCRZPH8146P6HSpSybQM6fhbeI
GuzhYaFXZrYG7yXgS1ZAkPm8HRLx6RE0LdfxGdY4t1sslGoYJm3J8EmEieYYnLRx3N/5ugMUNdFJ
v1//1JmO9fFwSCqMk222XKStBWe9Sbo2/TpuaW4yzq9xbr1pH9kilxDo6ZJL/IpDldojGWGN7CSf
dcMO8LlxEfdWU0jTnZBkGl+uURH3ZnQ5bx70MJ44/yaSd7AmKvPv57U+C5uX3QyfEsws5jY9r405
Cp2vBaIO5tJ+J3wrmmZTw5DxyrvvnkxdxHVWRpFgsbH+9dy6aLTTfM0pi6C2iQgpNb8apYRPI1cS
j+Og2+OchV70lF4MNSFf3lbalUoT2rOsVKTPE98qn6AuXeioxxmedYPSvTe71y+go5FqcsJQFRXN
ubuSMrJqQVpeYt4IWVDud0Qs0gAPSVpug7ry1JC4Nq7j0l1kAovt59Zypj/DsZa14fL0AI1S5Cl4
xWymkLHV66uG/MRWatu0EAAFKCdGFacCGQGmt/LB1pYTZd18QE7rhdjzuL2k8Ztq+Jhjm9fqm7Xv
hdOP/cYAIrruhFax069A7Vyt6G8ggOw+HT/wFzO8UMcud+evtOmMI0RhzOPdz4QcFzvQUg1zm/cX
SaDgNrin0vPm3MmMQ4GWWtygVTEuh1SBsj4ulpHjlMMzWBeUN33xd3No7/4qCfgTiRZOLbWrgVDQ
lj7gcRkdk7xWi9twP/en01UyfPO/WrI0Nz0Twt6oiEZGXROzF6FI6Uh1VW+ZGsPGEpdWII0INnsx
D47VEjVOM4gWK7CEoJCKt/gPYKy9r8IbOJbplmUs39Cb2OUaPmqKU7dZ5s2FF+raO+8KvJe1Oxmm
jP+mypa63/J4ompjByP+cS0AvP51muA577zNyq4eEznM44Qvo39m53fB1tSaFaIRCEXxhNaSDIje
JnTlMCqEbATGL9X+5LckmPntB30Sz9xX3nH7XJ01tE+QKTzS3EaH3PKWq8UbJmNtPCz5LlsLI6fp
pUUjAwuuOOa0fYHFQ070RGFyHYzYdT3y+MNNM1ikxdR6fYEx1tw9ZK6PocmeOVCw4Zr7ytRTVMYt
D4OCLQIehwchGoX/YHWGHk7eSl/WtUdoj7mxmkc2nvgWgbkfRDLURgZfBGDm2OPPfA1e41ye+VSS
9Xc5FYgBqT0hNwr7DX3uFCYb8+OCw/JOMjssprIYy2zIKGr213hCt5wOHaSTxN6u8PJPwYjRmpJD
1VWFhUOhe7/n15ytvP50wFmxQ8oBb9cnaD17fcoug94VSdZtzbhrPeBVsDS/f3SanVnvl5i9An4r
liCN96glh6WAX+gTUNY1cU1Pa7gJLN934o/MP+presg4YE2eR8UIJByayFFWKqSaPi5+Wf47qUK6
MlMJG0xw2sW70SjSpA3C75tV3UPmAeXAWchhoedaoo3yzFXOJi2rTb0MqXzqrZ0NcOL+Ohs5jAGj
jq+ZtkxDO6qf9HGphtoygPjENjoEHmO3L+Rf4MnYkjW2G561chjyuJjmB4jaKPm3zKNVvLbWgRQG
l+3+T5o9j9NnU/myLDmpE32tO+jNw9yFb7E0h/D1/7RnML7Y1je8Kz4ZM8ZM2KOSft8F/bjW93am
Z8DFUQljjGnsQ59DQbQiIp41ncsGPJou6u1o08C9PRS0xlRmRYttrWgqUPuQ83skZePLlNmkAdUj
fktXv6Ngi6Z69fh55WHDo26T5ntn7g7Nn7vERALyOfVsbdpkK3FwUAfPt7KFokQf1bmfF8OYFPEF
e7zCWeXaClZytQDlg66KWkVf20Y63eql3pvUM2ZvL8DwHmgcDs5us1ITeMQx5a0NOxb0frjyNFcM
hdxMoQTPtaMKBR+6cJJvpR+oopHpb9k6mlBML3VMakolRza6f7bNXSZd1RvHe6yxBZqpuOUz3/5F
6yvjxFAjhl70x201wg7bf57DLVYybOjne0IC7CYnFPPNZrdY3qcdpvh+PsJ9+9MLO7Q1EwXAfDwR
qw5madvYTNo9t4emhm6adCHGzZ2uDL1THoI0IAcIma13LXa6pEpiItRZorFpPW0QztmV9F9Zq9ue
tStuEMdXZnA9YYyCLrptlF8tDvZSLuuLQsp1OjgDGFbW9tE1MifjHC8y094jyAmDuATUyWFnQhFH
AKm+AJRC3YvhhVJ+ct80GqapcrqT6g2lar0/zzubVdf6GTJsSoBcP6T5jswfg0KnlUPMk2dO1WnH
OgSt9YYfRIqMrH5MMLwSdp1ZqCGSC3YyN/zS4Edsl5rfQjzugv8ATGWomi/z0CAuLXTwupq6zxpi
ETuzIXijTu3g7GxplsHqryRmbjm5sBy75+EbaEIPBtYtMqH1ZyB4Gnmofj9q8e4xIo/o9FgQVR6a
YS7+FaCL6mD/uTwcJmhGkRbfy0Ho7FcW9Oz+9TDrq3hNBdbBskUXCVEYahGj6AZvZxx3wBQpLW79
Ca1q4xjOEm6T3Qpt4kHRZS5tDvTUL9lWk4RRDmH9nSJsCBxkhNmiGLa5Q2h/9+oxBR4Tpkbq3slL
e1Iq1VkK/wVML88dUjAFWLCZ85SpQfFgWBR7QQcQjhkfgmjGq0BUEqgDgfbj8+xi6L8QKCWokXN6
bMgc+RkXgzA61dRGS81CJQcq1Bm4VWZIGR0e/HMbmbBfWfe2XRy5tbc45YeMjwEsxyamac/dgpT7
Fc2yoyXjp1lyxxVkodUf6/POWqXFO1OlaTNjImihKZN6jZ/naXZRuNv4GgVOGniWynrML8bV1klG
f2tvGuxjiov2dswLqbbwXCHfPf+7xsbg/faMbvMgsatpWR2ojkA70OVA/tbHxn34dUoFuH6XZiqJ
9EQFryTIaOntjX594Dthj/9hxizeZbu2V3rn5ILXapEJUnArrhL6aYK6P9Xxwo0B8JwS7oeNJHt3
ZxujAhH9qScOsImpQ95xnUSK/NfuRUme5EbQR6JpPBS4qksRAovVvNijhjjCbaa7jsbTvjiFFdUj
km0eW3KNa9ahsdpH9il1BMPvfT7VxLL1rYEs9/eZ9sOFPJV3AErIBKBM2z3EJx9rR3JJdKAi3yMU
xU4I9UJhsMp3oiWxKhSGQ/FVIhZxf9bRMN+1Xf/WK0lBJVhyDDYeQNgRVozd5lHoTeY0mjXGOK/x
9j+i9gllZbNhPHDr7qkVHutOsWXZNiFlZb4LMM6Mgb0MvnJTRZGNhymVFJAi+Px3xfs+Hspo2c9i
n8Dmrmm898PVlVEFSh70onzwoTRQBXGLKiNYIUNAkew5ffge+3Y4E6JoX1uqUjSlBEoleYdV+Kli
f8r4bPsCSVDy3eYujMUctdiqvPnaTWLayRSl2HOP1tRuVtEi/eCXOhTlu8EBCHX+AOOlORaqcxH8
/u/0+WwsU7czcdZ/NgnSv74pUJw8W9mzABGY0LURyh3BXZ2myn029/il3c68L5zhL/F3orlbYUcM
y/GxW5S3gJV+7c84CBL/iGvQzkRBzQsYYD8L1MHrZKq4Sqtrjbn+c2pp0ZPdQQnkSGUG52+7Fvv9
Rwz8RWDfvttXMHiiFkA5MXMrfdtpN6EwNsydAVQfQViCcx1HAfIJJJKMALPpY71P0aZLFHM5yJqh
nOrn/5ZVYYRkbdYoDfDj67OGIAnSf1aQmjoFroMTb8T+A90r+2HY/xftaxR7erfdDpePEOpqQvik
JKOHyffHPYGOWyMxrv8Gh76xCV14MO0MK65Ho6TIfMaoHewlqcRkpnBGTihSaBDo3CN/jv4I3oqX
ZaZnKj4sLCzS0F4xswc8hGUb3JQ7BmlN/1dFXAR55sdfGeX+C4Xl1wdCPPgh4NmIZBsfTMWstuaO
uMg4BL2F8r/+rVY6LRhTq4/7rK1MqKAiZpeRvL/f5qTojdH+mXDmw8UWW19K+jtpeEdv3VyMgsVF
cYWqOOjN2ge0Ix9clh6JZm38Qb0tY7r+8uFL5Xf4f4v2YA5jYZ/JmQoHu96x8gP5jX+gpatepzeN
jG/L62AlwlmUuCr/qqB7lHoEIphQcGTON0z2+WMksSTqAbTvRHt2T1Z9D1onFx7B3cG7cT0M2uGD
3uKuDwywGqjhPpGWTq2dBJB6n06VgGBcmMl3j1Tvv4V2c/ZirjSMVHSIeEsOr27/kdffYIY9Z7Yn
+zyvc/+Pp+MeHvv58UvovpFZRhBwEyxRmy2FjCfcuR+lvDIIDqPzyjjshm2K0szSe4sUs9YEJF2j
C3yCmLUWDPeahmgyhkSyB4OE+KPCVBNXzBIrAfDTZwxWtWHHfUzvQKN14GD7bHywoc7kGK8F+vUK
46/ZLUxqTpJBPo/74zAmw+AtbtneEPNBfTTyeKZKJ4QbyQKEQgkURSeVUzHdU+00xTj4TTeSx5XC
YBdgiQkbz0usBMlxbdLpi2ER5s7iUKFTfQ1ZjvoYL6EeWMQBxTBXJLUaiko2hMoLDHuOTmIQ7j1R
qQoKDkhkYD/XcaS2kZEFpjlEzLEdUOpOaivKMj6JfS2kmAuMSgzcvJmQqEYiqJHGDM05fXmKfWjw
CcSI3U9vncVc+puAHGhXowoRtf1PJvCUpYVq07k5FQ4otHbgmxs/nKFRj1ZSIOkz8Z4XtW4gWww5
55AxVrERRQl0vgP6oCyN59hvBoLHn5lRjs0/co8e3HFr0bxpu26CmNBvQA+rpwJzM7shzwbzXsp1
nFJKNOCGfmxYXnj3ZI9wl8cXJkcOxmxYGVkL/VJAyAdlk4LIK79saU5RutAONePfXY31RvzGqtNX
JddLBnUQGJWF5tfh6DBZhEftFnAyAEdxtisWLoDVqREcZD97aDdiVwMAjj4DEwkbiNnViKDfXBdE
u0c1DgjFsh4rWj/k2csIvmVJu8K8WN/cQk9xiCdogzKUZc74xlqCPBrXgOfRNs2IA/UkjfoZxWUp
9Oe5SsYt9S5Gg+1YM+Oxax87tZycg63ZleRpza6JlVDD7YUUChG5OS38jwKGMengu+0jcZge9OUt
yn6fxbAHIu5t9D7uVFjwW2OpMhLovojBoaVbI9VjjVuCgE7ArwYcGLT90l0VLEPAkYwXjYrwVCpK
+gUAEDkcDuvRDb9JELZ39Ol9OWFDe2haTciwj8MT0nguAeDp9WZ8S6nSpfa4MAxJXTG1WQC8BI1E
9iW+HhDuJoR5p9Pxl9LR6l5v49lCrY3hE91GjXDHeJIcBWLBvnOlNlvuWGxfuAQp5fUjZzBo52ag
wa6cA3uhQBjeW4d38j2vDsIW8xGZI9oW1pXqOShPGZaslUj2AUJQpONUUM17IGxVkR/eYuZZ7CYS
vvSAmw4H8paELVl7kE+zqetDNwuAVTYg7PSiS23pi/XZwKPnz2zc84NvVW4/hY3R3i2sGnq6dmqr
ix6EzyI/MPsQlAi2Dn4LRAzSwJE6rHndkHYaRpero5yp76bWkaz0eZIh4eAOVWusCBWlMPKHuUz8
zSC7+TP6YNl+s9oe0NogQ2zm3hHeJXTrTxDDmB53sFuYzUECq+w8sNBDLblYIHPCjnp4KyRO+UZl
FhbeTEx3Yst/ee4H1KMyeRnU3ztPO8bBL6PnRX7/LdCM+IdwvZ4YsvA2F/8v9AL/v0Bh0nd9oy2F
d96dM341/qCq7uI4z7M5qeeZ8a1A9B5l7I+hApmv2IQOynK/U42z91j1P7Sk1tNFGgUy/bMFEoTC
DLpIMin9l2kyho/SmsLegKD4KECfbaQyF9S5qX8xpMR0j77TYMMETgKiWgtz0uoK2/qRFcIdv7SX
q7O3zt5W5yhiTKM6DG+fQ69A+0VhezVvr5ZzYtYVqggDlxt69IniSiZip+WXKcwsBINCOxDIWrQD
j6kCXG57fn33s68evsUcLf8BZ0Jd0qrJHyBRvbjQeT7I3ll5GBbsXAD5+SESqKu5GGI/BUQhspPh
PWrPe3dpKWkhfMkOdmA3Q+NKk9+C6kn1uaYf+gshqoAhZB6ZsEJWZc90XbDf0Y0bIjF2HSYtsP7p
jjz0UkIDK8pTafTnF9EIpxdRBMPwHwObTl2PRXu2SJCgYoRT0v4KWZkref8jvHrhNVkLj4xoSWKd
uxSpsRCFzBkugWFhrC3yavX8YmxQzaretAOopu0i91oqNdAblagLrl9FYqGDgli0CDS5WKUPcFl7
03iXQlIc0kpnTFZZAWtCS494gDVJq/1Kwj8/1bIC2CHxa3/hykItepBShiWkCL2iDPn0HK/yRR2h
YU0Tzci03YJTyivWuRHYIRgNW4g8PuVGzCFjkZ1KLXlHRbgrDQFDetwvAxxR4t0oZLITn/MmrxLQ
sU7BSCiSUlzdsGHXzxpX8Kq57YJrdBUJLWJVMMKKdvMRKTM8B4bzBwPAlblZPKV+RfF1hEfJDAVi
VSkH2a9APLtDV9mZ2DK7dubq5YwQSvy6J+5NRaj0CS9OM3iz68I9ZU+mYk14TryK3xwclJaiAKic
YvfdwsKy4EDdayAp67MSiOGBfMiPzzIca9hbYuW/N5Is7zR0Gtaw7Sg6o6ljxrKXIlA3COVtPgHa
NY4hmEke6U1tjaVU06Mwyg9Ryay4N99bGRhFQmajZVBzuLw2AREauL27iTQw5th5DdvaDK9f64vS
8DXsI5Qo8PmOI2hffX5PMsbvII5QuphciEPrC6pIZ3Bhwgewzk0UT6pvZTYN9ok5bIBNt/aOg5rC
sR3HojMuBlpK8J9HkubQhoEzSFiAJlxuZE71HdhGULlb514JKhGpxi0PsfgavA1OkhxbLEnJJLMv
Zb8rwdzMN5CS4EyO1UEra+KY+KZNn4qT2BWfnpeuhZmk+Zkz14CMtAiIm82E/hx/6oJd0+Aq67jb
gb2ZAnLAYnKC8hEFh5Go4Jhc6duBWjHuxbXGkSScTQYEQwiuBodIlTRL0PgY7a7ZTMSxthWJcJz9
RHn7+g7w3Bp703sTQmOyMm5N/BWh/QWvhrJAdMVxbTPZMf6rXosMvSHZXpYgCI9q3/wq4yfviVkQ
HlV2+/IyWavHdZqSC4n3tVSjtdnHhgtn6KWZj2q4HRTe5fKOGbNJuTd62oKWdpEs7zrp6Q4Z8BJO
UjTCPvOk+pXO+D6PBOGhi+bsIIypPadLT9U/rEhlkKigl1dFNWVucB/sbuOsn/sZvvgpnMMlKDCu
QJR2mEeobuK/S2a+NN2l+p4qMNA2iPxwneRHK4cckSb41DtLrFcN9eukm63KWrVnTB6M14hXod7c
b9wBVA/VXL7lQXEUwdEygJFw1nmFn730iAjXlCcULfI7Pw0ptt2bJESKebdVRsMgqUvny85arhAQ
8F/gXwqTNogm/V0IrSpXnYEgBhwG5F89rePVP6uEiU3XCAt1BT3NEwrTgcI9IiYtf4KAdkows5zw
VDa3rspqaVcd5Rvmgg8jO6wYznQm3KiWH1M7AlhCcd58WC9MGwjOUR4QwGL+dNC/xroS9J1MNtRV
CeLLFDQM757Kf9fPPZJEPJB0R1iFeKc0ZJtDDHolqdMxkHMrLyRPT1hKxgOfVC/eW4bs3za9KntA
0pxa9B0uHRrZKLTIb0E9yTWn70KSyne2//DNy5rDb77HNtlfVmdIjijzTJppmRRUprI+dgwlQElF
6mj0QNSLNdM/3VREn00+cSUkLptmuV/qUafe6WpyI9pYvVFpJU31jTe5pwsGyYeBt2zPmAEgGMEH
qQpHl2mSJVSS+jKr4VvfSbA68HG5B1CLqtteAmjbK7icama2aa7ldeXm8lrYeitmfXZVy0MGFvjv
upW8AChgGb14pTDZfzUjAfTHgoP96Mnjsy3RyhhC/z7pX8AyigOo2LY2fYHnwLY+SJodEikzvwFX
fJWO7FwM7Y6EUH/dOnGA6b+J2we+Ew0UGoGzCFm8yi2z4v0dHrXt/0L2vF7XeLBkrhC9TzcAldxV
zthSoTIfzqWRrsA8S/dNP/YaYNSd9WlJ3qW/Dvc76JmK7a8KXCsC/WB8xAsBO+MhQISx8gdA3JtY
CG40ZvkfCSAesGsONwoaJJWpdUPODLBdxA4ARSwpPwG9ksva6ojCrD0Ds2oTl67mbqaamUZC6VGP
WsaBOYmPnZwffE4kyeI79o+CzKwDxzy/y9ZJ1ROAab0Zb96nEG2Sp/2KrMocM9t4SfTNocMsIOcC
fROpDIB3/BkBCDdcGqhxP0+bpyIJvmhyrbrxb+YO18YjvOye/Poe90g57bXCqtrpTEURM61Oako+
hmpN7Q28LvZmk/BRmADylnDSZ4TwaqSUDxqZIlIYtZfOm4NXVZDx+wsb9Ex1ddxnvmJQbhoBm3to
IVuOfhXlth+dGQxEMBBRRCop1NYrrF/nKyhRCG51YyXHHhezk2HQ6lbXveMQvA/OQWhLtEHqYj6x
eoJRUN0s4zQd7ZffN8hZpJhD6JQDJhDU3YZE3saKkCKRjLVavp9Mi8FGMp3pcSZPAc8NyZmrpupG
pscunnOGCgk8u6j+C4FXvaoKDTt+oeFGdYMKUyXo1jYfvLjvhvbtNh5L3muc0SYYhd62ks0CiIob
muuQ+l6SdSdSi4GA6wdUyqOQK7VSoE6rpuLHHo0RhUP4HTViiBfO7WcupaXkzCb9cSNBTaVBJjTD
F2vU4FMzU3oqE/Bm/fX5qQovNOULHq3g2tk96r1IYb83LIhCBgDkLaZNq+dMWZq9VavyCCkl1vF9
qTNzYw6MXzNYkOlRbNh1aQaIiQYlPUiJ+WCHLXLDfDjq3vl6+yZT7V9tHyGOpHS0wwAv7qNMN3Ir
xN8hWPXZRpT32V2ACbMcanRufSHdjnVxCoMfuhLdfKGnoEDjl0ninOqC5jxbo77qMkDWPUvcgSyr
a/Y9nPj+IMObJv8yCuFPkRPPIzkc5TiDbAM2jOek91oS9e3EtlDpzJ7n3cfQoV35ZfY3K8KS9Q6A
ut6OvrNG2ALGwyvev06iAZR0/eUTMvL6Jtm4BYn7fg5UYuVqy0DCgxaqgMYsR2blYPjkZBzrSFR2
aRvL+lSJAme6pLQbOK3uxwYibxj4TPdkINT+6zI8vBtD82xRifYfMuva2Xvo2jTTVBeggkSZsvVF
pqukvhH+n11UJGH2CBEVq99ROoOiEwxva5IwzlK7Md0y4DIPDfWCH42cGPTSA9xfwh51NGD+yH/F
cJcyWVkr9qkKkUZj0Y147cn1H4GufqSmXSrLZbebRP0WUuJIl0skIw2/s1vsSIkQtHj2Fu7HQOx8
0JuYc3SQ+UTQKTWq+wd/DnfcNhATxD5FpR/2LVg3usoah3q8x7jKqXhMYEz7NMqBgfrsT8jxFESc
yWrSz5uiCPCI7tIXKJJb9fjI9DUCIMhPERMGcLM5WqYUfcs2gpqPqrSpHVrfOzQQz8UpjwyEX5Ss
zaHqlHHzu8J4mZdNHcG9xxSxiClzo+yStb5VJEDheT8Mc6PHENYSw8aEt1MQnDkZ5pe1KaHSUNgu
PcPL2qu4FY2CbWxiYMb2LM7rZ+msdfS0IyG8AT2mbCBXocV5enrY3EDyETxE9UbWTOtSAmu44cpp
bMEZRyiw/trroL65FUVP6TApGP1cKhVhetSBHJnTZcYiSgCnwHCUnH8m5HABS4cnaEBFZO0ulJ46
Z10cqZKP6KvpZpTrQ6oaAM3EEsv+h2P0CObji8hy6Suc31X54FPuuleyuVa2RtN3MeWKqgmufPCp
utMJ3w4yhQGczDCVHkkWeBtMcbc5pZRJXHm9SEqMNt4OsCo1GpoUUwUwz0fGuSaCXUg/SYcgBfSI
FuFfJhldYSte4PiLFMAfukydpmGyTSQaSeL9GwUwMdxjvd52WFefJ26FM1rYGEkHrUsNmikLstvo
i3oozsjcajUpMvYjZbPaMaKRjVWAUNGYxGI8WbCiR+SXzfgbJzxxDraSoGF/liLwfjSZvj0O1cBp
auNbi430mHde5tzF/2f4fDhzN3yKCPsIMWRS0IMO9EKcpFYzI36N4r/TaLcZXmyL0bIWwhfPnujU
ALtNBAFwqytoavRf+qzdP9wVjIhX/BG0z9DBJMWCM51I+fDTWcukyQDobBdYEdYkDXsLSvrjbS6I
X3pTWSef0z/T6OCXpBJ+JB8zLBsjUNfCf1L+LS7jRvpxNf1gbFDeT4aQSx+NyGH7MC0bLKqbGHwh
EzJT24oYVqFAxGfF90jxhY9O4phFM5cxKbIzcO0d9tNz31v0b+nWZEpEHGqVK73EtQWhP3AsA0gG
EOSsuwr0+JMHBobDSdF/1VZb4PHij6I9lMZqC+H8W7U54ZPA5dfd+a2wnuP+t+ooeAD9lm7hH18f
UE+2csswKjWuGkiTrwdTKY1vXERF2coelYRgCjtCAiOutwAkEE9JLBbvl1fKo2hAoBqPowS7NNwn
t41Eg+KKyvIHysTp6MMFadnwLgqt1l+4s1Uk2y3jQYPV4uQH+KQYXbkUJmkfju6Nqk3rINsRO0ph
biesklJvl1ToMKFut+0kBSknrIFk+Uk397zBitfF5NHfiBzHqSEGPbKTXD7tFz+3q3BZDmlA3cK6
Joa2KJQBCdBZh9I5FY4qd2HQvvcK9ZPU2aqNRbcdV49Fxy4mJnjedSlPod1cK+JH1z5Ke11coJil
mPa6JphWUG+ow9NxG46Q6oMTZUgs6jokisN8cn8kE3qjdqWs+2xB+I7kkdoPm7kFL+C/fHN5rYSU
y+qZUPE4UaRDToHCna4FP8Ja1cDgrHlp0d0N/15Ys+yCRGn/sGQchukbMElzw2B0eRKYJd56205e
noo4PQsGWf/3rGHfQX/YM4LFSGLiCgKZ2XiqaTVNIMoghcGKKMfRm2ydQibvzibKHYIPH4GV3F2y
SWld+/lNRDcX+xFh4dymBxf3+sreHaS4oNgdKDaIF3cWW3lnDfxjKBVd5wMn5FJyUjKv0iBQ0Pib
niRZMoT/eo95AVHe38rFmuPqfcd3Be7ljenuPH84GqVL5PXxxZyMb2NFy6H6QjsCcsPK9lMTlPAZ
X4YnTIGy3nD4NS7u7yuJuaQWInuHYNfMW3b5d4M+Ag4SU+2E2E/I4wryoPoMYkqEUXr3Qa/cWg6N
QJ4X+3s+XQ1fD4C8uv+EVfddo0YQSpua1ZkPVKiSXHLErJgJwq/ri6L52BApAT1GM1udClEwZeZe
ouG2BLsms9BbfQ9tz2vAeVO5SCtu/uK8l74AlaMItxtmzkwS5lD/zzvHpeC9PI2GyLw9Sp+ABlQS
HTkdLqmHRHTy/PHHkua0hZKpQrgioKM6z3CvVh9N0JxSMm8T3xIzttkZy3fGGU5qi82o0lyMPl1N
MMGCJTN20/ZPiQoc1Lw4F1DVIYkoWH3zUUv6TxKI1x6gZiXmjBfWcSB6Wo1CwPVD1E0qpINJ2qpH
0xhnvkYNXBcsPSYlGNxb7a27ZMizmBLMqsCuU/Hkwme2NEHfD/tdU071BY5TbmnYfprtbYRWSAzN
GisGwFuDao5CdTm8skrmlGoM36AL4dStra23BKLN9wqkvLfC2Kxc3aKqR1VC7/SzcKR66dWAUc4K
MOUBpLh5U14uNZFG9Cck+ouU3tFrHMQBsSZdnoCxFo9AaWlR3uSy/ckDzsv/VX13kPXoADkVGArs
wKDYoVEwrxtFVvngm2OE5Ktu2X5Zsp9biNjTuImXjOi0TvRhU7pOz2hRYpZNaiuA6ZqvV8IuCEJY
Fp135VSldv8kqjsAv27W/6eYKgPUHpdro/FcoI1FZpXp+pNZYX9TWMu497JoHPlHltAcdij+lvKH
VTtLGAgYmBl64+7iLOB5OW/ZAKY9A66dPHl7nlD/fCItvfoYW56fSu6F4f7uERfqpqvgRMrlja3O
PA0Sx3EpnUBg6wUGXQORBmV0OfSo5yJKvZKpUMIVezG7b83KWcdPcj59ji3mmWFPxWubyhZafBo/
u08thFnZfuFb3UOT4QTUi8wfl0kOCsTvmr5+eoLSoOoMTkYa9OfaYpYREClBDcTWMCTKlYjIH3B8
CPhOz1iIFdsOJs1tCmWenDM8rAeyMVFlFsWyKFAn8/QgZwOpf49lqNEjgwtgd7RvrI07ngQMNVN3
kW41Ip2fiPMfgLBf2sqPZsaIASDHH2aKkc6T7ejEhfEwGghCJYsSarU2fruxgFrF+nQTLDmY6caX
qYYeQDwsEDS77vYdUu96O2tN8zyPrDAKU9AQCCQW5wQypm5n5YoHNBUtLYON0qKBKg+n7j4vrTs4
+pDaFocFwT5CMpCJ9tKfxPqPYhwOavMRC/zyArIQ2yFtz0Q/Rd3NeOctqJ6nXj2DXZDxdTTsmPIy
4uk5KpfDI7tadNceV+kWJqaM0Z4p1ELOCWcf2f9toi3PYUglvSdiXh1q8k8vLTde24KHzxe5JKyG
cfnowA8oYJ4AwVkdtLhq2SNEUgP23+apkKZAdyl5f47EcHttpKKnlvyUDZdANCAonjyUf/Tbq7YW
3DTjIlN6Oxq+BF+At662ZC8uTn7jEZ7tckYxNjEuHdU3QJMOjSTG68wyayXYyfoYWIVIScvSBtTH
OHMHC8UISe/izJKZy0O3D1t2k36qirrOnUxMWWduWUDJPA7XnXS78B/m/+lQ16yNR/1+RQJeeKR0
7yRBN9MumtlfTltdh0rmrTx3tXledHdQ182PdJGy+5Nblky5DI3hL174MuATOBBIWK3Icdt4b198
VlyWpM66PXzQzsgiAXxq15q/kQynPI0REZ624Bo8ZQPNvi/vRN+75GWi6NO7pwVW3GVYQJBjYgyA
FM8bs/hgSTk0K12DkKRkdY1kR2fHtpUlApZD8oRFhtIUB8+0Yo0MarPBkKvyROp5nctbiLz108Z8
hzO0nc34MgQMOVC6GPjtwB7xZC1OM394G7rq6Dgy4jdu38FvrFs+IwTSHMR7RO54QrVg1YxaKD23
SWdRvaKhKluawpVFqyeMOAT72oo1OpjAqB4zP9Qp1cvrZTHurYBWxJ9mIpxRkwamphQv/JbeNeUa
cAdegEYSrevKZmj/r15iRf1hp7Zm24v7ahwXVVXNaz90y2vtAELbhsARvgzmd4KooVmgQzZ4XYNz
uhj16O1InYm7iZpwqV4nfOG+1uK5pwdAWK5NeY/BdFx7fpEfUMpdHJxax/2jGtApY6UQacK2Nh4/
UEGYZWpnqhqz4+Ucgy17okBPucJdP4rGujZtcJ78vRXNKYuWtBe67A+2n67cq3oX+uzQFCXIKbrB
7/+WiOmvslm58+B4zcdyeXybK5xlsoZ+128pOg0TkTkpA6fY195E6noFx40HIPCsr7mWj2hI7tSB
AkUa6vSTlAI+0I0Z12K5il9bRdYzURlUYbtiVsnarcpo1qWISRNTgv7wonuIA1ETOpcEzVoZlK5j
Glf9WZu7OB5aWA3SDcE/YOJnb6gQuwNmty32SC/13gjHTdv5Ip3Ftf9KQGOwPyqfEgQIxbFbvrdo
mTZMd8B5LJkw5sktePwb1I1qS/76UZSamt1gELazDbLYW6dQzf3slT6MDjbs4HM5R9Y0FZMRL3tE
gTthHCN3BzYJE4yiRNlWCuqUHkxH//znb3U1yzm1gDlxFmbUfTX+vE0jd9HoVqIZL80aHLpQEvBA
8jsDwaVfSK0IlF0LXAHhngBOBQ1LaNHtfyle3ZmmSGuDkgll8XG3cBuskQWP9k35wSMbSqwx+nK8
ykozAmWkgo3BVsF8SvRHqSNdeVizgxf3uYEUBzACRvVK+oSOQkvrVkfROeAQzdynQ4REY3SDtVhf
Y2JetVHwoF4kmLc/fb1oePiW4Tq9M4Qv0trUfnYH/h41bhTCXr+fomTtVn/FtX8zI6JdfrcNlsKM
HIA2pmg0h9049VJkGDmg2eAP2ohNqIOvjSIOGjqhbPVbixkdYaIDyjg/hyOVfAZDsSJ0qzKdVERK
W6YBb7iwiDG11PVmzXdTPFiDf8CYeCLo+5APsiUsWKEm2dPAEa4LsBO0eVsf62vkswG7FhcI0Geu
wFH9R5ePkl6ee7u3gI7VlwBN0kDl3ubYn7rbZ6gGr5lJIy9aXut7T+Mrqpft55bqwtP0PP40O8GF
arzgFyDDfC5t0+zsKzQGnI75RJe4OE2vZY7Azb6P7GNwP4i7fuPbHfdLZkB/3kXZFlfQ7bUq0zQx
DuFSCFQigF6kvJktE1Nb3RN1O6fFNLWxtrohPmTS29lIkjOO8pIYHfbemVko2QcD/SveIS5/Jh8R
ecBMc5Vz2x5SHm+4RoPuqEH8m2ctUt8e51zAxyydolgDCG6fTIJp05KAVmY1DZImk6Qmm9IcEueW
vjL0z4SrwDLcPx+QLAOl75bSV9mLKuurnRHSEXYHf9Kus9X0rUk1YLEcdFSQF6gqykB51llvd4Pf
laV0dfWMbgddl10wq9gsXiu3ZmMqIk2z779wyAVlwT80D5DRnHIZnG6t8PeSyriF7I8/71zossuj
UrFg29mENIyun7S7Zn/zbKRhqE7lFPthz/cTRbYnCJ+kIGmqy6tOD8EQT9caQ/s6fY7TKHHE0ZnY
vQBSVKFuQIOXCQ20tmoDs1J9tbw2wfL3ry/Xnhd08RqU82v/KWxmA0iJoMm2APiWJMmIA1hDxqNK
+q8rJ4dAErlgCcl0BoxmEQ7rpfZI773Tyyg5dCeN91wU+RE5oGiw9BLu4Btxxmf6ySYbADhHC2hJ
oBXjTBTolfJynd/9enAuHAK+ahCyL3I3vtaOOXMpX+BzyvZ0Y54mY8juaragL3I7/igzmmDg6IpX
nvmkNfmUb3zNOMCBTBMDytie/zIU/3/jlnNTDbrstEgemFq5lWUxwLu2srUKl3GvYgFWX599A/S5
fzdHaa1aC6boJYxNCqFBlbC8wZv7jvXqE9TRW4YnC1Qj16XyFNUZb/9Ata86O0PJo+MvFMt0mBRp
kgMwU6AC5tjYiD8Y0NPzTjA+zwpQZqxVz1nuv3+eg1i5EtgDCCauyo1MDTjBXmOJzllUiKoUqzfo
xVFUS5xjR46cxhS8Z+mYkAZP3MBUP3f25Q1FQXVMimYiW/AiukozPwHqLV4g5eTolFpMepOvq5sF
t+i1V1zUn5p6qLQWUH8CRzUy/OoQRGV4+d3607vXSau3Z0ywt6FRbALre8UarT6pnIGjVJ1ErgZ4
kqaEMbyBPjSA1GZbKGKfBniqKwUisuDPcdQXEXrkd8X+AraHc63IJhiHgDBJib+kJUFcWadWJaig
HIKWzGcTX1OiWbRZXvUnOUy8OU/fnarY4pMFJuO+W4GSd98xRfq9ny/wDeshJE3eXbQW3BTENEWp
sg2h/1LvwaR0xGVzpq1G87A3RUawVOeEc2RokC48RVwTUJadywtcTVXZqjvWPvnIX/h9tNfBxBnf
J/jyZhF0HsunJG/U/bKqES0jbkz0/FyaJ/M5qO05hNAj2ArTrkEddVc6lvDCw7OT0bzreEtQa0Cj
4wIRB1+klQUDvTVS4NqYq/cZ7kLuBZRXaiGeQzr1X3uysod+vNxJc7a4jwI2uSUs6KggqOiK88E/
jhoBZc2Jaf+CaW5g9bwHYq8XlYGGNhEnWDJ5GROBIsOfOQ5qXvu78YYIF2rYJ4ATuHicxFr+1VND
D4tZQqsJjNOirBKJE/uuTrYjSPrqHj8IN6OLGwwvUNFrQxMBjr73M2AIZhTxo5noWufWkw13QxTX
Sl7J830oUFVrGkjdEWT+jwMg23zQkKzCaqJJ5cgxzb0FnUhVhp7ijDhUjmFlUyLTyRZ353r1qMfO
b7b5Ys5mt4rtQK/UGEJxa0iZDTb8u4sbKMlq05KmEJvlLeJ1Ml/47HgXhHOEX8DkPMyQc2DMmTWM
c7UIXFO1A6EonjT3WodXjE1aOQh2/jUvm2H1AHIxG4+gBNJn9mTLzPFhgww8LtwNBbBxLjYilsC2
Blmlr8aVwgCTc0d5NxdlSyXjNCg+8RqoTBdtDZFkBb57FPsNh69nFlHobUYFJJ2BytE3X8dcBbOO
PpGKY8SIlZYFir0EfFOV9BQgcF2vI89jqLWWpWeab9bjR2NLPw0oF1HsxMSgPZKh5CmAdtrNW4el
IxRei4yqx7qm5ybRLt8cufTWnXC3sUEPehiHLq13mDdSUKYOI8dsnQZSWI82N0iJFxexwzDmD9UZ
JddX9IxgyyfCDfOlVpXnwvHvg5h+qBtL/KiZFb2CJ14MzP4dM7L4AAUsURClj8ODqjnVrVw282Kd
8QcCmKQz/FA8LmAFZ/fugw/gkCn3BZjjMjRxyq00kcYbpvxlC4OyzvYFwzRIs1FLIs0UrJc7qPQ4
Hl7kRkmN7TpXIT6bQl4UxVQMaVWXqwGbjri94t8YlbRQBOyoIi+MbqxjHFphWJMub5r7fs6zPOyI
fqNeloduPVHAqK9Juw313uMyarQD833LOn4IrpqIkmDXazE3fvMpK5ZT2gXTeZCjv+1VilbM75yv
SczHZmhfKv55KGIzs28eaQdwFJl3C4v6zn7M8XTx5FZMknt2lmJ3r7C3ylAnqMrERIrW1u+BfYTa
EEhzjQaxhgySFydR6q2LBOKVcexa/vVQ3ygSahSefzqBqlMqs12s3eOD/RnjUAaPCvociPF0D2qD
jgakcWj9jZC8ho6dizAOna36JwAinDWT4RRciJZoCv3bIZFTQzSnc9hSl3PZGb8dEluqEOQbZbqp
IWqc5R6dUBf5h0rbWOiyV5G20j5Y8NDeWLJMrtdJSzUb69dMlAVaWdi+UB1K0bhHkLcYAYZOMPS/
ZSEI6BX2CbKqnPZwV17XmkHkScBvPTv2Bcs9XqvqGIP3RzMb7UGVn9sCk/YebUv7yySxHALoJTkS
xRaz1OdiX6s6lLms55F2gWdCI1Nio55lQ4cS6wOfKmYiVf1BJYBmFwm1OSar8EBFVwQ/h9NtkG0v
B4uDfJBA7QQdhBTMQblOyIAzN2H+pkdDOxl3Mz7G6s/ZklXXxhSDCi4+WWTwnVsyzJlossOdfjo1
Qk0Nr67zkGa1WNw6/ZmJBcBoIK4OgLhKlBDav2jKBupEZMWB8OnkNUsMWTdCOukVaFOu/icxf4kA
fJVha3QLEVlJinOdZo5imzhQ4sb+as9J1uFqWWAeKkAcTfdCiDQcJSLZ1UcGWAG84PlaUBU+yx1A
UCy6Z/WPRuOcLG6nXX156xGiLGqlw6WerLzu+vk78dwt+UAq7MAE/KZbv5/vjz0oy0dG0mIbMEWS
noznHrneXnQz2X/XyJkhz+m7GJd4PoySE1lZgctv8+wEwqJufYOv5eWbGEaAYPzUYBbjJ7NiNT39
iba9a5y0TRxpofgyKt38G1xvY9WTvOWxSKcUHwxliU8gNTUAjnKLf4K4JTjqxIOoNhXrCX8bWa4d
gQvGcb+7OyTpr7cfqrAnX4AqzhIAZIiMak1Mij1z5BG7u2qH+Hn07YGLxe3AVQw7DKImaOqW8i9Y
ZMH12jp06W/myydRZo50RYIQPZ5lwFu/JqF3t9uS1KsMe3k4WQjlRnoiIkPZns8/7mudlJesVis9
aSYNl5IXBuHxkNYKHuneMfNKxh2JGLZg060USk3Qt9G1qA29sw0v/K0CvIEstcce/zhtgy9oI0gC
ij0Du6Ht09/ifH+NZfVJWC7ioM0IEitOP9/oKc3sI/hktKPo8X1jv55W3Zwo//NdQnp41x1z2iyo
ozW6GEMauzTvAQatptdA4++HHLH4ql9BnkOna02gEpJX2jQSH8qa114hRSNAMHR4CRzd+osLbin8
K+8tfHchrBqrv/+1okpbTmJVfz2hiq0YMoIIvSPXPJfVSXY2fTa59DtvOFOJ2O1S57dPUSZWoRvF
EWC+dwL02gYtXnMdZiwsSef23kJKPlQYjLMtbFUH/IlOqxmw09RseIjuXC9NwMOoDNQCClBPjQDL
RCAH9+KVzi5xPmGwtOVq06+kMTzX/nfNwktemOOTKfeXqr3svH/ovKfCNDEZzpF3Wf+TocZ2+KFn
Mjv8Ss/8bqBCR0gWWUXnES1xAIvgHPrsVK7w0Y9qubMbvJ+rC376qzEcNj2R4MLmNOrDRYG7w/LA
ErXxiksIxkfZvTZqy2bMibHeKUBOTqma6XRC9OoNjQvvgAvIr6abfLEOdpMf0n8NiI67bP3BRQPg
00dyQI/DlNlEXUz58+kLVFqobrhOnmh9/Oc1dj4Q9aqv+MfDJ0s2Y/gHY3TmLgfJE/Hwa7g9l4I4
kqaj+2hgqdCByfprSa/noXtucwes+zh0Eo37hjJQ/tTq2hYO461l7UovFPliYdRasdEdNlpUY+EL
UGKH7XUxvuJvER1DXg+UZddPAqN1+tiwVWiANghcGj1ueEhaGK4BfRqsrJc7Omo2jF/Qlg1//lbe
jIdC9+yzctTbkjcfXktNPvO3Z+Acg1h1U1xAhBp8AljONuyHwlqNPI3hBwEr1ja1krVceCVD0a8/
SwReffq9gzd/N2VLCiw+GyODugm+n5J30xq3+PidManB2kIpEySjwfZxpvxCDsT2/EjP2J5ckrrH
ZGYJdWgwt4riJkdQV35WB39DjG3jbMJC+JIwqJQE/I6CN4a2Jf+auND9vHIu5/GLKRbGStK/+GZX
fzEPhMwJWTPjXtGXrJf8Ku79CCjKC42hOenpOj6KlR2SOyY3BCmlB4J4L1jTkBrzJkvw/GPuZKKn
bmSvVEqhnJaqQqg62nWaKeg0rjZGqmpTWpzX8L5MfS3dLcb/x6vX5CZVrED0wAJJc211zGUb59kS
UeDOuuL7kvy8TWOqRyv6Amp1mf6XO+N+haLLjnKnr6Vodw3kqJt6UDhZZ+8Fnfmkl09Stshbc28J
Ww5OWai8UI09JyutVt8YsaWaegQFYlHOEWB+zwKnnmvQsUfU8yNVRR1hJJMR/h4qLDx3mbHtJybP
QdEaS6gFY1OhrIxMbqJBDWL9dXJ5vgdARxciFfsPgn51/68NwLzwgcGGKXseE0FIr26xvnBlRLXE
wL4JJAMVCGBOfbTO/Swb9aNJaelxeKRb0Y2N4/1JEJPs7thPY5jxMbjJUGDEe2jvm8OP8qxoX7NU
50GDf44WyW/qW/ipUEeH/6ufgcFe01z82v9hOuhX13fBzqj3Q8DhMmn++zwMFTM7Z9MoW/5EN55Z
xSzc0/ru262AUHrAoOeZj+b6NXFDlnxENLYp8USOZDDlpA2SSCWG+vHsZmfzqbwMXoClAOUJSxvN
lEUJLyw7VpGVC7QKcWfmm8K9QOfS2VMZ7kcurWcJszfDs+1VBO3unvlxbwAeoKhOTxnQaKua4YLU
GH9Aj2mlNJmb+kKXXtmTMAb/X56hzGSGjxlxRnxRI/4DjGv/S3XR90rrJCne8DXVu9ZOvUeyvw66
N5WSoaHsOHmew5jWJCyWVcE+YeI1oofcH4u5NBUuCRemA/f/8qa5D78bZqog1DOCK9+Mz0fKZW9S
2z3nCJSiTKEE2OWxl73Trv2YLHQDJSw9qPmeeOgAmSEaJh7zpDGOuWIWYdXDFl7AFLqvYiHmm944
Pa9sE691hBNeOpMul94p6zikpanEz7yqx2hpueNb9htJPjYtf5gVMRZ8J/Kn39wO7hOWbcHkbbGF
15dzJ2gqdU+dmzcBvq1QRryn84G/c+JOOXd4oADcd2P1TQVZde1VBr+YnSPEhqVtOdE1cuWbI6i4
A02qQAZIsgE4RjM6vmM/wXwxMKS7sDqO+O5qJMaFTYVrQvIO1g6rSuy5IjFFK7LHxWwK80E7w2i3
gRalSCmupwF1BsomixnRMtuNOG8icamIGZlHrrNS1TJ+PbhjLYa4AhpFGgLi5sDKiHf082nVBq9/
vDGs3gObwC+LOS3U82VT3i4LqzWkwKIIMmVWHvREpz5u6G+w2le/o6ObOBq1nqeHWCd+GOvjXoPI
Z3yGCV9SALhAkSX7usl+1VcxaTv16hsz9vBVXT+/BE2WxUeiGTK4roM/aRFNsxlOmGt01oFtPAoN
lGah7ZYSbHLfh5KOCga0vrx1A8u3brYALOfjNtAHCUEp6jfTioB+kLTyI4cKsRRQxoqZOIcUxpzL
qUUMvqYWyzJL5VbrS5FZoa8J2RtDRqkgYNp6TxL0mjttTd8TiapB9yXvmWZKipBa8NpXm3sleXuG
Jwz7nkVbEfr6KJWB7mubEp6am/kizmbInkI+uGcZBxEjaVfE83brcmMfECHAsOk5I/5H7tgVDZeT
FSgZVoaTY9IT/GTjmuoH/Y17ih3c40hIZJB7ywdqgi4q4AO1bm6Gla570EenRhOSV5c3bgnFRXc4
kRYfxmLzdT9tDsZNFtNdP4UkL3Hqt3nAPqE8Ueia2YRZUuGavrOoUt3WanOeJaLsDijFBVDDgshJ
WKYXmCe49RsU4oGqLhKzYO8CS4NYwQg7Te85OqYClT/buw/IpLdSzl3xSx1mgsFbc1IfMbaPzXaQ
05pKgf0lk0AajzsbxIehiyhUgJ/UJ6r4QXWQwf+ibpwZbUXi1ravnYM2AXnPyOb+tUtfkNROQuFz
0/uIljI1HYssZ0WhZQJ9i1V289rRGq07dYGZANOd3/gSRO0aFPTvkDarN7jWMvmYfm57Ym3KtUCJ
XOEG7a9CdJpW1ZBxM8NpD9WTUT+A6Q+R2HK8oR0OkXX30TEnZ/KvhVg8l/UZp6V44aR02dnt4ZsD
4ma7gMQ1lBTXDl1dbS7WxzDc1Imuvfba3Da90ZkbXbtNUru7V/7GNrESP/2MwPLPhdlmkrcUTHV8
TBh2dzuiOs6cXRETvNexjUJqiJVtlUvCxOCaNjgzl5Vq1qfI8snR+avc0jchbtDRV2gGfvKw1F7h
33dxSVc2gnjBoSAUruVUkUt+2Y88ceTGBjknKUknUyPGSEZQ5PTo4rt88pyHLqmj77eLmd8rreHE
UUUdQ4Tg5hlTzL3i1PM5EhAGn7IjiU//6AfSvAcSi3vyFLnXsoNfkmTgZb4j6K+haDOTILcZEpM/
hUkYwOCL5A0lSXTv/vO+CTaDHss8/5pS0gXpFUIdJfRzC5Ern5Fnvn476SfWqLh8QoXaLXp6NOnI
qsDcJZdT1IT5bQmreVB6OVNDQJY1TM1nczcjuTUJTUEegJQerNzusCoeVhXypqCkM+TsAWiN7Mtl
7ZIazBeZsgh8eg9IaUohA33ZxYYbC5nK8uqJtjrsBXGSPxJTwu0H4Gt629SYXpy8EX+K7od+3e9q
YvienFmpRd3p2vTj7UuCR25/XWDeDLWIuabEqlQCXAvUx+sBLMGcAoPsMIIHJ/+Hn8c/E/sl/YZj
bHGuMyirurnOvRIKJQVLw5ya/4nXfD7Lme9gqdDrKub/+KS+QjaHviRDCSoIh/0O2hb/Rt/xdL2z
G5PT29kxBZXkEeS5JQtOgjid43NKkJjIyUU/3aSmXq/WvFfza+LtIKxOBzySC83Xwvwd/9Z3o4Ez
MTL1rzhraIO1Qb94ulsOr95+4Q4c4sCnuu4BjV5CUaowRwAKrMA5cUswrkXDbEIVONTPwEyQ7Faw
aT1i41WwlYyYDS1zlKDV0p8bZIyHRRO5xUM3ZAKJULtWuVjjrZEAQosRLD1cPEf2dkCu4Sw7ehzK
TH9J15F4hXgFUrQj3YDzvvzAD3bo6eT748lpV9L6GS07ONl/BEFDXb5fnpmGBszcijW81i/GJudE
pI7JBTFlNRYZxKjsBrAXapkLh4d3YVZv3ei5MFYHFtP0clQnma4Gr3uSftXYcriZ89Q5GW/JRWg2
uA7vnxBbP/lijlw4Dkdllt402cmGzVboPWRnPrsoTrFtEcfLyW8hojtzz0DXTk9KM++kaKE4VUJZ
oC/vgN9S5UChKrT1XuGOLmXhcByEXZWhMPhhXYcG0lRvtdw14ea91bSXr7R7QgBpoSoGzZbbuOq+
8lDZlRiO31CeJsXfvK1i79WplOo7DUE9CUVNmgybq+6RYRVmCnKCw5kTfgHqgh5lJxL5mxZxNWjh
Kw4dmnLB2OYBWhne8zMKOlKg1e7XeiQxXcl5263NKjhmRXwzQd99dBrQaaEbpCyrZfbB7NdAUtxO
bRAEMiYzSZUJrmG2cx4AmzpMj4UF81RuCG/FrJxybZSdhldzTeWP1g9w+YJI2aiy808/s/wHRfXf
mwgg8ysIDL3X6r7DVLxNu8zNnNfMX8SbWSEOscAs/Bnj+YPOZaRbYMkYb+VoBQbu7ekcaJ9pCV+i
qy3ptp4z092qM3NWpvp6NRLq3QWSVwG8DxXumZwrho5AoYFBi2IPRjRWCc2jIVffwkH+29o1BOSR
NY2SAhYTFcpfbydSXpV2ckBG2arvgah0HqJLwEkb7Sgafhh88IOGSIR+rh8HVnkofwygS8wQT9yY
giy9ZijT3r9lNVrRdUQimh7+jsIsVGLLtDr4oy8QBwP3nmxDuulJ15goNaU4KP3w078K4gip7TOb
icI7E9687TvWDge5ytlsfk5/uS+8fegtedgBUDksA9/pQVtrlvwv64hj+xr5YLXk05+8WCHJnqAT
JZYbFCthlz8aQe2oqEx2V1RNL/cJ+VMVtudmdNLAiN+Qdb5dFnh7JqidbZwmi+mfQ8qI18zQ6wC+
tK7hPBZJqNzer6fQCo2T9QOk2GJ7L28DA/Hankqppo2Bnt6AGC75kQJp5QXfd3bvRzy4HTr+wW63
72ikwydhEJglWWrNmKXqi4SzynVWP341IvIkuDi9knduKFUfwOi281eoZ9djplvvaDUXF50ZAzc5
rylsN4Q6EIhB118dXcEpsSW5sBLFuYvZj69kZBkiz+3ZtEWhX5peW8gYNBlFuLm2UrOR07NPBW/D
NxjbLlaX/LoL4TK38hZj+EBAl25VnvkXqZ8aUiF8Sg0pXYNm2Mj3q3WqYkUBYB0Q6NpPUy3sexr4
/Bs5yHv9vtezSTGGONYIO3mjs8rRZI3zFpgzFMiwZk/GyLahncPuLxgkJnok0dkflnqecBIk+8hp
afVSpHRfVBG/KsDwnQdoMI9sk1HsHfTIwaThc3BrqadoF8JdLtkfIfyo6Rom4zWSveNevoV8wOu/
Hqn9R7TNTeOGdiv5Cw8iC6RxhSYTtvfmiMBiuhiKppME/yGM43RBAUwcJeCAk/tV2OwcCpW1edqC
5sZc2cP78TpLSYE7x39GhS4ZeKOW54vATy+uoUDKhmqOUaHv+wniKAKmPSrutfw1osS6P3Wj/93p
UbFvs2j3K/tNwrn83IK/CrBvxe18/pupA5INIae8A6EpAQbgiq9JGLoGZKRRzmlnBpDphvz7hNa4
ttF3CBTIuh1wBwLo1rhub6HIxSSXwHSr7VlA4jh/G//jCXaBe9oKsFo7ElsOSPckF3RvuAoCsHMp
73N9Aaw7EFugGHGHfPUgqECcgT920NYvys2rlOBkVWf5hxo4kDteKD9QxhZCR+YLqyzz/NCbOuE9
RCvMLJU5AXr2EJUY9NJHjZ+7qa7YGjrC9Ku/78AsqnsGFsOI2ailKHFmjnOvPycyZLhm599JctK0
tbQJ1q8S/riMabtOSUzWrOx9u3twkq+f3SVtxJdY+irjLifVy+q3XHbG6LogygqGNFyXnivafO4M
k2eV8N7z6PZADkw6aLdV6deNjj+BzGuW/zEjVFo3WdaAzr/wugPtpA/+3u3qt+sm8vlhM8m6t/UH
TVMtKb2a/FeDKNMkAJI5YP8bgDbeazArvqMLdzC5/BaZCriBUEtK9HarHy52BA02dWSWGK6qbht0
Bigs5RZCsY8Ccei9KC7k5knk7fuDsSwkvXuolPKjWq4icr/Qi6o3hdgGf01D/9z+badRNUb+rzwk
Ye/rICe6xST/Wrkvid2rj40VgfeMS2LXdGCsIo1xbA2Qg+zVZkQaBrROV2v02waMCxqh7f+IwzeU
P1GGcNMyLgP/CGjCkHgU+rOW/gLMAh1lstPgR/3R1HYC1u6DD4NMBfTjUZjKjrZSmOXn0IvY2joS
eRBPJoHuWM5T9u7a9pcVEJivL7CaNUv1CKLR/q/m1pijypN6LiO+CE+OvgDJmpTz1c9KsX/b0bGg
EgW4ljqKNqgyGgSbhfq45Fn3VgqGx8oavXbDrm2MZyuTxPLhhuV2tme0YMYbody7E+MDfffDKpgY
sth8QcVkOR8eSh0+0NZ8fDthmGz/9UDW/xYqohU2fcjGPJAuDEbEyS8g4Q+clK34WYUVMo+lOyBF
KOI142dbW7uDJkZsXasfcbjpZqW9GHRdk0jsaviZode/maZn4F0Vx4G9ZNglzSfUNHUW0pTUaSEC
5GwrWPZgcEgXQLQXy6EbGUtjVowxETX0WCscZbEnVm4I9BVvF7kesEcq3bVnaFpuo1LsXHgygcMT
zBWMDzalKLBf2+TPG+QYrwlcMQ4f++NnSCwtpEm6sJKMsV9ZYET9kGC9IUI/C+9p0q8QMQ/DiJjO
LmR0d1uxUPPW2PBbOsgI5KePaB0Uuh4Lj+ea1UOkCi8cJ+TIO9DUwCxy1Bj+W82C3j4C9fSuPpvu
Nm9Oy1zpfGoAPV2OpARlRPzW88uX7lUD+istMZDUIUINL8/jDGf/1/TWUNcvCvuGyKUJFsuVXdGs
433fIkUtQjIlPeHa1BGAFBbkDbqLTMGl1Sq0Gea3zJOZF9kNZraQe1xp5mEeKMGlWtvLwD54V1JG
dLlwi2YUlzWhfWMi4b3JS/FJhKX6NFb2ZMnB6p53PCuQc5LKqmeOM2YEgLIxXKHt9z7/xL/G1wxN
V0wBismbYbxZRGiXMN+GGUMy7GSlGj2Z4YrGYs66VvslPPto9kOFHZrAlXs6cibaCQLo9uqCJtlL
iQeZmqTITz1FIOxlQZA4/36L5ODCrq0w4SK/hF8JR5wlNjEXZgpvWlNt0YGBAfIZvo+fZKvaMMvu
S3E+rJ48k9hwPfffNH70zgtsdLqlz4zddUQu1EGwz96k/zFZXEjHyqnO2YT3sdffESkTBG61vCoy
0Svo1K15v7wqyj63jzjlhcKCFefXdm/LpIA2NbJQfMYSDAXhMEPKMgJZLeK3lt9iqnt0t4nTSzMM
YN2IAon6JoF9oo+WXIYw1WtRCiW0i1kR2SfPaAuwpuneS7JixDiHYxPaeDDIopkYoVehkTlVwdW6
BAOCYd1FsyijNDsAxEEaYzWfd1qoyTvyLND8/J/tbvdr+Zb55zwg+W6o2wFZMLHMNcTwGnDv7SRd
/5mL8U3oUmMPZRRerxedGOwOlDXY81J/PRZ7BQ5rIvh1HlVwfJNkG17244qirAJEES2JYppHrAVr
+khlptteswpwxki1iVs6ngCmbl1Y9p+gu7HsKdGClEYziiv/zNIYu4yvq55i+L51NbLxVUThtGo5
kf0fYJCg3M3mZXLRBwYnG33bMEWnGwQNtFf3LE4wC/DiqxEBrpoEIn39Md1YrKzy5pxBjQl83r2o
Bfc7tkWq3vpGSDsQHhahhawAg+IDp6jHKuU/JrVRQD38SVFRDcoC6ScmQIwFZKa1Hv1fZ3Wrx2Yl
KnJigkGL1IXd9l2je7Ge0KALth7iobNEt7Kdl/EONuaqazr8TnzNjXYqfLSf6duMTMoAcTKQlWh+
sMiwfqtqGDOpS9HdLmO23ofidfgIw4A6QPO7j5x7FQ8Bk07oE5j+qt+qlOXMMGH0IZ1YtqAs/1P9
ss+bwUwHZvhmUmITNa1Sp42b4jdqIcRJT7CWe7yGi+LhvSpC/b9QJY4HHDjnmVBSXapTKKa5vjN8
gXPUDGV+lITj/Cr+eGel11nlT6mRB9UyRQwWQNjAg0+coiDUrRvrFfyT9vCfdlzylPSH97NlKVFI
JtPArIHLWYsu2yVdvUeqcViwrebex1j5muUzot+ggz/YliBP8JERJ0ysUst38O6tVMboyHjpOiDj
dhObOCV4UwCJYZE8JpMxbSI4wzYeKphjiP7hJ1RyauU65usOxPjsAgydFqviVIwHfjGtsRj46Y9q
fSyoMsXrpRFZAN1Vo5But+wCUunJpUI6WWqoq2NnMdFcgwNt2coq7gcH7svMbGLE+6jnA3PbGhg+
43X7LN1V1ZpVn7vERlz3G0fTcW6+dE43aPRUG5tBQwUm1O5D8a2GSQBnbYrKmMafzwwUH8n0IxRF
oJ6B7febwBNUyZef69ZBSAVqAU2RY2EjBXlcNbe527HpbEoCOa1MrMmTHAZ0bPILn4GGcKkeIDrk
6RWKCoeE7pwKCn58IGAkh1Zi7u5Nyaht3oo5nOWDAk20Ecfsk0GYluyeQJslCLKz+CyH5c3161mN
8SPy66L7QSJc+ILcW4yOo8v5E8DrnNqCia9gQCftGTUhInNTFDNFSbAoQ03+JWcncRpgu623XHA0
TfxpjdEIQAqhaeprHgwSdBRFLIm+9ZHl7TABoZfNbS13ZScRPGWcWH8QWsr0FfCUBL+kXgCB3qBQ
XuYlEqJTxf4xgg+y5xYSUEuNpLxKPvXAyCyn+82NiTczlVu82+7E+es3A5BizoGgcaukqsQ2p9nj
QXWF6yS5hSOUrkmvhk9eNpkuB7CmPQQQf31BnapdlN+G5T1cq0djy3rfnoPmc+TnZrHWIODMTDkv
lrpIjh7FwjQNBoBb4qGVJ0n9DfI7u3UGMvve1MFZVk84IUosv8io5L86g4k4TSco+zRj+D1ctdZz
fax3VkV8obj2H7sStJ7Xc2BlvlQeqI78vgNvDIRZhm2vpvC75bwVAvWJ+iy2zJvr3KBtlWlMG87Q
Qi2QK9SOJVmGFhrVHn3tKNRGljhY3VJ99l6q3DJOEckoBwD9s9qhOMwSOhGFkjpzP3CWjapjIgEa
kaEMskSXg0F6+QATlxO3pH7r6K+cixyOOcWqKukPk+SzeIeEQMlaq/e4F3AlRAvHhWSGZQr88am5
KSKmBlU5RvqeOnAAiOlLxzYr4jlI1h+PsQravP3Ww/Dgfj5KP3OaKq/i3nr3qhXIv2+shJmeOxsD
rkdDR8OmAQogZGnm5XnMnMvS3mTSoXJr2qoeJ5uzECtx4ZzOnq+07qeGzM4xmk0KmZ1cJunzPB1H
SzOzfSl8hhyBMyGVkaBaOaftgjr2taycxN0CBGe/3GI/JPC0s0O7t3c8ib0hq/jdmF4bFzfQG8Hy
m+Lq/5ZowDIcYjWqyPGy8BYtQx+PORGOi+JcpOdu/CwCwuWar7Lo116/Rud8KVuHDUs5K6Z469qA
262mdJToEpRSz81rPVY+UKOy47WZtmmyBCx5N2zCOq1W4DVvNYpHJISc1+ecLg8aAoDPzEZkLElM
+egFDyokAvIwOTn7cw6Frsbh8dbBrgjPFsDWFrsMjeKxwlbeSMa7rLLxi7M85rIkB9KisolWw/02
Unbm7QS0GMnjcRq7FYuO7q2TiwLkF8YJBbVmE715wv3Y+meUKVnUzvZmaULzMCKylvGo+qjrX65H
k1uWVoZSTVizGDTErLkiLo6uBNipw96O+IUrSx5RjoxGTy5OD1gwvh777+Xj9Jm53/5/kxn5ORE7
Yu3UgnUhk0Tkpldf271wTkao5cSt0chPUkv0Ra279wPCspFkn0oJT2Ns/RZGb4HJup5tBp9xlNIg
Bnr6t29WNaQiT7xrLaegV+2g0ITeXkwatEOxDrpdjmGqZnWryyfwAUsYIl7WMVy85CQtw6AAbmvD
6AZIqr0lFjkQIGjhyBw194XT6la1g8Ow4V7LNS1cfL6UmK0hOnccVbRBQTmZD2ozswnqWN1mVBo2
zzuf3873/vYlNWg58a8d+DqFhiT6tyRuAiONixZoecqY7szVtaBw7LKJlEF/iZibQeetQV6ABHsm
RrPLNoSM7zFnIrgpEXLuLV/7wsje9LgqcQgKaYeoUTidNj7GtdS2iOLkrBxPHVSXmUtnnPWbj79e
7v+7peXUee1bKljLVMrJelymQFm9M+08qYek6DGB1tww6h04Yunuw9rgKVPc7WvCWw0oylOkEpVH
zI9UtUjPIxyCypxVvPx6Dur+5+bCoZVb+6oU+fCnmoO+oDRrsXK0SVLVRYgsxReNdIbQtItBYkBn
MuiIT7PQiyfqsjBvc0io+K0+qkXhIy/PoxddyNVtkmXW5og2hi3O5/mh0VHsCN17+hUWeNp7u3BI
E0mlcm+iFHwOxMZCtsMznqWroi7ZSKpCpX1ISFug/FWF4U7YREjhfeWqTNGPSZzm2ojfqlYILcwp
kfCNVg56Kso2fMkocFI49PxTB31V3t/NQAfvgBTrRnTRVXjsWoAjhAHsk0uLhrycieoNGuQFtxxr
1SY2TL54IZiLB3f+xV4kKK8fKomi8K07zvZuCSL9XmcfLJLYL0u3AFq3ruJI/pTs6bqwmNRVVCLU
j0uK6MKJDSpWlibQqYg9nHshVC1iXa+wzqDHmSaWpoUJ0HUsy7bUjIcyuAqHUWCWy0t5AiEx98uQ
zyHyxO0lo5pX6uGlkHK0R6F0C3hW/pF40LMZahtKZ5i7JZK8gp/1V+Qi3UpVJP/jDEKKuFtOhCsD
3qhstFM1eSNgDzlvxY1SSRvhm2NHVBZSQOzK9ins3HGrnfXjzA9ltFiuk5eCDIQtnGijeg29vdaJ
fjR+X6rqtMMaVQIrFSu0TKcTZPHGqxJc5IOuT/wdZF1GZpWTo84J7a4cyj2sSb9/WbeAmnEECycY
6s5YKPStLRWqGVXvJ2coc6XorKO3/OHrfzI387WhdppLperGl0FaUWCnSOOk8n88UH64jD80K2Ce
lpyQ0BUDe1Ub3b4TQmqAdoJ5yHUlXJcZMipTFycbMY5cXka0EzZE0l8/t/jmAjVadaIm4HQB7jwo
c3c9nBBDA2FBy3nHO5bUju4ojBCJbHvruTG7UfPiC77k36VQjYQkEVrC+LR2+EViXSDfg6HP4n4D
/Ntc8xrrqBVxAlWVxkTABFsk6Df4klaSbKP79T7w8Uy9IMfi72tONSf65x7/yLsPNZjA18A2BOgl
Jonk6x1PcOpF9SUihP6kJ0KtRxL9Q89VHRLOn3PARrIIK07I+eAXOhvS5MbZOdruQdpMBj2HhSQU
TReJ3T7au5U7ac2X9ASqGMucpC8VBGHpN2c4BswZBMUeTCWrESRd/KyqrG9bSF+sG+fNxfx/th/l
9FK1BjhjhFU3XHAOHEZSaHcAPMqLtTzkqgwNGNb0G922TLHoiPh1ddHZptZeWego+cdKIeDd3sj6
LQcbrOjTkNi9XPZbk8j4YzGDVj0jBW6F4OotaCh/XEl7v3b+g8ZxPoYLFfuJNwC5JYtnH/Suwyzv
6nSFD5HMG3cBqW99RtesvpkMbXW3nFaAHX2Ta6KwxT9l8eF52ieieiwrNcs6EKsvnBOy0e4NEqzr
3jdVs3kdtKHxOay8hVXiBbbY7HUCS8kwMc/4uGmtQQ3Zx7GvgJs+WCw+2MuNSJw8I/8yJmEKh9sD
HH65Zm3L6E6/S7Eryxl3XAXd97LRW/a88GFRJb+SsII2u+c3Ro19loD1dhrLPt6pxmvnV4zru450
Rg7/+3y5fr84obz5XIA0ma+mAzYEmx2f0NnfFovdMeSXZ/jlLZYA+1i2AmAge6cQDww8grhs+m5Q
80a75pYMgMzEA59aLg4tIzzdDOfGD85Cz2Y7wCgq2Abp2SrknOnLeysleWTiY0a6gKeT9W8JiOVD
YiXmCL9yNaR+7bFJLYbNyH3Ayc+oM0sWhYWKrb+BdOIEL/Q3JeYnKWtC7689kW2r/32BWQZQmlGz
JF54Hhf/GqATeJy6/8FjDHyIynTZIf4edbKEK2OghHfLo48M6ZP2cuUZhysN7DNrnYkzu1KorAli
4cD8pMLnTTWPxGcMqSbuouvJ6BdI4zeKkqSaMV+swJn56gDxfnF77wOxgGU0XlujGtjoUqDer6mq
3fROse2YGJvh/OMTroTqsqrxHa7PmcvXx8k0uDkMhE5wZMuTA2+soHzKX6QhqFARfjKGmQ3Vxi4p
FzEhdHLLnw8uC7hRoFxq0FHmipSECK/bQSkGk1uOtUKNkB/Hgh3Q2MPFBavE8whh3QdKmWuQIstJ
iZoOQEyVjPOEZWioQ2oVskyz7Sblvv9T7vl25eHEFdCO+wAUEJjl4juq3ho6XTFV1LdW7cdzrEfY
J6Me7iILM/C4usTeasrQ3VsKAyVBGVZ9oprKXVN+0GpQRPb0KKR61k1BRB5wsABofzelil24w0Z0
anZ9ep4EQwvpTyrcIZ5LJev7tWFGs5iewvS54cTVR+dhMbgWSsVrlBvvs5Q2uFMpCumImSt/hGwG
WE7ayYyEWNqaVBwSiP7Sn/iWsI3AoT+KhgbGVe2U5gsDh5r2QE4P9Z4DCN+3FypwblOVmyLWa7OI
aBjUdJ5fFyOoDvOf6jWTsVYGRa8jwoza7If30CYr66m7fU7n2FUGNS/PldiNUpnQI/OXBx392q3K
QQeCSl9yuUGWDK3OorxgFSp1q9mvnFN/7E/bZccJA0i74DsQNdRxuha7jy63pQbvHLY47HPi5Jfd
/e1kycHBSzCjoo0HIccsyrCxeDWw+0QCu1aqdcu1Z0iJw46k1Q7GpTW63Y7SokCbwTcmAxggE+Ar
bX5Puv0icefL2u8N57PkOVnZcVLF8HWjFEKb2w6A5L7S46T0sfpkbhxfw2mFQAKVlS095s7VLUOS
/bwaQ6IMPXfR4s5QN+aEZ7qfxujaMS57LEFYXZLDijKNetp0fl46M6iCRq3jHn2WrodbdFOcaGe6
VeGHcjoJet+reEsDGhCnz4XjZCmf9du9LOOkkpiLkIiGUwhjM1a8+agWF7TFuqBZO1CfcAKfQryS
/pFBS/9NkOJDQ06YFYZEh1DHrnF04XucwgyJpj+gh5Dr2KjSBbzNg1O/8/NnnHyA4s8dK9JAWUG6
mcfV3ONiqiLSHjXq92VOJY+j6qzmoI5XJM9Fe9Q6R1AZpxkADerI8AdL0V/uxc2ja9uEMLCO8ims
dlEORgwN6xe5MfZI72AQjFE0PLdx42KiiuY+1t+3wiLn8t09WlPIM5CS6T0seYtZnS0zhroxuGAg
3q76y23l/V3/GCGFpNR7+pyISJ5V5VhjnjJrVUEmL50BcAaSz/CkTq/mkbcUuath2zKNHxRZ7sVM
FTHUm9EZFLdsv3CqS/CMhK6NZicGBb5HzORnQucSmbVOZUl8C2zvo4dWKpry2u2jYw8wffPLB7EE
R922pTqbEhRREnzEYpbIMzIOuttVW3ReIP+EIAPrH2lbe1LPUwrJRGCX5EM1v+Dh0wV53eD5GwQv
584zkWzgfBHz6iX1fzXtHIEkI3zwg/t9v7+qTkN/Z6yltxm9YWhJSyMFk73hR0XT52TW2j03uu9N
LKZkpemHsAMIahvs1+sPQK7d64M047vC1ZKEIdkuAFWtw/kGG90woiWTv12cAaSU0UZrQxaxJ/D9
hhazvL1QTNWTaYg7n6FeaUzkeDUfBaBDsIwB2Hf6ELTTdmMy1tu0vFuD9pAfzNxIOFIfgZY8cZVt
9HhC5459VgMNp1793oOJTBmPwydo/thrd10FQpD1Ta9tau5uXjoF8/nlxuThzwWjpTsKt78bvb1v
eJW14mWWHPqyyqUhwKcd68Dz6e1/gXJ8PRso1Ub2lEmogB84M9inyTOPh2pEeJu3yGMpEw/K16gY
0yhS2mj7P/GZNyRwnsibR3UOyF7mf199oLH7IphTbI/bob3v/Phmfe3THAPysJ6JjuODqAS9h0rD
y6tCVhjA8PFRuLlaUnqTRWyh7UV3wQ+6B/YCSIT8N9bHxmlp690xx6EKnR32tlID+tYNXcuNRvjG
1+vRe2pPdwP70mdEol8cvmka4Guzk8FErPOhvNJNg+mWo4MgX4bmh8q00wIg/8FfKkR42AHpMDUm
Fn2arBW1AcITdeTCKLNuyEICLBy7xaRiRcV0+fn2dENOxGgGb1kN+OGunDrNd6GYF3lur7b4/506
hmmNOPYVdRjF0SSayjUgICOmLfA95dC3Wop3Y7emAxfdG7L+Xztrtqc+H1Y4kDpPSkcses1w3pAt
RMUTo6NXsZrDTixuC4EwSDT0L3FTDXr58B/CPSDeOBOtIvyAyr+tAtafaIygrMC4PTCJxcQM2kaj
2y99VYmQIxyflyEoeaJRkOgbxZZgA0qRFi8HUFlLUCDikZgFHbUTMlYtrJ08BLpVtHrowTXW1f6i
NAQqK2/z5Mdz42xeFLybNh5RHGDGTvWfirb1zemQxyY4SFwWiPKE5NsB23bslErT1YH0gZLoWQPm
QuV/ROc9xU54e0q8LIKcr3+o/iKDdxHVX+MfZBe49reFP9umUJYzleTeIIeG0FDUfw/i+2sFlEwV
UZkENasH4uHKIt3KOI6icgKDhx94kQJxvwLg4Gt5K5XJ/Hppg7omZfZ22MqUf/8I/AxaT0e3a4HW
ZOeocVqSpajZ6F/B0UTjopGLXJUd6/x5jK9CfrUUa30Vu92SqXXbBr5dvl/5Wam6XxwZxugiHZ2g
grmTVorYE4bYBAwTmsYl4tAu7mkeyh5AgkR6f7A3uwrSK8aRrphVWuKZJmlMU109ypMqzeyUznfD
T1IWmcs47NCERCj6UyN2cs6LYDoXP6Umj+pcVPCG69RHAcW0U7uHxlrnBjUtbu+x/ztAG6pWoQly
Yw1G706vj6Pm81m3eiR3Kz8XO8Rmj8SNiZp48VPjRaTOYTtXa89/EoizQaXn32Ku1DgusRFSoqBT
jGgjsUijBt9tVhRcGW9f9qt5uQOzWrSN2venR28qTjbDTdPbWOJKxXxv2PbeuY73HMWLAjgZEtpT
yB+qMt9xfUd/l62vf4+NPT8+z6JY3CED3IebwsCrnXjPZyOV3Z66YzhXqGisvO6j6Rg1NZQ0B3zr
HWkvQ6ZHhR8X6EDcI79S28gJgqOasN6xfwB5sm4s+4yXsZ9TLibNXb/PjLkc4yL9O5FvuqPq0LyG
zAtwxf1r/SeJx6PXwuVuROIbx1qYP5grCsOdS86keUlRPQHPmc6KCovgJWZ/mivwBXwgWmbpgLXT
n+vCyzI9cePeewLX79ud+qNEVGuXnFghVlYoGYNueeDx4QpZPCjPR/Oh5motUIEl2xPXNYxK8TAC
FJIL68KpbaRcsz4ACoWreK0RwJ0//tI7SbOO4M69b7j3ljAQ6KsED6D74VXG0g8tHxQEYyhdMPRz
XoUEIPJorYEXklaj0v4bH1oT7NAgZMOKjgkSkgMbZZyu3pwYr6rHXJnQOX1FUuiNMMikXm5c7dBg
R+5iHWxIvY/xxlFobtpxArBTBknLqbrXnRXScoxotKSz1G2w7rHzM+c0r48Ms+awcCOM6bSVgGkS
h9Ws7gKiw2RS8xQ9UDnig+rEAnlTXO5LmeG59deJJIzrUDlI3HBPdBJFbZ+MKwYLbYDECOs+xCoH
5SJLP4f+vnYpo3DsbT911MfSaJk2g0xvkqsPjbtOpZd2+wcSt46ZR0/mGG2TSDEyvVIO8rHPy+lj
X98UTrwu0YICaOvaeNZ+gF2iHUaZa3eSVECLL43ZA2viMMnt8l6MW0XO8soBGRaywJK30cNm2S7p
qRJZjh/7BM7DPa3QZLAHHcFH53bbXaWipCicii/VF7nQBDo39nY33TWABTzH7UtS7hfprBFX60La
ydihjG0Yk9rRSvOkZf4/KPOgECnjJR0IctWuwSz8Ud+ZkabOLCYS6+sOwKbBge3QGeuVoYpuMVzs
jGQTIHMMsXJwLSuLQngZEv4s4R6WGeHTIZOMaedE2P/D1KDx857iddulfN9f9T6058vKTl1G/L7/
yDWuYdg1eoNDqUZLLME35FP/tIneyxurb913J/UFa24Y6YjlvPiKbseijolDGCqzs4m1TNgAfZVq
MrD3nz72NeAf8y06pbyLdYr7+X6obr0Qbi5v7mdw9MOxdR90pc7owPURYtelT9Q1zXuVah3fvQKT
AUKQ3o7VdboHQCC2h6dnV0W8idyvmvVSQ2d4q6ngQ9iOidulM4umwiRQcAKz0Z9PEEPLsNufQ27s
MfebrfyxSamHZm8/rrqf0Hddpsv8A5sk375C43HZPatNTq5TPuPZlQdW5Tb5wy6K7RuHi13EmVlr
XvTtiBJbjlIEILOccWf23WmCHUYnMY5Iu6PVH1TT2kpMV9hEyOj67kVnegJpnekaxGcMAkN9w5Ku
Vl1T08Eg4x6RRmT518fUMujliFYYY2VPIvZyoqGMypFcJAx0uOuSamHfKqXRzP32Dgd0OxZQmXMg
hj9NcVfb7wZgZbsMtJqnm6vadf8SfSc374HA7GEDMO8T+NMofWmuZ+OA5zV2ss6EhEVG+kPMj6GX
F8cNtmW9ZCjXDB2Nh1tjFaYjXgkGFJqqbIjwXnBnbwVH+4DmS2Vc5hoLrDCzfy5xUpFc/NA7UriZ
ezG+IhMgCxVF0V6OkDeiOA1s4TFBUcebQ4dxWSW02m3IC4zf/82VxMjQfqfizs1QjmVLpL1MWSuF
25f+uFQkuR0LE5bsaVx3QFirjKoyFZaxkpcsAMHwdsJNkuUW6ygzLXWNL3FtrdrqHPXHcBl1xdmY
g2Jc+2MraEuyGellvoK+yS+VqUpTQHuxMdqKD/8GiwkyboyQZ0jINDgi6UBD0VepHsOdvQtBbm57
nHD7JxYw3RkLZXOLqqCYkB00CBIKhzxry3Enr8EYlzgqbOw96P5yIsUNiXdlEPUfABFyKwClHxV7
Y4H5iVW+Nw4Vp6KjChlzDWbK6qfr0X6LW1QP4EzHTO6j9Gh/3NMa69Ouo/asQbNp+s2E0QYl+dl9
k0F7+Bh7lAjzMdG8l7FIQJOyutG5Qof25gramz8kuAEJdvQLtnQzQCnhiqYM2OFMRxWV3zw7EqKY
mAwoMkOwu1QFhbcQY/sQYL7p7n5gUACLa2DTJZh/vd7zskOPk6RNB/JehVQArzTPq+lGdjgpPr7q
POYia26jPgCQF4rJeICWyfVzkQLtHKs0N1G4DMBCWuNDaHVDKba6gfZB164ykPg9rXzO8ZkmNuQT
RXX4nabkQGhkTa2tYr1SYx/IQXF9D9d5S+s9XOV4u7rPa8F3QtDtdek/mxSJRQGGSyYCuK25/G5t
udmYGAVbcv+TdY2kvXX3q1OmIuFT3yJ0WSfHFstSlomwJsjAScPiQbVWQqfxZuEa+iWhIvCpLovv
XlUTUKTfUE5ok0iYNlXUeIljXvykAfi5NVVOD+w7OXCNk6gN6ZlenpGHOC8DqO3uEwAq/ZbL5fpA
kHHh1+kOHbauXxLK3Eru4nL07R1sDkglwKG/sQeMoQjCmqhg+K0opTCTA5HW7wtuvhMxhjP9fEWu
mRWXSQ3y2cZxwb1/guaMUy6N0FSuILoSJGzHLNQcA5+IPXNE9657LHVqi90kU7h/qoXWR0YOd+IO
UQ3Znagom7nbHECvHD22v/XW07WNWwsxtXX/V7AZMf43ruVneTX/iwjqq1ewvoZnW+sXvNdz1TyV
m8kBizmGfQ32yALKQ1Kwu1dtg1VtxGEAT9o6muzyRZWLA24WoCpfr1nyPFNq4lgt8X61PNf4o77R
4Hr7ng6CJSdWNmXnJX03DCaCxv61WxwcQ9Cob418d44K/lGY20ZgP47qEjQKeBkvX57WApmXXXNc
U6ceEgtlwefPx8/NRFeklwHOlOQOwQUF4ZqU5tsYY94nZg29pNCbc7jOxEP/ybpD+pn7kF3tuL8z
+p3W9OvV1kO9WYgaoW+Xk5fpN+br0VOqpMcjHKD11pjjdysfnPlqDtxtvUHpEeNNWsIH0851tsNv
0Ajov4Rlw/mj8W5B7036xmfn5JRSnrTcwDo9bOv9kHX4JXaCh9n2KmeMymrB8FIiTS/3H7/DitTN
qOmbiUWh+ifck+vT/uAA+W5GzuIs/8A/aahMKtZBAb8nuFHY4qPCe2cXl8RbpGp4Jlvugvt7NJT+
XfmWcWGjACKwzhzFPwbI89ApkL4832Hj6HGJqvts1rLjS/diqOpHr5fkxSYBg9mKcKfOt3o1D2cd
8okdaTLPpmi+t5GK9Yc0Rl74+XNv0/b+cJbkX9uiG4qavYLRCycq00l4t1+u0byW0g4teN2nxAdd
zODCLi55jqLCJgRrG//+uMhTaQCwpSlXBj6NYquO31G10BsbQF1ppGTDlrOkWUHQ5EvMWRfGwC5Q
Q+QkgZ/o+uIgy/z7QBh+S2hIRhjUY9k3OuWq0HnM6aj3YhRvUL53tTZOKhzge4A7oCnr4gxYcGwb
WxKzYPQJjfUw1Ah7iZDxY5mtTx3OlYpXNTG7Fa6Ik3s5JQgLuqfKLzhNCXpqnqUDr8xbw9Tr/HCM
i/7ERX6JYmJnmeEcx5SuGb5skcrnjmTa00HMMoIFir0AmP3FleIK4yZAEStfkuzXSkNOrc/Ri+E/
B996WsvUXRbSFzrPoJ3xGFLqndMl1ZQlDXV987gQe62T8aZRbzNcnqfIos479qxwMS4emJ46hpBY
odw7MDdIHbeC4dtHAOQlBD0KOzhVXrJ87wNsOke3vMfVK7lDudjOBAApL41V9+HnHzwXa/mF6kdp
eDJ/aB9utX3KqanOphpRqErVg990bIG0qoKS7tMi6HvtvbmttmAQMrHDRa8wy1dkMYd4W9fcUlVK
FEp4RWagoFI6/2QG49uVnIuqdXVXNImyFM6ip5AadC4SD6SyMK8LysADNJSHx1mYO1Emxvi83cwO
1TGpviqpuhT1fgaLkYfJ7NInKpMnTp8BTcAosVTjcNVhBxr16lfwJQWHN6doxr6clj1le50R4PlQ
ERfTvVS+CX4JXIqj/l47XOIcFaRZHmLIR0d1K1qRrIpI+OyUJ9D7o8HBid5DYBI9wr86s/repjTd
tahjP4dT5bUcCkZIRM+X+LZuyAzBlXKSuVUWp0N3rB2HAZ8+7agCdgXH/M5B8a2YPD2TtRu6s6WY
6jvzfEag9CxaRfkJZ36nLf5KxINsUsoCKSTNtCHVXsLC7+S3eqwF4MZW2+PW/h5gfhEPCJZJFiJj
I1QoWk8cBSIcWon9miWj5Ha/rt42XeWc8GT4A5g93AHpbdfvkti8naS0tdYvrv2d0cT1Ei8gUHeZ
FOTM1HrqMJtuTY0U+9VAakhhWLG90G4igu8VVz/jjDUBW4+wjFD07EIa3wppOUut2VqjxgjKoJzw
124JfY8Rb025TLtSs0Tj6zsaLTdN0BspykBDZmq7VANgjJH+Z66BUvEAunYw6I/AmvjJKk+/V8F2
2W3Ib2lpnCQSdyNxEAM9e/40Ok0hr63ZRJSDyeMusQJyKKvzYr3jUi4fPdr3RiUaJNRfw3JSOxuv
9F2u/j9xSi3DpGiIo874wlGpQkg+5I6izaadOBP60UTyrXs9M1+orRxa7+LxLtGCUf5PeXy8ljQB
SYf7eJ/SNyb1y3ldSDf+9ZenSdbQuMPmzE+tHUBD67prAxTLPkwmqyeueLbEd8awoNsM0Tq0WY+m
N4zUDRfJKC2XLK8QRPM7FlqanNXxhYM4k3Fpg9JoCv8JLUGYaZUzR8wTncQaTVdMrr4oxgzOzjCC
lnd5Gm1zRO7OZeiW7T1FUis/CxLUNZc3k8nug8NIhglUMUdQXC+r6+JyH1u4Sy6vLn3+8EdFiJEl
18lZ/fACUis3wlZrCoC/HCjVt8yZJFalAdLpAkGnDC/YQBZkYGgtpDgXxeSArZrWmGLj8ziP6qJq
ZhAgwyxmG4R2uZ5D+FSF0YCLl2MEX/NhoCsd6LAgqN06r4tpCbKxmPpmFxivi847Kae2YvW+4k+T
h6iagXuD8b8UNsQnjGKKv8R4m+bfKMuQpUh4k1JEsKVq4/wJ9vHr53pqZ6ytLVQZjoLqJgzVj2ty
mtdwJ/8q0VZjhxvEl/+o5YM3GiQZPJpA575m/JBELW5Eve9XBaEmWEEgx38CbvOzls50mHOgFlcT
rKinTfLdFsBruH3BjHR5LT28VLtLTpmx43JbcvU5t8ovnovkxE4GkBqX8JnhpTxgk1W3Ib907A9F
6RwCS0cXrd5cvmIlQfagSURBkiPlninozX3GlDHV9Z6mJPvKGFalp1P14tkgspUBU30tyA3eEU/+
P4dUkK8KgDspyTo4X1MWS97AVqwTq47vxFMl/EAhAI5VB6wqYRLT468AAgHCCFRZSHEcB4lkv+Lq
A9XVr6RFKYFOflu1ME4F1LOhHHnitW2yoamFDpmDOohRWLpTg10Ml6mfx8V7ZcwgMexzvOMdkI5R
T1o6NaHGGIvJ2fG5MbqZBz7kyDoH31odKvRMRB0F4SDOEe2MX30pu3mARAbvTWHjQa3TI2fmGTLE
+6Zp9PIepELo0AEBtQLdUDGkaAfTk0zXWAhNpayS7HAf0RxqezeGGjX/hzZ2+Lpe9fM/TKa0FihP
DdjE6S1xEjBVF7OjL87ybNi+eZwnrJ2cBA6tu1ds+xYnG85uHeM/CpxPdZHsaWqc+usRWGdoF918
JftuQwJrdsecu+n7tPkncRsgH4bOW66TLL/uHVtOBQedqnbfVacRleNxsCMU7Y854lspC5rVq7l3
Z9x0+zScRKaA+ewEcMPxVo1jtdDzW5H/01pDgtpDO1KGcZItLhaTyBdAMRcZ4CG15IibF4Fp4Hfu
A8OldNxSwoJeJwtrpnJip1TL95tvPkyl2+EqwWRyrPh8y7nFbd+ZUX0ZWq9i0EZagvzqtGrgPvfA
omY78PBbPH151GtM2cPjTwRjuy5Wk2p0fcpmHqYciOEELIna4dipnVScOEjToj5yi7k17BwRe/o9
InFQyp2fYKj0HDZvZ04I9VVspBPCLH1pnjlbfCsBd/fYP9aRa4/yYwruODzfJDW4S7WTS8p/+fYA
ytwOODNko3MdfMX3cZA0PYToRCgvuiMrZY/Ot4+XgA+ZR2yh4pSBiZju82AcN0HeJxn8PjLhJv4u
JYRtstZYIwYMyxQNBMLdX506dqyIO1EaTLLILPHiq+TQzwyXdvSuaAjupHIENNqVgvyj9nI1QyVJ
GpEjBNvQ5ZQkbdb6GVcnSfsfHE7wtkaRh834Tqd50MU2c4PBTtpBTNFUYArsZEdevRL8w+OjZj+K
5zBHjoLYZaaFCw7s2mmlCG+6AxqRoh/5kZvFY80l6Skhm6JEFEmQ/BD7N4pW8kyYpgqcdOXH1kol
DcSUFoz0KRVUfXkkwv7Eig9mEQqWt2wczogvs8jQZ3AnMzUyiSCuP8BlxRBkTv9MakduNju6dhEr
0VNuFleMxArqXbIi4ntxHBF1ZmluNXqWdM/PoZ4bd1WBfaGRIHFBUI4d07iqojag9oK9KKL8a9xa
vO3LK/IhphxkNSMIRHgFQLQ1V2qZA8P8Vmfppx3J/mawQvMx7Tm5Fsq44OZHpil/2UJb6zFMAGCE
C2JQibyqh1t7nu/1SnYMXnfLFcRUAKNWVO4Q0kHi1IOGHzXt3jSBPOVfe1A27nfX072XSeaMFgwi
Tgk9cDKMci+61hS9oQuKmQOuQBkG5EEz4ytxooc2Gql/vN92pPuzMZ19tL7L2yxZqcbyLckEGQKa
NYXRvDmqbC8ZGY/QH3hliDkg0B1LJ+C/iIW3PbAPAxzEX1PWeVIDynk+yIGv8xpVemZ1taVhHGGq
o7ZTeMjZqgK9mHU4FM+zQhBSm30BMUvTC2+q9vTtoppaz9KugoTz8mU2akwYibpIARFKZTlC7u9v
dWT/FFzgaETjzdr77pQQ7+25jjC4Tx0SxEM1JF9CyGs4oYEXWoPfGRJ9+gT6wHiLEoOhaZ91Z1J0
5KJJooo1W+Mo9MYsvr9EbD9n6kECboP4G105JDSHMgjnx3vZeAUfhXqcClV51smCeXRTJqtAHvyO
3Mga216cm1HiPvWPKtGK7CzwDVe2wMAUW+kXs3z0UCycFx9IhTpo1bd0AJ5wnSPEkGR5rULrGywk
I6Scf8Nk4/Nq9xGCnAC2OSog/OJkG0htSvGAQ0hj8yySpGRf5sKJEbJE9dWb9gsLAVX8aw1SU86q
Wtz9TV2IS41iUW5hD6XXgyVaUFAtRV3KfwCSg04muU6yT3sWUE/dTbqTel654BWAigvMzpN0AkGO
TjtSesmyZ5zRAISOYvZdoJqO01ds9iMpj0Mj04L7Kg4wn4Z9mrr24hk/tROYvFyRWN57pvqZSgTc
UjTMD5G6xvTdoFWOvgVDEqwejqNKlzMHDTmqBz3VP22jQbo8H6jNhB9q0ziQLPYWVBbQVmYCKmuA
aQraluEAB4ECE8LA3YJfVwkfWt0yrTwg8a8tmG4urF9/G8kPsLcoL/8BoPCAGrY/x8wFfVGEKmcI
nUtfQuc2b66dzbjkx5jh+hKKfOXEORgw1IIgX5jNV8OfI8dMR9x96D6lch3iUHxmeybxnA1okGHP
q1T1TfqQCojr3NU3es1ZgNlMp3e0cfvrUgpMhWsJ68YXQtPTw6pNaFMlg3Z2d95Jj/nmXWQVDOFj
+RDxw7hN4FkTffPRWaYfQ/8pE8E7vErBM50p7PCjm8rzf8UqhkSdlDE2FP1VVFSd/eYKL2PBc3jb
FsvpP/48oEtZ3BBUFAAjc2HliwsluiyIms4VORbsH7NrCh6FIbkL00pcqv/EZcpdKQ1j2nr2xco4
YGm5pc94OU8EEcwC1onVX/a2w8tCSuiCT4+bRx0OaZKcMdRILKnuEo1zGgPXtqWnWtyJyUmVBI39
ofjQUp5MhwSRObeK6heKVuK9wy1QOuvwj/vgXHag8NK219xnS/VrG+Lx/XoX0vARtS0PJ1Ig6Fcp
9Y6EljQ+cl+yMtp4nIZtZAwYTUzN1XiyEG9ykP1J1EXRHSdZguiDXAVqsLj02VLVJN5XsCHP2B8o
2Q3QZ20o4CfiDU5lM9iKaHuf2BwYxvfyiiXAY0LXTAvSQkPLA7YtKSDDTTW8yuhpuev1Do+70JSk
EKHdqxoMZqhMobky8JVL2JPR7Dvh2+VNJKMt0vwmerHIps3/cykvc1jJmx300OWWSOe5JdMEV3yo
JzD2csrpWup6/WPCVEL3edSZk3l9DJd/d0wjtIlEyKoYGbJ2ycwEEybzPRzP9Zn6cVv0XHmXo4nN
vno+vm1bG4anDelhSXkE4PcjBLFkyg8BIDAGZNbZ3tq8T6QbIXmGPQgVNXfVQzbfrnIBDZ1ZlNlz
Qo9slHryLGCW2yLcDa6oc+80Flvfrz9p8ty0k9fbl9XeA2cb8wRS13RtTz/dFl7DGkscxZe8o4KP
I62ifFZmkRVQXj4Glyi0qIL1I+IsCZJ/e+oCm5aDgOJCWKOFfnuLu9oFClqSJuTodqyxqFb3hoVm
1qHkhU1E9TIUNNPbJHTemZVAWFBHHtWrpM3KRrYlFeVdZ0bj5Di7b8qoNXssn+iZyHlG2YFyGcG4
FjJRm7ExN9XnQG5yZ+Ntmtkj8Mt+TCkfRHSXX63+JT7PsuhsRujY4ZRshhGAfbiAdpeUjm+mVZh6
RVULknG6A8xOs1Dk4kaJDrdMWnbS4tMxKlof45zxNsx4uZL8fLGIcWaSHvTnP+mCQy8MBs5taxBH
LaL/VSEFki/tpwMNZ1n1Lu7OyoWtgFatBKuRL6Mk9E97BRAnfPX7pOIRPPATc2NBU1w7Gs9sabGI
KlDLpdTFpPw3h8BqaibKKKNAMcOOtJue6q4oINA9ZnDteRacQdhSiTAleVsMlIP4fIJovdAdPH7X
UDhGRlY2XxzuciTO0ABUAY5D8CIsdUKUt8S9z7fDlXBOc2MfBtpm+NbBY/gjNOtLBoFs5tQ674A2
q1AYz2zlfKHV2Il7K8U+pNR0xmq1wPfXukiYotS6kLy9s5jDLG4jH0vD/Y5SlPeMHE8jRFdsKi0d
0kHDYpFZHLlIovFALC5DPgWMZzkw605LTZJI0SNYiinBuls/5MSX/jliLVW3+mis9tjlOSV7b6Ba
Q5eyZTNcUM3loZ+Fl9AWB/nh07w66xV8u3GXqm/qtLJcWUFkO4cfqVwnPPI1TRNWYMTfvvXTw8To
iL/MQ9Gcz3r9ZrZ45x7Sa0G+XY422V+xJ0B15rhZK/4zRw1qS0FlUYlkLthJSllCMNvJ1IhIV3Dw
eh0LWefK3G5AaEDETh9Mu1vNaNYtdmRmHvCNK22p4XBD3Rx8utr4ZwTR65w540ZYNcXUkv+YEOd1
y3nA2HCHoH4BQAThgbkTXLQuMif0FY3w329RL6/mh0pJSmjmPlc3FnjWVoxrmSmrPtZRO5PPD3mw
DP7dzBQrFlN5sCDWqjIEVnTzIeAcljf5v3exb2TUNxuDcUW5ISwIgtjw6N/xme8boA1svTbApVnu
zk1y4RgRukT3taM32ft2DGlYTipL9KHuYJ6Qhjk/tcWxSWPL0JWlWyTPWvIkgZykSdZS6Ppg+Onr
AaC3UttO+TcMv0jXx9NPxGAWt/Mjp4HQPFvKzfn4lC0H2HLBtSNlY5HngfKfD2sGV8PnCxcqD1xO
s/S3DLgHLQMZXcfo+oheHEGbIz9dKeH67lIgBas1hC7BqlA7EWZX8AANUhOYm3dB5bRof388DFjZ
d8TNrE6iZFN161Esl3QmirV22rk4R3PC5C7FFR3f8flhgBw4Bp49sLVNOEBMmuJO+0y4GE9nhewq
sDfJhec5bg9yIjD42+LgDe7AmNVTJDY2dqydA4WQb3/vh4e5+eamDHxoTLV9Et15y/e2uU44RZMe
tczhkPJ6ivPSEjpwUfk4Vmfn25nuDxGfU+mRjdx+9ANutCX4Fc9tia2BwfeSXUhwf86840ZyP726
kbisVu5mjaaFqDE6y5J/IiFAr5mGytn+Am5hY6M2PymgGJF0KfNdXFz0zTxBfeqhPS7qi0OlZsen
p4mMuEDTL1JunRxEfSBYx2jEZpQ4ORk8Nj3yOttb6ecWVDNnwicHXLhOyubq1smsOIB5oWDrpps5
TpXSX0Lnuu4oVfXuWTDjt/ky4dQ13WK55l/NWMDfvYDWu2t7MkBBNs4qkPGMiiWDz23CL8j1I3h3
haKaTQH+1J0VzDPkPcLpyCwt4pOGTJAnv1egVZb2qfzPReqn9RBb5jl3XYvYwnZaEU5VHsLwz+xt
Y2Gm3qs5rhO4XcSaO4xdtG2O6w4XblHh0lOxXbjBbt7WUFxxYIpkejMyvyp8/XL/FQsUDFb1M+Iu
iPgM04QK2ZLbHPajm7tShweSNsYdkyp9JTLX6ATBITCOBMZCTJku+xCoBrp1cCLR/Q2ICp6MX4zR
HIHeKpMNna3d5/NUDopjKZMvA8C5dv1Lo9QcJF3Z2VCmD1GKfPeBLukFe9cqG8SZAjnPkYj98WTr
Nek+B8lU03csYPLlOOoEI0lIMisgqIyna6NVgFvJ8ZJxyf30Qn++eI2GyvyCRDt6CODYNn1DeeK0
lPCv1sAE27rhYTWmIYmTLskcS0rdMI+9IEa9uAODkNeJtdYN3tASLFCog/VyujAcAr5iO1jHKGHw
4rFDT2AOfr7klGnneTMy6CHZynrfdkE+r4t3Acj1TnoydpfJ3/V6BBGkflsgIHGmnW/r8TyU1mCe
8P2rZaofxPcZaFhobFeMH318EZ7Jz99iW9NHHLzxpY24EI0vy9Zza2v0UAqU+D6faZqkqyLsOp7S
x/46/IrirQqqX44H0I3OGqrC6zAC8t9XWWXU7kPnCwXzXjDipD+TqBRcJxSBFI1LCyOUwoUIFTMc
28A57eyIzD4yxBJksQdbajBSmSAKCmqTtlRi9Ug+YsOouhgffhkAGEBaZF3kDlr3lUPZf82ljNBJ
M9xq/BOtPw99/3AOXoAVlIDhcJvi3utUv8la3SekYXLI0yYKsbCC9wTPz+A8T3aiNFfM7lhKpCa1
rn1Nez5BA1GgJOhec146pFt4dRWmWi71mtiV3x4LPDQQuwe1Wfnzp/lh2ib7+7JWjUbX8i+PM182
DoI070Nu9T6lOazOqlTVgK9yZSWr7tTvjPJDhv1banMgatawkBPF9CLvpEGhe3FN8S6JMnCG5p5x
Ety6N+qaLsTPSFPiD9nh6YPQAfkRSv4sPoZp8OSnVnhvRGTSACitxeoPlEACW2XfLmnFkbKfy19b
to9fIZXV/+G5m70Ljz6qCQslsDU6PnHLVKvthmdkiTvgeFCNRTMZMTCfBxoLqH2KpjT1KAoFDvuo
cVCVFwsaTZDSqa8JkS+9iO2rWUmU1LHkQd6SdIeThmvfwVl/RcJ1xIozVAm+L2yKL8p6Whj+yhJ5
f/dw83GeBF7uiBGptT6DS0lB1bGMQbSJWWjadMKyCg/Hbny5Dlj7ysZb7/0cxI9/GSE3+zjKBtSf
12FfYpsdA49WKk0fLwvhCDVB+rgI6tr+y9mY9qJytDYLgAMCO9PQkszL0z7BP/FQIh+2QiD+xgc7
cVcC3jqdU/DfdIuPuVU15K+E81zLBcn0brvobibRkEi1wfw9t3zLbbjOE71ls1j7UKKBqJT8pwWu
l1gq/XMhVC+ixQeXY35mzxzPYHkETKHNNDxF+9cYRAcOju09czayUZrCL1uo3HBa0H/wT+yDA3O6
rmeIWk7lKuxsN17SP/E3AKW0k438FZVC9IBhGOlCaUaG74mJPU9IzjDVyALrk7w1kFqycxGuhK7D
ev7TuTjHaSCPNfB+qffkXQgOgkV0lOA8PzFd7u869sBH10s3ZLiyQOyDSW8svt1TccV8rDF5Tw0n
GjYkur0cYcDNht6I+5iS5tZGDWN5BF//v9z51LB45Zjlnh5DqKbQTi2/DZIQNsuFjNQQM676I6fu
Xm/wYhOMewLTP0OWeBRF9SwpKOYU3SiB7Ot/8ozQvJD30ykTtH1J0cAK+N6DmaOcoroLg/FVl2Pv
H9FkVfbP59JHp3BqSmsITYZ2hOcpWMuLFwBLtbVSn2jNThNTWoE1/qyty+09HOEVttASqi1l+73I
wxsgsB33/WrNDrfyaKzHOHwwKORD0g5FXDoT/3xZ4T2qo3cOcm8MifnUPPTlAdp6pQ6N4Ey314nx
W9mOO0rbf+Cc2s7pmxMPWHOmmSXbn146N28o8kR9yFDLYDPiCTU5ygw4clASbJ0Sa8c0nF1aIFVr
GTNIkEiEgglBNmfGuz0KgTwI1+8zEookWEU0brUKqi9E7IIxthOr/4I9OYHSJE3TNbPSyFjeEF0P
W+3gOKAifPA5mLSa2IhG0BiGIiMP/Uk52vgv7hC21f0EFbbCuhwBJoFamsTZY4Gs22IHqeHZFbs+
AvAOvhHXaziZzW7nt6eTRMf3ljnwnWCmaoC88rFCgul6YLUChKwYbJ3pBksZeiWN8NJukp4+lYoN
hRhpcthF1mLV1s7nGd/z03qGg0qOUVYC96hX/1kw440xea6W2jT98Hggd3I1pvCaNPFR1cJZ6MqR
Wov59R8Sd3S231wTXPHwpLmF2DcEMXSNkFmVZsACGwfDEX+sj5CeOgmLgd1t17+Pbwri59dikZFR
6+VzD7BInsyyHUlG7LCjHV1clz3WbZ4JQ9ITMrbF5HYSxBC/qnWsCc52YC4RGagD2mPOGTIBcwAm
rpkLxV6+Rh86sXTmR5bYzcou5FVPsz65yzSlY5EuVp2C8/wqvfpGzRxaxy5vk9ZFAInuST2V7ntO
Waa9hZ7yyP6lTYk+jVdkaFr5p1ZF/pfePSB5x3QkinINJHESgXa/drM2uhVQSu9y/bjvZQwoyi3p
A6ZUPbAs+jDUBBMVZK6diXi9Atg9NlaeX3957l+uAdh2CsVo03uAkL/aeYEF5PId+KJRwwX9fucJ
y9aMIz8SEZJ/awBx7TRqh48Lu5e413+OqvU0ivQaXiQSap385pL6Ua3A7H4LbIUO46j82sGm+Fuo
Dub4U+lbkbZXalHvIY+I0Gkr30kmw/Nz52YFQsGt6Xa7KfbZHWeojmnFVWu6Jz+nVit9njdC4zzs
48/0puV0rw26jJkqxZ1KxFrfNZHlFdlsFx2dA0CrNxSGKCRnrhwe7CeZwC22SmDMsTfkN4fMAfaU
TgAjxF12ZwAsibMJjKwBxBcaGP75oULLJEHdN54NmE22tSpWlhTb2qhTY3yXKU/t94dD9c5GEcez
7JN+aLn+AmxJfS3PQMNIojzdtzl3tlFiMupkVEtcEi47a+Heo+xTR1oWB9fcxzyaN0Mzekv+Fwj3
d7blZ60zkt3bkig/0Nxpe2k8PGxab8t7OcDVJZ47AmAC7NYEPXCYLsqqdjaSeKqAktoXDSQWsHbl
bJOAWi7879ne3ir8oDodSvUC+3m1mVlTGxxfb/FfpXDWMpEmMyT6Ff9JO9vlFZVzgk1ANiqA09gQ
vzSKKLjsdjInHaIWgMvw43CQP6RH4snjueFpfD6NAOXN81LZR5sbXi5835PzwqG4+k6iq4qhNKO/
obzDGZI6/cCo7qP28RA1WyT32UinF+BkaETjVRebpt39umLLYqsPf+a6aL43p4LK2JwHIeXuNG1P
Iu2BxeNXXzU/akS90zOo7rP4j0bP8dcABOZ0s62SFCuYZwAsr9JdmFu1J+/ERdKScNyJHwN5H3UP
ItDONWc4wli3+logKsaV5VcZptjQez0zf+0IzjKayipWVTS/3dx0kCzAQv4+qNYtK08dCNVE14+k
Z0t4c7FDJdzaaiIkgoSTSXEy2GOguisHL/Tm1KmE8ENx0QIfdcYXrW9qM8DgTfl7qNX9Idpsl+JX
oPoVtYUuoIjQ5bbNonxx0LkZk7fVRW7sqKP2Ko3yNxCG6wkcay0E3Cgg0D0jfBdkihZlPTZdsbyU
x0O8TyQ9sLN49F7axVCMblxCnru++YT2xzudtGRaRR1md76rjlcRqNGbVd3EGQPgRjw0Gr3si5YN
+R1oTIe4+gU4tT41WcF2nL/uSPj7iPgKhIpJINEnqb0/Au8AsmLSyZUimG9BmGbXW/eoRRY6P34T
A0p4jOkQwfWYK/UT3h0TDZNCh/w4C9MB2HWqNBZvW4pl3n7QMhKHpD+MKT0V6dVgpASuWmTTdpA9
9sWNlhmbEptIyI6Vp7KDNR74GpipEHxhOxR2J6zaw9jREbOwTgvPDMS6t6INj7wsIpI+QJVNLwux
Ecufzwl9TVmul2V5NKxvrtmGc/qu9UCslvgnmxGJorJDuRcbMnxigwwRWgs98qyee8JQFJVdvnSp
C4NhJ+9oPpUjtSXQIqGov7RxASNQnigTOS3A5R1E6edLG9MKzNs4VWfKUg0wT0w9HBb+oPq6vXZk
FzJkfQSMWOiUYEHpo28p+zjE2ndspAbhprcZOTNmbO+02FU6+/ATWiZvD6XihQfUIZ3Ng+YrjmDD
WqkJwM/VvHzTu8Bxd+AqDuYxWd9aTfffOFv6N9qKrEv4ydy0AYM6eqH3zKMBDYg512vw5oN4v3Ny
1nfxir7qRKQCe/mp3pguWPAO/S27q26Zq2R6BGIYbYVzk8sMGanZw/LjzsBdRAAGObTyguuhX3V2
0z7UMSXmv/PpW78kNH4GGUCbMgCzesP8Tq52vbzZUbrOxz1HpxqOz61dFkx0l37VAME66NSr5dPU
iDGhNRMalwGpizUevkkCvBAiVnCPzC5RMSY4LMdS0E5Ic+bVmkg76BIBz9XSlLzR9fUMSxCse4y5
dK2X9sw5B8ABcTbcFLdEn/gV3DThshyLbrgduiIZ0v2/T90G1JELJvKhl+fWg9FI9xtydZ1ocMGS
OYtVgGJxWNS+LRo3XTionEJQIl6RJsjSuy9N2w3nZJnX74otjzR0epHtIu8ONAdN606ZyrCSTUud
nZMvXyj8uADlpshS0qH6fbkNGonyXdzCQ/Atx7IUtcbwSURMHRDb2SGY1YvNPCdebHRTsh1QaGii
ljfF/BfZFvgO5S6j+J8J7bJ6NJdOceCwClGrAWa92rJ2+4zo0TdqcSjG9nar6lArNht4z/D8/yq1
GPHv8lCWZBchFY0aSxGeJDhiY4mbi9XMGF+E8L4Zs9mefAr1eH1deSFoJOJ05gBSIsUW1/C/plWt
vyXcV7PldqjXx+4UvK1T05L+LmOBZZ5IyYY5CwQQ9XBqZbba7wLTjW/eJGWmGWOohxLi0Pa9YkCj
QlgWR64piixIWj7NgrWAofl350vKiK9tQgbwHIOljerOVkgl5XNhmDrdO05EjAePjsl76EDfwYn/
/N+sL4oN1icU0uaquArtiVpV2kU7NrwG+gDgseIF26NjTE6FUVAwGIMUUcjiq2fqG3RN1XlAKQPf
CEF5EBPZtzP0uGf/KeUNq0vTEwEeHl1hFmBN81fdeC0N8BkDUcgV6DsXNpGo7Kmz7ijtu2yL5rBH
WqFKxVl5z48kZhnZkVCvfQoxa+CCs0dKyxAdq+j3wwFKn9PLyHuBZsYVI/5IuQDmg+UmQhMMxm8E
HByh3E6p+KfVQKgSGL0+5o4Dgaj0b0Ds5MRgoYWG1hn3VV/ieBM6d51b452FmNcH4YiyHqMot9hN
n8WTye++gLmnc4UkyoXGkUCBFtuAPjTrcIwK9Nbieq1l1QRsejnnKT4R0IUTkXTRU38/6eTnKDLe
ToMAepYlCfUiT2867Cj3OIjE8p/UZP5J0YFd9ykOPs7VLG4BieC4L8qFxN2fYJZBDR9INvNt0UnC
H+xivI/y3CXu3N9EVV381tlMDN64GezP87ehplFUmWOvrxBcNnrct89WdDDcB8kuEv3BoIcOVRr4
m3Wg9OGN2Po0Usk1nupVLeXqnmXi2+/jynDT/Jhz4SSZVED4rkzp5ss0qeWITzFwu2asYLOgnwBP
gHEx2MnT3UdctFtGrLFuPFYC8CqZPUfpU6nbwhwwE5k83BqH5f8dfurU6kUDcXYKEwYt9sg+Baku
PRrwDj24Lu3yFoRHCQ6QFgPRHL9eRmNnvEGdQkkhp79lBjGe6nsf62V84ZH1ktcazHvTX3n5+38q
aKUqJWCHOPXFGq3uCbjUd50xFbmKF9iSPTo4dDZif8Ksk6bn/h7nJEzTQ3cMoqKUNbfHJeLaEM1r
xJ9O071g8ghdUbY3RmvgWQi/QDU57LnJfmV1WdD7Q5m9ENPpnUrZPbKH88ZMoTRZbxlXdY7EWtgB
rIGUJ10tfx+P2DsQZ/deXfc40jrCE3tR8+TJFLEc5Ny2UbPjfCVmi2TMNbEX1XBrJ992Q2Jsq3L4
61FPF5sNKSiwDurmnO2zCrDz237U8VT+14RIz5fiT+zcc0nJBlOsgwDZyzLQRR8vQhbNaoORcKID
KhNySyXJA8ItZA4MdHYKzO7PkoAyL9PiBTQpZ5/c8u9mN0P0g1s0kAQX7fRgdJhnqCKCV+bfgF84
nkLHrX++mE1gcMkdPTtLO3hR5NrGVeOGrrq5FkAiVbG094WghI2tCqcNLL2b3/fmUSdIsmGJ/bmi
nvEUM2o+CCrNV+tW22VStU0pG2tiWh8aR+5UfLJE8Tg9T/5qrPhgsSZ9bjReAHercDBwAgDXHtVa
SzuUWI+d7ed8YUcUtee5g/W9dypSdvaJe4Bd1NmouW9GqIiEnmkSej0PyD7eRmsF3b/w1tBpla7A
lmSd4izTOwKn+Tx95QmDJoTpJbNqgv/S98Nb8UkZ3zoUPr+Woh7D9J6B+IJGqeFTug+qE6JiGoon
OAfdeRw7Fx4HIZDsfyeubMKAbu05o0EeiNSw9BuNlW2/omEDeHyYod5oqmvA9z2rBEKHPt6UQAAl
g/TpFmPwLDTmL5op9FYb2aQPirvO0SIB/H5RfMsIzl6xtVgJwu4WxaAIHfrd/nI1h+WCF34gDYYd
KOMxt+LVS21CF0dzoOyaX5quLLFuPkH2jpi2kkySRcK++h8MaHcZjklQsscGL5GsWsOJ9ObTM1h8
yQbVLMtgMiKMxPRXkZ3PFvgS/g+1D44a7p2FvaoKmHiBoWap5CsslNi2UEfkIw+r03eSGJpDiMSV
vw1/wRTBTE17bZkqEySoily41MFZJA8ahUhht0X86KhPG+RuMUZvDQQhhBC1mEpw3nrxkgAFp1/9
VaYfoMOrJ1QBWtKbfuvXo8Hfi0pMDeGXl6H4qmUaWXTBdH9sM6aMzstCNDreqkYLpTCiGUGN6oRZ
wqzJwEuZ7dY0r6VLLUhRUovvm/iTUYd/w8ibYDAVdbbZklYbg4+5iEnIWGo0LkUTbILChr/1nD0h
iVH3wqsKlHks2r2kL7nK1dYlw/Pp9ckTTXP+0GqWGNP1fVeqF8siT81cGRdfHdmiNXoTW825vtpT
txTnO/XBLX1A18s3RKE4woMaBNZbFNp9s324qgd4lYPXpYhhA+mQFW2xxonzl+X5f+vjXoESz0iX
Ow6i/KfdL0/3+ygrsB6wHPY0cMbNV9/XnBp9/vLy5x4keZ7r9wrgcUl3tSv+uzg/9AdodL/Ae2pE
lncikzJAb4QPkbAXhojpoldE6B246VcLgDWO9Egt8RBASbqZRK9DVfd4YB3bf+Lmg8JzJobwwXv4
8WXiPwouprWc2JVf2t5QVKvO+d6LaN57s8BSUw+L9YbOw0iTC0ilTsr1sznSNdMgJBSDyZeaJaUp
beKy9E9F4YtIV6IRZgZOoJGw/QDUThsIFtMcobYhbTY80v+vx9qITsG+rFpIaY3eCC6MLkVNUXdv
fpsexVM+5Z9O9XKJMm+PCn3B/NNcoB+KmfQ2iMeofUafGGnKBKHFsh0u4M9Es3zlY54wYTrXClRO
OKKmatdR085oz3stJliAVEdqy3GsAGSYpvV79RIrWUNnDo4/VuIZYq938P1oWiHYOGBzzsbouy4R
II2pTCqObLBwty/Gtsnf8VhguDZaDxzhOmKw2hqnT9LCSfN81KLCxC+k3V8DGS80R3tWanIATq9s
JAsKspr6TIUOmoAdStWiWT59L6bjrqCMTpZvwc7q4o8e6P95ZEi20J/dHNGCY/7uNOSbkpxmECta
ancxWf3+nQ6sNb6wV2vsj+7pYHl7scrZSnvZ4sNLJmg7YpccFKZCqyHW0uHInimCWsxHZC8aDSMT
yG8sA5vRaC95mus7wnwexVPGo5mEX/91O491JoMlJ1XPUml7kC7FD25MPIYUeICCH9yRVJYcUYQy
61HJzRuEcC1ggBOTkGNYvOOMekfoWjBHVdR9hkzizWPgPh8oD/G70CkNLFlPnetWi0nUmJ4BtKh0
ZDuskeq5C0T8YoiQg7eKTECUoHU+oz/2OzAC/Hbg56rUSo2uxHpsuK1A22JRujrXuW1hyfYS9xkf
LSFvAaoWudwb5PIC4Xu24fck46g/WaWp8ZPiQOHoha+bsphjf86MpOFv6jj0FgqtGHULgmuvB9zC
gFvFnTRzOyzUKKZlHQMbpfXAhhT/H0JghMYml/GIoCBQZPHyCuNuxaWQ0Bxzc/tYVSGeN7ogoYa2
UNLqK3bKcOBzoOegiH4407uW89Jjy8oG9yRX8khqkViO/q+cvV9Oo0nnrFVpQPfulueeQpCLSe6T
qFdFlR+jSLyfTRY8a0Oe0dQz2hAREhj588ZM2+nbkux1LQOfNRS57Av0S9/gbYjZp2uXWERAkjHu
2I7furT4VOwTFknphKE/AD0yz1RH4q05sqqGNeVxQH56bbBUeidsEhE0In1bCTJheQca+f91bLPR
yJ4cHjKvGKd9FUgtcCL+2qrrISSgjlz0u5Hd+Fd9dPcZiEjFvsSjFFXwDPyjqajkw9eXMVa4e5WS
6hx8ni61yUgKuKldHcF+EGdERCwKizSWispWMZO7uzewkyVrKRcxGeXWblPFRQViOuHEBkYUAls6
fL9fw4TvvOconTYRbFctyVrIecIjrG9i/qpaLkcNWkM/U3X97f05SifJw4VkYLyH0skfDunL/8tj
W+6SyzaCHuhT9MoueNSMJryf9rocmWLX9biLN1F3Drd5/SW0vrPcxHH+q98SmT/kbl87y+DCAidX
yTanKNvqgSlXXZNxtO19n4TfhtCmKejxSd8zJwxAymGvoPBkcRatAz4oViuQ/I2Ht7GXKQ8up+3I
ldTSrSRyrnpt3riyDSlKwgASzRjKscjK0W+PzduToizuQA20W65Jd/RRNQWVtd6MmyqMGGfhlMan
h5LFwqaJe/7PyfKwMRC16MjVj04dKq4wcAfaGdwn569DIOBu7EKVodqYDSQNI9ApFskUKVgzBSR8
Aq2EkUBXVMn4gC8AXXXGbzJhlRM1X/fRw7FCr5E5MyRp7rNp+PnUZdsjy+m4s85jYypl+CTOnOCp
1Ah4LEZouoC7Kx5IGBK5A2gV4LSQYDzeaKqZoDWBTNad6tz+yRzkWgmCSHhWGhNAKVP/JyjgWccl
CSe6pptG6V01dFDYe0DuKS+XwPtxdF95MfZBEX8xF6dsRPHuh/NpvRkG+CldHY0N7Aac7PwfjQrw
qGYfxY1x9HLv2FU1GUfZhHrfwhQ2AjRU6HIMN+zGZVdN6NWhD3VJ5KKrNkXsVjf0I33DsG/GDrWe
vyHbHX06h4dfqBarZXTusIpMwORyepZV+uzpsaOhJuXUUhLJcbKr5VtEYqbx7/j90NmJGLX7tjNB
q2LgYWsFCYFF1e4wmH5FgfBOYezi/zMRGtU3qG7ouC+7K0YvXXilh82dGltC8dZN1m99vjZ4Q24D
NFH/ub1dW7rEsCKNyBs6RWl+W26Ycr9de+1oZfLj4Nbl7luRf+XyQKhuwDvnvEGBWLQMz4JVt++F
oJC6zmpcT2sUyUk7As90vPuxphHNFZntkJPQXrykm57qNibourTfMrjwyoPfIq6jYCi/rtJJFFHX
LqtXJx7kNrIGgOIAVLmVKZ0O5UdTzZbHDt5UlokfBBsg72ci9dWM8s6U0CDzdoiYaH5lluWSHs84
+QAjhSMxWj69BFBxiAhOHx6zCJc/1LBLmeVEVd2dRXhB95vycdzQbYQ9fU2uQUDaM6VSTIid5iCg
8G5uI/9Zz9m+p6GenfRwZlM+aYqhz3y74yZx7r8giV99n6Eb/Sq/8Xb7Y3rpnQ+Wa9r3KDkQz1/M
5XnECiqWR/o4sr0KKXd2Qgnda8O3iwhC4LdpPm2QwhUdRJths/MqRobc6gLL6KR0C7SJejBH5xHN
+eSrjKdw+NqhA8cedrO1GKBr53IaOtJIZ9eKkdP61gimEGILyS5jMgzx+hH3FF6nZG4Wr5/KjY7h
Rwg6oWTPUSZuY74D7T0MersvRNfymnAFAHhHOcQjwLT12/8jro7OqFjynA0A8ADvPfcqy4qWgImv
RilohPLz8WrLwKBwdT1kJSiejuoO42/taIHoe5A4PutJkcGHnBehtZPJs8tplZ2zktJuw5tb3ANT
gOouOHsCtEIO6XjAV4ZzrUJ635igptWp+5bAjmcw1pzKn3sdr0Y82mdFOlJjHkZem897XTP7l/HS
DMTWe103wp3YJtP3bQVnsk8RwU/ByJegyVbnnqVsZqoNZhOQA3Qj3VLTlx5y5pFyOG6DcwB1h6vc
5z0i0JT9PLUsPuPtvUDGyBQyPsLYqOYDmIhpolKERypEM3/yw421SYlFIgssLUnNerO0/E4dAjWh
nzyYmZa8dh7NtMFl1Buk0e/44XgWYpGkxN2PPT55ot65Sm55ev1h0OCwPjl523bklPrv8S4HRI2g
qZ9zzlLnYJCwGBOYJJ/j7o0+bQx4zBzgEwg7gyQj+b2WHqWW2L0qqOsD3BH9l143pqAoAeBX9PgA
QjXH6XC2+WDsMb3OTnkw7e57vwcNIGp7148k5VxULNPYB3BseWyOhwThUQ9ZvXFxig5Eb8j/VrHv
3nKe2QaFqIHO53sAojRuUAESx3vF3K/lHaogPWbHmvsD3xGY5cQOVvUuaBbFar7xOpuupNytPJ1G
w14EZTxXccAV2oRpakBnIsRaTXCV/31g3GAdowVz4lg0QIZKTye85k4xnSVSmHzuuMEukCuJOQsl
n3SNdVHCb1m1in+tHgb51fO5p9t5Pm41b0nKnjGCpCmnJBR4BIXbNGJklorJirldo/phx+YHqjmL
zqkP2MCwoCC3/o+o8W+SHHg/hIKwvoLB6/s/XbjlTm7E2LT8Ez5DZ/2sVKmJTKZEYFUh1sK8XIGd
Eu23DsS0lT4EKB324rhto/YVkq4PjNhqv5EsdJejfTORUZjvAzuzdYqHDxJKs9IzHcjmtrAj9Yub
PEXcm79bD52DwrlmB4SGSVRgiimxYab/4cE9iWeZE03L5aCprAS39UddkjvccfpggwplA3ePVoby
lB7T3OP++asJJjDrRh2L4O0NDXq82zV1AGL9MJhExRhMlwqFpAJqrHKgERQxBBkS3pYXtL2KD2iA
EPfTLdwNyDL/EATqYu0VjUO/VMKWKnbAXGEoC9/3NzELByyc7Bwl6lvo15YrzbCXRUckY9Topl33
SxewWqmNX241WULuUl5oM7q2F2irxPHBGsuKJ0GVy2zCGlumPWFEGJaGVjEuy1jCqUe80PJmT3YS
EMpSbgmaSZhSAlUKlgghEcjZsD24YKWMaLtrMKpdnCo/w4eoR8TzYmj/0qhxW2QsDMEdfgNIq2Lb
6fDiV3ScFr/2CYnl9yPeuHSIS6g/T6NOFA+rz1v6oyRyXS/o2EWLXRxXvJmFzMnQeGniLW9y3tBy
Nct0fyTYo55coaWHX9//Kv9RfAEISjHW6VPXzQywPMY4Q1LS6TxgVOXBCNKBFQpClf93KoBHougT
Vv4PaGzFTfA8Va20xWgN1nzKmF329qUs+azd5Lx8SDMzvGU1MCUsNvYMOdbp2RaLgIJ8rA9yKW5W
OQo5gBHRuSGFigGuuQBFWb7o1C5V9cXDyMnLCpCv6FnKYMdIkRv+d4La4ieYvgaTEGHOdUkfL1Gc
BuIisCdx8rr3z/nRDV0xKEGhmtgFf40qhznA14juN96y6h8tHTTcsRpX64A8pLkrqe682pCTqCjp
8+NDUjo+5jkUWjygq5kYDgfLooZYkRimN4dq1R7JpGVjTdswin94+QwXJCOzDrkt55ifatrd9pyk
/rXQFaWFR6/2uaCO+BT+2lG5eS28b4YBRn1Sw8FY1LcZ2qGCCy/sxKjYvEE63bndGiEXtrATTv1+
NPsswOTZuBsIEb9qoaCK5RGOHj8I+9TRtGiQvWVThZHC6RRN71k2JnklJsqGihijmahIiGiTCUBp
/ITnnDmT7qJFbeo5sFvg9xe/4TWf7KYs8pd5ZZNed1j2N5rtWT3zXbvh+Z/GUGmyVmiNeovii3l8
ascg2MmswniOcFtEEvNmoKpK+xpQix0E6fvIIG6vySKd5weQJKv0wVo8U+wSK/4Cl3e9EAG5Mb7y
Ylg3Ztw/pKZJRN+LDnLoGi80H1O3E3YwbKJlQ6IN6x3ulxOp20vy+Ee09V1dqyIFPbeGp8FkVIGg
TLB+N4/5jjl2PtKK/8ylytqpX7kULz44FYMeAnQEG4hU3ij21iS0DHt3va2OM2ZJlEyn/HBTyqWx
YwfHd5CDWls1S6do5ROA+7Dn01FhOiZhjvX/syt31ZXRO5GVqtzf/I4dtjfzfsmcimjncNhbU4lf
M9eyZHzFOpVThsZWEfhlJUx9RPEYwzXkxo+bBOXDrmCshon9exHU0nquLOioWUTltP/I5olDVCo5
HEdZjsYxs+bow9Msy5bbDrZVJMNeogg0OKHpp9QjDsoIaCOjZsdbgU2YVamkRrXj75+INrBGpWs1
A6DCdEtya6hhOTsWheNXmBbNznPeq4b1T98boNBxPB6HwQ/wiDqh6tNqsOvmUQrzoRlA7TjGXLnz
T6wSlPxnfgpKYKbWDUg0VZtCEBlVDecpznzdHYbbk85IDpGn36DCAp2WiHhsdOK1EUBjWm1lmRmX
kvREmy3xEb7Z2e7vKpc/7UpFJBgcKkLAPatXrofv/irvx6JO6BWgYtOrFN3G1fIDsjVVhKkpRe0l
dWjfut9mOq8E5yJ7fezndPXYt3kDYI1smQPecnrFyrX+Cn65pAxA5HG/O3+uQuw2ndgsLUAyy25c
gUT5pX/zMrAQpPfCTcfxqS3wi0+ZBCX+o8u8btPp6RP8tyXqyAvrmeKbYA1WajTFBsTUwg2EC+yz
CBV9jfzMw/8vTJtqZp0RVslTV5sElkhC3mz1YKIKhUgejSTjAMJQmIdzd3P31ECRXw2i8on222dH
w8VTfXchOB9qALq2u8OOfst/tYJ8mqKx43BJg88XAPiWkKzRLm8Se+vsZuysWq4vgiPX11EOTFyU
Bbnvc4n3LgYsqbCiJ54MutCdFKguOW04JzRnEcsddflaznL/9+dDC3I2XtLfqYPu2nohq8mGRCdf
8PdmjcAoPHuF/u8DJzJ05uYqOxswEn9CwAfCa1b3NuhDwHptsDAs3FGpbvm6/unw4vjx58XCU77N
NUeUxFS1lQDFWF4qGntz0ybBxlO1qvxeHHrFdkn0NHlNITdj0GyboAc0o9xnyxKY8wNS8036E+E6
2uNqz53YE/0DHEm5kliCKt06uQAQxcG/unusAUpTOaPC4pezSigpsTCGk0WhwlwmoYtNxRCWy3yU
YkcMeHitaJCcybsqxxYtB31eYES5JV9v+6QyGiJ7cCTJpN4d6r32+O5KWrHlDwx/Dz+T0KfHk5pv
jniUvBBnu4ayUYDebzs2KDdVHdLYZV1dAJBX++ID0WBUooetPvItA49KdCsU/2i3CiapcAidgEBn
RIW2wUH5a0BowiZiiDj2MS517rH2DijpZKgmSYG06Sbnh6RsQ3Qo0qF5va7B57C+pQ85i7lsldPh
GLdWMQ0oAX+yoEdYIn5hji2xjuxyvnYCBH6XtuEqYB5Nf9hi06lKNnHDfJ4/7tsgp84bNt0qXs+m
xsMZaN3bGPVOiyZcVcS0w/SZnO1ZmccDrDdIjUrdgafSsppdjacGu1lGqM0B4pQyOMzwSIAF6nEU
80ne8qm0Uexp6LHR/4Snbl1xY5rkNUqgKm0cYbXteQjMuCsAgCkLzQp1C0R+MXDt8qNs6ViXZwEL
28yetKwk0T1zARkjKQiJ4AcFpAuRJ0nRyEz2C2OvWTxlvGMRwufFKG94npnYVCxx7azzUj4lqL2Q
IAjdVvkimItkz7t3t+gln6Ehxx7yPytBjmPuz3Eyg+eKI/s6+BdOV9pHze8G8vdnKqxXjTmqsUWO
LcYlMn5kSJlXOgjYR70MYYxp0e4dUXyyHWFb/Ovbq9Fgdfawm93RK3lIKUjtsSdmcf4dSMK08MxQ
IDrgRHycrraEsFiLfd5rredPtWc6BbM/u49vLyd+FHdXpqv3gRCuny9aL+J3Hc46dJu2ldS9dbXt
bBXzGkEokfJ+TejsQ+koszyktUVBJzmtBzIFCpWBlYZvj7XAtNKQkHNo4HQfykQZgexuqAgT0hdt
8u9/e2tz6bG4eRlgH6v+zh4h4b2HPNx7UMQNYuaJdnnsM4QI7Vh02dqBo3bAUwCYTXhWgXrL1Mj5
BzY27uuIEWpAMWzMMfChhjA6DLvYkTsV4iJpHZykO5aDVnmC4owWU3nE0bGM80zHJy7v3US/1eqd
J2SDiHSGvTLagrCX2xV0E0FEJY1gb2JhcuEw2kJTZOFScTi9F+MMeOj0aozb23FpiZ8dd4Eg2sOw
gSogH0BIo1K0uTg1IOleAokecWAAbqD5J597gJ4naz6hItl53BpBzYgWHjREdTRnylbB+HTGIGjt
lzusSP0TGcbM5jiiGGP1+N0T6T7Z+Gt0+xqGzxUTcEI7nIh9frKj3CyIShDnBaem2ECkSwEGnyKP
NQ8/yrxIiwZKy55e4CZriw2ZG9SkfHl7tH2tlPwmzkRQeNRw52/lNZxfq+dl5gg1xoHA5UY5wRD/
kSc82b+/geINqDjXBvkfzhwu5cGkvxRu5b+ySJYKwTtpUmcDj5sOgNDOUMHaWi2k2Q4xmwTf9hRZ
QgNIYDSCTzZ7Xysj/F73NnwdPauPGhq7Sm8nivRFH5rj8Ur3kvq81ADVj4LqfkOhlfBtuR0Dk+eZ
Fr8QbM5B2910NF4SbyqHMlx2k478f3/x97L7kz/Y3R1vG9heI7FKtZHjsggCUfIT7CQZ/Jgrlonq
TuSdFw+IKKERmwAt8Mrh6WfOTJfxgnPhz58iwOQh/k4Zza2vGYUlQU/6Unk8wG4hSaS3XXRuam/u
TThWYoxjpRIcAN7UmGTFTKMIru2kbdoybWl+ghLq7BNimQwnhRWDJLfvetKtbZY5ByZAN6cZfrgz
cSknmEfRhIkeGx9AWEXLU3UN5V4vR/sinFvxTcg0mlOxI7eq07blTrJviDjdJotbB6Rrk9YcsKAi
LLw8kjz3S/76KAy01dIaHf7s0VC3AdohlT9e1QtU1kjBqYMK55ZhZw1pmhIPS3k7iCTpME0110qc
aGprdj/9xlk6qVe5OGGdlfRhGJVNHKkimYzVvwICeRb8OAH+XumlYrNAaYaUhA7Mzse7EXKK+xy0
zU25Z+Ewwm+yOMff8t5sFIQGuvr+dMlSTbCMGsyQnGY7IubNPAlStP9h52Umrw4hTu1wu7A8OYaY
tNdiw+yoHglaUH3z2BngF7bd+0kksYEXAK1dxpclivGPDrKL34AlgaSFmlGfvmyK9amF6AAAHfoN
w7JljuOa6ETYqwK5fASHG+sdySOcYXNTF/cHnvScUPQ3y6ZmYeYFty64hYgQ9nC80X2DVa4TWtAI
dI1I0dAHbkCKE+qaMc4mIBRYcKJV4uzeBrFJzadh4NeEqBHdVhdHg0UYs9Umwm+3gGpEJkqVGHzW
TE+NO7C0KdFo7RoCtiv52zBAGyUF7WFw9UYvcpEmPu+aM8dKZqA8DYPkciA9uNAWBLJyCWr7yLIv
oYG4GNSaUKcjyL7eDG32VMGVPa9jUFdYtqoTDsq5Htf0zgL5IVLB9x6/HbJiUJP+8ZgpHNZEd8Lj
QHSzsreOFFzAjJ+EWgYLC0s8SrVQ2S+zV1ydXDHTnzZRc0TvxLOoC5MQFuKv1PsMi2CNfzsF9u6R
UFAYxDAZko5t9UQ+sp8c5uKrU620ydnvcMFMsbmlK/xj5CzGNFrv+hjm7FG270PebYg8DrF2sz2S
ib8m3dugttvzNnT9sQ6raYl7I79590/U6UG434hLvhA3GnVil5bb8A2HXNlgmTDmVy1+0V4yOl5i
aIXDpy1p3p7azU+XEyY4GqCuzJrLiVJC/0iTCJ24byPJT91imBiD7FYdsGegriSIOcqTBbjIejtC
LWdCsHtDgVFcz7oHZnXiJQ6xeDryPk0i4OsaHJsNh2Chn2urbXgMUttqT25zbdwnc2kyYob39rlS
PZcIRpRrUK6+BHuFrKgOAzYurbJGrXEmPEvKWn3S2jP6IOYXfG1eI+mtv8/ESaasMbQck0RnODXT
gokPhdT0lUWDuHNlNjkD7gSa0RPdyBtLg8Vyad6cxoN4TSgMs8PdNhP7d1gHudkORFpdyN1FiCZK
yyP0NKNDtyeidbnFFSqdZsj29Jh+cRBUITsuKzVv5aS/NzAAdHvU6K3cDEZGrfjQOJjPiaEEXGjT
dhMVlXTZ0qz/JjLDsQhG0f50c0HshDUnkcBhNLY1apJ3b4rqXariSoDmcY7TcAbuk7RjYsGtLa6g
ydo/1yS5BJIqgmLODPKPc3ytEZThBQeSTR0k9KdgW3rv1ocgRJz+bTSz6TR20JsPU9Q7EcuUt6sa
a+v04IKJBEqtxKSVC/bxnHORFsZWHOgBOXEAGMVT2z6WptyM8knkUdG7EFfEXlIdv42swPK+jsZ3
5b/iVJ0SfFrniYqN7jGJHB5n+dl1sPBC/wftq9XKSjYPW3B+BYNQxqKZwehbJ4a4D1phvorhNqMn
WmsMSw4+U9qjM8HevGmbCCpLGtXoD0+vEJljlj8PtXFWzPiB2+/lsAX2CFR1MMXFKnNXXtEGtVvX
pq7gCgX3u/oIUA7rVxDEu3MXVnJwDXQHwEORnZZVG5KNdTBmb7i8J2wXshYokorCGE4nwZbGZ2tn
1V13045z3AvIdR+x4ZAA3i0W0jmg1uXuNExRHCMdSmJC81ohrxq0Rk9rbGt7DzfnlcStWnEQgFxa
KWlqu5euKznSn8JRA2aublS6Xw5/BtDr6SKYUhuLrrArouvD7fxdDDkd2N99Y/dVgradjMyvDfV5
tM9/Dfl9IbKoWg5gujtuApH4oSd3Ejln8xESPqYRIoQMcwIvjld7vlGgfiKGgDsbfMaOwzPAr3wt
vXXeLuUH20hTVT5w8RfQ6pwRIWE4rDpK8esXHPPsLhtmIXilSESyGYZY9IOUjvc7xi9R6yYdD7EM
d1u+MoII8IJgLojQlWbqbyQIylv4FDB4gjEJ/uQVf3zHG9+Uhe5AkOGKwe2Ug3nUlbXk28/wsc1h
2/M/f+s7bbku24opczNs/Lx1SyHco9VV4DgIsMHAgb2yHXGqrV6hCT+Qke0AIsmlAHPp1OLXRlYV
Im1iperF6mPy4+QOOo1u1SYZOiLYCjYmar1OnGh7irahP8ln212YxZnNrm0W+LnRX4F3HvpHff8w
8aWzyO7yLUq+y43rE56SdJG6Tg/KwApeJqxxEHuQRLLn1s/+YMQA5yjNYDT38g9eWYL23SMFXMzA
Z9HhHcnidkf4hAYFjLy10G+xL5bHyH3/VGLWY3VUexzqBF32g99k5lSwSGIC0dMsuMqEv/smRlWE
ibcoaKIrL/W1o+Hz9qU1DpCEfjyDpYLbMHv2MR58N79s4yAFZXNzY80LDNwRtlD+WXMIpqcAIug/
RplynTfDIsIVjIk436a8Gk4b/WpYN+A468LaVFCu6hyo+5iCJJez5gzhDJB5QEXgUT+Db27m5neq
T6H3fpx3GrM8yxp5clpIfy9ySKOJE5flKsLfXOUrzmUKx9PXl8dOasG8Qmhki4lmXPYmjaxsBAD5
HSfVEyjQ0FTPQWOmmyq78gcCvx82Uh1mhC18oobl0DVZMlPAdqMWIWdilgphQy3rHfdpIKAKVzJb
u5X6ftKeoKAR7EcO5nsIuWfcinhw3e5TL1YfuKd+j7krI9ZhzGeuHBtSHYPLJ9L3lmIB7Op8Xp7x
yY73QrMRLbWbEJRIXKOJeHNiQypqmsSEL+deufTlMzHpTaToFUnbMykQXVpUWFub5TOAMVio0LgK
Dd2DgvdH3beSPnQUhi0v18EW+ClLRsksCXQX9At74sgN+XCLBqryZzadiDzOGgBGEc+/a/LpL0Ue
LfkOLDPdLNf27Q9cvd7CHnE0RTPZGgC1NY22PJWu+7H8FlE/vyMtcJpUg5nmvm7bL+Vx+jswadqY
cfbxXepnjwu47ptDlMoZay6BGGaajIft54EIHfmpCsOPam04f6rGDyBmRZJ53l6NAv60UfR+AFIS
s9Q/el9O5qzL3a2AczhlGajdj0RFoarnz9gBcLLXNsfsP9GQdOG+f8+N2JPAxk421UnHyBK2Yo9U
/6Dgx8DFWzYgEKuArpt7z6whiSdV8DXicgL4s3flCaW2NFgFoXcq8HUa1I3wIdceARzwUBuULLe0
WMXNMa7OJoyyYiKz2q/z27N0NjYRWV2OdiIzhCQ5IXf+TAoC83rtrCRNv8cEUZr6WwQ6WkkYNb57
U7HkfrppEw+4QDvE7JPC+iTbGmWObGA0nWtVwgDmiIMYwB/QzgabW8jSSk5X4xwntnO45RGjGCH+
N+Ax4f638gKqUjOohIEVVNisP9X701GOq1vrULEnITxbfYglVlEm6TlQgzETzglrP+xtwCMhUR6V
BTPMEgHOifprlvMzhSulyliOkPJ0JV3gM+ZdHPYdQ1q3hTbSXeNjAEBnCMge30N/NdfdUD3Z8x0a
7Lh95qQhc7Kia7HUzx7mxPARRSdBM7GsHkgvy5Rn+0+iST3/HgXduU8sinVZwk+8UFfW5N6v1Trk
R2iQHUx0t+hzCnt7g0/H4V4HTu90ApvCYwCw432JhqQxxjE0oYxnKNJ0M+rPFIN6EVjGOBVl7BUN
p7JOr5xFJPr2vebosga8hLjyo0orX2KOkelY/On8MW0r9EriDMYxR6fExOdvWkm6/OSEy6jgOCA3
qm4f1/Vcq4+SgiIv+JH5iFJAhPqN+JlkRnATz2u5COCd2/BAJVf/YokgaB4xtpFyypr2sallNKCN
tbx8GFZAUzQnyWot8Fqn7f4+9ayn9PaTnu4rbj2WFowq8TeeD530gi5RaUOtoQ6xENQtNyHIoBpG
Y5ZqSgiGCsW9k3TfkXZq8iVPm1zMdJTiZvolv9HgOLlKwHiPXkkgsDbm+NFjT2ze6C4tJEuMz92/
DSXlCNmLXFBdDqZQ/ARb0vCU3OBI4dGv8EsCwDbeOsG0+B7vcamjY9iNuQCDSrrUZb4CYZ7a0ozw
EWV1rgyNN+hMlNMaZrnZV2nFKfU6cWU15xf7QQUrCr8JwcG3IYVG6YTmJg2C5QQxuguj+wCB35OH
AK19VjrzH/lUnTg/yYrx3rKN3wJDnq9MK5SbJxPT06tbiqYDtPHQjGTFCoF5DxQ3lbgLrs1aeOdN
3oefJtnSuRLbqt+bu+J6dlgZMAvZ6vkf0EG2t1SJsMnB2Jb606lZGgj404fn6zcBvRTQg2fxpF/k
iAbgu1prpKl8sMz5n9loojLznnPDamJEirYrIi1QGAeS1oc2F3e+mq3qrGXOdpUorOc4j1hoB5YT
UZ/bTZ8hos/XkY3sSvEjxytHACNI10m9MSPRlOdO5G4YfnK/aSzlhMsj0K499zm7JBegFo97yidb
jWem0lPXzrPwAjiLNVbvZUeOnJHrBZz9GWUg4uAgyKqLSTz1wo+/5gsv1+kzcLehtyfb6Po1GFwV
vDRw2k+QZt/LIYYVIgAOd3iPCUABMmrU8LK2d+a1th3nLT+eGKKISWCVd3AEJE1wTn6ow1e4eXKQ
7kw3nhpBuz88SbOvMnAsp9G1csuYsmnnFPpnpD0MQbh8EXtDM70DOikKHlLD6db9sr5xh7SW5eyr
70sVI6fU2NbBpCLiK+8ItR/n4E/J7uV9HvHmoHgoLfa6vxt7lkVgKBdwq+GkoKBiIIgX/Mt3gHIB
nP0ovulA8F2Sg36NMQXtISY1iqe7eUQUA//V8ma0wXK/t77sWRvdr1hIEwDWAFCsVvG6pDXAwIlg
2M8e2XCU+Ee3hMnoGnQQzdL8bvlGj6kTdBy91iGQ1ZAQTeMB7Rv72w66tDSqqj9+LhJYfCYoeB6f
soWaHCqyYpW0TKP1CtnIZFI0Hfk8In5GxB2HLIZs/hEZ6QpCsNQRoHpH9iqvLBa+MOHzgSqMRXJA
jUj8jO6ZJEUC6FvmUoahsSGNv5svEUXGtyZI791rg8W37nwzhjVG2AoX0z/+lgdpQagw/jRIT3Vm
/Lokqo75r4zzthrZASk2x74JzJ/Iqo3E/FAAMjoWHvMVuBA0MRYRWjjnwT0pU7PtP87AVcH6M1E2
lyCmk8nfMPS3ZMWU1v+8bkWbTmnt/uT5KNOLk06VKdQR5PongOv1bRWai3jWpVdhVvhSBDFNV47F
/5U+ropl+shFHyr1qYo6UCVWwvHpEPgCTk5M72DdKoe7j5bkJaPLNcTXiMh85xhtG2PVfLhfgW+F
x5GtCJ5bWDOXGr0Bluwjat3yaiGH9WqgbKoFHbmVjFjKu2hcgyYW5hxMjyJIrDxibmbX0Beq5uhM
eFA/DQqygzOibnSE+EVB+a9KH4OuSvDIBqpu9FK2sk5TCKjcTaZapZURbtsblc4jE76wcUoyLdsO
T+Y00kRL31Es7vRfCt3t1H0vvBBBvScmrv3z3q2kk6W8WN9DHzCYcBkx66Da13yflmd8Kd7O8oE1
eE7DLuK/UjnXuf3aK+Liy+XcpS9a7ZN8lApjPvSKywx7rejr4uQGYI3+RpdVEmvQ1ZgEHlFdc5g3
I7bJdzNlgTP2Ok5uKizJLfnYjEsvhSRau7S2l9iM2J7GM5MzLbMZLG0xMylWzgDFx5rYAN3hOJfo
C47AWCR5UfNUi0BH7z9m1dTWZGSxDDa2T5Y20CIOhDdF3wRXUbzvBhTzZNyTUIS+WpsIpsphVRg7
Kq7fd8TaUejx0lI08XXgc31sGaI3mlNES+Z/y757AGVb/IQSMWjzg+lK1TRh3g6E11wd4vOOss1X
nlZsdi1Iy1NXz0uIUZhTerHH6ky+HxcGpfbG67HY4yxi5NxJOuiW0Oqcea0SeaJ1AQU4zWynlwXH
tWxd/qoshrWzxFt33BbgEf6KN9SfcQ4+eUvSxk+NKTuWK9n0fNjm4b0SKnP/yKZ6h9gx5MA3rdiG
3me+9Avna7ansUyvpIBfSNMtWOyhsQ8y+sv4DJvxchtECaczzoXbYqJs1fxcH5sIztr8f6/n/DoE
MzubQQ996uzTYKwKduBOYzxkr7msoCCqlkFqWb0MLc1vSgZtUN/iYRk+cQsyfcbbjXYyGGdAybV4
lmoQhJULjXKT/mOMxLb5l3CXFmTRqvRaxxwLvKPgpDkzZdrSF0EloHzzD6LPgaqHaftBDe7BprLA
LGqK4ZuHXI05irstrU2xGWhLY4dV+RwraLL9opMgC1cRY81yidiPP6ZwKfLnWQLeVNKXsKriP6C/
Yt3XQDa/2gCiU8odkWDCxmyW1oOs1fnWlYBnF6vZwUfudWq9LrgqiTGdkGKNHajupbGKGvLkzYkx
9Y48R+O50MH7UTt0lJOuKSoRWthC6gzNj4j9aIOAvrwKXr5XV/kLoqbhymABDJaA5Y5vRSt9Xgjv
MsuvUDM3YIhtI4Wh+iz2i4SCpqPd24PwGKHBx+K7Nfdzkub8nol3AkesbD4+QH484monObFfj2wr
HEPc3SQXnFgzkbkLkws10kuwmtRUH+oKcN6a+9mtoZI/1UPDZJQtJ4vW1isbYQzHsCrGQJ32iUmG
NJ71HJt0HpXAEXR9vS/c/GaH8IXjQoCu3QX11mwVE3qsq5TchJklHjZQbtfJHWd8BLp1JcMzmomJ
WSW9YBUD03aAF1vS5bO5fu4HS/N9nu00MhhJcdYiGXS/NCdczjiyJ6VXHX/ccSwZ/3N+H+4xCu5A
lQCzsFnDPYDWgfELRPQ07gnQtZpNFeXAQppCpBCFUCXBxB+XlOv3lx7L8kca1LexDLZE08is2aWN
Q6LpelpPx5KUeEJmj9b9u5WLCnkQb5YkKo2MZHyutyWs6+ABKGd3QO66dCMp2YDP4IK6AfTcK/sP
NVe4FNDBu9qz9AsQxGyj4nedy6dn+DEZkAJdCYDTdf5Lm/Q9FRz/vp7Q3hWJ1gk1cwgDRj3Xa950
W6vURftAJNdA1hzW7JdFXaL7zuKITuVMAld3k8bSf8k25fs/k5vH8SwbdnAYbDwYDR81X1T8S3an
+3+rMYMh0e+2m7gudEG3X9TR6jnXi3bzYRGXwln0aFdREsHpfDbfspkV8tnrgGkkIn8z02zLr1wv
7NBsQVQ5ZvQsv7eAuefUt/ftrT/TsNhomdcVCml0xkILOnKDo/L4Mgjwb42+VPhlsD/wrvafIu71
q7EaI5ZYdLTFee3FMniZRxCtuMFICkpCD8wpod3Zfisdb9Yv1h/MbLBvsIhsIrENOl/Kk/Fpgi2c
xZsSqP4arUSR35GRsbKPtJn9pTUtuzgCjtbunc5HGCXhIx9UV9+WySihLsGHbGzfqHjGEDi54w31
DjPXsVMz2NgQpNdDeO2DywPQsfLVejPEaoc05iU6vFYtdf+RJBmqy1yTWbAsv2a+RPOsCr864pVi
L32U773TTQTqiORSefjn6Ukv/oSg6pf2EMetfSGY8olRAm8isfUWpYeFUcsD3QRo1NJAg7ImYBeP
AcRIW+53Mp2NtRVR7IjwEaUWfWSOIW6DXG0cHZHb0kDkkOTMshKtwlPPc3+i1UmQNeGqJpIi6NMT
leBO/NfmkRN0bu0xIXZcVSGinIUrxAqWdhbjhAcEVtrB1iUiI/ARGvlBK+KCt5cP8ujEBS53tUPx
igqgdi6/zDHNa418jdluQBVeSrkPtIDTnfSaXu1JX8gO8kroPVHUyIhD2gVjq2C82A2XY2+mdKnV
NF3y34zsOEryrTRWFXrSe4WDgHNi1yGpo3hoUDbcsioY8EGIy8kBZuvf2zzW+a3hn0d+Bxa72uGe
lsBAqi3pNBQHuyHoqk7c7+0FVCFsGgEEZWsiurqzLyfF27EHl9hoiCKXMQow8jzIrQvoMG0S8Ozn
3ELGzeE9/kfgtf+tTebjWU4vRKNkczieszh8DQxcmJu9EV1EAcChlpYMM8ReaTPuyMPuGZuSU3jb
9qjKABaSgW3BXUsSrePyssZ/u1YC9/no20RpGxDZPffSf9egUK02P0WqlBbJGy7xqVaHCHuHvU+p
8kpcwCfg4hWnR1Uk7NggHcGUB0sHG+st5IRln0qpmDXBZaaNnXqbufFlzOyBU4nge0sLyUzHbicc
QXleQVWi+bQ/TaKzXHo67pDs8naKqN8qkvCV5fA5YDn/tgoH7vDa11+bSe1qbHSUgS6x6/ZLY1GX
9Qb/9CFRBNYY2UMKtDp1sm5QMOQfHj7elJMqhCP9ayNEKG4rjRyvfNZyXxE+ylqJ9FEi6aTEpIZR
fwEvKjCkrKUCcO/YJrBJRhZf25X7Xia5GwUleVUM5MWKB94T6zHpDP32aa/S5gJofeONtZB1BcAi
cVJ8NmTrg3HddHLiyaiBrW5htVCOJRH0lDi1n3wC6Vm8xmeEgLUOPqoGV5SQ8rAbbxnTscAM+vac
ZyksPQY6APwvhuueAXpGuw+Ri2vbM0B008QH68j+Mde6fM0tZsY9lZYpIj4bAG+YWlFJ9PqqiO1T
LIP7t6Pedr6DdpKd9gkOM2iQu/LIUiGOrWQCLCHUF8pWYIrJonwbW+SP8UYsam/sojGbIDeTPsZY
GeBVKtvGiqv8Bpw2jSEybcUZsClLODBIGYIko+RwJUg+YTDeD1WTeDnH5Qwgc245mgeYIog4xwCJ
KjhHcijgwX7jHo8wnreG2y4rxLUuMkGE80qmDpTsjNMSJv9H1mqhIxI3oTGX7l/opm/knJWwcoXu
KGm54wUiGzB751Fnw2PHzsjIYI+lGrOh1WgPCNwbh3wm2P0IYavBptZPaCXrIhrGJ5sJ3RaR1a2g
UJEJjT4KD8EZAX+H3tZPkHHGfBAYDmGmACDAhwEXmczUe1j3Qx9Dho8emmZqOIh2izrQq3MO3Opv
7GtsZvtDeAz1qUAGJtHmyD3zv+jq+hhOO64t6s383nJJpVUnQ7R1jVBPVDzx4luKOV0+7uGDdCgc
397skNVJxbq2T5YqRhLIrPT4E8yPts4a7afvhUdgDr3fCg8khvjxGcWuZsZ0ujxxY8+ObZVSs1gH
F/yDDMV2zcPZpiWadEneEycTTRaD6TxJ0J5+DytmWtIs5trh+BEaOd2wY2wAnrM68LOFZyPjZwsg
bZB7Lpn0nGpYjtjCuQv2fmqxQaoptcJj+fStZN6Zg5TuTVchUdKXuWH5tDPkrGrTGvTIC5QqIxel
QbMDaUVzABUp8m8bcIn1A2oOKhhydrhFuAgouICt3lKlKDYldi4nyZHdGlDuOZerZJQlGK0rmbOQ
oXNyetmnJWxmF8pa+yr8lAqvMngc3+yOseLxP/6zttseorFzsZ0kQBEw9GxC1dlh78ZYYrSYBjKH
5gjpfIXHlT43iHVe3oNnCJ4zYo5IXXX9QchIcr1fnsuySvlUcpLhnNC21Mg+ofQSktTA6HF5yq3b
aboAebhuOeFqWrBEWIwC+j7M5DtHCabwN74FH2a+qsjWjYTXgdzUUng2Tl8Jbhxns/ZMD8Dx1EIM
UT1bg7vSeoF/qn41aDEh2Tp/EvgamKugR3i6s3tCMzquF+6FGzdoZ1uNrZthWFHDW5YdP4Flm3og
ykgSCbNG7KKQU1ZZW0uHIno+tTR56EA4tiZOaPR92wiJGpAHSz9GVXxYVclpD7I9ovADsiEysfoR
qn5H0Hpbq5IqA2MXnHYtu2k7L+k/Jz9IVH6+P+h5dsCjLbsVDzzLm/pbNOlqTyg5kay2DbS7cUMm
zUKn1LQ8JS45o8K9v9A3FfjiYNy5GawCwjv2/3poLNT6PLdWCvRJNtXv4/TsCWB779uI2Fu+EQkQ
Pw0fyKZpnJoVGdwL2tx4oE4kfwObsikCkJFiY7QS8S1+xHDGleQGUm886PI7r3ZUoQQy412paCxD
t9iuIhYYOP7FyGj8HyKcE3fvGAbrMzdr+wSh7p2ZTqpllADV2WB94n7sMarFXJCDNNYzmDkBbXwW
nNMpP2t1kO9uJk89ewgQh0gDEOcmWPuTiAUC2/3tIBCBUspnRaXZzXOyJ2nJzZl9cyjVipOmnO66
Qr11jpNtJWTzt9igRLN8twN2EzMGyYK874WQ+UBzY4SK35qM8tsByAUyyq0XDROoDctxyq3VKGrb
jUUjuzsfyPOePaf8GETDuieeuWxNUF6QaDG8T2UEjvcy5KxoHAqeQONY9HUZivG3rjU2B4RhiPtx
k8e1+5nJoAuNz49YPFsIG/FT79NLMEQWE8xxHm+zHAGGZR28asvnLnJe6FlC0DoWAC7h7vrzq5iM
fRm2iXn5bLgcivmMPGYCjP4E+Lh5fr6cfOQjT8zZIcgOhnuI/yuo9flNX4sISA5+DTK3wbK28pXr
Lnrrs9hDU9a5rQ2VxGfCu+xjU13NzB0NNLs6Ink63FuDBK5SK3fZuvh0Lqg+IK/Sii7ap0MNFhah
zEjzfZp0svka/UdcJTP2viTv4BxKM+ovkZNfYaXOWWcVO6avpVrZuKbvlrVhofWyfUsW7rozDZ4Q
Ujq2kPCsCKSe0Qdj3UuTgyJNWrAoBLoK+D4yFE3rBJ2aEhQIbGAvbrDCxpdxNnl0e/J1XjOJ/0dK
gcXDV+bbU7s6jvm8Hh3oGNi13ZwjbnqR9K30Avw3xUA2sOWVjeH8I7jAeCmH6I7qraOjwV+tVIhs
1lK0HVu+MtsJ4yPX/SIOntwzTRhLDEuL9e6e1vC2G0886lYjrtXPVHqp0Ia+LksJPv29bE1ug0cP
jyQ5dySk9YX6+J06YbMdkt22OowZX7vzCEMPfhEZ6ZzGGiLEOp9le5f1w0uAyqS6ijrwDugsdXoP
sA1irDloa2PFnlxMJNo/z76dMSXubo/9OZz+QYhkbmWE8lGJcR+WIbjDox6BMUV1KmZ0Gnry4JT8
rXqAdQWu0ZsQ+F/eTHrY+8xTngx5dT1da0XZ9Z6RnkU+Y2Mkq3T81TnxZ8zuLqGYTM8T2r+Xn3KO
rS3p66mMSRxR1DfD9vOMQs0YZmt4X1lH4BPnsew5+ucWVnLNe6TyMK5Z3NKn/RCixqqbhR9/O4Ne
s2pFmUOB71tvbnghJovERkTdihBXUCxtFHWQzocVkn/gbjZXVTBVZnKIBBLq/PelavC9glOIUt5x
UPXfGif5onou8ivjzvbshniYwl+V5SjDwnFR7AaehNn0lECaBnRFT8mtcp6y97omuagNFbBvpqOU
IkA5ig7lOakZ5jOZOrYqw/JOpNw2Kv7yV0g2qJS3zn2I8ksacl+Jg73UDDnKHMSFCKNmk04a3ia6
ZB48qdDbzNMAFaSK5Rg2//CQVR4Jv800GwtrDkipc1B36Gq7gP9JMoHK8jwOCQmdnEQY5jLTmpY5
h1UWwlaT6MrCC1EZ2Zz5BgypEPeVZZZGq4p5ZAGQcowV1kweI7tWYpwTPqtkooIMb69/PVZ+WwIc
LQ7vQjK4IgN95MbaZQoAyk92O1Ia8Xyc0N/uNSgw5kOo1NOCG6sUT7kN61qXff3HtZIeXJADIZvR
6xrv5qPA8jTTwZ4vNEHI+Gw2zfdyzbDXxbAH6HNYJqSXDec4ZJAwf2f47WPJ4XfZgTo0SbGgWNe9
SymLikW2NlYiW2oTVyNyOGZ1QBO2Hs+hMDir1/+3zUNTPDKIXMxbPh4GkKkppEplseTtcid6RKZX
pta3P6MFWXidR1mJ5/RDzaq6WnMj5SRdAe1opqbjnALP8M9w/Ld6gmxWMbiwvojv+VWf0/VvhDoq
zwk6ISnCrsrDbW8ycOtjk+an5XdaGDxW4Uj+A0SSTPvLM1lYREclEMm8MnnW37aAfGC5c61lt/Bk
kmsRMvvEzF3f+00w7x+rskspmp+x66e/aapPppKyEzJzWqhMUTrk5M68bDisewgj4xAmHI/UPYFZ
ZvPRqLuddEVrmmRXZMVO86JngyT2M9o5R4IWvzityizuXwdMcWNTotEI7jLQPg7tWW3jxK2yC8v6
F+3kdq8bTEzmJzIZ1w3CvtF8S/rwXHHUMryuG8PK9RfI0ykf+H0GXc0P0RQxvvDVofY5WqLRH4em
sV/tVzO45dt+2RzuDe6k9ZX7F18SvJy+RorNIXkrtCaBMTVEvQOZVzZgVfvu0nR0v7zaNUfG7irm
IUqvL898XL32vJfbNyKK6OFpaBnI4opUoJttfY7XMa8atqgpPrGZp/e/ZZ6GrfVOZObqURdMGN28
SgHGQbpTXS4rBJ4EjJbqGyAA385VmoXMSnFsB7QWl+cX9gtay5qSbeNZwKlBV9Z9+OU5YIxTpjCh
+USLX1866r8wo24wLy1ps6wajeGM0c1NVATKTFJauiMxT/9e/A0T7tjbZKjrucCCW7bYrvcSBjIN
8QX0v3+hRf5u3ycNH8CY4mMli9uq3iXZdAQISUU7Zu49Zy4sQyJOIrVqfcuX0gz5yYTFa3iQECrt
laInSqxtFspx8xzI962ibWfe7h1cYAbNH9ehZKusCGyb8BJ+cOuDrJtKqjJO0Do++81ioRfrvudK
Y0525zZ7iSX0PTvA3AjvMTSKn6l7N0Bqd2YylaV98TlejsaeEhlXgz0ZBeiBhQE1asNIWMjMjhFo
VUOtiyak/NaM2B16AjJ0B0UIDkFYTpHzH1RfNYJbZUZ47HUIXt+/0dJ/KpHoBirBGdRYXsq+Oeso
mfeeetMBB4uxs0C0SM6Pie98x8Iy2DAtRf3rVMhP2VPLes2oD/Ri0IwqfNTbeLzTm5tC1yukFrz/
yffYdCaDPOQ8D3IiSl9uZ3Ni0FUdICyrLExb77ZraOBM88JSLioBw27I2FtE8nXu+M+nuvEkyehK
LPqlDxrBiMelPEJthO3mzSByizb+IsdhiqYjGlXN1OUy/0ZUwEyDgFUIwZDSpKdsIWBkaT0fG5z6
4z5y7+JTWyuFU09JV4riL1Az7/x1eVDC2dLJA43pAkIeHE065pp6TQGriPZG9gQYjSoLnlT3sxqm
BKnHtCjGoLuFQNoMyzeUVTfNJra3Surr+3NCO+tUf3GsFzhp/pwy6+VZEXjONhPhrFNcPbzH+nb/
fMKQqVDsluR4MCiwubcpJUyWFf/WgNCnU8032XjlXKkvXDVfEp6EZx/S5L83Zv3QSLMklTw3MPj5
lP4jK0+BAvIM+7TyLUruKYURyz3mlZ/U6/4m2BpzI0RKJncEpJNI+XiSUBk7JkxHZR4xX9dc0Ufb
BnHzn7ImX4SW8uN5oibAHe9Ezbcb47Hny1gJf7+1WNh+ta7LRIg79qes4biZLJVZ5jD1Z/R7+JP5
lvr1HzAMwv8WEyToy3q/j30S2WvOIkU5HrE3HWauS/J7fa6/Bq8cdgRp7DKVdOBS7/hfrCxIGZe1
7zdsOltGobCBY5JiI7R0U0b9vUAl07Q6c8Ou0Ndw6UW06A+IqeVaSpklQIxQVQ3sEgcSui3U8d7S
VPrXxlxbk5mEYIobG3d6CdDKyXpIxrQWeOZqv5+HQk96vsGCpjerIxAWUrADLUVDb8ec2OY16s5V
8gYp8WBHsdFELQ9prSVjOklFarv7thID5mrKS743ymQVZB2TOK01csZWrChGgYqHj57l4quzXjjp
41XpxRCfj8mAmdtl+EdMLl54qpEaJ5j/dqqIm6Le1dfTCDNU+ccgK5xZAi9kMb+/nS23TCfobHf2
E/oX4uOrgHYG1soHdSuc0eh37PVYVJStdEDmYwOEPATvl2o4rxd1sayRwDbQg+z0X9HH1GF2/T05
6E8Dekdunk/OR0/UDD5SRShzYJrJSX0xPh7G4qzhc96DTcVNivybPW5MYjt0YNH+HuzdW9j49dcI
4nLZn3Zj4A2cPepfxV7Tz/82tZRcg/elN0TMV36AcTwsCtMV0xmIKXYyTG/hbdctCMvwrUSuAi3d
GaIJoEckHBWDDEgHMuPyIjldrbrIJzekKcdtMoSQ7ImSnFt2K+pn/zmPq+iSAKW1Dwx+VciVhZY3
GS8ygRrSg3fkUAN6jGQDNArrkOPrXYjEujC1vQN9ub2pwrpJOIimI/Ghabj/3UrAYJEBB6Vq3rRA
IAtIqwaPRenFNUcgUhZj3xJTrcQXugmvC4j7BJwuqwzkywJyOWCBw9qShReYlKEKTTGT4qM1FS6z
dnbgg7XytUn06CYLVZEtnduzOc18mNHHeGzoA4HNV7mC7+biixskhff1fR1hzHySvgnmSsYqmXz9
FIVL7bWrxBMjR5+g8KJVh81q6Zjvce81Uk+fhh0lSRijJ0737WumsU14+g2DKGla1QQWpntW7giK
aZuC3yyn+6ytcUeSijoi7XUBGVlvmhdt1Otuiv+wkFsneOVqIbPEkj3nLo/y/gE0OYwOyithSzW6
lvoMC2BOSmvM353xD3po3pxt95O4O+dIvHeylF6veQZJadUfOEBD5V4k5D3Hlf1KWtwOHreYzN6D
oMiwLLfSMX3k/BJ6dPpK7lOxdiX1r/uHx7lVnJz9rPYcFtyHBCehUsxtAWPnCcX8sfGHEJ84rrXp
1KnH+M5FmmNSd30zcqT4QFClVyxxXq92bCzDJxxNcuHcrR/w6DOZPumLTNmvYV0vmhnzpnHQSfkO
4rgPJRAf69M4E6zEf2sxN9tMVSA2V8laHEkS14s8X2RsTBCcdvCH5VkelV2AGDMjl4eQ8BFL9osr
gdmyTkY8jT2fDbmj7kBRo7OyhdKsgRwg0OQjvJihGERpB+cXum44yHRGXVm5ZNDIzzwNqFk+jj6E
EeJ09uw8wu2RVb/k2LjCmOzjCTxx5ZKmblOT9RE+F1drD35qOsDUAJgdeEzz9jC4cMOxVttq0jma
3gPVYkyDWWXq2XlH2kXYDHAelSVPqbdLBQZ6+wUIC06HhjLxZzYwDLad9PbOGzbE3CHy/GQ+M/wA
s6gyVgKlvcXQ3Zp4BTMmaMmENkxb4xi1WEKFhbUCnpFJxLtJLA0jzyb7sfXHgeSigjG0kiIEQDcU
qKGZBxPJ7hx+3jLBacjIsRmiZ4TXBc+y2lJDmK1IAjjgtAZ6v03Rh2NDc8Ox7F0x/mPMyVDaC/2G
ybMAqTN/QpV/DB9ub/AAG1InLwcz2Fsl0wMrO6nIR5jX/a328xEgIbEkABlHjIBrueQS5rwyqE43
A/2GMkquayN+bZ4Aq10Lkq0Zr5XB/tTl+Zzfiyige67yxwu3OM8xE/hDSvLue//URTRiq2oX5qFY
s6ySx/XpKFBl79/bmawb6fys9JgQzdrpXt84HBMO64BJdbrzLsiczSJS+O7xEb9UslEDxWVChKtT
3G1eVGFBc43FoDCB4xsmOEyJwlL5rnx/dkXfJV0eK0e10V5m4xnkQd4N6+N5eBPBc3n4HI8Ftx04
QORxdXyYkuiVorRbOThM142MlsSX7iOa43kK/dxyaSfyAMVCO/1HnMTN8MNVL2vhCIbmezaExPni
Qn0iWsjVUYt8GoOJToebcc+WwOgrTr4wMNcPGFjRjGV3OUGAPCX95EJ3v9FyuVwVbINP3Rp80rx3
WCtVR+YVxRO9C9/DkDgGTwkTDvu4dr4H1qb7bSYyjO+8jd7T8/rtvWL24tGLUnmOeNbfkhL4QYKF
ekTe9BVdfeAtpwj6M2tw0EqG9YwVxZ7cuiU7/wAhemfzCAoST+1Bbal7gcTyu9hqIVsMyUlqxp2E
2lKHvQTNaL+ktOIMjo5104mm/FKPEWHB+c6qHdZDxDPpLYg7oUeRRMRTtx5m447x8xfuBr6IT9Tp
Ct/ukSHssTYEq+ldNogpFFpu5x4T+8PqoSkueUu+ogT8lFtxrSROxMUijk2Vh5qywBPUOd4sQZ3P
MMgYH9MV4ENtCrvVXx2RwrbjKT3i05K1f92Re3ROzgjWMZZ624CB/ZwMary/cAH3m63NjSABUsfT
uCLGU39hesqMfMfW3vwRK4zbF4Ohy/3efJMacanYcPTYGGb1k9QhJzaIP6qroFWNhise898yqlws
YzcbeBcYP8t/g21110nuyy4dupbBfjUb6yJ2GcJ9GBp8kBhD/WniN7DD9wnOwtxHJaYQlbJwCiqe
xFEyog602kQ+rC+HWTebHjt1CONMYIBD+uhr1BV6g5Yy0LIf6uvrN8Gv8FHy2Q1gXTX3xWLuah1D
/Xa9jDPFt6KByXbfXtFVVcrkhyPzN3b2OhkUF8JHjdXQVB9Jhb3+FSJP3lhhtmduzPoh1FrF45eG
+jLXs/871WloqG2qv4sPp7CumsnQ4OgVJZmHFIF+E+Io12U3BAL+qZnvdIGdpLr3ancUkzE3TjV9
h+dAd/je6HdethzbKFhmxWheqCwPIXRhiU+g3HSAqSCGVsbwZoZeI1zjwb+OA4NJnFeQwE8DvCvj
JLDvv4kU7y4gDg2za3rbBdypOhMv5ALbMROMLjnpwY11EnXbiWQ7fRZEa6TrSUlz8lmoTgRZFvGj
MtFlctp7QifPdQtUTy4XMgTQz6P5v4vMn5uuM8ubYb1VgK0csqWBHhHfg479c5siam/sEdIitVC5
f8qsofUr1MvazZ6uZOQVsm+FgpFso2sM0BaUkwPNFfFm2RNU/mlqabZMRcDrlN8zwNFB+LD7+x1o
3Z1a5oagWNpRXZJ4QV8xxgltqm6VcI6aLeYwCbt3TZEltSzG7hOi16393ZhdcNLNbE6ReiiiFwGz
j6HHY78taCjo/qB8jtFoKISTapx94vDTLQCjdf62nPPrf48bmnlva0ySCYWOaIFCApUya2FN3QUS
QGhNabgqeI5qVWrMdGEJN3Vy8t64ZAyU+ec/YNnRxLC+e5roqr806bcawwzi4ei6yrOXvdEtFzgn
pO60pEgG/JS+e9fRc8xfE+v8C2kv90Tqi4wgA2Dt+tqgIKpyfbIAXCv8VRmCHZvai032fMabLc/t
FvYrH1yanXBTMhoUehA4nKJOeysxzwpiU/GEP4iMOmvO/Up8VM6bBkNngalS08jW1LZCdLZ+6psV
lAnx3ZPtyI3kecKoZBYICzPnfWt2XcFciQTe6tBtK8LQ/6M3R3fKfVKeriNvaLVedYZmnAbAfL1F
NBM0W7D/eyZTICy7Lvdj6MB+ozYW9VdyjskfXSCYaGsBNmRN1m6RBCpn8cZtMpvQ6gGOGY1BnRTE
ya6yx7gwu1aLvMY2r7P6gYVsCUVsxw9g01ht79VXTVRRRel4T1oNPb9oWl1UgjMWXL9G/7rcAihN
tzjk0wPfDHq2KqOixm1Lz8sdw+MNd/c7VXSHL8ZkTRW+M2SORd9obNSlXHd5SNcJImljFLJfOamU
AIs7KPqFe3nK+LJuGUmJUFfZTv7dH92xYXzAMMHxSA0uO/RZod3oTAzfTaI21SaOwJICVWdRrF5B
AUVdCCvFNB+ji7xm84t9k3Ffbb0APT9cCYtBjP48gzCH8YqPXWEyTDqVtqVSGxvkkiWYQpMgZAgt
zDafWJAHO2tYNSN/mA5/6ER7Y7thjLv3Lz+COj529rEKgjLGBZASWKYuVpRI2j6U5aqKpWmJC++i
SYcObwywREU4ZBiGZOXlY0ySClI63mzGtX2UTiezSCQb3yL9fN/q/hlh4rcSxxo8VyguVAPxdrr8
u2z6yZdUnB2nYJO9rksWvhj8DaYHVgurb7EjS05TC6UY/5awV7O2LD1rw4cEHMgvRtkvas4Z0cn7
JgyZev2SFTcN9cojqzJSizHJqq3ZZg6ENHKSN92tYvUcLmxjy2/+9ZAeKd1G2/L2rwk4g4KBEbji
7fBT7XaV/m1j/VGLHkOPmNcTBjVzz6ImDpTNohZi6d7zoGYwdrFidWzFOGka0BbzofrbO4rszbtU
ywsNsQfdzmfa4RIvLQlsjqVRjCZ0wVg37vHRl07J+OBaKV7LFvvIfMLpKODcm8fJRgmFel3crJ7M
lyDsENQYbZNBjyjH4k0kJ83mZB3zagNU0r2f6ddfXcfMh5W4Ep+xyKP9N3f/brQ+YRpiH9ZWbTEj
9xvNVZi3PsUYQloFmN+Tjt1BtCvLiOTRHHSzNRccy24nEmLaZutsgmJcGbTUoaS3dMEuTZqq6Nl5
aGVgmDVLTDdU6kErUtHJ41LAx66U2MxEAnYiDLJrnKgeGYzT64KjOSnYi4aBi+uQSjJcvUs3bf7Y
mOa9MJO7ExrfyJQAUkJYJYh3KyOjZ62HXFcwyfppmeKV7H4t4Or8bKSSfzITOXQOrE3urRWblhOV
4v1MjCkCfFha8uLlTSb2VXpAW3WSbxAYXcT09RUbI1YwgjZ+ctNmzDH0D3WTCBV73VJ4cPvxHfK+
t2j6PWJrGiCBJ3I2HeiQDxm8YW0CjD80jKaVshSZx1dhPXKu5ABsmOgFML1Y81uISkNwYHBVmbAv
QPRInQvD0mrqjkbo/j7EmHR/oFfl6TwOtus81AQ/NOb122SJ+JRKXqdgTmKnKUPPy/f+vTl3/ikW
T1pTBs29eB8NKPXojXH8Jn6Zd3f+1sj8gpUod8au1FzXcn37qKGZYqSDSkIwMIJy4XILoa2w3oC3
ZOfzmEiYeCy/tvCfWzPNQZhDbAtMMRibWelHdsdpjnKDbIM4HAQCwtAUq6xk23LcHTOrdlURgnAy
I0SCCePH/jUWzM9EMmN9wi6vUxMRY0m38fFIRCBAAd/pb7Q78KIjwi47AZVDaKe224BabMcBP4mb
ytxCpxdpP1cm9jd4yGIBJwzfQ1U0VJ4hJ1hlUn/yptJ/uSncfOoNblgMQEuXm1Qk4R2EXVufPKHH
OI5MwKvg0HvRWxc/dUQrDxKvKfSdPgnWg8fs4OUoAzN47y+RRT9ljTBPkvzEOEPv0zsZlDuT5Lr1
WH92hdoEYB+/+RjRZ11uIr7ZhR/M1v9nkd0GEK6PWOZCCU30W2aBnY2g4rpwmhtLdBE++c4AGHh8
JubR1bqcrGsNXQrcnLe8vzjyM6RmOCTNpdNsTjFFLNllp0bUGKqzpNkcYjUgzdeikizl4Ov+Ux2/
RL62lnEtesbI69+FFyJclIcABGg50iXmJi/tzhwU4a8Va15jpUqoj7v51ocLZ6gmXjVN7Dpz+a4F
a4Vlab/08hXnYW+nkJ5KnMZ1JKfHkYiGX8JPfRW4TQi+AfCuTr77yjZr0bYIvY9UerBVb9p/jKtr
z3az0ttkdV1Mcyf7RNdNm8ZvnkhMmVV5ilkWzxUzHhuOEcO4F+DovtCWUxT+PEIEUb1Wuf0BJ/yy
HgDQSyhNkf03kjVwKcrdQuE2S/Kfm7NsIFQutyhE5AYXMfMAiB2gtRh1n430PxJpkElPdjivR2eV
8URQyjDh9yrFbLGNGP4BPuyVbj1M8Tgq40cBfPSBz59ae5GFrdLxAbR2wEfdq/DUmPCBZTKPHJP2
V/2yGARNnWlOSFnazgQhygDaMyCqep0tFvUv7FqVMxMeJwnWjsy02j/I5mhVljya+NG1Nnb2S/LT
tox68ZjcqcgoG6SinE0l1XWbumamZrw+CBiNPiZO5LBH2WBfO4VXROQ7R7NLgZTBwd+W+mFtpIAU
QPGOslwx6dTqjg2yTPtu9reGy+zJf5Q6kGw95auFqwuFOEUrIfnOIOmZPptCIELEvEPd208fMM1e
MMXX4SfYmbzwI1Hy22OiQcflVSbsSI2JgUTe0fyKbq7D0Kg6Vv4FEottcl8uFtTcQaS+uC1d4nty
rOk3K1/IP7yxi58fbC4r5PiHIKbyNMqD1OVcN24TmI6wbjxOcpYf06K83u2d/ApHOH7pFqNxEJCl
8rG2le3ZwSuHmj0iW8zoDxhKxSnDwT8t1B27NoE9C7e+77XZMFGKrHsouOfP8h+jOMnja+o5cT89
2TmZJ9fWTeueRUHeJ5/vMDJInNWNHRAz5Ds5COlom7E+L6LB8J3Xf0ybpuPk3VA37KGxGPF7Y0N0
4JXzvrHl0Aht0fWg/ln+JpG4Ey26Mdwp1SzPC9wrFoDqMMz8+R0mdI5Aa/KjzRHddKqxTWsS3pJg
HAv8uwbrovginK1+QOjmMkBLKKivdL1dU/QuIMSAOnUeyomrT9FdknKqcupZ7wqyRw1mVP6hrCK7
9/aQcYzT4T9QzbU3IFwUiyu7hyVT2xlp6uB+iEFuAxRyXUE5SmrykWB5JKAdzomlCJBbiHCh7RuD
KXlyOlc3+KzZFrozeIO6cB97Baj2xYW6HumA/mduJFqL9aRvVhOZ2d8tKVidW4ABRvGBLXLZ/UcO
07Oh2s2YV0JSNPB3px+eQKeOubxQnh6ftTryzVUCMXcQlFfFEXi5C5R4zaFmY0Reu2qUaZSN9gdZ
Gu4R0UQVJZR6ai31R7EcoAP1dX9CcnblKAY50yoE73TAhBGjkVwjSWULsNqed3TImGQYD6XoT5v4
x/KH828CyFRZk4ZLFnP7weN28EocYfEUM9CEr3yC/uOPe2MdA0UEBX8RC23n1KQCB2Szuhc+c+2K
v1o0vFWg/VHdyJYrkM+8bkIKgI3nH+Z925hm3MPKyaIMMZnpJ942rxUw58jaFWpJytGXSdq1HIm/
eBQv+4jeER6m64ZyVWmlUMnSMiSZT/1ANTUqEsHSyaxt9jDB8/+AZTiqop6ArgtdWz4s2JEzWRxq
HfbLVHb2qIh7PJoQJ6TX/oKPotvFCf6jEqz2PsfpM7p/dSV7vj8++yUqjdaQMRJrqrlL+EPkTdxd
ABRCXi+hC221m/8Z6Yh7BGDaYrrYgLK3yUkIYx99sGEcDXMHHoVvKnYAetzO/SZr+t8YKThaLTHi
FIDqhHKUZJ20OM0zKXJrNuI7L7aQGt/KwitBLel0Kl76Z7DHiAlNqVod3/vuWAq1KjyrVoZnr6xQ
0X42MBsy+aHjxQMblYG8C7zYOMn7sbvaLL4A9aaItSNMc8mTLI8NZSiPW5vPiMCWTl5vfAjhkIvl
lEYBnxRG/gqvzlx39Zh5vCWv3euqHNUzJrbLgId0mRWHK/dBS6LgtFNE//5V2/MaVeTRy0fQEMQc
zknkPnFbAt2wzwPuoEsCxCP28rHinLSp8ik0RyMf0S5LQtSxWfoOMj7Kvu//SNNA9AKKqTmg1h8y
e935AnF0ND+ZA2E9uzxPrQCYCL7CHWdqb3oy4pUR0KR/ZJuwoYO7Kx2T7rKwYrsnS77czFOxLqXb
BpHVEldBD8slDMbwkw6Ft7kmoooP78jC4dpGuguMc0DoXLK9ym0C3nnHwEJkNYwwy5NHXZwURGLG
nhDQRxsK0kB+gjMx5ta07P7lOzcq5GLXQvpP23HM4wT+oR9xVBLaHDDb6cVdpTBk6BgINYTGUdie
apy6CHNUr4x0Q/pSdgvaVT1+/d2EFCFt/2hMsUDZhgvoupJa9nNaRjMDzEe8ShZ4LJpWxAd7ruds
WiExhCcb0WcazPWGCk2B1boT1iam4kA6/+lcoOJ8Jlf9uHwN6pQCQFkvx4Ff+8IR8WXLTr37i35O
rfR6f3leNO/ckeGYc5CxQtpXpitSZMC4NgDjoo6DxK8ACykOyt55HwySU7FUid0Th4fXtgXr5k1U
Sn8U8o4N8H3KqXkvunaREiJO9bFFrZLh6sHG6SYYk9dJuubN6cMVFSSCPtEXdZMlDwDgEaJe3wY1
jjJxxbJYqM1RHb2MH8LMrVRWWONtytTtCA7t6TS2MAQ9swjyz0XkroreX5D4gtkksPWJGlqvrRtS
NIAKGVHvqCROggyZrrNphnb73vjvWo/4KVnLtdrdOlAgKUbXk/M6R+laDaQavum6AbvicLT3EyUq
V9P1ILyVF+kz43zb0simEWT65FWBrBer9n/sgztOdNqxsFvcp3bW86zj4zbrcenkH43rbYl5mW3s
DGVBdVCi0Ue7nmI97rD8ZDiZKeZrAF0vE3jZ7fpEc87gatXi4pONO44iSIPFsVtjUJDOuXE+1nYt
nlBvQDyysFLj41rGyxznBMvCmC2VGfsU2CNQR8azBN7nxlvZa2+K9v0F0F0CGGmnHDF/3mLl1eIm
xx5PJBXzKP26ulFLOq/JADUp0UaHZdC7K1i2iYPwVTWdYHwqIWpLpPsn06qluufs6ePm+HL7stpI
C+a5LjxjZvC3n0ibPl8p9+C9ZiBvx942RNkrN8RBZHO6tEqlFf6hFVOqsT3KjJ4uFCueBhMv1HnT
PfTLUirPBca+mJIGTuzTz3labEzdEXnOAFNMyD6I2Go4a9NQMV18J98K1moH8kRd4fm5rdx4lSzg
BuaLxfk6VUQAA591AChtK3ViYPNhJ2WwzQGBPaaRO9IhVi/NQIPyLsBhgOZvf2r6YQNcNHDo0vdr
ByA5iGFfx3dQ+/pfnxt+FU/imzJYUhItL+0IsoQLxaxuKJKiGzOYgTWrXJ+P2dMvCs//QbbhdI9R
WoD8XEW5qZCePrwJmu7mzh+WbE3jUijLi/QAJ5Roevqp82ncYps0K6S8TyQLohM2wLAnoh7lO89m
N9ZZ32cXRZa1sAwhrk6lubCxgG/PCiBqBCPHkAzkwzQaBkGf0i7pX300DC8W9KUpXlzV52VdeIwj
bj3iuIqyBEe9eILNkVRBi6TQ/e5LqQvVpdw76UL2sfysFudf8O5fyVppOmjOImdSRvvuvaMLB5PN
2y6BElj7OFcMBDEuSsYQWSo2PIzseQZcNBgsNHi/LcSM/engnLE3VZJR8utYSifuoRC+0uJqLin9
jQ1z1rsjbq+GKRh0w0pVP8vct1sloe4PlkAch/RqMXqOU260HX/aUMzlScLEnpoYfs/+sjCWaYRN
f6Rxt6znRNNoRIugIPeXsY7LuJOvSsdYkc/lA4/EmtCQXK52zOVDBPGVu4VzQOmBlOHCMJNdq8AS
SlFGKrSdWOgb15rshnJuDk8tbbOroYafC0iXHKDTghMsW9IM66fxIN0aEtuUqA5dEYAx1UQysb5d
Kz6kMmf/56NDTi93Rs8uGBJxFJgWUQRCGjCNU+UG+LKtl4yjLktaVPOAvHM9m5/l26yDbXMG76zm
X1zXWBiuKrkIN9I8ElY4oCPeOqCAKUPHriOsnh6EqdZGzu9Hdmhim596Tn2sGDNRDUCW25CCi4EJ
zQw9ugVT+AsXC2UJXo/QpC78lAMc8I/pDMq2vO9eucLY0Ofp7I62tHA0iTHBIJkeHnkSS7mh7RCs
2PKsKgaGWPi8mun2LAmv+XRilaFl5slgduveE26RrIqPKanMTgaCZCupooY1BCrBEH478z0eA/Xk
rD5YsD93oUVdWxcANmAUgBDs1In2cjcuXyZT8imEaPnF6Auv/eFz1S0AnEQKDZrrHTAAdqjDMBmB
A8r7UrvDQSrjXjjYkTisYHCQdvS0wZyE/ZNIyrtxvTR+GlgiF2KkPPNW8L+KPB9Zba0iNsmalPna
K0mD5cmhgkdUUKVrzdbS8EYyS5j2REDXy8ghwYk42kQagz2wytJKdDEpX11JUa+FkFyEeArv36BU
YpUQWfiTagnfMNf0xshNKr/znZVAhc5XedjaOYZYu+dbZIRrMhjTWmOkT6bNkWgrjXc1l45DI3ti
JnRliS9zSapX0cy/n3FR6azIVpe7STHJj0wDcp5lLxNRI6BaPd/nlbmDhOgl326gSrbgdJqCHxUU
pZsA3+T5UIappt4EVJ8WCor8Y+K6MSYbQC+s3gr3K8MMrz3HVIgMgwIaY22IkAqIcQ9ydyqHUwWJ
e8eDETEB/7mB5NSmlXzcNPQhPVNKCttrVD2+/6z3XeicYNdn69c/nvHNtl9EMDEsJO0eTcqBgZ6q
k8XzWKkQyeAfg+fQsgurpP+CVpxBbb4738Q1PfcA47bS6lhuKkkqkBXXoW+uxXtwIcsfkA1ty6t0
MfUg6AYpt9Ivb670DgjW3gcYdZ+1p/hvWQdC4qUl4Rkd4o08MhSBdhowmfFHQIZH3+RIrVK7P/q/
+T21uaE1TJP3iiggXiMbayh/85v9F9Mt9f25oT0dw1JRPpyChyFm4SuCodLcdDUCh/ShZ/zmUHxy
ZSvbYWOpQRjfuFEHc8M1E9ksuoet83zp8ZBzh1ioMKLdtfuzvs37E9FPd5GVgtcdtM2w+o8e4qaW
ySyaIgdGHoC7gR/0xuTU+9AMjKEk6pyJRZjg3G5KctXYu97+fj+VDr9qAnznbjhtdhdkT0poOI0d
NogfbyKMHa/7+WaLsmefgtMRf2TTA1Ys0jR1LcQFe917Gd7fwwf3NvdhFcuO0DdWXq21aa1VWfUd
9n2VoHXbJ0yMKVXqELYLPF3tKbsadae+2UHQktJ4hD3PXZ59ZV67GyBT30QBHQ8oDs4yKzhYl25l
wu7bWq1Bo8dgF28eWK0JNxw674iI+jcyQk2qmZRRzzxFNSAdlcNwBfY2ryri9AhQyGDqjm4ErJGj
P85erchKxio9ZJzIqEpcWK1Ey1kz23FQvEy5zEJfaOkwyATSS7X1SNyuhnKj936HlYf85ZvbiByE
l4XwZUFjUyWSEGNF6KbxYspoUl5W1ZdG2wYkSkUOYEDMJyXuSjql4z8b0IfSBJIr44Kp37hMwigp
roS3n5UrReBZI314jBxUyoVsNU31HRHXCxpfc8xa6XSQryNSGXcI/1Yu4xji46A3iXJDGGLC14SG
bRShGb7n3I4/YsUrlK9L4M6hyw3zn1Zcg37Uu9VqaIoK5/9sRUUqa4riaFsjNp1bBErn1ReI3Ux/
QHtzCJEvcKyDRhRrC0bS06xtcbvD07IRmNd3gPccdp4iiEyZEKZliDnbcB1BNpRKWKFvT42BD/7Z
beQ1yrgDLpoUMl+CYazNLMam9PcVoPDVebxBPE3yewz62+p4Xa+wom11fbXS7PAgaHUEU4VSEGka
ynb1xW5BZyrm8FH9Pin1SgShKS4BQP7kKXyyso3aMQRgYv+TT7wYh2cdV/XNYxccfmy6Gtn7P6Nz
rW+qO3NImoQSB4wpw62OykUUjp2LNnOQGqdLCMFSu51EcEUfpTacpwoL2wT2DUpa/HOy/4o/sSLK
4h8nQEJr8/j+EkEhgg9DIvj8us8SWmGLC+se1/MzZ7d1PzxMbeYcuejgEB/kJBe5ney53xlTd3SX
6mkCK0nw4D4axfCEkFQeGLiyOUlND3vLYD126r+Xm5vFg4tyy8ecpDLGWd6lwSZjWWP2d5V8To0c
rn9gmAclGgi3qA+RxuFxbpMIz74igLH8O5pPMI19bM3XMrMOMWsdiLfcxfcxcly2OuVn0/pR/zds
A1r9wvewwv7Lp+IKufWNfueriSZZI/vFGYlY16/RNFxV9yG6vv+kKaQIUrYa5ysopNaDKf/d4bpm
1HmN3YDV0u7xiU6FdK3Uli5OllEtJ38RLrPRWZ+wLWjIbpX5OKeH0hifqABdyK8IR+XaRby+sPWv
H3qrRtd6J3q2u34pX43/ds9WemcPnKl7kh3Xtk705xrC+N69uEM9HHDg+/1bbpHBf02AiBkBgAJB
Wl3JoXMCtHoRFkBNvLP7OPKqUotWKnW/neM9lmbmM1rg20rn5hUc0YE6lZO5AgLINjx54ShuYqBr
yYePYjT0SbNroX03TvvAjPXEOT5/avgYlTnS0ihBNKJnYvqu6tLX5f+SuUCV8heVdlB5BFl+sYOZ
ie3eBeZv//i+dhRBxQVuc3pgVEd3GFU0H5JLuxfhNnCLR60mIikn4F24URfOCcdU2OH7uIaeGNhk
3WXHsnit8B5g0P7+BQyBojyHj5ce/L9LFs6EDgW2vyi8eIZSRV7XWhRK9Aqdk0nqS1sujwRmJxBv
XYJk/mT612VeVjfUo5xNaBb27gfi8oWbKQPQvrZHDXaNKbPo7s1nFCE+oUcVXTxVo6D81is1G7wP
eAhkRIbRPyfMAUgYbQz6oRqZjw4/cy9XzX1+onTgN09ZM2/iZOyYpuBy+x/Vm5vomFIJ9zwfGUpe
+th7BhzJJXPLsq/MCeFBkuGRpFG0x/3JbzWtSLxrbVPVz0vXI7iS1Fl0dNkriL1VknaiC1CVC2LH
ZSsKyZpEyLa1adZkY6nFKrknO2v1DBHB5m3RZUDhUS/ujfMHF+NzmPewFfRKcKHq+CC2lYke6epJ
5PwxrlDLTFgNnCwIIr6lfpq8IyMIdF6okouPFKSO60a9K+AZqp6BWs1JUmW9FMK8S9gRDBxSAfpL
WGCTCOiTSyNl9Pno+lpx+7JwwCNSuA5oxDasEhqrcDjZY1opBKkNRW60/1eX1KfCumxsak9DtuN+
eLSpIa6DtWoLBSqR1JPXagbGekoQ4+ivtYX5f3fFd5shC7Af4MUVOVYXtgLV2c6LLvls14ZWbxYD
ijjt2eWAi90r8/mkxFyC/NWalVeyb03Fk7tcwYl1bU7ywGNfZPMLY6PsJneuspV7YItIPnbHYlR3
C9gWENZFUTCQHZxZ+llPvTSxLXU92p2km3ezBJZQsrOdapu6qxif2iLEI3G+iKJg8mkGa4Mamq/x
RvIPgHGh2lzRPGRkdUvtOaJTvoAM5Fuj4GK3yWbuqGORY+axOJG0419JrvXZl9x0dN5kz+IIQEs1
ZkPdmWkBST/3h3ZdJWOxTShszxn9OzV8CnTX6X/+YVgLa9KwtKP4QDXHSumJ2fJhn7re8jZAEitk
Mx8p8eNDY4IONdevMqIc70zbkq30OAFNzIKZMq10ZbJ6C5Wo/7WZKv7eWFkUilFVR8Ob6aMCxoqH
ofd64B9h2nA8E0zZAC1yATn4hJBD/lhfNg/ml2hLM+pR/VsnqmkHE5w8OLAp7Hdz3RtC8RYX+lGm
Ip9eAXgEn3DRryMKbNX0oLHnRF7hQuVgBFdcGLY4cMPlznkHGejPpPxNSs+bFpxySEw9TkSjUg80
OjFmiOnqTsImkBCZT+uJz2SNUdKm4Cao99ev2GuPCDoRmDly5MJ2oVWM0Bt9TALU9nGHZdkUmIGd
382zl1lXx/OzkxF2YA1+hCFVXDtzttUceV4ZfytZ8NNw7DYe0y7wfuxW4Igy2eP0P/LrO5wDvs1N
b3f4YeGdy4EnC9MXgnD8YRUocLs18T6Kd7WfH65+zz89DA2LOdGylelNkh0IshNAgigka1Nqrl1N
+19PRA2ukFPt1CIf9UX5cdp/cVdIb09NbBJanY/WTzUtYcIznFkg8yr7/v+WV2PmuluTNfUeDV2Y
V0BEmDXfLmJNofmaZiE/h3y9oPSE9nSqKq2U+kS1FvJphjMG32CxW41od6yo/6wDofD8t3HJ16Lg
S4RWcGKp+XZd1tsklLNi9aEZOS0Y90JbxPV+D7OjSKM5j3H/KQPdT10Rimn7RSazLqBngPL5WVw2
y9VurOQCXLCZ9rwxvQEEEhPaiX4p0WnVF5G+TlTMbEpJHFQu9qedFbJ+AhaiE2Ly2E6L0ommRcDE
xg6FFO+q/dIgj9eB61Ob2RQ7Gt4IqfOXsbpUtSklt3cQjz6eDkOVHDz5VVHqepm8XYhaT6pB5ip/
6cAfVt81gpzYLnAmwU2tr9Te5nx6FuKi4eiDb93bx55yZQvzzjlZECmn+zV9qPbIxPoqXwMVQWFS
xKFdZzE0o/m3duOjNwn2JwJqMODtFcFAj5HNWAXc6jx6DzWmWBn4Cd9LFTMpttI9NjPdoVApi4s0
YrGgzeWgfAhQz5dlwWxTd3ggEtWQ1MWrHFBKlV6PHF3m0fR+/q7Na0TAB2rXrIiOJt8Z+Lo+pHrq
RrLf+iPM41HHPQ2dXwMVcbomyOKHVU3DrRsdPsVIPj964ZTMs3ZT3X4/PG8D90UsO6J9dxzODo07
GOQQUPzfQdA53PJrjey+CGiMROXFDE79z3v1AeC1SIv9vVVpD/APceJ9Is7A8KJ23ghuQMtOgSLz
mss2BJXOvAy1H9K1Yaa03oR9zEV2u4cbDdAV02r5EaKaSgLD43hecULC44P/+xBCp+MeEL2FT4Fu
2garqf68B03Y+84uStJdcaElxYfFkYgxFcazabIu+rq41uOb8UXJkidhSAzZsYmDzuAZVmlFlPFe
FRskVe8jMLZ+TC0O/oj2aFk+Cl2Fd+A1Jk5eF13AGkq5ioOHTyt0EFQ3CXKvvCmj0yLUGgUAyhF3
z7tjb7EGbPj82lXP2l3dCHDi381ah0wcBkTskegiMJfE1k+wH8h9a5i/q1YEkfFOUI8ATJ9AciFm
FI+JoL0zs/TPOE44VRJCx4TlRGZ0+VeFIRzMd3CTosWDV+/2fbiqwcpaGPcNy2Lmwzmtp2QPLU6G
C+MGVJ5YZdGB61Z2ks8Ikqf6QTOsddByd1dRh2O3EoQKkS99EdGqOLUyWF9kLsp8qYMtj3dlXAU+
B0+nxQJXHaHG6+3FB8gRfSVi128A/eneX74ZOTa7wfkTNFr/azNzcIZddqMqCL2a3Nr/v2WdD/kJ
UluTBXF/57zzdghifvLV8ArPGHsUkUTEsn2Dyk4jRG0TTNqY9yWpWGoAqXz+RFZHIvtttI++F16W
NwyqAxoHZWFxF4W+Y2hlx4YMebLBxh+flFOdv+0wJVU5AjR3YVJA86N6Nq4u4OEYg0HGSwPY1teT
zRO6tI2Gc0JpPw+w3SjvKIH+00US9CNBS6n26GunCbc4wbEMhDjz34WkAozvjp3Pv3j01f6ik/Oy
YdCMNFtutDJjoaIQaAKcNRBBOn6HkoMyxxliqI7zCR0grlr2SS22TNhEi0xmw6BVsiT0twjjoJL0
EjH62tf0PeNLJf32cvz5Gm9JHOr6ACVf6K5cIJNOAMVZ6Tpeo/XC4q9eqJj0crVUZwVaKBPmw9CA
KHCO6xS1ApaJubdj53gDCESvXNdKlc+/u0On26VPw7y3t9pIoCRxHPqVtfQtUHoZFqRnLti1AJRq
gvP6dG/e/yrzqLr6iGR1dTtveHFsllDpu9DoMnWpbp9/VoNRBeEQflIb6k3dZLEmjkQxHFpR5oGS
h08qeONJrhwlpO4bOwUr1qlIcSL3kMQnhmNtsB238rDtZDE4aTTAf6cWMAveI+4oG4/3T3b0mg4b
taIakeR8GSKdAJTZu54pksSmXlVNRHMiKI8noi9bUg1igwYYaaBpxgPr8sDQDtQDD31cTjHWOspA
KF3RnyjPlYFGuGVxrZKkaAeJLxGKDzNq2C2i4DLHVCacVXtQlizuoC34HQbAl3fqLIYkAsG69T26
yF7vbBvGU+0/OHWdvbhrXlLIXSKQxfWaJfme9K+apw29lgy9P7lL0P82uW0nsRlCdtTlGNpelLNh
jFar/brq937Y2Zw1mzANjkLMjdXLl07+KRa+lPiPpKqp53Tk1CLUQ6ksmE6yowCEq1XAE96DutCl
fI2B2KIq7DD2nb4h5mJIOLgR93Y7pIA7dlFK6uGJ7vKDi3kbe7CndxK8JlMG6ZlUtF1DyH0PIOV+
QFIWdmqlPEBQil6p4nLiZfIBzKsn/2uh+mVs8UAER8qqRiR7bGOl3qo23JdMb0wpSnYOnOktkUkm
CNUL4Oycnf8bHi+YLnSyuTxupcbLvnnZmcsj2MmYcgxd8oUrnnbelxrWRzOp1GY2eCND/fx7NmDa
nimOPBrjbW7ZSqpnM4biWAox0p+KXH7nKd1in/tw/0CV222crYn7ZfRllbqJ/goCp3yaIcPYNRe/
ANkZ1shUBnyyMC/N2OBybQrv6AOLAMHkYhGlX0IslcC5J6EMiXBa4fj7sMFDvxJHn7Jj6uK+r35R
2BrpA8/jdsd2MGRfE86ajGNKri+WiL9m1OdfVJHINiW3ol1j8/tH/XHfA4DzrHX7ehgoJGi5GcKm
e1DdBCZmRN5BfitVPjqmuSosBvcd1AUFWeAWB1Gr9PfNahYVYyVgvvRN7qzWx++pzTybjtAfeqQa
3+JK6S7HrQB8r/TnZpKyhhmFqwM2wgUbvfuRgPkM7o46dp3g5chjrdSCM9H0JAPg5Q1GF7vzynbz
XFkPgORq2q3FleN28tQAKm1zg37lLkkNrTQ6sYNhh51CCrssgzwZCEnexlMlf4kbqFBVL7HBQuR8
ZR0NOG5ZJXg646KSWcNyZ2VUplnlXQwV5mrzGPBzhZS1arHCjRQb8xczDH0TDw6umf4ot8hPACEM
md2iwHVJxfOBxsbpJ1fRaoHYikImdCx2gpiDyLNAhI8Cfnhcu215yQbTAuSJ7va5sEfXb+nwkMj5
CN8wNu4BQogCwBS9unl6dxXlW7fUTZcS2LnjSPJZij1kVhUJvQvJwwyqj6LJz7UdUYKgTJAqA/Ey
xHIrg3yaorfxdk3imMtZXkgm4ixTMhBFTD7IZ5stru+UYX38mfp77B7U4B9/uQrBk8D8kOiIaRIl
zgqg6ItAwLn4to4oOEkCDpPD0MjVSS2XrI/1GW9VEiF3cu2cOgm6pZxRBp7cUNtH7Cdf4SmsDUyP
/iRuoO56Mdx6X2kZSyK+w3E5ceWcFR3WEZmBEdaVOqEdBWJdln32KHDymCqEqIPH5r5a2Y9q+jFe
w1BTSHZSnzPvXdLc8rkCrZsyj8V7yKRSxwfwy3QctwpoyQknbAagplfs7MEh7jx2XcJVIpPFQWmh
pgiyS6lGUtUVoaNWvEGBYI26hiIDNjVsoaVb+2YUDv0EG4NJyuHzm8zvZ8WAEX76AT30KXSByiu7
BbXiRZPGw1K8qcD391+1LazS6odGcQuq58vjUm3hgC5Ayi3zgoSDoOFagPlrmLiZ11ADjxC4F7Qk
oV5opKcab0VDzNUTb4wLAQYXL32psrgIbHTyxVjSVuC75Ht8k6sYj/c+UfvEzQHXdiLwDVHMn1tp
uZYsvNzdHrtHcTD3SZepBPfpVxvQRqdLmt72IXUx+UH6Hg+LJ54/aMODks9sNVDb+mOS72ZjlfUu
wmYhcVxoMHFKIMa7EDcpra/sFmvsDtPeMY/1dv0gKqbOFj4VKndM7IzXPxn+uVlwcH5b0QDuRh9r
9C2aUi7zJGV0x0FRRQU8Lon9l0qmoS1q7f8nTtXExtWdGEmMuYv6l4JcyrBvkVFS+LGpVNtgtCix
Nrp0BSJLWlHGY4jDX0X3HIcavWCZVNUIFmp3IinFiN2Zkm7m0ZWiwwzcu54G+n7q/gS98OM7Tzv6
x//oHmUBllVufYHnVTjjNxyuIJK9vuOaj433c2QOwYvgEitdQkvUNc+1691b4lbTJ0OwOBfx6oGr
KMrtEHjingGEas+zGItp18zR3QKYzcvyXAZCn7bSd+1DegR7oW/7r7PuYHjbyrk+IFtTjC5a9ArG
pQiL59Bmrq3HAzaDDwHY2nQvWTMrHtnDLsz06ijkM5kVrFNKMefxr0YL9L77YgCFlVO3kZRV+Jxl
//wGpEj/uBIvTnzEXOzBqSUuklKKT6IKOxqhqas+cyR3Kw/hDhJy15GgGTuF9g64Jm+8JxEVyzuZ
s2AsoC4Gh8zQ/fie9ACgFHw8tZ9/aDl6J7xGGRfJUl5ZORwyTTkeKDzUhe0YNwAjdjIXbhDiSoIx
mQcomU5JdDFt2xi12ZA/Dc+0iee1hKkeFz4zXFeGh7jnbj5+mBNicfX+igCgLNsbD2Wxp7BT271A
98Y1eBD6nL7IvZJnBY4VT6ddJtbbcFGM4wd6qNt8EiaoNhKhbyUlXhf6qZw8PyC2DBVFjoGzYnOp
L1f9fsPaV44vklv9/Cf25JG4uEvuMv/Ny31sHwC/QGHaS/e4bzZXHlpwXTGvkFm663AH4cYbk+fD
gE44Ls665LFoZB0yC7OpWZZq/5BmU1abXgLoSxdnd1nkKsGq6+Z32H05PpKVsll/p3Rnqam2vtiT
VKObVJYdwtc88nDowhBpvCY0iLLe1vUAYB/m2nGYoXTfPzzE8fDIbp0EmwEJtH201tvKFtH5q9Xf
kgA25ujxO9z6uJZ0h86VESwGhediwZ2a04xgR3PI5ZblDG2bZdXZcwPob0hBVR54GwvihG/tY2Yq
rZcDxl9/U6R4rTa038QyD91PlC5o6/5Qo1UAdcXJGZHEax2zTQNvcb9sWS1yUcVtJOdQv2giAYDJ
Y/q9nmyAK5dhsF4LbEac0uh1QzQAUvH+jX/sj33o14HURVA/Uh3+GhaXx2jlUQaXCI46AB9uqSc5
Lpu6Ra0jt6YbP6JzqJWptZju1aIOm4ipVx6Ll7jNxQcHlHOwCWtG5dX/nDs5BXQY/WgBy95kdWjE
NqNZ1mBfPg37K7VyNsLdu2pj/udvsRXEFpA9Rj9ppKx6AMQt4r6YmuGiDQwwx21I44LAPziiSelD
crxG2/BgcplHhqk3SuE8oQVl+znnAbNKGmbiMmB8p/8PtpV2Zc8xK3m0guw5oZvVEsSV5C8eNTqg
jwKFgUl4tzE0SXK+b5nV75RTNXPbZvGbiqaisQHx4va/uN1ABBuJswqPkxBLkOcfiw7+HOvgCi3Z
BaMdjnEJLraRNhDWSx/doqiEEGcO59/QMinSRpQaRgoIqBVkyw+/irs3/x+/TuzwXM6EErj68cfC
kRv8YepZuxV7NS97141BLL0eyrDeUBAejxYIZeYzDsPpeVeEeIK60p+ygsCFsjCveKU/3dfuLW/K
scqmZfOgfE+6Yz51NSQN5gqy4kSn/4ZikJkASMEcpJA4mQwcYSudOtFyDPO0c5rX5PYkUH5C5A8C
nhd+UlZYUEZ9XterBlgdfU6UPZpN6SCGLMD7GQWHl3U/6N0gZDRkpqK+gKJnqW7+YXMjdvf5VjsO
XCPr0Efhuq1EBqlimBhtPB+tVz2V7nJcy3Chie+oNkvHpQPvyz97JJNJM32nl2AjcvP7Dh5ZRzxb
T3MDfCoiwFfNMTWfeWvcHCfeDBNfk5lIouDgiFkk1vsCu7CI1P/cOr0+SMDlJoSghjSx8PWJMibv
1skwOJpaqzu+RPeQTiSYsQj55oA4VtOIexXzd1VIa/54VdwOLEHa2347+nHoc2ZfT4KQk63apzlM
zCAiRwbvSCP8TFVMcPruEYp7XOADFrfTr99EG6EUJorueNyZhy/hBh2kBV/eebOaFFbYtf3ts0LS
xN30b6DlIyh11S691zHvqwAlcHw2WzSkmfelE0vw6AxweR7Coe6zjbwzfy58N35xk6ZlG0IUN9mY
/dtMNy79AYbURZU80ziX3cnc6y5jub+apIDvuNqjeyMJSxNQp4PsycFpR49WkYcyHB+j1889THfK
e0BGG34dNG/nwEGfOEjApOR8Fr0lPgTliTCNpefsnjK97TS+r+Xqiou/jSHroCoLSApzCFTpQA1i
uIuNN9B2EEsyom3pET7sMjEJzEhMv2VWMMQKy5hg69tGiJl4XNXGnf4FpZohjqz656hHaZDJFh5R
YvQbD+Qh7zyw9Z32CRD+0iccmTNnMUdGNBjtBTP7iPxmiryoId7GH7qx57vwg7Eg8SYmCifs5KPS
YPLMpI1C0BnCjA6UqymizLvig1LQeStt0z3PwmSXIcokwo96ncTYsofN7lo5/Hv2b7gEwfg9GyLR
bk0QKDliUIIpbeCoSmfovbo1/8uFNHMHdN78gcbNN87GRfJcjhXpt8kmn7IdBj4grHTTHrrj3ol3
w3getUwthwVBZvA7R2oMmOw4obobFoNqofG4R0QXlKTOjPoYWUti4v9TWdyPVQVCRsE/Btb9heFA
UTuzPXPoNJT7Qh80Jbw+1f1Zvx/G6ShfKqaw+QSgSGU+IF/W13ut69cbf+JJX0RRK8gvSoIL+Bot
X0w0z9gNOPuDXDj9cRBdLD3FFZqhSHGcvE+bPQawO34tvxIuP9sE38HUgDnI+orqm3LXGz2+PSjw
llC/8i4E4SSlO6M9EkBYJqZm+A8Ha4iBng/mJ8Mq45JPgaoV6u4A2GOi4p5as2Lzu1hzhTqhCRYv
Di2m3+/EIUoW5l6hLKbaoXpjpzDWU+PfE0tbtHBOz3PzC8DdMqbq/yZhi6K79aNdo4rSpw7n/DJI
+kp0wtlKgUHwvDQ1lccx4UKiQ019IR60661pe9znAgQFjNAY7l7aM5SHvmcpiJT7ZvCNfTr70j8i
hXPZVFSqNCrio0P7cYZhgna9R6a8sLyxX75sZfRKvlznCICzyg4dsTaHy0i84IqDqNjZ1A059Unz
JWFSywfj/eALvHv01dYR3iS1TpSIY+VoEMeOHBMBRS3flQK81hOdEQuDQDi7lhEWWZEVRvdMsZCt
WI6NPURpCtSL8YuNtbTi+G9KRi34KCjKELlz9VRRlfMab1MboX381lsjsSkwa2ta70N8CJ6f/oGT
ZzD+kr5se0cHrhQ6nGxa2XstMuzBQpWTjGYLMRrc560ZNj2SjUHjR+4/a1iievcAiWQO3Kpfg52K
kT72+s6SR9zXvqzBsz1TZ0y17W1uSKk2gfiOn4tQSJNE0h0YBjQcmWZ985Rci42lUiI5Qq7XClX2
DpIkHrz2j7hdIvADr9v5I557mtF0JqZh75GxVaz8j1Q2TkeDUstIL0iC6YkEDaMuRl7PP2cs0jwp
M5QcItXVAaV+IqGo3eOTccwHzYrNFQu1VOz23QaB19PTfOIWG2/HvPtNtD0Bh4midAN6db2FLagz
zukPEKvoikAQ1r5bBGOy68CX0vymDP/J9ndlgsmMMgyvzgmzBaxcPPnroDVb9IbNOlxdQLA+AnGe
LNPIA9To5GGYS/jedDH8CfSHJr1+QNr26xH6rhCcFJDuN2d8Tpk2JYqPhCi5jT7AK2p/H+K6cAB+
QalAA75JymCpM8BNSOAENOgPs1EoU1raqF+vYQ0714GC195HPO1F5QP3XPDYns8pB2bNiUPa7gfj
4EJXURybtfBgmG1hbTJATw63w5jLcb/RQrnrTkVONkSALyVxDp0Dul+XhQqF9ErSK1s8ssJd1w43
5crbk6XbRk2vjEaUuKMaWBfzA8aEdmNK3SIJbfsU4EOVey1XmDnLcBKUbSMN3QEIelxntaxCdDYI
DWhCYdsKDmciL0NQkTWbMQfLEYBWwt+SfLzGdvItAU6mNQDSLJR9pkoX1AM2B88Nonm7JpnWV5Td
YbhPHFT94Is2vRAWUd+jQ3rdny4TWrLuLJEFln0oYx3G8jYNir1ykszD8PTlXI3iVDxB5HPmjojj
qFvbizTWd5qULknz/fhZRe2NM8DPFLiTusg3czr3PIJwQCUq+pXc8KrGWPA8fZCMCILczMe+/jBQ
xXWlHIVIZUOiInIx3cXBuLYo7nSYnxNuASEbWBER/H5CQnasTKYnU52pMXH6yFfAS+3qZAcGT8bH
Tb7x4mJbXltO1Iin7nkk+wMwqP6js4UlxtHv/skjCGZDnQQmh/Q/zn9R0fCMXfIMgk1K3gwfelT7
wWd88d/2U3mHgJSdApxTDKwBDvlOv6YyH01EBipoj6pzIQfUyi2L7+C7cjWFM6dTsxGpdYVqsJJS
e8XDR5LFNHh1B0jRUO+LdXJmdbi2WMzBrCFp/gV+J3GbKolqC34LLipw4M9HESius/8RfPExltMl
ylR+DThSTJqX8xz6vS+a0qfP5/BQD09lj2jmQhjxcRWvakFi28rTDp2oBLDSUCxCFoepB8gdo8Jm
ntBbLcaP85Uwfkf9l0h9riECnIkVCAvUkSGC6L1AtIY6b4/Prck1xPmflNVhBP/7P9P6JQSSEh0H
7oL08he0o111jonDEyWgN5UveJYmo2eQ03z65hunHGs9VrJ3Rb5UCYZjHXgo1LhrmcQDCOPHPe/8
V0vcoloPhSwDvZp0vJTOaWti1ea5vBS6aNjYk4YAufeW6uW9btw27tUoUa4u/ld9YSOw2iFOrCrC
SH4nqAYBAsf23xi9pwfSNA5WeZwAZXg46FK4j5SMr7YDpaa3hDch+FBNg1zJqKHsUiQFTgA6K7wW
P845HWrTrOtK6OLBBiwqmk8XmmXvL1RmWncoo6rUSkfOyW79ubnPMZZK4qYn59nu3EbkMCtSwNW1
NuzOxXrEer3M6B4bw3DYjsxlyfJAhxKKPAZZ88QGC6ICs7oyu6fFSTaBm4BVhwCFR6ns06vDIQXf
uKkBzwCUrFLjsw8DLkCkhxMaLvo/ZALFAnTliVrlv/UPWUc5MosLAer2s/D059khkeC3xd8Md5dw
6+K+mB9WS3x03tL7dl5igs2j2DgKvQazqC1r+u0pwTknsH490LGPbHZ2eXibiCc/6dhPYsVRTcQl
hKCcR/X6f4qSPSirzP3hcTm8ibqRhJFC9bv5EPFyp5++jxwHYd4qMeqZUd1caLucUpp1qBzobUsV
rUYJz41+YZDcrKHcnuAIL8A4m+MNDD/or148GsaJoaYtgz9FfLwGABX+MwbH2gzQ+YlWhATuuMXI
qvbqaAs+ZqElZMKhNr6lbT89P3hWmVx/KwrA1MuZrsLTgHXX2IlBDSOh1AoZQd6QK2wnN0CNJZji
u19Lkwwyc0sWOiaBgywsZsVcigBavqv6hslAjO3CzdP5ktAQDLG1U0I6ztXRe9I7lNJ+CHSo+HaV
/3nhZnWuo9QoQcJLy3xI5ZzkyxL8XIjCxqaUSC7ov00l4QuR0bgZsafeg3mui41xe+CNWZw1VN4A
Dwn/umjJgwIqVIft6N1IfS96DFnCGPSWrv6gEIdvGRC62naaQzmu5ckd5icwW1X+hgm0TPHDfb4a
u7WTdZnWmBtE+td1RZ/Jluwteeg39+CZdqN23K1L4QWVD4FPK9B8zl+iLqEMYRlShLC7Z1nrba2g
FtCJSGQAyI9JMtiIkLBzDwFjaEyRnuCWg8OI15F4iCWzUtOFltAMlvS9wFAvu0hWxBdooVpJUpyZ
4bVgHBNnigsKiN1rAYVpjkm4nwPmM64vaUKMROBDGi+1sD6CSkY3jQPlsLy+YeSTaCk5FnDHtEQD
CpR3FQqPoplpkXX7dV949NhqQEsdm1CHL+S10MEZG7oD7bsZPIZHRBcxJ5KnV8ZxmzBKcUrkiFn0
4ij2E0c6h74cckYS/qIWloQ2OS90wBgC6NTDUTcp04zsvnsJvY5Ucxgn+cQWisNN0r5dnJR6v+pV
o+NUYY4sk0fNazOPO4tce8OblKOtE0+zZUIC3v7SaI31Fb68c4M07h2OqBAlZhlZyE1B+3m0ftXl
txBRQJli1YOZTRU25PEdaTufn21tchkoz8+FTXWfLwpj6KSstOM0oZTYWPl13N4u8O1xD7fRf5JU
ZX8y+93FzkG3cpvg8lVc+LbJDaHj+XAb6qMYNcLRlFWyu4VSMqeB+YMgJ0n+am6a93dBn2r9agY4
OkAsonbkwPAaPZHlPQ+wfyoWVjPQ+9qccRSio2C3Gu6Prxaw6euuk6v3nT0mdPuXujE+52b4VvIl
H6Hk3QycGs7H+Xp9taDYPVwZffDR4K3LZAx1h7+tbtYZsMBMCkjyV/pgAVDl/N1UW45C4o5cbVey
wtIWpWe/WHkEvnl9eCd3QUUM2QHNNdWITPWCfcIHNKsrMDTZgRf65Xtww3wHFeKJ+SlU3pZmQutZ
Dvd3S43rSCgibazGan2zh+HTN9StjRr3Uzke78H9WuEx3c/26VL6vPwGm5lXDTqVYgvCY9nGT3s+
LLsjSKfcFy+xZF3RjyhgxZ5G9RW1H0A/w39nZrq+Wce55St1QTrJQWdBCd8WwBVmifvxGhn8GtKV
a6xmbE9S1xJhfoOIBk/WUgg23u3aNoNd2rU2bNJNDv+0M9G1K67LodvNgHVspUtdRcStu5DNWLqu
o0EAR3HPPoh/rufDU1YHdUBYXJIjcT6ofG2Ftmk9i5Vo7JGZMVP/1XkGEv9OIZ/CvxKcM0G+W6My
BYp4LZWOsZDo1OZy/p1n6w1mqAeLqOh6eODw9/yovHen4RlnR/Pyr3XsLaStRb/eSnaJRV1n76qz
AUpvlv4wiwsSe2aBd54RLofRVyJ59+eHrI5IijSpD7ZN0uqEY7BO3XaYkiQQlJbrszgw1yfBsGaJ
gRgtaUVFIf1gsRZxn4UEjV/ZfmeSK+e+a5vNz1lNOsnizfcwmCHR/u5x3uqDGAcuriIduJcu0nbX
UpEI1sFhsmNzopRSuTUb8fizU4I3xiouUTIlI+ArLbh5Ne81JGJA5MODnm5bmW3/4DL8aOjO5oPB
8ZSaLNCUX6ROkJdt5CMaaBQjgTMfGZeoGklJJ6lRVi5gUpUrI9QlzUga84PXoLOcSPX8ODy158HM
FO+ABqcIgGZc/+8wm7qCpU6gl9DYzgJcY5WdOzWWmOrnaj4NJlU9NM0zVjx6bhiykzyXri6va+H6
3J/QDgZQ6z9VchXsaPl6npzlvCIukVlmqHk8g8x0wFcUMyLUbOAL0TlT5ZbPcweXuLr47cTVM/r1
W6yj7U+xd2Yo8xDJueDQaEAvA0a9nza1Nu+dTK7h21bi+MyxeTumEip8h0AMj1zSv2b/w2d0yU2z
0rabda1ztm1X5GraFvV6AJpFvCKwud3/TfRaA1b+cZuZxfxorSzRymWXj1M5rbswu+UljrNvkSXr
Bbb/Sub/YC7IepliTCLiJXkpMxi/45atyFQgY0LJZQ1S6RS0NufHrpuHeJ5pQPNcp7RSBb52SHvh
Ezuulc0lLFiIi4pzkvZBewpv0v1tOQ7XNu17PgL3Lo6o1Nc83a9v1fasdSYb0rbWk2BuSvz6TUhi
bCgusvwuJP4gUdYeIogEz4fg6W1mCEbssfKW/WWXcoJS90ixqLKUiCbmOLEYJTRATcmW58/Mh6P9
pEWEkcjmNf4iHXQwlyJnRhlnA0CIywV/a0V5NZj+fBk64bkpTUnHMwwHYn7gh8k1ITeZuNdGe0Sw
Ew+dFLxSEKilPiLW+EREeR6ZoLjLLbAFDCNDJCtCbAwqDl1N3pRxkaig4Gv0nu5wem8ZuNbHYS/r
Qki6ZGLnMt3gq6Hrf0qNXfUcUgnNiYxM1zZ+EBNWGTyDsDSmyxgQB4TX9/PmhqNnpyuD6me78yXf
SpVEIZm7HcfrJufGdpZC1R5IJ7tG7CA9DLcXKvvx7I7bmGHumo+x+/JOV53Xnc2kE/VwseThXmxx
IWp1LuzGhr7xu0W5znlsnyZz7StUlpok4ct1jsSFpfRg9MqrBxGy6Se3APfuIiqZohG9BnjHlS1J
Rcv0bEMZwdReiP+0eJOKdoD8ydN+LgWLVsJpevai65K6Yc9ewDn6moP5o+ExzcHggT27/5dr2MTm
VjcbqhChPUlnytA/y6MGMXjb05CYkMAL8YMgzesnCKFilAFdfTS6Q/IGf8MWpTdnDgP81PZkFRym
qE0ikDXVmErVvKDsOqEckdEiLfyL6EEp7Ux1/BdmBamRbi33eX8r6C0PvzOHtc1yE9j//skfDl1L
z02yQQJwwnQSd6leExnKnKl8zfM0ITVJ22S1nsfeolzULCq3h7VgO9gIDyRr194TdV+0kNyAqa/6
4s5dp6ZgM+3RplCK3P+JktTVxI4lKORKc4cweeBMnLONwLnOthOHxHC5/KC2Zkb/tr9fVB7586wQ
YdBu9XQLwSsS2pKrNsWoRDWNShg0gwA+PGRRirgx7N8lNqA3iVki7oHdfrDaebEtMB1W4I83sd/Y
OqsdzcErG/ChfTnqafCIEZhQm2ZUYIwDq0UWkrcLdtnDTjv3ng12bqLpwLA52AmIvaGeupYXP28d
tdCtvkH0ZGq8/yVKBfgkAmlhQd3cGIDd3JK1xgZ2dRmkLG5fwHMaEE04ej4r3o41eI2/k4nytngD
wklDWLmSaTodDaJKjiJyBaH/meZo1Cgy5SzZrN6N967CX+vQ1/c4LpjW/lFyaWqMwAULC0fyUDDm
p9oP3GjpR8YpIyUtUn2CBKkqMzkKS3zDuuShME7AIuTnW+RXe5ozLL0TTIoFBQi/bZEQyvXEPuFD
r8xn1KHOpZaXm4lmYDIExxag/o2xLwICjRMa0xAC04TVLmEW4IMGD6FbfL3/+XeYfl7uTX2Uolk1
LUnqjhGRoMkac185PgoKIRp7dRTn7rTlB/PdubBKYIChOJuGHhSDS1IypuFyItEkWpvvht9KUlvF
Ud+bh5q+MERLqXxJXQxeCkwK3kCwC88BTbf++9Ao430/CsJVoIkQIB8GQ9cJsxvETiRToO32yeOH
q8sZK9vh0Y6ErW7oJXJZ7EPuuwKuvtUXPodcekNcK/4IapNYXpfv8dbMmEjEgJPXx6CnDK1To9yX
xXFkQAsX+5vntBGigvLgzRMr7WdaqOZya1sC/lTTyAIyncW49j2/djSJKoOoBgk8T/S73DVYJhZ4
6N5wygJwBB1+MscwROuIRLGqI8R6sIPdTHynejVuXcTfsgeqkwwk96ETwNCAT0ROBa7cLj2FnT23
JNdVgPr2XIVZkmh5chMIKc0bB1g6HxGzXfXiLw7CRTu0fj5vsO+hRpudTVk+HSp3Xxpfv4whJK76
8EwOMDCIuHIMOXFvOwgyzOEde94fd1sJM6cZW8oGzEwlIdJUatI+bTyxc3N4g5qEigvh5XK0uM8C
La63E+j5RMAejMsV/KBOJhNUdLffCBOnuVyM0sUg8Gt5TA944QklrW9oEmd72XSbo9OOstqfjSdV
hfcwuUDdnL88321OKLj1bP7VdbhZmnnEZvoHY6CBWjJO2Epec3VdoPMt7rY6pcMgZECInBpDLvzF
wuScZ7/g3J33EnvvOntbkPebuUESOBfBwRDaNfuS6dp4ZOd7b98WmYTjh8ZfMd1bJDg+bbeiY4nt
S5xrLu7/KIHE1NPmlNwslnz3yKXI1hXApNFknJhXh5YMGefwjK1BeORiknhsL3sECSwfBfVnP0I2
CgyIcCnAgd34yETVP/MKm6z8gjTqWCLWJN5gVRnhdTqN9StT8LL8apy01+b0PncQavywMWSPklb0
3sFa+l1LhC/zSppJtlCXoZx/dQ4LS8jYBEobj3XoN4i6kNloqlPTYK/smt1mHYCQ/LZuTNmAlzt5
hT/tVACZ64K37LmybOIhy4VPVycqxueXfjueMy8VH8hDQlZIJDI7zPkqhvGXbjrXGQDsSexssRKJ
MTNuOOVDFPj7TQPWxCyV+Fe+tdd+jBdAI1/u13bx2Nvy0b7/yZNptW4IVUgUKCzzs58LxL475B5h
vuyotH9a0L4YEO0/6WTPtKkWUD9Uq0bMIYPaTo4CYc8Nwmo9xvagCKBTe7Y9Q4hcZbrgfhVE9JTN
SM9+MmA/3LCbXUXW6hb0Stt1fc+V1LA7BcRXLFGUCU8AfY3wgt3DS5iUJ3XGB7qr8t0koCbPUG7U
clGOepPwnx+6XMRFCorZRm5xFT10wFm4hNsWG2WYLzWKKZOm00AcDC+wc1qMVqT/xOB1lfwpOcCY
IbqAcij1kYydlPoS7YcCZRVDBOKdxQFlBZdU1lYG2vyeJkuCHlPGaa5NDkjQxxjOf8FrG6YWNfqG
4bFzgdVZbjHICDcdCuR33ocICiEyJEBG5DflJebAS5nl5hiSBOSfm2CEc/mseUhpjhoGOJTQkEBR
GG5WKxlUa488jksrZZ9ydielSHRov8YdBw5+GKoMAPeBJaseHYSAjiYLgRALVYlS2v8DkUjnUDl1
HMjvG+//Za5PwYhGbOA34Avxmb7k5Nrjgwe/SnbL0dnaxrjue1ocBEKI0R9t9iExPGBVizVrdGcy
CRuGuozZA3Jwn2fQ2MzsdeRtsleryiW9QWNHG5/0O6SUAC+R2O5PUFN8qlBEhF2m+poqONrGq+pe
XzhRbK5JI+Q3BeE3IPNjv5hcirQkXQhH4b8zum/AHgdboPPnRfxvvGIsgdRzCLy5au1Yf/Yx68Sy
CliB1JJVZVnaAZ2ez5zcDfV2J3900HmbUHdsFbUy4etq26m871kpHdhbn7a3AFyNxDqPyJbK5GyJ
SVUIINaA3OxJR71c3DK7qfvzfR6AaG0/pesIxKeXNwiA/y2PlMgRjfAebSnMiPjaTobc9J5YPuGK
31CaRzup+SzytS36JPquR8jZZSe8KxjWqNNYUKW9fhRrBF7BgiRaNSBqqc+UnNlmADArfnazOhFm
iJ/QMejwsDgX3yWWclvPiWLv/5Y+KLrL6mdghaGlS2x5FW/s0Rjr+oYETefXVlglxYqdMHgRMgRp
YBxSVN408w1bV+dWSq8m9pLk+/1EdZ337TCJMVVy+XdYUvvKsvMKZOUFkGkrr56ChaP4UHul6RaM
1TxTrVMCOEflSyZlpM6Cbh/0feISDvmrqB7nULw3kgBG/0skSS53s6bIOZVLZ0uYq4D72VagXDIL
NLLEEkeWiXiIre9/Pf1TNU5wN1ddhWms+zb+JJucBXC+q7TsHkWP0WueRwXPTd0BRK4QKn4OsKgM
hChHqtBcz0FM79OIEWI1yHHbIHgL+ocRdOpxIu4yv/5mE8zekGyKLsM3AYCN5CfGXhj/zknoOq5B
oVM/vdETbkGrsGi2weXh6yiONhSxIKTxovaUstkEEKpYMJ3k5zW7cSTo0wCep0sb5VKmOIICLkHr
WaQO/G6x/VXH2QoS6ara0Iuw4QmDvihvD5elRcNMQBPPaxR7pVJPe1I3PR9IZ7LRI5aRGW1jwcIE
U/72CYc9GywZGHm2xdjtmxaliYSmlLfxLPqssLFA4A8SgxbAHtbB+wwH4FjQoU3zz4h+0nbiZNUC
sjaVT3vmGUm0WJekptQpl2Epj8m8Nfs7iO2ku+b0eZ5V+WZ1ZCbd+RcFBiAAMxuVVAKKIOWpcxDf
2Ld2385A1vcR/ciHsu2/26mY65IUq6Wu1n6u9JgMW4kZsBdqWLjwU/BZCGQlXUM/qnPkUT2SfEOQ
392Uy97Dl5gjBcQ0ZQMX6v9UAraZcRu93NeCpQYq7BmgeAfubkrk7YPftsDrab0MioH3Q6lyiuBc
xorYVR4eDKoBkq3GlZ/igyRvsn0aZV9oIRhiPuzjcZSsabEq+fnJNiyZlHXEE7VrgDKUkD1ohi0c
1P03GTi+lZG3XeiueVCpMBx/IPAbvZVBcWbSwI0zUy3QHLgnPyoYakG4LEPrN+/WgigseNqFZdzU
Tr+jqWzzIxkPNxcDfnuM7qtYtxrwsb5DdJGD/2KHbg6aU/ks+lU8lvKLGUe2lyQR6a9PWwOSV63e
dAPnMpVdKCs0kryGAtb5JG+yRyB7Eni1CGlzjXymXfkJuf7rI7StQ68Tc3UDTOa50lroodyCE5Ft
0S+f9LKUa4+xFdH+9EPnbhwaSYbHQshxOG/iOU7mqw6GyscuPb+KwUEOkjhpPl9yj/SyT63BS/Nx
Y/qFIipgy3b6OWYb0zFn7ucqpwIG0LI5KLA9KNagyt+IT3xLMN0BTk4ekbMw+nw53n6yBtAl9KSh
HBohuqg2+IQE3ke+BhovOB52W4v/Ya8bNmFNyEcWm46MCaqXg+uOpaOwU9dKwdjAouITGjBavbhj
VWlXb9sgBXfSibeuj1nBH84TBGIjKRi+1G05UJs3M3n5zMQ4R2Jhe5xJ7iwobrcmGtP1c67tNh7m
aM5+O4FzEu6i2KNWbj0sPoJuBF+qMCcRVUFm9XWT/r/TFLRl15coQf7BPvgRQjKJj43fKlnHpPcP
OsazZvP+kyNh9PZUywCZ/BdCQw+dY8xl1VfnCsnLGA2KST4V5MonziCKQQvYraL8VsyEhI3yHIq+
QmY0x56XOH4k6SW+B6R+9Q0c6k7WcBdRbsORD+0IZWsQgwjFVYgWdBubx4wANpKP82IReh8P9aBv
OTBGqtykpcERjUs1GrULoyPv1Xq9xhuRVJ/ObRu4NTbYcbMw2EEBXFjYFqp+7JMyvcYg01qcakxD
5gewqIdrpC0jG4frZ2Kiusbxctqo+AR99ujem/IuEvM5vbZAUb/jIqN3PrhtM+CsCZSmfkwNPpmi
99O+K/6yHq/Jne6oap+KIBe+mbVWWxoIW89XHJH7ZG3hvctsjL8ayf+w6x/ZpSAbQ8HJGY3QPXcB
UXf7dmss6FtK7cTiLlbXlSJJR0bWddR3LYNeppA1FjR3L5wW/IiHXid6/QknP1rNnkHHuCG0UdMS
Zp/FnVbSaQnI8kEq3/kbukpkEf1wf2sF1AwKh8KAj1m3eoF1vZlCTj1ZY7TNu24gkAt86CCC4XBR
3ZE7WZbWVwE+eZgV8u1x2oQPCGpf+oeNqyy7trA45lqG5/ZCPFo9hZjNN4AhPbq/c/AL48qrbzTg
QZKP4FN+O1mbsxTO+mVEbC4c+rCvDZErCSp4Xycm6UmdVhu3vxvlQzgR/9wQFpJIL9DiJKmobTon
6bV2l0vHBa8WS0r+6AV41kIH8f0fo6DPN+czgdD0dhVZE8ohpzgR/w+HdQpquI8jYOf0c4alZaxO
7YHuv1Cr6FC2OTBG3eUg1b2qBUHqS3Jn6OSpb8NkvbNATbyUbFDax1A35DZCgXBTAqt471YUdN3q
1Jue87lzcEwldgG5yv4iXoYvBSnr/TYifXlB5W+RBM4XOD0hUL4UwWXTn0YHFHQJBrUM51ulYL37
mcC7HVQdO8eIZBDVkGacZk2bsqXBbzYAALQqbt+HbnsLUvMvg66Sw69sednyGYy287DvcK9AJaFf
S2qCsu9MpJSStZ/IU96KeTCY+X45pk2kEz5mGenaU3j/N1rTdBzgtKJiWD+H72fGNY713Z1kAqGg
FdpusGGV06NN2j3heguwfHbaOKv57c90xvZkbPXbk77T7aOtxsv6tB6nB53vwhqoArGYu5vtYS+Z
SetqNubhUYv3Jgke85mXTXTS8NaNiG8BgdHT1A/x8z1VCHlOA2+v29zznQFFDH+l0FW+h7WYMabj
/BbUl/L8cESOD1b0NUiN1gHUISxXnNKP4n4O55hJZrHn/BaRETxnX7aJAa2hiDKH6M7rVFw/zxdE
ABQmA1yKxIuO2ESscc8AzktfdMhBeLldMuC50UJcaPYJf87bNORyrsGTgiKNn0XrSuacgxVhvsFz
ca3/J5pYAQWM3oV1CzxhGtXn8JjkFBMCKZMKacp4C5/PcXjHxHBmNIuwzGm0ViQSJmNhgHjYm3ND
IxiFncbshdqz2llyrcpVC3UQ6yVM6RNvVg2T6Is/cRq68iSm9zL/nPY+3yS9TgjwLQbw0GLQStLy
RhGKAJYgn0ospznPUK85D2FcwRBZRnQbc9e/KVLEDWwiDF1sKNIotcyh/T9PCovAc2kWiqGJ+17C
m1gM1hktlGHMtCONx7aEftuCRaYcSxwX3aI5jFENuyamGe9scSavOEQuREosooXGmJKDLDdh0gqC
ZOlP8H2BpUixlNBPHJnFOCYLexsySYEwQYscGAoRkMSMHiEI8czgfM+UMzlhLvFeK53RHSWjrkLw
2sRCfXY1JI8gCvX/ekHpR2vONIC57VCa7gTDPdIG3/2zIr67a48dsbKTrSC91bToUu0um4Li2ssD
S+/1XmYqSL5OUpcVUNzWpfn+oyOCYKWCPyFb1vK6pcYnSDyirAqW5JQDsYweABZ1ASWu3R2tBHxP
2S1GPMp08gnZizsBeYdQM2yPb0Qu8soj4AjghXPB2kGVwrCKvsQcICjcqp6GM6NttckF3oM6pDrG
D+kWQXMGGU0WHNvTVJVE4YZFNZ9+LQQCVKtRp1D8JrCBJCa893Z9t77wqW+rkUKZ+refMHpXxEVi
wZdxyqomP5SlHhk1CuhfA9e5ADlhYrwGFJhqq223gqk9LUJxbJF9Uq5y8jMQR+rYWlBtUJ+jo04Q
9GHQDz+tNwTYrZQPEG3xqtWKdin6+k9A4ZFJ13Tx99KxPWNc/mP+LihuYLbNdHKKgfos7kp0vmwB
YlkvH7T2/8b1CaUMKzBITc4Id6JKK7QcSLbI/sH6AUpLn0fQgQ9aOueYlxLAJ+X70by/FdiK6Ik3
qDz2tsSc7UvF8AFvU/Nrh4b3dKnb6wK4ujQ0qddc31TTix2t8Z23zAB4CRQJnmd9Zwb9UehXU3QB
iA2HVktv6DIq+Yz5Jicz7I5LYZ4eJ5F2h3eKNrWEaK7MKmRMs3ZlVAgRzIGAzzsKS/u3h6KuOvwE
16KwzrHf9sWpf12kYY5V0wS1Mfb0cfGMrt7j+UVWK2DpqinDEknfYEQQ74jcuTVPeVvwUCgB3NiJ
76H3l8SdOK+Wffj2qq8qV1t7S7xwiY2E1+SrVbxlGgNsQiaUgBtyLl2g+ZrjEf2znPt/T8ekzWKM
ND/2nPgV+gnZ7BSCXTiZXcV+jGrR/2M79c6szaMoAAy+F/tslrSB/LxDmWkL5zI5BZpQ2Uem4cKw
GdmhJ5jWay5KcnQgv1DW8W5DYOtoiZJn4GAPUN7vmyPdurjdNnM5ARXtp4utuweTRXnc82DQIBAn
Dl88U62cFyA6wSibcG4id6WFwffwSpbUS2yVthZtwXgpT5DYZUBY9OTlwZszFe/30VAXrKwizI4D
vXr1yCIOmBX5+bG16/OCUa7ckbuWQFs5ptepd5Z2HiBEW4F9YHWgAJXmGruZMQCIeGaxR7p81oFc
wFd4hPKVnx0o2mBAYBZYEh0pAUQfX71+PbRpmJHM8Oe70mXK6LBGY590crLfwzxOC0pYnTrHnOsE
2NdCtwdIViKihdYsPKGGHgQ89gCKeJBWjfuLCnfuioDzGczsgvNXrR0WpXWx/5ACKzotALR4TwYk
jZdX4viyFrXa/VP2SKuL8SS5wczIvC3UIwM6dYVJZJUxgi3cEeUbB9YyjbfDR5mZXffkZYvvOVc9
EG3TDlSKdDSlX5yGU9EWn+0XH1Vg69J+zeNUe9mAI36I6XyS45ZEqa4fWSN66MXfE1laYkwgd2UP
qmE4IYjz+GinSlV+rtuFlff6tg3Wzq7QjOQRFc5WbxI0ZLcfp7jxbP3YceGfKYxIFhrcr7rEl917
YtzVUlpEiu9KEOVNU+tk4EZmJAqIfhlueB5iL2kvOALTJ1H/xWnQ2zdBQBcKW1bx65eC6qLo/uik
NDAzPKSInsZgLTDCTMdAmCHkHTNkrr86ePOw4pBAiAy8CU28t9ELp2ObfOay2xinVb18UPkOaPL6
7CeKEXYVJXvH2E38a/lK8zeWab3IDqfiJ09nyAEuMpfkzvGlIxJTsp8u30rAhfwTDAlhcZdWkoZr
HKT2MkYWkY2ZRL+8gwW8gUI/yIyKkaP/KH7e19gYrxQkU+6buMlMPCq7zeBULbL1BekRjVD552Md
c1y/VWc7BuTlV5QD7yhXesYkgRkZ3DTbynP2lm/RjPh3TgIGgU044wgTKEM84Jw93dc9JO7R2QqI
b9RKx0kb183NRO2JyUBFMO2gSIOkAn+wT7XQiuKhky+dSeMjyFBweuUYrE5U8ZL9xoy9IcBMaFo9
YSQpNtXtg/gZqDPOl2IKSxWt6coCNr7Wr5SAxo6YAQAdMtthSSOSpA+EWQasc2rQu4ZCScl9+qXP
AY8QH1t9cH6cKtqZSZLUtlgDYhFIn2X/2vcg62vKUfaSDXDNF4uYxOoRzPP/ty7VE28X5/3rTrMj
LYlI/LflwgLgGlZxlRi06USTAqAWYBerCRowHOr4OH6Eup10idAzAAW8NyRoDkCvRU3feAYx6ssO
5bEoL15FK2Za1EDizcy8L9Vr45S+oPkXCUFyAXC702PiwzZEILSzO74dCdgPEQ3EdaKfgT3Qb30G
J+0F6u+Pr+tmtpPlIrEtZbtqBqPJkmgKFxDF64aqp5Ca0MA9+6G/xdDKivmE8K3xGpbeXjvy7C/4
FHVQ9m3PbMNkx+M+dEGdiYTeElWAvYhB/e1zA/KTL8U0WuJ7kr/1Q2YjoKfs58GT9QghTaEhvezH
LXkRUi3O71qdZFIMMv3BiF50Ww8DrDdR4W6mD/D0rTkDX7uB31D5akjj0UpiLrYWuBX2FL7jXwLD
6uq75/wwAjjtZbVHgMngNOaOGjE1WM0UwdKhoDzBgE+i2q8rX4duPuZArcNMqER8OkH6uoNsEb2l
VZutysW9DD8NhikwR8Dnj9KDrGmp2ShvLgUv4ntSAh9DLxY2j/al3rYya4lgg+Ne64/8efyFdi4m
WoGUTA7SeJAxnP5TE7S+Bl4YgNgEt1HzuNBpGBVgW0l+F+CtzPH8wytaC7ff03pLzDDzCIP/4Uj6
E2hIJjk71ceH+8u5rAaBRoFKoja9SVuykWe2nV7n+JbKYhWgn72ikNUfib2mSr71TRv36Y9tou1O
iTD4GzKTbCsmwI23C7iL6pkrZzJ3tS5NXh8csv1RQ1GuekgJuXDAqKVRBCjAM+A08Fw/MDbJxaKN
q0ZDw+70KT0rBsSiaI+MtiUn2Rj/R0ne6U1zZMMRXmPOtE56XnbjSnaea+gxyT/z91fA3lnNUJ7v
yIytK5DRQRHd7FRjXm5VAZSEXogvyXlAIvLE5BrdoadVIFCbQBc60Xc91RruVg9dUkVq0OcjBeJt
YoOb0f54wbc/OaI+zg8rogJEEUe3mO070wx2LRFvcYYLrOehDNbEWpNJcGN9DJ5j1iLGxgGNUQoT
r3kpcuNPbFp/x4zoZ3s2zAkbZA5kveA/mgXyAk9978cxke0SA6K/3heoq1v1oy/bRg28FxpY2qqm
T8Mhqactz3zhZfbLpn9D+xVJG4ZapUZelvEEd17nlYDRXGxvwejwPqVM3LFr1hmq/DxJKtLSGGJf
STMQt0IU8F7rZ6YlqJv0qSbSg5PCs/UE+Fb7ujm+WUgbi82ckaZq2OoV7SBgZl1+c1xjeFt/v2zB
vTZpjPDMopoVHQJaLAGGffq0oMtsqgjFS5HMysnfLv/3oNV8j18LxXpq1ukYjev9Hlr7jwZF3Knc
T4zltbJBI8kQ8Ez4PUKOQmO8IzQXm+4GAp1JX2iQHewhLDEKeK3/mIHbugXkEiEASPnflE2mLepH
7CZ53MWRgl5/SVl545LBYUteReTi3RNSOY8uSez945oX74rKYBs9aOqiMqqyYlFHe01iHvF+sdB4
hLtTO02glt1HRsQkfDCWitlT9npqYSLEjNpJyUhCELINb7R+d6cJ2c3HUsdS+QjvyTzho3e2P/mq
Dq8XPknpZpwNTqpTx1So2k4e9B61vTz/LkOCDIyrlem7Ljz0Ic2YpkCZ8u8eqB1tIHdhYicByGYH
agiKBCmGxd6hAwxHzAyK4K8y09kBWsDhEbtDjjJTWJc0UQXsMSjjUyNSGwI71lLil0sptpvc3s6F
+4eewCHa7uPoprqzHuJHhakGuwZQc2hYJ5lOfnu5KlFCfhmO8esJBDYXfnFlraFH6x7EI5+Sh2jP
akznrmZdcKAcGaK9z5+H2XChIAfS4Kfg3Jepv2GYLvv1eYRMARl1C1ASaeD27EwboGC7MkOnuzp/
ALYEFEPJ52YLhHL28KPOj6r+zhG8gI/1wKEz5KCdnT1YtG36acFYYyhY5JuaPl6RfI3HSFjm9r3Q
WbV34xHsQMSWNlC2E3X74En2J4KW2NIC9MJ1DaxwW2yEJx/8/zpslbLXwEhCDFXn6eoZSUXfi5K+
UgNGJ63POKMs/3q0PJZIsV+3OVnB4BGZDoxZfzAJ26jB098qyZyngLgQ1gT56IQxmz3WbzIwhxuF
V8qT7S6d4COIEx9J/mtGo3qPv5crunbqA4dzVGX5toa8dxJmaHz85mB8w1NnZvRpEgLKJaTX2NX5
wX8NkUWiCZcEUlOjSfH9xFcHxBofjgsfa8oP60G5bC2DgjCfoQ4BsDJP34f6NoC6k/aLPk+5b6Ev
bkCjXo+4ebtKWKRSMow5AjeWXLt0gT3wp3z+kCElrTg+eQssem3hTS+gn6TaUVUk6ZQ7dZnUbLSs
d8L3+3Z+H9uK/5+ZWid5TVQNj+iA2roBU7heSTmvfhYPA+hq4+DjDAfz3bFqfmSSEr4HrltLL2fA
jrHV02nhPRAj75QMaP8356x2XQPBc+syT39zJiv6/EKNWEyi0kQ7XTM6lyQaj+w8129MA9djteG2
wPzmELZzPeMljHEvDq2UuPaAjG+ul/U28OV2g60gUiM1IIjfrmVpLb7Z0/etOMbrupVFS4eQ4nCO
eSu7nv5dSd3BvN8S+tjCxfoc83HPtwAXQls3TjZz0lsyisU/4mu5PGBzkpM0Ex8SVxFNbfDOK8dQ
JQgQZYlaJLvv7+uMqFbErLCdVdXOCBlpQPvOgr6tadBUUCBJkNX3mhpbQTPckl3GyBMy3K/Bqc7K
OmMl3P0ryY2Y96Wy5VEX5KeAhgSlmZ50G+epLmw7tKo1q00vXYqJ5CLXNrkhuh1W0RDaUZe/4Kn8
ZpszbE7YYcsI6Ld8yjCi9CQTNBSRPa9hyNOhYLtfyKegHZtjnyx5ZYfI8bSU5mjIvvvKA5cJ48rO
WLqeOyWorf0NqvUW6zWLYsPzQ7+kOecFBhdMf0xKG6q0BahU9mI+QQ7YspxhcUkSEupMFy4ggtmv
aK9Uj1kV3NfVQNLIlEyi9vhIrsZkyjORUVoZ1ru9rln41WxUDFBvgxjpWoRFJNntB0iR17V7+B3L
/YiuP+AE6AxP9PPg2RoCgPbrR+EDP3DDZp7Zyv/iUAhd9TtG03asEdFdh+b4Y/8m3B8IoDPN5liN
+CCbgypDBe7z3zrWhNPUcsVFnpg0oc0JTwZoWzTX5HROQs0QBiQXN1Ua9TrpZUpnJAi6UZNlZhAv
omuuJeSYD8gtqXG3TnUnpM3a1t4e5sh2M5AuTTxcn+fc8VR+akCgVQRUou6l4FYTzF7PqmwbSNDK
+v9BQUe5KvscPXXQcX36TRDjvyYRLkJCYg4GjUYzRxn90T48jZDX9ZO0qhq9eJWWK/0R8ov1iOOA
lEJuLrJt+ZZAPd75OsLu/gkO+zRPdSd3K5OEpu5UeJ8p/3oHTjSOxluT4yj0eUXSOd9uj4faMGGS
3cqlS/QZi5bNkIwGMNBfDENCq/FmBbucQTLy3yGmUWdh5hbF9S7gUHU4gD8qXrBuM0gdvNPXdsU7
sAHnusprsgg7NCNg3vFOXwVqZgptu03QR7BEw8SsNGGI2fyTb7Rjrq8NCHG7Iz9kE4amDLRZqcaz
wnJisuLzEKZo50CoWbUDlPfayjmJvoecHC1MOpBYg/ZX6wqwuEBVG2sBXrb/G98Z3AnZSjfGGpzp
bIdvAx65DkSPOvVsa7KjlhHd9oTn33Ma27vVFi8V9LoFKb8RGdnTbjjxnpjAURV4EwLwI/gC61EM
MvWd60WgZom0NA5FMXVu3azt57KhcXSucJmTt3FyPkw+iQMN/RlnMNcpKOiw7q10neyP8ixqHku4
OR7pr5x8G/j/ZeRgyKaSym9WrGLAJ+TAaKyUTOjItX3ySoPT/WP/2Awo19Usrb/DAf9Y2NVMyIR8
Y11QStYOMlZqzDolv0KWcjkBKDusy2n8vtgwn86vjEanXB/E2btFKf8uZZFzeTIn80CO/xlnldS5
mtU6zBZg9jBdbaaGqNyDjBy9hmyL5G77vnNk1UAE6b0010YMwV1p+P5/T1+8F6LglLBsvLUMkRex
dBU6OjILCtMf8u64gBjwS/7rEcaPSe9PfQU/8N4TE/2J5ZFc7zqPWEiJofZi3JXudPoCKFlRvonL
F/450ZQKRKl8D9AopSBPXEKBI82e5YpFydfQWDAdfibbRMEEpXjUWXvQ/ISy32qJ5rJ8mvZtzknW
7CbQjYgazndPSO7tWMAstpKML6yVIbCftQIdlVpW7mkBP5SdS0yxi64o5+e7CfIourmn9Q7orp1d
IJRg+hYGxhupX2ZPyUDNZRvVrbFFm4bOXAD5WQQdrx+CaFD8H8nW8/Wa2JuX28ZRa6X8Hhr2QAAL
3zgRGeB2R49245U9DHGMLCJuqXW8FHNqT5K6S1669b5/K9s9Ki4iw8GZdMRdnqjt+WIBXsfMq8ll
ODxHpgtSJVC+fz4Zv/CTCDo/zUdvNaw0opPIVonIB3ev7BvfWCxBQagx6nzS1kcHUkaXWB0i9qeC
XH1EINlrbbbdDrSU13ngp7ZpYa4rMRW/+p6HJj0FwsvjbQjOZvc4BVwuFuDqgsfNk4Cauql/GN1N
tCvEyR8AlU4gxiMJLUAbCwgsREL+m5QG0uLSil6eQXU0VnMwsdoOFSFcgiDesBjkWIfCxmIA+6Xh
3IqiUFEKjvazexR5u99Q0fBhzJxcXRjVYBY+KhkpsiImeqtskrv/RndnRzknNO2bj1IRq8TJIFfm
y8U9vnw+Mby8rmPZBtCv+3HZiojvnYgoiH2QIz+dEdhRqEBvdAOT2KH+3erCD/oKjFUfU0bWI+Mv
i4twDnWSEHIbSyyyMGnwSc4P/3X+7zXn3/Eb7JgJL0STsj7ErJYDkX3ycu4BB1/JGP7gqD6Zg9gM
5FlSxv8+/YbJ9xrSsFztPQ6D325OzdV6Ke/IjHPLvTtLvQ+zBiuPkfTDZjcanN7xJKB5o1Bhm0s4
8T2AIt28PTUIqlQX7uabKU6v1oO/t3GAWBmEl3SSZczUgEbHuXPioJrJed8gMXYKkcmU5aUHvvp6
tp70yjgh2iKgsuupPpsagv42WvZX3HIcTEIQmXIcPByLmItiMCuIuJbHRkYusftXF6i0o7neI4ku
kmfM6yR+cr7/+mu4M1JkNhvSKQCNXcMUCEIO0dYmCC54v8QB5K9CzdzhMr8EpzOmaaocdnLLiKUE
Zhrfbc8OSDWo71xX4emaAaPUV2Y4kYHtg4M9b2QBVhDsq2ot/u0zP0A7Q6hOb/XNH0NYr7Jjpn0m
pef/JtvndQ9YqPmE+sXV0t3lbxmDQZpTJJYplPB2XaYdO7tW1y0/NRQTRt22pBTGLDkOAsc0XK7d
8+zJ8x3AbBx8K2+mbBOPkGHM3nsdasqXZaSOCpaZXZesJ+Al26LT01v4cwERCGDAO7RBkS+WtfTn
KMvwFpIHl4275yzeQW302fToXJ/nSLQTDYkD5i6U9Y6T4mYowyIYjRxHxp7hf858fAyHdnhQL15+
d00n8TrPWehI3NXqDiftHxrgD/oOhigvW5bgUUhlwGGWqCZSxii9fClORVJ8zHk7kLbm/GTM3Lu9
2Qtj7jyIi8rNY0ivpH2P6KIT0Bs2TYS3r8pG8YFChbTdu5gaOYzybXlLeY8z+qwbEtgaipsfMnbZ
86m2igk58ivnoEvlWwRwQ5Dni3utvLmQeWTvvAcEVfxZEOm6q6yDPluAzuGqyX8usz2+cdrhbCoW
lRdHYE5fJeWIAUaDiIbCanGQgEAhCPTXY3OKcslLlFM1IFqgyfYGdZ3LOJrYh35l0vGFLP2W6lIv
W05siz07CU5kINsUlJSx7+ZwlgXuv52M7N8rs92+cVNz9Le9dXFBXHcv/qEBiVqFxoG6DV47mLkh
N+5sMSVO+vZj/Rjc04K84f+cXVYLVsmhj0IElPSipYH6WcAp2P4H90Q1hR9/7cyxsb3l3pYe2W2F
j1eovIrZOHPvRN9dUxiZD8PWeD46HlJ52/l0EIDC850PbDcwoeGDdaKzZeuiojwNhWjqf/8sLSb3
yLNPAcxMk6B+fxqhXYADW5FmJZLgg6Uu+K7rm9x988FuPuT++TtfeDsQGvA31v7+8/wbmJ0V14cA
QBzexUfleJRx0gAjBUMPndXz+ooEo8nl5wngQgyus9HBK4LTwLj3T1x34vf0x2aKFYh4LmqTnEDU
y8DbhSemqrH6ogsJZn74VN3YhqqsBzx0bDwhg2YCN5KLwz7ZmRgHXA4Y833cEXNy/ohhaSD9+uC+
x1ujMq/gaRKBnK4JTNH3ggrPxnN+oC4ThaiANYesqThgAQm5c9OU3FD7+slTTiSkN/6bS8MLoTuq
rtUi4+ft9PRq9NZW6TapvHAbBpWdRFKifvQSLpXyqSghHQJ8tsk97CaMTBzJBTomKLh4ON0En8EB
C0kj10GwdqZ6HL24ojvXbEqorUZ888x0kM2Tj+fdxzu+CKLVaiF7179cqpul4DZHQYf4mRhQBpvO
j22UDmXz9XMfWxGlwaQM2G0Wa2gs0O0u+8OT26U6SvHJxkRV+x1kEWFTg2e+X+7E1Zg+aZ9OkMhg
f7jB+aOE66MO2wDTD2q8fHJPIMYjOvPhqNR9pI5JpQRZ2zQVA2CutW8xpGwg4bP050oRgjCOX/Sc
cmPoSPugtQkv6Yi9nwYOJx55zTssRLwkN6iCwS3sqZ7wMxW+xIQRMfrAjCeHII/GDGD91SL+XuLi
G/O6PDrC6ke+73u8NORou5etsDDrc8WQvkUfKjurMPV8CR5r9T4Jl8I3pEFXz5WFZF2UnXQq4tN9
YKIN4WX2hJgE6YZWxvroFk5jfpWZQhQANzpCR4CZk7ymVGHpJhCT48IN7DowjUAWpCmrF9WB0TYv
FudHpiFOiy671Kk6uQT0DTZ4u8pUWhwrqdwnaYZISYh52BIPOrESc8hHUoSyHkBzqKHydrPSWb5f
37BGhxFSC94bpvEhTf+Rqg1EkGF6KhhNcpMB8CHBvHiSpdeRk+76SSC5nJ2X2N6NtUpVQFtdJWLV
I50qhFqNOF9svGSVu47tx+j4NDyTK7JsHC2OuMXBw4N/t4OP8ZjQ5H8AUhQi16hUsSOx5jv9jxVe
Z0QRW/3h9gs1PiQ70tCHp4iSuhuEPczo9n/GzbQerdLrIEQdXo+lxmBPVuWFZq5W/cyuI7ptIj2K
0uD+xhRzDeT6xRg0mFeh/Hfm+a1l5lr9bIspnY+0bbaS5Ennua6N6GqSL7OiZO7LRgQoCcOy/tBc
24viJYYbHSbH4zqO+0uPWjqdyysYkRd4Ux3vyEHzN+5nSCR+T2TAhgutRWLY99OflUzjbNFUYcVo
K6J9Em6OpXNAwV7FbMyFTTWqQVEdm4J3rpJmJ8D4d+k4VWssoiQiQk05MBUK3ZD8yYt4ISLC/Vox
xweACZPPsGBxbIOPsqpYjMVwN1XuT9SHgvvZ2wOcZN1ifVN6/tvMFxpLGON/STzHvptQIh+XinKu
0cJqGv7QeQNrtimI3zX1lUYw++b9cn9mPD72WkObPQyavazeh61oMfRNiUOLfmvmPMvAoDjCMjWw
+o6cd1+i6ecRAKOk0qlTkBBxIY86a1y8bn2n+p0cHDkPcDPg/TMYBDZkx7vHD1T/JUDi/dBzUHF1
7Qsk3q4ArdimOaZHsheok6kGtjkgIyeYeIOwMCu5Nvw0O5hgIbNxeLIH8Nk8KidT2TUkKxxPEAqW
4IhUVFBl+Bh7Q74Qf2F8Bxk0o/rii8MrmIhlqJCCLKcqP9+L5ycN5lcV3FnAgkrPVG914gH84Hmp
UFuQ8/iPtynnS8f0SgQenIe8GBMLJmBaSrec/fvzTTlKbyZqQybP6Yt1D4PLHkFnIYfUZa80UQE0
hqrN0wm/mkvxwRu/yA/vNCMoUIm5nBbzo6TlskEeotltpnvDE4sfoPB3R56PNQm9vVMmRu3DQGKn
Br3qwgLd29uh6EyqBykqDxmUuP9jIo3lQH7nyx/isQb8v29659752qdRYq9CzTYGdhk8kaUj7bL+
jbNOq+8t44QMfVWiosZ8tHoFrNatZq/TouUgxz0mbq0YyQhBhlKQ5VcR6aBFoOmrPloqAAZtYZwO
Wqae5JA7uUxHuMjafLoeJK0esZ96EX7lkIJb3oL7cp5YLlrKdS919RmFkbH2Q2B8XRLHC9ghBGU5
U4D6+KFf/wi2tspclNAWmqHzI/dfCIQAxQAfBLcC8z3ABfyUNnrWl8XGlDTbGVBQzV5WIpuSvzCQ
/3EreHbjSIg/2HCyq6jlqKvZYQiJZhRrmLYBAryL8paujaXpAKm57DGcVZNMwOm8FOVaOMN8paoC
sGrGfA+0RuA6zq3A0nMleJkyr8aJjbvZwtu2zqookNbLN7l5Qfc2Ok7rPW+PjlDtKpWSPr+LEqff
7ZFnkYZLytUIbY3kubGjYkrZpz7f62+VI6T/ivD09/z11fqOLnaKPA4dVwip+dhMd8ote95tI0qs
5A7NGz3hy7KBcPzS6QWGKY7ktBkTgH6X005b++pHFyfnoEzNvP5DVqZ4o+0bVuBzfypNFhWWV6+3
sXnXASsgShRVcU0mxlT8nDcbr2M85BspnLEuJFGC/cnzCQYJ3rXK3TCMw+BPIJG2rHTVq4/Py6Cs
HPFmsdVZS/3aOj7cCZuMb7btH5k9a9yLCQjlxlDNgJnVr1rDtaS/hpGO9ENcy8SSYZ087FUzO42Y
1ORks0EpDA4sVOGtIuFwo0KhvQbuh2gK5/T0Y5gguHCD+c6Y1WB9/zSAJaB0wMlB8lAWxmwiHmz9
Y+uACUxbf2qkdc3SFiZmjYhjVR9vXZ6sZn5M4/jVJ0Gnp+axaWomK4l8Z/KlJrzPLgHs8TdHIrAY
D8a+zcdU2IOuxi/4HuAWnZLoygxmrA/fNjRmG8ObAwacuSJ+ZAIkMYvRJSDQcWT79XT+Quww7EUv
17XX5Y8N9Rsx+MDQWSNvDgdlpsiVOyPwqzg8BdOQuxd1hWimtSfgLGaRqVe2r9JLujjjTdZ9UwQ2
wgNIQ3pakNx28GAEqAEN7dPZwZn5S8gK/1ayXsoQAGn8b+vlY58HtkfI32hgaaGVqYHvDDnk1ntB
nfkIcXorNBaAcC+2UuP5JAP70xnYtJvoMEnd32ubX8aY6eMY9GSbEeXgEgw8MsZu1qOeLhQXjGGL
yP05uwFyZjBCNGLnErgc4fTYa/VR9XQ6gpdjx2h4hMPwNktJFlg0fJMNSCTlDqr/hgzEPTT1ns8U
FUTIn4eXAqY9cInSrvLDEZWF4pxI7RYpV2RqloIkVMY7PzaAyf1GNi3AnJqaKRqhyY0g84ur6xvm
vO+GNQjn667UpIHbptvXQyrkBHDcSncfyYKvUkxBGM3ZwSJ57N5wXyqN5ctF7I7DcefYegVulPax
yv1NiRPiMIT5ZUbftsbWGx5NFxJObE8z9jO0+u/BFSqEuKVodpS/oBQIoeXHUWM2/WofOLd840GE
ouxbe1AnE1bRyZPPcFQBq75KfoFgiGgjXEFqMu5eluZpjC2iktQid90YdWsBh9gEJFKFo38aaK0a
oCpgYq3wwjKqnpF/J4SOgkslhqebr1L9T6iwYVZbO8+q6PJLR5bxXn8C/I/auaL2S73HNhKtAUrt
hx94LKsoaIpbWmgnRzc1+cFVdtP2AOabU58OH1tZ2PdkiCgyytB3n9ng4g8pOHw3A8TIulKHy3HF
+HRjyLpSHVmG5kF3bmSgPIo225V3boiEDF9/Zs0a09oj8u4SmE/k7AmAoeLjJD9w39DDZs2ONzp3
0xviIyR1Y4bUMNwoxaDEU0CSgswNkFkOAwO42WphbqlMLcxjT3d9pl/ks/Pguf+zxNu4w0FMiTrX
MwWIf4rhETTv/K9+kt+PjnrfoMTpm8J7z+EPaJuAstqTuo31wV6Ub/gr15xL1p3LQ4GGrUQppisG
XlrSwk2cwVHnPW2gQ4FRZp0SGhDvbtIJKjY6ylBaZQvYcmb3wlRf8++FEL9nDHltmbt4eRSIe/9w
ZthmNKOdHfzN+Ih2NsQYYruYp1rwSNd+Ky6W0Syvg29KuvONFWT5jzdgI4PqutXlnUeGGn9NTARM
gyFkiidnCs53CSsiqh67pGILZ2/nexFapQ2MZjME8+EvEB3kdS+rbwVIgRsIqbuReWV/LBnyoV2P
H3kDooo10hu+VDOUWbM+TNMEvx68wKgtq30LJj34bLDHbBig/0iYcv9Y0LmiORKzljoo24BDBfQe
OaSuu/lW3m7+8s0TtCoE1iPy6L3aCC+ddqUEMeTvbTQUHicZXr1118JRyHRLSwawTpUExGihtCpy
c7Y4AhAVMwWPj6rlSlgFIofdYo9oOnBRBZABe/KIJGzxY0ghlpY+vwWfPbUEcMC2KyaTl+BP41h4
DLS6dNWRsoUsZc9+UK9k/3IGrKHUDcY8zOjMAP8iVbCWpw+yDi6J3tb/2XeVSwJNDyitDjPo/Ire
67MWBz+e0zCHXm3+rSEHr3bTqfJqzvFsgz9BWBT9AUHE47O9Da30nU/7FKhlAs7TZQBAEjyf/y+Z
TuKNE+Bw6RTvoVykuwxSvXOUI0C1v3B1ck/GDjjOzwjhW3q6uRX+nn1w3kuG7W1IL1o8oghpMbWh
+AS37DwBdEZ5EKFfaTbbXCEdHVIuWDu7LeG6hIHh1Js2ZEq7Dd62dapvNkFc0W2FWN0rv9UNPVL2
KVwUa/ZGCHPkqdPBuUkcJW5eHbD0ltddZQxbdQcKxzYVULDlEmhIKqYoSVa0LX7gfuPCehHbu//D
SA/JqLihrJaADNNQ7b61lyrCgK4eI/nlbNM0ZeImUhMmjwK+381ULjj/2jseML+Ik2VM8wk0dTqY
ifURlFSlc/sEF4nvCIF0mJg0RaY32KPiYWLvL5d+ckZyYbtemuqeckBtKIiE7qshkB2S7181EJJx
xyNbflJOutxZnk6gr2v9bBR0jwriwUz+Zhz0PutkQedqd8HOC+noNHVfhxEfbwKXFmvqWMUA2LRw
VKiMu3SZXoZMGbB69+7zRow0xsB2AszkuaS1WprjAhfIPRowdv6LuLR/7E5RbusVqvaO3JZEzt3h
x544RPD2k59ssFVEmyVVcSEd+HkEez+DWHqDzEchgslROWSs59LAdoEs3sZdo8rlrfZO5bVm1jet
3HrhkvH5c6rzH79XR2ORQ9tm+4H7pjUGOzMeCQh9C3vqEbqptLwsEnq/Aj2QkQqWHmZ+Lv2PNxc4
K4aCKRDqOPHZp8icPVjeGoKX9VMmXL1ZtS5Vu5WYe6EL3gii9aOpIQ5J7yukhzQwneM9Q7UWV7yM
eWYBJvk6eHuhFPdJKpnzGcacVQ3Y/0jojcCpCUvtoVcups/E7yFVDIqkOXZSkemPhQEtOaItRrE5
8MTqHFQZNlu1Koai+DYGUNnYQ1xtbv29DWZvUN5uPF0UOu6VUzb6WxcK+rG3oVPXmoDTDcE8dA5g
M1IPiWpDtUYZE+HqoVubivkuqPk1st8JeE0BSO7JBw3c6tSjmZMaZeLxTUxkrR4h5CHeG5HQm5rG
ddXklPG/hWD7GhuOPLCiZ4TttG1Kjp1MUvPblZOutuPT7n9Heci+43r0cC2Rw9A8A7M1XpZPIt2N
75A7ZCS1ltCuZfiSOqyU14/fW3SmLFbg5tXBueGkrihwAlLlReivOkVSYyw6g2p02V3VQWhlVYn8
V+9/wY3jiXh0ZbTlOL5U8BMXiLg5expfQ3hneojXxw4mT/ruqrOCJUM2jYA38LRjkFGf7I+/JpQY
pZdE374+UGb7KuDGyppd78w3lP10N25UITMuL2tZUVYf0y4+pfYexUW32Ij4WUonNVirLNKfpePM
8fAq3MjQ7qrvPc+NzdrRCknqlfhV/fNx21P+cfhjruh9tkSzy5qeCewXNuGp/g53vErBakKYTnxe
h21Tw3pNi8nrLBNbQVnkiD5UH2rLA6oY1tp37+YElwSO3hyHOs3rjppFo1DngYmbT+mUDvfJYwm4
SIlcb/4vHsNZha7jlMTEMd/n/PJ8zEnhQQH6JRGNeuWaSCHh/LWPoL3SKPRYxiU+tltk9a+OX7DQ
UZn6obGTneRN8Xb6h+cA1nmFFUTuH173Po7vg17iNNJ2J7D7lEswNyZkdWvDe8zwu17cavZH9/v0
eB8emogtrosrSGMoyhkaQFUsoxUVmLqGulb7+NYbTwrz2CUQHzRs6voBSgk6H7ViV1KCbc3Fv7Bk
HS8diW3w7E+D1cy2LsqDeLWuT8/ARHuuEM5SUQBwUyj6oD6FiWVQZUBMWw0rDx+ffRUXeXYXSC+8
AvKujFRui69jqBhOsIJ4YIG1+MftVlgX4Q3WmGLMV5C9JNp+NxA+tBbkFa1xTrvUwN6mVS09TEOA
J0ugPaoprpCN/r+UF4V3KfIOqL+FFTP3o5rx7iSY3rTTvUhqX2oo1xKgPJ5sYO+mfYqSlcX6ArBn
Sw3UMn8UL9+w3TYAerPRJIDiTZJXmeySP/9tDQSrj6X28+37OjYc0+ayXz7WU/+srHBx98AZd6Qh
b3z7qCAUptd+pJFp407ELCgqZhoIhdmVfdDbgasLUuS5jZIY1L1l1cI6Qv8Cnc++ETK2xto6tg97
od9Xt0CTUqX2Ie+QOIDa8qKm9jAI3Za8aXBrnqkM21ItCGVvOBeBSw9VethIlSq0xgcDGhL1QrL5
2fEXKdzRolIgw+IL3QLv7kJCHdZ2QVFmZNRZGRTYeh33CTm+IkJaUSaF8XzLk2GRqmROYEEM1U3U
VdbO51ZjOXgGe3kySYnrp8XgIQ2Ua0DO+DCu8GAc2FgNPrNn0h4S6YQf+SOc3A2Aaik/jTZyZK3m
kQtCMAevqGCyI80nXhdBnKEdpvMSmipNN6hS++AX26q+STDU25+8fzhAuz9ZzRJNEUO3qtvBqmZN
ZNTnsjS2LaelJhf4s3BMofCkHqOZ+S9ELaCHXAeRe6Nmkev0WP8oewlu1ylmlWnt/2b50Tre8wuN
FJv6axXTPZqJ0bNoHpQp3ScJzXeOd3ETrlsQrgGRsUe4Whd3eJUwkY1RC3eXMzJuExSBfYoCUzNL
IoGnLtisRnGNdoQxrT2QclHlHRT6UyllfrTwDCqzhkuJvey5RNMUpTbrR+nb26fyMokIpRP9HwgO
JksOVdlkRJakbRMAs7rdsuhv4fsYPRebgoaghXKY9i91eqI8Z32PlUM9dloHBO0/E4gVvprycZhs
ueH9S9CP9WQzsdlh14NWWATMeqHLM2lUQweDBKOrnrYldZVvBnJFdpoBaSN7VaXNtZUchTw9QP9W
xj1k/NTTWHRiw5TdrfWwevzsLPhF7b7DsTLJW+UW7FxqEXn4tZOYs29LcI071J7n1Bxo7Ut3KmHR
Tr5LtTIXtpuUgep8TI3OqTIFkQpu0mzfizes1N+y28RkBBwf7NiTc/50tSNJW8OBOd5YC4CfB2Qv
HL9+kAych7NJGb+TI98liy7eNn1LNxuDRlEPWX80j3TW2tCfnRwT9Het1hi0yOtWJii7WcPoHT4D
x09P0Upwxv8SxeaBg2zClRCvwlMbyslQr3JR//2HFOptgIK88wnlAy+kgJEznAhpqHwHSVDokNk2
Sgk2nwAaBQusch+GH2TNFZ5KTOtSMOV2CYm4Bj1N9t2sjeJPkiVBXwQUbciHkajeZvBIQYF7Kimy
OkRk3+r6jc+N7PaGQT3tsPjbS+Gx6wpj/3xlqhvr2GehccDYei6MMy20MoSptV15M6/KpoU/sKc/
+Zs1Z2A17K7nck4jQ9Nd93/gfvmeKk4z6L5qxPGI2C1NTEgf/+xpK+pRKcrYN3W6V/b8fUEfFim3
ZUMvHZ69X3KHiTHuNNC5sbwx0Ytwoko0dTc8rNYrheY3r7LoCZ+BwsUAiBl8Cia/cGZ0qv2YJYSx
iGoq0qrKtApoJbBHeTuenk9NPh7RRUgoq3v6Z1Lvc87mtFei27nK+qZ2ngbSLTW1CgIBzg0EAEgO
0IKoLlFQnkNJX3VG/HyGC7tKJLlmccNRFJ4SgMio9bYB6GURnAEhy2/uunBAw2XJDqDWLpDBXfgx
nJF2b3vujacYTplfRLLxMOM/EYtZv6HlwO0luSxJu/+PuqSbJe+0amEMi11O/JHg9woOqjp1Lmj0
KjC2BtdVlxIU08pHiBzfS3vOkJNNd3BNvjdoNvxLVsIP0IYEk5kULZ6gslQ3tQ8T15RPnQ3EmW6j
aGF1+ab9wzSqf9fTUNR33o0/5rtX8UZ8NyDO794VFreZ5uUlfsXB14rOS0v1h9Mlw3oYEo4n7ELY
kJdoXMDH5dZqUMaPLYpE/ZqGwvghcIx4zJGcgROuNCyJyO5Sypv588nG5VXMicvt1fXusCFByYTN
py0eM67Nf+JazP1T2MfKPJCN0CulgQYAeumY6CEQ1EOuJyi7FAFbxcuNcLVQt0jDAKmDSWYTOCy/
Ejuo0i5cRpwN8gjqiZC0COiNhfuhcsOZV6AN+BFMnkahRJIOK4z/YJrtj5bSh0Tb3LVfY+y6JTRL
D5sCWSyZdfdUBwY78E+riBfNBK39NVu0UwIHQg5TEIBcB8tBHdytZGAYyTf3FKAmDql7uOpuMH8s
JuhZI9T7cDetmcO3tpkaAsgOFppjPFfzXv3NornjfcB9Fkj5Bco9D8Gq5S03lIxJKyfRWTv6MW6j
mko4nbUrsi8M+KYCSl+F9nW3cfJ1zQt7nSU0uMH42yMo/BAuIfLQVIaJSTTpfr0JgxBKV5aZcdBC
GLWjfWfVjP6tAHNQKD026BXj07mjco/NS+J+16e6W0rsbOHTeh7PVveKFNsudtcKwWy/eoqfGaP2
5UeXlySc3kOf4pkyuxxBIQNvIT2FKmaKRka+yGPth01TC5F61hbHsGMMPUILbqJjJFXAmFYgyz1a
QHEJyC3N9/0Pik0x5VALxUjKI3RhF0WiBROyFh6sny/N+4bS7clUvLIgGe3634+5L0DjPjvJbUzA
Uc+CbLJRnklvduWgLpVq+oyPmdfWNQzh5zWR5RCKW+gcUTfZq6G8RBagPMyJmLmQfMYvo0nn8NtA
4AfZdKm21e4iHlkZYXcejAAEPbTFeYdVxFYV/AsVrBb442Li55q2Pepw1yjE13yn83Z4QoQz4Ivc
dLBFdhR2lJXeXkn6lIFh8NoxLdop1uHh5p9go2GtmopZsTmB/wbSf7D+Ae7Vk6oNKc4J6YmJnOQ2
dpGkDJYnNkpiJwjV1L6lMDw+4G+vO7Cihs/mVYvXEsBWlL5L1acOMotygX1HXdVFPl7wOmL/EHmg
O3zyhVmvTjguIXX1HL/uaiiQIT/uq7SxKY2l1tfG+ePtb3EqZFj3D8sdR+jduYqB/3q/K8ag4y2Q
XWi9NJ0E8O2A+TOJVDf0qWSHH4W+TyBbAzR+weFxrgtG5GQCYYB0oMu6PqsCcrSaOxYclNLCxmGj
nYkeaaxQSTdveJTFTMz3sW9cw/a5ovawhwu4ThnFgKjrfz2h61D5wERREVyacqCgJwM29Z3/UOTv
z6uFLxI/rCQCgs+l29C4nKSlrbuHHVDKLZiXaP4P6EOSrcHCBvzoE+pmetOHMv5e+Ff1IhGjXQxn
z3L+YyB1H98Itam0LqT1+P6EutBcREALuHOuitWwEzIWSy07OPZXs4+jpRqiEwxwn5MqYUXMWjCb
3lKjw9qqJYRtV0gmEuSRyHwHe1kEz25QhTOxhzQ06uccLJ/gzcYgYWKiqq2gFOzAAlI/xTk79MKT
E2LvZcuwQM6sjLPF586zs6ceqto0pnIwuNvCixPlRi5AH9nIisqxaiGcY8/RykkVBsWx/b6UUh9o
lZo28UhoLSu0qcTK9VvvrGkl+4cWpz8el2yk0Q5Efd4thcNd5ObSNC0YcNmVv68WSAMfNWfN2Gj1
m9tmurkkzjDSC0tu78x/mQv4BYidE53GomUZYVEOJloLqxF7M2VqRnYSYW8LsjVaqlGuBa1Wx1j+
SlYZ4HI68r7jbuDkYP879dNVzW+l3cwvRWxl1z1M9w1TPJWld+fdz82ZZ33lvKqIHwqjapz0kmI7
OOxwf3APVfWAyXyNxLn2TJpEQDKWfvXMjcQhJn17D6sHqjrvN7L21BHYnJm/XHrcN3wjfe5sO7bC
oIz0OTarHHWXOfAW41RNupVNvofkFkB3If3CGRGtBboF+cL4Sk1DlzRl9IurH5QDmnXUkjSFmqnk
kZb37vC8RsVVlROl6baW7Fj10vB4ogkTHdyeidH6apcTBgrOMDChTMSTLPma4Xj9+HK57oQFa3hx
x2rJMPBvjQi9svCAm8PCcOAWEuYpbSG9/IW8gAxOp9ZtflDlRGz4+oxit4CQ1ZiXc3alcJXJSxyz
6VveRY/eQJCY71duKSQTuht2IuiMrVIb3+OY6fE4EdaOlly5nZ3AdJJuT4OcmfvfBrnB9vIV3xdi
9ZNu9WBluTlOi66WdZt6SzCGl8Jj7aHlLlcVOCXsvBk2WHMvyTwL6yZKyTz//AsAe3hnf7I8iEA1
yi3wyqvUipf56ktOkQWzUhYHZT7dZmDBNzJH3OCuHh2rMdybBH8rnrXfG1uQrgJkteASg9B+u9R4
0nl74D+UG3dipwx5f/Fu+NCpzGoj7EwSJrspeKj15TSU3QRG/VVOyO2QdaeV6AEjhyGhymASmMNk
gLitrzIYp3k3p3z/CqZO7SRj6fSIt84Em4oqyqO+9rBB3/T0F+585EkHiRrjKoOVhC1/kLse/Ckk
Oayr4iUTQMwsYr8OQmSdBhyRpRlfaRN3ukNIJ3scwS3UHHvZw/nwsAzMQbVHKNadWwL9ddCc27Ep
sVB+gErvRc7jD6SndA8yyz2ZZEm91XhTdI6wJOnz2ZPJrHlz03KfoedhlChsrIQbdqpaFNFA94YD
L/XG2RDgsjLapk7Drr6Pwf8kAU0UDQOXI0cZT2q9yN+QMEtt+7H6wQme1ljnn4YRKMPG5jPFkZm9
PZNyaBBR+c6O36VbHeoHMeWvmYGQoEWQl1KUBg29OsdlbsB39iLVutuUwKfdkO9i6FWPRyS7LosC
waEfzrIibg/ORC1wbk6aR1kqJG1QzTSsx3CN3iIw9zVdD1O2kXXxRYpk7cnIIXsJtLpFoagQCnMX
OI9EohzRhZPjD29nsvsvsHsMznr0djv/j65HNZTfX76ls8BeMhIuUdtckUoQGNqwQDHUXUrVnHzm
v1N4jyO+SYAHYTVvsHXb8+sncKkATQdLcOz4zMXZHDx2/FstCZdocbhn1k72l9rlORa7JP20nRB8
NWHeA014eEp6ClbxFdqAJVUzfMWh3vPag6jKC03Ho7qoPsbBKxSU8/hCbiYNecQH5ZvylPoUOu/O
X3Wh4oPqIDysucSyyWVhTL6lLqK2v4BpjuKW+Karq2hosACg52KklfDr4JlEXiBNUwpQEWU437/a
EDPgAz1iWPqVT8ZqvbGMFSsNfDzqLOBpKuRIeVDgboxdVjLL9/AV7XU8NMCCsHq5mPkGioBwYONt
NKMtCrvxEpvHEg9Ttue0tCQnkX/O15Pfmfx+L8c8MhnyzBUvWEVM6dwTMg/KfWsXX08a4/oECHR6
ZtyrlaFdsEND9ALFwc1/mf5xThWp8D0g/CHAWWzTMk469YjBjRb/nDkfq5UOTELr+8/PR+WX160h
h5gqXDVj5/m1S6i2pA8wY0EDB8Zs7NbAcVlcg+ziJJASkCNpo4iXUllN6NFFzF+jqY7IZDFc1MlX
QRjjH234olz3DXbf6oKRzFMvu5b4LIHjR+XdRlqVpx1wzE1G8+9s8fSMW8KgfQ87NtVvTjxJ8ZpD
Xt57Y4Lx4W8fHgsuxhxbKoSSbxL3uk+vwGttS5VNjAAXhUfo54DWfI5VbxPMI03urog4JbqG/+zX
Hq3CFkLZ3johEm7FLqbOi8pos0pXWGA1HJZ8AWLY+dVqn6RcdHGG3SjsZAZcoL2/aVyzo8bCon4b
5Q/EfTPgfpD4qf380h1SlyWF6LokcoLVbqSVx2cCGkjt8PFkeIMmjockKwpjL7lJflB+D/rLS0sT
R1sXgnk0S1j8zsyNHzGfmIUWb+mx67dc0JXVeWDmwvU0pa3L56e7gfCXhikmgt+poHPQiVuTkkJU
15EkH/npgSo5TZ6o/ob5ylLDqQb88cOpSMX0ka1LwRuk5phA1UiYFJFWJcV8GI4A+f1KqbaJ/oKj
sp9iPzF+THMxTVmGck/I/6Jc8wZVerF51UHX7LGHgeDDTiR6WwiqsA9QhWXsvYlaaEv/hPdZh6rH
YJoSQZIXcvvX9KhbCA5BFw+5VQuEvLL17I8RTRo4BOHT3jbtbhU6VCz3lgmYUwVB2K4hzidT/GOh
ZHd1KQvgJg43A5LOquqi+PmZZLOZj8Km1m6PcN5/4KPHHSEhEor6NdRvAxiKP57lp1oexqKsQ3Nn
6y0j9HrsKiQ50Fi+fuA4rrHA56Ye+GUWKMxCSZMKnSCCzVX7pFvi6Hz2q3+5W92lFxrjuzzNx5Xp
pje/9UaXEV/8RKh9rjPFIkLpArfDGVg3IlooAm1g8Fbon8PtZmG0muoQfABtLhl6LjOeYLi3loqa
47XB5q4EJRLDD1HQyzjlB9sJe6/wQpQysupuwKK4bcGCyBKl+QVkxoVJakid+aowjuDQgtqmsf9B
RIOz2OLfs0vUkIwBzbjAmu6ekH1pBcp+kckFjkam1uJs9QsD0Xfh7fdQdAOOugkk19kO0UPvN5ii
P2NBSeBajS+rD7572/743mAL8INvvrSxDhNtnLw5u1in2ZatQwuOqhY+frpR3lpEpPcMq3RVwyo/
4FZBsnKeYtJXQCJGDL6KqJi7qnrddFWxpZ2UTMlDIu/SwbK6+O0hvYJmoSLEimSgrBUlzjdSFL71
rxJC6cI3+OuLyPTGJkcl8KEquHc3ZMu7ZaNi2mBLiWOdGuuonl8pvZY5p7JzBHW/mFSy5urulnnH
c7ww+2wzFPLt9AzCTgnqgTOSaH+cOKxmoB6+JDrbnT4f0GbMNtQUl1jZm5g11Hhw1Mqu3LBbX6WL
CnDvBBmjE1tg9AJ2C0Qwt5OtCi0S424ulLKH59NSGgnWWLdF288NiHQPTclJJgZHbZUg41IoBCAY
nckd8yD/Ju7uVsMNnFaftUd8M6RXK3yADxZDaXZtQSe7YOErGISVMYaaL1m7SoDRx1slhx4Dlcl5
d8TQa07j+VyauhRaMzvO4WXQ0tfcIwA1Fh8I75hAzCzSfIf7JHabOMlh0odw2+Hj1BG0dg7xRQGr
Pm19DXKHgVh5Vu7Eh1ylfqRq2aAUmo8xwSHqFRHrqdKevzyQkNDG23jAyGmPoYI3vOO9+RKVKPOb
/KIypGsriNe85+/9GK35oDmhYgBchFmDCRn1Gg8NODSt6AvMP/Pm+3sScLGoCcCbnfRCHMkncbWN
2tTMpCGkY5YQP2cJtxceDYrzMgW99ySQp7G/Dv5w684oyjR/tHTXUaW7SF3JUByVxwwjhachGfLZ
cRSoXGTmLaSWdpwUhHjLNLbn5bRgOUCcq9ZDrapIsrmoAE1VmGL2Ty6fNVQpTSudIhmMEABLmUj6
zSCI3ANjXteh6ozmW5yQcxQNYhN5Hrgqe/bhfUA2LR3ylLmoQBkU/e4Na1KEv3lkzAi9TTltIaSN
JsccPq8ZTHlUqrB0BRQ7sBNl6bXmkjozakHNNPnyF3hBLV8bRaOZXExLMueUQXeMRkRpxDBmdYjO
0/i1TEzxJAf2X8hcVb1Xlgblcq3xC0lrGjysjxy10jZc0yUjrwAey3uMGXx2oiwxeZajk2/5Ou+S
5NEbply+Nkbf/yrnCznyfPnLIb0V3fgxiYT5S+nZKj++LTsrComRjoYMATvn73FaD6qf7/XlQqhd
GIfF1yCrhuCegHkQX9ROyN/2ytZCoa4J+7KGJF5I6fc+OUuGAV8m61OMDKRFctUs/k25tA82ECnZ
x+gH+USq4XvQE77F1S/Nvt9OfkMBYeSUiUFbjwbQfB0ER2nOJvTkCBShWg9niDbyBqYtxpYrYbOp
1o44PUy1wG8ceC03FXqbnAR014X5a4Zccyi0k3C67qSXD1YHPdmo7P2QcRPL+7q990SJPWsBg9tO
dH31kFEdUjfE9O3G9RXrl3bWU5RnCNdL2h0d443D4qkNAimrgHyWGHO4CbxuvDC2tWPRgesbx6zW
chfU2YeMJSFiBZXDZUG+56Nic9Fg0Z9sw740TL4r63uKqWf+aJmnFMBdGqD1l7l9vnepVGVqQ6iA
9j6JFyaQoTSHEwMM8/vc/aCUzd7LoKmG3ZRqFlB0gPwsclcejpUZL1BsOsr7Edzy6NY1r4uMN+gA
/b4YIRu3oyTwGS79fwS19BGozQ3sxy7bJYNoIHiCYv9AgYNETOeFlR/Zj0mHyWAPd/6coh/St8Hm
Pefn1qHpV4jz1VuJ0AHqkBBm18UUcIuW90/16w00koL6lFFgufwCG/24FqbwWfvWMqZqWQ8Q/5sF
sASuaW8YuSnPFNZMvX9HcsR5vfgSRK5V0+9yX4EMk0y0JzmANbnShVctbTYwjwTEU2UVhFPLyIuI
tTSy4pzhCtjB+n1vuqp1Kk8UhZWOfaeqAMHfUSXFgwZDqTPBgK+1lbTOGd9iKeCixSrbKl0q57u/
syn+dDuS4eWdFJ37jRetTtEwTjcuBLBeo2gNX9eTPM/bg6Rf6bVxtvhVbHO9qj274BWle5XBsGvi
QdYY1u2MhM2qJkQ7eHVPPmw6kpYEIEoSs9q9U3F2StEZcsL0KzLqYYqotKkqy76Vj8UVzA3SICuW
uDkNGInriQr92Z/OIvRVOsbdQziA/EhAakiGk60DScjo7AHrYROlv1gA0Y0LSs2IJ6LRCh13heeB
9JyPf9QrVuhmlFKuleMIvQcIoIYGA21FJjLt3Bc1D+v1+ZXrfqxprzY/8suWPpXks2Np7LRZpcOW
/kXQvxv9uslqZrl68HKfO750jwjDqr2Rto8QACX5aaKN/KHs5h0L2LUdL7FxITZzY5FHO7qnQZH/
RFf/1E5DFNyD3bUaB7jY2FzP1ZP4h+XCDo2fCH1PFHkK6CM3oQdlhL+7na9++nU5U7mOzBSunnP7
VE3NRrPE3t7qbVMKFawf+NNCOI0DixFqfJzVzQxvleFMuaYzpGErLwUXTte+SYBS1D7ICcXb1QLM
rrnMeI14Lg9WHRIMmGq2RY4iZD5UBsJE/Y5rhToo5oVpjpE4nDQepa36fjMssI7z4ySPLqu4c0mZ
O3cG33Ti5f9Gk51i+2dm0J0VqdlUVB26Kdxk/dWff/oTh+bEp9PL3ILj5Mq3vyHb0Wl28eFyoesK
2mSRQNonNQ7NTl1vAfbgG0aZiWBX2VN5HRDw7boK7EZlghKFqj89DGiAWX48ajKEAHLONIBqBGoa
INOZX5iOu9wlNpW5mLDTc20S9XrgMvV7WS1EOcC+KcM3OX+40HOiLMXCUUNS4eniy0IGY668t9gy
ieQPjS+Tbkdhb4KMgj1BPz8pB0LR4TO/buBDN4Fa6VUP0qPV+qbn6rROA8Z1LsaZUtMqjk6Sf1sl
z1uRG5KXYCQxhpVzC/GXlec6HzLudyxxbStlb9f2g5wlsOTKF6gOlPuKQHat2y74+BTRaDzmNZMS
WMWtgDkOFOWrN+PmtimfKMlK27YesGm3daCgM9kj0ajA9JeklK2fIEC4ivMbTIlaHsEQq4/y5Etu
hOYYtvc7PCrthirqWcMMEfkL0M1bluM1wHGSqVu6DTMPBhqGA5HA2BE5NlRbEIIyAKXJmJCrUKHX
go/HjNXMn8Ae34hgXxjL2/NJ92hxND5iegXAj7DIxp/eKu3gSZARoKyGsJqGM9aCLKp7nbbnBqKX
h7WjEEifVhvAgBDYPgRyMf4TTSJRxQbJH5DUOm0xuET+rqWwDExEiR2r4YIWUU/4fwFL3lVWRzPD
w0AMuvjz1mMx9pOKpZ+PfLwpH6hNynDfuJf4fCmCdd4yeMdBnDN7bAfGxU5qDqtvbDbf4TnCG2XJ
9+nHOuziiv2iyR8KXSpEHsZbiQivp3cH5h4ii+yqUQcZ7LT9IFEihyNeKddbdUvhydlVuZog1SRx
9a7vQYX4tLB41BPv64bCT9wZ4/b6N1favyB1stBjbHMCK6tGsfgGbbdrVEY1mXyADQq8xF2G4Xyr
OeETAwHXjxV9LewcX3RX8w5ONuUBQcOkuSmVpkV1fLjGMVxa8HgqFrP+6moPmYPtXie84rdjBpfG
rBNXqhYT/PWseCPju9+/o+Gr1E92QO0G2s0TSx8t/znSzsSJ+dP0TQSCVr+lJFyOLYxsumMBc3vn
U/M/ia/7KqZEjnQSA8X0YTdtGn7Jg5M19l57wXDWicp+7ahIxTbgGimXs5YLiLpsVGklIAQP36T0
6bGFKI7+FZwRx7bQZB05LrqNEySs63d4vKAudqFzGpfiosX/K8F9EHB3j4h1IddM/0D1oPX2M/Fu
2ksoBicEWCc2c4jt5xRYr24tbOINGrsBizfacVH0Fanv+hYa4nsBDpicdSkuDdfv5yRA4SwBQt0S
2T1W7F/JKDd+PGb7y5eYB4Hcp6DLPA1+rOoyE5dCyoZ1OxF8RCA0aoUAWlYS0vCy98dPkcI4iilk
I8VsThVSilXqFdpIWvYAqDYDH+AJMtMOEEbsUXyEPftG6GdYDWBRO6akOIWxiyhCU9bYkRkcVQI1
gedGXxa+QsmkwLFMrXM0h9RldwrhgTdIpf0t14Exncp1hRCs6vJlI0IR/q1Ewt7BzHBdemBc4Xqa
26tCyFQSGin6f+XVi9OsxK++tWvkOvV7QNN7WyTu5Qaz+sSh8/T3HFkI3yM3HbWs13+zOhFtvcYq
Tup/NUwSVrvLbq0iHzI1dAgTYZ3hBBKmH9OX7qsmT5BgFnNSF17Nik2KJoj7AdSUKWkqdKRrsAzg
9WNf0VaLpCltn2wJAo2I8Cu8IngVPxqOYUlrClAjJrT6EwGAl7zs60nnCKvq21gA2iwMK7IBAdGM
xpfJWk/Dsw1Jn2hwfmvM1DoWGhQgFVoI7nroISoPRoJbqPi8m2Esk5K+5lfINXREOJ9e3hG75pcC
0MfVDUeMi4CiiFuTsbOlAR7rsblxMDJY+zYUKsfEvJ8TlHbMdFAqKPmxVc3U7562CNzLZgLpfJ9c
10Mc/4YQMcvjP9rgTi9JUi2UkbIVjobtYiPLI7B9V8kuL98Et1bdmxnStFmFR2zCwRwVNRjeaauq
XOw9WExEj9zCNnp0F4aGD51LFOuulHkvEYsbsbBfDWQ09BYbZFJFo+ZlZP3ybImf78vGHh34k6If
KmeuJIkfTguyALSaAsfyQgN3MQlZ7z6pTtRwGzZVK6p4+du6zLF1bkoWaH7coirZzBJWJdNdUcm0
DCwl6Z1rBRnRDFsvJn/ITg24C9BWDcZBqPpigAjASZlizNMm45Ef0XSjmoY/O01aqe++u1xE60TW
o5bupzle90pNHgih1xdjLlj49ZaZDkZACmzWoFUrTIb0jL5CrLKGP78CK07sov0e9noTWTp37CX3
asgY0w9ET2reVXxExvypYNdgHE5O1GBj0BPdWwgXIF4w3LOOfeZN6lR3rtaRonaaC6cH/mn5Kaxn
COFio+N0xh9E0AX28fWTJ9uX8rmUTkMkIhUUorIx9PEs+Ndd2q1MGZflv/VfFEgsDzTqbcwYYgEX
5r+YiSWpiak+ujXq/VWu3RFkKeuxWRK/JAAKtv2QRZniyaieDH6Eo6dr5lyimjNbaQ54cP/EwbBY
W/MuyMajodba8DlGR3m6sU8PZel8+FNEVGoU/jPOaooyWLmw5S2RSMfy2gH43Ct5aO7O97YXMqc1
Sqvlexnz15ml1CPGisRRL41J4znRPqGWobpPBJZkoDQXDrGgYMI8yFaFLULqdYbptnzycfUH2Ow1
Ey6p62kK8EjKFPPCPU9UAxBsJ143QjdYodb5+1x4nMWDQc7txLrONKV6pK6KjPga9sQKWYKulWGd
My9dUIU6V87CTQQuZhPr9xTu8Xbzw5b5+WGQQchQlGHmF/IgMf01Z1PUalSSdY1sLJyHb5CuituO
j2efEZtVs8D7+tJRim+hV+Cj4ZHCR/NrIkj9srWSuTP263ICViFQbCrNe7WZR650CnCCPs4Hv6Qs
c2t/PrH9lyGbV6K1jkJxnLl/w1qbpiaVwvbgH8F6L9776QG0z0UEGh5goF/fC2d64NcE78S2z281
B13UAK3SW8kZ3uxT8gQaFG7uwSrBaJfrwZnV8we55JeINFTjxUZURzxWelHMkxicyYM/pJCi7faf
RmJ1Z/T4pnMcywsxDT3axNHGiyOjPHLIEO76DV5GqQIONtmNvwslOgc2Wnqb+vsKZiM1tG6s0kHe
egl2lpJWlMwXWxgmU1tlRD3IpeiGiTGo5BqFV1POX2Zka/M8RrgBQla0hb4raIXjf6s7x2+aWdC9
W5W6cfJ13IvdIIZEeC3AUsh3sp8WzGxFWkjpu6erWdKDyB6eBn0l1hF/AEak3yHbgHsezcWQaoG2
FrF8IRubR+lGxkGXJDS1xOrQ9n+LqLoNH77YA6MjWuiJ0JgDWpFdxmWAmdhFrCps1rTjm4QtRHal
c+uj9IgsqSUvmbv7G4TFgMJd2nsUz/W2WUzN3TSZajAX6dopu3Rp0xeDfeyEVkT7ss1QMkV318oj
pctUdCfa7kOp87VB3+8R6ll7i/R1Il/xFveWFNd1a8D7SehG20SMmfRx6vtK0wSZNigGQY5vHsW1
HKI88xF4V9r6UJsi8zYccWwXrvuCJmViQUxwUt3GHITauzp7ARHNMCDgphAhT/nTM/7vHInBjH6H
sHXmyanm5iI0GgRhbkTrsFialVyL4LOX7+ZshH4Q6eP7Bw2or7nMgkrE9bVZ/RxgSF8DUhxu2GGT
q1JEhLVrQWpxiUg6JVOzbS7DhTW/VkIRkCfaOFjkMfLLjavavI1y7L8r6ch+5iBcItmy4gTKx0pT
rPXfIv7SHL+dp2R7uelzm+3GLP54FUMiPo67j3U864S6SX/D9T0uuo7YAA0JL3WmqefXi32SqQ1R
oPwyr29iIQQGyMNF9Yo/tzXx7Lypo1/z+9gCHQvUnXI4i+fhohNyQZ8erKQyAXyDE/4kedFmsf0k
kdWrjuQ8qvYm/9bBsI/A2gUhFk8snniZM9EEaNmAO2PpEYlJblVo2PcY3e+5og8V0jegpC/YDVK/
pbIfK/eI4O932h9ktEO0Hb5r0mM5C0DuV32/+kccNEsqOqQQGTdUO1XAcR3RCtVRyrkKO04XgCL0
l+yu4CPKd0Ycbo5wo0XtL3xw1N131TZ6thoAxHT8kFMuDAjiDvx1PyjIdqp4y7nph4CAjdV5sI+t
eLPg9id5lbFdryXdq/emegKmK+EDb/R5dDQ70RaL7FAJko7qVMZSEb9tYgvxoWh5ftyBHvTKHQ9j
zXNwkpg5fm8QnFzx8urvxVld5h+Qy1CXyBzUG5T5oLlLA+FWegc/8fUa2HrnGuzWjukg/No0uoyA
aHhXR6SXCiIeg1HwyV25pgSozHOvtpj2vxaFPLfIMRZdALvo03vM2SvfpEh9Tj/hEK/6aZrqXqGF
eFpahHSnwPIg79RNvPjoC01HoNqEQVXRhy6/dhizOT8a+Owni+tqTX0Kr2+KVvz6zNkSfVx/Eory
r6yqcu9OS/a4HFLsyf6Epbx9YHnZ8bhTKwNHLSTCuyXZByWKTGwOOaO1AE4X2T18ZtUWu9S5+2Zq
y/t26WNnDQ/zxclaT8/dn9UPfpUKHYRaSLJ7ANy6jV/zEmQ2pjxz1SOvTN/XX9sSSjz7ISniH/mW
V56T3UZ2jIM7h2FlVWw7eYW1nDVxZ7hn5zDBRKvqREs0gK0KDjs9OwXYFzXfLsm/XyYsjJqZ1BjT
jV7RiJMUEzYY7TUfGPZoAHwFlbAtizuVQQ7lZwH6DYvwkwviqKYAUjfwYCYe7vA4H+PdpwoBw0IC
1O5QsbjnbpoSJQSvpA+W4M0IrZHegrfWXPJcYXGtIlYRGZKSbslBjfKZ2mNbW4VJy7sdTHHD+8Ti
Bt9x1Ro93W16FfXUdOEgN04rcF7y46MIGcClXch8Amk10WGp+KKQBKGnp5AMmNCYAay88C9WyK6N
dT8KpQyr1RVGJo2LeEqZadwudLDFRMj4S6RA9G6OlHtlS4aAzcrDOrFddlQwUusMwJcnyvk7+LGj
5Ohsp7ekqnaruwYBB5DSY8XQPv13/y4pykjDXTFH5bWK2/zmD80wcn0eD1LSPj84O+jRgxZ7eZJ1
0IPJfygojW6vIbRHaoe6ES5HaihxuJFFRhF2DLu+3Mu/WsKgcgzDbFrY0pavEibpn5ivybtvA0sV
CzsVZ5at+0CSk1QwuL/06LHLqR0m96OqVg7VyrBG/adXMNQn563DrXObTaf8llqIqZIvrbzeh6od
plrgvtarnrAEw4VVZ8f2XwY1XF/rpAqqu9yHyTISl3u+PTFCsTHdu7d2aB+RPYOfJWu6TbGP8f2j
TxxkNGp2l7RpK4egBdVr8nYsr/PcACdb7VFdrNfdb2JlQhWudTf6a0QpfnkPb5FDv/0x2bI3KG+h
zfsZ9Sfde0txHzZIXmC0kULFEBk0yZDYT/GzY2+zQIqD5wSEjoR9Y1yj2bKZjAsI3aD+9+Wub4Jj
xZs30FpNhJfGtCB3O75Q4JGjaWzQM3gN0sWbSHQFjsmiSbpahq4F5825T29skNOi+zYy6OzlVsyX
ych6Ggudc1yY34+wkyNPhMvjkof3h9hu6rpwdc/BQWrv24DF2tr1Kam0SWmdRr1EZdQva2AIzJFK
O1t3k2gZd1P1FHfI5nQP85tihs4HfMCsMB0tUxy8QmLJHciHaqndEbNz1jjccCMdqBtxUwqETISw
jFtjH9HgggYzFbsmJojIbUOY3vAcBn7WAfo3VxxLDQelqzxBC6sCl9UuRNqJUQjvzalHn8KqUL76
/hm6QG5J7fRxTIMPDqubBl5nApGgvNVm0QglRsMEDIFMYxZLqBGIzlOTA9MBcsWedrKbo+NFUZao
cT87RQuaX01SQcxcTrcocsgeR3tauOOSFJutoBKfI57hVBAG2aOG17lZYFJ4UnobddUZQd4zO/aZ
uOQZgRUNbnEVFGc0RLdJDU9jNMsD/GN4ul4cat2cRBuWr6wDdqLogUBzTLv8QBFNyergMk4ZiP5r
v3tHD4N+u5YF7LnVQ++KGzypOyU8LXE3B67KLrHmKE8PVU8Olw0cGH1VRYex4ImZ0Xz7Miq6Ynz+
HBaGruitQIBiuFX2/Srhgp1lrWIfip2aXmYoM28Jyc5SnsFaPPJ+qvADkrR5p5G/4H5Rb3Xskdex
N+Z1tmOcMAIy7yS9lEdmvBsGZWldhyHpoDhx3cqTwhzXIJgiQr978GwA73V9BtHyO4Vs+zZOct6z
gbtNszQKZ0jSPtv5l8dKrg75lpzxEBg9YlcKco0rz5pTB7gDkU3Qw1NNk9Y376AzZg8IyvxBMeiY
8cLlVEjkSCDOIhDaKydO6IvzGXNlUNyVEfbUGrFxpPtji02KRAZccpSd+G1LrbxHfCZhPrH+hbvz
UcCB7B4WyDLhaLb7AUAgFqldaNecRbCYXTPZwlW0KMrT4u/2Bgyppo4gCqgV8/NBDOJngwTJNI7C
YSI3GU8l3u1L1RCRdlDNoVJCktmCLy4TzfRakRVvE2pF7mRTDlqWfGO9uXZ+tYB+zEqyOaWKlBHY
9IWhgHlFfmxhRHj75r9XGbMhUYa3YBNKY+u368m3Buvxg+oF3lqPNCJi6vKSe1Rfvca94QldUk2J
iU0Zwpou3fDvojvJzswFz/L44836cgxnVdPyiVMn3Rw1Fjv80cP/S3TgK2cyzOUx3Gr02Vasuh32
xOibdJiL3+Q+XSfmxBnexAxy5w14XSbk/bJu/d27Sgr3PXa4rfIPeHvkcqgO/9W/2d/BRE1OHqF/
nrcjdK084gCu55NT/h2ujZrhYpGVSwu+pNw+ewL+niOtwFTCVBiZ24yPN9VTs7ig+SmyRXigvY0g
UvVxGNNGVerGD7qdudOZNISGywSkAngwjmW3VQxyxUFMQc3DrDYBBDWEjC2fU9hpvd+LYY0/55x3
fQtESo6weC75Ht4mS8kXmfnJ/u2+hkTN1p2HUU0VfvPvyJx8r5BMSa/JTuzEdoqg7lgv0lD3FbrV
qWJC0xXRtFFup1EKVZHbhDHQP+KYSKQT9vYDwmPTIbVHHxnG67dnX6HXogzia6NubA4TeJn5hM/9
cFIxQAjmYG0WZe6W8ytoL9u1HoP0Zh14h2p05Wf+C+b741isa0yeJIl4nHbDALhaCmJUIYSlpbYo
mozr+ow/01ZeXHLH4bnepucoPB7POzM4eILph3V4P49BTTDAmfrsgY4lebZQsa3HLyOpRgilMy9F
dLzA8WQh8rFo4SKb5esb4p4vGAtL6eJY5JrrCfhtXzAhEkriWso++i0dZFUDgv47THt8bO8zF9mh
XJZn3xJjGdVo12E19OB7Qtz3JH1TqwpBcjR+SrqkJ1kOd25ha3b2/t1PkSUlQAT6Kos5znWAOk7i
ioHeDMbdVE0KlemmqgQNyp5Myhc77ExX+K3KRxNATUHfERk9GI+l9NNLEvFfd6VASAbNRzaYl3jm
bFRHubtYkNUF74dc0xb8eYomzngt3RTuDm9qq/YOi+wGpPMl+iqmJKtf4Y/oKdpWDg5aR9h0lNS9
5yXgBUg4l0vWvd+86tMXxPK0v4/YX+aV74Rr6gj0gCe9NBK/FDuhnYwyoMXTd/UwMkx0KyxfQeZa
ct8k5+jRCqzjxYfFMY7vZc87CxGwoxlDhuLCxow1PE1BwR7R6hwuVGGG5ruzKmzMPEt1ZF/p2Pdg
wW+SO675v2U7Qx/ogk3EuRibTA137bCDpJazYBUykHdUakh+aY9qFPaalVnBcCgSNAH0a9kkgg75
8wfi2pcvInmbtvLx2fPNCyo+KgfTydzv4QPl1dRJm7/vI4eXBMEWdJRxkZDSvZTh7mMdB7CM+dQY
jiJqbQxxW9uchN6As3158a+JaIXpHDCa3R+U93h1KiSED+/r2JSndE3e3u5z8LIWNHZGg25+439B
jXDKUCaU7+SuO+m5uoFmlcRjnQKtgMPMVZw0/Y2X75g2kJTKhI327S2DWxHNT70ix3xt7pBrYmju
KtG3dwXXfCZPHOvhKH7nq3UETO6wK5cFV1t3BXYQKuew0PLED5TI6MTcH5M/+dSx9HNb+AkxUnqO
5O+OMcnHPBVha/3XDhpCrbr9oRrYb7FTkWMAIUPxjEAqWW7NOSR885NQ/X9KZL4j5riffiChkfWg
meCmKykiPbe1i4tjoH920lGGKZAg3nHgPhe/6fXvMv0vht6qgWcVPtbw/brCOHUW6ErdZBOePdCK
AnkXNuHWSc9WrPV272awqQcj4ezvNX7hqO5RWt+iTv3tk1XdPTDR6N894Gf4iz5hoEmOQQMoP5Bx
J7+utINr9yabQTJ+VB9NH0H8T6yFW/RVOLlDjPWk1CORZ+bA908r7qLPJRfg+losHozO1zAQIQSg
d8VVkQBSdKJv04dftp6sYasg9ggIaomHFMYF4MwskHsELxEYwXekkw4QxxMWJkPRJHGR8opdTkC8
ULMDj6tO9SIpH56bh6x2eAd9t290l9d1bBUB8HrO0N5Sw4WcrPjhdqsMyt3LDNlsy1jUqkUMRXJT
AyByISvqRCmx+Zg+6sPlJv6p7aTx6h9vwAwjcQyYBza7GOocQZHyz7N53/aXODpG6tDm9z8rj6+p
Svnny0lLriVL2u4DhgUJLyWoxiub7eb16Ayn6rBWloMtKHRedcXURSd9M9WCx1DfdbLqVEVZhNLL
L6kMOvBHmPekpxana8KynzoWr3ZDEZd99xsMnqvlJoABSvMPH83eCbSupxrEq0L1Vb1wzQkkcSL5
CzeOy4dV1BwIT17DY0I7hl3q2ShJtBJnr2WWSOfTkBWctxsAoOYqNTAZi1i0hBIE/1uteqcnsTLJ
kDXZeQqaGMCWIoMg5jt5oVGTgynQBxxy6QGAYxM35OdZ/otn7kBOgGvkxbcCd5L0qguYpdUfgTr/
2luuhLWl06U/M9WS4fJjnI4S3nPSi02IujpMlnnvjRig06uatphzYnlwCb2gTs2Ox9qaOgvpfjtY
lQWpQdnuRNnYM7SKAu2KC/G8uK2RrOmeb/YhRxYMNfl5VABuYgvs0eYiu42aXpG8tJdJXoaVYFCG
dwrNgMqh5sHAwfYYonp6M5oonrzBQIrodeNsWpo+Li7zz63pv1vD2WG3ZPLa4ySIGOUms8GQ9UTq
F9gwq+EjglzwcEMLLulQOKD7gF70cFOebH89la1gAA9T52gus7TYZ1eXHzNWMFRlupZEu6jPhbVr
NzvlMIM7FIf7GzqSO8+t4gz1P9QfK6ghGtPaRWs7mHTLUOhneJrFY+zDd8aOvfSu+R7Un8GNK342
dYST0WuViN0sSqLlWDsJ6fht+3QV0u3qvE6ZgyAMFPOihjj5FGiM9wdcSZAsS5fReuOTfTeCfO5E
ir0Fp/ZSc3J0v7njH2Qx9gVAmMZ/Fq0CEtsP7sexnk7Nrvrdh/T7keCoUcDDMUolYFKza3Uqwc1K
wVfibNVicXIOXHDRP40IWTM1ZIQmbdq0sF1Vt8Vg2i9+isngPK4gamNchw3LQ+XUy5MvW2mqEn77
orSmpxq5GhLpbqJzZNHe9aO6QSRFBhD/48AwJyAEUGhzsownf6QjmC30GCrDdVXCI1b8jhxTNBPa
aBVn/gqtN0p0kNfnSHwNpYLCJc1/QPy6e8BZ9t9WvYavWF01yuC3W0YD5aFCZXqpLA0LO8mu/fsw
A3Jq60kiKZ9yQz5AXusPMPhXBWS61vIsw3BynncJYonRxLLe5hX6EZ4K1Y5JJK1IhLDUdabD9b3v
Lm9fCq8MfpWCJSIZWGHv68q6yuTzWTbh/iWpeHUcoitiRLsLs01GiNPrSBmrg4npZLRhRnqt+6ol
YbsNk0rDsBNKicMWkSiJuibqAPiXPDHEHucaS0kdU4hxQRfBBUJaEAseOHgNq/HV0Oduk2ESgsa/
J1/1Sqjr30F+B0umW4Cxj6up0c5YmIDZJBGVBmONu1mU+wu3BpKjg5ZIzqlZG32bX0wFR1QFGEXt
pDjvsJDCvDMrbrwxR7gY1N96mT/cJArJivpx7Db/Eh62xE9cDwWQyC2r+Nd0Nkfqu5ApD2bRq/X8
Zy3/5NYqQHNhQ8TBc3tt/zaV1inWr+/0TSwvOfzXessH+FkTQs66dx/R9DfVq8+R5Mki4vk4a5uH
08nU2ylydsQo+6tvwTNIb6Z8PjuoegzjAP4zFxO0BJtTYT6njU/8eI0OJMBf5BrQDDf6sS3Ly0T2
gLg6aoOKc3siex+6ggklIhoSkcMydnZzWEAdKgTryFnaOEyziN3UUzhGRbceeRFJ+oRT/f8Nncop
LJKpcE+y99e6s+KVu0vSPMOzr0DGkF6zfJeWkScdxShEzZQ1+CILtH0MfedqSdBPPaTHua2swsGA
V38ZZH+02S8zw1sjDl1JwkBvLqu3lfGQPpJHMQuaSh7mBYyT0FXOu7kxdwBNKNJNTbuv2tauViuT
2fGjcWQFzoiIakNfwoTzAohzVTvArJI5whfGTg1tDqqhwUO6jtwUpxOKJk75BkBpPtz6WGg73yOX
Xn6QkuIhiBKiERYhxGzR9PWXRnwjPNTVTdWrylunsAvXEo+9T7+F7PdavIQdlbJAmDyTMIdsLhpn
043p0gZg0v5UWwk5SlYP+CegEOF62N13x5NO20XDMt22LsDMIIV8sa0xJf/iixkQpzAFJ5a7fmaE
UuFGDSXVEPYw3YkdKAIo//4UOsHQU51Ak8RhGWkOASYL4XLaR1dHufLaQ+BDZMRrSCht2xsbP9ZL
n6DnmHJyTqjA6BiJU+G4KUe5VMN90zuCwc/De8Tm6T4s5FmSl/t6RxXDWhEJ8uNbeNi9x23gGdD5
mq5172hKuPj2U92gJDbPzYFDl4dngw5mo5QTrUJD2g6Y8S2jRVvkeH59nTKonD/ztxZzPqDOHWBc
sBJhdi+KSlqsO3rsgUbDqFv8BLfKa10Napn1Wsn1CevmK0/0EeX2fPi20S01PZUuuPFMoi7uQJp5
FNMT7uSEuM/xLOC1WtoaA4GjQVY0nBj9SHby1/aJewV31BB+eng+FOx90M6VhoIc/nDpWgZUGREG
4KvOCxau2b/mTfVjF65x3ki9XaeOOap7t6Ukc+eIxf8B3hGmP+DQ9EwwuLMvkvzXzkrqlAhnL/mh
BlPqpPZ2a83iayyxcZd40G22H72D+rxc9Y2+0/IGrJ1bEpCnKg1dRx1iiOLXWwkphtQJJSphofSo
9rXR0J7r7dq3Jp/tHBjyInBfVKSQIVDQzjfjdMoooPG/mUilujm1ifpn25sQw/of4ZDaozT09ODm
NzOU+/HPCSq0djvgYCm0XnnhadetfYSjXr3O7RPLR1I+Ze2ifOrXg1OCkeSX+mbXyFiTHnPE1kpU
ejaLgmmweD+IChQaAO3X5St/R9zkL1tz9BoUPrTXKg/7pffoaA00jeSvGodvheq2ZVPNHV790hff
+o+XwmFgKWVB7OfU2zS0c/Raj0jABHQwGXUetEoAgbFdV9Muqb5K24gnRX0KT9f+g+KXUJH1I5w5
RJWKF2A8J9cFj9RvHFuplgtOIlv6k/JxOtxuOuMEd0IV/WFioFZmtqtWdOzHerqum7EQq98PNXDZ
BaRi3/N81dYlSH7tZjhhGyBq0DDFiYL6xgCNjSWWYZq0sGFp86UPcmUts2l28aH2DybnO305uMlH
WAE/kubOIzReLYaQxPD5mX6XAsrcoL4g+oDtCUjE0LxZS5Q3BIhbY4/CJ+jA6r8WxTzQZk6BW6Pu
lj3dw3Q+0xTODZ2+tmLfw+s4NIxLb4QgorTDXMXGDzdXVDXp9eeRasowjcxoKNekLMJJ6cBq7ZPa
wR4bd8o5xFElS32f8AnXYW2K166Ze43PFDGa597/VXQF7ybVGm/wTusb8yaMT4BT3Jk8RVwUqB3l
eDB9oknPSv/Q1mNKjkwJUQLpOfHrIqu9jBZ7RtYqUixfsm30l0GAxkBdjDiGuptQTboY0yIK7TAu
jDZcc6jdkL/DhW4pHFK/Oi/R1uyuyCQJ0Vk5oGN2frwWljC/LtQs9Vj8804PHvhfAwKz1JWEOw4F
rghUcybZGqiO3TT4CC4FjvLpm7ekQ3u2Wf5P7Dw3RJD9xTiQ7xsUDUSmVkaX7Knv9cupO/X5N1ha
KAthnVwXJRnI6WWM4a2KnsuaY9+M4FDMDhAu+m3V6xDJM5rGV64DEWgWl9s4drVLHmuWKAy01Cge
RrkV3UL8nnOkkCzWcmmUshbjNX3jjQBXrk7g3+XVFSdcGob5THRUIdohelcpIH0RhoZtQJoEqDyV
D1d1TM7Qx+LJ4T/WQcFEJxqbuSoMForAZWapTTuoWLzcwdObcmGvFxWx9hqV1wGNJtPuYcKQm49C
9xsPs1dFdDz4GCyslv3dz8iLl1MwYJAx4MWgPOjjdjEh4KGp0/txEEVHnLaxSIfsF5VN5Xe2NjT9
Qg3WTVdIX1HlnuuNCYRTojRzS1H+rFhzG1oHpabi/K+f3gyy/7paogulW2X65d2TXCKV37At6fHl
75YXBX+YeIUwAI3QD4deC0yXhNVjiLPyRcC8jeYZLsFrSJFLgzviuzpMyAsYx6NXjhdX9o7Gl8/2
8AbEhFWGvCQbbi6me7k21g4GsL9fWIkSBNU0pKjfC48bgjg9N/CVvKI2rWXEP44zu4uN3lje45UB
FzWeMkNvwPFPHdvE8cWGulF6CM7v1VroboWZOf7ITSe+pHRdp3e2WFbHdy1mGCfxWw5EtD5kP99J
qbpw/Dc7V9By4pIbMi1atfghTtz7oEm59mTPS1A9xQtLwi11R/EKAd6fFm+wV9cOCcA2z0AFUjAE
PSGzqSrjgfFV5UNl7TDFuR5u4t1/tOPyg3Z0GkQeWRga51d1EQRqZBvcRh0YwZJnKKwK3rii6+da
lBFQAmlguUCQBVqlUlc9BwZNxhNPMsTImPHfbH/oofOeCpvmWpyge4wTiqV/h/LP9zlx2bs4hQmO
93bHdbIqiSCDMNshnAomyMEnoqwTR3JplS+8gUVFztlJocGojUz/lOrQwfll6l/kJ0GyyuE/bFkn
AY/SbFJ4qKjxHFmOEwRKFstNGIWuUrVtcdqnE3YfhGwFzOYE/oOc5hY0EnPVk43HFOnD93fgf/FO
cnsGzEXw3ElFNMPofwHf5/9kk+8L+gpYy44VzxjpV81VJ0wIgoSbgzWnyg8c/dKDkVinnym1mDrc
QwCYx8SWmnWMyq+933ActwLDJhN0L7e7AMptz7dhGS1qYQlQj5tkSuHdB5Qr2CGVn2Hw/doMndej
hi17Z+A6q07tESNPXLDsercGG2S+WfBJt1KR1X2ZXNpX3lYEV22ZSBiv8k5aX+65oYC/KZaUyBik
JYjLVQr7XKYOEF1OScdhSVQ1kIh9FB+qIlu39P5wcPpDKcZF799kHZeh+3/8VfhJgB2HOdqTJ/up
XkemarO4qVkWOZQeyjQpP4f7g1YQNN1fhi6j3JSovx8XYzmsZlgMPRHf4fw14sgrIxgDi2+414Zk
k3/YRpt23LIrIxdg+BZkKURDeGEB7RpiP0CvQqcTk+kDYHu5tUea9nkQjOHC4ZrTzbB2Z3KNOHKa
J0rcLHLj+d6Hc5D6wU/EP6Ak8pQLGxubbnOQjeh72krhFvqFFQzyvfuaUlJVtVd2THfC4Q78uaD5
bxwxseqTxjtUrgjUoCl4sc+SBatSe4a32NC46YzPmw8r8tyrkQTCldFlwNEr4csiLrloPhgrt7QM
Vd9ZRuXpCHf/YIAC/tJZuuClmgLu0FFH3Rcw7cP1SK3TT8Al/K/tu0fTd8gjb0mnUbTXHtX3YtFK
9cKu+zihLn23xb68/qgq7vnUbKpsXNCLmLqy2cVUQliqWlfm8AeclFCxBLidaBy9jxsARPuNnwCP
sw1idU/4x6lQDXIjmV17BBjdyAY66OB9U57JoEleCYtnIMOkMs2+TXAfTQCGw+Q4yGw8pQBgY1Vs
1b7vfxfaehS7U3Nb+DpkndgNy58mw3Q18b9k/uYIWC4lpPEWpQr0imkMBvgN1U0pP+hthUFP8mlY
UmX5oP8hykNarj8C9DRyA2O6n56y9/1OB/kaGdDAeurVEI3xI+VP1BuaC8j5u67a83BqBlPucvdj
miRAKN6JIUyV+i72ymLlHSGLqC0NmuCJyAio7ucWITiyttsgvOgIT2+8eHLXO7e4WngF0FNv5u1V
BdWiclYJXBcw0jxyrvYXVHFRpcJZN3vrmcFVY1M9C9GMlj4yGokEj/LDLdzFpSlxq5Myictt4OeT
Zh/eDgIVIwc6YaeXcrqRloPbuAIuk+h0790sqVUhC1JXRO11A2+6PSPkS0QnKjD++pGaWQklczkj
FR01QuzGNxSB3TbpC1mCX3W+k4HriJcarfysbp8Cqnq8KFcnHYjgP1h+fQ7ZkuRpwOXvb3ZA67bl
bJgEhNbL2Sh2Yzrqm9sRq5mqrCYQMOst+6a18aT8X9uSqk4ARq7z6bDL5DT2jnELxzPpMj8YdFK+
Wng7G336181Gig2ebKiZwsViwNChDDfZOwSTdUcsZRNP+Vd/MFfzRVNuDWlLer3wQSJRKw08Wt6M
klDlBc8Sq48Izj24nbhrFjIhlpJtQ/mpoYEOeRoi95xx5D/IRjYpg3KIuGRyoxuTf/OPkvk9wFnC
u05zfIgoPvRLcc3oYWqB/fNeEwi29AkJ7cS3yPl2djoMQPaPHh6bXdkMFh5sg4/q9s8yBm0DFi9S
Gq2nmKplSwZzX42dAJBJoqKYjIm2wYCyJaZ+Q9YaYo3bqHVtvrPwiJN/Fp9KglW1Ml6KcZ45m+/X
mcpNu9tWBaeEZ41Bd14a4ocW4Lua55BQRh1TBm6RHOHudSZZ9DXxvnSa4rFilWyy3mblkNg3Oz7W
3BzbMUHNa31fHbekQALVRMPdZ++bBL2++972ArSFWRKd1al8S0pPzJXDMKbvbznZTFW/rFe9nEYq
lNygWA8CX0eD+XRS1DgOZzUZdmnG8PPiLsXG6FUbFJJZuQehZ+Hd48enYDchZhQYy7ctVBmVzJ1n
QVrXudnmGUUd2s/qLwxT0lGFbzchmP3OmDELdeYNuQFS3HKw1frpczofIiuH0/v6Y2clP7lj9ZFl
VrRiXwGRRF3vmy3l6cDjVYItIH3AEdeDKpllSZeTadEZN0zG8Bk/p7ZDiICwkFLA8Rw0hkpn9kVS
FsYNWGzvWl/Pbey7p9qEW70aQFmLiLfqly4Fi6eEZ5O9dJW4XvkJbpb+ciQxHovifULkonD5kFiv
zHg4QDlRD1LtFOCJbX7lxhUgGPyknPrK2TFYIcHcPIBqIvp8Lfg47knlyMAWJZj028p4f6W9UTaM
mpeghMN9OpJA9DLfstmwpDfw3u2qdE3P1YKFnZOmZockegiidBQeHe9OaTkIC4i8qjVMrj4FgowM
Q96NOCHW6XyctPAqjis3NpQWYI+gaqwl7PjNlCtCqXRhSPuzs1Waf6CThzRY4Fb3JeJjx4Xa4sQ3
MbX8rBHT0Xy8ehR8le68sCBYksxBZp5PERqEuHWP8U5JmpyPvNu6zOS8tj8x5ljd+krE1g94vI80
cRyOczeGyy1fC3qUK8apxp5f3b+d+TrpyPbJ0eqyuumzPv9/IAzegoJOQiQdLpvG2poYxSWeODqs
x3UKuWvCXjsr0OGbrVu1qtgKhj05n0cN4SeQF78sY+Ai1abNk22ARAwJkS3yKXS3V6KkwWCVu/Nw
Q/YE0l51LMQlRpfNubsKQzHuqtes3j5QPVNiMXop/NZNG4+i5KqbyOOcIdJLqQv/E165wv41ZHWE
KVwUTaHoY/TYJ7/BvDNbZulxHffW0E+jL/BOIvXMsoEWWWBQ6L9f74uTOKMB4enW5UpLc866ipbV
2MTAUBcJilwSLkPqiVaPiYMbZTL+FN3J38n+tVScWbrRvGoc9XmTykxzgaP+lTIb8QNykNNiia9X
iaYd0/gzf6wavmRsrKspi/cquhbaQEPTf45Ecc+tbn3vYyzM1Go2xZb2T5gyBi5ryyWQrK2Vpckr
xcZRHYDBOFzRAPzDK+dVaOECHAOSLoDYxnJAfc9tKHg3uExXfbp2oc5PGhbFsysSVF74/Wd2fzYm
kymAyOx6uqrw2/ysFb5R7S2+2pgz5rNRAreI6SEuZz/+mMdzuxsbVbPwn3qf8zprWBn3QkcKY9lk
Ui5rImGEwfY8dl/8ks8f0a4JsBMOQK0s6CPZwpZjIuujSVWHtK9kaW+9VeOLsUNETZoXjvV3X1N6
NDFpkpiFL9MpNvCvWoYjLkmskBTBt4HYzflIAtaHMhpFuXkL7qDhSbegWcR4EZSsMmf2ynf7dUkS
frzA/JFnr5UffhHkQEU9mABneDeJG4SObKBPoPbH1KLQS4fsefj+z6bEJPsBHXAeSB7sfgItWCXm
oirPikyfL1AcuLRejpwXvvxlkFEy1xx0ypadeYdtiZ4a9EZ4BSMrtPCEKyPkHU4g5POD2n6lnbH/
ToeV3aPxwALO2Zj5jOhX5oFYxYSdiE/0zwPpiCtI1wmz+b2+H0HibowiDPKOQ4zc4IEoj7gm/vxZ
RLeZkHcQe6+1Sv7B2T+80VJcYConKoLhNO4mi5LiPWsfswKgRXvrCFwT+HYzem5I47jEfcniXQ1m
JA7awzcdrUiO/fl9rSZmOCkZsVkrSgBYi9yUwUTPN7uCQqNwi/wYZuIh82paAyUdaMtUAEq5T1WD
g5OGmHvRPH5KdLBDzMbn0AEF0fvDvARgf3Ucjcj/HvC40Nid6gvtoQ0hxpEJNzg3IQE9OOujqWff
Wut5+RTLY2IelrX4Q7e90AfQDjnmfIufj0iv4sVbtX68w2QN2ujPrQKJIl3wDfcPyx6FWTzslC5m
ZFK6c5CSotAvcsp+ThNuLskP7ednoAkBmycPDrfSJMhOgSr7/5ZOyyaVR72xzW9NVmncucO+T0SY
5DRrWrFn5aitU+8Gof3yoCQlg6I4fHUijiHZ7Sd5gh4w6qIitMcdfVa13y/h3U2m0pNRR0swV78e
AZA400z2BmBpPVllVdl0TQX1WhAqbxM19HonufWHLmvu4PzNOltDj3QiO8Yd7ybDJBrZFo/nWBve
/dX1wAQHB46ZUf8Nx8Xxipb+F9Z/w519w2tALgWCFGiyjFXxJ34BzlNKN+7qbF14/QlpTo9Dxxv4
bQ9szTghLj29Vwr2Rfb/v5+1e3yGxc4rjqF24ANVLnuAgl3NtN87IxzQoROxJyLSSy63NBznDu9P
rvDiwIIIrMcm0o1B7Q01iu6GO73ENgXb/W9F9FieJEtvuOtVTb6+FhgKjBG2Qi27JjWim/Mw8kKF
LCbw0vtKbRQJE1GiSP3c0FacAxK2YOjqP0oprT1FQ39KGpEb4+9ecNM55X4tvLwTH+oXiRNjmBFM
P92gQPjttUXIodFqbnQiEdbwAthZt8hnFdytf0jDCodM0kIFaG1WVjj2/3YnabXKyCXKrCjqvFai
ghxoYPqjfFatkoPs0wUCp+Ep+X0s1Vdl/HeJhqFlSstTtTdHT4QTyY/QFQ2HCgXwaJ8Hu5cq0tJR
uqadT1Z5mtDruc/hMYHFE3/TV5BPbnOUZYVRvH9ZQOBNCMz9s+2TJFwdSUQ3flpAtbGMdnuq70+2
QaP5lmJZp6xXg7yzJlVijdcEQUYJ2lEAgH64jQLhYdRqKBWwtUSyrQZv2mPOvohVwSRrkTGX+Abi
2BpQJpZPabCyW3po98TOnuUArCUBMX55xrprgv1GzLRH+1eNtVvpnHgPJnuamyPqE8kNXAGgb3TN
0w/hzRjVXJyoD9DpozTfzMJucsiA7v4zRPb7PkKf9/7Lap4VfilI6B5ToQgKTsX9nTKRO82N94D1
/P1+fY3I71nOfvlhLDLMFtNgDVI/5DfzDStDKwZ0NRDrEJ4olrWDdRNow79Z1G3s7VvaqGqj+xVi
V5hEgX+5Bdf4xs5HuTvHPA8W1N688BG7mIeBDOmheYR1XVOlhb+l+RvzzJVT74GAHxoKzh8C4WYf
GhSNQFZAw8m2tHGydV+opaXz4svDBEInKu8tczfGfJAiPw4LYxYdJ4CQDqdKLbjk8hKpqM+nUXXa
YW/T0mdFMZCrCTKz95f/ZJ5HwFlFTePG8b91t58P23QNqTsTnBApRAdpRysn3RbOv9d/tniCvf5v
q9BLt1WhpuytnOz4sf7IGOiu0zc19A7cGorR3jo2ZPwWfB57rdefmiEB9ZqAJYNPRXFwXuDyPhVc
aSBwzPy5qMKnogplS4zNs8Sfi7qqNh4ZVBUzp350t1knpggb8MxAryvONs4y59P68fwpnnLBUkxM
hsm/gpjzwjLKnnMU91XhrrsUlOq9vHN8iSZeS0CqpTTzz9BtXBUCY9/dvP303n5sQl6Uc39O8O4n
3BU7IhKqXgB/7rwids9uXENSMYaUoSvjA15m+Yaacwc5cCFQiO/UpydfALHsb6nE7o9N1ziaMNhu
p00tMcTmg3H8y3IGZyWSqcuRlJVl2vLxVJfSScJuBgBlItwrcfTovE/yOGuiD7/rj3Pwax6v7NaW
BZSeFkuXF2C0tHpRKNJzdwnO5hohKE9GUUPafHMKnbIUWRsUCUGjVmgV+z+CwdTFjsZRHO6PxAWk
US2jci176vNpmAk73FzbYw753v/osBLE0mQ32kyO54W3UNkiubTMl/xGUwLM0qnrDVDFhlvmY8js
pA4GrFbxggrmRUgGdmkvhbrjiAq+qnCiL/5kr8S5v8wdhYtkXv7A80FEF9IarMmiv6tciHDuxYFs
cs1cem6rHTtCBn0J0TImQtVA9oT2RmXJLluKY6G4EAMHHPLxBCtf4cdJrTywyjMCmC439aTW1SFv
c25JOFaB7GuJ4LJT4NcclaI4I5VshI0CPd6mFjGLdGqvpf5QOU2wBdk26RNcMPvVdfOgWjhZf9i7
V6kjBetNcnQI8FlZJiJno+XvFwAHKngHbcNmnKqawfUYu7Pnn2wOHjeGDEgc2QED7DFVxiPQRU1T
NbmHPw4oCjqIUoCh9oCaDM2gS78+XDPS3s1z2c7vPvOzrdX4PvIwC25s3XzzZD56GZLJy5cSkp1A
RPBygpwrmqAsPkZPXh5l3VZ0mJJmi3TihhflbFcjqtSj65+HByl5BNpa86zeuahG8s9j9E5PvDlK
tKVoTTnYUyqj0YLEgyrafmFqMI1pUHtAsgYevGle1eYIvmtEzfgujn0j13Mr6wiiOSjhD3m/UjIv
tqXSqy4J2ZMz2lYipLnuugboLe6YFJa2dBfap3sgiwENhZseOlYQee0xb8/z3vmNQTF8RZOxLu5O
tZ7LxHSzn5PpTGmeUmJerzUYFV2Pdtyn753i5XJ0DZ38Q4Z4AQh+YltSmEqUX/3XmoqDynlAWsBa
VxS2fI3X2vyMhuqLZV2esfZPezKQcZ2VeviPtqjWJjiumo2KseCgsrTTI/5MUxhga6EJE/vbpDqm
oK1sUyHMZWvVwTM+YFr75TS8f5wCUJtPrm4QW/8dsMhdnJJ/PLCb1qiXafOPuTueEOJ38Zv5IHp/
K8cT+p8aX1cxw5QNsP0rf7eubl4um2wws/dYgidblVkGeIvR+TIwbfp0ThlBz66UwqFG2T0kHoLb
cPGaQOa21G2axZ0DKQvDd3AmuKNlC3ti9ugLsIRT71WZ/DhjDX3I8ahKP0KTK4OmPMyz30uS/URM
4Ulj0FOeUH9Kb0ABsTpb60GtEySHgXRqzoJ0GAx8EXB6Th0HJaMltuK30oh4LtGPe+4yLjfC3BdV
AxG1LaaGRw17c7CfvC1JROuPZSA1xsCqTCnHNRtA/7QL3WgWGCzBSUHftJu9mG8r8KCBOPLJzeDj
Eu4o8m9ydiU3AYduOhS5EzBitdPkmR8/ooHiky5vAdB3Bf8Fvd9AU0JvGHnUQN1r3po6N9Q/FA8Q
IG8duR1RZjvKRR2QRVN0R3hfW5/Th8wfHwPCvrAejVi7JMjigvF+PmZtUWEEAcl4/nyK9u6nz3fQ
u7Qmzeuw1RE0AocMStNWIejYdtMhNmY2N2IgS5HbUANX1chCX3BibuKJW1VP3Mjuz+TvWumARNLW
9xM9O9h81zYN/rjNzPQxQmltK75syAvsN74ZRxo05TpVmj/cpdV/MPlwO+rTID8z9OZNU3OVhGlf
bZK3oQP7QAUv4xxnnuRBLA8kXlyncJ3cPqlIEhMOUErHjC+YnfWTqxAGz21g9xH2S6TmLTzvXzTJ
NGDjPtibEQ/gJnP40lkHDv3r+6lIWQ9MDdS+TCaLgCyr75dLiQb+CS5LBCVz8JylsMGbCFIAz5zy
zCS2lmpyOXgOktzDXMzIQBI1InL0LPJsSVlF63VbKfuT2M3FD8K3CtRjGQw+ng3MgIPYGRvuF79u
iwzHb//e0d/37R2Oasf12exhIw9wcpcY7LcPO0RFjcfWTtbdeOkZceUZ8hahQhk/OoodQffm+dtC
O9XS9OzGPmAptyCKZJbxWdO/ezmbhtGfhduxYouM7B6sdtOX9cwfWFX/Kb7A1rFVdmB7I4Ol9P50
1T2Sn/lZLDbolYvh7DUadBAJmT6OyPQVg6umOdrwQl303I6VYrXqIhTKcwUq/M+iIf0V3UNLgjje
fLEIACjoFNNgryrDxRew7oLrJSqbgF9rbGq2Zv2+wncyJxMOoHEaqxGT4iKnhgBxFkZHD301Pyar
6brW8dl7mvBKR2YjFiTtIVzwQi9GFA9WcWNVDz8Ff//PPkrDpWBM734NMO9nWU5i2D4Vh5jf1G3H
BxBKttc10VjRw1ZYC4NuwXLzCa0N8unT3UaTI9IenT3n+0jwXhl4kuiSb/16FsT75z2INGs7r3UF
cn7nC4BU2SetBttKJzUPYv2mtdeJFf15W+IQTFm5D/GW6G7LPALfdaem0xTOO18QG8fSyxX4pF0R
Z41XI/D6UoISU+Y6BAv056eeiwCrs8p/zbQ/SxSaK7qQXxL8EHTuhhxOLbgN3s+kE4kxk0dRUcCw
LuefhgGAuHNfGtmbgZ6mNZf3YvXdCS/jFgOy8CFDm+0kWLlKaljSrqCb738YztIWOqc1RJycG1Xf
j1tKu07dk7QbiVzV+3/FCPuLiZpruJBn078tsFDBtiyUPYU68wEgZTCl4J3r98UDDgxS9mWdQzhD
mNFDxkNwBKPljcfLU/zBmPVKquYU9gEpgQgNM01K58DB1fTYNvYUE4xA/Qo+7M+JYRDQIlcbaGZ5
V1kLZqj0YMAflW1YGyTkdpHQFCm+QFSFx7TpeRT5Y4KnxTOws52nR2wuKd0zR/iAbKJrJIg4d/Hk
LtkmjAoIVftU0U37Y8xE4gp5vJm86jzWWKpYlr3pfjE8WcLb1+Sar/0jKofxD+CPWg4I45xxlZD1
j8Lnfif7HfdTdGLmSwbgrg4pgZtPoisDNWgu8IbutVahdF4385Uc+oVEEoOUQD8IYmpRb5/BV8f2
uI2tpm2bJAOdinevpPGlwSl1KBemmyCL9Exp2a6xjBZTNkEDl0wJTRvkK5JIZtX92YSI9mGDm1gr
ri5RpJMcz7j8kbqU7AfVLPEPxhLdKamQD1c+HjEN0ihsZ+O09nbn9nFIl9aa9cOQwVf87WJgOHfx
T2A+GFAYBqXuchHVIMuGSF4doeg09eyjzJHPTCqDJoMjm0v+P8rc5TEWU2YHFAH/9ctDLt9ZkwyC
fNe+CwMVdlPvEQAtc5hBGnjeN+V+rmvAdAn/Xa7lzRTuowHaARtNw65UyBLirgXWrob2el5Izqic
tY0d7Wxw/nhrQvkOTW8iD4jQKd2+lj/yfscA2DKaoo3Rh3IFzYkyUDGeme1wY9Qeu7O8Iy52H/H3
shnm8EVd6HQSBgIEFqCjlc+L6BehCisHhUvyq+RRII2JFxdPvLZaa//yp+JqfkFa7nZoPfC7vRvk
Gl1v0cybNjcCtvFaHYl3NpDqptMe8hPoS/c95R4sCJUmfqMOcxTFvJu1qtaWuz4EnPI6HM3o0ksw
fF6HZhK5DppQ0vZ/lxnTSWpknulmaAcxlOH1z8uUMewu/9T8602prV774NPKaWjCJaH/+yfinfWp
EMv/5TOi3o+UuVuyRPvR+qHuuvehThOb28a4slpCoQcFXw34liWJz8DtcswHAtnYIIQUHOoaVJn1
CCRj43kPMelvAnWLCnz4AweQxq3F67VbH7ZzwbFEpB7ThCXrhq52jKUzD5eRGsFtk/NyADWA2niq
+fjNjvbU+hLUQxaOfD9FJ6NuMigXoABTFcAVbL2NUu/uuMAenhjZgbjKy2vB3d9O2uxXM3ZcHLRS
reQ821dBa+HON0/ydROLjwXPlGpjGS/V1hGruDTUaS7o8F32f89GHrb9UeqP/giXLDpaAx4J+Lc7
FQqKFVwbQtogZCqHt0s3hFEBAsBFrQecZEWz1hgheJRqvokUJQimHDJElBKLSiMCH/6fiWgAvYoJ
8JTmRjK9DpPeiI8zr0aZL80NZ3ODZrec+cdWaC7kaZMiQ1DlHpA9w3irHgSOL0g19Bh9TnwLSdpp
oP+fG92QEG99rwSdiJDjyL1Mcs1TuYuWWQwBZT+k8QNU3jakVgpE8p03sQk+QbbqpoCbFu5kF0dO
gCCOqlNa4lTbmFJg6C/wYG9zT9JJC/vuyq14JWajPAOrXaiVzLcGdMpBq5U6umek2kBp+b+OuwO8
kYKrfcHmDXzXAhMJoD6WLUSKwua5VH9RwuDF3vPXOznqmNNIXNW8TeEq5YbCZdYUzK+cX0nLvgg8
1ZSPt5ZTVHOLjF6fHuvf5dCTHH7MspT/GINZXvFm0/+uDgVuq7YFS3v5hX2T4c6gY2O4BT2/Rvqh
GPX7GXO7RR0iAH2ATit2wofVwf++Dr4t26Ik4AdCfUBTGuXyGVLTivrmZZPeJaHy/htIC3BzU8hp
I+x9pLFgMuwr+7BuRCGbNLcEbmY61FVYs6W0oO1VScRP0+H5xSDRcvU08D9x2H4MBRlqVgpFnuu/
NcolF48v0knGthaRiLfni+iGdoBho/AAvtdq+Jf8kqKdMw02Mys/Gj7M+M4RRa419kP1l0gNJIAb
u7sqyZm1lObAgWHnFU791yAsY3L1OdCYKy4JIuWUT/2JMJBXyOX5rRpHqZAElMai3pqL1BooW4cB
vikCFYUSf6iIfX3637D3pERhWbwt75GmBND6zHbYY3jlPKH9i32tGKGVJ1QSfrvYDXgE+BwVm+R/
DPjhaY8Ycsiyk7e1TCLx2ZvjKGFXhQhp0+74gYV/DW08YOFscdGHannITtMtuBGfJ8thjer/saFq
b/9zCw2HcH8gX2hgRkSyhx2+4iHG6BaabSU7KTwWg/1tYk2k9s+X8Z33VF+lsnqUHOoTSLkYc+N7
beA+aCjsIemBKR3gfnkKjn1zsKDIsN+aLuPEVHvURnArkdUoIgDyqnCpPOmy2wc176ItFpNJ/jKG
Sk+9TIKzewgmW/pnRbJ/j8sG2XKgCyTENEXXSOYp6yEqKBaeLQTSZOtDToDboS/MNYdHPjOLIA95
biwMuOeCP74hfMErfOmjTZuRrBIj4mgPEwUsOkJZgrHPd+oBMiqeTP3RL+ExU2emoFSZY4H59Z0m
Oi+toYBlBN5XX2tM7epHGbB1wTkB97OW6eSyfNN3t4/JLREkOxpA3riuKhzqjFrHfPnVVlyORunO
GY+8Q5tmtBRJTtPRP3/BUQ5sNNJMHUlPEm46+6hon5m8lhKkCIeRWe4NjUzTPfX67XKCtEDX2ZvM
uGmhluZMAXKfy84FUOudUje9BXwgpBQZkig8udtmv/0uHbv3s1AqtIHoAtEZ547SXdPTQADNXvgl
R9VfbZTHg4PeDG5N7Xyv0W8yUiMpUl2NocoCbYO2f0lszRJKHT0KnWd9iizNYP+7h45uiGHmq4jI
Wwexy28trMJ0U/vIr5TzKgUpkqN3Dh17dItEizekj+b15EouOKDkWa/Qdu3MfpbELR1WRR8hLWhV
pSLlGpPXLYnFvcbjgnG4ueMv/R81MGKFW/aPdycYIFBPI8fIIHmNJK3PJLZsSgrNSYKAEiC/Wgi2
MXK4wfe6G7IST9MluxFflCjbgFoHJz0B5bCvMqptZchlwfIlKY62FW4HbPLq9C1gnUskfgxTyizF
iCXiJ8tfTuwhw8ACSMmbFmSChnutkKsqMWqa7TH5Byf1cguAE+V8A6OaRmzU7wX7KRUdYTQf7EQn
A2hoSSFBYNna+NodSOatjFVPYadVafEE7i+r005vQhzGoI6kPXWw7XStWhLni6hxUx+r+pObO85x
+Ipl1ZKa3gCRYVQ8T4PFagCLn5Temj5XE4zK2Ix69WlnGjZ1PEiTW16RBV38IMZ7LUyY8qJnj9o2
H4VeI8ssqLm1Fz6ZkCuDHLfeeq81hr0tQTdhbMILyletttpFSdEr01E/X7T1fh1UkCTjp28Rp/8j
Ry+g8NmaZV4mL+YOv17W2brOFEOSU/0TGbt5lUmEqPmLUxoZ2SZ7pjiTqNK3RkXCevbRBO9XtRFH
kJehgsxLu/37J2HgT3/pXOPnpTj+gbWG2xDEgyyU/ReeZ62249+KZyQ2O1ZQ8HnrmAqWijeutFih
r6qb8xOD5HDY7ChJKyPn0Oq+afsp+r5rCVI0d4QVfJra4+SmE/eu+Gjoh+Lm3o9Qw2T3+tDh5JYp
0YFTAv/TEYNEfcCDjezu815Y4JE/kxJMmvWbnVyCwRvpoXMek3xdipwy9ZJQXa4WCGXXwaaP4i9O
IoRRYgACj7WmI3hCwd0fcCTVkF90MrSb6ct4MeX0fh081cHTj71oh/U7mKWFHRmOxW0L98qFA2pz
JTXkaqHkgfuwXcMoec+DDj6Qtod748k8VOeS1Z25V7s5maetmDy4DbxCekABBlu7UfEJkmqgszac
cPxnW5eAS3zt2f6wL6AYddRAlOKKb9qgE/t6t1PkvKy5YLQe7Uj93UY6/FblYFaimY4e040joMAD
3p9O3OVHa0ewDf9OWNsB6jboedjMtTtBs5e3CO+jIs0aIWCS5GXyTd3Yi5FCXG5jGNAQwXJnwcEj
GrrGICetib9fv0Nb6LKUQ1nvnWEYO8z96frt1hqsZAq8PtnjipwryoYxTOaTGXDoUoS1tTDuwjH2
Uz4ZjR2m+ebS0o6lC/jQiecafhGaxPubIt+r7pma85r5X5VVbPVrjPtaphKcpDBFv4a5awc94dFj
dASx6t+g4XSTYRplGfEisyptdi2L+9UgHcWv2VOLBuY+zIqRBVtpxXZoOH8yyarO2wW1JYy1K1sj
VZy83xsSdmDKbtb0pV6DzMesRqupkd484Z18NGHTzoQVDYfuqDMJ/vdK2NjOvPgg6r2IDIYbj2+w
TBPQ+a+/902qTur88+ZKh0T16wgByp63ZdmNWHoGCopn30TCkiaDDz9Zkow5aOZ8mlCdjk8N1Knq
snOSa1scYkeW/QYaCi8fL9axieDEckNW8KjNgdPf5SojJMvY3dT5s0k1ayfEv+2ZJTUKYzBGvXZB
oMhISw57Diqmj8k2u3F4lxbL3KIQQuJDVVS7STz/EhITPCd4oUT7QUqIm3X6Cw4tVkN0e+7vX39q
NWXPTum7hfXVXFXfL+NMj461B3rSZ1ImyPUF2x0D7tYzWDXDbKdSP0bDfikt6r6f5n2t/hsrqGfW
+iCVqRUCYmWCEyprO5CYYz0SR08mbDWBJqYot3OrJ0W7TZJVH9oNK/1woGYEGewLl2o+2FYow6+t
5L1IyjdicNE23iGbCULFYipgx57DQUJhrdXOhLQKmVlE2nm/QrgI62xRB2ZGdjvChJrNxpZf+Ns5
o4tEBWyPrIoG/KadkIlMNeFZMrWwqtKE1yj4K9S1q5d8Bw/EYGjUu0LujLYpHR+iwoD6CRP8IrDE
/+C8HA1OosT2izldu3IU1yOsHsXl98rNBPgyKFMr2cMqgQfhNXq9h640CbZsQW64ef+t4rdU9X5V
LXRWkBZmgyK4eLLsMRXU8p2Co2839FmCBx1VzWNzhgrf15kXxKn/vBAvONFVs6MUx56gCztxRFiz
FhQrCx9RSx0V96OZGWcn7UqRyqRMO7BkCZPSe2ulLjTS6s0mtkdRzrb/LNTbGeFgvlnAEGVVf2zx
RksKOkTKMd4sc8bUfsK9pspHDvINcmAVM5U7/LneFEWYzvUMZeUHXzPD/V8ypqg1gwukCDtkA14M
xvDjTRt7ltc2CGUCrwWJr3KFc/6tTF5TSXxdPveQMwvdfFX6/kBEnB3X+D+2S7o3YllKAATeExWp
hIP7kVczGAhrKcW5Ae5CwGd3ipbDz/NdeSQYPAIVnvSMHOLor7wfBofyzbuufT8IDKpQjRuRv5lC
N39262QDsMYLfUNvzv4D34MbgWWKfwdx4at2lssVUJF0HuayuQHXrJ4j1+S5ETtijitYtYbxlM5f
IpD5bfona+jsxAG4Lvmm34fISmxUWD9qUmxKqFfdmVv6r9jc7BlGyZcegjDWWP4ZS4P5bF6yoPEo
BAJJjSCf55grIa6oIXPmhfL0VwxqUuX+QftsD2DPeHBNjH9HJMyeDVEjpBDDL9Gv4fNoyBfWOjwd
SR0OMl5kK5kclljjJoaSBMlgTYLu8QeUTf2KPFoQhLf7rgTBE3PBcdwXQ5rs68KXNbciiFOtYnIy
OJD3sjRpGZwbNt1qzyCcum4qAdrFsY45K9EEaeYps1rx6rO2CKU6Ir9NO0+2b8lXiLAgE+9TgYjk
BdOrH+I/TDvh59OXZaXNc5aUvRaWayOkpRdp8oIWJQwZgx/VG2fobt2M3niQdL/5fYVJWeYGNOjx
OkGiD7Dsdz+6nerMTvQcjyDOElF/zHa5U/in+pDWD6FA3LHXT0P14V/tEL/g7fINPhOwSzcmAJrp
CdeXEdSJbHMDaJpISSUHGKYk6Bh9GVxUA51YUP+UkgrXNC8W+/809u2q33lZHIMz2mYfABI+Npzc
z0HYu6jbnEBR89/4H8XrhPq2KJaG5DfwZSkNYXUV8poiN1qgJC0mH0ZN4S0P8D0Egj73VoJZItz4
CFs0A/vNnU1cXPlX3kMNa0wdXEvWvoQbE4dnoWI4bHGKbMsblpX4AbIO1xFFrCwlpvnIyDqFkpqA
jQX0GGLPbj6bJ4vgH2LQiac7raLgO1u9g6CTMQ8McxsVPWzsjS2p5z4eobmFZZvF4+HdNEjW711g
734gaNJiMDP+EgLDfb082GT/Lj/YP1ZMNdThslg0jCjIOALXQoXKtGj3Fl4YAjjS2w657cBxAkVr
Pl4AmzeqSbehEqFBQ0SKyqUuUvnrvnKGy70nsceyIesS8R53UvSKlt/r5JRZ2whwjKvYzOB5+aoC
IjOJP29Bbxcnez8Z9Qr4j22AG+U6W3axNDIVv5ZwXuR2SHj+rheocxnLdNkp0vQ5NTkhfljeeJOA
6X8Q9ESj3Uo85tpmytoIUsq+1v7MVG0WM+oAK2bcmFVBHC+NInhzlLnrhDN2Sxhys0G6SpwQYXvV
pajWHJkL0hWF0vSgLRAKCsTPLeAwKAf/Pq0ZgMkD7mx77BoEjAYtENivJjDbvxt5Rq8kvBwmCoKH
WZCQTRJx/dG3gwzfyKN6IeEJNtGD3o1yIaDyV2mc9AP4ruefXMfXYOgwxmi794HeZ4CnKONvmSXc
2kYJThkfFWlg0M6rj75RxAACtDwDdTukOQLQ7uhRQvk1GHtuYNFkZGh0tVy24i0qES9lzINhXslR
qtYzat4gVOfyn6tmeijJs+/nX4+0j/5HQWosZFjKwLpbTbo2SGqJFeDd6VbTrznbXPAli+oIMf+y
NxKvcYhOa6mDUPEbvQUENUt3wd101oWmmlPFdjpKfyMNOR1j3VraH9GhFbrhm6aDb06UJQy/zbOn
w8YvP6xo3mfiLl9/pRnmJ7sUKETcLgtAahsV1eI14YnQJ1PqYKUMzHbe5BXHeCZWLzAvyWc0OD1j
6ggk3VrtxTEluCeNeLKO71HLtE4U6mTShlMwzeXDYQDsexefuEwSVCrjKxpzHzH2zuWzWXWjhWui
GV1JUEnvHoF6G+cUuK8Z6JsY1vGpgGDwagsa0WQwYmgMYPmQd1/MPJK4rvLft8/1oFmZcNDJbO68
SIOI5/dmX88NHs07uIzNJu6CyGYWhMESQvXuskhP2fPIb4dJd3b9hxAxR2uH9Z8jz8ue2uXrl1FH
yeWsy15j2gXuKYU4xF4g6xN+oz0qHV6yrYbSFJT4YtbuSBrToknacBkfT5v9wODRil98VGP9Beyw
eRFZawXg0CRHoirrX6/f0fOF5cqN8gv8HfgeVLkAaSqs7Xn+WxhXtAqkUIIqOfNLDpQywIFP0syW
L11R3kZoBY3LD5rhUR5KKZSxMPfNyrip0OasZfkZHY86AHCdNPKK2dSv75HM32y7PyVRzWZa15uT
clfTWTylSbH+jkLhxuM0Sb/7aroj5ER5nr+RxNAcD863H/duD/1ypKZF/JMG05Nay+aH4/TJuqOG
HhCshvCgeBqTHMEmWjEfvvwP5pAmYotRdlGPnrTYLDDYpC8/teV+SqQtg9h4mjwyRyvSXMeSik87
JEVb2Dw6lmOzMpRVKAnlkPlZNR+upvVPs7/DwBP0yt1me8Rm1f9ZdscO2Ep/yw2e6KB74GUIrblT
9iuiALxBbHA8knS4YEK68FjgxH7GsOMwXxDn7dbDnbU1V+nH6HRR6bV/hgUlUHcA0LgzKM9l5sSp
K/1OsQ0daIknnYsFZmxcpqoeYEmEs7BPVl5fW7zL3iJW1SzaK7uvkNr6LIv5uFgA/4o9TVsSnQMY
2u7O75bew5Q+NS65dDhLt2iIBw4lEPlN92ufV69jvIETLqJrjGfAV/tG069tEaE2tbV0yZmn7se5
bts+DYUa/YicM6t6yVdgy2NQBpazHBiaT4+xk/82reSqeqMMvjv/PfxM8uBqVVTPYVtH+lQennl/
33dpDdJEA7+J5GL9+HDHhPXRPF2hdlbLNdRe6wMf37nBxDUN+GtbuX4is2SYg21KjeVD2S+MxRm6
JvaeUSqjaAw7Tav8VOeFaj3YGsVsg0+tzJAt50w7JgRImA6vgMHNdxdEbi4zBdUmUYoPKsNXubpy
AJGvxfP9coJbmrckFGdgWUzalzDC7fDoWCQS5nP2dwEPg6spFm9emVoDsl453XiJmGaOjZbLDQBF
0X9XVMaernxvc6bwDBd6RqRwZ0aVBsMt8NB5eWqoqsZPiaK7HvzRY/Zg7x9MDHrbrbev9mBRB4wk
MmkBgr14RBAaSJ8LLGBR0tMaWWPnGaudqwQbsuxrweknTJngNPtd1iy9/h0IZPQbNoyG6PEeINpl
HFQkpGRebQa5YYQrUfBoXLpYqCWbQ9lTNvXxTiFKyJVQPNuDzcU6iUAAif9Iqyc6Z38mwU7lAyQh
aRVxz5SJkGMl3I3GFEhSOm/en5MACAwApXslRmzX1cOe7U3pQI8AiA/yjwB4IJRgQYIQ+fkgWYKL
bYR93fDniyJ23pxSzmapxx57WFVQYUkKHL0snE8ptbNa3BIM3YGith6moJi0tSK3bw9g2Aj1AY4U
+TFv3WwRIyPPf23R9o5niBGRp2aWS30/gTUHKZG6dj0oG3hWkaviAG73qenCby18lr9rhmew7iym
Q6alRY9h72vFYmgQxFdk3E9zIM2dqK9oajc6W8V/R2gAF6o38tbzH5jtYxhkxz/zYHj1XKi01PeJ
YRMQmKZ5YllPa5TAhKOcaGW78KgvpuH+vsQmqj//Gj2ARbZexZRQSoCOqBn2vo4w9Zp0y+2AVoaw
dmYSUcfKfOfZKEb9FAgVA3xm6OIaHSoINRnxa8D+U1ARCiHangrVrw0vC3RYFkwbGXa0bgUgF3Og
k9Rl14pA1wpUaP0KFghVJH6RSeE2K3twtfU2KLb58C7pBeuHZ+TWUIrBpYWeaoD+AC4zEvd8AiX0
MPajhz44a91+XlTLtM4fDFFY7wx0tWRRrDEu5DO6IlsL5vpKMJpPvQVP3z2onQIsDcqn7c7oz2cs
yvml921GkZxK+T8bRmLSITTQyn9vTeZGIar9qEyRGIje+T57/3Fa1rhTE7tbC/EVQmvU2cLqcI6V
SktzimxH/1b1/R6YVbOv5UDHp3G+dKMI1CvFSOCmCayf6XlhgI7zwikKHHANHTJmJMrz4Vyk3msR
1wVqlhT+dhJ61BuyfiN0EP5bW2nbZiwRIs5fNq3I4a3/d0DqKXTV8mLwFiEdWvXveXxgwiLOMP8G
SibTRhUqFd8Om7kZrPfuHaz2GxqbRbR+pJqSc8q7yuMOjZYif8mv9Uf1mMCfvDVWpITKFaSzA2cs
OjvKtxbC/j5/SaoMyzeEC4wmrDVinwVFqbahQN+48zPJ2p7Py1cYFTyfwRry7p+TEVqaMUjAgSlE
HS/YgjQiUR5rt4Ck91O+VilQ1O0C/gvKuABLqm59M8lpfTZ+hbi4FjdqUo603Z7r3hbcjN7l1rj9
K4yspiazf99gZRj9pkTf6YR+9zEOhzkJqX4hmeGLF4X/VEMOD2eT9VPEfJAjXlJwoUlV5E4flrj8
JlCiF0rNzZw+y/4tUOaQBGIki1nSxVPP5Og+nRudLl2EuhAL8MQSSM651P7h5Aduf4GxgotH+W53
GykLGXMvpi3qRTm/YSZiXPTNfMBHm0boQCOxOQbMIlPQI8CM4hF5FO02+wVxA682UT7cOTv2MqRj
xL7cxBbSEUKZvhg7Ql3QXKCjnDEKstTG1tfB0+xnOqUpDOYAHwYWiVWzsh64dT89MpCBtoxqh8SF
203js47n8VudvlSERsHVqvIZhEV25havZIzP0c10QgDN3UxwlDuaSkRJCU8/wILVA6ilvOhVBKcT
1EO1x8ZnlwdMtwOeKpNIH97j9HAZniDJwh9xvTF+ePWQkCTmvdm9uli2krodKuKNwbzl9J4WmXnY
6sFwYErgiHAc2au7kkXCmdwRHBwLS/1Ks1oQh8VS1f6jDbnAV06S30Dklk56dcyxIIjfWiycDFIH
U6QfPW26nyJfMrQxw7LkIkL5DzatfcjeaHMoTLHJOksjrPUebWid9uNwlsCsZkTM0ftlNJy6Q6UZ
YUGeBhl5z4tqAqc4nZOPUpPvcllBFRVOZ/adLTQ+l9IRlLsbzWHyJ3r2mSQJ0y2dnIk6v7ZNTM78
+grn7ltXUzmwwksnyTcgYXyCNF56zGYCufJwxi/DHB5RZDgGenGs5UMR7IfK/1NPBRqeZdr1G1p8
Pm3gz32UKVrKJ3+lZcjxnzbjZVImbapKIi874s9lbLM68cLDaxzBOCuPC2jDIixTt42ocWPkDhEC
PXTR+ufw33zxJWLG/6b8++riRkbWgGlxYmd15KlNDlL2iMifLi4hn6nTpxNzvbXMAOBH8ZdAKmU+
YGKQuvzcXMAIzZ2IlKZsCXkVTbgIYSqvUra9F911z2rpbPM7e74hBwuAtvCX5Pv04xHWaYV9gO0L
sVqj03VbQo4tB7iT9zEW19z3zKLtjIGr/ZcJHKS9rpyANBu0OnNoSykJvyRdNTV0MjnpY2Vthzhx
lxAyPF9tlMI5dge25w2pPHK5lmfXJl8vEe/jZNvAeJ3KQjqPinNiSZlXLCgFR8dZHJPzAud3dHl/
sRc3yZ8Nn9stGfj4D6QOeTBQE4AkAnztkGhyYInMg3xvhKrV3amkcLvQ+un4XmeA4LDWQUw4NhEO
cOsp6asHuzXvzjlQiNTjqdTBiqVscqnqtQpz2ND8jpnYFq+VgZ7ou5R1Bd0j2u8vlCl7mjPvHEJK
EQKTDw7aGa5O3R/ueZac+heM4QxrGNQCod8DBFrBj0vmM3D+jqo4tmGQeMAn8YPsio5TqfNJtDIg
4ifZaGSFC42FA1QfoPyWGC/Tyma1TN7PQR9QzoN1/jm3QhuuRL2BV51m8I7mH2d74MecwrLyOyHj
JtLmSoUBOGyg4upvgXPZ+f+wBzR5BV/BiC2u+3df6vdxGF5st120bbk5f2a2bpexNkhdFVVfhjTc
8gFlNpXXBisWaVzCBuQAezOoJCGUOQ+qVMQi4FPDEEjMrw4G3dAtiAjnG3yvZe0oSqr//mnYLOtv
J2MYAKOUz246w5DajTnt+DiJqlSKVkgx6GZR7MfS68IbvIeb1Q7tmlnNY+iC5gxp709Lp8cd0H5T
0Gs198HubW/y2Fg7KEgLRfTigQd5UxCRQwOInZv6+FT5c9RzD15gbbBRbo62vj2fvZASm1HaEX0I
l5C2p38gdegTQV43MkeqlDxCTVundZkq5mUqktjFiq9YmN19fgIrEuQxKDixPOPi+m7OIcj+S3S0
dxjBs9ArW3q9KLk2whv56P50sm2cILuyxh2Tqy1Op8Okk+hhsie/r43BeXRo1fu08gUPfej79CuN
/R+Jniz0E1q/y7KjUw+aRUSp8Uh/7Ny9Wc2K+/VzeJgKB00UTCDk5+VwYLrHSiL8TGiVLdelAFI9
4J6iDVmM3k2sK7OnfFkj0QAsB9/ZIaWxUmUgO1SnoQJAdvoemam2hk1Uim2bU6pm04ipodiXXFk5
Zyxo5vKw7Y4CNHT4pzhC0VzxlHnBOu1bXNnFyaOtv77k6G1KY9VCQVzZdvlHT5pxC9h7ghHbhs1v
pHvxq65k30pCSXEz+KZI/SyufLqPM4JvhZAtR4JroSCTKlrfdWgGF1z+RCoYcailPqh1IfXd6lE7
2prrE8FLUejo7JI/ZTI/c6Pd96k1uSJocaSjdF5wkM7w2iGY57UzpKqH9v0On1Fnq3EmX90OJf0z
YJ+W1D0XnfJac9dPcAXBm6/KgOjI+/fFUN9qkLg6u1c1Tq3gvhS2vdzbHZCpvYaPmyfudiyUUbII
vWOAJGHfGGuNQFc3m+QEFHP/9FCBEyY7YK1pwkDlN3NydkYckmrQzcQyqTX721Rajwgq5/nEQ+E1
ey7S/DydGlWCstSyL4490yT1eXlf5epHyFpDZkwWNs/LnxMRqdaVNquwTPWAcodaVYaizh0qxLrq
kbwQMshBXWyRlKFA0+dZQpSqLg8Sw9d4WZQPIPExgOfH7tPhdEbDLts7cyc4BG5SJLsvuf09XZW5
q8zLWSRfpVcANMwAXh+jGhtOors+3T6eQ2qiPoTxKmLaNWKBuNgGwFis6vkc8RxWh5BzWzytO+QL
LaouKv+FLPcsSedec1onH5mrdT9CsBuFiKjOPAu/KpnzlQhDKpUwhr21LcJa/HsdIwOye/nCtPrA
jpK13QwTLQV8ge9c+eEIyGnB/qHDZZ82LzE82G5NCApgUDWIlxg7SxrXbJAl4n69d/KZQD2i3AlP
fbhQJfGXXu5st9mpeGMJpETM0FM3XtVjeLVp+i7+YgqEcWhUaTj/VBjAGhCrLQEUlc0YE1X3Er40
7eCg4pX2L2OxA1BYKrnuEwKuoJ/Fb+6AzY11hkpUTo2b8OZc1G6z03/KVPOzromVIOjJLmnUoXh3
IVg8AOS+0U6uYWgC/n5L0AUAta5sh7aCM/3J1CQGFmWiYKx4EqjJxUyJJDZs5rSOucvoswK33fty
DsqydCOMizwtXq7I4Wrgm5yJfEoAqGXRkgF5DU4Dvtinw42wgbuoii9R6ymcJZ8aNLRamBuclC2M
qQZWSaAqkVTaKwXaklYIBNKGMUuNACt2W5cjR5t2VSAr2Xct7KGtvuM03PmZmkqR1dZ3/MQNUGjh
+B+FS/C1C60HtdSX8V6sSUiJ2GGrY615d+GfikZ4NqTHBw8ZoCF4RuwN8r9KFL8nFoWZlqCJBBAx
6jO6+g+zS2k3yUrnq3JMU3mczKisssK8E7XqUsgAfT60WE3EFeN6FyHHQ4eT6KRFA56zz3gUNNzx
diXkMJP6AtFqU/8m/Fy3y69qJh/vZKi/NjcufqIWHJbKiP4wCxFzL+BZ6Z2dFtJ81psP3qwc0NVH
H/wePamRDqXXwqTkB3vGl6ql/YEu+yjNTzwhPhQZszsg4RiNYQEZ9XdVxM5KUjk16Mt5/awcTtfV
HzWSEOHEr+3oYQmUtQeeIkDm1OaZ4mqgf4CSe8PuvPnHyMakEcKs+snV2V+svYlnf/+1514rn7YX
zOo8GzNViUYU2hze8ZJfzH3f5ZzZyVspIVKpv++DF3KA/mMEMZnZc/w5wBIwpfQ6xfQ3Y9wNFnF2
+JA72n6wfIWwy2XnwCWl9v07hFrb9KPXDHwdzz/zReJmlS8vs+FhP9gb/kixhUw7XGdSWn9Ok/zY
e3xN4/NdSD+LmGxZ/kXsrL4uaiMo7kQ+EnsCSn7+1E5B+yDdiP1SpkY0rlEi0z5t7iEwbj774RND
h0Bqt4QMA9eJvvE7tIlj5NJxFex89y+K2rqcp8TEp4fdA/t1yc6eSLgbiNVajYuaEFABhPC+lw8+
2Gi3T8wuFuhq0eiTyUOhQ9vQkbFzBOxcmB6Bwgbd/LPLcQda91UeuStpGwP0i9plbT6gOhcSQhmn
IEMB/9oqZkjdbalTLwHR1lVz2qCUJYW1I2ZCaN6bOs3Quvws9R0Y6lOJsFU9uj/AAmAzcipfnx5V
knKl/kyvunP1PQ0YDlDIXmptIRCZp5U9IgCJ9TwCl72vZV6Lk3AYP/0GoSme2UZBU0GHArUFy0ig
GJ8VBynN+IBQTJwG6mNbAfFDjhZu0NxXmOwiz0C7fc1ksNrZsg81eEchOGt7RYyQhFN2qhlL/toh
UL8N93o9eOgCBQxu18Lw/kdblTRklHzqlbcLdur0dY2sunnnsyvV4OHPHawexJ5PfahnBU4Ymx4z
eO5/+de4yj+ZiLj8PdgsIz2Yg13xfSqvk4PhCyzQOEyo98TX8RUvjF3ej4tZ3i7xrCSzhnoKmQK6
Z46d26C0FLLpRptNfzVWvKkmc1GRqrjzynj9R4vNNi7FWof04EYw8MDLXN8lH9O0vlR/6ozejZv8
ewFjAyD4j8frhmj1N7rnV5czxlRVYPxj9/L6AJf7lwWTxPb0zD1zshZ7BJ50xY9Mf2Fi+o5EvqTm
tg3y4RWDNCbPgEjM2bF8wLHTN0qVtKwYqtNega7WxbZMwImGQHHzQMeG+j7TxJEx6lyBu/IVrVif
elSjclY1qwu8lh7ed4IRX/GB1T/QVNqpXddC4ca7UImVtKXdcVm/QRvd+w4+Ma5/Uj9YEPnRbDfW
hrzOv/l4uZzWmTtasNb+xeyC7N/kHl021iikkPckyw5lL6M3b5y7JlWfxdS+I2CkvXELNJuPrWXD
aQZJfDx6zhxkd/ER5oMQ01lPPFKT8r+TDV65DwgpLkEWU8L4tpp+35C8DZyoMbL/7ZZeOGmYItAU
JT8PWW6usSGsglHXggAWXJlq0xKAnDu6XDhluKEe7DJvPPeuopTzyKklG5ZiWHHBQsteg+uCKSSI
5sIAuuOAxawEi9KLiv6kFKf8UeKJmyK/rRCwFOA1Zz8tYihJEt9KppW/fcP0nklofDtVJdRAY4BT
pjTcLa8Al6WF74eRqUAWIH/i1lXOX8cgAJaIlB4BxrH30Ik6qFC+5SA3/LdBZDO0RmrzcrbxLAnx
4kk3xjQWy6vPvkjx6wnqCWY9viNi9XhRQcvDarR7OD3Hf6/zJMH28xjdWo++C6secMVh4qtsJDmQ
pY03mDGfGogKgI7STDp4OUneMJ+XvBQQ3el8WiCDuMmLsqDzyRm6tk4bkcgw+DySTqblbCvH9rl9
3Xddj6jHmERE+Ee2OFBhb/bdJ4QO4Xce/7yZKpcEy4wJ7IzJy7e2RK0lX65lK8XHcGIxgT7+lra1
fDYb1CCH8m+aMbx1Z6hHxu4fmHrjesVHCB4qpjxqnj0qKPMOrWAYxjZkqO1PS6QjsDXL7r5KANf9
CM7rjMNmf3qjZeOQL/g2VGtJ0uqsbg77dQSwl217bihW8cLSt7Vvsb+S+vAoYIvotPhK4qzPXda2
xup/dxDnhrAHuStb+hOIvfHEYyEXVBJE78oTqmXnnO87GZCPBndrOPT9D04byQZYAJRSYqQb5G24
4whIU1lW4fK2bZAXKdVNIXVsOboLt0qx0IywGqUMCHh0s97INCzo+I4MWF4u6P+uSvAwb8ApM55f
17VteZt700teWQ0hodo8N/kcynzQczN1EfsMu/4WjBuIPKYQd+Jgf3mvk3A2LKns396cTQB43fKt
wqolUrR3pVvTBtKF69AxPKJFOeAWo9OS9w9b0SCQwZwghc6rK49uwV239AdgKRs4iC4CtSeaYSZI
4ZtuYcpUAsC6LvBqGfJBbPRmmsyKMbrbZkXeg4hRwzauvaq+JzjmDUVd5KOs4kTNgnz7q8H2CbYL
nwsPt2+JOx4zJICr3AiK3DcM2OnTR67LR4kpD6Tb6bKeaCk5rWuNzWKzQsfvnn6cKGjdBl2ZAmas
U3YmdifQrQoCziYM0fGGxl6eO97M7R3GAG0Qgrocl6rnk93QAYXslA9LkcMGK4z4CIritPVKMLDN
dgTPSXB3tlichua5u0gmPP36qMNyytz1YTiW2x2UXU/AMCX9iIkCUtVqIYXUrxjhRfy+id6eVLNN
gkDyamGbl3IZhwrcYaOKg+8TVlCVT8WB5jx08UQGJUhkq0nH4GRThjp8o6k2fiN+R1zuEL/7WaYQ
V/Xr56mShMZGVdKnzkWVNHJo24+uMgVj/XOi1relwvdqS0K6YlSLsJiEmprJDjkUQ3WEUiMRcxqq
HjtOvJkYd9oKLE17Vngs/kejjcl2MYEgtAAGNkvBhPA7ZaXAGjGBYMQmkyMzgLZJEqEZ27afebdq
jUK3f5MdkDGaSZ0GEO8+SplTu9au7eGZIztg59e+svFok/iwVweHCAES7ue1d43tvILGHlhT9sEo
SSGeW2D7DjrM0Q4rBq3xnPn567X7FSs6srk/RjpczTH674RgFkUx+xeyzg6Sl5wt8pECsolUTEP2
tFm+5K6tIbtfNkoyKOynInR1OgHZthmLi2+vY1J7VYAvg2K5HLzV73Vs68zqI1bnXwJmt1wuvnsF
CHg0zwZJJtbgiJzSbGv/LO+DGW4mCsTtzJyrUmr+zux9F25ZBzpaTOgYABYAVLTOJcwhVr7Dlze7
FHszL7bWL9iHqBrodazy/BlLpD7JDzMm7zseKT6koLhQH58m1yw14S7DK4XvYDpCXcY2KQ2Ig9gH
P5JMScL/77u2QHb1PJsB4V+r6zJSqo4F4fWQPWm+aK43e87kV7Z9ZgyZrwsjdXujYKejPF0teeky
89mcOsmQO9Plx+fkbnQb/4mbjd6BobVzbWJCL7+aIVCxMSBLdC5P+4M8J+tiSJQ0DX7qzH6Ogt0w
v3wVEhWxwjyAbBUSu97OWYy38cEF76P2798yKKKwz+8mXG1aXEf7RM+5d4OSZms4akSbrpJRGr3H
Dy/3IhvI7yQY7iYZnPoqYMFaH4ZrdNeAG8y9tK3ngjfhiM9k02VZDm7sDlTc9+y8e3YHWuyideIA
1L2UQujRq4mo2YrtSe5C1AhzPLzddX6PFp0VrgYF7Js4w/nBt+X9MUt/QMhmi2aq6JQacxSLli/7
6Lhp8XP5pT6/AZM4dRRYchz8acOzCaf/R1T5Aftxzs0d9MHI/uaYq61m6FeSd4RMWPKqtB0n4seQ
rDb0Dp9+OpXe35TlqEbEAjpEw3MRTCDeAZyK2wOwBkzQrsQMOLp8c+8KXikBQznPFAhnI+fNJsiO
5PViFESmg/yer/+XSsRAlC3eOPwODLH8HEu9fhxJMveIcglB+xcKTrjR/vM0CEtuYju9ujrVgMTG
V9/GAtcNer0M6ghj9Dg6YWYq6BdO+jQBdyogBOiSLZbOWYPDz44HFOllREczDlm+DEMaNuPZwsbT
Bz5XUt5yVG/WJbI+QXFluGksjgU8qC1sRFofovryLJ3t/ZOdD1RAMEtD7YWB7ro+f7tL/vMrfyeI
KRHBvyJWE3yfI2O+oiyIlX3oGPKaLUdJELfsHDyjfa9IQckl/dyXkzhE3bOuOB+n/0Wa3sK9q0mi
rHljrblozgbJ0PXHTYdamtkC1qTRfwhHwjhlTiTE/ZtegEFWuaYDsorU77l86V0b7EiwG9NrXOiv
nQoZySHFmMPQRIk54ZYSJlxFjpOLmkc+3BvzroRri99Lyp1jEAOxmwEWI5LhP1Q8SqH81b6cqquN
HCvLs7L08bnb0S5tOZcgD8//Gu0gH/c7iIRc267KfmFy6eZa1HkvKNXnuNxub3Q+E6a+lYZk9FGx
i2noGdpTxZzLhNyfBCnF4fxLu7Cd1CBcI0kIkR/q3jqrAVQJHUYciJIOGHdH7bc4RnRMdCb2xTKs
VMSAxwZu281qJGrmxncYFqpgf7oNG9PSVL5ayxbIkbBJMV1Ah6cQMvvjgQjtFfHKLjthGkrtdnPn
ojsp6JMQR9ba5BPiIOdofNeZg8JmjSGd2eGbt3G6MfOGEWzdbcf0Dhn3E/Y0IYblFEnfk5+gw4TG
vE7585U74XhkpxsEnpg8Y1MHGHMcEaDJ90A7uGlJhUS1NX4YIop/3BzP6HcpmMbbVoD+Bo1ZLgu/
NX5W+jW3AeiYweXi7TqFSRdh2J+XnojNquuqBog37aUI7otFDt1KLvxGoHOjs/x+BxMw1gN4fnP+
pyJyVxpj5m0mRGEs0ZIf2UhiOT08ikInrQgviy/KUGbehk4/N7rMMf0JrA/D4IYJwD/Nb1FpUxzg
Lde4a+blZikoS4BFeJlVPBgvNfI1hOmK2YGn4g3aZ+ILRt8UGKpSUe5Mo5aCSrSfc0emUYCHssuB
F1apFWfmCLX9necETChisxEQsnLgJY2hZ4jxfhbVaAtP6JckVzNlWsHEvIctpEBmffalS80FCOLX
5OcVQ3dgK2gSCBnVwnwsCUDaHw7AZaa7O7y9BOOp9Z5UHMb2VousZJxrC8oWuGlOj773/odNA3o3
b6AS84DcYsHRP2AHww3HenyXP/fVbByz/VlgEetLlHd3sbtDZpEg8JCg91iQAxLZaggiRCGlM+H5
3JNu4671gNW0vzXKMmpAkzqlOcV2FnVnHQcYQy/pR0w9fGV63n/yDWWbwraoTICOxn9kylBfEIl6
xlCWr/U4r/whqcNR2irnquMq1wrPmTKkLgrhjxb7xzb3JLqk6wVLYb0/46NmzeH1V/YSbUiasZjH
DtpW1QnP8DUEa7olh0IajjxQQAWTqihP+Inhse9jxW5XXpMrbHTL8V8xDOxaWpw0Z5Xmsu+Rgunu
GSJesn4VyHkHRrBwO9dHlpOt4S5SwkkbJKC0DFYgK8zLqH9O11qI2vXRXqHitPMVEN5Qo6gr9s05
6/k/Wr308TD1YHjLC5lBFMqReu2V+84h0+7fBFFYX6lzQ+bslYLXsYP0nL0eXYDKnr7ITlimx35Y
Zk5qJcUyYPT+3gRlvwXnYQRlywsBxNFokt3TNB0Fpxw2X/c0r4bHM5hy6wUm2AjDDInNf80DV/yG
3phrKcHKkMxgcQ/qR4nADmlkk/EWnX/1oPbzQnP6ypGNdbIkcX5UuqRwC1lavRGBlpY83hdq4w64
f77AHfNCZbTdGlhXOYP+zlEEKBvPIjMfl6231UInzbhXlzCLBYfD1tJuV+spJYPHzSiR3yRiR4Jx
bXXpjc11amNE26Dr61K9m1Q3FsDpnaLeHAP1U/Qbnx+WEwLdxD/Cc1GgNxVfM8O0gOyw9CWT9sKy
5zkl4D/aUKi5HliK2RqCGC/tr0lYjtxdBr4AMEtX5bde/ZXT2VCH7zgxdeUyLaXlOoryp0CBknF6
v+wN7TyENLj8w1U2j9SiAVyTObQ5betvGTL3hpYciNYBCy/jOohRZm3MQbcwOYMXchRu5uKTmfYQ
Js6vF2CZVIxg4o8PT4I6P80GglIjx2WO7kEjkLdP3KmvXLT67YvUfT/MPaiTSEbuUfR/FKSKstUl
0RKGi7+f4kUncz/+f+cFNZn2yZRNGRf4BStCMBj6MkZx71kKE6gZWiXSRoE0rg1ixz65qJ0zqsFQ
9td6nKSpYUu15Mwzx5tcNe8qP9gBZkluwraimT/TshrEZufykPGxeM7+U0cNpbAnTrIesGrOHFfF
M2s1TIOsU82HxfHZcRbSPhWzjlkHVrYyTuHPq0E8OlUa7lNFnmWb7/t5+dOf3SI5Xpm/vZ4l1ZEG
VS2vaFeAqb/SaNjxAb3WlJpRZOZc4sBSfxPXUydpEK/fzrAqo4EGSacVFsvnrPTJyxpxAaFrIDtd
VfIec9sqzgClQpRsWNtIq9xBFIXwMcOnzen0tLXP/buKMqaWqqaoomF/DmSlzHc17zVlOdgfbOzW
KBzwOAtSnoiwabL61Ni/p2Joqn+LqpJg7nWD0v/ayHvghaX//LgmgFpTRlZpf0Hv4TN3kuLwfpaN
a7nu1j9laH+FBJO0ONlZ8dOMOjVpaP7vrOsOs2kIzcFw/Z/WKLb8uKJyVD+MzypgBE81fORfGomS
hSjrl4WpQ5K1EZuv4vl8AN+ysJotgZGHEOTAj+E/79qZvriFvIjFYSNCKT7G6tgo0Kllz925nkZj
YiGxCkjB85JDR7NzKnyc20GHQ8rirErj+o15YqTLrd00shF1nHZK4fugNuawl7OqTHLxAK42aYEb
rConljcwBjFQkFZlAC1u7wnka5iEMYGUTRn6s8EP1tlRKB/z0KKGvGwqmVRP0h+I35Vk4D2tp+HZ
EHCO4Nvh/L9dJI/a1md1phq5buPNV3XkBSzEKc8Q/jPFsdYvgmyGU8aX9iheB/lh5Ypa0GC4FMBs
xvFi9ticpLrMblk6Asneqow37YUgOL4tpOHL3pFN3ejpHFp2SfBlA9cDS9/MCXT+NjUwV2meouru
w2sEQN0wyIsFGQEfZLNGXf/MWwq5GYk8HkfiIMSWsWtbH7oNXAdXiWHiRJf4mLmsDqBWxxmNuqXS
ZrP8/Gj8FhH0MA8NQH1uygL63MwaOoJrRpAmBhzU45s+alzwOyDvJzxj3as/2HMia5Xh2C2v2E/n
85Hi800sFnqgrl5oRkjCkGt/vPtayynKnfF/BDX+ncvC7ct4gHtoMnOVS8bnFx8MKMVbrul7BuKZ
6GX1l7Ph+83vogFnrrVihpUryqc+m9jkM8aDGVvLy+FY77BLN1rlNuiTU8WEZH3MoUcCpg+SF4b+
g+/yJrmyXTIhAS2h/TzBUJnh2W96bdVbDSFBE/MYomrm9GRKRlIZHylMWl3cSlGHkv2f+xM42vkG
JNjLcCdQwgfRvkkbB400j4iqgI8pseNFwEzEJP7I7oLQ1Bjw3PQxP8jGElOSxh1E7ZD0lYtRU0hm
zfy77l0LvnV2rQkyS7vIzvkHfy7LQiQoat4aZBvnj4Z9xNo85KGxMW1broftIDOOHYQtySDyuVem
Ws8QP29Z1K5MtcOdPx5asX685SxT+UaWDS/Kqmlc2bp9QSIJ1CbblSKGrtIi8XJZiDC0PTNq9DMZ
DBy4i8aYv8aci5EOtpZ2wQ/T3DbZla/5uSHkR+0kT9gmFY5oRipTxNBm+nU9yEYIfHcJTJhqJo5k
oYjDhooMHe/VBdOGhODgaYE25Q/XYQ9F3BZu6c1hMfPG0k9l7TWb3JMjuc+scBK9qtWHAgqM6qKK
MX9GfZIle8ykmcOVIoWhXRKr/S2QmoOqK/hjVjQyPhEHKxOigUvF8O59qQ7ppoTxV8P5uSfaLhHV
7magvtoRipq6P/em32m82pDEQRCiUEg03JL13+OLnR9hDWG9CocOKnKArstsOpIwomtmFIiXf8sJ
+20XCsRlHxBjgWEPE9kG7GR/tQjo5RLOBqFeHfeS0lWG+i1p9VXj/Pum5ZHe6s3pbPw7AdgOtad+
jxOGX71QWaJ2gqATfF9Am8afOsfiuat81EYZ5eb+G/sWNsNXpqpnpFg25qTB+fmdNtcQzRV1FBnR
/gJwDaV3TkUC7l2zJMVpOZw1W371W2D3FrkP93/oPQTWH4t+AGl8QTCUCVzDp+tGbgRsiHo8uR+Z
W83R962ni1vpfKhlsZKq2cZZo5aSySO5guVFAM2hsFUkYWU6kbvAtsASnvqba0k1Hq/56lB+QAUa
Nf0ylduSPTXCSfi/3A4fXazU5Wi9g3v6720ZVG7A1nGJU52TRcScohlyEG3LuyFbopDryNd65QHo
5cY+23ChTnC2QyLdZ5rirLR4Vma0oayDuDYw2TdodvinMPCflaHrE9Vy2ESS2VboM1beRv7YqrP6
hhoSSR/JHVmrCLqm43Izxa5v4zuVytBAOlc8sYhVJ9tv3nQbMqoJ0blP8VcO5Q1YKzcdyizv9EWd
Ye+s8AHChWYStzu1Dnm258Jc94x2yAcQgJ8UItC4adeJh+EZ+OL+cRqH9X+mWoggr85Qjoo/V1l8
PNfTmHAAyAprUpYSEk/RQw59LayoVVbHiUcDIBc1VBW0p3KOrfzzUqmdcb+QQVunB0WUorZgkbzh
kX1tdDnZAQhqXVPJGrfNJm62adxDg3W8cKf0YYgQ6gUtY8mkNN0s3DRcBWXb62gsLS95HKokkNqq
et+7bSylT00xwyEq9AjqXZoWPQzkSX0u8oPwRqr6MlocCx9ROpnp0D4QHyHUCPypNZ32eZXSyPUG
Kf7I6up75dGCdTMQEIxLZxCheDsi+6WuD1SF4BopDOsmspfpJQhlhWCYdboA5cU4xjNLjXngcVbP
II5OYKaaWdrmq5AeZXyknZTap0zoMnARwRlH4JzfnDzeZ3mK6GzcRPUXzO/gMd9z6up8mYAYpdmm
gylZWpSh8RoE8uOQHQcD5CWCs9S9cnf1dICK+LETk35wcP4Jw4tJif2+bqn9aHwGPbFx/MkH3gJs
8BuSwKC6DBModHXWoU2Z6/valNpxzyDMUp2e9rz/iD254FZtJoIsUEZB8EzDz5lYFak+SPKrnlBg
2oiUQyJPw5HZQv+jRjHsIzbDMgtu8TR8VURWDc/aAIkLhXX6I1phbm+kr4+vGlUqtJqTJisp9c4I
QAd5zNPlcgAVfxiP0mMmlqIbt1NRTvDemkbgEs5GoHZ5B1mcEhViR/9uPYpCQg1ZmguzhV2oFsPn
ud5bhkbfiTmxZn86hzyWeWngJhlzTD3/j1tnKyBUF12W11wd+p+AVhHlaTptq17Wn8nJTGYQiF0t
LIxDvWGQtw/O+D9jYwKrV3HqYGP1LICo5fA83abEc3oEV3UMVYdUdGFTgcu9UUhPx6XnPn4EJsHr
jFbP6BLa7vTXUmz+dIvO3pfJv4ZGHV1bXFOIbesbe0ywxESdfE8USi3R9SXNwKSWq58UvHJneTpG
EVP2DXzvGbLVLhvCHVosG/pXelfVoicPkEFxITBAJ1XoTDwaQzJ/9f/x6AE1USft8iTO8f7PILt/
nRseiCfjcqPhIoywgR+e70EOrn0Fze5ImevR6MP2QJOV4bzYzqyHJSeuAzQRZiwo0/HqlBN8kNZa
gmgeNlcDE3PtNIrEB66HP3z3EY/J75tBbqjq4pD8VjhGGK61Fl5MTQrEajpFEBOMBh3RK9r4OwvZ
gERRB0V6FHABif4aZP2S6xH8ACy4li0Zb1URk9LBiF2gqLfPYaW68fQasWmJ9MZNYDsGeD/duNOk
uUYwkCKNtcN40uouUzRoVT1DSWzrIkWLfVkPHa32zvxPCOd7k4msF3zePaZg1sF+jUbgivk9fATt
5L3tsnwhLBUZ61mJMfqgvfQsFpSXqJFUr3dZa9UpQ/1KuMVhJhgbLQ/nAjLaYc3DpHyTvB14na+Y
PLuTqVnacwk+vzRPlCHicvZFM6zICUiKcvSlEWBDb2+Dk9yymhCBEz9iNoSZtMb6hroY3Mc82EhO
V5SSSbHfq7YXxxzxsJ+sNmNgBds2yICuWn8q3OzC38pBPdFJogmQjgYd+6Ti6l6U5uWDEvCROCyC
rbWjPYalzGm8zH1tI8tA2dbnCdJbzpChC8HtBcf1a7MlXJtTYMvycTpr7Rqx4Y57LUD9fX69wmy8
68XUNNERBXxrNH6cjiUWi96Yv10/u/0LS4zazorZij2Q2fCOwzEMerXYwoUnTG7tdSolXKhhXi6X
xlYR4AFsV+1Z7fL7vJ3vQhacVbQjqJEwhvSY8Boj01B5CafSZDd1dpyQmQ60PlbfJ6e9oCA3MUs+
F9HYH8SknRkJcjnFucOGRzR+sJBKLkJca8sa0EbhqCR+xUcHieRhg0HB/3dKRUw+SoebDUkKMv6F
FlhRKaF/we+fgQVmk7vfnzpN/NXCys9nl3Bc4cj2uv5ufTrys1unhKEG9l0kX8mkg8omPp7INzsq
k0sEKPW0uIHmITQhWMb1q0lSRMCgmABy5/HjRi8eK+5ZrlwqmmHSCL9q7D5o/IW93oT/dg5/1HRD
zmx9sxP8iiUJ82ez4Id7Dj68a1XExXR4XwnJW7KdGTqFa3itkdeOQBlJi8focV7ldprRf7/C51l2
oZNEefAj8nOhzEtZA/dJESu3GdqHO8LELTkqjgol0Q22UBjKIMzCJkbGPe179aP9TSWOYDYbCtXI
QVyJIivPXkUmaPXJnqDW1gywRFZRLLyYrG9nmVywg2qh+YmCv4OQYsWsrE/xlFNFZqNVoinIHsdJ
FHaB0NC50nLwJznk/b6ylUDwimWuEwaHi04rwTVD+qF9p9HQwGjjekRvrm9jqt+PqkFQsXB6UpDx
8zgHcbYo5hDulDjChl0ufOnpXw285XMXSValg3JgE65qOJJ9skXzGsIz5HVik6N5/WWFs69Je2Um
CBYF7SiDPhiIL2RK5LEo01I2HOoWTd3PEi1IObV+DfwhBtBj1TJfWcZfNjcKxABplT7kg/0An4+8
G2IlLXp0LAA1x14IQMWjsNIibLT+WsIIjZeDrjyjigSQps2R8EBV0SN7dFEInPrBL7PyK2tEV70C
dPpSg5XROxDph1VOFB0YxioxyKph4kD0Zl+SZicg3CmRSeCZ7ID/uKwQ4Bh4mEMHZD37dP2Nb4VE
+lPJOMxOVBjRDERmRkOi9bm2eYpSDeOxAW63xXcbUBkidKYLAoNEjMHGm9FdkBkYubKobJoEMiNk
YIZFle3ouUOxELDJ++C0x642qJKCdZnIUcN96Je6I0+2wjvS5TqG2Qb0kHbRdvVJ9cq0V2R8017k
QcqWRfXIgGPMRq/OJFaxhd4L7z5pCcm5MPOPEefRQ9nJPW1KeWCXhuCLZzRT1qfkjBMVsNZAbLvQ
dnHmC7psH6eEfQVeQJKE/B1OHcKVF1ygc5cBZfnqm6q9hpa2KNYQcNHIN44wHJcLwpr7rCf59nWT
G3ZVutnse/jxb9vlvr88S86+1db2Tr04Jbb5NuikPfHLVPJQv/x+kxleXzlFY31utZcCBxfQ16xc
zpqLE25IDVmH0sRHgMSfvCRHPghXNFZs8MgoYeD0WFmcvLUALHzELdeel6j4Ij8V794xAX0OgRZC
MnIemXZjHtI9Enqul2S6lLJnzTzMOo9wPz9SUyRqvIBMvCqlyFe/IsHTt8WCtMwww0TLUy+2ZTQL
vRF/2RoTga2eJl9P9t4HvFHTRdifaS0xvXz/rF3U4vGnGWemQe4i0nG9LiXI19Ln+rwVGb9r60TM
13eUB4d7q42BzHMxlWltrIhdT0W5vyUnyTpJIm2aFwFJOJ/2CDBIQdWnqZIStedX3VxSIJY7dsb7
vHbojox8qqlDY3Pk4WNJJas69sHGn3hS2qowGkmw8yoz0GwdyqTvmBXFhKbLRIf2e68UUTn5bJq0
f9TlVFmuy9AbZe2idNJt8pEozVQbi5BngFuRlFTtruo7dmRLQEiPmzzf0AR3Vn9NrnwtzJQYouHp
RJ57DoYM010NnF/egc7aZmL79RMl+AWW6HQWrkYe38ynVNctryCsnS2Kb0BcxG5y+sMYlz10gs5y
PzV9jQOnMy1zEbFBEMdcQvbPDBmrK2d7SZXoRfMMBQBeR9GZu6pcLc38CZ7ya04kYT805k3BASmK
Ums5qWer/9aT9rFpwJsvyz5pF5XL8MxIcrdBLtrdUQTTBkYDpDKIZohiK59BeWvtuvcF53sMQf69
GKmqQdgg4iAkoOEdzCym6JoQdaNn1vFsBjQIFONStWIlxsGBUvvKrgOpfccBcKPnl9IGHmDa+txl
uanbKg/BvqF+3Jr3Lqjt3W/ugBymB7IfXeAk4p//0eLRRHccrKGfmcHqfr/AB4vBa94TJJT27IB6
4aVA2ltBKN6Frr9TAzAJACi5XnvAxUffOCPDU+0orMoiSVxTn5T2LEnS7teAWmfpf/f+uorZPImy
kR0CSyd4HlQ3iGIZrA1Sy0jhwszJQ280Q+Wy3U/2+Yzemoe7OPrn6IUnYvqVmapUDVzZFJEaECAI
jnE0JrJZyBMMaYlr+pwHciHIPIsuWyf9ZHis6NjVieuczSmsO0LVPbFq5pYu2F22ZGVflWAhqOCR
xX8b4wF/xI/qB5a2+S1wihayFUS/qnXn3OjlTTtshOGjD9ypNa18FCR0ZDab0MSL7S8sQljPNOm7
LUynlLncUvJ11IuiX63Tba5UYbHiVhe/Av9CVtdUbulzSoqedgMdp6wym20JF1OfZ5985SMFXy83
nTbOUTJTxiexFzX/xbWUQ7QyNxFS3llynY0T3EmyKr4Cbw5qMM6nQkHS7+0b64QRQCUHhQyzTJMu
SHEVW8wflg+yJFwB3LN+W6Vow4OqurvPKuRdE6hrj75tVnjzOTfEFIrdz42+PT7RtPh/DxFPKU6C
03sJ0AQL6Y+o07+PhQWaBcMuRIT20qKFN9mKx9xk3IhoI0Oc7N0qrn+tClmiXVUasq378aPRPqu+
NabiS19eZ65aVo3GQ8zBPdv3u5HYO/M4MhhN0Gx2vcGhDIAzgkDbCZqcrrEdiv1ZEvcMgoGKorwi
/uc7pwhlkza8lWXVKG1kIDGMM3wuXBinFd7k9lg8SHCvh8qJAjdVC6OfR+3BcHKUgak3eTT230NL
ln/6M6+IBCuFteaqI5JmLo4+xopZDuiatPhZgg1RP8+MdD1XzgNGwOVwE6niTcS/XE19GGlmT1LD
y8XOQ9CKgy4bvnW/NSD5ybFifJaPTOqLoGtiDnkR8G6h+6CmLzfqrnI3eTIwu7njDqLWlr5pDed7
tNBKOsKfvtRhvKafZCF8rQEEfXpIYDRDFqgPERY7uJkvaGMMyHyAk2luMkrnO7tCosCSzZ0+7SFa
OIvXyv/59CVdhJUgN/7RlFVSU3EbJqN16J69OuamU2OYSZSpx3auUX8dlN1nRKLVWRXEfi+CIDUc
4u6lP2UI9WXMQKBCQmZj5ntZVTEBRPhQVYoALROHtzkrecZ5sbB6yyB4IsBwr7KBuf5wrKT4M9sI
OABifTE4VEfk6swp2nydc+PG4ZRyj1hCRd/LjIu7WvCl/BFysIxF0KXqr1VtUY7UJSBptlnXAYLf
6+gd7PHpiF6/BjUU8xQhUZnnl19+tSXb5RRmGa4sZWiMgmrZWH8IzkeLdgwQ++BGr4oY8tvdQK/v
6tvCyliB8dPBWrUxF09MHzYJKesp/GgDK1sKQmA/IEhYnmUCMI/ZPNiU18rKJ9mREAD4OdJHwi03
/ODV85lnBpQ62j8lfrLD+MlVEnMVzCECQpKIAEmToxlYZowVCkinYUn8bP2Ldxu2zSbosqFW99n0
/zi8Azh5HgBjQhQIh8G9jU55AfWZ+83kpHxvaTMiDuZ57056FFZRzbpNpHIJ0gCsMOJvtejrAj6J
IvbWFHezfWYBWzVjhcKf/UEhp5Q4qgQEo94pd46LUoqs4X4g87vHI2pNMhg6DOCPulcvpN24a7+8
taWNBBcgBOoBQSGUmJpdQAN3mdBUWrHVYhnVkDIhu9RjGGBb2LoHG7tWIjuml9ROnnxr1hM2rSqy
JLNPP4m2NtaX9HS9xqDUSSVAZRwYzOfm/6/fIz85Kgci6Q+Z5K3LjXV2q1miE/R/Q/2Z9Wovpe30
AXqSOByrFGHkeHsGgFSVSDf5gIZSyIr6yIOnP9f7IAzU7C96OiJqmM5lLOAbM5KfHnwbtzNdbZ69
fdy5hXim1C0Uky7Z1rTcxQHZFc1Nsl9MQxNQ+TxXsqJbP1d01bBPglmIcs+ZBXzSIQh6uc5NRhHS
/1Fs2JC4XEEFhO4BPk+3DXWWHtpojaRD/DKSh8YiACppBfL+OyMfURzJITb4t+LzCPq/VdTQjq63
6pFB93E445IMPk20cj1dLrUVS1DiB4X4wJrgzJVHAoRD3pxtuT0H3YoB56OfHvfkWubMKINahlq0
UvFTV0fOwq9V5enoMgSootke/3mV7Cn/QcpnDbUiOZ6ryPcydYFvNhuSRpWz3cAyg5jOtc8y+4Tt
XR/CW1Jn9zxzmFn4tU5cstlvhIpOZ1CFUNpPufFeGUTrK6W4/eTXzz/LDhBGt+JCSG/zHGX9k+iB
4Tgq1vKpv/i9NFC+lw9CqBzWlH0H0CHV9FvVRjBGe7AoAx5hIsszXTOuRDsILuQBwtnxgAV7zw+L
qiCKpZ+WdVEYcO670duZNo0jdLtKqs6UhC7ixzgcC4lLdNXi4/p1jJMgjrQWZwNIMEvvuSZcJ78Q
cf5HJPXEeLmdByyXHccpbniS+U5fnT61VUGlva2n12YHZpufFo8XGKe32Ioier9Go1Sat6pjVbe1
oTWee+0BPwIQOfHttyKlt3pZAkOOO8JJfp2kCCmL3qmxTD5l8g/l9bWgzfCsSAa1NbwmzgsKXe3V
oVO3wAH+NWzKEUHZ+k3mw0CgGmkgFLX1GozFdeJIQcpxr5BBo2O//eCAVKkIm5+rQ5T9EXXDpvTH
JHCCKlbb7Ix7MFxlYoNwvt8oTh01gtJ5NLRsWyR1BsDp7fxl+X76mh1Jo14V5KMFPIQWOLfiLHVD
Qpfdu291HYGH8BayR8iPxluB8dnCgrhdPE/c2NNeAM/+AnbJlITrDia9PVqTfIXhArkghRfObvBr
pklZlRw8pZYFXsdd3SaNwGiOOuYFaXhJ78kdYvKQe/Fr204EzjLtATUtT9Xg4i3JHxw5jLNH5fmt
09Xns+HTY8BfVx/PI3OdISf4JihrhfH3CXZQuPKYTjPPdh+RMoygtWa/Vni/hXjXuXCDXm+s3I2y
xInGLSkHjj2jfNXyO8QZRNpEguglNTYhU011dK/xeveAf4Fj8OV3kL615QRl6KiZ47ME5HFXHDcC
u53LoczNZkb9/cC24zuJrcxp4NzdhQXGUZHLFm6v5BG7/0btNCP7np3snVEzQsSppF1IGqVgQ4iQ
X1jXlwaAKljVIBMlJTVPDmA50OuL+mRLt9HdERV9xG1ao2sg4ueT2vKdqI1TwHrtdtOgJayh5byx
oAIly6xDibttdKt233g+kjEoqAWmAYQsQ3YvESxoJ2dgG+z1ClLnUzKXoVWEdIiBS/f8xKr1ZnkN
Rjt3HOXwMKaBC/gzkfsVpvX8PD1Cxw+hqT3nvFaJyrIUpX8vq8ye3ze/sDW9OtKRMoSYGgKd0UKB
oTEOitHkxraLRTtG8u0HfNgplLVqz5o3kv6VmgX3qfvUZ3Iemb42mjT258+qlL689fBm8zk1ypzQ
jk7SdDdiuRyXNIFeKTmhTs1pzHeNYNQ0CBL2nI1apqtlu+l4W7BF//B4Y5lKFT32EC8DZXkP8o5H
3X7WXqJONVlSbfCRfGeeaMvdGJb+0mes8BrnAf/2iEXT2MdwG6PRoytfA2noD1We6l/CxxfjBN3J
ak0D5HBkTQ7O/3zzGIudpmnkzZAf1G5twzqXMjAYhVm/6qh6gOmsIoVNhK4/mbQ2YGcyoV9Qyxz3
TvF5yLh5fYkGzhF50d8ypIIPYk7XQwLjRGk3LINfVzdF9M26uCK6fpUlPkDyFbifgvvSRXHUHATI
YrUxGApt5bPuz5dkptXLoW3TOQbI68knK6UiKf8nL3gGSDDIp1dRtVhviMcwoKiM1WFnccE56N7d
SmmFFrlk5O3l0niDp/37JYsWqja5NFpkc/1iZUtmwTIbSPioCZYW5+XC+qoon5D/xImuHaeO0e9E
3/FwrXzgSZ3g6PRri9cTLwQfEhWl42D/CvQWfgkdCe0C5JDmLW4YpQVTCRpDrgOUX32SB5MHpwFZ
s6pYPiw8jifkXlxYH/7efMVcLD/BI1aQum8evn77JJbgnuyAym1TMZWOqtChn8rPMzwnMOVPo1Gu
++DNNOiXT7UPm4A7ggu5MbflcArbwM/sQLbHXXzL/t8EKMPjw6qk5TMbQmF6ir3D96GTlcQAGtVD
GXrctS9Xf17Bpi+lH2IjYhgZQIh7TcR1DpE6vr8KZMEr6DI++lNRnA+0k3FrACL8pL/MO79f+hFS
/kqdsGsLR7MTxwVrT98I38BGtfUa9idYLBiKAe3hIw5zz7Hzv5AGNi6pbGoisF77LA/uu1YKBZ/P
Z6anAkZo8CZ8nFaAy4MUuqMGGMuHRmAKLc6f0aZfZ7C/0QZ/egrbXzZGXe3GSv6hLJ48ETu8gBGY
70kEE5bYYiufrv3bLXS678Y6TZvg8cOPMy03Fpn3qYxBMEeUwf/HS0fm8lgk55wOxtEAj8tyGHZv
ssI0opTGa+Y69afMuyUUdpHIHHvvMPJpyH/PU1HxAse3HK6sFUKnwskLlDNDAUw302Iw69l1bOcI
rqsTJ0RO1h5EBOivfeHYldhjZwENVa5QTkgwEO9uUQjXEE3+6HLfTGnyIECzyxycP7SqhJS9Fp6y
/yXm6u+T1aIRVLAjlbY6O1/+1UYKzWxnJc3eyA2gk2IsVlBf0D5b+yikObtUI76+FnFhIeH2yMRf
hoEtZUzhX3v8YLCZ4o9rEJSipXGYyrfELDolNkgHluP/tkF6bqUEMiYVEZ4JuOySBuP6+1CoJEaE
8KQcbTWPmnG8YG1R7ocf5QezhdHCGt/CjVLpu8UrtajhRX6ooZ2GdljKDGgGA94k9Linpc84Lsbo
twNhglPk5ResHI9MbgCz5BRz6FVXbdQli+swFa0aThzjqn8oLYs+ZTNFAdBKHGhuOr6d6VIeTYUf
6jbtaC5xqB0ypa9UI4bPjIH1lBON9tZ0wYPPIafIzFQM/s3F8OWkTIV8yuO0bTKd+HvBctQOLZIe
z0vhhgSlYiRd/FjYLDIllUgsF936tZQwijLh1bF8oF/X6nj/q+UWQ6m65EADwxF/jFA1jJQK1VXy
l2Wq4U13Rr4VZ4RLCP6CWy8utQ0b94VHp2JB11L9H6L3hqGQrtpqB2Zb5/lZJ8w5xj7xvGlvN/lx
5/1jeabPbCBZx064BsED+7psAQN2YlV5pFhNxRHdF4FQAQ1RRRdRbzOAm8G+GYlYokIXgaD9ObEe
7yY6ihJR07fSXZqWg7fa2OPjWdZZ6KKoaRRSURADkixbmtyLuGOhY5/ch/O1UWGhymcLfAFxVQhl
z4jDA5C853oybbAnhpSR86nHVd3DaDKL701WVwQD0JFM9clp+7/k5Vq40cNH6X88Q4casoUZsG+Y
fILzojqgAkZ9kuP/pJB0xLN0d5CZcDVyTk2Ou9h5Vp5I0T4t2Bhk6gQ4eEHZ/99pTyRea1MJXE0f
YwRVZ/kazeEna9o3FkXwu+Cftx1j6iblPhcM1o0pzgw9RPRDrpT4rYkk1NEK7e4aSRe/5vlAEUQC
wmzVmqBPTZL0I21jLtUILcnuVCgr2XY4sg8sSAfhxm9mUH6ThkX83OFGkCn72gzShcPb3ZbGs8FL
OSoEzIwRp+/9u9gtdCWkH0Khm0jZmCX3gPIAUI18gAX2HYRZtscf7TJkTF8uJEHVBbwSnog7CZi1
nA3SujIpLstzt752Z+mBl7TI3mAHVZsH8agb4rBNkRigYaGQwN8CIbuvFWrd7Q5YEcDEzPfOwOeo
mFbXBfHTjIM9BltS4lvLav5Pios28NPofElpEcxujAUkI1NZ010bjJe276zIPVr961w/z1HBvtjz
Kx0wZJgpl4U1dnPQyJiW4zgLujO4rzyx50cP5wtzMCu44Fjcl+9gmQuJhUuRVuTK36Yvl0kUhPof
Ljeo/KmPDMJSFEL2I5WCyuI7z0GJ3QZICdiKS9STPlV4JSoiKDdwUsh63AKzXSfpsybNIE0f00v8
EOcN+YztIB0D8F1Yh0+jG1e3UywTjmIulNXcPNevdKnOatC28eAkX0ZLbKXRFje9o/HU1zewbv1u
nch4deMupQzirA7Yaq0EDrYjddXVr1MyzBnbntYvoryg/utKkmbLMXCwkrczb0IXID1A2bXfOaYw
0OU5KnC2vY30WXgMFoZXEjunWd6NlubdoA3mnp3jg484XasjYQP5Dq7vLNtQWlRCTCB5fudCb3wI
2ONUXB48IBeS58nm8fQOv8V5hlS1yOSEP/p1dSGTx3HGk+A+ZH/qcL3up9AeTWtzj8K0Cx+lKh2F
ubfehaFGPOEc9W4iqUOxOy3UZdM6O6pjcqse1YPOE+PRcHAQDdLnZah/1tigR6BdoGegcqNxRoK4
k+3nV13fXizYXp0NW+OQzEtafr5+XdWSiAS7VtQqxJI22pB5NYHIV0Jvl13nc/DGVnjEiYuW/IYP
pudC9XL20Vy/6Q5DEcS4Lpgze/6/4DlORl5el/v2QSLYEzgWbdjluOBSfIHjhryW8EiLuMqiRBoY
x2hb2PHyRQfT3irE1kgh0UR4nX7JBA+NvFObMOqqF6i7wjEV223ylGfSLXHsvG+fYnJQYlS0yZom
SYPOGUi5fqKhYz8d3onjVko41tywHbEF29WngZVwhQx3c4qma4YGWLvDy0OatMNYuTdL6sI5LZH7
dAycQyyqsTk0U6AEx7fOKtSf+2fwFq26espIlpuF/MIIpQz7XMXs7djYmP09RBGwGV0oguNnw4e+
bP41T8QAlHwqwRsW7ywRu0Ss89LLu/IeHmzwpf+Gj2GIFuZGXXExOqkIpEWkC7U50sVdShiYB/C6
SuEXl6aNXh/E9wn2g4IYcBLdnExSwh+BHZ861NBNctLbYRmCApyXYAQJlbW3c/xyZpR+CawM19Jk
d8wKTMBKWAMWkgIJxWiPM2IFu/t/BOggod11QY/uBVPVDYKyGkyGQZ/OJHnhbipw5DsU12CHK4op
fvtObwM35hSg/9CQvf4v4I2RKgcoJZIWfKgECxjcfbvHRDODxuNmRCy7ybzUVx395A8raUCxOIML
AY4FYqn6WY5/5mBmX+wHbyyPqJBKxLo6HJ7JUZ5z+F4hwgc+YULc9IgxLiseErprOZJ/4F1y1g6c
yLdZqI1trC5ScdikTxITRjLMUIGomiFHk0i+DYYAdhZXbw6TKXuLANoGPjkDxftqAJpn5jcQLOiD
WNl/DlJ5Mi4eulDhLvGPcNsAC0fliwoTXbCrD4nk2AEN27fuOfS4zXfld/M27ivz0sK7W4bpXb5C
dq4zNsKRIDelo5fSvGKbgL7gtirR1AhU7KUIHgiQhDBHHLWTcy6cHrEyO45mUvlTkO9sLmnE0MBh
4rz7SXyUE0OVDbLl5HthOt2PNJtpGGfYZR+OjHl0Ob+ynNygHsdT9N2HosfXeGIMZuAuIbS4k4dr
cGinafoG078QAPtPmRGt2T37Ej5cNtNRjL3XKUS1iKiTNSSgQRSc8LA9dWIn/YBr6JK3Z4t48/rW
KXA/YMFCyihHA4Z02pAWHtBkTWmEICuJuBJuvbknTIeJBnHjh/wWvmR9gTv0Q+ueboH/m8OsPgBM
5KhVW45Ex+F1voJMYirI2t5owYQxYXBohVf5m+VgAGp1QYxLq/ObWxnDAkBcyhbaiWzFyWNdBht4
l8mEwRC5ZQWQm6qKt622T+vj/5CmVSVOWZQh6hFiqls/lFI+bbA16UtAP1/vwdFf7fYgiRu7TmeH
w1vnB3L6oXPcyqUTuhXSBgVqdKo+zgKQ53Ufxy59W+z/5R2KsyK0wCdM1DQxNzGz0oiXhmqKNoAr
4hoEtT+4CwZ2oxndPvUfp976ec9+gAYhRhqXh+s8yPDq6vaxi+ACxKJOTCYK/defRCVs12320EeL
Voa8AxFGx9DJ8rtDf+iScD3pUraVW8E97CWlqaoCU0SRAD3020yC63ZNQR9QDn7HpLu/CuTFnD32
8W03amzYk0magEZQvsjGphKZGQi0oEj2Z8jke93lJb+VI0Vgqd4DPLlOI7tLl8gsF3tLMRtzzPRQ
TKut6fn9ecgRRfstsyUxgzt2RuwoDpjldTMh3A4HZ3DWhIKaoW5hLICrP4q3Vi08z2rqbE76K7Ch
fXj5KTtaFjQ4twW2cuEsg6PJp59SrLO7uQRo6ycvFor4pwSF3sLHI9/vFrD7BlgFTlfs32BeOkEu
KboRIcLgrY/U2TDLunHw6s+aaXBwLw9rgI+RBdN5GDizo0elDgYGgvB0rOCF0kWRaV+6gq5gGUj6
KoEFZsetafOFY8EECVKqTRIvwZyYpy8Pp/fXa8IXdUA3UO4Ra+P0c6uqy5EiQBsMvO58ACg9qT0S
yhoxc+meMTHxstlokpcVlcYGuXmOsJ9KUeZO97McdBhtVw9wK9DF3PrHOgXdZVi9AK13f1KKqENj
1jLFWsYXBP3SBHuQd1rDUesAAltmvYNtCXf7nxwe7bIgQwDDbZ5nQxAfHcAwVpTIW1r10myo9T1T
Ia/9uVev9kD7USb30K4yNl7f2jtquYjUJ+0UsvRg5XRjd6w3IwNfDbVETFNByuwmWxViKIpWSF1d
HlJOteekKN/k09ak29PSpSQ04Q7TCpbxdObvjItNZ4ySkDYgC1x1BMzCv3w/y5FN9105UJBL1J9g
rX4o7/uM+CXu+WbewT+IVHgghWTmym+qFoHRVwzmjSd83gAg7K5LWMCKpCT0uHc4tzHYZrgSA9Hf
wOSNktux0+1pNH2+Pxd++pmS9oWz9KOcfsQiOjT5OcE4l6wsyPhcxWqGm651yPxOqWo4R/J0VqLy
BtjXspGbH+yag9ejE+typpGMdpEtj9pqB3Lz4ACkti5G7AaAO/IV7MDpi6ACFms19xxojANxK+1T
wI4Jm74e9jq6+DHmBmUl+z2t+HYUEQoW7O7l7IIxnEk3K2v9lf0xZsTXq8Ld6//n7qIiuQ6TjcRk
TsEFjquCcrIk4pLlK9DMsYP5sgrVZ2vGflB4Al897oRw626Uwd6BGu5zGdFk4DPT0d9y3SmBED/H
rtJCBLh3+Pgxjbfo4zQ9v6cW59nxTUdeLztzLgujn7S+z+xy0TiRDsi37gpX67Ikd4OEni2i0Ha+
VZDQPbRhV7UAdJC5nOKVA+OH6NTbPLC27H7+0urCw9xu+G2dTvvVLLVP4qmRPPF3JsGWRfYsv4bu
9raYVZtBvFII6NmiVnYhfHRVIid1zOpzyHWTXFTpQbNShvH3JT2wRyeoKukZ6r98TWPKQmLxuye3
TTTLnipPDXaRYu04BLEzFq8AXlTuT4Is3YOfVbCPqzg+02YBcxsvwM1f4Gi4oK95HevFIYAODkuO
fchvvetst7GonuX7q0Lu6zZBUO9L3NyuKaYlZxy/CUBVPMH0unJv986OEk+jOwb+253vN8HEzcDw
+vGlO15b7GIw0UDOBKJDQHbG676ZGlaCcgV4072Yy+bEuz1zdBzgbghJbPI6zyRuwHWcqDEJSkXf
tlF6c7qvapO/Uk5rM0pR+eW8ItVuBE1GQPz/9x8qcnCWcKWigbeN9q2GvrkUgZ6KZwm9zh6SwUsU
6gegTcbKbvAKea0IBe31tiZxR/5sfI9JtOW184SQaLnWOJG31cKhD0wSpdSSCIidbioLDDutT/wV
Jj2tl9+qpR8Li0JScCEMJJOqFcN6KkyltLwqD/ppYDnqTaJ67lfq+SM8ZUeZAIJGeViZ7qhBsSkj
M7hl0AEGaLRy9OHTb8qvph+gZpsGoG3hn/2lLJCSYmsLB8MLKqkTpaugnvgjm3qSyRiC12YwM3Tl
ljr88OQ9eZxVVfrbpYSntvP5Yz8mVW+6Al9tc6QyVGPy7CVKEpkk8GAvWfZkPwMdKGHwJauh6Hgd
SElraR4PUYZ+jXaMpHiRGuOHcRvgXID1TrY56DImwClO5gvuRL65qmzjZ+Zz7fK6b+zbuCuhd2RN
mQ6aCoRb/7YdzECiRoDxD5UTyRMHJcLe7Yfc4ffhMe0p0WWtnSohFnOySAx5bkpTNE+mFjNoafyM
qz0VTMY8PKxBDRDYYDYcf/8pmdyYqCDQ3aKJAHrGUHlJ0cNTyUjAiCxm0/+H9m/WodutZeQLAuPG
xuqs8oEN7Ua9vhvRJSDpECxIw0asG8hOh4KDpZ58INLLy3/FnfvzMhuUZgDTlyDHeARyKp54srYR
i+W4p7W+jJLoopL09sP6cW+V3TXr/iO0a/w2VC2PM7mq9MlK5OcjjmaPClY4JjfAYRHwIsZrqY9t
6g81VTWbiIzcQZDCL9j3joAaATdSyNzscCt2gr+cfMctg+4yT5Y/gYsbSImFWOZp5lprySqXBg3A
CvGj4nb4CHHLjnqCN1zPljudV2ojGiwbFSfUJxGrAR7JXMkubkZqr2cjOq1desK83xfXRoCwmNrf
p7X4ih1Oz8GoNN0vvBzyetE1dEq++cCA2LB4G3HVcnQ4gaimcehsoiVMKXjA5CgH44EzH8Fn/kOW
8NIUKfVuc6hYLtUjq5CO0Bn4Mf0lCeVZmvl4Y/bXOf+3OJDQ8Mez4qp7maPA4ifsccaylbAc2x30
B6x/m9/ZPADV+YH2HkvAstytC3ZQtJlXvVJjJN8O+p9fsfq1yrvp2AN/3gkOiAe3ElYAYgbX0pZZ
x0D0S+8o807CxlU+CujrFkTPmmdUGdakXzlr0PqRS4ppbNd9xPwvMw/8qvMoijjU5LsVAh0YMa3S
23jLgJzbxB0nMWjidKd21iMqjwfOoxoR8EqF40AjJRMZkAEf6S36DKVXM6R9gyx0ZmU/EgHFVEKe
3ca1XP0UmjPNOYho+75p/YpqCWfrRV06tXVOsmXAHD5BI/Ok87ox/unPfwPANABo8fKd1UqZX4PD
k9GTj36GjuFNoGvjAXNfnbPfZGTuIU/ZvUOYFK9pnfMnV7CsWpcq+LWUjjUVph+V7iwXw+Hps0a9
OH25wlwS8kM4Qn8UUyU3UMaTvzde8iDAi5yLy5WaoOVIEEFaaRgZGoiVILkWUeTjZD/5jftjta41
MBFMHZuPCMwo3CcImG24/RJSAfsNarvXY3oTcSiPwHb4ZjFOUWFCRm7/xdx/bTfwUmgML00xPfdz
nLsqM+SzI25TbfsvNysNKeoWb8A5AEZLD4u9Qq2mhpl+5j9omj9dW0cHlOygrL4Bb4+hhIzd+x5R
QC3qkZKJA4ZA7JSazH28chjlIRpEfdUZ82FVWFFJBOBjvCALMg/W8+m8nLsXadwFjLbSOYgwwKmj
iygGaQ+79GNXOmYXOa/ybEO0e2zehUqR/Z/LywVaFL0jDJlzg3Ikt3ATzQXtaDfAZxU2WcF3ucYg
OYSpcSCyP9vuZyz7O2B+nlLuxUpgvNnFOlLWJGu3b2PvaT/EMYUNaMCpjtSawke81oU/qPxVn6p3
odIarpBzYdoqE9Gu1iY1mwu3XwxfLZkqnJN4rtH6cC7IDIv6AGvc7ejYGr3Nj5oIbCTBIQwP0cJu
na59b4QlWgvRDNRor6X/rP5FhxuqHLBlD6Rj56GM4NJ5XtC2HPNhHtZ/ltF0LwH3GSmetdSJ3n+E
L3tEVYqgJ3wRK0XEZX0QGk7/ondgou9XIamrSHGvXH5bo5WxsMNF4SFvjf77WjqKV1GqPIxLiIcr
PriPG0AlJ0+WccHj7LWS3qlJmugV5+D56uMjB+UxdHcnFefTX09ox0QLjEWmL6NNkuw9lB03uosR
T3+xshAGnhN4lZIRGX4uTc+x5oDmpKAujyuexlVzcPja2w7WhdfBHtPzxxeuv+MM+CrQX4ehO44P
KNTcbxF9MfFI+lNoyG7WrQWwSHGdVjPV81ui8pDyJlIW0nJOPR3Wc2AMNBLsKGmIOilEyUexlO2U
sifOnMdfCo7842y0ZqUGub6wXnKcIhuWvd/fSbCoj4ngTOu2a82E1dLUI7PlXXxH61SHFRwmoyb8
woAtn3F61Y22LuDvJExoOOmi7oG2V3kHpkXvZJEA7PkqEAkT6brMevPd0GIpWq+AFEpGYL5OgfMH
IlATBHpF/9bKx9FW8NNojC9sO6mlKtyKy/nTJ+e9y0+cqPniWU7JB4MypHqzGimAqrLz3etValOe
KLU3uIFBamWeuZb2WQGh8jV7enfd/Wpbh5XFxyER6/fcS0zkvIn9NmY10D+ETbTPUevyKJsUh8Fz
pulLKnc5L2RYmu+1TOqHgzOPCCwZ+t7lH0ZtXvK0769YhSyXYU8RO+ouLGoBIVkaDpb1yIVuGY2w
onJqI5MmoNK/jTcHaDAc+fZMwY7Ls0o6lZ1h8Uw4L0o+obz71TM0Q9dcFftMj8PzO4buZNlOfIfq
ZYhEntTgUTrhA7oN+7t6Xb9AiERYn60WZ0Cj34UAH1tZuQaVptCtkMnCdx4dMeV0DnglHjr6rSWu
ezYB53fhKeyj1a7EAVU3rX5v9g9GgOYmoMGfWQa4wVqt182pzN1a3LeRpTR61ntYRuKxzWKr+wHq
umBsNivpaVwJBPuBHknJHwQfE+xfjry6WilH2QY8gJx/j+JpRu2WkDh5KDaTjNsatnh3MeOtsqC9
0uOMTeVl2RCurzxPQf8IwA6EJ7e+0vfg98+jmh+m7BGUmlEHQfQQ+uuL3oBfqfFZYzFpsfQv4tuM
tN2W5i6pVivPbb69nHjqDlFwTSh286pHmtxBWaBNctwpFIL9Qyoz24/yBfg1cTD+uU07tneR3mrC
JYyhpnBJyrJW2i1X+2WvDrJAHWtEA4a31WcZnkX9DIIrDUIahaC1RFNhyw++sT+tv3riylnDamuG
JBy0dU/3YhJEeMxCrVXk1kbp1DmusNHznuK9K4u6Ejgidh85hoWxX0OIjduthuoGI+XfWcHDuhbv
e0ToD1OV6x/Y13C43CQp9X8qkf0V9XNtblTjPy3gZVvk0dIxDk/gIceOSurqOE0a9VpEmSKIEczm
e9oUBqILNUAIhpn9ElbAn+klQT4mG+uk9rVCIPay2AHE+gc195ORZfX219NjSTKYgloymln7Rouu
5XncYOsFi/LIwGj6mTojSeIklfJLHXqufXdSWLoSUGW9b5i4qrdaU05djwmOD9bpoQ/m42Nql3qZ
p+gLjUXUMZ7QcTwbnb29FBxr4PXrWRheHNBasX2CjLd23TpJ0lrq/Zfk9vWb5mEZWqM/Z2rza/Bz
tf+EFdV/XB3/ZXU2OZGw6iHLmMP0pgKJsAgc16kloAzZQ2kPOzEFH6wHfqehB7wDRE2jrAc7z41W
i/7C4wNwagizATu7wLUkw9uY/hWGKSlu+qhBhy16+PIzA7WnZ0mczd2xpupNqBklG7KXn7GMY+be
Hhg1Fj4tvMyUQJ1owZ82LhcaRftxZzk+vHxxKcRtwnK63bSJObPj3PAr88oBqmV7IIAvwLGhdLU2
RJ27beB6Tn3IkdSbHray+VGB74+Ur++TRJNk0108Ek3lmsSpU8y4qhxm2MSiOSIL17m8DWQ81107
0tT515IXfNhYagEh+f1NKSKlU/i0mL5GWXeKc5y1F8D9B2dEG2MIH0qNUMjvNiudKDzyWQsAJCE2
LXEj49K7LeIVWlN7ua71ojjsrrJAlWbofNUwRh1LWuvQLV3TbDSmVr35icFT3oEoRYm4RDEWjMDu
3dEXhSSKbl/FBrr9aAlvGmAupZ9gj37FFbKp4l9g0bAiX29TbtpunYvmf4ZHIST5LMMIcBVCFrTM
H/jciWZQF9IPogeRsG/kIFhW13i67M2friuNRNMHccdVmNi9l0md28urovkJv91AnvypOn5ViKPe
7mqUQUIWh9X3RLt0KioBEyGsRX6CNP3VYKxIh4RTmmKt2nlrR8GTHSow5jaKj4zv+az8eptIVRIR
4w2QFQhB206gP1x4VlqllEwhU33n0MR0xHi7bM11MVVRgZ+HEVJynX5l7VeIRt/4OWqVWfZ23szr
SQ9sc4YxTRFov6F9sdlTJT9a048uQP7HArIYH2y2EDMD1LRmZ7LOmrizazqV4DRHMDVcrD4jNI1k
6r8XFs6iBpy02dFkvT4SjFwq72yfP1yKepwCdkXBQZ7fPbLKGDVJ0I5qJ7FiXd+nyFlhWw0SU1ZT
W3AoZuiOF/DWnGm9UVu/1ceE77IVDtD9gEbH5amQahR0Y3ecJ5fIfEIDbQ2oad5CtQl2w2sQT/i7
csK5ZFc74pUrV7gKD5USqNsxttAIFtWH1/qxy6oJaRKeXRApa/VB0sLvXEbYq/7Z3NenNsnjaa9Y
nllkizbtAIoozA8j4rcvV/14+kqNRI2N0UO/A7zZ4fToyVLZqyy5tEPDGpdNUConfnnBHE9z+aoU
pvl8IY43u57GqZ7MObKsbdWJLtlPikYyZaqge8CehHsY0Xj+cMln8fLW+etuPgzGvMzgpmynoDCQ
01Nws3fFppWqyVkgo/27wALx0JNYkknp+zEzWLqHEio700UTeHmdYZS+blypjO+MnNJhPix6peJv
ZBC5s2Uc1AgHNi1DZWXHxv5X7ofobrsB8rbUWJZcgRTg5E6SMoCsDoSmXYZdtmSuI7U+BJ/RNz1f
WMQlItxRjfaWtShY6CZDd+ZUgg2bhkwEMxm6vMgP9PshNTsigrUyhTx6iUFNczVhL7XO5eWS2WLF
2Z3mhwwo0OsX24MoHcNohnz1CJAoM2TsPeda56dr0BvHO+8+YgY8odAA9y7BxfY3PXiZPuXG2ye9
OYBV78ZfU7WVq1I/H0sOiL8XHWsEG2iIrC21hSGpa9k4/LAWTOc8RJxl0cxo0vEhNJoHlwYA5iKI
lVug6eEeSv6bsK2GE+qMbcRRx3D4hh4UuKBgmcwaDDql0FcgllcyjCLlhoMI/LqPqmjgcdvy+H09
StZmjjdjKWTcdTMDMYYOGXrSZRg0ErntAjvj6TYqahsBvsv8wuYB3XgDzUE/T17M79NLMrK5IaVu
DBj4nl1t0DDEg2TMqoSe6ijkGXSvfvsN82DVLzSy5Cz0dJwePfihMvbPWQpMWHmQS6D/s4mC1Ykr
nOVHsValRlC72xHY6yfo7Sj5FZFnrAZ8AmTmUJKjK/f2o8zo1X6IEL/3+Xqb/qgJx1bcl1QAAz39
z5VRnpUw0ql0ZhFSLNsFGcF1OZ86jPzX+Txxn7+8BPvDxt6/xOpZa/K4fR6f3NG3NzW0OzT1Pkm4
KxCYzabIt7byERXVT+PjtQFo5pHOWul5qlpwUb/eHhzyfl5qKp88Wl+T4WElNgIc86a8RvaMnBaT
m/kXL2sJp/7Y3ZcEtwOTOK+p5jkVm4m26Q/mUrRwGQMTsHrPyto/sKckoPOQSNUx3z/ogId4/uG/
mbDHPALdEgiPhrFswkHFAnQ0VcP4uT/j9okhDaWfrGA6pHmuJoXDVc0e2hBhZi+ugAvPZDuZcllU
K9gqROohVMWWpgaOlCYuokpdeyato37uWFjpV2O9jIuGiHxtk40o/DRqOj/erXMt3CGOsQlMaAYC
SvjVWqoGKGrJOr6+Lh1eXaYM0zvaQ+YA61tR+WNm1D9TLcOD4lljGffRfh9DN4YBcowSQY6mAdCn
wTaBIc3/RCSAD6E4JbG3tUzKfTrSLfNTnsrDYOSE09H214VyOlWU0lJzSGk5OSwrLwUNqy/lQ40B
PAos/gZFQA6J3Krylkgv1wEDc+g7zThRiTYUnK9lFLp55dN2mmMw9M1BC346G5SyGX2m+2xvV73g
ARXPY/inBnTM9WkCXJFGvx9zQ4kfBRzxdz3ShCg74AOxXdDQEUXiyYvt3DMYTSlNRLhIYJOIOUNH
o5Zun8MQs2iagGBvYCWzRz2amQrcuqWhi37+bikGRA+ogKb9beHhM8f09UPM3cBfyaikUK2TI33R
0bd2dbEdZAF2jJDy+aDehEUGmcUbxWenHYsQNQ1OMyxKl/1FxxIM5Qbqyc2aha62alw4KoJ8HOTn
hqTquXjqZia5nHDZnZshrW5S7GszNnG878VC7L1S7fqYihnaiGCWQbuXqMpjmzifSzyIeLuakvnh
8NZx14CEv+HnAQdqlda3VUFYlFh5FaO9RqwA7UaQJpTtqCU9QvxIOMGfYoU2EFdxRemNDtqN1Tx3
yRdpvlhNZ1Cy2C38WBfTsv7EG3yQ5upgkxfNSgmjLQl6USXwo1/wLz8cpE3UY6gdhiEsKZz9fEA4
laxR5E7agexIOEVDiRwi5J17Xv4PweHqZFZrD1rSFBGOM7yVS4TiVBQg4PrWMexgjAV/ot0LJne/
zbVl0zQb5M3+ACjrQcMxt5pZKV+VRQsDYPT097YxzYDHPmt3OiGeMXVxfdw1xuIGc+HhmKmLrC3v
KYcUC9ACnCuQoQKRZleisFxGpyARtr9mpmZI9+R6ELOrfYt2LvPDlW5zYwsH2mmUigHAi+kFWi2P
ugi0L3pPhdOJ1W8/tMwj+bgZjUvtHp/q2oLIq2/B+1LvOQniFsTSlU+nIVULQc+i2CfKXEPU1Aca
W3Hz03WHOAYMQTPviidexY63eZrZpMmIVmO0RoUkAeRtOs45+Xc9rzwgU/IgMdj1qXIrvQ9/YIld
Lv4bHHLpkQyVwgP8M8EIbAcq2zNXQ+ATNO8nlTUKXW43f9q2KdKiLMpYlHdr418wqLm+6jSdMvtw
+UoJnT58395MCJK/sMCzhaF18s4OVrAe0hy3+EG8aNy8jqr8VaBZrdW94ry4/pijBsA/aUkwAXnO
C2dpIjIurKtMnQpH+Mb7IqWVd9gmwMSORgwlJu5up24j8mX94CCfo9knnhka5WBu1faMBYzf7Bw1
qukNJ7szbC9fVMUMvqPwEBIXYg27gArSX6Oth+gN78rvruRVi0iDOy1wPC1/PWZAWqscOWxrEXLa
wHNrDeo2J7A6kQMiEeDL+5UDN796kg13E+0LxJQjDE4/1PUkU4pysx5PJeuXfE2NzzxP4ILVHUXp
LkDnvvVlxqV5GVLImcEhdp6YHUubG8IpAdlbeSrKYOFj6GjBkWx+I34ip3ppIrr9+ailOdsZpWRd
cu50RStAHC6IzOPQWIfwDS3JhGmXR14K6sgjCKNf0hed7rZyIoQvauXh6er2yKmwmE2dEzQGbgqG
zi7BAdsiPYazlhcR5/Geul9YLSU5F3cLHlYj70pSZ6lnXogU1baRKaC/f+OlBmguTYSo2WnAOci3
Iyp4a8Oh+0NmNugRZV7KIBVCUHO0j8nN2dTkdzga//eyCcUoRON/GEN3LAAocMzcs0xsOCJ32A0y
LI7VlG+JTRczrRlbB/n5//mf57AO/qwqIkbSQ+cdr+dE5hpUOYBQb5Z9Bf7VPNiBzY08TckVfL3+
QpmA1toGfawlM9XMUbCnCYUiCXg+Zq9NGg/skzsbot3FLGlCmE2SqchohGDzF5T8bOKFR3TjMQ8Q
omX045pVI2Drbn0eD2FyChz4pdFH6np3ebvW3E8NA19D/3rYiIIU7yG8qnYoWq6sk9Ux/hPf5L+N
Zd0BegkLruJC8J/cKMgmNmB++nfotB0i59yGxLJ6A2XEA2QFuFRIR4OqYlad0U0h3EQ39AosqTtv
y3pGy7AJ+ySm2TIuFBUQg8w/+PiYCMgT0IclvUM0gb1+xaShuBWIvNBY+Y/qSx9bDdrC0OXjSB0g
HDDYMj1dkLfFqSILDQUC28VRCtE1oi+6iznUEe9m2PibbF5Ke3A8LB3rCba84dCJVg5DDfSSBspE
CHt4JqpuGXEj4UIyzjQDwPhcTD8ETMWj1H4NEPwJ1rbwcJZ6onB5Gq1U7mJDYemk3gGNTV6+Rwz/
pBDrlWbMGPZMkgP+VCVlv+sAnbpMGM5xtF8XHpHTvyB5p0oPR1r8yGx08szzcNyVKNfOy+RUmSKH
oJ0ubmGmpXCslDeImxAxst4Z5gekfO51hd0wZWQceqjClQjYOGn4RvncIzYVN6BAZ6asdkitjudi
jKazqQVMln+4uXUnZUXGY8oPWAXj0bilWD8G+yYymJ/Xu1bWHkSobB7q5wEtY9oZaUel/HliIa5r
XTljJ8MUjjoK3x14s+SeF5nuBo2BOQGvqK8LME6/M+TGC8NFYFc2QbzMfizzVjUHaYJqX3LeMsON
vn+WnWHkS59HnVWgRY0PqvbJMEKL3jGoKR7OrdMEODK8aZEWohoxBHIemuUpBS17XMI6b+6oAzND
OCr8qCDJGE9apcxnbT1Xq83oLr7zTIuhsBlW7x8cmjL02odbQ3FgW6MDCsgDir2IW6ZLTFULz1UL
JdrmGlcAXBCzE/zJqTH9QLVII3/qR4kGCxl7QNoHWCTE/6CErLk8uAa4II6gIrgebhEcY060eA5g
xVDgauN7If7RVZ019iXOConbevk1tzUNbOLeco2c2/ZRPBt78INKQrih3UkY6eFkWhB+mdj+pAXq
3BkM9CMWONKNVqPgDtXzyOn5lU5zJkf7NSABda2Ri0YXEreZ6ArASq7DE3eUoe3iESTp/e1y4opU
veaKDnpjHu5wwYxW68weNjbsGYoExfrVG4YrSYAvBzzfnYwsxNGC+c7GBLsjDfpfvHDUAKp4nNT3
y0lDZRf4gg5rppghNlZZeLpRdfE//3UQPxIJCf5zf9Rg6ACYjmvKUkqnKhwMQAfDNpsSeWxpPQt/
B37q73r3N9H+QGA/+V4pA2z00sATb6OZxkBNq4vQjC2CJTaQoadbGjwdSPTludi31XpHEJpcca9D
/COQ8U6wHVGRvLwEIhxFk5MxIZ1M3wwb049S+K/CTTi+wWCYDAIhrndl+O4cv7QeNJR3PSH7GxS7
IvP+NlkQrOjO9O3RZ1XZzbaIZzxPnXd1DuUYCWdhNk3BIZDB1Nuy+sf1bnJmK5iK24h49uoUXG7E
jW0GGPYi4AkRCJaD7Q6TpjWztPKWW3wWrZNcoN8PLWn7XWv8oMRQofSNNgmYwoTMlbztT25M9jVI
+vwUI2wnpXuPTLr4pN7tPOPZ3uzOWEWYF5/CMTz0US1vlgBtWfX9rA8UXYIKZNU9piE/o2Wa4GwU
XLudW5MDOHmBPoIZIi0DJ5nxAQOL5nbhHGHzhh/XHR4AtRM/E7wFlizGfA6z8ejOZPYaSlqSk1hU
B7Hbupg3VzT0MtnDkIKzcUrCPQuQPRvmlPVA2uqXCW68wAuojwshOyxDKBOjGv3+90lKoD27S8Y+
tHGu1JlepiLFwUY5f8Dq3YEGJuHJavucPA68P/cMK1HURM0JdTH+P67vp4n24u9OPemZIXl5hZf7
wYhWv8ArlIzhx6NbUEc/XUOushINpG6y00Nr6bykdIpU4o2g8tTh31RoLSvu0NaBp0dEm/1Ba9N5
39XyptX2YmHbSa3AxFFtbQNgE30jG9JRGOUUz4Q6QamTJO77YvEKp5c3XsN2t3RWbHvieWeKUEEg
aJoNN7oTmQ3v89rmhNd+QBM1l7HyhR+7cfV2lNUsEUSBOLxiT+v/TOzSE9y5HIfoC02lEYo1SNhC
Fi+Fc32e2WwcJpsDGQcSg7fcFFMd7AJLNUbl1VMfgf4eJTvXWV6Ker7x7Uap4ApacCWyjEQ4We1Z
tsnyody6DTgIXvTf53XrVd0UAbO8oZX1c7X1T/GO4V57nBhO19/6iF4xG7fu8h/5Zu+snbh8COjv
qJ/LFanMCkMK8UA0adPCwEf55G4djt4woVfV2bw7sn9i0YnCyRvvjq8/k+3OYX6T5ljAMtjekD2p
fRWa+7DunqGG2RiAayexD5a/SFfkcDZcXse6j+28gdYypLOHZrO3YFMh/pc/4ctn4aigzjKkzhAT
MILojd63lSpgk2ksDGtcsS8WYDhScRqa+bjXzZsNEm2EnjiMlvU4j3BfR93hkfBLd5FIPfLV9aeu
2Z04zS94phAOsXKbdUdI75R82Les4tCH+vUbXOSBOF/Hs0jhLIiBn3qzP/awUTvixU1VKGEjhIvF
EkftEG6Ooy8u2376Dy1iMv0WbG41oy+4OVNyRa3suZTtKRkhxh7x4LkxEAJkS4ogQn0WU05Q6tOp
eJJnDtZs4Cmx70BW2E6dqSDYlTlzc0rCVmzZOdnQM4qxNCPFFNnOlVsHdmFyR2o4aUF0yH1HG7fb
Y6uSw7ezhUfLpNLJ1To8iG3S39sYztLvoSokyODWmXLcLlRDRGnlY76HrbAwkHFdVuq1xJ5fZwpp
6SOsPsCfyT0jyXfkyHV7F93aL0sHl259mBNoWmIf/z2nGePXDvV7GhBZNd3qp5Y9N66wpwIhATIg
PVE/Dfr/AoYNNm5zO0Ao/Ol74IOxC1JKUmdpwPsdEofflhBc6evRz4DGXPPOL2AjUXoK5lm8K+sl
WYE2xk+hZ0UK+drLTXbSTMw+w8IQ0W9e0/cRUkckyvDEOeuei5YdlLYszjcWry2UfdKkEhjQVS4s
77lj5Qygy/FQnkwk9j7GiYksfyP82yThDwTWEg1M3xJ+MrXil62ukmYDZ7hJO8H24AX4CQ7Kb61e
4G3MNVjr+d8LcrMSZdhQpoModjgFTyye8BPeJqcEG9gYiqMdTOROryjR1osmCFocqZPVD3ZG9sXv
UxUPLkGFDbUgjJ/orJAU078HmzAjxv3ZX4U9jCn1RhfU9btF53D2AhAAceA9NLsXGHvrHLpP7wwE
/5TUCa+vDgw/3cvK1RdFXNPLzcVwfZDr6hJSEwbKUoGiJ6uV6IpomsK/VQNg0zJPpW5fXVwN3596
wvxpfFbtwYgz9fq/c416Ap9+LbYMQdveI9LvPMyARdgZI14PC77ulcsfc57RS4dbm44E+Wu6azvS
pnsLI+FuFaRqLIaxiN9rTCw6zxr63wot1dQGBA+e9Y3jN+FEhU9d3PswjhgshfqzSmcPEDJZ1nf7
RHifBWhjz1X8QAA0J3g7nJfWcbdavdY8TBNf6jNsXJ0Gf0hnMGzkYOvn4B/8hg5tMKIJ4ukvgkwi
VsybDreAuiQH4gm5oJQ3Xgaob32D009LDQpPhKZL3k+ECYkbA+ySjYOWLczs8kM8GNAEg+WdIiyS
AJC0SCdjhzKiV7Sn+jvh6k6LuXoxJAzH/v5+/rJaL3Uwbrr3EgERSrrXnGLTQ0W0XpbRMI9cSYdu
vSagxEljqluArTj2GOmveQifJ2seaKal1cd8rDihHb9Z2yf3u4Uo5n+EoBpEuisfeDxkd5z/4ucH
DAt0L/zvtqLN+FirNb9dUp5aMkXYVEIYs1pwdiuO3QULpWRJT52MMjWd/dgDt8urKO495DkeQSKS
v6wFNb37pkZR0fqpd/z0gypWVdauwGUHGkIiJxT0nsPswqK7HIVwhw4d4oivHV/gJWQYNG9kTMKB
QRYuVRNf0bv177hiFHnUc8iwvLH8dRABbVFRcTO6wgOHp7X765GEVFGtIntATM4HoMz4CM1s7eBN
qt86fUX/f01u5Eh1tTXlmmRjqfljOw/7O0zIguG/BcwwkN6mjwiSrCJF1jxsNyKF7ks2hcNUPM2O
ycEwt5CprgfUza3+k3746hqTEkcttdPc4JvYOmBS5SwmRx58mYTsZsF1nogImll+Usa8EwxYUmVC
KTSuDT5QFJK3WiNi6ZUr8cKSg6hXBbbSgCZ/98EivbrDRbzFmasDa8oweE6EfZrbcZshv41azgHF
/E+GlYBo/X/zMdytNE8WxGBd/u+Sm+JAfnaodNiBpRNge0x01rlxSc3296Ple88hyNrKq4DTmM38
6jUDw/o1+l3+lJgyOuqK3bFEZdk/Z4LdzST9v77pn1kBH2PthcuTK7jYYOumklY8DGRZG65TVcKP
Kk9is857FSffiiFh6X6GTyB+7sVKdpBj2wKMaf9hAO/HmtUxSfuB74w5g5eP0sRXZ/hSU7uEnaL5
WLE/o/Dsdx0wDL7bol/dlLVaz67JPqDBXRByT2osJQDth24T69gypGDuF/SUjs01jUEgIIXEi/xX
X0bZXKf3PM7JMDXRzpYbyRZgMvqehpvIIC4L9cxTAfrirP1rfO2yC1pg9ZqovGm8rxyFJmVGH2Il
/GMC+CaW+m8jvzix+ohQkwp6Tp84IOUWzx+Yu7X7Sr+8HOzywPxd5mAxeoNqeTMROxuRTg/MsJyy
DdGaTh91jOn8mogysmyKCHxtUYm2Ud3SIxj6eLx+ZbWBMMg5FNOs2WP6++8r2O71WRY5m49sqQ74
BG7dSsdvB+E5y9+k+MsArB+sh40WndDyKBpb8dTVz8s6nCfgck7ryaE0Vp4AEwh9M3VRLk9N/aMR
F0WRbUfGpnpS+D8j6qz2E42ysgqofxc/iTbaE//DTcSstOmHAU1dQ5ugNT7iCTcrg3LEdspKisCA
lvr4EyLfwB7C8YhDLcOKKvhGcb5C8li3RhSI4yJXNYZTl5ufc0POajO/Hb6n6X1V3sdg2S5cBJL4
4U9w2UFKyMRqlZkCoctfG0SxZIHQRCiDJTDzJYrU5R14luxxwwRVwsnPiXADayjW8v+CYXVa5M9i
BmtmDJXVKgE6qQFqM+D1WgrhN3wWa4i8W09yzAZLRD2jkZUbJ+E6LAUXcIi/zADUg95xaCY1h8Av
qcdb1KxZSNaP61+Js76wWOrEdJC1CYLyDh59mQGNgk4o0zv9SBqpP3oXGmt/2lDYlY0XMmQsEvcA
pn8kscCS6+unWJlatIxnnr17E4qeJrycamt0i13u26Sm2um0ICpne7RYRSIHnPjIH6iktl/YIMyV
4MieFFd+XyUTb3AGA28El4irLy0ncjplnlKtbOTyMykfpyKzchQkaqvWsRU4wN1TmX5g8Y9ZeZzr
9P3LL9/ysyIK1uYDiUAIMtrYBs6c4klDg+xnFOwhgjWbiKco3OB+S1CJnTNlU01FxqEBRqCYJ1c1
qdAWqL14SZzpQE3IOATO++ivhix61WZ5rDZbnuIwdGzivhDADZDubUDb6d7hH+5QhosQmZlBQcRl
+/RszlU20DQnFP3hzPFgF1DdkOM+++JoeqbaBUZVtqpOHI+KWY5OdpJY4jbiKiIsnWjWjNIjImbZ
jYhN3ClpH7tvHzLxghIrMPtwr31zVu0WyK/1LsNTdzmrsVdhfGxkHvfKZHWx1OQDXYGV8YR7b96T
7QnJRpF4c6s1d3rxJsaWcn2g5aWrCyLItQrPNeFOP5e2/DdLNAnWubvcRFcS/ufbUHK9DBNi8uGH
tdVCWDS8Pl5Mi/0MwrVaG3B8joOlyVlU4riDpcj8uz6g8qMQdQNafnlE9SWnMXTG903oWAE8zJcE
Z1RHjiFHIMrNOjMzySJnZhFmMUPYbq6jtCLzn0c9wKk2n1ySMAOJto1LzuGmBU8hcKXKihVE77OO
PIae6NGkqPLf9+d49BRrCaHLIJMFTB1W9rwX4ANJ6nta1QuVWVnFpcWrdqnWMdYFOCJfAr69Yku2
ep5lZjKJft8IymOzzL04jQw+SmTl4/V768V7tCsNjHAhilnIcGpbBLkh9LWUvp8TU2XTkqWDcMXl
9B4TsE4+muYj8INTB+lMpuRB+8kPP4F8YnaHGPxM3I0icKGL7zOShxwllhNhSM1xhBlLRxK3Dn6w
vkxcQ2ZQ1o2LwuWZ32R9yj7WlMYEK9duANLBUcrluZ721TwjqUhlfISYOZAZplKBfRIOfXBEPFVq
Ndxaw31ypz3D2KZUDxbk4BkvE9QsmNSwp1bRDI+q96GehoS/sseqTkpk8DRwKCA9dbtBTEjMkZA+
DH3wKdurPVoaddY8hmKuuP38p+/q6qsagGBT0yjDA/zj7qBvOXJdk/Cptyr+9qN+81gOZohW4d9C
/P1YscuSCEgMHoPhz9bU+oUBBvrvdqCe15lgvzbbdvXx5dGXILcEKz+Zk9Gdf72/8jGN22KrxPRc
hwkyp5bG6TxIurq6KeGase9S8jk4KCIWmm9ts17LIx/8dSqQ/332P55P1a1rp8SmUIswZfBlh5H6
B3K81GBvz45CwUFff3xNESqtJbwBZ6B3KfLXUwYTmFRib2Z8hkOiHplAk3EMFB6IdONxJ/mA0OvU
RlG07iGxVZ5AFggOR/RuEAVAYNypYEfngFWe/KgUuXEjPtlvOdZ83u3f1RIQziJMlhkV7gPSY9b7
7lymFG/ERgHx9uqYi5MeLQWNRC08IeN2UTZjAk9MCWYIhrLUQAweELoIkOT4/80Zf1e+6q/Mpdvr
mNMY21WCS4IidEB2C9f6mPEkzEOCyqa9i2dj4HWLIYLgUUiw6oK/KCP9DbKEgY3O5U0zUxRVSaCu
Sz0MQsultoiBVtxw5qJ5pn6hQNj0JG1VCoK1h3p6QhY+I080BTpnIKAiL0N7EaN2Z/gGxYdlyRcc
SlK+jmIh2fEHe9i8FoLVrpGLdiONyyLvMStA+53OHpbIrSnYsAlPCEg3ytdyt44Aj6NpqphRceqe
DI7VGxP0vEPB21RhQHb+jvQilN+kwAcZPN2sxS1n0LdgWx16sboXVbubtOd0Iaz8XHPPi4kFbaIZ
EiKjvxmQ8QnYr7pe9kuPQrZH+ZN/0FmYAKMwy9EPyicWkkWnA+m7MYno5wgx8aca+Y1ni4K8X75S
4j73IyhKDJJqYExUP0aQnWCU16PRu/Q4ExHzyzoI+dCajjP5hk8hcJsIHWIJyDHvJrUtvRDBWJ/F
33YNrpQxAheJYg5057D4Lx5iQLWYjhXiJuH3rPuaY9y2lZM3EE+aluFLaKdmryHgzcfuiyUZBnU5
KmQl8g9EljACYaPVORPSR7M84W3Uemy1qAa8qECz4BtXuLubozKsVoLI79YNdMZaJMqgxVg37XIi
8+7N0DKnCqYOJ7fvk5y1Tl2U8lXlh1D8ngv2Vl3AhgJiNvDLwlLf23x1PoishP3PXZa5yZr2+kLI
XWsJs1aoTQpwbnNaZkUJnOT+YeTsm4q06kKNvlGeBoHAwQahuCCgZUBt34u8s1Er0CyhXFn6UgwT
QKDM6NrCDZ9PbEZwMB3hp0S7YkK4sYBM1CJupOe74+gENIN605eOtHGjuYEpuY1Qs5yKTsos6pl7
ZHZ/0m6AvI/MBkeCzt8d7W5RezYEYqmm5XUfIwsHZ6ao451wAKwxr3gLln5Ke5x5MGHg6Td8ZQLU
MlfqOeKQQJp5kMPbej9RsKtZPTVuJTclTvUpGfTaXGpTg3YsCgvUVZ8cZfnZUviC8ojCK4bCHy9G
i5sdnuHHbuIQs1//6B2D7tCu1s74cuWynomYubrZHBQ8zMoDPkTsEEWbKnaSpRXl1VThZp3jc1I4
bRdxNSPWtIMPYIXnvt/H+ZxIRVam/eWi09KZrnk9GndILWquGaMJe3ejiqfF61crDAdKlhubbYN1
GAmzv6RfVJIaSgxu0FCYMgDAm4ackpdZkKFJqA+5d5NbtSIF5qrX7TQiSDXuOmVVcJNMlVM8HX9Z
roWA1kJmHCkpM/tJrrZB5zdGi5k9JLJ2rgji0SJPacLLW99aTPPExUqajR/7LxvxVN3uEHuZ3dOx
/yLzYS0CSB3dFqpau2ZDNRs44n2svKvYPhYgObwIMwpA63JtGoQetA2WRFoiL5/khn075WWvpLKv
TMksGriRwHW+6xL8AjKf4P0wy8OCQqqv8pZX/KIcblWS3DAlih7z/RN74oI7YwNUCrgen07MB7+v
My8yReWfJ4BSHYXvl/s42hi4qJnWVqiZRCld18cq011x6fXc8pvyavh/05emkciGSGyF/l24urKh
F2v0j4mqaWkeM+HGbMyXbq4Gu652iq6Ub9mk+sxTY5NXxv/CCi9StpQmXZORyqEvouAmnRGiEHyL
awMfqlGJzf1L64fF41R6BUHWOjMoUzhsVxqBpQx7PBZ9yeTvcZLJ3dzsh5DxnA2AnoOjT39RdHD0
lGJy4KAyPprI5ynLpqOAAl3+LTiuiyy62+33I0PuZmqzgRPRE/s/mRvJWdZqL32ESLp8S3c6y0vD
hoNXJhnNsurtpX2TsZhrA1ot8HPGjZvlVw5U7CIxUCp3zVdLgVikxjvEe8ewQrFoAqEiuXPQfkAa
n84AdD1H764ydR2OsGwM+wi+4a+9DkmOulazK+RtJrvvK7VpU1ExDQhTp1vQv163RZX3Kgz49HkA
EGKWVkFcZBKployXsSgPqWwyneO+As5UB5+v6JmmokzRR0OF7Gqcgkleg6TTsEFNkqw7m4/1S4ys
Nlz2fSbFOtKTCLjEPDOuFk42xcOjbE342NNBBcneco3dQ+r8L+QYt2lUbH8W+VypKHE5rL1T6395
vrb9QhoYGYhfInl5+y2MCULEga7E/k25aNsWcFJegllWTU3J7XO78XpOEXJSJVRzUQ7yWj7Pa3sQ
fuoq2w9Sn/cqkvos3p71Ds+OlnEvkCjg4AVshiPSovqFFg+aq6fsYKxLE1vS3aLdSs0akjhofHEX
qnTDEx3mg796mn2ees5dKcsmKCv1VTgQ66W0wfpFf92hzo+Ks9Vq7Ea9ZCiH/0F+UiReipXgNt8s
jriUU7nWS+0BAJ6q8eLcod88rZLrCrZkIcco5OfgFAbZxdjds7fwJoeH89tBlX8pL6XWbGPcGFNW
AWceJEBppKyhfme0KcmcD1NLhkDWM7ErHoYDhH6CtzR3xKmJIQL/Lwm/o6UR2BIhrsGsAShh/itR
DwKaDyvx1H6CAK72dwtAipnTcDGJeIeGpT/hMRt+5lsyPYpbeqPfxzsXp6r95e2cDAcohh1sPxtf
Af9taDcagh0TNR77cT+a6xpT24rTBmYfZ3us72NuH38kCwc0D47pPqAyjD5iE2m+zUDB4ppEbtVa
vwglydhTwnw4egl5gPdFEJxrqTrzP770xakVFPz4AEUQzOOVXl26ahtB4Y3khqS+ZgXNLNqMCQhl
Z3r5tJx0+jsjanP+YQp88L6v8O7+9qkwGcEhRU2eot/XMXqvnHSA9NGfQ3wgm4cypo5XIuAVXqbj
WeADUcCFCgVC9ccbXe1nGmb1M/v//Z0jewkglTn9UYFBWEWAGQiTB/RbUg067U8gfa6ghJGwFlgB
vdaZ7XTm/6KL4U9+NJKHPqbU3LukJeLUJo+oggRlGH8WSr4FQnenTKgJSCjRA+M/RUuL4JPfQbfP
5ta+sancvTkqH23nPUyPvdUSn8hJ1eU9kAKiAEaAH7QbhZRNNqA/ONoe2DhZRjdgEeHbyJrCQ6p/
pZVm/ie/jZ/WkfQFib9kPG1iIAI4tJEStpzoiNYGofRELX1Dw7/+9/0rOEQvCA4Q2AnlV6wkzAFc
JqfeSMPshH2t/be72K5EX6ie4WU25EBdQHkquyWHtHv9rhXAlqhYXYZ3/11g0OH86IjdwajRRXZZ
l6DXosd2XgNMpRNhkTYppAToipiD0LsesRyCEoZOYGu/sp3tqSlpRCvYPN2sx34N8esnmR//AOmg
+ryxERmb8tU91s3KFFx5jAyHHCeUOAw9oLnoxFNgOkNp/ViVCTy18TBno34sU6tg4+OVu6eR/SfT
kEHWVk3Qaap2Eb7kgTC5stln+MsobRexJw4i3HFGoubkCDueJ3rsDLtFjyB2b0ce9+JfpHhaNBEQ
AHcr5/RrFKnrDGE4bZYy2xLXEmeMrytT1GUn+16SySjFPvmr26l44kk5KCn2CWraLWn1dL46e/jJ
FfDaeyH4hYEdmi94zIiU1W1drQdyn1YBs4lNRAkR5kaJRa1hB1JoilQDvG+fKr4avI8P9zDU7e8/
O9LXW9fyGFIy3gbo/C57cR4bq1lkjCSjEOF4Ef1v4ZEH7OpEWIV+zVufpGASGMpNqjvY9QQs17x8
vM8XQ1fwrXG8rPgX88xVT9iD6/wCl92D25eTDfUGKLHme0AaU0CEbr7FVwZEh25cfti3jRJ4OB/A
og6CuBDqhSmaohbsYMpIQEIVy/vkfNu35CAZS9I3IrlGo3lznt9iLat4kMaEz/tS1IUkSOcyovDN
lP3SNuZA8EYyA0OPPKNcw3UIqvA1qtV7oMr5NEQKA6vbxJghgkVt8/FRGkJ1JglHm3Zl2M7KltXQ
FgSiULBh9UJ1nFrbTn//I2xfUy3o1wZjJRxZn2ciA89ETiy9NTkhe3rzX7YuB8mUWQQ9nPlamR5G
EGZTmydq+JY7HKyDVxOqICAilpNOm7Iyv5/OFs/i+XJB25x+WGljuZmbopfuhxLY3EpTg3rqrL4S
2SCscFoQRqfdtVzfACEu+M8jZBHcfN0rExSeaqh1efjrFqpJfMHmpnHdlChuHKv87I9Cd19vCnik
3lBLqyhmgGi1KeCBsTfNZMUsASLqbah7Njxz0KcVAQHe4MDCfphnbYBbDa9HaoM4qu+gqccGDzBr
KedUIlDMXkxHXvdsV4U0vHY3zlRPQF9Le9AqBPoyyyj+be9R2mpp2I9v44MVyKYzMZW1GrdukpZi
wR+wTTWs6ja0XPblGN8UlasfpSBbSxDY0lKcA+smyGvAdzg53QedSNcyKNDwPpM9qJ5tSF1IKr/W
zOn/xYq0zO1dQ2e2yv/s+Y+V5wj7IiQHQEKt+/Yr2tG0XR9+priVvFkIGt2ZQWC+eh81yRxJ12J0
7nj9XJmvtqFgmWd8to8+XcheIUW48B+0bMg96N1b+LhE34Yu8IyV6wkUgywSGxPy98eUzzNgWDh+
O79VWjZ1yQOmygNgkJTyQSunGAgFuzZV+ArjWpUfnlMatRmhW4xnc/rbQhyRQUBxby6At1umDTpB
N0ZH1ROE2YK/mU9/GjlJ3Dzfnxipic3HkxgZlU/FVesdZnlUhsSQ4Vj8rUnTZsJRTWV0OyqzOnsg
X/TPR8saHKDw4dZXfRWIUqIXWMBO1vEDgcvTSwCVG5kJex9qES/TMJ7dA31u2eo8SY47eWbtiJ4Z
P91qDVL2HoG2Y3q4SM0H0hlVUWxa1u0EabTNc2H2Wti7YXeHw1x+0v16LyFMAz8BEgN8fgQMw6ga
cHhMoob/7t84E2tFvBooqcGhcdY/IHzVjk3F+ANw2tzg3jOUg/QyNGcFfwzO7ccstLMzUBW1XcNd
rcV1uHYXyPoL23bs80kVpwOXcIl2xzIYZVOwL96kpvgqqKvklJQjhHeAuOtb27yke1q/hsSWWi9l
mRLP3SUEOy3MMAHxzhnhOsvYem9xEjYkoOZSZAW7gj6YSBGoIt5Pdz5XmxtOdY7G0B96oB4Vo8tj
baA4RsUjU7lahHFxf87g6r/Xd0o/E9+xYtycUbikbks+sCxMb8anHHEw3fp7x4PTLkFXdXBrlzaZ
4LC+cy86J3qxfqa6I76FjW8v8lGdSpNjxk2bp6TZk3pgWMwqST6DpOliNy9kZxNYy3GmweRkpuSg
AXYvsH8B5TSAKJxezpLtFD5sLb/61KaUXJzKfj5CWHZ889Yxe2popeWQRdB8t+iGXAgb3A5KCLU4
mX0Vns2Z0hjaD9k/f3uUrlebtDcOTRIieomVZJ47swblG4nAdPVkjtRe9eBLe11bPPDWqzTDxE2i
7p+0sJu0MaQiNq7Crp5dn9v7aCo5odvzSCYT1lHU8zVrNXS0IsBNglgZvIjypAQjiS73rxqXb2/P
07htJ0fn4ZjqO/SjYB+onfdU0cBpF3O4muRyfnjzzq+SqCDWQVAIgqC42ieS4IWbsdtZwbnUBkGs
boNiP10CP1r4Ct8FBnQi0qzTfY7N0diEEQkEVGZLsNW4bKrlMf2Oqo3OkouYUuBBSJf9PuheBvNX
lfNM+dO/FWBFz6v7JXmz2NJ9MimpxDWdGknGKlbq/v/7t05VgDE06YufF7A/W8ZGIjPRPMhBaawr
MSzZHWVAK3MwkCVhPYo86uBtgJN4aTAi2U+/UD66Fhm9oE+QN7yFdrZ1fx8/N1pYU93tJvflV/6m
9tqCd3fLl1MfgCkTTUHMwdFQwbnkwPvjXl/dAZis41AC4O3dn4QJVPOsF5mpse2RtFFpCKVWwVku
KBn0geMlPwzY3w0S+eD9yGMIgQGmtTu61VzmxEolywtZpYk9ZiMhHoLKe2Xd5qTqmBv0MqNGc6iz
KxPWhkMC27CX6SL9S6t+J0Q9XRvtebwkV3ljEmv2m+tmTmnI9HtNDzMjAV+U0yymamecSffHPArp
FvF/lQ0SRA7Pp/89Aas/aLBa7g/+v1sNDX1i5gLXtMdCBnBRvOzd1SZCBUfel5qk5uQhpjRJOUHC
4+udTQMmURrHhySptjRIJQRcMTpKnw5wk4l7vjlgLT4Oe6oeuc31QhPuHHGWJhuJXepoCJf+AF3A
5rSvw5JHnX0IPAhjM8wmwbMLso4pJ6JePpNt8vXOXTjwSUnWG/gGdCKi2yhwGFdgCKh4EwEKChi5
eql74LmJ0FfCIFBfgwyxlrZBlnMJMen4rCWTNlYH83rmPtxVm8GMZhaC3vf6ukDqPx3YjJrJZgeA
lZ+dMb5VkJyj6HDT0zAO9LigOSMvk/4m2Qs67kMASFWjX4jU8o5mvwEFC0Z1oafweZcL3tsQnELq
nP3c29lt5SSHtfUMspGTqX85+v7x4E8S72R1/doty3eCE37PHX8vHT+pYXXBodnPZXCK5ISOxAhV
YJOW7nj77oW7ZaLNxu2uFSBgTYBwKbtuWV8sprfLnPIGMG1oyUrPnSfVmy/am8794TnmbtQwDIE5
evwYKOqZTE9Ce0Iyg4VJ19EVeZVmLuc/5Okg4jc57u9g0KHANkbcQ2nnLlTpZwRi622vjqQhjhNs
1ODafbTekpnBubRnLlRT/T5l6K7VmiBXh/2pKgKyxXy9OxyAUE22RxQuKIMqRdBgPQ90MM0LTAaG
Z9mUXSAhtNBb/ftHbkaTGf6ea/jpIDnoS0UkNjMWyuOlflPN6l/iNddTlWz6mLvrmNNVX4AMV1iw
a6V90mnZ72zmyKniAwoXpI2BMjZzup9S7/BlSo1VfSTUW9tpG7Lw9+ZPT9rM9vUTmmHARZyq2pAt
ZapixTEQf5a5wGjkTVbR9+AGNtCEBQia5T7Jr5RbacuDMHGVoUfalWf2LsthMWtxezXN+0pHN8pZ
j05VGmX2KyWN4mpIePzw38UwCu83CDYUNZXROiuF1/drkiCLAFOP1cGH2aHava6nDcWugKfHhrDA
n+Xvx2bIE3MtbzCCJAFxBE4WlmgYPZzP7QBvmwn4s/KYneNvBIItqhTfBZUZxhlMH2Fxf3ydlCLX
FaA26KOaHNBRPLQAL5oQm2u15TGLmhOEIJU3BQ7n/YN5M9+bH6QOI+leRsu/dTwc2HiSyhPrRVhl
1YujmXuj+ssTpFu7MJMZ4NbQJdelO3pfNFtO/OJOYKP0Mj6z2Xr9nAmWbNlTduJzhBNpqrWN+lav
kSNTAc6dbRdxzRI1KCPeg3QXPWtyUeG45rXu3JdRZwpFvwGAzzK0aTbGctxctRiPfjw+tXT1ssBZ
lxtLG485d2gzT1l8uOa5UuDqNdfdcZ9rYJYhPCzWGU52rMYqeyRkVp1LQ6aKHfcUCSTwBttGPMbN
fw86vERT1oc11wKSfLMVffYTNc7m1lK1BB62aQVLXfHWWpPH0ztJjPm17kzmN0OEwlrHWAby0fId
PgJtxYkeACV4XWE9CQDzsSXxiXl2WVHxuvhUfRUOBVWZN2mJFz/yg5hQeWdqg39uYxJJlP9vswTx
ZnXLdocKVMQtMi9f/i1lKPYrRhfz7stRWxPG6TUQkFUENhbvQq1F5lSjlolDhYMzUITpKdR/2qBi
1X3W2Din0RrQCAcgU73xBIjdvKrzq9XPNICUPva8Irmpn0CJlANZEkMT11Z2CX+4VZx3ehtR1/E6
lEAfzFDdfJLuUtdh+VqjXpLXYbSNfDG4Ni0MSJHucoskJaYVvfbTp17GLOvA1T1PT+1UHCJuxzYO
4sZQnTBYePD8IJt2Yp7e/giTJkkIr+cPEIpyC3bUlGr+I7CPmrCL2ljCqtYgowWQMshwmybixDeF
wozs2fyF3DatOwZp28XVcNzkFyS7msAOsArSbXcaH0KBCRmJWw3DMcSXDUxnlTzk6yubEqNTaIT6
Xuj+ghSE+zdAXGgPYbnhSY2jJdbhQ11HbGhzv0MHMLGSScRHVrp63YaFbydlM4XAKbpvC9qMCYgF
dSq5T418nzml/SVyI7ph7DFWmC7NRcKtwD6ZxphXlB2WLZD7UGnZnRSnKwlD5iTOJElFDNpRuU2D
qTqOFluWiZOfc9VqN01WefPlQVLFhGVeu35Gs3965f5b8veCBlvQAcjqNi0EpRAczxCqzwuB2syJ
4WkLYlmdCIPHYStmErIZdHxMq4RDGoqbi9aSopDzKK5WYeR8LAfA46lcqAroQSBwgtVURwOvsHFa
+q4LoDiYYbDV1YSZ+j9gKwRE1D19KIrC93skgR67Nq95qTxaMtGnzWugdPG8vxZjUwarpiwYM51u
owirlt1P8d4LilG6U2ZXvTYI6RMbeiCF0EcW2vlISeEZxyrabmuFBMzZinkd2MiDFI4k5thnJ0QT
2h5smE3GcROgmsNQT+Ahu5BU9FxY1aWGU+mHUnwoajoLvOiOuSFa1IiO20sHgV7f8vP+PPCJJyag
sPgIL6FSa82Y1i1ds+R39TOysdGD2hOfUPwkZ7uRRFKNzPFHCbS49kA4+7hYktUD9RzWYIhHTMoI
0brYDAvBnFjuAyukyWe48ZB472mIaHY76zbS9EJ955Jv/UTmtYgSGkFNDHWekOWFPUqDF3obmyZd
SNAnriUKoAQhrdTNgxsFZ1AbQw3AKHVBVBY5noIWsWQEAuV6amHzgOawKfCkpvzgHTeW+BZ2ns+z
JscA4RQ8TDCdnCKUU/JJbtuJVMpINOEIAk2uq3y2gxkvKeagNxhZNCyuEH/NCFUbrdf2EbKUv5Ch
LvME1mLwdu9PO+bA/4EFn53lddrOnbnrk7BXgo70SaYZ2fek0oo9uRMRCee9m3ulNPSKPYIzYv6h
lLD1TKKuoF52t0iJRDMJyHMVSbGOIFcd3bzBKCABnXRV1fcy4z4fzWwYkXWypEsBkrg65Hks2RrT
8N05RkcVLN8E9GYz1gQccy/hSTOn91cLUDYdlhgrwFlUUCtKEMQ0Uz1KEOLRdFiyePotmpswQjnL
NktSEvvSH6yz/hiE4sI4/7q15z7qjb1VvMkOlIGjbxAjYSfE7DChTA1CST/chhBW1CqGh6wuB6LR
U3ZNWZVVRAo5oHkTYo/S6JhmUTk9BKSTYoEH2iW48ORud9YM26BOLHbJZXdAuvmIZGvqrLemscwo
KDMJw1/vB1YEGeZ2EmTRzJAXSFzInFwGGiXnbogTPYaesVnnJT0jgfitqB2KdzSA1Q/2WpWr54Ws
wnclinGcJrRnewzCsy+wSSpZtHuOfyTroL0wkCboOBai+oCkvqigYSXUHEHtpIHGIJl+PcZcacS/
SCMqzGr/Fu46hoSbREt056y5v32xBu8eIkMe/jwbKbm4XbcN6rZVN1/He/k0igwt9eSL3Fd7MRf/
BRirDrpKVXArRHS1m+SXwoinOdZDeBUf2wIezLqgiByG/3MCs+o96ZeELEy+sRqLayPkO+riv0Cz
Y3R5B1wXVYNcEm7bW/PovTkDeUNIjJc9BSVikH7yMVPqJdpgQw7l/XYTkASous7V/boRIHw0UDTP
e2FV7dC3D8ixmd9ZrhK9uceflRMCXOTqUbxaCQ+Riur9Z1LfMvD3xBKzXWWb6cz9shGKczdVuCXT
rOe4A6ektr11Hww+js/Ti9EdZQ6q5XXqiOx/Jg7TZ+zDONyDv7b5oacEnrzB/HjyH+u3E1kSoby9
zYq41cH/5RdF5P+B4ts1RFV/RgfHf/IoJzTshee5pQh7AwseBeqYy4r7qNAHugKOw4ajr0vw9W4a
d9TEP9UM/lIE/G2rm75+ScwR/cbbZXQaAck4mQMHw1xDGok+VJ3Umo8uAZex35obfBwFP5xTHycx
dpUJhWnZfnaqEFQfTnRDm/ZSBmlxA7B4OEb2UR5/ZDOS5T/w1KcLFGPA77RYkgpm4HiZy92xsaX7
jr9VLfDM+eFkty7Qec7hmhmWnYtP0cCt3saAp5h07wB47ORoFfXAmi1+o+Tt6nQKKsUuYDrEVaDM
SF9BtRvfG2Y3CTrK3do/TP6CT8mqv7JAIfdqt5iPhA7Nb3iEtsaYnvpJjp5RzWZEfDlSjuQ2YCQZ
IXLV/1TV6gkzUtgVVN8XMEaBhZOYh4YVnbMb2mAPKgj5gxYWZBvFnW7AZ70JOPzoNBgqCkF/AILm
agxXSAexWKm8vZGNpenGki35QdJThHLWgVo3AMxllIl84jxrWbd1qmct4OTyjduix+Cc18q8TdKt
M6UXoqZKbF6dP1EsO4b60TbKPu5i3ADQikXO7df2YaSmw8tAUHjk7WW/zeFjDJcMurcY0VcGIiOQ
QsexU0EyTAZR762+0aglGCEFHW9pZ6ujdueYage83OgFdrcuSykN+eSCkpQN4cbtgfUVSdsHNRFL
FC+JQ/Y50W2j2Edll+XHeqo9+5xGFS4iI6SRCHYQmY2tMWlKoyHBm9YoB95vuPPkXd8RvSMefoqo
BcG49xWG9q32i0rswzahwO9eagNOTOm+bCTg4kkP13LaQ6oen1PNW/Eaff296K/KOIGtqj/YQRfy
HoRFCM2UV2T/U7Ygh8GqJ66BhDNQ5lk6hY77IP8Oj5I8yvE15mZCK4+S/aG1CWgBKfYBQMzPRD4d
PH1OErnMt2aVhJaaKsUzYq6aM1FgfXnHifo3DX2xgCL4CLNjlAPQidrJGSs6NHX3sNJlq9163SEf
g2PIAVfW6Uv8BgbrZkgYutOJjqEGN8o9sp4A2ntIbV45fZnWf7UxSTBZKBGURhLQLGAN/VtkfdJr
1xvOsgPlvxSctIrPHJxRyRehXcWVoyATF/hgocwpMExqjR9e7/cZd4b1keh1K97hlrV7US40tUx3
rCVbmEs9MWulMQmGhWfjDJp3AltkxiTQRQC4Z2arRwf4QWQ26u1XX2FCa9bLerwKybnbeaCOLHEF
j5A2VDBfZ3p6bYLil5KPOv7CNg/dWFZRx5EMYA9wxVRhewxys0MtY/ZPRrZ8pVuaZZxxNC2TkZHc
XqPkoV1ogbJ1eCatdt7kWDtwC/o7kHmXdYkqApIuGtQLxhbcF3pGJJUuK+L/0EI3xAkOEEPhki2E
YEyX9r3x3UiS9wWdnjq+3rYSmh9l8K8NaCgDE01IyewefEd34ake33vkMBM6JSlA/eBp2FfRNx3A
OM/VRq7d0UREy9eALyUj4BJ+oTAhoo6XYJBHbCT3QdIp+Qel8DAkO1Vx1TM6+ct7/QKbImgmVjYv
xK9PAOxkd/hImNHHzRb8/gcjJQ+ceonRbKC8wxigC36wsTsesfNBn389Crk2xR/DUHykb+sK4gzI
KEVFzRcrE9ZpHTdCpzTtsg9JKC2T0NLifDI01Iz/GNG9Eib0BNbE7mSwG78QhFRjn0njFSy69+Y5
y1Ibhgrcg/N/1x3+32gD/geRkEBylmjSyBBYhmIOzYD/c4R9MSXHYMPjqtbx5oRD3X9ZaRAZU+JJ
U3GfDcxQ466GE9cMCQxPO5hmFmXGhPJPfVY3+E1KC5/jw+idxwzKjwk5eQJqHbiJ71Ds2rgpdjcE
8XTCQ4psz5yWMSQY08nDLedkwiGj1IshObmKqvt0erf1uETFxS53BoBKakgwUYVfDASFSKq6hnJ9
F7+dh5ZZJ6reiacm4LF/uVhbVSO9+9xuwfRv0y6NcIjlxAM/I5Z14wckswfphIfiFDv2HnXSayXr
HhxR4610hlSrbsJNtmaBbGCgmcy8iZoChegzCMThk7qtfw384Uks/hT+51v7Ne9U/v4TGckTkONl
kNz6wnoAPZdzUkZ4GYxMB+rZEQz2Ct06AmW4P9X8UQmMvcOAj3MR9sPVPF+fri1k0wxGKJnGsQvN
69cv0k7Uaku134C4fcFAKkB56mwHo3NdHAqpzqdLuytQuJuUWltnCqVu2ttTFO9Vg0zoCZJWCFtH
Gk55438lALv1ygt1vkJAvflREAPhX9PhqgwiXdiRVoo0/fCPthqep0QMNS3PjMnv91OpCzkBxB0s
EcoGIADQgrniVeknQspnlIPG7y9gNBXfBa2xT4LmbgVbLSiArPlIFoS3SawgVOSy9o4PLPQK3x5T
+ExmLT1VcATB+ucQJ/LMsv78Zjd0kDsZLD8tXsb5IWhCL2C1Jyvm68s2nEUj13ZOaUXGnSt/cOof
rZttXsb33S3VjNOyDLcX4+GLj6w4DnHIAa7sL8ljqK8vi0WqvwyVl/y3mQyvvL9IgSl+kaeV5401
8NO4AZo+Yls9FY5fKw8FRme/40bwC1NgxdjxHPGw6je6p7TXTiE9cgXDcc2nmFCwOWAVpwjVVLgR
e5hxzJU4aPpBf4agBFpGZ264Tv87EDKDi3LJVI5oCMBuHzJCZgm408oRV58xhmaJJGiMOtqAm9ij
0jIpqFoVhAk+BD0gOsmoWPyT2+Cl9/kz8o+UjAM/eIDWjQK7YybuBu9snFXpI+OMKpEcXtYLuuxU
u8ZUA80l7j7oWt975XP9oFM8KVZTTJavao3fHASijWEZiu1dSTDOeHT+JLQcLTTttsW5dgFiGG2m
fHjf7ohnz72tr1WHzyKnlfU30LmVjn4MSb6dA5bLiCex5mSnNSq1oFhuFN0PKSNqW3gXIbkjuUjN
2Vq/7U51+XmnfPsRLaZMP9tUG/r95W6SEJq2rXsywmlUamBwX1CZe4R6QdNPKxQ10dilb4EBAeCi
KD3lVSI2OOhdFir8hwSGyNe6C49yfjd5sFGsGP1qsOFH2/rQd1sOXcq5mVXCBdgvYsrsRpFuzROT
Du/r7NemrMkhGOzOp7UoMk5VhCGTffWGHCrrad4/GjtxLetabOlyg45lR6CCoYSsILVWYV+8YTno
QJ+goVHiIHapi6cc5Zb5B+tHD3pUFH/g+F5/0ZpgWqkWZS30HJuQdb4bNG+f6Zt6i9a9Ve80dGiR
6LAF8E9zZJPvyCB6ivbBeq0ii4gTGztaUps7WZ1jkvprJOzmoMT3zCDxnUUWXFJ7ummuYjIe4kbS
ZTNwaEu9uLQ4xzoodOLTT1wq1JVf6pxJqFp/Laq5v6XjBlEvAzgpWrOcn8GGoH3dnS6O+hGEfa/l
CQ/Cg+nj28rjMCK3vl5kZV/xhfh2j7n25V6yvuXwPEkPqTlKPC27CHF/mmIi1X6kXOiGSmEotAUy
bGdJdTk6B8hejJ9K9VKb9CeRkdcITnPdlvQP03huiTJCQeyMlisSLUmgCJj7G+E23Ms6/WosyZzG
a5OOodXwR7Y4e5OOQnOIq2lnMGp//EQOFNRqWLGZgdossiWEih3gC9E8EDLjpqQTy5/Hli2mLqAl
tYIHpYwXxuq19OQ0gtTHVnFnH2De2ZfeOzAnHpVg62VpbfBtqfaA7sliVYSWSp57DcT80KPdY2CA
FWMQUmL2QrmynPw7HGjCrPszikt77uAnN6iIItz8GOsFMnEkWfSWz6Hts88RE5JLZvF3wLuhPo9p
jxXLlD0Z4dMTAk71oohFtnWz01plDb/qfXZUK6TCrImY0KuRlwAh99bte5nQJYF/t7dagzc3QXDb
xVx7v9bNeUSSYHBJsFhwqHSkhUrnKAkE0goxnAn6FPFSUM3MdH9I1DqmjJoH05VRuB/pR69SIKis
0vte0XWwhJ+pKUII8xxMgk3c/98ibigexv4RHEqrFzziQ4YW6CJrlifkEaeqZoAIlIViDgJmFkdz
dLchfa6vabYecXOKFy/Sl/SiwEeVpw5QYfqpBVuJG0Mmq0nXbjtFFvlrtM1nbD18ZnEDI4Lf+aZE
NM9UccKpqlJt0GntFI+FG1Ca4lbisSXhf1CEZAsgiVhOKu+saCqoKg0BgjAQuDaGkYr462RLKEzn
y/1s/LaHpXvmzwJqsz0i7iFeVleO5NPCEGxAV+x9ErWnWs93LMklxBme1IKRneRzSS8obvgZ1UBs
QEP2Wy+u+pnobnwm0rRJw84BYFPZUZ8ADwH2Q3YPa/TK1FV1vdU9TE+kiP+SV4zT0wgDA/xHs6cU
NQ5eGZHUJ8VeKYeCxm7rNISbTe7nZpBo2TMTvsXesa/FONNgG3DLuusbEI5Mycztu0OYSbfCOekv
HdIs5BpNnmVM7ql0oaS+PhxUoQPYpFuSI37Bx5dFb+g8v38ndfbFBo8HLVuvj00pqQp32KhjkzS+
aGlBhE4cHaddE+GqyEogCqCWphFNvyyLnn8ZsiAVTO17Ug1gtpCqqOzYSw7PJi+AprNq+mF26RMd
87psiooPrWwGtfcAMrY6rv2n8obNiQFPGsSpm9aEhhPHYVjQ0KWE2djIazuswKa2Qr4nXhI3I6YI
nCMJU7pRWXbwIk9qaGU/KIbLJf60bdZbyY3UfNbtNyv9A3AVrfZTg89WCSahODBhQqFubEZCUTkz
8GilIKYDpRE5oOzgp6wwpeKT5qXtSNdKb0tbUwKe6gUc6tu3ixVweTajkGTABMumoIBP05hC3HlC
bJw0EGEwxO1R0sg2s2D6oiKoyfn0Y7VLHxsuL3gY47asknXARQimCVOODjH1ADk8biZ97uK/2/ml
ZBguC6fzwOzn2ifBlOD3abtrXZvurYrZsVvxFbTq8YUsDkhp/035GbugT3V0DxwffJbDc+r/rFGL
CWLbPLevBMkEJN6CMbquGdjOMX0BdFPhUAFoVhi0C41PZl4d47v6anOsYTE6LwQ/4FskWz8WyXD8
tjICfI8NzqQFW5hW3vF5aDf8XZIeTZE0C+DwlouYzv/VDzhPBVVKGXAgR0lPI0caxSqMwvOgcn9T
sy6okaP3AmsAxXj2I5QwkZZlek/vnEtDTbtP2HPYs+NpO/JmPLs9fxKozx7VBsecxjqgSaxkBKuF
hdfNauQhZ7qhv/GmUawlq7AyBEE0Hyok4eKtaLoi8m6YkW+ROh8n+vmOO+FUQkhZ9GbykBh6VlAL
IZ1t5MAuspoQT7PAgWHlr4ic/ApuDhCKT7IHmPvnJZvjK9Ox6d1I3V1pP2eUjdKEMV/lOGNpuriP
7RVjNJM5VVcltyoAR2Gc9MgGjnoQVr5T5GDkCkFK5YYhrLvUjdQwgHaiGQ3uods3v3k6lKL4belN
T1iQE5gaBKWKZ2gW3ZrpfkuuFdubq/Lqt9/2q22qiXqZtCKcBJKbYsvKNqgHnNd3AKWDrTmI15va
60As1nDV6qEQ4xgZL4AXS9jqma+kmXQKGVzWcoXs0WfbwVck3gqa7sfmWatvW1jPCLrz5CmAxZt9
SmLRFIR5vufkTJS9C9RwUds+iQyrSFTRYU4ogaACJOoFHgbQdsXmMemfii9AvdSTc/0mypnKpUBV
J7diqlTRYTNdtPlZr/nrKs/qq4MzjbqAdCb6G3Ljdxyf3NCLZCZY3ry9yDjlzHYck83gfMBeMwc+
iewD6+gY1t18hGgi2v+qlSnj0bq4vQwwEnNDomlv2Qo6oVEJudiR0GfAN0ekZQ0myNJyHZP7s+/R
NKI5NPEWIEAQ9x6CSx8sMtVlo6ac/3hLngouMd/ollIBphYvTomXoTLoZyHLbQdm0a4vHiIr7vAQ
Im0KrXZR493vwZq2Rtb96HaNCKlq19sQU2dC+L2F9D0ZIKqawniottbqOVA/ljCVd970xHr9+yiZ
qjwLM04BEQZsnw2sVnzbXDCG7p+cb30zak2zm/BruVO0O0TvSy1sQwNOlxNz3oDFZupZJn8N5+vc
kgPhFL8H9/Z/qDdi61Rr794JmdzLfJt8Tf91bYd0QnnB+J5F6WC1ciu6ePxVwKD7aXbB50B9uH2r
6MpU5wiCqjv1/C5VMEbbll+71NElezIcqLfOQ2OpJb3G5U+cOPtvkJgExREW+zzblhw9aXU3ziHJ
QEXwJRcQnv2zZWGn6EZCtv0grU+5ZhVYTN420LPM3VVZr8byJZP1Hv0E9OiwKPVi6HMir1Msp9K1
iXVmTqrdTUJqH07vnWQdM+7RDeZEuGcZBYkHSPB2aq/lAioXPBrZMwFYLZ6MYwd7lVxGRkSIikLz
zdAtAMQwCaRGe8fsFW+ZI75EjI78d9rgKLSSCYraOUOYiiy9VOVpibeGFvmwOXKPugy8YGCWa6dy
M1fVothEwllUqQSiRnUeZz0/q9E8/ie0lfzieRn8CYtPNiXGFeW78AW/QMbGSBE1BVtcuuXRElt+
3tSEKmXW4Wqh2UCpRN7KTgcp6Ei+6vnMlSXn8kqOtmCahynsbZL+yD3rfGlua1PCryaFpxvESZOk
9w+wrXx5XS0ObVx/fV/yb1g+oVhFeSLJqmTE5e3nioBUH+EEBs+ZhVnY3fTYXyPCMKrND+/FlitM
kaQUQJqxj5ZPjUNvOMCUHfE1RONitqH04WxSUcsrQyE5uKMCPnUxmM1Lhz07JDSjMnWzxVfCL9Z+
/XuQtpVSJkmUiYAWGGuzcPgp91iYT6epaL36WkwNcJzOzrI5pYjIA+fXCQn0VesMEjq3zxplYamZ
zz2QLL5rxoV3kTeQaaVYB5IpN2CutMUgaFzidc9WAUV8uVBaAmXpXMHC5/Bl06MX3XSqRZ8ytjUk
4ca7RSEsZlkDOuEdBslKh2HyHEHdsSi9wl6CKtaPB3Ug9AmuOA9hUTj+7n6yoQmEi5VZ1sBtoYPB
PGt4lqDZBCOwHgtf9LCJm6vinPBFrejVqibLgGXwsZkiv2GNJVvlbPUYYvTStaUryDHDN0gwYXQA
NUL03aJ+LzrnOvXGZ00XtTGBY1EfHrfueeYoQ1CNnC1MoqjjyYdwfTltxtcNDR5YclrxlKgv20Ig
AxUokd1etM9LaKkxqVADZlHzqqghI/SHT3iR77bAlePVEp2nWTvFViEJyGfIVJd5jdrvzJP9bzaM
DuWx+zuQH0igA6Xc9CUNI7qCTtco2AiEtcJIrlhwgp0g3Y14gXZmnjoVng5rOe3LCmF0oOLgAfE5
3Qj4Q/bxqpUOpVc9MUWh3Jy11zHWo1CufSn30DcsdXA50AOtVpwB5ShjmALIf3Xt7IrM1tYuKfhV
iJoywHDfEEmABHK/Qb6OjRBOisPrGfVAUtEwMfyOadLiLOEmQiXr1aSoK8kA2bv1rM3ysEQ3Jzcc
IIncJ0dkes3Fv7p1gYciiQn5s1o1pENUJan6+bUzpjPN4dnGauhHjoLAl0WOisx/kirFCSRJbhi6
2CXB+0Z+Wf/LpA+8suU3bganH0ufIXbkgx1HZ726wfLIfW19HNW3WbFyX0IU+WPq5OB9XaFF4gPA
G6ckR3VRrvrMWrC++J9z32nqThk9YbNauvb1IOpRLoZX5AVLJXA9xiT/fLkUy4duJt8HVv40zVzd
dn2uq/QfeAGB8nnAEdRw2Ff7lD6fJusjadYxWOCwPILzECAqRcqdHovturth8bzJJiWsPXch3ZlT
gQfSgvYA8w6bXPP2MbaW3uHOE0dTRagzClXuWybnNkXOGcSCmoVizhKNRGYphSGyLA7pEhx+CVTj
5DYUrtNYhPEGBs6hdQn57wn7Y4ATqJo+/87zdVnHtGjIohki6Ds3loc4PPLR/rLGeyZ9HYM0NbjY
6xskPN6/jr2loKEcsoe7Nmyytod96o9rNx/ZJkDuM3w+giP/k7W/iPjHW1ErNbe3XffO1C+z4Qy4
ysS3crTWJPrmqiXvbeXZfQwcWCM8CKUyrrQ4nP0BZYy6ohnjKBTe5Uklh8AJ6ZKIrTriVfaWsnMg
7jn3ZIiGU9v91mGkB4gmeYdO6ImMrF5C5vSpERYqScUUVJ8lDkEvo/U9f9PliWHWlpMMdyQhd+bT
0E2aJNRzsuOvY6TIgvNKwbi4Q4JeVnzpouLq/Fp7qhV2pIA2C+l5oKhsL+7pSZD0i5M3yv/y48yG
7RVu6lfJvS8t3fjQswbQptsuWOmUtzKxKd5pdRbrdSi4k5pYSAEk5QKNduav8kPnYth8PXDJZwEY
/vaSml6c1LJ677DUW3UuBv9LdYTWl/t/2idxpP4WGiadULGEf3Jc9b8B1uYGlH1Y5QZq6oCcpzo/
tROAb6yAmjjrpZogUBUGSJAXaGn/5/dpGbQg30hVPj/DgPMVVQ1o4sU5L9YrVt6HAaNN9GyNLvRV
7Ewu9peEW4TuWBBeiXmsgRteZFtdgeBE38LtL7PJFf2B4sv/bQvP0RdbeRuUOGEyHSAN2gpVpP/S
sMDRAztt+LzMwTIsa87iSRfPdRZfWx7/TlxZ98GycsLM7IvLHfN8SBFOq7QFjcLYty7ijYbnZlv1
mZ+CXM3m63Y0r+PomDEJGzJ92QnqUTJubFAmIpwfyhsJ0F30MomFOoCLWXROHnQw/XclSzAjhcLY
FtNHt8cuLCZ6mije00dlykC4BptuPWfkDOTY+U+VSrBb7jDVJ69nVidrTde2gd4qn3AeQbN4ZWYC
SDUWcIOSjXUqBJoNvvxE+XE8GGGvMe5ngalue0eHumzhh38k0kfGVLfArmPlJj7kHQT9s02DmqDW
LPb5YCbMalhSRdJ3bA7lzf7fy/UYcsctarJ87/H1Pig9VnpYDwjcwtfz4rokoAVWyYzj8KJ5TzsZ
xhyEJFAqHQ7Z1UXFyiXAsB9s5Z5SPg8Nf7dS9mQJRwGCMM2U7BHN2BEFYFXuMLuKYlDRqCgVqRsO
R7Hsm+RjL6S606bRhjab579sjTXJ2D40bgnrKXDeWRkSeMCSCmECaARxPMZd3LCcb9s1LF6j4XQ5
8qNlhbIfUY8yStcCyjxiTw5ZFH6Y2L8YJ0rLGkQ8pdBMRvkdKCGQtZWWNeSm4OnLzE2rkHLC0dYO
5e2qtt9kSCM3EriBYDSP7XhpL/ohVWXs0C4p1KVFPDedbtKZneemoC0dMIs4/OCn8NIM/inMc20T
iIbq/8p1ayE5F3lMFsZ1ZvBD61nF2nWlDkGv3HCG/XuGOKqBAjpaiifyR2CzRzewY1u72+luVlj6
NJfKWDeRPfGfdVPmxQTCVHq0oPW1hWKEy4Mg2a2ETo454Xd8cpa/qkL4LX/ccpTTz/mP6+XjOZtK
gpo1KFU57T0J3KvETTcjlplnvoZEiVapfyY97Af5Kq0qT03wMuH2eKpNP2pCUnjotKJUFxIp/AUv
PkgXJvaB0xI9+HlU8eWCNmzCUMHE2WvmAsTezCSOitH6TwYIt3bV/c5ygMNkarzwqdsSpDQPjL+z
vWtWWww+/Cpxqq9W/8ZKk967RwVAgnZ4SabwaZD4ZMMSvkKyz9caoowojeJL7zQMogPfXYs2l+C0
QXafyMowxiyU9zKArPyzlBs2MiiDopJpGEcH9gExM08QbbV2cFicVIjbQ8flrIw/6yQtbb/ufNHL
tCjk0A8Bo/ih6zKeTskYEak1IMLRv3SfF0S4Y72oTUJynW8D6VSSLF83fODNoCSFTVAWWHRmCd5P
VDJkjZ9YPrmGYMwpxnkQ2vXV54jBtxf5gFVRnVW8sFFqsVM8o026KNa9/G6Rl+YDtm5TygOi2u5d
iL/IzgUnSij+TV/o/jA6SVhRIQF6go+C7VpuGjHpIOJrISAqajpa7Re4WxjDf0PAWy9jWQ3dFeMi
jfJOPNMnkTrszSARNb76TL9A1qmeHjSvV1bYqmuMz8f5Ol9IvPz6hLAEqwQIFRYYXXBIA1wxeUQn
8XAgbvTlx5MKWrHqpxzrs0xuN+n630CosG5Y3+HRNmDL9uU3hlPOxPO0l1v6jRMP886qjQgOH7jc
/RQlax4sLCLwb+WqiBsfkA131IkaZIeZ+ggWUyUC+IiQXVp9mURA1TX5tH2+eBkR045JKmqIiDYE
0+lqffVQAmHBiuN2BaRxb60ZqvE6XOUnd89cvLRVUad94gzNQHcGSmBRW25HL885uqgJunlMs/nq
ZVGnZeb+oUgEx2BqzEHteoDJ3D9i85e+ogLWaf49h1mS7HRFSK6W4c9+qykNdfVaI7GiH1nL25G1
be65u9w999fbe37YUnwWe+xWN7G4mAEHgLY8mZgfh3KyB62CZVCH6WMGpJVD4eePkOZMEQKQrKtZ
VSBeMg9P+TsmAXRcVWYvD2tmXxr+mRBzTN/un8ayWoxc0Qpe+j6S5y3QNvW7V8lo0CuafwwujOch
BgbbqFpyN5S2Ni7WAYeZCGr+iAPg8gttOSJ0H12S5PJg4+sRrIhSJyyyzV7uDmO59DKpOr3x/4Bz
3qeoE7AqfPwXGRXnLX41ZWY+0Q8V3raF55OONA8UIiB0cWLEsqgnfQLrwNn07I7HWY6K4lVQAg2W
Mxyj3RufCaieXpWg4GwFoHZRPpBn6DhaGe9pPRoGSeM0K71AGp+ysKApDF20Ccl/N7FS7WxxzOLH
Lr/UdjeKFTeTcpck3CmOsHlu2lxA6ihHNSxCWuD5CFxYQlVAGJcfWhE/ZXaxg1buLBBqcrRHAdCH
kzCPicDKR/yC2ojy3u8EER5iBl9WTDvDmSki894v7ekjS4KEg4kdniy8lIEkdJOS0Jaa5CRWMDe7
0riWMOWQ/+QHrB0HRlj4jgpR4pAxsgnJRx6E9a9oRqxEXoTzHKhf2aXbMvPN0PVI8DXsY3cf6+Z7
ToUhhOgyX+Ra2Usr2ZXJj6Hwul18azzSH2qrEeEG1jWzhE0Z/bm66Fui6bJ7mij+tIBN4N8nHP/W
O++Gk3C8gX4lfw7kQRLljO4EhKYvxVpkU2za5IEFrYi0LhS4bVkGopaiK5xrLp9sAMTF0jqhRRhE
kXFk1QlOjU251MGrQyyvp26j0mQnf48hUQr1v5ROrecA4o4MrQlzaZ0o1NKLNgFApgOKYMVJZMHQ
vAgLsm1eUG9UWNnz29c3HSH8qtxTr/5ZHGVXUMazeBfeUZB8l0bKT9yGKAoZLuQ0TK2duAiCRBKm
YTYRcvz18+rqnnyIAs9eECOY4YBw+1yrCu93244XP6y6EcoAY/uWLGuF/DFJqzQJ/5uagti+27Uo
kt2PzFdYMMGC5FXpIrhDpfoyIoIDuQZbkpLsE6gXyJbL1ggLZzjAzhnP0r5srid0Nc1L9WhzlJ8p
V3LWXg9TMnigUaxwL1uIRhg60uQVpr0jBr2IJHccpDyF+FvtvN3DIvbC2sw6FIUecO/lXTTFTCDc
YRi4GkPMz0EkE+h311EhER1T9mE1S2dYV8OCfJ26JCRRR1joCSTe6JZuZikJHbOGeJbWxBmu55b2
VYfhNwHeYxK7j6xRAWEhBM9RdUtDejhu1fS5lyln8SvsyOU39Pzkxwbms4Ic0xM/hS4Uakt9BQuO
eSKMsNm3WQAB9B1ZTqT4uhJDQxBcFFAHqAPNjTxEbb7u6WebnZ/8EzSBTWfRLavsJw/Y0sIYshHE
y1qa+G0T6h/EIDIfilL8zWrRivv1Rv3djoSmuZ5XLdCjdmCnuS/49DS7oMXoFdT/nxDDiFT6Anru
QNjBS3DnBfhyvPhAes+XNgMdF2OM0+hRgecwYh/z+Y0w3FCAZl3iCYMg/BtRSmBNxf4ur2sZyCyo
T3pIPZCfElNKyf655VsJmik20TL7iTo3bpakLg5QiQlQ324S8QLF18LC28ySDOl7CaoKHqMuDlv5
vFO22nl62vacGdD9HOA6xdI+HtIv1TxSR3ZW9Z9nxzSLX5we8rpsL2rcVVHDF8V4NODK5Ygkbwlx
71PnQXB/vF1kK2yvZydvTe7WoUvopQPqJKkmrNrzWtyjPiRLHir2w0uvvARYlQc6BkPJ8t5MceuX
11zLFbDD/iRSCErkLrzokj4QFW+bfIpvDGlvcEryYrSPca0hfyKm2K39j+VDYBYSTDZ4u7BdL7eQ
eUWioWtSV9ah/GEFhZctEuz857ohP17+2ybBbuH8+VyT+sP2Uq8X/K1HRMlT4Iq9TiSj5Zb2QSbU
6HvYRaaiE1KkkM9PtlLc2Y7U+381pnYNfhjGCO5W61XLG0L3EoV+pNRWVuJeaQI937CHbhkraphb
Wk07uuEgzfFDiNBZSKKpFDhYz2joInngjyXnwGJ6iNol0aLIEJZEcwwA2Z4VC8sriep0GyvkTM/C
TDZ3PUzBsrhWOBPJz8GcuG14/NSrkeqE2yNRJcdxIoOsCermP9fNCUIqkH+Awq3Xi2hVkv4JgWa6
E1OUSqEKSdU3AeeR4WL/1G3fqvouzfnJzQzPzLMet3zOoKoUqLe79fLYnUlF7ZnU+8yR9TQ/wfw/
Bba/QZNRwqrFA/ss956Jky6A3psiyINR12pzA+8tQs2/pGjg+ZcA97k8CD+ky28GJ/9rRbw90w6o
iGreI927lWs0+A4jfyNdMOOSIlrYItnK3j7/3r3RBiqcSG9BQYu8vqtTb/wq/ayW9mLflcEoD+8E
LuWKu+FkxbI0zUvSJLfp8nofbLdaKJ/BXOKJK35HcuJRYP4KricKQdhBEm/DfojGz56qMm/Smv8l
Tl/s++cLwB3qsyQUgwcCILLI8tYYYsk07nAPWIBDAdqVDaA6Ut5UCXvxkn5Q4rW82KCSUzYydgdQ
gFBEccY6RvMDcC1MyVi4KYm+ED96LTKVu3pZkZigA+7kohQIwNMAk+vsvX35W4d50KKiY3kkcI0A
5TcE7OznWhHHrxO0mFd7SiLHEupPJEoPZqNyKucggcg/gv46668YZqBPbMCbZfWVoEY7wIZxXBLp
gXsOGYCE8KIT6O62fTP67YZ8S0ZMIK0EXiX+vVfp32q/ORWSCu2W73JBHTutmli3xSUIExRYM+AE
M5kk/lAaWnaZJ09BlUNL8isZypTmZWLju+Zh7MOTCC0lx5M2X4zdKy/r/bzEYHdZ0yYR+BJ5Q4qZ
TeYtna5CnnxoPrKeTUHELbrcajaE2XGzk+RoPM9EN7+2hooILr1E/sYwIKChS49a3hNPAup4IovB
LRVGpQxU0K1/ZKxD1yY6lLjC0ngzyvV8V+i1p1mtY5TeFzbXwjr0o5i3+fqYYFiOW0INuYxTCJ71
ut+1p8AR+5++t+eWFLmUrZltEaS0/n5Z/EAwk/OzyBwpUtJoCnm1TIf1A8vr2on3KxjpBytyz7UH
E9v8BAugi+4HLsVFTOVj6VnT5TgcQ96Qupz7GGljh0VxO4EZ2cOiIc6OfH2SZEPaKdPyfhcD2+55
0BkGRkPplh0ihR9lJHLoCWXmp7QxXwjEy61xtOKsPQyXZJq/a1wpLu5PE8QV/HBslfxQeaxhfQt4
i2aU9NqTMnffUBOyq3K9+aw+wVcvLyilZ6s23HYjJohqExEUJGE56Pb6ABiCfgzbmqfBb6FOf2Dz
+bZAqaHDB9vmVKOt9WGmnLck2+xtSBCzOKGPnw1FLLkui8uirztau34JfmzQGOwGPVGlHWccbdpm
RzitRLCK4GYRNgjtMyIned61KMFh3DLz/J65PW8lI/6+ZJjZ1lbwFNLv59Og/vE6nb1aX5PP2EvI
3JZ35kEAFyRdBtuQQ+P7SfWXwr3jNhRyKRXD845r9vEx9RNQT+e0K/1Dw+V896S44eRClFjR9hzW
Yqxc9EprNpDjGp8YDzlvkCkSGpuCF78GN3CD2m2gH7T2cgxepEa8dIMJ7gtqQg/YHny3TZLL5wYD
vl+7OIUB+skyPVzE/UniFxnsOR4Okv8MKwbPp/jyp/54/ZhihcxF/pBfYus+nGvH8Diblm0KMQpd
enNOdzqzHFiR7W408Z9F1L+7tSX7nNthwEDOQiG2JRD2miQAfnAoYDQLvkHyRqfy3Ai571E5KeCa
YKFYI+WLBzp4VCDQ7U31wqU33qs1NdtjOBTxoGcjTdlFhnPu7kgcuhNN6ccLdDjXJPM+y/7jFVcF
bM4wqkzgX9302tnFpInZn+Qm4EzcLttWzOkSous8E7IGW2CxTzcEhUHDsuZ4ZdK+Q0h8obWyo/x8
4zN8J+C0SqXCShRkGzrcwQ1+wfTAdcqZroUIdSqXHKfgEEQUtqV7gOsIFM/hKwQx8MvPc3yAQIEj
DksFaPUcdUplZ83kRTMlObpnoyK2VWCv+DSTU9YE5iKyvbNTJUe6rbotqT9XCZr3GSfGaHvtYyoM
WJPtD+Qq6ntMhFB9jfIVLxgrTEjvLjbLSYAMsCXvTnaTtB3i3hik2p/GjBCq2sBlwg9J6bbSkqNS
tTcyVIUYyQrYAMp4ILs4tbYWQy274usq1Y4SCdtN34gi7lqr/8xAVuc6v9Wnl39NpD6C+4ZcSpxZ
K9NFgSw8XFmoEAxVxZceoUGSyBzr7wbzoR+pNCUU4fyA4lbQMpwP9o39gwslU0RjIH9Aa2cSkCbi
PJjJXEWlurO1U5eS0H2lwtTOL9sNQK6P8hlWjRlC5ut8fjdjw1TFX0V7AUFA0FUk3nD58cJvQeF5
pVxUnsk9g0YzpMbEFbvdJd+OGdCTMrmZkIxCeDhO/UWQVf4+6rJj1Mws95INCrUxtuT6DbihXUie
VK1DUlhB9hLLvnjnUavYwJN+9Z4izZHh+D3ZCPsW9Iy+KgyseZg1yhILvp1qG04QqWm2Iog5Gq6P
y/juDhO7knVNv1I01kPyNdcZFYFQ7yKrEqCgDCSMp6K+ZfkCRTvzg6Jn35SUX1pT6vS5wwva2tPP
w9qynKaL0a6v/85/XZkTPUe/OdfYEw85fLcSNW7x/WfXCgciVCLV7HWHmc4TUDBAzyZe9L2hxpc6
V+7xim/ZE3cMNFiRMwJVh8WWbP+vLfiiMqrqCiR9XaPu/sPErvvu2OpqxRDffsrc79Excs/IBgjq
NP9kHtF0wK6oXwJyCLsrTtJlS6jB62iJHIF0lC1PhKxO4kj5XtE6n7KMVWIVGIzFZshEhBifIKET
5sOO1sZ4KkgjFlnFE6X/oZaVu3slpMdgApE6r/jRapGQVyTetv7CWj5F9e7XYuC/INVM0Axvwt9W
A97r8yWzI8cLc7M2TqsAQA+Y2vvZ2cUQhtP1Lvm4tqbWmkegxGAwGLFsMgF2uHbV7/MTwB5+zbob
PVQuDfpCZbES5sBSYOhEd9AdMByCo5YKXUpB8IUMUzXVGtNAKnSglwPWptHwvx7nq4Y+Q3LZFjzY
7HvdGBkTqu/FCCyam2wiCMZQf+sQL3cgTqvjSM3dLSrWtsmaYLdFvocl+IF0LqW2JIQaw0yggadf
4hPKLE8CwJjJ+RFdXIFfsM1MYw0WiXLJ3bbNpiYwBq+1e3+oOMOefypEqN0hmo2e2ScXEoboCMis
YA1ugaOAQ8IYz/86YTqXmZEwxfstI0estRvD7u6qpDvk2+lwWyejJ7z6rd3j/1c18Fv848xH5p3b
lqNhdlR5PIVWc/vRQProges0UYvT55uxEfl1HZwRP15pbmL5MelZsFu2MRYzJ5VHhjS6bGoRNtB2
aekl0V9FXL4c7qy25ZiBaU/XYXRpGTR4+50kyzbcS1tZJ9CNZijlnCNs5inOJxEGW5e602JcAd3R
qW2KZMpK1e70Ooo1lg9MDr/Aepv1BMe07PHDXSl5mBJuwYyYGEKKnNnm1Tv92Y2itmhYw+lW7knm
aA7jfyXAyFx39DOnhR0dZTbNEWTT+A2NHLeZJQVit3XAxk5k0cpMgAmS5R1DRdWEdqoQYCd+DCZs
a6KBcjl+GLIE6Bba3Is9/uI/0aIRRN2X21x0+D5yK/APN6yTuqaTUrDnZ7cpzIEju1ofvjKfGKKR
8ZMVnB1GWEWZHxdVtFCc+bKwS0V9E0sijXfSh0T2QMcCiUmZ4wl4vWLsJbU4vhEybI/tQ188axb2
zju1smzDmuImwxAUMMQb3wfh+KvnxfpVIh4ISIjtVq8yMvgwgOA1BlUtRp3gymhwk5w3Pa3yKtpd
f6e0+G9KqTzmqDLnKbOV6UaenEI0Ck0VT1D7txRrcsGWu20LH3Wu8GthuWLrYezoKIz2l0QqWVs9
QW8g+lcvO7OMXuLctay16BKUUDJkCYv9W/S5pUZXtoT+aoaWNntTMAOkz2uFiyv8/882Osi1uijt
6YzuhNC0MkFJ6bp1YPoP8PeP2Qxg7LWdzAHr3cJMD9HH0fXMJYoAVRpsJUMU0nEAk3QsRCxj7dWb
7LSfKK3js6mlpZLFTJnPWcOk2rluBGUx412GCP+ekjIGtCEK6AReks1F7SmDXOVFLmiy1N7uqDr6
OqJ4itLH3+XGnIwnlZ+lqSZJ5VNNhL5m8LsQ7FvNH8sGSWyUgmaVviJFyPROSjsstdC/NpwO3wbf
LhGZ/UloA0vs/W3h5O9DIGjldiRVLQ194uHcz1+mFsvski84qZ3fw7CfqZr5DAam6fE0fIMu6PJw
4I6fXYbaKv1WlvVaMgL3aXpgK1Jic7kdN0MKTfvYR9VbtcfIZgCG46SuAiOpFyO+9jPp+aITzESS
sustNsQ1lvW1m1tJkMPBpeHpW21D722ZDMxJ7/uCJItn2PIqh2smAcenP63WGXd84XwhEwlThsfo
qUwTjOLCMC1nNxahukCvft4lLqe0v45hdZByVPgl8yWYglaGTRzZSREbSTLj/vXAXJLOrM4T4vzT
39LtX8Thr3LRPOZr1zuakRcOooioX6FmxUsji37Y7xDeHq/htiwHEpwPpT8jpt5KbPkL6xLJwkoN
PCE4t+OZ7Cjnb/6885pq7slEAERI5JgPB6xl3a6bjHoz6Csvuz8JU32GuFkLD7ryG+B29nwNYx6p
3caancVTu9PmyoIP9xoTSIskUMNj4ujSfHS39+pTiYWNCq84k6grtNLANPXGyiho61YVJOdQDIWE
t4SsY7/ViauoBRCdFbKQSk852Cw0Wx4H8OpqlbOcJuC46XbSytzQKIZSEelZrhqHaaCe4/y8AkWX
95+mUhDLnXj5iRyMIFXI8mNoceKaMy0f08kpiadxIrgIuvQPqI9zXPIgoCWSY8kt7GVVATWmIaAa
OwwUNdYKMasUYR5E2/IpDgxKxCgj+fNbTRu5L+QrBi2FOEOiFgUhn6vnpA0UYEUAPT8bB/w8ORL0
z65cLlNmV0M4M6ScWHsLH95Cb4j19MO8KUkxsUlpt5qz8mSHkCc6INsW9dqP9JxQPLPoN6aFWxZ3
NZoU9Z+0gGKW/eVo72KCYbjYlvzCS6E5c11vIaC2wSW+j3INk/61TKWX82mW9ZE8hRnrEc+6hd2m
n3gw79lbY2Tcm40prsDUOEImzS7X10XJZgcoIfe3Sxok9tUQClERGZHLqJffu/Pz8wd0mP9/7fkB
0qU7Nj/iosQv4RRh+wveOpWS3tsO69H8OK1/fvEWkivINr4pzyCB83GngsuD3EMoC2fP6i5Vh/NL
OL24fsnDlKZfpF4DiSZ48rCubvbR2yMHuNgj4L9ZIhKVr90/wwTcdc0fEY1o4iQT1/C6gn0nk5yl
rTKoNHpVH7iNIGog/7oe2TwLS8CUal2iVmnrjPNXSEdoM4hqFcJ5+h2mQGXvwbD6MtiEsKfN30Cg
GtpNTe8BFoKsXr25mD+PDrzV3S2tmCLKzC85Rz4Jqi4nMoZ2X5oa+XJEGCF33KImAVDfowLJ53xc
x2UuTKgLdShZLln6808JaStJCeYcxBPdrYNUNWOQo55T3lFYLcTrrRrFGSa7/iajJyI6/iVS+ITg
pDhA6BHZBzTyyijCJbUDmB61usFAnwJG7nLciD0hS5Eb3P47O2/5Gr+a6SSskCuiyshT/Eb7/Y62
W+//zYii8EiyKFlno17ypvQP7HSKsjmO7hT7UEgKsfZZnjChYfT17WOv5MzkP4Tn+z5qoFV69Rzk
imgcFYtYyWaOveEIA62/ig/08xmh9WsGxD47ohJgEKEV6+pFe0IQDv1LIBeOH/3uvtqUDparaAEv
K7xH3idWXulC/3BWLRte/KzXC9+b4H4m5TNiANpHqBR3gr2lQR5kq4ZgHeC3B4BUlVmzuwK5ERBf
nR86/+gVrqPBTWsEaS4To9g1Qgf/fqnRbLtiJPzi4ke0IsOIGJmHSSoGQILr+l3GAqhAjp1TRlue
zALbl7DgKo/T8AcIIRbW50GeVTYDwsqS3ybdzbb12AjRZfkVGNhckXSbfhPOiI2WNt1JlYOQG6bK
g6tY+tIdHAYhp/WGg/QHV3DpRmAv/rV1jk/pZKek27nBdbgdeLoSr7JB+wi7bAA8At6OdS1DFl/k
hBZcTw1LyGZFNRsQvSvM4vqRc69NhigxM6eV1cVg+/aQaOgOMDS9l7VOrTIkF70Lmr6YYZVLKBle
cubOI24reK/IKL8DKFfMx6jPq3Cb/T4SInMCAY1l7lOrY9Pp7VbkFd724wqNmB3XZ1AT+057mXVK
tuOz52X7pvfa4Z64BFDzAJMn07HGrAc+v4/lKmrZFW+HTtriSsDqoi/YnWir7HtsKUpom/s2YcrT
T4PFjjbQBiCCZ4QWRUEfUy/mhZsKcRbmIKClVqHYqHLt9ilelqAqpL7EkxK7A+66sk+iGAJoCmlr
Y5ZpU4Mdzji1JhnIfdw/t4ZEGfdAWvjfdxyhO6u9rBVxfrJ9bqELmql7Xg39Bh+8UX6p5C/vvYSJ
YY+G+j16+yYPJ5wpYWC4ZEaxaYGDGwbGdPgntk2KsBftSqIcwYAO0E8yIIuUwBossT8l0snt9c2E
lhCAbqT9hkXAktY/XVTWBXwzuPu2kLQbrnRSHbqXyPvL/NQNSqfqrb2Dy3fj/u5ty+fIp6948fO9
3joAlgpsHYQpliazoCah4FWV3Hr5acZLRtTBOT0uc6Asha9yKChqfy+7qPUzW5Kl4N0Lo11D/smR
07K3IkMAWDdfHwRCMgCUJWPMEW8efiThUupIrzybiMHDMPZDvfObXm/q8rl9X93rxzFWyWY4ZHNy
7Lx4htaefgR4cVvCGgtV9nsRtuq8zFDmrL533ASrxiKlku8kuJgYWvVXiwIfaypen3x0sKD7/2KP
EzY2kvT+3voLQy8gEOGxg7T8qBxPXXRHtTWoooRb/9Z8kUQSEzBqeSSDArLtfjzw5Q/1AfYxE4Y9
hvSZP/aTJvui5L/8pU3JviXBYG/61pbauKeOf4CRdwFE0F2YZ3XjePPStbx4ujs2kYI+P5ueJ5at
LRXseZBp2OvtuXMpdI8hZI4QAzaIvP9yOWSY4Gxx67XiuXlo/XocJxcsYqzCxg9/owt21Pa87CJP
nzlPa1ydeUwHAqfEzyVOEqJ/0lR53jcNT3bKU+0nsb9/Qqp72RzR5tZM3ZrXl+3J2R5uqcjgd+gc
0hd1f75vrLlNfRxHVO4LChwwXyjFeFXZDFJDIR2DRD6mC8nTZvOYz5Os/TOuxG+jP3/YKnUnajwf
aUcmuSCB2hVGxcTguybknTFWLhkGIX6aDca7SwvHuxdFhPXQSSKk/FIRf66oaMscyc1m6mJxbcLm
dQaL2weeuFy0JD4506LP9MmSGyVGMXzGCIjYzufHrTqN+/kYeaQJzkayS2uQiUl48w9/+KOTLNXo
+3IzV78hvLWfj/WWpy5Nz3rH+qlokis8aT7OcmivYgLeT6WMpi/DHlB1TdZLtJlw2zUh2/NxFnIF
A/euVSu4ZbBeDqQraIwVP4k8kt7TIVhDx9rNk3JAl1ZB0OW93x9QKDT0cFn9xRdbu3uO+qHTlEsK
qygO28FoYGFXVq2mqPSh3T1WTp8mwOfmen8vUaY0wtnl8EZR7ssL6hy8TYVrrJoEo81mlKI8tnPp
V7G+zNYcuEY1JgYcrIzWHer6RHrWmlOYpCvpw2u9ZepujonDwpAEZJxTieg6DdmF+I62/99XzqxG
JiiF+FmIvUNdy4nY0srYcQfAHKy5Ki1PTcodLAlJHKJXFo9Olypvy3GWShBIratsHNPHNpOosU+I
pEiW63HEFjHs1HX+x+x+E6t7zjEi43jleXmFLiBVYNOyserbYDsw3UaSvKrcmdTLRdbO5O34w91V
C/0imUKn5AeagSSxfqyYhOSqRuOtLRhdo73YKtHAOQtyEdZaBjnzmxW95cIgAzmcaBuH3Ls7IHcj
Qe4sG7P43yGpRqE6J+fPQZyCJq31tELnEU5M0xCIrO5A/MPwSlzD54UqAQmW/k3n31BA8uuBM0+4
iBEIhQwfaVpemFXN4voX4FNct46bQKE/mKg2mOuPps/XX6XhZIa7CjIm7lyT7Lqn4m8Nee371kuQ
XnLTJGnedYbRrK5F8P02GXiASuzlFBCEJNxSmw/SEyRFysoci8JXoWx5jZ7KjcX5h9X0rsboRobd
XwAnYcDyRSU2pZKKU1uLJsgOSFpmM6Q2SmN0zFBrP6nUaDD+LidbpOCDSztO5Vlhz5iMvCP9ahNM
CB1vowOA+UW3FuNeIyDLdM53sBNbvTCl1+k8fxWY9R79ltRbQ0hI+czIdY66OBwTuXSpYhPd5gK+
tVzGtMAOmw6sBWog9oNFXk6mcCHu6oW4yRrvJTLjm3c9d6nNLow9DBPjI2GIPLdyVCnv80znlNJG
rFXnXPOlGhEbbrky4hYDoycXmJ6GIMYNKa7aYqiSByCOoxFy6d7O1BF1Hxr+S4StXTliq4Yzrt+4
cytfKYMIonzTOxd1/xAItmfDJ+dOUnANGIS40oBmrm6FoDYRHooix/lIJB2j06svA/gkN/HPWbde
j+xpZt2K91EQ60PJB25c0iWfFeDFLqE1g7Q3STKwS/6Tdm+x6y6od9klIcvLDSpuqMuqB3BR3zXx
j0sAv9/0wrlO7eb7H2M4z40lkX5iI5DN3vmtPGL8n68dXkKJH76Ub024J8+cSkw+b7imYqwzSyPX
Fx6zZ5fyHHqcSM72PQ/oOIlOnjCHvidPjygrMf3U51/MqbA5SYG6651r1nWmRX7g+3Jt+/Ayc0kv
0on2vCXWSZ2VMgorhAG44YNONqZVj+ITj6wdCLB3eqLKIrQb2Pc+CnWjjmkr/zeNxFk3tgFmJj0+
QQ44OF6ahDrhXGw2PnJzJWjJx1eHQ9jm5stt7J4oCjlLcdjQpkJ7qt5XtwPnEJNUdxl+w3WbdC5D
sSGbWP1CiLRoAelbRoujp1xROI9xSSXmzT8D6mbt+Sf74COkGgAnQLGqRENWrYs73zuUt4ni5oTq
7Yuy/i3H/YrnpexvDZTG7kQ6bl5RqlvOQe8ixyQcbmAG7zMBJiuIz5o0dsr692TEXkK/TUdIlQa6
c7YOk8vdtpLx5gXm/jwS0C5dx9yPIkUNtupp36iSVhD8xrF0ib7RyWu6LhyXXkhDZ+B5z7VTJveC
Z9D5ort1hliGekMrSl76VUFJzO5zwpViwBukIqImPDEAx0wCi3g0kR4DY3TcDIEkKLWyLjXZrzF9
RPqjEq2Ek5dZ9/JpYziHN//yrqu2L8Lr67UvFPfbKu/Fb1axZyD4lscEN2HAmbs25ViOJ3f26fMi
t3SR6MMaR1R4uVrF9VSAiIZ7uO9zNs1VslLV1pldJFhnUlcK/14ELL5ltja1Du3MEfl8BLVGjqyE
TOjXeu11ugkd/LS4epPBRk3EAyuCuJuBjHiuNoYbCzMKuwhNXvII8BM00x5SI5123YLEVg7xgOHP
LbIppaYvNYVRY56UIMSFbWlBmcI+Ph6pShi/Uwy4rSBCOJ4TjDRKqWflk2buegO3dPO9G7kdq76Y
L3wGNoMZi8FfGQnOTQa6wto2Xu0CTK/6DQ7ot7dVJzHNgur5DaA3zvqQ/6dLW9E3u2r7FGahX9ZB
D0uLHdGHLtep9RFEFCKgSf9eojrHY9ZMwYuqwtd1vSixG6sefPusIlihRJjNqmNwz/SUQTELy3PL
7sEmvowwjPpmDwjYy6wZUE9bL6TPoTpYINcQjo0sryb8zeSpv9mSoHLpRDTQpT7qjgLwxSbBrikh
j5QFZjq4RznFQmToXZqFVzM/ZEVWKzkra2qqrmDNSexWd7z1Dhak0eiXrtMDywSrVwlIzEH4I3Fd
gbmdCn6162UGZTWDDduMr3BqrGSG/4LxyoBlKcFqF02LwobPGw9866qlqM0dajmYnyXdqhvmVAYe
ilBmtn7z/9xCdn6x3wF4lg0iNz56rxDS6rMwcyGOWEAuTyfCXLHJEdDDGpr+CKnuL8DiXeZRAvwT
6SuBr+6P1cK6MWGpeU8v26kX9uIB1c9xtPfs26k7e3PmgPcAexQHDmdg+6vQBpsIk+YWLdHyJP5W
rLgj4jta1AgQAHs4lJh0T7clJC6HyZv98jikCIXibWNNrCoA/2aPv4ZtnJvWZ0E2a3+Nj999Myhx
M82/dJ9cjKNl2ae+/cjqut9iCVka83kYy6dnFqI4l/n75xWkpEmYwMMnl9kiF7wDdAXHGmdbsDQX
zZSyrhCG8jjasFGq/DzAsHYSGiYAf5smGuLRzzH6t/J/hm5QxVhbBLxyIQL8Vt4Vw4cN2+RD+SOO
R9b/kcGkrcGBtgd0kjy4CTxC5zK3BV10q+owGzwkX1dvgd3ednx9u6YYW9EeV3cgS2pqozd6zAHR
kDU0o2yptIYivtyQTs8jD9mes9FIVV7BR5WwPWltlEXdkzJpYwr5HEOf7IprIi0F33sT4raoM9L/
LTFTitI1Nj2KwfQB240Q9c008QVjcp73yX6kOzsoJULbaa3nbDwnAV22l2MliizM2j+3asp/Ia71
X23sINM9d9ieUSzv6nT7kSxYFx7+ar6DRmysq13u7xFFxdcTlred/ajtT9lZavJvINdfLnO+5+BS
7fYLT7in6WXplkUfpCFgSe5x3OTZpyiJjITt/pMHcYqFEJLMAtU13xN4Tki0ZzMj//6qScsZDKWD
FW1z9yqjZmm9E9LDuA3C0l+hlvvCerOEugbRsExYSQH3loiTUCD1UJTmi+0i96sZx0llQbiKas3s
RXEcIomBul2p4gPHTd9oa24n/Joy0zCGzA9m08PYuf4vCP+wlI05r5pEuFAcqdFROLvvXsYfg/7S
RhijcpMJRfzGq0GPv6xAPfuIgROT/3nImyD5DvwJ3CAPmUlaFs8vv6AQx0So2jwFTeqU93ZSU/hq
Tj409lTWWWqYNdmHLn4KxoHAGx9VewJgh8jL2B4uvLHhdSFoShqWogg+uUPD2RCVlCPY3r6C6fDw
YlHE/dBL33MC1vGi2222CGdBdSgH3Opk2bG80aCa5n7ItxUsVwAkpoEX9h/i8ijxTnp77h3GR8cs
zl/pERdDQHBklRKn41D1FJQ/O4YSbqGYrCFzVAoDkwLD9sQuOapRjxeUnV7+Da2uKyqKfZ8WxQNv
LVDu7hUrWc7GcaUndFOj0TyiX0VysQ4mBRkZsLAcC5msDU4MdCRnZZg1X+wwVLtfA83b9ODNm9/T
kkGZ/bE9yQUYJj07hGr8NgqOPBLZezCdyPQ1mVZLpUiKQJv+htyRLPCwWMBW8hJ4RItwV/KYcp5I
Byc2mXR8A+tjhT2IRyhOSC8TNIZxrq5x5Zs6IJSz0WcwpfyPVbqT4B1ze4pp2KyEHsv//+Hd6HqC
x7XKSUjvucNa9UWua+CgiyOh2IyBzwmdfJxyKVllBPq1/Vj2wVpYyd7nhFlTJOrykd7MPjBcQMoP
1kQmVIqCD3+OpTx4ASvXgYRupf9gHwAgflYooIQyn0+7dlV3wCmDucinGCGx10AVgnIUttfZhRLP
+amR1lftq9ocqrNspAG62waSDJgHMkE8hCtagrLW7NpDzz3XQoBNbDecn7ALg1t0l4SRUl/cR3jE
z3FboIWjHt21fJCJpcw/HxujQXkDzlkr4x/Xwh+9nFUdCj6Td8Jwj2HmiuQprWm3djAxlQbyqMaT
eLepquw7B6edp7AA2JtriOeJjRQG8u7PMXMYl6t7stGNTpHBSXkYM0/9D5KdMar/40Mc0ceX+yc+
oCYcfJs3y11UdsMpvbr6MMKCsHYH6MJkI6E8O6gM8p0CVrwsug7CW0FRrDg2CrGkgmHb8bIEqr7b
io4o8qBsN3kyUjpSTb3bVni6bvIqrAK3JHo3VlVhjw/U+uSAHQ5tFwR+ioH9R/cQ90Bc6sekKgHz
S/T2Ch0HHtsyTkr9eptQdrc2QtVm4zOUvKolsEH7Bxqp5eBb+oT+uo7SXPYQG5Bn8bpa5TU32ktf
4WuBeuMmWKP39fjVYhG7v260rO6vhBiFN2flI7e8nmmbUGndxcVcPJvDDEfeDefuZNBwg65qoRfN
sZtRQVylMPCXewt5B3t5RUlRQ1lOUod/LYrD09cudCkpszQXc+ANIJSzIZiQx11VVnTw4TzH/zZR
a2TaQAbYZgCDd8BNS9GsfW1V12yNz6V3WMJ/O7fYkSmz/IuwCkgN8GmVZSZ2Im64Zu3SjthLkrV/
iMwehPIzU5Oj4+sxB+jkVs80ribNXvdu0d7Wyyq3XCrgajnDsnIuIlDY6ZDsMXMvydKaxRzJ5s56
cORXEmuHTYouGP5GUMGzY20rCyI//jn0WLdfICLFHqbb57x0geb0woOtX47sAUP8vhyDdXF93BFt
glPzHEHB87ers4ENwYcSYhb98jtJs5odRoJaY2r1zOKvfTlGcl8djDMFy21SMwhkOORQp9Jicgxi
6TVZwYnkYry3PYas/hvvXKHJbcyXpxYrI5EgioW0Ze9HYogO/m7IP8SOCedbT6Lp8VQMXd3DNgnO
jqj/+BNvzvT/YbQhBrnjr4wJfN51v/2bf019NJpnz/rMUyMCjZvlp8SB/vjBp/y9uXu2APPPq50i
EpiE7Jl++pNWTOjl/aWR4HJa/OHgAdMVU0jFx06VXirVUxPRy1R/3LxEcCCCPdS3ZLn6DjyXr4NH
9FP4KQVIe6qNgRhSTZ3B0koJ4C50P1isFsqEdFdIpQN513Dqwk8O8DJQwVxCp3Gf+KXDXuZxfO3M
XPwNAi7XPFG/cmH/AmxwDEzBx3FMJz1VLcmXVt1CrMWVh1FWwTal3p3Fti3U5Zt69l48zJQemVdI
jAMuqJFYPge49ta3p+k4jKPqH4EnV0GbwLe/+CbkLTRqRK2xTluoQDK6GiMxs6C57i4ZVEbXEXpj
XgWy8VUdP28sc7NeQbgEtH5LLKWKZp2C7W9mGKcQsBW2lx9oWCNBQPdC8WbUQcG4fbwhreijC6ko
+Uu/59o/VCKtiscawM+rksxPW6LukUSYgQ8KmyIRoBg3zzDpKgzLJBL4icNfl/XSXhDtmePMhK8n
zqlHxpjy+5pKqJ4koD+3D67e8656rPIs4vx6Jlp7jnnZWUzj2mIHdR8E6VaZipEB356OxPjgfMnZ
uZgFdKWbjH+8SqoPUjd+0kfnHy9tAeUX/5BhtVg+QWfA/Lu4cVBDq6uv3NLFxMXIOgqTo8ULFbt5
5a21d6jcZeFAmclyTOinRtQpFxJ4K0zLNBa6azgAMGe2Vv+qmprH0us/QkLmy/0mj0AxcgsWdxkm
Wa38F0lJWkDvJ/TomLzZc8S7oi8SyrqZFt/cetS9gzwATCwQhNhe0aw0jNALOE7O2+aDKR+MszPW
OUJsrpOuNGWwCG9MDb3lna+URY3KnSeHu6tnW4xD5gNZVp3N79b7/G/62YXneP6TWIERXbPY9v6x
WQTzEMfYH3vG2PQFjWECG85LnOKayTWEI0QlP7EOmjAChJcz0O89AioE7DGvr+BWH3ClyVIsrUIH
Ewa/5XG1x7LvLuwtFLYY2M7as1T1XqDMs9Bq2+0HoXQLspZ03D53dRuwYwa+guAJuF1JGh/KTHUi
rBD443l3nbvYTjn23xGQhKel6wwvl9bDK1CGXRPIqbvvn6ipFv5OJjlFo4oMJmR/B+fkw/hL4c4T
JmEwdWv4YF9tsfdq/giBPlx0Tnr7NbDNNsvY5fqVCBv4LGyvEGihWYoWUm9TcY6jfnxoUfb3qFSn
WQzioBUG83+3y3r9byMp68/VO52a/2+/Mx6wAN7ZivTRd0YszB/D2O4WtyIwdnNoqezApau8XDJ3
bPqqO0XWL6OPh/ntJi0bUwAq9AeWiLJpkkC41nP+BiKoBITsy41zuiKpNPh8UOybyI5h1pOJUtZv
evajGMkHbxD5jiNVJGazcKSfhedF6EhePNckmDidrNSyX14J1hduqdJziDqGn4NDV/mqMea+ZL1a
8rWXNgOfd9v8oVgzgwMiFC2x9zpfWu6jju7UzEjCqKdUNx8kOMnwScJYvsUyN9LR0NhKrQG2z8Sc
2LNH1kQpx1BH8VRwn2jEw7jkS5EeFBiTRYHlW/5e6WOr+GYThxdAyOz3ISAhh15tblGJgY1Vcc5p
Mx07dSmG9ipoHxTHP9L2ccfKfcPELwKseh3qvjGuxxvUdnSs1+1rzsb6AEF4QT9nP3YQjzCl+c+f
2BsCi0dL+hUa6Uwivo+cugcwCXA+F0zvid7gShRgTrxtF1r3wYjCeIYofmsP6zeIndXtu8vVV7qb
HI4UuPkjlglXeTDR9ZPZ63DLcbhADmW/v++TmezijPlrxCt3M87ah3S3LDpNPExXF5kYPw96ttm2
LNCqNzWyoSRVy1NQrX+P5ffToLQ6joequ9bA+jiSNCL0I0VE2ktZuedIA7cIygb4VM6Nl94sLx/N
fvytKVXsmP9oyXbUb8IOE/5n31VrWf8/O6FbXcRo46wSWseFTqVOHX8taZX/Cbb0HpkI/F/Bk23Z
jxVNkTS2daa7cYKmqxzIBvlkQtGNRsYJ9fj51QMS48+21iYyBjAamRM9IMHD1BwYLI5Zdx3SWkXU
pRAd6ylRJMtU9VuoAcCeZzdmjtjb9Ex4Igie5tyzYw1ddREUt06cPcxzUxy5IdKtSTZWaKC/yrc5
rzdLQDxaIhkuK+w/TopjSVxGyD+rUtI8+knCs8optbucmbX0Z+4afyQYOB+ClkYq2x7AqxJ62FTz
shVeBgbnWL7J60rbLab4qOVir3iPqo9IlVrtALVQfzIAFqeTyblNxK0xmXDt41uHeuB+dG40ZhW6
g4pLxC7BVcZQt1H49LQW7lNUVgxE5S6qG/vQpcg1W+OEUpAIgxKrXXo9yJYt38DcXMGRKrODgl1w
jofltZdzQLdVWKw3zyLLhgYgcJpAM2CcwOLYltzWK+ckd4YA0U7fvynjExcGyGcIADpDyjeaTCcI
2uruP0BYqrUsm5FQZ997CuZ1rnZWLzN5laqwjWId79kjEoRZzu7j6ScKwkYyzUKL6/2VBtnxyxxk
tePdYF+zW6xbFgwH6VyUivwZCrbsyxMJEvVV1aDXcoDlCZgB/WD8hdSP4gLxadfLzn+Kw0oc/7Hr
Zobh8YKlX36Eednd8AlhPgHNlWidaWJ/aPWNI9nMy+8SIdZJl0lbmMQzs+vq2GJqW6XRPCVDONWJ
541dHmt+Gk3j0POQzHLz0YNIX8BacZUhn+ArUD33FguGOKjh4okWcMTejm1F67qJnLSd1MF3yy2h
gk9I6RYueBWGsUso/F0hx3KJqqdxLTilHgFZDFlz4AWNz/rTsPWtWo9gGmjnPzT0zsRUezMzZW9u
Es4qjR/Y8GsbJt7Xdq7xA4Q1t5aMbfKxYT6vkMWnTi3ijsh9NErLbpvwWTnB5R4/lL2nj0FKTW6G
UjFPUfojj/EJ8DLVDctHX9nA5wPv5eR7XwSvKqrg0j4tMGODlNwW3b0kHJ5cgjezyRkkza5LELyq
iNkrEFpGMl4iJSUw9DGMXkUB25mUuave3o3v4hzX5DhWOoP8gzELtV0Nq1T7F8tQt0iSphEawVv2
tjzkwfsLYmBbg6CfJTMf8u+GYenQMSQqnIEzB6/19u1FIU34F26CLYNIvUFnESsAlj8xjYWyEeEB
l5hGKmCnR9irStG3RbWQ5kxiyqo0l3JOI7OeGtY8Sg5bcfNlXhHBzVZ0yNAFKAQ8Q4L7Rio17g6K
0pyvg/p3ZlFo+paFVOpCK9D5MCFmhiaO5tbCgww6jL63jed73iLf51QRfEgy/gb0e77a9/uLUhPz
kFnjBniiGlC8OLQKQ36jpdsOqQmuCQNPN/5ZR3EPk5E5veVjvK795t1/qv1m6EZfQvdC5ZxY+R4f
ZCSMGSWlv1Lsfr0b87vfCjDkxPrsQZtuygAB1QTjzkulIa+oqBga2L51jDm4k2/F1+2gq6eGBgD/
pUFgzjc9rS/ZZwbgBPeDP8rdJfmMoSU8GHQu8Gg+sbqMLlkpQMwA+da73OHx5h05H5FCfoSaeRbg
Ceip6ckmosGEKCZ4XcJV8tVet40flJD9leVwpgayIcU3i4usW91gjQ230db+91WvcmfmCSbCMwRE
BH7/KuEZv60EYB28X9sO48x+MTGEYrMOeUHpqhkKprqYhAdgqb/aB7uNlkm2ocKIscyLVN2/ynjQ
XXDLDLpJNzRm/9C97gPcuHYxPOOhsdiyWRSiQb+FScr80ol1KxcPqb3/MFBrdkM3oLPWMyiW9Wzx
mfbMwffXZdx25Wv/wroOSy3g4IopIosJQW4f9m7O/E5JBN4PzlKJIB7X4KU9CXMuCKI9aRJavK1G
J6OrVuYrTXM80tynJWJXJxzrlWxpSJEqWzXYf3XwVxRFHpLMdOixocdNq4UMbpXXNgAcxjZ/Oyhr
Zaaa4+X2ejQ98EsAxdb0C559HkVGdKVWaoeLGeUigpGnLP8XG7bPtMYN83IJbMt7kOLSUbv/n5uG
w+F3gpXrAkSdt9rByk/Jhy1vZ4jMLbII/oGD9M3S9Dd4AhEL4SoAGO17LnKYZizbj2P4z3zItLcD
5Jm0lDTWj9LKUfhtDXSBhvnMIUPBPk4o3MpzViKIKsLxsP7RyVBb2Q/0hiXFrAOj6zne9DS2o6Nm
I6YrdPZpaZfW39QSiZjWSCL8+h+WKgzE4+KBDT3XqilRRe+86xBnUGiuh3daZ2cWQQaTTX80DzcA
2WirqzQQG+ogdjFA7jchr5ZY4qsLxQQ3vnj47oSFP1yDMrbxjmuXbmFL14yrobdFbOi7dzltcygF
Y5ng5IMnd9upnORdh5DoS0TFlCQeZVY5bCPS62VzB4MB+bfTll1Tv9Dm1iorzPhIU5CEL3INOEdW
S1SwmLNE6NR5lg0vtgq0ahO6swP00J5skUN0XyhOi+U2ZDlwAvl+TllcvQZYmS0c1jruZFmKQTDW
HZ3Ru7F5JLba2ud/ny5+6NstepksBfEr0Vluhnic+vK+CceFHpDhD8uTitHee3Hv2JUH2MyR0czm
SKFAucZBi7cx8WCURcjFe8dFt1J//aWR55aPCnJjSSS63oQsJjswAnmHju2ddmemWWyVJx7np1El
l70mmR9rshALqlPnbe1JM6JoYX2iPEcewqw+AVvhxq2osKuSMrgWX37PvuHEVNxG82iFCYkl/A/a
Ee2jAyB9axUBJwcgv+wdiJdKI7oZEQlccOACnSBiOmRBn4j/Mivdq3+zu5NAUw5+nbcFxC1D/PNz
sz0zPamCV1ef6dUr9UE2s33qmEbaMegdhC5WaiJHClzXOrz7GFlgznZ33Tm02O3vTNFbF4thmloc
FpT4TfgSn1JdlGx2OeSNucnTq3MvlMvV7zddx/seLQmIlyRSRFRn4jrX8Lnt1MomqsL7KJ5hqDQU
0JbtFqmTxSrhYDp6cIsICsM4rLID8hVBUzMsX/RdlHydu2n0shpQyiYMaPe13/KyjiSd6Kbr5iQq
GCLyonbElMnb+GAAT1koE4h8BsquMUX5ZkvycBQu+jzfwyp6DgKCclCeHczc4uSmD4sPUkBba3Zg
iRQQYSHEB4vL4YIxNlsXrFQ1TMUSXB/9RoZxd9F8JbQbvrqYjnO4Y+4HCku33jedxEaHpFqy5eSe
G2dkWTGxrjvpUCK4fOLKxNY45LlNpgrjTP6VIETuOtDD0PqZbV0w1JZo45tGVbsLa3Cb+aeLkfve
AuvO1bytQ1nX8BKegdFKFh+smhonpbeUic2765YrAfsUgmM5sgZnVBic9nbGpRYKpjwXK9wcHH6F
UxkfA/+aURgEug0pYhhEYHQmZMWRk44NEluqtE8Olw0zqnZ/DZkP7MFKEfEiDFBf/db94rIEyd8v
deTCCLZCq2+6Ejitq1y6cdw6cWNTMTJHni8sGBLs5rV8X2sNxNyqc4Yehcda3A/MsyVTKdQvG9ix
DbQQBi5T423u/HX0+zvKfaFJQLZiFAYSOi7XGphmQ05pxAQVbyhh/GWvszAd7XhLdsGlFBDkB870
Tn28Dc0dMSoIIwWJJO1Qd8N8nUOIqGL3HtaYx5eyCjHkG/V50bE8ingETqAWCrSSyed+NvMQKUfp
DxhoAas7tNGvQI0dZOG2Du7i4myMcG++t7dTykwLeGoj0Ji5rGkMQASt8uugW1NTPFM6Bc7vSYxm
pv2Tk+euWPNA88IWhhIE3mERhQJfCdiClETN289xu1yDI1dga8t+Ay8U9p2gZsj6a+OjtNlE7OD5
DNwkaVA7AWoS1dKJ2u/TSRVi619OO1GmiBsZWdZVbXGTz0X+53qypP3J1UIH2s3BABm3mFEIZjjI
5brZaVcdgkhgKUXol2tVzwpcmrsYuOIyT2vpkxAym7J0XxeDOHBeLAgm3b3LuOdisjk2eg9fSjMQ
QQOelaBvh1hhjY2wXFO6ux34CKXpbyDUjKJrFvjMBA+2BgyedING4on32lADLfJ1VwwG6Iw2YUp6
hE8TjRI82EJWdlmKDvI821bIcs+Rr21q9eIO+3DLz4IM52OCWT90mQEXdtWNMjKNWpR0b0uiLmSJ
GLS109ohkNYAJ/RqR7VwKWBAxs846mg1di3GJj35OhUhWfvY0xuWk5Gul0yhAbwQ+2wIEoHe+3qF
/RNCvkZJX2YOfEbyXGCaqLtILDBTHandecnfD9QjW5YkbeJwVp/NeYk5rZDE93mvuuIVvMjigAwP
RUoCgFgbuZ/eXII7H8gU9atn6qrZ17cKawPFwEblQSTndHqioPKFT0b12vmqJJILeG7C1KIhNFK6
hi3YfSW+Uxk75F5RHYaK5N07v8mtprzUlbQSAmj0q+P+e+oBCVJ92PCtcfDbazxvhhwD6suoHEe2
99nbSiRhJcSQCW79nM+esNGcibjBjBqhPbyGbVRG7d8jE2hEyGZpZUVh6RLtod/4E7DPq6EUbf5l
rg64XNk7TPkbWUr+AVdzdPwjPzFZlks2EqU80OskdQcjw2yE27f/XKLD2RNm+ytR9qH2xpXT69QD
1zlaC7KuBCfn1Kjblz/NiWqYVVjIBIx2tNxvugNBibkc+RfdeT08tX0n6qzTh8/cquo7tVaZ7WZb
yewrid+x6j64d8Gk3AQUzpNCPK0sEu6bfCtLSBfHZLd2CDDaRfliPa4Ylw8+LGLk/iQfUSNxEXcI
exAUU1NqM0F+mgO8EgrUAKAbqY2HDrwgCIIm1JeypuEle0JbXM7z2tcYRU6XDCayEx1d5HcU9DS6
xsckVrtGMe/dtwvG6dqT3/9YMpGLeQ4O/qaRkBL4RBv+nF+dbzWCM9+ZPI+DmCExRlXzsGV5Hyqw
Q0qWvPTtniCFeiksGyMscDnlPzM4NaAHTH95/tVm7oj8ExBBBmBMM90biT8ChNBZID37JetW+Qm2
L/Y8/nl1UYUeTMJ2qmlVEtDnHLBNEuf7u06mFNQYrYQUgoASZQwRePFrnFo1oiQl7ZENsGovf4jn
opRSnFRD3bSQmLmts+kEWiayyiREQwH4MUmjEhXKdjuo/k77DavQwrsVxehvo2kfy6IaHSZBHMdd
dvnsPhXM3uT8Xol0KUVHanmO91j4SxvMMD7tyoX34MaI7ms1t429M10iafvEls+Dj9MWiHc6RZxz
oKmnX3OYGFItb+lfsf1thr0KUCturgA1a88HIs/cVvQ0VvGL6d6etOEEqC5BdK10JOWcU0rV4aJW
xhgJN3hZlh5B4REHbsExqDEkPnwkj3DGROrwn7pS8K6s6YpxoErPbw4Smym+YmF3p6OWPY/H9Z+o
J/eNjirGk/AyCCn17KeMlZyyhNJ79kiFfqkGTTkya65KcqOfcd4Ck01yU8h0DBFst1otNhKDBveH
BFtqssYBkmAAkY6Od7DamVn5EpFs62o71zyajYFUHVVQD4t9U5m+oyKSEAPxtwmRvyToFLCsT3LI
iBSD3720YBNSFEco05kpF9Ca5+GxhYz7+Rjl96hBye5tkvDaTATsZkaBINLaI4Ng2pS6n5Qlly49
bWIAkQ4EpThoi4Q4B2enHhgbUoYp0VlnBCKfDo+0NBLizWbzhme6HaeWt/4Qk6eR78o8GmSq+gh2
EjLyljeMJFT+5Gwug+vnZHsldYKvOAul4lh4NMPI5GHHZ1OWZtQ4MNRWxame6RcjqWID7RwutlIT
G5rR0/uRCyfr8kWiE8arcxlgmyuPnYTwIcnHPLJP9F6zQPeBX+pFddd/ruo4pbpjvnwAoSZxjjQR
KZ9qv40NTrugSgoG55wdXZtJg2qa/a36YnNUAn+CqkAKjG87RURXaTX4SWz4z1+U30K1nTLnirJO
UyCrsdV35+/LABDk0/SSooyQkE2ed0GP7vbjK/C6SEaSNKHs2LnvX/OkHBLwexPYJ6/UWXMhOlAd
p0h57vZ4Aiz2krjPzSR5cOPVxPHlISSqaFZclJ+/qc7G4A51NEPAO+S360CQ8XpEyQYD/paSTjN+
96Yzi4URAEVVilazL3A3LA0gxQDuxiTJZ+u8VWNx0gYNJ61HqcW5i6UoafuXs3oBfvjnspg1sqIM
GyxjbLv0AQlpaG+PE5Gw1jaaDPWzrt5ywCXjzNwixwj7cjnfvRQ6Kq91+TDXygzkkMIom2wvrE9E
t3hkk0wnK4gqlDUowgp/4FTGdwCSU1vXUzoWqZExroTgLTlSKG6DhCVJRPicGkgUN/xOSdvZ4SES
4mYhVzQrNLXMnB8ZF8ARD9ywoRq5fszZVXpW0cYgW7WtIW+gt6cwoevyPRfAzSmiGggVeNb3qEAZ
pUaFJDDWdwfP9NpuJW9hzissCAF8Dcikf0fxvigNYXxrcVkTtqU8QDjTDmWGpiDO4MyRRaDV9wPG
r7ivW7cOSYwZiw+PJi/4hneHvWqgZfPzEy7+yjS+ikk63qHn0pL5b8pvGkg9VcW2cLH30kpz7wGG
ojYDAvQXr0knktvVVvjkByS0EfGCIDYXII3IRM0AoBcSFZEcVzrsZ0MZDZoSR6pyv4NzHGvuvOHN
q5aZDCt+H5T4pHpqPRIXj05kQm/7j3JLNCkNKUUuaOf/jv+Q55z4pLJzpOElfy1IUt3FAxtAErjm
SJObpatz6sjh4JwHP6vI6y9qgeoG8k1++fsmtjX1boAUfGEJIXXv+1tMz1BWwUuVidYJIXXpHc+I
3SU2z9Fj+uIJYQLpv/e2lHWTDX2w+DuOWYXpogg7RULkAq3aUoAUBnBwRCJildkWMTBDXYcBJvTk
5MC/SyKJ1kKn4uLr10ZL6HN3ih9Donv6Op6wCNHx/6Wh+Gmmt9YrwsaRWg1J4TFWdLtA7xIwQDiP
WYo4pLGVlpRMn7xH0UyLl74k4Cy0nAAWWxy7e5OEw/F9Lq254Yj4QMj3/56e8J4bvoYPs2nxMqul
ub4vwxUkU1r03t9wd0HUMNMRvTW6f6HCNrG5KyWKwc2iZFqg6OMfu+hCZ7HByRZrIhyYhd+ctMpo
eDh5qs7PNP40xaT7YlwjxvHmSRAX2MngvnvQYLoe68jQpCCm3Gm5d2iFwL+AdeDz5NGt6LlmOQ3c
1Mz6/uYLC4Swa4jKarO3FCbAlQPzm2fqBIR4GT+cClSOkQNYW9tM8Jv35yOzgQSSH8+5ebfRzcbW
QYCCVb1Y5541DO+x0Dkorag7xUMTV9QfpbLsvKgBD4xTpFsqdEFZ7jFIfeiTD5F/Z6LdnKdHSNC+
UEwz7D+3AATeKGqoy7c6cyEdDNsobip7Rqo9ihlE+SHhK3m9YGL69xloPJX7W6mzenAeQMe66l0d
dsyttwrDrBbBgdJuWalwxzEYzIx0HxuwYxZqJaQFFGfLHU2RFjBg2DFs9rflCh8EQ4pv17Jqjln2
xi6MALDOAyWNT51cwOx0foDif4cMlrtAi3v5lY08iE6bydNpJyTcIB8Ugj+oSbyxMDAXpC+f+2ty
JZaeynrCuXnzTXBjfpAnPArmOU8wz3ge8t+SzaCb2y1zotNnyXSEplGlOBHiIeAqC8MMvlx2CIqe
5l7va6drji9U0Vb7PSjWagLcrqzV+2zdnosJfb8PTP2aXnavoRikeIYZGrSog0y3eKHFXdq0MdF6
8tEGO+kluROajv5igS4Wp+6HR99OWHkmkOdr3avD595ze3jQp1p/z7tAP3tqaCjjX2bD02vJdrI+
fsPfrwTqu7Wpgb6h0fBLxF6qmmnJFfByseITC1ouEpx1jQvNPQ96NWh9MtJvv9CX1NoGiGdQuOnN
LuTPziFyQ58tY7cB593FFfCbAsoW4eXdwHv7AbzO5m2MORRAwd0wimTJIKsFtlHCQJHcEhhKoxCI
qspsMDyz6U5cgKFdNHXWNqxW2HrUWKJkJ5kul9cg22+IApnxxKRjUdSP53MQlyM/DwAE72ER+zB6
xxW/+rOiiFaQKbwvCzWFVE05wIh+p36OpDSFNjUb4cMMgIHIy42spzKs2i4yRxIp/gFHo1iqsake
mlfeOULvVHMLFXITdTkb9ANKL2oyfCpWsTxs3/T+hYqlTF4y/kZK2u1g5/IxXGY1DDJ3Ty932bFu
zHtILbzuYuZwoONSurf3mB8PpGQ/n2ovb4WpxdDhmj2MudZib2DFYM4zANBUm4nWF1RTxe87cgTZ
jVabWH0wTREvn7QD82n3VF/tGyASfSo3ezLHEH/h8NlO17IQ6TlamKh/82CETlADTAC5dWh9SVYC
uoPSvZbK/88umvfA/ZvsrTLM2Dm8buaSxXrWh1WN8pLe+EvBcMzIOOKNVKivDkOS5dQfUkIrIsKA
TKoBl/UQGGVFqqCd9Ar6BKxsUniovFkhklfaa91onTeHGHiRq92m3i3/8xXtcq21inkzSDKM4SQ6
8lVbjBZP4Sj0lrIbw9NnoqztAUFmddNNIu1roVOXvvRQ5iNPWUIEHYoNuU86FqH9q0+5t5kz9t9g
96B4qNB47nChVstwOJHXPZnZWc2hyiQGD4gxpY/frZqKf/NU+zHzgQGKOuouw+4h5c5nnQkNE3at
rieIv7/bhKC96X84Sy/RbZqmbK0Df8lu2JqXcux7A/t4MrKWsP+l4hqciHT84rf5tB2znrOpOD0w
FKzRecdcpzdOuY+ct4a48rjUSSf1YHujMKNJEPP8qJhB28N3NN4Q2mBTs2mtUeJlMZ0ZCm+j07Ji
ogdPT4hZvUcRZNcDNivYJDwNPyOLKDXyR+AxRbksrWHVqKg2t05J888rThbnXtFaJUVMXjWVl0/r
JrkBrkRTcEo281qnd4jqXDWg4eDE6TeKOsaDd9DvVgox2WRi05szu4quV3PrLVnRU/hHfzuiIBAP
BNkoEaes7YDxYsn9T22jM5hdvV6zNm/P/pGjGVS2nIHeUJ539BuxO1OYCl8RBEjhgLChYBeXPDw5
jB2hZtgc5lGsvBKSjMLoDIvsiXmt9kIPFa6MYNweaXNdynugVtfPvqbWQhXOEhf59Bgc8zcD4lNk
cRx7dROUlFKb1vSR/1QFhSRkwUJg9PQIfyKOm2+xsrnyBh+EIxKpTPk4Big+tsFL2Y4+nfBveA5G
R3h0/SH06mLDwx/pOmFG5dXM/W7+9bpnswcnAVuuWnDsqverhZs2av03hFAy45He3Baa8k6XBGpJ
LwzGAiltXHEPLPcPwfxXJLOF2U38Rpq6lY4e7JN2KwjfXhJ/0XOZDhWUB4F++NK8G/s9ZmXvFv/y
Xf7mzyQcdfl1uWAlKYXsmFVEPyIv8oYXhXQrgf3UmAPe8Mf0bfq4kOV2TV2/BKPjujJDD9Y6Rftk
DiXmHnPeMCMmLQersy6ZzyKr7iFxlMGHGT9ZDeVRBnfBf5mDvBK5sr8nSvP9MgdAj1RbvP0MghWA
Pckmjkbv/4rQQY0p9YluVqjAP4+zc+DRAuvxhAylt7ZSV2ZP6vzDfehwTIchUFZvuzed9Rc2IjoG
iOdQFUSeg/uGha53cw5SZJdnO730DdJJk+cM6ttOfs0PQGaXSd5oD6bkJWd2ZrXRRw7TH7jDqivU
jZvw4jKBAq98wkCuhiiQq2YU6nUt8IUQDnWJ2GwmTp0Zo8FYE9hoDWt+Q/aqTNJBtj6e4TxgIX5i
TfS2//+IBOxy1ssEHX/QP4l/ay4gMY0ij1vWsk9gGo+I4YFf1dyOB3QSY/kJXCvRUsji8Du0c8OW
7e4+3nVRm3sDpUPy8EMX4k27eYQG7p1Hrka+aFTnFVZS57z5Ttx2ZyWl6gengvoYs219LIj8WjML
xlMvsPac1w2bbeasBAbRdaSWAw1b/l0k/RBwTOyzPLYK571Vlim7pVicvewffcmMlJ1Jmp8MZjst
Np4FqZitxYTQq+01vJwmf6KVjE7BRvYa1QMMKieDWYguf7+p2hMKnTTFsKumz25uS7vx3AfhxpcQ
+pYBH2VEm1spoqCWW/gMHEszeJilJQXWebjBX5AP7IAqYbutLB+jE0RZtD5N97CysTJtvAg4B0cY
O1h5qOwWPWPsY6J6Dvau2RAPsPpY2gEf/SPJHOuqEcPZfPnCyuonJii4J8Z50AMv/Bus8YtxG6Js
0AXpYiHI6Dn3Q4S55wg5teJNQQmW2HdHUqIFl4wdLSB9dvRx93dowsGKkpiT4DWb4TS81/zHdfnJ
MvWrBK3NHUsvSxkDSZ67vrG9T/8JIEZBTWr63hfTJGkrWtVDrhvwgcdJuDPV27No4EJ5YT10Iksa
5zknWVqwybzG1AZAOBBAs/46mtVoxFbJGSUkHVgmJqYSjWSiDiYJFoWnRgtzfudqaRW928XSciVY
u8G9nhfKoDDQAxwnGdKaspuN0PM7Xi+jrnrCoLxfncDY36e0r4NscCQqI8VPIexI3XBWohYZSQbN
C/3Wwhm/zUB5SI+yZr/GtKHL/g7yjnhz8BEhSMvcLsI1Q5/txwSx8c6ew2fMHTc/gl0Za2Y8dzOk
gWTtZOWfn12BuPNOUVo2XcqLWOu/kezFFly0gxNc6/x3oWOxIS1yKjvASmAP2dCMDyjuyt0Fg37a
g0k79H2Zci0JinHX+SfZN6imIXJnS9A0d7RP3mfsPRjfOTcW7ZMAOU9EAjRb8YK9Pgsi8XFZi8nH
r851Cwvjp4MDs1vod7/vYoutx8s51cxu4S5SLG1hS1r7BCOZEulRTL4hTUNjKmVJ75EtvPv73TMa
5zy+G28ebMuaV05+Viyd9otyO5k1zDiXQWMnndi46tE5sqHZXgyEkE16Cc/0N6aXInGgv06T8M0c
HY1nv3S5DnQ9M7urauOVh588bfkpDeFupFzq79VcujvD4MqQr1ta5JfBl87F0pq8/xCkGV+ZXthY
d90sry39SujHATZLPHCIvNwzLDWbML2UejwI5t9JNqx/xfwaF/gZZSiG0JsmLi/gXzR/T2hqQlhC
YMbZkzLHpkjJ6QtgRsm8xwlf7B9Y7qh8Y2OM+nQNewszbiKTQDL/4bO5t3WLVJbQ6C0FKFWDET51
pz6sJwmp2BK85/bsJXhz3wpjjWsnXSkOB5w5IRmJ7T/JJ7+EcjDN/eX6KRUrvBE3lRj+Kj7PkeRE
BEjbRV3Xn0qluCZq4DTTG5sWxVilAY4dgTaeyqBUV1zP+UdBFsVUtDtUijfGMy+jkxrJIREplB8i
x9RkWYC696lzPvZIszHA38p/7XoG316cakE1d7brB9XzJ2fljJz5Cm5KAQ03xhvF/oJ0NsxJ2s48
d/lsZhFTHzaJMB/xtiMZSWtPXvH/jJbR9UqxW4TkQfhaGk7JbWR7U54LTTBFKvdyxsyTh6fVeSkK
vNsj0d6PfIXXfWj2l8rMngplJjdiE2EclPuWHNr1qud/vx2tshAakPjP1LW5ehe4cjorD43Md/QB
9oFJUqp2Fw9nckRFtrOTXkIx7lJpnFjSRC3jxtYXB8BxiGwswsAXXwKPBIWFmNWBg7XIgyZ2X6i2
EMswLA9lc/6DwOxZmnQe2SgNKbdW/ynHt0QP0HWzk4HJA+ah4welbZgmzoWDm+of21KBfvYSUT0f
QZX1OKxSUTsO6IKY9+R3FASLDaWmCPJmElSaUJd2T6pyn4VvtRKcbwt7O4yJcKTOjD3vJaVirVcq
gpi3ERiYnpoPEhFC7zcpeG5KJY8CAY8aDiE2vd5D2yCK28FKr+7qYqSj3Co3eiqje90pK5esEaAY
dbXuEdZBxhckFvxueFnlMrtYmdlQQepmMchO30AGdhvlJBUsMI7DmZ90xwgIAVP16cq9S56hb8EH
kfjS/JTZYKveicCkWDXjewMsyVreJYjsNb0yJ0MJtJjXAsLXtZxES1a4dSUclADQDGql+aOPty9d
SPsGpRrltEZgCerJRP5hiJykAGbrtPCHXl6Harb0ikC25lr2DZNZj34+WRISlhukoLreeYfZlE5i
DAi4LKyKnidMOXq4gEfQlfMK/vbtKDFpmxxhFJV9TJc5dO2gFM9uUmZRowE+lFN7I/TWzwO8w7+d
4AgibM0rhb4XqgnBzlyYjFi3/atKRHIpXyPj2HxCbPou+NDId1u6FMetg+/aXWs1iy02R+MO8pMN
vdusjw6FhFVJv+ruGsUuE4GDbsA6byPMtCnx7psZlGv5cCW5+UKx769X7WBGe1pg3e1W/VtjegWQ
CNCKoKoDNMorfv5E3pKTcAQT0WJ94Me5MZACXxOkyNfvyIDfV20yrBU3hGHUzswT9BiSFNf5CjoT
j9YVpxKLJED0PWVG4uVAa2RRyt/KCkb14seJdkcsIStQZBl+B4d4L1uUcyv5JU6AWiTT1TRH87CU
sNoMw1LJ7GgvXjqZ/mOm29LUVKjC5cPTeib9D1Ym7KISuyxRQaMjkcziestoJ5ZHUpuypcAuLhxj
QBmVtb/QxQ442dU1X65Qeulb4gRSEL/iFjEIWqa/WHQhKc6gXvOSxf9OkKozsQtRNdlvo/vsbdis
4da4NFnnwLaC1d3Szg7BfT4344VIJftw0LWEuJ3e5iJdPo4PvPS1zq8q31JKxkX3hBXwVWaUmzQw
Jh5g3QGDfMUOxFCgIrmaxcDilA3eyG1TfSF+CvZk5dYmqQqFF9dTudAEiHFuft8nnr7s/UUXzxc2
X7if/HxnXNUN7N1Xh7zFMLNMEweKNWWnz6U4lm/GFkw4JgeVAvUuJy8urhpCMQlPRa4muso3vS64
/SROM3jxvds1u/+JDCX+o0z93mWUTJB3ve2dPAtfciVKZ0WfeFSl3OoYup3tGcZGNndcmoYNMXFt
pfvXT1sTX5GBP4RazuvIfxU9oqCsjVZd+9rHEiB4ktCBhd23wLdtGpTLUB0V6gj6IX06r/OF8UON
RMYupeSMymNwxwKqMEl8SemZZzq/y5IgV5Ss/RP4YjasDUNl7bHJUpzKuY5T5PQSt2el/k1zzGHA
0XjpOcoY/6f04Gfg9JzHj/3Qrr3q9C+IPCftNxm7xmsQTC5lNJ/E2460B4LmO1wxyzHTFAYd88bk
bh8ZgPgEYc36hMdPn4sYcbSO1PaCnTZ+M7t0eIoOu9rfC/MH8RZo7A+drzbgX6SXU3lqm11X7Xsx
pEaJt67LgCJA1jnfbN+goTIHQFnwuilBKwyNVPpRW6FZQJYZRKSV3Qryrwp5PHXSy76CBlCxLP98
3zH2gaiGGbOzYLbEDRDoiFOznCD1YEYCnBq1pnhTwaTvM7H93MiXg30cbnsG/riJzrQtIjswhNwi
VewbomlIWizRBiAPTmgL3S5kWcQ5YpsFoDRNdYYGGbM7VVkUaqS/HnAIuOY40jgBcwJP1ll/UljF
Zgdze8mmqYigY/EVavAMqqK8lhmyvJbY41cyb6+MtX4Qy+aPOa0bx2Y4wQGvCNghB8YAgFETjEG+
sbKYpW7vDio79G4V2KigMg+jo8UOeRfd3s8W4UrptzjdnHPoZvMqGT1bilukoU42qvXvZjDElO6Q
Wv4akO5pyPda06ca8WJjtyXQTR3HSXkLB/sAPYuuYHbkOF+kYS0cy35xOylVNLRVldtvl4Assozq
ElHKeAtYURurpttsaAGfZ6DcdiqoHHnoRfhc2ywM7cHmgIhhCmGI/SYx6gZYuh4vN4Pu7sOVsrXH
JA8tWpWH9jQ5p+nvzV+ZIY9/9NT1JDG5TczIJOVX5KtgPs35J4NlltCeswn+SH0YXWbR9KA92LLp
zFekyZJ/cD7aqKfLqyREvNsUrolWomE8v5h/0+vzPE6Si4LP/wlSv1QVrpblh1xypP3wvbZpK3Hy
SY5XUe2yOxTwlcK3vm0pt4mJZflE2W9kLiElM6PsP72jZjDll9rgwCKC2H8FTxm0DfXotjI6ITwl
pdQZ9ak3QMFZsz1+fd6NP14OUZ9pbKvEb7bSjcreIfk+cDqKpYgvfLHUHlQVp2wXizyPK2eNJbg5
3JU/OVjY7ELkWC+kRvWM5U0sPj/K4QeabuZjKnMLMSl4Jkk97oM9wJqVq0pWOR/EyM0bfgKUiet9
tvObv5HqbEbnwi354GnWixR/0FYZSuYoYAsWPsEAYOgIdcjswv00lXqYag1f6MbL5q9y5OHzI6sx
0eixxO0oCFfxr2sv+0c6JiAf/neldaqnyT+2xsTlnZzKV04W6wOCXnG05+4GP6PrH7YFSlVcD9kO
mU2sr1dnNtM8Cq6r84rX42fnRXUpqakaYgESmNxIHlzUlP7YlsROYA7GHbAZIcWB2pRO//XH+kq9
x2VrlAbPPmpBlg+0lXg7L3oJQk/f4Ich/Fw/oft6/8IDjenfFpiBbZBC1KPx3nIHOG3P5a/zd+ib
7mCeHyn8BkVADfl07RY1btDJ2s7aouNy0nZ0HsJR/n1Wrhojx5QCM+Z2CH7mlw3Sh7N6wjQDIICg
YAoFuHnhjQreOPZR93f4sdCFex6gRh5efG5LI6ilM6tNLYHa+aM1gIKaihQcRi9hD8PPNa2RmVcV
jLILm054Vau9P1Jm2oEPqEO3D2V3E65yANbY9vAi2SYYsol+dEupLpobOEtWXMHTEYl8nlSQu0jy
lO4HM26XBfL2MbqSJVj9KACD+1nK8qgQpcP3XBXqXEM3yXxJahmgsojjqnxz0vDRagUQIQAr0U8Y
bGIDxshqjrko3YEiB7qlE1idHq7fAP7gxeTKT/bL6PYyGjGLchOM8Vlsi7VpGYQbcBzsBtRzTZ37
4P9lsW2bn255NZBi2j4YvtakREZDiJ0Y7Mr+bffOL/Uf33R1Eo0Z7lPK2Kr/bO8ZIJ3O/M66HdAj
D2XmU7h4u7AIoeyvmkVgUFLryxVTHd50DgOmoMR+l4h5tq0XymjwIsO3HeYiJVtYtaF8LRPhHvm7
oMGNZz9aYyEaCT8Mec3ACDrM3fLrbEF2RlM7oyifUNkgh70vg4RdZWKzC018DbkAGlPUzV/uQaQj
c646Cxluvxn8iwv1iAikxqYGcWL48cm1zOFAPQ/lTsbV/mGtTy5+ZVgSBVwPtdUhJWgqwiQl4WeT
jUmlALK134MWMIyrZK94U4L5DWIXjJ2k9a5UR5YYPMvsstbPB2efBDlwNlCJv1oBAQBDU7a0RAGR
lOWjfnU74/mHYpaaklqhJvmHZZhymYlFuUPAmdTgusvTAYW2gSpVWTzIhFclUJxZMqClg+LnSAPt
/sNUT8w2UpyeIBcBhLCcubYzFI3TjMeVdLfAmto0/pY87zWlnKxn0TF+oV8Kr8AARcWOLkTaZOHh
koQvtqY+6EXxqLUxYmVjR1uH01CB5vsXJB78Ktv9/2y1UZBZGYfQoLPFXqxEqlxp6NuKxQ8fJWVh
0LayIlLlwoIQ/J4377Oj5GDw4Gk171XE3ujIF+ZKW/YaFBuz4wJNs9Um6vab2xlh3dS1MUYxECJj
5O3NaxzhOYWnlbl+EXLnGuKuhfsQTZ5Sd8iCSQTgSF+7R8aicxFsitXNi2YP1Zfuz6agrEZxXUQ5
2Inr2MlrGAl561Vj97hPpgA+tpCRn/khsj7a8Hl3y2Ubf5aP3Wa1Q5oSOx34ZJKjLagpqW9zPMkv
QZFg2+Grytem9EwU7rJOo0U8P5H5h5/qKNX5fmGe98NJteBNZsmGxWUTO/py2XRl7EFvlulncx0o
ZFmshm5lUmrjlLY2dZ53Fha1NUUWa+owtuwO25Sc2ZOrvN0+6NvoUI0EITy7LcC9ct+AxmSEZZlJ
5QYIJe1fJJ4hfVPCxBU8y5JsjacNt9KNoYKZ9XhDTCfe7e3glYj530W3ozz3kmuMiavqrBsX2Zy7
CWTtarudt72FnYHOKYv/g3q/u6IHgOrbkf4q8brA9SdJMDmSAoBqmOWzoE9i3yCpjHJVVDAP1DL3
XZAwyT/ta+Io/sLKAe8rLZ6uDZDhJr9koHbluXfUsX5QBh0KWS9XJHeiQb1+oDPNug97hnvScO6W
4Aktnai2fLQFqmaPW+FlaL7jkwWa0NflmSn/FdxK4Ou3s2MNINHYSn7IF3H4YlMa5QdcFaPLnWFA
MheBcZHpdJ0Bkyv8HyQu8j0NeLmz/s19yLRbpVbOQwP0k5bvxDBz6gn9978dk/Es7QGOp3+hQOF7
9jC3Crti5N7Zh75WE26kzPXQn9eJr4gh9Isg6Cyy8SORxQZhUMu1+R8euFfAZ3tGCDVKuqZ51hGH
kg2sFjPSQJMlSZ/nkAy6W673XAdwRY6zmVtut6YmIjHAfX0FM9xQe8bagp4qJlumpn/0BG1T7MLB
lpbL3IZePbonfoAFA2mJfmoD2tLZO1w8E/CRMFNZ9KSN+5w0GbxkSiCRThMhnAIxU/Lfqlcd9VOX
kbTWgJ1zksB3ObHV+f8HoL0ffLKljRNNt51zloPAfj1bzHjpm7jf0i5jk1ouHpbq4WnLZSOGRh92
2RmprSq7QwGyFEwVfAFp+EGwaGVAXfriOYG8jIOfVf2Qvd1WzTqRg/Zoz+D8osTSts/+6RF5C5ed
PqQ92y6dSfsgCKQ6r+s7maz3FZTZ9yU5Ev4fjKueLDTOJ/67uxvZ/sBKrpcRoEGCuldsps4gxYer
mL2ehKayVnq6E6Clb1CXZalxaKDvfVyPMsopeiwarkjuqrhsdf6jHFAigpoeYiswPlY//Noztfpq
Dk90mYfXaRmZm2D6DNCcVArDvv0Hlz+JY//rkKXyftDcC5IeJjsFue47LMu4+1LadMqaT5ohaZOR
zQnoN2UFmgwvSKf15T9Aa0/lV7/HrWgfoUmX5WLUbUmtCXMeYA2xe5ct2AVxSDZrI1PZHZ2KUkVM
crwXM9CxVNSwffHYwLU63whcHi+BBlR/OqOR5LKcSY90vf6QEp1V6RXXx+0BEs4NuaZjamSjn/kp
T+4QGPFj5iD1kdqouze63Y87kIJFWo5mZ9gMaAUjcZaO8PQHvvDiNgqjhPdo26ZJuiuRov2wVS7u
iUIDkU3qgrbbw8kyqT3xx3MJcCWslynkd/TEh6GnBfFR4KVZEN1Cwe5lQsN0aC+TFsh5Yg5RBvJZ
gjxB4weIxLs3QqCBY0KhtfpZ4UXvfj4ZQe54VoXz4Zbe3Cc/vVmX89HUKRswwiaRsfVes7BJtCcA
QJaYXrTomEMcnYyWKv5ahA2dNGtwMyv6NRJcXClkADY90DYUnfNznDYjE/UB48me5VNH5w2FmwR9
BHTWX5b1natauGMsralupmrDqVbeLavNe95f97jYmhZzJdEU9FAbY95KAmKqN+3aInKbFlyObe09
tRzpnE0nakdI+BKGOH2aeNcC1kunXmH6nyfAlUCWXmkwRdFnfOcybH5ZwuqOR8uo2PjvHnyaJDi7
IKW/piBHVor3ZxczKg/FqCxKvd8IUGM+MgE06MgIKPs9YHyXeewNQAf9RiW5UDTJuohWNaEqCkPc
ZEYpFNzkTpYAqZvR60h4HH7GLIsYvg1VB5MAvxuywYGrfkTtWr7t0sAlWGzY3LjZZcBe5xWAI18T
oHITqT7aziQgT02JZuy7cqaMoNMzupBYX68/29nvriz3d8rt9Pv/bYJB/U8+6ik66vYF+R4scybP
gm30z4JLB/Dc0kHWVKiTq0XSvTcRLE/KD0Twd2zxEeOTusYFHrFWdkPxpXqJZv4B78F+zyZ0dN7s
2sjSh98SPr6+zIgGb/BA9U8XHg62ZVpoabcnoej9m7R1vnzV9dDfZHpUoTIIqCg8cmA94fU4BXCo
S/GCj+iSI7uInL4SkcfIQ1EWs24QSY8lHgfPz6taeGbYHBzOClZCOh1M1D103W3WdvPXlY8vSxDI
778aIMzhTmfTCDtFMfLIRT4OHvIwg7JSwGwrlJrJtOBVzX9qCiNWpGErrGT81jnFrPD2QriC2NjY
rIe7Fk9WYZO4e3nLhHzNBCMTPwUW75TWG8oZkZQCt4DWSYp/Kce++vk3Z/2+KhYtoNlh5+NhNpUn
nfyeJ8BnMp8e2y5Qo3AAbo/PBQ1yqItEjnsUAMHcps18HxFCCAoeQ17bwAbRST9i6h7zD4L/Afu+
cv+tY+/fywDw82fBEfr0jRgRJ7Ky0PHXm2RUvANR561NIYKE1H+TBBnLpQzrsfKRPFtsbV2IIXgR
mDT8156zrd7pHqdG+JJbdeZmeKbfWe+7lqOdm2rXvjSP6tNHV4PwtSvr4dbKRElSGdsaU3jHZNSE
fzS6jiS3SmZkHUumSpPA6iCrig1+z8Gjs1f3LxIP1DmPADDuV8EpeAoy05JYun8DVZPT3lJPRDyw
9b/Lv7MxFQwqZ0yedqyvznWGDoTFfJadEW717YvuG6ktd1+zk3K5l778VeRUnHXj01AZC5NOZNWx
2mV4xBTqODI7P7tDz13McwjtsQiACCaTKVNpzV6RGzbDFhaS3mo1xx8k7AOJmDnjGwFh68JEWboJ
f3adHNqGsGewYICDm9JnLr8HGL+FeLn/ZzmVuNvDXvPDr0LRmgmD9XQuNRJEnuWXKiia8y7qs6i6
growzZ9lUiJGTeoDtcXkD3+xnCCfODzk71doXF98mTlA9i1rrcz+3F0rZUXxA7Yu3WUDSq3qnnmg
z12hNpGEhTtWm4e0KyclF81kCD/KVfWdtQzI/mxmxf+wmwfTl+xqu9pR6E8bzG0iuqLAR2j5CHt2
rSkwa9bBewMR8NkhXG/RdZ3a68ERtBER8uGjs6dqzpJDz7hA82C+Tk0FuJNGWfw1cBM2WowzrFt+
JmXZE1M2r8kFdKiqVSYRAmwT+UhtjNXsM8IOeJGUjPK5nEXbfOXWtTN8C/Fy0HI9fhmTioh5n0sz
pfvmjJesz2kH41ZE0fdbyn3Pe2VzGiWfBJQTnh0vs6bcGKQCTRA6lfsqMJ/TP/GiqBOEo5vI6SIu
qHURCJe1CYi7fPJtuzvNjNrnGUkJrsBljYsQIdlhCFgZgduqyTnSdOK1wxtyDAj54T4OGwwFv+XZ
j+PH5TocuEouB6OS/QygshCKM1a1Laxo1RcWrW+O0Q725h6Vt+a892un6F3rysP0H9BrCkdpdn63
TepVbrT3fLy3iuJ4hWP54jy9u1cXTDYaB+J50KJE6xejj2Eno+nWACqknzc7otZNg9gFmfY18KBU
05wSg+8eMXnAJQS7uHmQXjDne/Z//rxhStlafjTYb11CiE5I+e+/Q0D7OCgxU70aoV8ffh583j9G
07pgWuv/1gmhqQft7dA6sM8nWqGtBs2+SpZBd1KBHF8fPW0Ln9pJHBNIBmnHM9mCEtGZ4EY0V/jS
s71Ouyj1sZ0MbsBpKRjCeDaz6nJSL6PaKUWhsd8VQ1NumxenAXU4Zm9hniwycGWtaVkF8+dEtHiG
l7aCzHua0OdXsQ0A8I0R2xhNQKINOPJGGA3c/s7lhoFCyHr/amBQdz0wrzPk9Ed7ptAcN3c1k53i
NYq6dTrtT4ipJQjqfgv5G0rYjeG//IzwDTDOnxhFsXOZ6OgeagnjZCeApOtLlpQStlNdLZgd9aqf
j8PjTABbYRSlXNGW2ACzztKkeA+UqCMKzG7DRZAt71/q+5hAWd5mJkk27TTO1Q14PZ/VKuedeTvM
wR9YULglmApI72ANbUFPNozQQqbD7jsSGVdNkDct2QhKaJkiFR2o4qNqzNeDHdVOZjTcJFUixg7a
0jVVdV4e/KDiKWx+JYV6v0NsYx7zDdRrDfAIlzpEFLCTRVNk6Lxx6CS1msmAJTtlMYnrig4PfAYJ
hXIzPWzYDj8w7qNdyLA0HCSHOwgnM/n3ZvY2biK60sZIdvkZCfl/NVYgfFWujDEOBJWLDGn8/V+X
fvipZ4+1GqqosXkRG8byB8QNp/Ea9ZJm8uf80a/gUUdCzuTDiIRsDRW0SXGgC9p2IxaqzINpF/Tt
Xaw7J58QJvRXvOlW19Y+J3vqyBjy6ShAS3NiHpZYGLkvckrcUeKueabxjgoPE+htHjaEy3MtNCWc
ed3vczaQunofDF/7XeCbOOEWZVfNWnrkMGQmgKCylrS3ydZjs5PqMG3F+/vgYw04Ax7/bCuDRrbl
9sJcvIPbVWaKcTkxILr/A5rQnZL+GCdHcngaKJ0IyTlVY44WB96AgHOqHcuoAPhUzRPpTLxovr8W
5YTm4kG3zWi5J1U+wyALq7dZG75FGV9jl5G8IcYrpRXXSfmrPQb38W4OX708EOkMmIaV2j6AsdGH
PcvvvQM5tfvKHTZOZDfXrfZVnrzhx7bKBfY8m7wvxiAuKyOKOz0jeS58NkEHRGXxVZMzOYMxAakp
YIAbCCTX73Df0rMHqnkidrAWf69qsW4znrXtpGgQNv7GBPqoz+3mnvHP3YJW0QwMY45kEwItaREe
mOFwt79pVAMGhSMGT08p4Bsi9JFLxu7MgK5112dT72aOkqL+PLPTbPOwKLoECNQgOajpgbYiyX4L
aT8JKEFkyxJbi2GmfDvflcyXTAG2uHfaAN7W2GE7zpTifwB147c4kvXo0FpeEpOP8R8+DaZD+Obk
QVYhVQdsGiQX0ltmYmUeRpzG6kX4Uz+4jTn4UWk5F82uhIHy804GNZjnskoy95i9Z9VeAfYpHEJg
bKL7l9yZaQoUaA4XO1P8d/P/Tf/+yOWcN5laYEzeN+509zH3BxAcTziUydDC+9z9L2rgg1hR2pgS
qM8T3dXVunQYi5PvLOky7XyNFf0e8dqxN4IeFeVrdeAPZbG9Ut2dc+lL5NdTQEcg7D0xRP8P+Sqp
GAEapGfNwp4SyWpyzp6lTX8gYP+lY1rIH8BolEDnSMCVNrf6wvMx88g4nAf2ji+gexE1xk7STLvw
8j7pgqMaFHyXVKAaCpgnp/uqGiQG2gznGe1nVKJAlxJw5g8IRXxqXpH/UtYBnZbcYh6TglEHSapw
Lvd0KL6GOL4In80ZRT9ksPWw2E2FuSnqpUUVGkL9Yj4tAnluxaJ6wA4MzjqUANXWXzpgPQnVcOv+
Fbe2f1H6KVoOm1SN2lHBKZmo7W/xhJEk/pludj+vPUZ3S0mdopmUhcgDNtb4wGc7ktS+BLokFi19
s9qK4gbMEuKzVMeDGNaTkdRka/qUDFF5YQsU0DRdRQucqEsk3B+/zi0bTGM5YMz42H301vysnIrs
zWn2vGxvoxr8/PvVFfGSqlW78/BmmT2Za3+UqQncRrrdkGxzXWnmNCNkXgyLNl8YaB/DO5xNXNiY
rg/wsRhUwWX/++Vwv7JU/mqCiFTmcw9Za2i1OT2l+KC/I6wxTh4Ozikj966uMUd9nuTZQUU8Duao
Gu8hGgyuAYPOZsYb3M73VwMy0LVmq/h3e/DfdPeYlzVnItFeHYB4O+vmU1jp9E6ytn3ECzBBwYin
v1SnrBg23WeIkatIwiLtxdicOvEEliKe3GAJKiDyF/uCFYAZDOr+BpQZK7/1gJ8MdoW2LnXPHZBE
Lw4zsybMO0z5cUsDPfPVo1r0gjvjD87/1vyxWaYZj9WkXi5UkYnEyIDFalOoIvVx94IkJ/qyDRyg
u0bkCpz/sO+a1B+tRLL75P21VrgGoj+wC1F/WDFoELLXcwDmEOBGIZzIqepkVo12dD9G4rRC9MDG
xXrJoVdHYWPXvrAhhxhw83cDO1UZMiIMXiQ34DcSv7hPzwXzhYYb8E92OrT3EjkosHB4z9Qz4U/m
YhUxqQWepBlVf9YrjHcFhePoeEsBoTSOkeYqGu2jxHo+BoekfXqj6emEaYwNcD0a0MI+/w3aBjtf
XyBftxXDfurEdvmS9Y4KvV1wlBfhoJcEzPM5FlAsRxGW4TpctQO16Oo3PA4fBWleZyktHnOprjGw
JbJs4fsiIBQ95dZBjSauTItk+vy7lurrjGBqC9PKFBNh6KdqWadNdU/Ir2V6Sxs3cA4j1eDWUUNO
cG+l4yoj62z2Rjn8i8VR6SDWu8e4nCkHuIODEjLx7zmcLSDqahLJdPlIySc/VQZGorNhp1EoG7tE
iiFNi7bGb5vVNHbnfCHsbFt7Z5KOZ+71awrGjggFTigY21q+2auNx8ywcELckDyITZ9GDvNGHL37
iFHVzlEdqRaXcOCB9QTVs/xOrfpVG1Cxi6P9Mn+mY2qopN3kZqM5MMeiP166awC7L2CPGhvCm8Gi
18PiI+BGK8YMohSwgHv2/J0ibIBKqNvZy521JT7WvrT1Dp4gXCRtZSmNBEiv75YQtLoDoAk0FQUE
BmYOhL4e80qVPE+xkXwg8qmY5uGwjFGyTiKRMX4vdOCdjKZQahfQ23dbJ3suHSSpH4fKXiLqQRkW
V5Y6YfL3Vp4v4+s3ew3oGk1QxHO2U1lQ3W7lcEuwdIlPzA6/LpUVWxi/LFCMDkzebpTan7vlXypa
anwqLY/M4ezf2Mkv9uxDONtVwpwo/gRGVZHc2BCYFxgLCz4JSTCe6BZMvkXgxkIEeuXm12cscGpX
O1aTrpc7RfWeCJuUWTKlQ2dDJlEzUKBfpUNnAjKbCgcHkp+r1gkGhoJwvtdJnDbHNKn8wvLBB4/O
xaGb9SK9KQCzHHeB6H7znTStMyNyTMMppmeYdRSfW+3Y7IGNCelp66y2VnQodtAYOxeJBN0+qdtH
J74hmt6mN4eIlv6Fl9E/lYSjlEaUT1pLKfMTIeLK2Q2IebZYBlkF9SQwB3QsMq3RbwUIe9pC3f8f
4SOASaAy/+gp+izW8gWrV8yPDdbEBCAwdWkXs2MJtOHce8A+Frjp27p5orquJayvEV7Qc5D4YKVK
RMsiuEH56yWTkLt0rEFbOwy8siAwF6YrvnMmMUqYHKvB6cinIRJFVJO65nEaquln/jSfuzNJYezs
sNiCs7/Ik/0lHMve5N7sp/TZ/XpLyQ1VOiqWzGIMQmwfPD8MiBqPhwQdQBg3d6R+RYD6rxXVGBFd
q2U5iJQ9aoSVn4xitc0LgYs/1JjvBN/mPkFW9CMcJDmJOpU/q+Ybk+HvtPEQJz4Vf3YXuZqIKblk
+oiuL5OcP/7x0p+jTumedKRUg9pEVO8Vg5Dt+8gHB8qyo9I1FbriiOXQHqW9XNDwwHm57aoL+k+V
gi6/Dncird1Ebp0HfGtmCGHYtcauXWL64nHJjHVVeRdlB+vRS2S/uW2/Sm/b2k78GtSx8jmNth5a
cHoiigN6SUDcGSajreZXnJgkUcgGMkCCk1iMHJyKDP5Eq114tRQCQAKXvfb7q0Qf/12oF6GyiJ5T
+Ah+mrfcii0eJn3VYtJlk3YFxYgr0QBtgEcLOHT0KEEdQo/JGFIuHYt7AcrrZD3rRqefEVV5Zit4
jaY+m5lu3VO1otvJNxL8ElBhezjptITJ4fl/dydsn+I5SMXka+TQLS4Aoo+rkPUtttDtHXloDbw+
5Qnm0HiAyfiRy+JEkw3QQXOA2/EaLosWtQzdDEBTZwWZqOuo++T21CYf71uSMyefqzpP/YrprZW/
kvX1m0/twjC0gaZ/r1v/oyIO2Zxf51pBtpktUEKHB2KY7gTqb1kZXh8ZqrIF3eymHPxbC3Xzogff
aJ6Vv32aLUZ2hh79DfyDhlW2b1gnqjFzMcTl7K26wif6hTtpK9xf969x2dQGTCxysAOk467HkGm6
j2wKPMcAbt3+rPmN29w8A5WlC2toDXp8HW3R0AIuobpU3byqHqYFzXHRsWq12grQL3Rt8klvOpFK
+UorhJOefPNItanOBK75pRKC7OEYsBMnuPmnki3ZPqIKMiJ8bZEEM1/ROvmPX4faWkdMLXzS+eET
cpl/RWRq2uu8hpz5knpQkUx2vDTkzPviSynIPtUUwbcdReSm9BshL7pYLTJfxrkpZP2c+4+ooFJx
LUp2Hx7dL/kfaPZeXe5WPymft1LQhtmHw0a8tfdey0eE3d+At0uObq80xCKxGc8J/xoznCs7utYo
ha7JMOP28Vv4GlVeQJOgxhjqgDHnfsiLqHMPkXilMogF2ddUFsQ5iF+wlrn2mfNHUIJyF3gA/Tc/
/kY2UBnarq79tnC1JQVDODVIQvLWL90pS7picvt2NZTfQWx0zLWG6aQ2tE8IIR4Oi1mjFZlvfHcZ
5rrc/q43l/rNdcxaBtjW7iVx59xDySy+/z2m7Kc2Um9E5mOzHUqz4sTeRCUkEztecnoWuOJFFUmC
4Df+DSLxdW+ANLwamGwwm3qa8tkNywbrww44xBzZERFe9144CN62MZTvaxYhtFB5tF3qXfEcVYoC
ccf7qwnSV23+bWI3ZIxTH3IIreEdCgK1v0l8Z8H+qR3HjTiPbeK4N5Uw6N64UPPA43HZEKnm1iz+
QWFSpIm0fTPl7f9Ye9RfzBDXiYruJSRtrL325Jb1/C/HZmoT/aC61rLUuGlmXmohxgXKDggg7OOr
v02TDVXjR05vhoDw3ysvY2jHrqFuhoRqS6jejxUOEyAW+Hvl2kILTUZ9qO9jTEUWcZMV3RG4uLK2
126HN81JRBTZFxI7TChubBmNjhx0W3VzF4hDNMcql/pUet61V0k75FIjU87z/c9SQYQA8Dfuul6B
B9q8h3PfsconHlFfU3yo2QZtIj6wTIdZonyoN2gJyl7yjpC+1OK9dH3KgK9i9JoQq8XgdQ2s1ZBa
rxY8lM4SZVrupEo4MziiO6zEy2WVfPodBVo03okl7DDkwcOZVJ9sGwBMPU+BkF4+OKCUp7bUHls9
KvYKm+OQ1p6SlkKT70w3LbDFhnmFBm6oxHjIKJG2oHLT8ttEWxwIs8pGNRYAR0mjr1g/J4n5lK4F
h5V8lmumpaNgBex9gasNdQv1ldQLOwDPWRuNpkDSuLv1aJctaG4JU72lgRgUnCD6xuw2mS7xXq2f
yNFXChmkB1fet9j9X5uvJyf7Oj5qtegvWWbAuyceIwWTUj19YIr3PHLVyUBWUuui5mX1EmRgAres
G7GTPyxDU7n/Hh+KA6qX50EaOLbR6f1F8wJ9m6D4GMjDMxT4Jo35PLOg21zDErcy0e4yjR/3ou++
mX1j/hfv6Otdh1pQAEV5aByYdaXSmQG1ugGXNJzggYQLSJ6A2/JTJvZox2nRFKLJuCTbNYmtzCMB
CXH7/Ksoc2XvS/wCpqcJDkEFJYyyT1ekoNuFacNigJwE0TsIzuHz8kNjWMEO5/FUu9FodDyueg54
qWThVjIZOYsOYGMEk8OvcOv2GCNMTHSJWiPfxPK+oSlyppt47dGgai2NGDL6PJC9Qt/23sOd164F
qb3e5U8UlOf5rPO2TSzmueF/ZWksmQEN+cllOkqC4aRPDAX5qm0/hwn/Q+2uFHtLvBZEQI+L4DXZ
LaangdoUUJJNCC/EEAdEEEjDMtlAmtMPL8ST1VVx34WVqbqeS8tt5ldMOe8FSab6qN5x/9YnfIQ/
Tu008GrCo88abj55lsqMjrkO5sl3U4AU9vvuffLtrbKIwARhN6QNYfo6Dkd1yZrWD65VSR+r1tnv
J32dXJkNkZRGlhNkCF0vVMb62qvcAjQD/HsrTE+caFkeBlqfQKDU1ySJulnMrbead6rnzhHJSicE
wD6MCZOUFSIvPy1VO3Kov0QBUbWiLai23jP2DCcQimO5wfLFuNhVtRAYwWlVXRzDkGBUwfuOX6xS
NwtjFujHm8/UokJx0cUxYskC2QGYELC9Fa84XwSbhT30DBQiX6eE1L3oZ0aGIyOx/1MwnUaONyBD
LTY55xstvLzWjG1tW82Hdm05hVauSRUxhiJQ8n8jytXhVZGsnKXPYjZ/JRHT1/wgwwumGlZZZACh
UlKwMrn2KSNBokWh3+6nwMDTzyX/Lgo/tCc3JKa1L326HiecBC+UoXvcLsLUhleSfdcIMv0OuT3w
8ginqijTESNJZ9m1snn9UKYfjyuyASI+EUk1xAnQcy0hSFP5XZMWrx1ocIpE6SJ21ZEhmPdktAYh
SqfpqhxR4vQEH8odzXU91o/DEVJa/QyA8nyzvy/XR8NC+t8XQYJYXb2JbxIq4SGUSNvbu2/zdmNG
XV9x3nX2CgdiXPBa6WNKNcEyCZeGxlIBp+qr9yghTEMbbkyPdhzAReMPU8xnuuvr6gyDvPu3Mycr
OgU3LwBYsNZrjk93SvWh0wr1qWgja6IV7/Wx7lVGdP1ulK2+P7J4zr3Qx9bxfIWPswBJD/4xq60c
8D2pCq3ekb4lCV6GeYoyCHCuBu7KJ/0B/3B6ZbefktAFR61zhTa8SFhcRTa6YyWkWacBKX2qjGnX
KR0HRKk/xcu314eq4bxV8gZYEtns28CFzU3qtZn/lXnROpz2ftvwzghrhNUyr1cWCTtGxwr/nJCW
RIBumshQ5wC8ZQPIGmRA6em/FNKPL/RLI5spMENiL1GzrqFF6xor0E3PsSk/Jpbj9eteKPVFeU8h
tIubAo40Gt+33pLSz7NVGK766NKmkxEilMNkV69NGqf6v56bKbm22WBwsTtNs80RxSMAkAWrU+gO
bL3XjoFnaL5m12kuUgB5DnNIg1K+KhklYet6+31P7AtowqC1H0Aij7caJgObyPywzyQpAb6M13/l
ggCal7ySd4BsmkF+WzrGeu8DDnb5SdOFXnrNVTtXj3JQQU5ZeS84ibTaOHqs08R/D7lnUQeTF1Ni
TyRGITRmy9Ya1/tPNFtjqMaWBnhsujnKC4k6kSWY31/WwN8pRqvGFvf3AHfshY9uEXWaFpm5BNcB
Pajbp9eOphVnPMp/J237P5pMgysVFUENdoCp3HkOh0S5EyrlIhTJ/2s9jAohwUjzJzSbCwl9KNdg
eRWmGhEtLeI669ZFM585ZhtQ7mCYtRbv1Y+vhasX264jxyNTh1HSNCuJevN0q4zRoT+DgTfzzAqa
w6hezSqC6kl5UMBXCQGoFMMIOREa/kA7KWJo8HCKfAjdA+Lx5HquYYHBB9n+L8d0CHaHgJ68erV9
G1kAGa+PaR7wVvR4FGNwnmETM0x+Qe4COVmvOY7rDRWdz40JH496QnJNtxzLFcWdixdTLodGm1Rx
4YMOGFWW2qsiuNjIXVnOyYK5zsBfLW1HiLxARuOKrTE/P+LBowXg5flXKUOlpJDL8gtq0wTA1qM6
/sNAk8826NSlVQgz5mT7XflCnVf31HiGsbZBVfcmkxhyriGzvEGB9pktuagHaNgl25z/0+uH8ueY
tZFlENvOU2ctKht88LgEjQHJ3AVCmX/BfqjvOZ9rKu0AEldxPZpBgHFzZyKE/LNBPnN4Hr4r+HRu
klxj2Pl3vsl2ayrmaKWpOUYoHqLgEwVVJoo+tgYwb98oypynq9x9PBQkbhcZfwggz/w5tCiY7TCP
C7gnP7b2qyHPpecsZxJQj81fjSWPb8a+hlRBp6cXBm8o9eALx6zxIHytGpz+9dHYnghnokvc556v
yUWeWi4OS0qsP8r2AMznNbv7h9KlusNMRVjrT1oh9ZQqyqoHedVTW0wFLDT5LlY7KGu+mkoF11Ke
VRhxFp/F6T1cydEuRjZHA3vH1JiWmT8xb5EjMxwdgUW3x2I29tMuyhgMNk+898SrErQCbnU0QHL4
lcJe+Xs0ROjviTY8RoDROhgp/BXkBHi4MtWY7waMBMTxHjD9KMtvGqu5uq5Q96w8la3Z9MPm1xU4
yjVLupTzynXMiejzHXbp8zD06Sr7Bb0T8gOY/0utSdF9mYmW7d+/rtXcJ4RhwyLXesQjeYrbsD8i
Btf7vrnhOTYFiA+eOiDgI2p2ZvUemIhrC7Muj/bOJFHH+KF2lX7FK7UKjtvHgNzPmceUmDy7a0tA
Dh1uP62DmYv8vBIAy6eIdnZPc5xJcUZFfIOwt0jQ5UhHUrKMPnWfUCA77quhb6iAh8xderFE5qzF
5WdY3FxE+IgXl99nh1TeDaqVe3D7XFEzV+p4KNsps+TGPqyTSEYnYqsmtZr5RCH8InnKIpZM0ZeQ
b/s1obbEFafhpMwuU5CoTq85Oc24ubtKJuhilifoYsv7AzvEc+rjBpF55tM5wEmbM19Zu7EFsQ1w
/l3u6+ztn0CBrwA5ZM4eD3jfmRPPnJ1kaFb6WI7Q2wFX4eI1rVyQNHwqdI0l3JQr5DBxBTRkm5Tk
1pUvJ68/ZhCut+1gpCC06UlKKC9Oc+AZptqzJevBYZkG7NOXto6F2EY4P161+SGmi8WIu16dBnER
jTQGBoeFIaU5FnTstDk696Z7ILFWSPgiCowmSHaAxThHcYclJhPD+JNNNCrm94IwMhJ2FRUGcSMv
KKxIPxZ/Nz+Asd70m4D2D1JKo3fBNyWL+NTIFCVUtJQYAf8irCjt5J5FR61zngT5saQ+ZS42cPP6
XuY0ume6MnKxYkoCKfhC72+wV9419E2sdePovXPBFOkLTrNqOQzUzR1UHsSmCd0WF/+SLhcaDR+n
bxopW/Ya4amZcLw05V7xTxMDy7gaHCTz7PcivnpUIhe4rPASlNKqAZQGvQdePkt7BoIX2rk9uMgM
J5pgH1kiFLjKRYaL4+0zW19ChUxwxpykVpF8wDgVuG2uyV94/RwnEP9hI6jHxM2e1GaAF429+7TK
5yaJv0hZM4ywiTqoFueoobmV90EHM2TZZTUjBHREJXO41uL919nYUVPj6VOlc1bX2pFK0pETJ1/7
txyBY7yPq6dB9mSYsr2e15BBbldiDZ+7dP9qmn540b3r+RxbwYAO2MeRE0fUFbo/qZo1G0pUWbDK
Ni1+0Fo1WpGaL0W5pfS7Upx0JU6LOky43/S7AvvhGJrnhqRtAKTwG9eOmgj6a1cQiWfSVx02nFWa
Nyp4r+oHGFKzZJ13VOlfpAWV+rEFInX2sNmzt6+IS/BB6R/jZcrL7WJOwLM5WdfuBiMZk0s1SUBM
CJuvzVlqxEAGdCJcuo7aev+SHNyXQPL/11ArlN0FsS2qgZULa5267r6xuZFlLyBfn3ZkgvUcA3er
19ViQaCDP4U+ep5+/gCtgSc8GglzuJqy95DjKhtK+mHECvH/6JWbrwA0XrJ4xVjx/teAp66Z/CW8
jxNZ0XJDb2tNhJ8uFrGh7vO92Z6lcdFEuToOhZGqbYf8x8fcvuC/Mx2abu7nRiOzPrK99L01gAU2
Jr+IGqBOvkh/6DwTCIz7aNCedfBstp1YhXyx4DLL73y6xa7v8fDRRq+RuZLivF36mfufEwYlsre/
U8L5b9kmeY2hzWWEUwxmKTLiRyGUT7DFI021kXrolJ6jo3YPCVkI9hGviHj7pf+OS272Hc0mUplJ
vFIVHY4G/A0wKQNbsk+I0wbYXzu3aYkGSzXYH8mUQ7Jl444zEGo1aQ2P3WmwrbcpHaQjr7Q5sqPh
y2qvf35Rm12HkZGsvm70La4losnCcpiUdIqFbC3ejfJvZwYNSt+aC6hNhWZ35C5DPYDAKCTFtgwM
OIV3ghMAdP2btBbN0TVIP14KPsLhvB2HYAk0LTefpexlZbJ/CXvNErMgtAJ+m94BYPelgU7b88Mp
i/R+NR71NHMtnW8VOrjAkeYjmM1uHD6o7Bn8hV7zZoNFn0FTDWxUfbR51HSs6DM0vAYNR4OhVmIm
/mIMxE/+6MfzEByB7dH0AQxQ/s9bDj1wWUGdes40MasHXFBYvuPuwxWW4B+lsYTKeYX2v3nE1L7n
lQ2FDLtcgiEdRlWvT065IGb8s7QZD+3qJAK3A3QXgdGy7XUM3eAmdhyZJnxG8deK/vjSwGz6voPK
b5fDqE3BoS7a+PhjbpGoggiyhXBMwQCZJWz9baFgL4yBX5PZkhgwHlrv0OU0PlZkoPJa/M8fa0Pg
I8OdgirI99Mq47ti1/OxYI3WH6xg892ci2uI1JK8rkxZC2eXaW81yIFb4O6ZGsIX1wAZeeBW6zqQ
UZi3+zxQZ/169CR90wx0FDgygQaNhN2VBF9KKSTfZAFGwMR0LSX07ca1ZcVl1c1I5kMWoIAqOUsQ
M4jwU2azZBfOpQnL8TgTQ2KKhUQvb/4FCkw5LJ0X+x6dWfh6laPoQjpenShqf1kC/GuNbRfImi8I
NRsntqBf1xIywIGT8D+fWItdYQAtqp1ipk09oBKtDNMzXxccs7ACUIQ/WyPvFUMGlVl5WMXR/B2o
rk9qjBchguUOuLw6KTgZ2UC0i7Jm779sICBf47RuKWc/Iv6NLC4wfAcfmYu2Uf2fNZLWzTQwN0Vi
cIeyNRDJQz7nZ12QBuMJ51pNNrIs1IxafHWe+885TjJjn5pT/E68tuNaODmctOnC/aC5LIM0e7Yc
FcUAElIeeLTjEztxg5UywHJJVSwp3RAUwHiUk8CJFl4EOJcFbbf9h5MkN9jBcWN9EKla/gON5oFG
Af7ObArhy5gjaHlaoMRzdoiY9ORebm8z4olFRYCo6m4pCrp3gC8l0illChznPMbkzeC3hbei+Xqc
/idMqkOOwhCvDVhIjVzEFZ/s6dyoGDOF8A0uHeZMmtzyC3dnjPf81okoMQofAdQH9dqqNAR9ZuGE
hpSIfPYm4rJ4cHS+vq8JYTTimDfIPIdgV2xT0ghH7tOg10W7IRIyLlZe2X2T9qmnex3ozaQWYyqy
LVrpGiMh0Gb7dcJHFBPE6IwgGsFTQK8xBv7a0UMGFeygnxas0xhKG3AlDJc1SEutuoQ/bWGkUtPi
CQepNZDAWUcxb+w9tuY42G18MSUlNHNpwNPQnd543tL1COI9oEPVYewctgtBqLCCrCxODVNFOi05
sv0v4nS4UesqZLh0KxyKHis7sOtXXUFiiaPFzbW6LJ3oCoeFl2n25tcMsncRyH+BNLnsvnuwugfV
k+ttvoKj/oIwVLNxoU+FfAv58Fs0ZUx1hfQcjg40GWfuI6Rs61kKnkoG0UEG7/sT1KPcd5DUOQqo
SoMNrc5d5KbBRZ/L416KeYq7kxITh4/hfbOx5Ov7UltAVJnB1pu8szIQyrmNjE6pZjXiU7yQHsD2
0W1vtI+Ebe5vPTAFzrf7PtQup4XFgcOS0qfvL37BGCFyS/+RTyFbpKq5AbIZ4nngWwdZjXxoE3GS
RhvRELRfCqmdQsVUJ8vRQs4ViMkMsgXIuRpl/IqgpmzZ/FIerNRO6CV+8TbmaGMGXeoGE4OKqomW
r7Q9iYYQsvmPXUJ2P73t8hdgD3n3+0zN60PY3Tsh/nQ+UdIVC+hhlhzwTvL5pv0h9Q2c2dbGvLNO
A2LWegwcG9O3KKv5A147e1O8qyWeEyRL877Qaf5WUIVNzg2LspJB+76b5VD3ESrVhrBaFSxssR/L
fdk1qCo3XsAIekdxs3EOBatl1ciLHFu0M35+6F3p2u+t8F48Y4ademtE2+g6l6DxyaGQ2DWTrAZO
CSA7InzkEuuef2B/dgx4I88I22i5WqXkheeGXmWy+4RepfxbxKR3GqT0vc6EY/qSO5vkoNlez2Ey
LmmhUvIKtqhC2rXnPtfFskZvhkAd75oC/rXM4+JZJr+brKVJUzhkoqN90iMSEimcw7DrM15cI5KN
l/aHctMmuxyqgm1+Z0bSXcgNQ7IVTXoxc8CQWlKndm04Y0etJyiZcMPTFBCurdD1DGlk/3Aw041z
sbIQXWNfPL3vROIQig6wkpJGF8kSx2cfxtPRFAwl9PGkRvQ5iT9i1J0FJoZgXt/cRIrUH48OFIUU
oy9pHZceKTbMYJCVTjGAFA1Agvz4N+WySxJmzuHG+R8XOV/dJXQTJw6jYPBa4kREPR4CTQizxY1P
nxSOIruvow9dxbLQ8aHr3QpN5/r8W5jF5HkUSg0T1lS8VAinnB8asU4CCcFRZV/UPZjqp+ARSeYT
zcSPm4HN4kozdSP793cnISxPyb8eywcXie6vmLAhss0gTqOuVEHzMo/5nhnL/Ap9PsNO3lR8Mr3l
HakqRWrz72MAU9dVaznsGxwAv8rvpbmD6v22XRiimoUcumpJtcG2O0olzMQpix5jc3Ef7qxn9XjE
Xkgb2hQS5RrK3qhw1T8fCZRChwKNAyNRxVTLcmV6p+hKi3T9y8xpvVJUcWYezTsjZAJOzV6Ooc5G
HKbKD69zD87epk7/j0DBo9VG/Rluhfh3F6Ky3YxwmZ8QDksQtTzExpQJG704cwaIYYtZ3WA+2EsZ
mO0HGAYljb85c1yBk8UuA/al2LY5KeUwte/2Of5irg1WkuDqfOkG21CXLWHf7utpTXTopAvr1lHB
5WDQIxhwW+AdvP0IWR0qCi5pDWouLAnuupV1Hm9DjF4AavxZuqqQfNAI+Br4TrCA+MHsydTbKTFB
WxwmYtG938kYL6JI9X5/HzOxVAPZwuMfm4wNhEBbbgdJsgMY3txlbsKq63bw4k/On1uT6ujkK3wi
ozRMTIn9vgwgAZ7oBd1o2gLhzMSrwCw8FoITALBLhGLh8fxBGAfQPgr59qysGhrMvhc9AKYYohLZ
RJbJAp0z3L/xO9+YkdH8Gnp2+SE9HNQcQhr9/e0Hus3zEpyOOVakogQCOGU8GwPLjRi2XAX3rJIB
FCs1PRPlKt2LFB3XF/1Ervjk4H5vV4ZMWQsuHCE02u12MNw7HVXMwAjLJAUmy9W7m4bu6pGKWyMs
3YqJPmkPfdUvHWJyZnSFtgC/VJjzuAucw79psKNaZ8YmhWEZ3kFY7FJV4crtA/TYIiQUFHdWPp7g
2l/Zd97vyekKKSJjexxgUGlhKlJfD2rHkdbHFvxrSg2Z++Zalmhg0oUg/fgQM5TFMXyIjx57KR5q
aXmSV36dpKkx5di96Ns96+4a5l5MF2bUteIG/Ep63GLm6PK5qMzTFmMqwp95jZGvjQwz1KAVRdmV
zEMg9lOtYWMOtuBqjnCauqT3Q9YfsLfURnZLEpmbCkxrmRT/NhquUMJ39IMm9BjrJCx6PgoetLUY
Lm0RL1uYqvC1/KjUaDMpz5fdPqgPLwUn0YnJ/S2fUMXAWSzz1VwNAp3BjelelrvhjDhPsjtMby0Y
5f5CXBvMYeM18+BWfKEDEWxmPh8JwDLlQIt2xxFkUdFlQRjwvhnnKvVqE77f3J/nS7tmEmBn2oKI
dIHIh2xMbkZS3bcMBh4UOYMUf/yn4YpcVV79AhPAlOkISImJJah0GnxUC8fYIDwSyJKUpVwoVT15
p9g7Iu6hQIDH8qsBRnyOmweVlVZ0Dlqp3R5imMBDwCYR+wbByefCKZs5WwicHOYuBiEos7L7GiXf
qkqTD/c+prYxcU8F4V5KcArDuAINjcxKbAmJ8ROaiU4zN30r1lpLNb+wnB9W+ZLtxgOwQerl9g1q
yxIsGotWVQBsdkDhBZ84DZ5/peM4zgykQy8Fp1NDVprnyLVuAlzeEREmuRLEAG3EeFQwVRH1lKY9
6Ds+VfAGpFrWGvWFhoe1vObOnZm0GXk2DxoKhBFKkaUvWnN13Zae8lgj/o0eD4P+m/ckXXqtSzo5
u9gzkgx1uvo85m6T9+KIISFBIl+K7MViIBGaEAfEHFywUbHY4zP7cKpbTJyoMeiYb/5dJUZE0h/B
Ue/jrQsFP9LLuwQaT2m5cpAgwZWA4+oP8dydLmEQJeACi3dvOIsVdyt8sKgNYe0S16jyc9LMZjnL
demKWHSUcBS8CzhUOds1RmybjJJUuHUcDVriYoP8Mj2bGFpQNbHucsPI97NZGt0rjsCruXWQbpvC
Z30sAGtBHlf50ovUmbtva9XYHpJNORQNOiT9MY1Kd+BBLuuawUayW355o+uCny+lMDP1MDvII5+0
FFIKxKFV8IZ02efV6mHO0D7ckmt4DMQUSwNrdJ2omkne+t/oJnPFcOUbeGvjMgcY+PEhTGlBf9wy
FWoO6s8wI3QfSfIbNEzaxf9ynOtfoyQDI+yHCitOP9elo6OJNJlMuOKrJwb5fgy/PHD5pmRI71vJ
NThMQk4f7dJs+ilCrOKM5h+u0ra3+UGxb415juTxReN57uUPePOYwvtqFUPdLnXVjTkW/yO/psQo
FqVK4ita4rPzlx1Hxu4u8q8H1sKXulABuyxym0g0aiviGB0hT5Hr+h+6V2xLCE0Ppi2w95d0PPZH
kBLBmVqEegQCraaXBB5DvcXBgloC4EoYnTjic3OHV8E9fPyN5UwfMgoguO60TNcrLlMGXRyayB48
m3ryZvJlzVQbBqA1oKu8qROh1XOv3iPKnHg42Mu8XxDrJ4aHHU/+arBlZsYpe3tDn9rHbdoEECrT
msBmRtV0BedD2FQXbqb3T173Y42QqOq40R+UMt3B/WJbTwXYfqao7BfU7a0Lh4cDwFxaccLX2l/y
CNlQ+aEHK0ujaNsKyM1SYTpoeYEYZGrQOARKNqAMvuxxYNTT7IuJ3kDHZ1zg84MOhht5NF8BfM6q
qrDlFiNXcmhRWKbS9HJmMSGMRt4IAJKH5ADTet1BlN+oJBVo7AWVYOhZmbVpXP+FWXkX6r6UYJ1d
Oq41FLP34dEMjrT1pSMHCW8h/uXQw8QXUOeP/5sQuVGCT4bF3KgGDnvYil80e1JJECO5RUrQ1d18
fOoPpFDBJ0qG6Uc7PzV5Qg7tPBCysudcksuqaoAGjjrS2+hqeHa2jVE2YvP2bEG1C4CQadJZ+vvV
mZG8HtR3KNideapGJJiqAnvUPLkq2PDTAJaPBCM70nsVXgUayiniqI2+h1KHn+UmbphapSBjTFQG
xs29sK5VmSZZQ5Qp6wo1whsyd1vowWxTWKRpDwYyExZmsQBm03GiD45VSsu3QA2aaLPLoAvBK94s
CgeiPdqSO/mw5wtK79WRsrruYh1Vvr9sW4CwqDbC+RTYocqd9mg6UGLzlHOcQ+srOCp96xUhxHSz
SOHquFh/fpdwrVNF41slxQXd7BB/ytq8KpfUxBu1PwZkgYZpSg3Mcs7Sj7an1Q3xkgJmQw8VU3F+
bUp5lU0s6rTuB1Uc3mtZaRjilJlUKSLwYyIUeCCcnJ1eP2wVJ8bJO3bxt7Cp2iO32ETsf8G0tftb
4BlCGPWRSjADs3YoZpc3GkZXftw4l6V2VLWsB7SbiPBS6LyYkxvH4Hf5abE7OpM3W6D+GtJZC3EM
caYhjjvzpo6d376lNpWNcKYZpWN/GCUlyfov/Se2EUADCJws/qvODzpntkwMOUxGOJ1MeAhbX4nq
XTNmjtx5+BiecWJuKefXJSA5EPwYOQtz9/2rJwf+jnmkMovdi9b4iyOz8kmH8/e3ILoI0u49UKbZ
MWJmHKRNi2FlY8j0WdoXJe9/2Yp4xdRl03aWXCBwP2hnvoGV15ul0gygI4dqshJnvJwcsFvPtSVh
o9rVqzfN82yU1VcKgQDjM20YWWVDE4kMh9bynl6+PeIjjcDwT9FbGPTK1GKRfr4QdKauZ6qZYmz1
+OJ5L9xg5rScxr5jObmH5WuHQBb3zHl/kaFWF/KSO2mgna2BmZjzTnVQEVBuLePLts7UOLj0ocuC
wCss5We3h6ARaA6YPr8S9AHJ0datw0aRR5FbpUZ8osS7lVTqm/rKJbK32DSKMV0JTPgCc/z5HFK9
1PNkHvlD51ugsOLvMUKMBivaFTbr8IgZOTrjtxlT9PVZzNy9FD7krDsZGkEVKT/r78fw6DdEKnuD
o3RstYMakOmrQqmaIt/+Lb1Y+r83NE5PNNW8lQRg2A6X543H6qi7jltmp/xVW1dBYEViOL7JuWjE
GY/76+XrLQcLFWzXd+sHlOfj2ef+QoIDwHXAZ4WapkR747H7Zbl5s9gyBZBXuZ4PH7SGL3SI3rww
hbCODiYdZ5A/bEN93LpRWw2AJVC4BfFuEpHuncMr1Ugzd7YxxsOdN1mNW0sqK0CxvGBGU69GdkCs
1VLBMIu0mq9YJkFgGzmu8hcP/pgz6prggiHesQfDfKTjJ4huvz0O4TnKsC39IMx0weYOZm8ESg6i
/l7/+9iPLWI/yPO6mH2yE6yD0e4+oOYvWgaM56/Hg2lFnyxtTJBRVDx/PHpF6tUrsvMOe6iDMyys
g3HcnDqoPVjGuo9CQZ1/a2zZbHuyTo94ga8ZGSX5qKdaQzh2lwQDOzLn7kMz00JJj3vQuEwnRCJi
EgfwSREM/+LKr9lwGK4MH5a4m35iAgmeJQAl1rT5D7fp9j1W1JmcpziBkmuzE+rC88/XZ/DDUyMN
3TCGlBhrYGjq5HD+9pBs8JuvOT6qRr/gEL9i6EBNXCzhF5YC4HbW9AFABJFobQaTJiujCfMhVJ/L
nDu2dcvCXO/QpPLlr/JD4IL8W6hp8yTBhVttmzdRVMdOVfKcvYWbiZ4QqJp25YsVpbNKklqFdzvD
p/YQetRkoTM7wZQAhHUdsqer0IXIZE5Eq6y4SecdN4EqphYYD0eFHWbcDBSCbP45Ux8NRV6bzCYZ
C37vZF8eOh58/iOy/cqz/RNy3SW4+9kx4n6gSd79lUJVwNoT9L/ud2V4d5Bm3jyAy2li+QkU2g96
EL88ORAaTDVnPDV/gl3xfx4HadvcRIoioX7kfPfd9Fuponi5OHVJij9wx9WCkuRRbHKPzYQLtHRv
jgELswZrTzDCY0HKbvu9l3uCCo6Y0mA9vcmiMvfgjHXskWi7c0DGVyjqOJrYvyAQyn6RmKJf0St+
f0Oc/rEsZbpIbZHRMX5CUVzvYfIbexSxl9p8yA7Qv9bG5ufdoXxkSUm/Z22Z1l+X11jFEFyZOs1+
FvRijEdfvLWThDuFz/fVZK+lVSCAZpsWTHw4i1ijxrMHpdMjMpwh+32UPbErMKdcvXC30ID46/C7
UDVcM5UlIZY+EpxzL24pvVl7G3U8myx0nKdXBzLU4RlOOk3aIRt/M45Ss6GMR02HSd8NEGcUR6eq
Xh5ZgkcSbTHXkMi445//d5+/5IE2XHPhANm0Y9+4UR3mpzitiEkcxnRPAL0vYWgawRa/Pb2BsViv
9g/Ai1Rbfkfmncohn732g/BdB+aJTwTsjjOJBpdVru4NeR4fdS7T8XQcXRdcwh0XJyGxohYXJLRD
2AVqifdWT36V01AVbIKHJkc82WG9XZm8wLpwgYkLPB4w4YDkGaPGPVrzQfB7ZAXccZo9Qb5rL7as
oEV6SdvgF5nH0wz2pAY2nWG8rxFYinArm5/pp7PrhjEzkFCT7gU4wnfABiwCgKwABw73HlMx1qtI
qCUg5O6vHQl4a0Nfl6BsYKjjcvs9lIboId/aA/1J2Lx6nDMAWma1dp4gxPemfR5S5RPBetP7yjlJ
GPKETBVu1QArtJGPOPDxfAR4tHRFGWYHlcU1+bVh8Pna5DaFkYDzc5mrfNqbnhnT824S016jrpow
e2irHjjwsu/oFKnlA2QZ40OAH/EYdqHg/aSJIAt+q8jgFxbRNa9GjhbevzEfE1l3qIUWQX7HFocl
6JkoZE3ZiBfn1nDvxNdXJGcTYUuYzNd9IjdcxUHJulejahh/g1wuYeV8dzIHqN7K6daPg56xf5IR
VQH3C7fNWihjNVg8v4JOLINreOQRGumWcLfkXfDpyjuImSA4Y5IkNw+SirD5922MTfYver7PxTQb
3BPG2bUcgKhUV4TVYYAWGNAxoSdfSADJ4hfJm+Pbt1iafZ+3FQcKhmtlXMbfE+8tb/t7nXn4VkUF
DYyjqpKZRDfjul5tBgiOrCzIJULfzZSh51QhpVmR/3WC/To6eXNrd634uvFYomAVn9Ob09zKKeps
M/7efP8g2pV5M7jAef+b2pCrZ6lpOtnUihiqMyQcPVqosh98HDn29Z1Jcjs48nP/t4Ga6uk79+aM
i1QOPEj2bg09vVKmKWw1SXKjRYW71MEuwXLdN8JL1lkYnozYO/R3nzTQ0y31oHwsVkDUW7ayvp/8
LJCWvdwD/UlxRJjzqhjfIx4gJZxxqnHdpzQ6gzZ5kzP+0kp0e8QbPmRNFruSWrv+QYan5tHMK2dC
7O3Hdb+cc3Qn8c+EgiZ9z8Qn8oDJKDaCXfWNV4T2J0sW0EAbBFFPqZL9vytkfnFyAcLDveJ9GQ89
00VD+k4mhmFIKlgl8wCVpw5C788vz5cNOqFqUi/iTBbhbNdx7/SKT6kjsl1lATiIGbH6/mZsSraM
t9PmhhtN3qv25uJkTn+zPqw16S5V0Igw6Sk22lr/v4sMM8eKT0KSgIJowxcEbtahymLdzoH0cHwq
SJGrcNvrm5UlurUXaRNOWlbCWAzsMPlQDgOTdlIPzE7BrFyvPh3w4od2a/ivtxqMdpmTZoNMHT3t
rD/kgnHfQZJ0tGVDI+ksI6+apOOAWCiGBXv6Xl2VE4uN1APsaHDO3k+VMg3myi3hfmY1TzBWTfD4
Rt9JeSeBAtLe8JQYGhV/xtV0veJn5eFkNll8gLmqgzxIjk1MRqs3bXnRrokoNq32LB+ORNcwWbTj
nmBngvl7uMI+WJKFi7t3TA33WgCvy5TX1q6cPQfBM0PXZu11BU5yXSTf8dFEVJcvx31B2JglItr7
oWgNs4jzR2CFCh4E5Nd8MbrCigLHdUn020giZtc3nBby44L3j7mzMadZqCyaWYoivk6SZLL1hX+J
9dvrzUeEf3pyFRn+hpeea1y40lEs1iFLGwq4g3YDK1ZM4jU9/Ip2wslXIV3RnUYHpxjev14Bj6nh
qnqunK7TXn2QqnQPYl5JP7zSaRn44O4x8imXdQT6+Zqz4zR5Rb/vZl4pPk1YuxSKFWubBb4Xd19z
qUJOwApkhhGyIm1xhUxN4O0QeOrdxu5ovDrdI5bhDsF6etlq9jWt7/4cFYucoxfEPuUTSQDbhJcu
awyYNo3wLgzDbK7CPeehUZML4K0oIWcQQtvixW326PzvtmYj+rJv+afWveLDBndeXYTqC3B3InVA
6jJpIex+POks7tpxUyQtzT5DQdXl3npWBMTND7Dn9DQWsoPAhoOSeH3Pgt/vtHF6YCLYfkAGgltW
xrEykxcPDHIm0hYGjBRtGFWvHJQYDj7fTPVE2vx+HOZSywIi/E22qFNP5jMI41XOeR2MfyIO5O/J
kVNI4HWWJJbAKkkXcHCv2ArskeXNnrS43/xzOVpETS9zLNCE2LOUup5l1rQYkfGfvUlEIio+6UQJ
sW3CjXdNvxdSGjFsRvHwkn1melXb2+CgJ+ZyLBFy1GLRjiZh4QKevbTixDOdKuCFDlo2N84ULoTm
IL01RrliLqn0JA7y5x7gMPP+t9glErpP3R/Z3g129l9431nf+T5JDmD59B1UNOYK3leuACOD+LzI
K8/BQdFv2t6ongiM5Zh66DpgTwvAAx96Xrdf6WNt8ESthQk8Y9Ff9CGFA5PlOzJSy9GJxLIXWmiZ
EOoxjojm/LvqfX595O6Oc3xMK2RGlJgn+4afBZQART5meebeiOFovll99fAIl2l9dyCG768aT4Ji
jwBx+F8UMr16JvKd3PNFGNbkMWd0ctXgcdG7Oi1njsWedV0nXIi2lELJIM3cfP/YewiGCrDwoTCX
4dKxV6idYsd1kTENBV6+Ici/6LqwOAEMRb2QdRXHlUV7VHi50i7SB4M428SmtGe6VLZ+84DXXykH
FXGA/9K/Bn9ZglVhWRc04UxT7LDKxIL9TF3vBd7T592zhvpohfuMnk4VGKyyrlgBJohNEVGh3p6p
LDSfNT737rpxbN+qRmOhU/CPfAaLGH1IQHNSNka0tW60zSoWZN4Cix/DpCejHQySIjjk3Wj9jPkr
H7Zee05OX6SBT32VRa2FH7f9+hDqJI7tqmc/1YNLzs+oP1TCoe+ZBZOgZxvdlgtfgPFsrIxpe2RV
xRd5FhsxfL8YZK5rugUl3rJVgjRET+gsx6X/VuLd5iNoVSGzy9Y6Xw786D5wZSt/Z8XJW8np7ucN
6RC8opqtWokKLIIpwASE1jQtMcFfzLTy1S/JRqK/oLuOXufc0Jh/Y/ElnTiCcV20VKm8WJqe0Vzt
KaGWH6o4Uc87i+n2Md3/4SH0dHF7WtmVX7MU/+BvAKRMLbutghJrANTuHSnE49bVbS351I9bSGPf
1FauTQFH6/ff3kN2dH4PEQFL1dzhcBqUg7ZWpnOCXY1odEGUToaGjXqV+YyIPhhGttAJOHn4561F
AEnQ7kmZQ+8g8OfRI6u9J0iEfQ1VKiajqIAScjbVKRLaHYuxwjG1JK624ctRm/tCWXLQ0NQbDHUj
RFLZchiW+WclcyPEXtTMGjQ2hFYZZeS7H6gXn7KeJqtMo3BgttqCMHXwnEglm/H/0vSUAFdNjgud
itcDCTgXspQQ/cZsszRr9nH3/5nRjq71hDX9rN3hnelr/ovznwXE1UVJfttdDXEv7OA9+e/1Y7p5
8noXoZLgzNToKrCdAc4/5j50w7i8IBkiS+tnQX7iHxloQzahzM8QqoftgFIlkmyaRM0L+P0OrPx6
adNA+/9IT18GqemLC/i1CPhtyibo/MoCvLTXznsAmbLZkmTGLg4jl4WnxPSZCpPwPcv0ZQK3jwf5
Jwar2jSUWzlb4CGwy+os7oXPuRhAVSaz1aXEFjT6Xufk0Oz06q0AeJCpGESHkLACXn37dg6jCNFx
Sxp0MocSCkR6bU03rjDobRKYgMzb8et7Rl7hsMsvHSH0W/00Z2JIhBa4tWipqxIv5d/IjlnZll/K
7Kk81MzS3DRSmaIeBlhMrTpmpFKze5hebhSskDgikPDuO7KkQ96EGSNXOGEmSEUqGfTPdVYh06CT
ekKAMuIJU0Xjt4piS/kfZ9BpjLU0TgIkkbhOagXx6Ngsf5d/ZAnKSn0WmKSZRE0fBWQpR3Jjj4qM
LqWoBmxpG681/wxSkDqnAb7qVFRlsqmfjxqKnmAMtTLpIjNZcJeeZ+POl2FyQdRQ7Y3TEbaIVgOY
m1wuV3E96iU4a22CH8hnDBADrZOb+VOfOnJ4bPeqM6Y/7hBi+9mJm1FJeamlTzXW6Ljb8z2IjeSg
kqHsR2JBzn4T8ZBY412Or4N/UT8f8FwcwJxi5qA9D8De7R/rn+qzVWQ6n1w/Sz/JytD0R/uGqyB2
+t4w257GcR6IRkw19GPBSf9NZB4Tm+49W6r8EUQdaj2EMVIftQax35kWPO0vE+5+GW2A+oLpUr4t
y+BKhZDQ+W+kfLR3pgWuLZ5wPu9I/1TJdMWRH5VFl4rWxnKCePvLzjzW3zpaoYTjzoZAoqr3rWW6
ZmGFBAET0JqHZyjiLWO8saTHT9831Csu1Hxsgc2iriFAfdMvyDuyAeGNVI5ssflCbhwKJvzfLCXz
02u6uL8j9tKUD43gCjDaDMrn1RqNcrlHb2eAhYfjaGo9kca5Qaxym08itD+cYzSJN0ID/XL9uB+I
LTQYsq0IHXx7js/AbtlMYtp+gUhMIcxXE6l/LcP8/10rAAhBCcgadfsvNTtIDoj/Mk0wx2IGeGmr
gjCQFeRUvRkYNscukjnPmqsM8Yl6FMIXegIIUbs9NKkIFcveMFx6YCrUrrIlAjqEZP9Q+zX14oZt
PlhIbz7LVUcgmmugku/GdbkDOGCb1e7fB3NvTQMs3ywjYASdDalnUrOQkDOREHxXBiOSxY/SWe/W
H0xNvxcNnBK6EA2DHEuuswPSpWnytl1azUX14KshJR3lLvZcfgdjVbxA+atXRROUcA9T0rw2psEC
pFARkCYCkyh0PBFMO5aT9YDg8bvGXkLgXGImDhmGSvc752e4JyVqNy1o6KZ6rEXNvtNEnRN+tHVQ
nHy1M7ZF49yncrCH3QOmMpA0qz3t/gjgSixXWtBdaJwEkOrXuSt7yhi8k0FPXe93hJAWG3c01iXZ
wEU2iEeLYkFSEnkg8FxSV5SAIeFaLX1vqboT1+/IKwsa/PjQQ+osT7lv+T6nt+jU1HkO8u3M5xOu
QJdfcIho401elQZ+h3RBnAaxqSX5qNZnNvlrIVUUBRZmwQv5YoNES6QSoeFRR32j4M1XkV8eEbHW
PSAEuPGHoD9YU0tjOeZtIn2UigG1dGOYvS9iLlC6aiTnEIc0aUQvLtnqV4bHBZ2cu5UmTdUq3/Yf
FBNZ+s5B8ey1Sr9GecnpMcJvABAssCdCOyFE2Ai/B668HYAVYsZX9ntXkoK40lO/pXurS01BxuaJ
FH/Mz0+4u4X19SPSsoitUOqprs+2p7pYv3ZhI3krEiAJ3nLmc7zqlnMefZwNqIWjuH6OCIaOJMPg
iV6IwGPHR4CDs9qkw6eLoBqzukv1981ZHVaqcjYz6wOdEXGZOw5QOl6QhKKofb6oT/l7STvq9rhS
kHeNhaMhZZmO96Z9Ry3SRZyqFrPi3FDWVXTo8qbzY3H4oIDKfz2MHozbPsP6p/AORwpG5gPlhv9Y
JsJNtAWvnxLW3XcO/Qaj9WND1Mfh5PQU1MqXFUEnMA8uQCfkxuQTwSHRHoWmjmhp6qCObJ+6cATm
G9nanKgWN6YzcnQ5+lyFHlVXk+/YDlvcJ9EFfxVhPA6gL0Zhp/vYed7lMJv2MvILokhXXpvT3xkf
KP3uq80rkBC6xVOJtZpbSgfiztzLTF6uUjkBSlSaIcfPRAKk+S1DbgFfdgkbNE2tOH1rA27gS3Wn
zG26hkkuIqk73PvepzTm3PAeAmIrG3j0aB1nsso5zjFPy6Ewu1Um7GsYPl6/V/OgK0KrkJTV74a8
65FEqK2ooJMtbqgHVNE45WBzbgYmu38oiZBeIv/Gg+YATamJXHq9XC6ycpFhQd4izTecZf3tHr0U
OAahIo4pxkxRoWf1P9N0oDXy6i+4pZpjdQQCTCI/IJ80b/Fmr8DgiLwXSAcW3oEpr6+6RrlG0Jux
zTBSxYfPt4Vfuf4PXqf6EX25EMOeFsgnVgOSbZHTyTgeiNfeE18BMCmeIKXmCRiK2z4LVKLMrTuN
CkU1hMKmSXzyfHgJeBNiGmJpQYdZBUeTFbOxzq1iUnfEix3esI3Lbs9bOd4mymywk2qKFb/RYYjm
YNUBdvl+1Th5iJhkSgIxOeS60sT63gEdEpBlATvOXu1xXddHFmEKcAsfBElzVOnyIR2vEA0uXSFe
dTuO8fPHQD3Kmk4YZLv0N7cdsBHAmcb8X3CjhjmgUkEvgynDny56OPCFZTwAh/3fTPXeXSUi09+g
r9whbBz1SvW+1j926VMuAFAyuBU7Xx+akH/InKFLJEPIWQ7SJZr4CKtMZZXYePRVq1tI3J4gPn/x
BEybAjPhYkSjrAGR5Td/nCNTT9elG5tz3GjN/vscJG8ffnVmjagJVWAkDwhxDekU+ZvHmjXimorF
w8cIoA+WZW6KZc/stYofmmFEO1lNtJuH/njB2gds4+CM2crTPph3+JphEmF5lywXbZSlV6urbmZt
lF04aNcr4QfjogmxTmLNwp8tBnpYtuJH5xVElO2lY9dvaJgVgvg6SwctXkvfGHhmFaBiaAzbDrga
OQmH65NkIJf9m+8xclvkmeP3mo3fBPahiw0qde4UU+NUj9yQ2NmJaq5blGqYjmtjgPcnDDzHGVDf
SSefIOF4b/PAcPSkaEuFtlNgHcyo0MGDXaYnlnNe2sQcxg5M1Yn6hyzk2RcSflZovbbSPtEbSuYp
e/vNIKakhKmAysDwYMSAOKkjFkk3ZrZwRkdvCS/n0RykJrBy/YkQrCa3jXbO9jza3+odPmJiDq2V
7faAYtTu/lGCoqyRm0o/P5qdGpSfFUvwmW0VJjSmG8BUCp2nRnfcJIScYmMbTIEHTB+aAAsUD/Y1
8BZwSjps58ZcmPICATWjuKCoz9Jl+27YSsU1jq9z5uPPSy1fb+U7CN6dGNJ+HH6NyMMY2krcKdPe
s9YkA+mfyzZ6TMxKAXUsZANf9L3/KrhjYfjnh6rWT3nkLtcr27C3baQOLFAOnmX25jYVmIGLkS3W
ZrOyoQZxiSaL3GH42eWRwlNzFak2WkjAyhs1DKMA1mV4dUwTAyGmpr7YWyWH16VrTe1LnfHdVlCX
/WFRJvuTG2Xw2XDaO32ZsdE/3rciTpUpcq8rQZS8sPsOB9+Dy18wmlWZ/2qPhJc4Vye09fShZEI+
jc1iM0Q6Xc143DkcBpK//mvnZF4ystxebMsZciaY/QzUk3SOoPR4vbtSVqI7FQA5cNGEHcuOn4dM
HYDelffSYJoNwRqGtrrVNkuAlz5PPgfCwThbd6IH1RbqqBlgvMderE9WGYlk8Am+ld1dbyatSKMK
Avw6xfsFoQW+NYsy+tMSjwHciWnvU5imNgU5jOBcWQppAg5NAdM+o+HsoQoKLW9JykNlXGtUFi4K
ogUbZ11TvsMSFhByezORgiUgItGjozKlkTYm+lsIUM1ELIbplOLlG1GUfWZuqQXUzVKWDahLy+rx
lO+nhbUrSzM4PeBpVSR2IAdMlyfNusbD3ea4UHI3vx77Bm9kGWazTtdRmx6I2z6vGwmNu/kfMxkS
8MKdJ0RvtSz8EfpBNjfo2e0u8M0ORW5JkVSM/x3aVShfVT80j/jSitlkJKxetu7FcgFRHbkekaD8
NDrCQDb4DbUdV42BaO0S2ZllIOChou5l99SmUvJiWHxvauXjUc2j5DL2SE/RIKHASaKAq+FggbWX
ewOHv0GKOuXbm8ch10S4P1Yu3AGyg5m9VtAMS9l5ofKl9DLhCJe8NawI/c7Jmd5FtlQ8hjnoLAeB
EuoSeipmYtw/69a62rBtOcBBBKvTPcauyNtwWcf9aS4FiOCB24D4g1c9a4arV5F/OLEFggpiwJOs
nc+EPKnnSbATDO9v6+N3HtqND0Zwp2vmwX06EaI00U9wTXVNc7jWKfsIhwrWD5vKwZxdhZ9VBSQQ
ACfNJxeTUzYl0H6lzGsWs6kQ7eZ2c3Ue7LrYlEtXXiSUqAktl2glFwIp+Lo0kPkr1wFJjUc4gXgX
dKGvOfQ0eajkXxemQ9Y8cl+bOEPy4gtAb52jUD1pfA9bJBMaTmGZJdcpcMJXc2HbCzSt4D7kkHFR
GGqRwX9VmrdKI74q/JB4ZwHtQbJBSbaESJ7q44+mLRODQht7BWHqBgZyjbpF09gzKv9Di6fl2fUu
UQmyhfkOnXpqptO3TDJnOheoW0+E5ziOxlEPA62KCSYW/uFk9sDA76g6nuSgVIogolsl+J5Xx3FL
1yXRfd5ZEYDAO0eQSlLqBjc5Uza0zxrrrOohvXhLX1e0tXX9MC7wVQwePdQjqdJGU6aXpZyIkx1t
H1/2atzLm8THAiK2yt4rE5npSRwv3t71AEI8NAWTLc3bZjNx90R8AF7vIyAAINQDv/EFxBKjoQ06
cxCTh78M3AWVEFk8cB407xPx/8LydFXA31qrhzXjomqH+EXHT75+DIKoLZDi+Y3vOpqUI4EQbnxN
vmhaiqSeEb7gcRomfrJS2yVEW6nHWQB5UdtCaVTPrSnTx9xV4eKnDpZIN5ebk4YOltuQnNYJ5BnP
z8xoiwV+h0js9DooQuWd0ZFg8lvz1Pizy2iLUIaiqbaFRUBB5Cv81oTojPwwQXmulWNq1HXv52MS
ikn0GIVYVOT0hbFTWZGlxaVj9V0VtoWt87cZ1MJatQkoIuSJ5S5cxrSRcjG87JCLFx7nyVZrwhqu
ZmNOSgz6AqIYXB7amQTybd5DBjTPomEwtVzbZjwfLuMfkuVSDWj5IW28yjS37F9TWMSRZhe+md9+
oJq6fHxmSDXzROGKTZ5I5iEUebPJH5NnxgsR3YHwJZ5uQTsrd5m4vuFJxnkkcyzqqCtiL1k8/0v2
JKn6g05WIT3vwkuczhwvdulr9DKZNIM593+0tqzz9l6NhNtXiL6j6YM8MA++bwdzCPbZaPoMeMnj
deNPRHOsITbrkfiiKsP49kWCExTor6ZN83eevlhjKA5NTmdMX3yaiFD4MXfqBF9iYJyxB+1Zex/7
kjG2MVCY9dKP+ZFE/ffyYsQlPASUG53Y7DRvwK1LPv/Xi6NEI86LIWnihDKAPY0GywKu43Hsvmgx
Sspht8FJ6zUFu0i68uUht6JEW56mM39AyTcgtIZzpvjRFqYIkhq0DqeDuCO3SrhPu6Cc4dhT9XEN
STpwWyuXBwwZ9LlH0Ju3WnWC0M2zphTUHdk/wT1MtU9lSO2nTXS6jU9E4JHMu93sUwHZ1KT6n0Vd
aFm4NVrAtcL9dmkg1gxj2gEUjQcFEvxnCaw+LRPQKhg2+q/x0Hm6CXYF8Q3yfJF7Em2L4Y7Kc0z4
US7sGwydsSuo2JLlr7js7jj6xV4HX+GmLUfFDJKgguAP/Q8f4LBqvxvJvi4i/TxNNoFv+c/UDZ8D
9/wSLXdB29PEcfMuxPRcErfDwLFhVqQB29Irt13FRdXUCwTvFjrRZvxlwdQbV/rUYcTUp44dW01U
93x5vxR0akQvg06T5ra935e9yct93Ndr9EUThGETYUZfNpJ/3MUxYlSSIXELLC7SHcKalbMcU4QL
exuGLkj8EFsxp3uYsdrZ+lTzXUdkfnKPNCSMREMr5vPSmCVGyG6bS9G35DUTqEl4hZbtqax6GaHy
vNYDB2Wej0RdhhE6Oz3ODf9Jzq9MqO56Ztc+y97eqo8XomgstPBD6abaJfR2ZiOW0O2EGI+L+4Oy
1NPf+QoRHa4XlC0reDRs2UOWIwf0r7wFDqaqkBBXy0HH/zcy2lQ8xcVxg3lVsskqbeyjTaYh3RyD
vXV7WF6/XpjUUsDWNCUpzC2/LPHanrwgBurAmLTSznepnPcOVRmOx1S6qEUx2EALiYlXZscatktf
zusj+EAjaSLj48YZbAMuuWWYvueDuvcL9PUUxLpJoiMTqvUOrKk9yQNzF9LRRLa37uEqP7KsMuqG
eEuGJy01SVAB3PTdLKc74uFr4VMekFFwS16ATyvrUAwe+djcoOvKKrWlBQN3pzW3+k7MyfbPdDAO
vYu/OUDrwEPAPMDhEPDVKH1kA+f9ieEAhhNwtaHIIqz1uxhuOREjO2ckEaXirXFOgBgr+MgkNPD6
U3SWrQNfabLxZdhN/wYEsDctc0bpAuz1am037rEt3FL3Xb+9L4BEZUR7xI8biJqTzupxTNAG1Q33
fnsvUM1HNhwFueR5vFKKCbnMp/mvfx7rGxQiLboaOar0HJqtZx8YK+EWcYHxqMBhWJcwoNCBxiU/
OeVEGrYfTCQSsSAT+4dda2az4NYTmFUz16Qr+oBz6Z93Kamztc6H5/nEpNag12VHsqlJpfjQEVt/
R0VBBM7YGbgMtzsu1RFHLEoJTe3r+Wu2m8c3ABbM2GW1+8K/D+fbZvuo9xyP0R0Lbu4lLnmucm+M
R+quIO1aJzErkiHt9YifUL9r8mavifQSEQzjbqaLh3vxJ81ka4zvOC4GM57MN0ezmB/apl+uT1DK
+Y6l29ljCeGJSeNob/ZwEG6o7NWO+Q1B7Svv1c4x3zCkVwDXud3i8DpBTEmcvZAz3mzzrec3bL25
PJBw/egjDRthUFfB4CqRQ5m0pjHNuK/wvfYxrYjse2cWP7i1OEk6OjF3OTtM6bIyDX+OV2ZNteh3
3nD3f4TrigKBric5sCao1Tt5geE4jLwAUxh20idGNDIClKshsJFwS0enAJpJwgAC2CKTkR9VWvFn
OLnnApwkzzWp9hRiTKfumYGrEPpBHZGXBKhPyZAm0yo8vKhc7Yzm1TIxyVi0x/F/2NgHtC+5ATcC
7HQHExu3WDHV/UOCtYaSuP/9CVHnDp/xPR82hFTjP+jHtBotAVGh9NIzrFgYieD6Esw+LAcJKRuF
KkcLANFsWsSO6oBJxIoow65/VjIKNmXP9u6S+Rl+J9HZNT+6UY76JDlgw39Psuf8YkTGVujYXjd5
/75GqO09wPpkSYaBORfvPEBbGW9N+TvvrtcNedgtq+TIur4vugyOKqyW1OnHj/WeDDW9dFlWGdgx
1w3zwkbERUaEH63MXl5jhw6ZgbjtheB0e5+Md9/NEQPyNpgyehYl/0BeKmKtuoXBwqy9T4NBGNeA
CYoHASC47CPnuu2FqfpruvbE7vhjx8JfiBH1pAn7tZ2hiI+vtUbAE46sxOwjNegOJ0u//VX+5bBF
PPmYi3w+9Oslms5Yl02Mwy9T1KhBloVhA7fMBlzrhSUL68TJou9JWv8gNtszjf6BWBf5WLwWNd/t
uhrAnbYRKeMEthKTuo6PBktiiYfTTFfviJACvC0giTPJ4/LOMMgo3Lr/zYmTAk9+BpYuqbW6OCCW
td725kEJh3cxytlwnyl6N2odnYWadwPZb1JwBvd4yOVSzlRB9MCebMnRSnINfGEH4WE0qhNaQCg9
ynhqLhIL2pbupx96dtZPCxxicSGtbmCHpeklubAIfFZmpaaDSerNJbKSPhRhKCGXKeKMj1kBmnRH
klZM0JkogZ1h/kMgqHLFkMLdcc8VXB+Z0IY6rm5kshVyo9Dez6tVd9kBakcdvz/KI34+lKYV7QZm
qan8W9xcgcaEuN8kD/5XXp1GY4Uqs+A8unRNDwLv+vetRieVNnJC84xK+1hhIkVR2F+2NM7vPVsj
a4MYViurljj/t5kA4Oaoy++PGgcHPHOHfSjvPZ8Oh4zCU9mgMSugSUuKPiHs4Q908X5zFBWdHdbN
ubF+TAFSOPNIeAt1jHryOxY8F+xGDvZRR3bWuslnGRnhiNYabiiKGQtvn3/b6TpMA9e91wFhaO7p
wMRS2yTIasCEVx/9cIGhvOrE4aKBbgrCVhIOtU3r3O3BUQCl3OV7WvcO+UB8jWY7R4aWajTAWJcj
2Tzc82cVfLgm2OTET9QCCaGog/8EgwU0udEuGQ/44LktBEA/lioW56CfzA1ST6u2UDbjy5Rv//vn
1wpAHdi1v/pTyOfh5UYOrAnNrzt/1vg59PBy/55WH0i7uShPJuAivULhun5Vb1w9jvTYUVMbeAK4
GZjC5M21Ax7Ou28fONcXvk0IDOF0FN0DifR71IpO7a4+6oiA+Dm9G/SsaqWmPNp1fkotANweJ+fC
NLYX29bJy5hNZDynOyQGmIMfserx5P56y4aOySKXUUIfDN+bLl2Tpk86OU0f6LpvhyycTTH+agYp
g0dG/b0Cm0laacHZhBaWAevPmIFCvuooXTZiBUTUx6GXzAY60VtT3XXw2WDkBFQMNNRAPkJK+iCN
nMG/GlMuTOxVvnt7CvcYJKLNsSAJ+q77cO1xyVOqdS/vwlSKBR9ZkW+tXvDESBiZoXgmznVptAXl
kmIr1sHNm/1BGkyBrbqyd18oNFX28GLuaOPihTw2iEevC5IaV2VeAhf2L6NnuQ7AZ3XfriPFfvsU
bBEmIDpz1P3raLqqk493/msky1k4twL8eJfZyvzy3ivF7tZXPTOUQbOLCJWEXqsCPEYc+LcfFEgI
1S+eurZV7BgC537nQZdvANZQxcs7eBMW80KffSC6uVvVCAYGXrSBXXAcF2Bfb3roZgWoNXalYSOy
ftDdHJksYOmfEsUfVpo3vo8Awa0oUF1wS6exwVDkr9Mlc4FvJgPU8ZqA29kQYQWnai5JGm8mf0Tc
K8xSFoY333K3jEbhnWz2Xtk/Lgox8Wgr246mTaUuApbFH8KsHnxQKiqbe88y0WGL73mNEIdVohv1
PMo2s2Z9lXkd+dLhjJ7S8jgtWyLRTkY6+nc0PoMrZZBigx9En+n/6Ho0POSU6m5qBr80d7xyaeCh
ltn/7XZPsrAjDVtL9icAi1TcdA9lOVEWjc+3hu8XloqJ2fYCmulnnxwSeFG4csxnNV6b5ewTXGyo
N7PQMpEsjap34NqDyIrJdmLPOTdV3Zf7cvcBcYV9u1zNvR0JhqnKo2WISVx95Dh45BDlVFTlC8r7
u8BToFytFqA0CdQ9HN/cfiZUoAkmnYzE1HzMzDBd2lD+zIclNT2fC+6wL53mvnx1EnUPzVjk1nzk
7QVDLQ2OeJAO1xh1+fsDtFfM84+rTVSZHcHstfuK15tpWaLwh91od86ni9n/6g29apmfzc/TMJA5
uwB/knyH2068/bkimhFBR1WIp8VIU+C/hEnkVMibBi0ZTmzctK8Ws/SVWguymAi6zxrI+8wpt16p
6+h6rSbD1hJQlff87YeTFX534eKU2Qjzf4B9rbcLUkYHCnfUcR97Vm8aO2Ot7D6IR9TrNr338aR1
b7RGbcbcoVy7BPHBKP+2raMz39DMCGpI2JdvE5g7McOAiWkT4Fv4mlmnTcdrYMxYe23ls6zZMjgK
vmjEYEmQ/CKqM4sX8Aa6MZah/+04UV6Por7g7U5i86Fqn8b3FofD6/WUDIwxBvZCAL9K6ECDeEZu
a/cv70qsPi97d/eO09g8Tdj1VikR6yfA8n3kHLBiIRaarYzmDPgh3cPiXd+OYjfgiZ/LVMydCU8j
rbGPCvQwtNQJVRB+ngYAPX6/ZYMCzsi7uVzhLAc1Pwe5QZBSNQEZLu3TJgbvSeRmWLSeMfsqefSh
dwUuY7rzxalqRxhXlxwNOCu7m4iHIrezm35yprLrzqPoECBgA1OFVqRLnAkGibemP0AAUho+iA4T
N8YwxoyxhJBlBS/4dQb5rQXnDq79XFc656RM5eXzP7YYPKL/sRQ0stX2HfivHVia+dFTFuaCS7zd
w6y8yMuF8Z73PRZVenKeFdW4dmlZU+EvCH+z9SLQLS9tph9uyrxaDjhlYKFkTVLKtx1/rx7hrIEC
kmoFHAtS+WdJ+zqfWs3vUdRkGO249N8Ml78MzsLTqVbwEBuc867qVqX16w7DON/m7E8jACj7hE9a
SHR3mydqz470JX+4k+9fZneD85Q654z5pIxd3cjnowSrJ4fz/JP9zYfcbPg9T+4nyE5YH80sjCT/
qUl/pwy6CnxN0JiNCg4d+uHLsqvq/AOdjwiTyPcAyxJKyPF7EobXcLK3UI1C3ax+eVXlfCndcGsW
KEssxYmH14Sb6DK1NFeYuadiOc15N5sUPNFS08H+ytTMh44dvwl06lvpj4UjUwOjO9vejwKU6WoD
5PyLavstDP+ax11wSNNhT68JRXsAFVD7J9+K6e13IUoKeQlnQu79Qcmp8qBpgFAJMZz9eMqmMLPn
Yw8KjLrk4Sa/kCaz0wM2xA5VUsY4GTp+d+jXdCWsJ4pYNmjJrZZGa69ttJscS3oyRa8BbCs8x5Sg
63Gj9s8L6qgjj1GzMMaMPfTgWHUkrF/PwbEraJPWUKYEhvqS/yVNvwJOB2sEm/GG2mRF2l/Xa295
3dC4VYyGKTUtDKk8xiNXZ7vh0KK6Q4UF1xg/viMvbcqaoqRrN7igVT6uvVBe2W8iughnf8U7vuFP
xrSXrqaTYjIaeg5LTTSL9oNwFMWrbbjOpQYa6rG1m4+GHuU1B/3ptRg5ho0p96N7cYAkOI2IWxZB
xM0pVtJDeve+NvWduzf8V59xbpY5ZdbwRSUud2AZ2L8Ozu/Uh3r5ZJH5Swc/CbqxQ5kELWrXF3au
voU6k/CfweRUIV8OunPbpzReA9zOv/BdThtth70DCxNsg3e2Dx/Eco7tHm5UIDElToJzTIfeQn4P
/gCcfHydUOOfVfl+TBd/nVDdwDdhzmwsswB6DuE8GEpNfVUvs+CYksH9tXtOIXUl2otj9hFPVhCT
YWen6+cyXVyCHsOGHaKdsa50ktjzK92F1qbgbow4qLhwYHzP9M07jzCOyhZSNfMRPoEUeb7unwfi
wKSqpivpOukqjPye3Mrh/jE26Kexbgy/iA5WTWGamO6MASc/ABLl9OhJJhM/MS5xbFsAJrAKDKvz
YSw+cWVOCzg3ULguz617DamlNrICovy9LfKoxbIKn/P4oRUoQFLbWIGRneISK5upb3l35xtZ0UEq
NQMXeCRtbZ9VGAyllmJMxaC67+xYBc1ZPu9cHqA10hJ/6PkVqTiJiJsULHcbzgs/SRdWYOYLUtVg
6JgG6067NCi7zkwoPpR4bD5oXWjxuX8Zbu+AuRSs3xthK3z7+qjqx+f4+xVY3Rbioau8afygFQFm
ZMNzalX0jcHkvuI+QCperJE6JpJVHjJSXPffb+jcym8amt9RLoTaSE/5VxiBE2VTgADsJMz51Zeq
4G9azGSyqCZ8+v0QqEv2PikBBIEw87nPqpY5e0z2X4HvjXrfVOsYKBv+FYA5F1O0U2O3YLxwyv0g
KTwVnZU9HH3PdGaUtcgQvKdGpKC15xeiHMx48008NARRu4eHoDwE1UK0z1PTeHvHNcLwDkGho9jj
GO3uxnXmnVa0olPqBEgmRukFLiwB1rTHtyayXA8Py22ORk56HSz6P4sXWFpNF09R0+tkpIfpdzmJ
l1XLx8ENF8kJebsvt4yXC81f784YlxCsUygc0Ac/2fdWN4iikXeJmOhzQQKIUKUy8tzbpy6iBPEF
tDQRhWmjW7fg6P9CgvdToOreRzgZfMQass0TO/hd01Kgq28I7sTFrJet53LdaKsJJveWda3bxja6
hHTQybNTs9WKUoLKkR/OTfHkB6ZpKgHoPWuBO0KeNHmoaiP5+9MYGkFAbPA4V2o2JAnc2nWVZbnp
6IDyhFZJJtDqmwsiHueJOF4ETsr7WIB1r0Y7jsk4T7oq4PozXan3WIf4egCGJKykm1cXRDpwhrEJ
K2P3b0MrEPMVplFAFXq4fS3dBZvgp37hd+TcxMx6a4VW/i5WmfFoXG1WfFupOry1Swwtmbm0G/cM
A8L/XIANmbFZYt+UT5MhynvGxsfKsI5uqTg64NbbqTGXaa9BlKG9e5CWDOYDUxURRlPjO9qc6+t8
afTyMpY2+Lph8wbRAMx9T6Oa2HyvPGU7eMbVrTJBDQdZlXNS9HKW/F4xBjK4PeHaq450+tZJNlWJ
/wwwtS//gC0JsaM01TfKjnu0nlGrSAO013te5nNuwMAsgRT11A3xQR+g8GZ30JbkgiJ0M3cUS7xC
LojBwrAUKWCV6vF6cn9m+gX4xW/v7XF2UyVYTdjpZATcHzVEv10FfQcadBGGwUXUQzLQflrHWNoH
mOIQr11KgpUiAvRYV8oKuMR9a1d93Tn19+ijeNXp7TNbgFE6NzDRpoFpv2RJAxnVyUGslsDpJ9GJ
ZiiQnbc4ePQ1syFNgcePU6yAhyakVafbFiLY6Ry54f642rtM45pCiWIrVdTA90YUHL5K/FDVQzTZ
PXi/3F4zBl+20rkHS4xo+zMwZPcWOHXhk+jGPP7WzxvRZco3OmMwcbr2EVVnLZPofXA1fdtC2hQN
yv6AsFWKpS5vtig5DjriHGupziOoXT6Gx1hALbkBoFfJjhvyOwvaVN8XBisdt1tKifyM1klLvL2Z
fZ2/gcKcYnia5HYjVd60BKNyGpD71yiRzHIabswCVEYe+gQw0WTpFSSwQztoVbhIzkoqoG7ge/wA
AoIWXg9qCQSGlyF/a025Nokj47Y38HeRSqJXCjmcEWtVTvexYQL3rSL754yNTY+7ug0LE1lJ+Q0X
PxhRo8LZ4+RLnIZMKkd1gOF9gqGoOvOnCRp1bw39gD0iT14tIc2jRWRFd/B/Bt14QL0Sj2X+RIIO
d8aq6Y/lgVJxWX1ZjvX9++BAELWpBHYqAf/So4HQHtcfF0VbJNssfmQAot77NiBR/4lljkeiOAyF
M1a0pTXfFJB57n3gG9QA1AwEbYefDC2IVN7E/lAg6r6yZPIdmEASkbpwifkmooJdAoYehUEAx8/g
qE2DWVS+XHHk+UzsKhHHaQIUuMuMJZTYS9KhecFVrjTlAMLgE6pVA64F5Saguf48KHt1Bx/YJgOE
+ZRM/wW9JMNZj72jM2F/jMuGa915wU5NOqABcvg4WwvJWm+JQ3NVYFVY8S3wK047bqxHeWtKDr4a
OhQ9Txn0JijQXzCF7tvGrD3o7IpM9B3uZbdzwgfq5sbAgwnehy2ynPNOGudt7SdacKlxQ6RsnhHn
o6cipPPz1jJIUe1W4c7U5qVOx9yXgWGrFGHsORaT7gtKz+2zPt6Q8hT8yIDkl75+1ldAVAW4zPRK
Ck4cS4va3Wc9lb0nTX6GnhWO4Px3y+vl76fTDgluV8rN1qdQec4D6BsU4MZSWeDZrthRdBt3wd6a
MOy0/30Ah7K4stTRSwXOVjrUay1VtDKQlfLu6XnXxKn7agkm+kAbgbOyl0KGeFg4NI1+lctkVMDb
AyyFRk6GyOIriGx6v/QAnew6aeW32HW8u98HZPgmBM+Z3joMnZUUZx9T6Fab8P+vNETYsEcSO+bN
kqQIW2/4TCUsIO7KnckRS+Wo0fl3mEy4dyb9S4F1rHyg4p/kHM/WW3g3tm07NZPG0HPVYvmieJmL
zKR9sNvrYhUZrc17GipG4u7Z3ASY7rBHReNz/KoEGCRSAMbbXAz63T5H9WueUj8ur6Eq1Cw0hY7X
V91eGa0ljs4A6foDa8Uu7yQrOAxTRt+zUgWpoE+jh7f/yrwaStxl8dVoQonRp11a4VUq+9/S4UOz
s8ppgcI7CG58J1I4rpkBQiEmQWBuu32k5JsMKECIMRzkLJn61EFwoH3LCeIbPM0ph3qmFdkCeSjU
FoJaq//gS2jbYzoRW1y2oeOK+/PofQO8XOu2kUxLbfxnQSfhPeCwlJldudRVO6ukjICESS3h5hrn
/BdoqZQmlWQPp/ZKHwbNWuoC5Z/zMjjP+Z1omftRM8akwH5nctBVz0/CeZEI2Nx06NYpeNZWbjHe
IRz53sb2M+EaKRVnCbbGtinemMNahyWrerTC5nbqP2U8TjxLomhMWb73iuVXYB2DDt5aHygA1gpT
h+2r3/wIOSbjGLurplut2DpVkatkqZGEnXXAi1q0uZa3DinElyE7mWvke23PUA/Oc328DEokrElC
bQGBeJ51MDt+Oa59xwwU5BwlRHgtqO4NuJAsljz6pOKnHxM/Il+BG5r4g5TfpZd7mnJB97wsginN
0O8/ECZw7zIreu/W+ajkrXVY4ufb3s0mq3BdVbxhz9t0YcdZId7V6kA3CW4i9FVpyawAByYu1yEw
HjtLOT6alQIF5iSsW8E2+s8zaJGq2Ny63nI/nUUljTl5f/EZowJp7KRTPUvjHCBTFvVrQKK42+fR
LSUojol6E1bwREb5HrnyEQa9GnF/IJBDcCYbLQKczqMLRm0ysUPdIZ0cIUdXFRJIBF5qwmi73OSg
xivsRnyY+ORuxhllT7Mk0FtJlmstbt8m281wjdLhIyBkGPSPkf7o+ntknGviFho08S7Xj0OSQ50k
TZZbz+CIZpVOKgbDvlUetkiqvQ28nFpK0pjuNg2b3JzJCxNJAViHR3Z4OrAUqLj0V22+2dB3wIeI
wrqLGGzX3yIQhMu30Rev5e779Jl6rExye4J4FYg58vyo7OpZtFUXUI9wOvnY+3G+up40+Ym36ZUB
bLQQSC1VxIgLpLaHvAidNAHSsEvp7OAX2gC5HxeNA3L+YEMAZKvnUU5VLDTH4vD+N/Ux1almn4GX
PWf1Tn9i3cscUp9i/+kV9Q9X3GlZ27ormHGsI/HDFm3NGrC2ynZBuLji/xWozjbVJpr7QISO61+G
XJdbXsOLdOzSDTYl4hmEXuHy8f1yebm7LKbiVBsOcuCvCkilCCnpqj1qAzya0KebmeH9rhLEzWS0
HpHa3gAonW39JaQRsJoOG7Zy5DbuHkJeK7JLsbndUcLNGLik/cxeHz1nHmRzXkQKQEoBbUNvvAgp
JjI9WgCBg+rbjQILRIyj3ng8mfTcryFSEbDxLsrsVKUAobAqvagAoKiiLqmjtStgrOd6Ulpxzfy+
GIB65NXtYpDSPnSwYgI3YjZpBZB1g9Zg79k1+7WuiwyUfw7bFwtEOpZtuYJGlxoTz82wXw1JiX+J
gfrtY4jUchrA/SNFDvbMHfpGUO/+ax1BFeC68V/SgX9I3FLOW5wmHbi1LkP9Ur/blOEPZdUlLRo7
V7Cw/BhHEpKS18eSUNE66dbUrIA/B8A0fz57XiQvQcV5bEMJnjDq0QZevVEXl7OGAc5etMaGJjS6
Cfo5g2S3pPGySI7S3Y5t4eUsX8AHTNM+vX7RA9+SF6z3iQPfW8+7meYNaRRmJncZnlZzThZTtcjE
Tt1Tq31bOfH+AHKKd3Uq7sAkbG90fyH4fdoo5Z6DuhoxnGqiq+WLCPgaJ/X1MjfPK6KmMfMmxVmz
nUBFcssXXGBp+vxJvJ3LYDFQa1hHXGe9sOtBt8+BsZr79MUs2Ck/XcW+8zxw2AevGiaqR59NfXig
kLhb8mwn7so6ij5fyDj7xXe6qtghe7O6zUegq534X2fXxBm6mHiLaSuJFyArDvrIcqAMx/HupMfT
GThxrRxt8SaASlfJksXabxZJocqBgR0APzMuQ5ZCsodvEKRaZ+73rg4P+pahkPbYnRsSe7hH3R70
J+lPtWIiDNErr09waYoPUu+aV4zSAE1rHUDpsQl8J+V5yROyEmiN0yB2f31QAgVxXNZ9unaErV75
kSBI/4UqW/jmikcTqsz7p+qMBmQoNw1kf1Ar70y41gK0ZM1cV8XktM1IfPVkjNzzgtMRCDfe6L7N
PqmU4Q0oKBjxCVB452Crg6r60i446iBE87Ft08BOtrFu8FFRga2bD24lyGHDjRToA867sCwZ0Lth
/lzct3D8CewCBJTcUAv2TadSXe8e5BafG4RRSIcdxcyxva4kENiiBFRiTnhpfLIbgBiCgu/ebO0d
jHkDbwAsoxzbwwzej74ZU7GgVN3CZW9ZuXgbjiv10oBNRuW1Y2adyqhJSDfCSJDwe2nbMaWs15cL
nfKmb78XB0xvd5AC0TP1/Rq6ZoyQZDg7m1OKDj0A+sEPtF1+Gjy0TX+LufgEtbXDYdLkmM5Kn1US
pi8hT979ZkINOzKB3o1tzckjTQDijEwqpzG0NRZxYFCP6R6ZpGUaluvbRaR/oWiNY1tyv2LcW5HC
u9m8OF0YDvs+gKrBl7ys3x4Ev0+tFPIUNPVOwqaXJ8t8bOvUuPWK4t9FpIt089h9OkvychquW4pe
iPBDjC3hgjwOzhJn9Po5soTs/Oa9CzpqpZHvOZz4ERNHhpXKd84+Fp0h0Lq/OdV1E3KH13l07oRl
uJ4JJtfqkSSuzXxAcO72xGXP5LdaPP+alU81kiGsDikoh9u7K6+KQZ8rPj9/ZpCCghNIEW5AOI9j
D2aw9dh8scxRu11APlfon/HXnRV50dVZaorZTIuRLw8C5DNhYGZW7ktsQP4OFkt7rKZ/+ea0k5VI
Kn9bpkTZcLmsZHDi4yFgmk+O8Lvdgrw4TVTXTFDxjzNi8YUCgKjkkfoyOEdNpww/gZTKFbGulgvG
BArlCihgpcYU/exPbGsxK9+qNppbxDvuvxyYOFWRya5LvN+Dhy3m4ctLKT/qGzV3yvZ2h9ImGweD
vIVa2sdU9cnfXgvlXYTz4fksBRn658zvce5A9xu01/PEHoCEJYTAX5JvDMMb23XxVOGflBSFuV/s
OpZ5QzTzqNbUCgHcMGnDIj5PQD50iVKkVgkXYws82eh0tjiWnQiAUhLzWuO0DZMhJnCdROenqlIX
nV74+G7Glwe/H48F9slwA3901T8i7LRwug6p2UL6RXH8t6vfgmRmaKZNu7ZRCEamhuGx1l4lQX3O
hvAS719I6OgFigN/UN4RPTdfODkFFpsn/1QeEWU+hoCDtoNS7BaHm5shfzjZcz0uyPsgR641wYgA
630vm9MQR3Rpt+tx2M5UHe8Ba3T7BkXYTsIltp+RJNrWu7l5mRRNqMCuk/uDmO1JShjfqw2H3nC6
BmGPmO5skT8yJifdowiNFj7Z51z+DBpHHhPDPlakYHhdwwZ8Zaa05g3v/iOg3qb/ch/gnlR9G8zN
Pd4Lc57ikrZ12gu/6mPwPuMorjzhyjMTZ//XCgXxyrroxSOr8Qar6HwOS8hk/2Us/uqdyMuyxZ7B
ytpG4zz2dmtuNaPbG1iLQWwH5UZDdJbm4LB423UQcs0AQGJcDs8eRNCDxeMs9H5FCYPQDw3cLm6N
XN4c/5Jf7UwNB9QH0Zwtmb8IGPq5e6u2q+mbrj6vTdKUmYiQv+hTOX0VQNQX6sWUarw2REVPvP7U
h1oTn/vdmycnkUXwwcnWnqxyE/MQSOGGjrIjUA1dNZudjYIpIw90+5WzpczcX986xwf93RPaMLV7
ZAB9MnnjZUncxUoqJpVW6IuEWx5/OsIXGe6N7yx1k+bciRVind3u3vQgK8OEc1pFT3fL9PzAiLmd
YZoCpliRfPq1FQWzFv+XY54dOUsva7lzSXGtDxy7B/+BJxYC2xRI+WPVLMTbU9iFBn5sajK1fuzH
lGBznfWaqE8gODVxQk775sb1de4t0an8ffO+aLBWu9Z5SqtL+HIGs++6ZL9krfKTj8/jvKKQP67H
WIIUNS99ffiDE5ro4ymj2BECEVzwoBJtw8Z0XC50A++XcMdDiBL+rl1KLQJ/w2dbRb8lU/jLdVk2
XviCQmSgREU6JHCxPjphuCnjYMVnnzvQe5WRrF54DvnzlW/P98TKORBnqtYH/kbS4r41fM33Z2rA
5gwuEgR1F2WGLXtKIbd3DJzPcskJdVm+kKZSQcQ4Ny7LS2KEzKj/Q3nzMonp963U9heo4J0r2dwo
Dl+oSHumq/I2eSFLO01zNFXDWKtMVoXRZn4/6vYEeerv9zRLjtQ/5kfmfKp/YC+/YqtAYvJSekJL
hwWg2/6skoPNier6WdJrnnu98INIdDgvfWXgy4lZ9ymwjoE2/Gm4ZbDF3WFJdo6NXD6WvuxeOTuQ
FRawyb0aRMioeOsLLxk0p+FHaTiz4bNTOHSJBNAgLo4xBn5lMplXPjz2MvyX/3oe5dKVJyriB1ER
dGcLc81QnEF6X2bOiEO7NxVBQZMyceCH9G6C+qRtRV+7igIpAKYuXCAFui8FAeeys2Orh9e5qYzg
cEeL7OCkf1613QUnh3awbbncNSpozn2Vkpq/WQH4Ulup2kjTnFFsEvL6NqA3DNxEpDdTh8fZAVD+
aG01FNJQvkloGgngTkUubYc7i66ah9PtlJ2hrHuDeIJrdG+E4CnHS821NwT3ODoslxqJ54JH5Gew
R9eNc6FsJfBRlN7wiQ3vdqcisKgCkvKYcBIL1+XLzwxCxA6UhbrDteHArYD4nSUh01qPkXh7AsW8
x9sjXh8JO9CmiHNizpG4gQRwDId8Z2PDrHC/rLGFsTsbNg4/68dxOYB7+PEI9sUrHcawEgAqA5Cp
R+hXMhIWc/iPYkZ801L9xPlpSBknkuFflTm0BJ9gHZfd7dLhCtZ+kFHJurPt6GmwRUxLf1bH0j74
iFs9TL86sPb2Kh6iCudsBgfgl166gImoaRnNajMRPlpQPYTH4NWucsi3UuOG4YnQDxe4NzOxEd2l
27bPWPB8YiuuZPzos/HR/pVAWh10ASIxJsmz2i/gj1Us77M4brJxKqhdi717Dak4M4n2FseeWhFd
BC8+Jtoc01F4ukj96uVXNwQSZ+6CBuxvMWpvHGRYM+51RX074VY61Pj+e5SI0jBVrp4eVKxLjlVA
kfkE4uW2L3kIJyNH5x2Rilb3/nuotjWOmYcMAR2WmsGVVk0gQL2OlMWgDyb74X1MfMfhCBXTDRTW
RW8kad1BocpB/fD/pRhGF0ejRe/LOE/dnp8tReCX0cqF8G4xtFPiOOrWFGi3iVwfRMVVDAJ0RSq0
BybNJ362TZ7aSJWwFrtuO5mRkO9XiMsm6lFq9/aYIFY8rPHza6c5vkgO1CT4h+5EoVdlRAu6d8ho
EG13BUZoWwzA03MFvPOMAQmgm42dtQRwoFHmGKUeijEileCMS2bQHrlRnBfVIVk2KFtdSUWHpC1g
ZK5hAvfCw5DPYmUIeWgEDfgP900O0yRlmmUzHpuBnAPGXrcdfLy397IXRboHiowG0NAz3VEx7vQy
XstVMBCLenDqSdijqvcJlqMCjKPtgPOMeVCH4TWvcpHX74BIMqNaXDebrweizq+SHXxz7GhPu1A2
D2gMLuZrmdL/wuerykRCBYCXgokYjObvvNrrQ3cWrnT/XVCWj/Q2O2rMkuY6+eKGyPYjxILJ7lJg
GAboxKoR/OvNYTTNoQNOJ+WxU18Al7yREtVF72uXEcGkpakd7fzbi0wTH9gpEZyoShHR9cOoGhUY
KJq5ieVBgS95ZVA3FrYAEVBidkYYO0QHmf3rkX6IcyvlQ0slsJyXnoeDhOJsHdZM3bOslUiNIZes
YHFHb8X7KWyKXnE/V06gbPryIjgpLhGwblgEJE2DXIiiLAHKy4nScqdks8FUYvsEi8xBUVkEZnUQ
c82UvYHJf/FepNdznR5Ssf146SSGhVYcUzHvankpeOpK9UYYU+gY25AEXvDDb2J4ZmuXd7Zramce
jW7OUwHF4FngNKzT0Mj9dSz0BfohMGu+geRy+ohgSL2VgwgcQOwu68P3d8tymkJZN9eMb9mAyQjt
T15ZuDc+cYCSdRceN7cAsVfFFnwTUs3kk6A4vcO3d8Ecn/5krFZ9+lwbE+Cd0hxJcqtTwpE5ZEHc
4eooJG3UDNmGNY7TS5OIVFoQ3tkS+x1PW4HaafwzOAfFPQDANk3Td7pYjCzu7XUjrcb/rrlMKp7v
wpRWFEamvhph+z/zMeTkfQ9dmFiMOzUxSeiJjbZXbMbdmwih9w+jlzt/L/bkUpuHBNmLGbTRJApt
25ss6lyMMzz0wEDUO8VJnQWva1P5hb8IUcUE3SvjvH4tAJhyQfp9gd7wR2wEIoaMOYYj+NNG4IK5
hRxXOchzsPUnQ82erqfb7Cqhnqif1KWy1WLroZtKheUy5m44NLQKiogVCVsr9IXKgtq//U/VlnCw
SY9erkB1zqNIVRIdlJFGP+vJ8CqzzyZwFOdaejI8z46BEYRWpMPB7DI/mgtdbncP0ilEVu2gTV8O
iMReeEENWCQ8PbzzixoWLJYsClOigpZx8IJVCxIiNKVJ8/Ocv3+dBddZnt8I2P+6zFA5m81wGS1J
xbcjW5dE2+RnHOSvZVLduz3z+cmYsOvJPIXqLq0LUENF7sela8qtkK40o7f8Nl6jzqjzIgjYdMva
XhDW+QlACKyPj8vHKFvGwkJA3NOGxEFIStTGnWB/B8V//pLf1dnRVrBOFtmwVqYuIlT3689mRcNl
DW5jsB+AKo2bzyisEuNEeY+IjBl2PNRvJ6CwXrdGJT4IODZzdSB8FZt2y0jT2ES1Bd73dWRfrX1R
OrTKd9Ugndde8Fw/T6hZf2g8qglnP389ENI8H6i/29jfalvUa0GWcW8KbX/VJlbshHI4g3ljIp57
TWTiaZrqFXVl6EyfnHcm0kuolAcDHOWRICZJlfoXw/qf1BNF6+fzzJs9jRIZ95QFe5sJqudvvhmC
KbUNLWggUK5qza7w7iqBCclcl3ae7LFzw+SxRqp0s90tq/cFiEv+vtfBS4BNey1FOuVUBMwFi9e5
0fmK69gQ8JI69rDyKlh8TGyl20nhxbncjiINDoLIxKOGo6GBfPoS59gm0cNBGRL8uxgyivpwOLbE
S0QdrmHlzhmtEFkgmV9+DzDKIVZa+nKCTxIuECF7xe7zseF1zonjlN8u6aVVIeaHamiOqi/wtqTQ
HeMPANRufiY1lHskvikQWhPfxssnDSoZo40YP3YlKpP9s/YPJzG7BzpqWL0+7+tstDun5NV9hjdl
2r0Cut0fgfFhNPSzbJwGVJtSTr/jMJom8JU0wqj3i08kd2fiIyQI4Oyj1vYEJ8r+x8kSP0BNJGN8
mGh/a3RNT9XKLtr5pSBLebNiNsuCad5NqpsEbP89yUnU4uW3lXvfU2tzLSRlgr1Jr6OW4NZ5Yxci
JKXfXh1lePWR4i1AJ3QQCXXFFYONlE+fzlGgSXkvvtfd2ue2SiUTpkq7nxv2aSx2MahdqTF9xOI0
yCuMKECywxCDLftFvmnXhkiHBpym8fU9S/gFxMQhzC/KcQVE+XK46BT040HxXOqP7gkGZCotxcOO
65teJOqbEiAt7KDImx+wsTaNr8JPEzDEp/1C7c01J+gubAbtiZaIIXeVvyzeuuxD0EhG31dsruDA
OhMhJza577GGpFC84ukfeql2Lp11jfMQV12xgkAxHm0sjHe2yNwEVYWgCHxxbul7JPzx/dRFlCdc
IO5jykFoBwN+E0X6CIX6k9UeyiK/EI3luXJG3Mri7drJPP0nxnbRvKFDuA/SGpp02ng2GjaPgp7C
RfplRpTECoGhJCEQPEF5ODBQhlVCFheNUI5zOGveZU6kybGWKmAHusuV/n9BLot4qY34/Qlt9CCz
toHmg1b52nVUKEx941skNVp3b7f0Azg15DDY3BUc4CpliuiBp3bT6Ec/HzE5EGejzhpWLuZRVFlV
K/4Gx5IKKKQiosRKxRJmEMe9VsMicSb0HPcxtoscG+zBXl48NUz84GtrGHyclFGuQzFVwLFJfxmH
YRX11SFIeqX6xaa21mX4GsiCbSiQq9BElh+jlOSvw8qhG+cg1sc6H8PWvJbRNsTC9/ti/Amokr4O
53kGMUOdcGPmP0V2bwsJwgd9P07SX+4tHdG8yu6vLWQcKd6TMlm9dIeIkPe7JEy+Uy57L/J94C8x
6Ow+5U8rXC+8rt41wm3WPd5pGYRTNzDrYl94za4ApDDt2dIKWGNTFOkApknNvn1ecju7vadaIUwL
fpU3LfiMQip3KB0HsbTjqhUxWde1Hdo1/XqOt41jPWk2WWCjGBQQRGKIQIISAejufCGzwsMwpNqL
8lC6XQ/JdyOj93VyM+xJBHMEmVlHvPr0eo6YHTovSx0sFqfxXUBkxh8hHlXMs61sa1qiQ5o6WdP0
FUGS23UNlY5SorfdxRUIwxsB0do88FzFtBxUlzQ9LCPAGIEFbl3x0R+TEa1OI+T3GS5JTaU+8x3D
tFavw/s5P46wwOYhce8ovbtqJIJ2zUoDihaxq2hSdFtTOnZvcmCcWP3XBH86MdZ26JjjqGNb6J8D
MwWksBttxYrewdvt5rp9SHZyaUwkUDG8GzOVWeZ/5jLveCzffd509hLCfes0tDO7iVkYztmPWO9s
6n8RlwwiNj2rn7qE/aEhxSzJW1O5nWaAAu8bMZGmeu0TQOPQUu/mV3GQw+9EHSbzDSPP3Hi2UfCd
1NbVmzNjElHbz6+wZGW+vCR/6rYvjQSl6Svi5gQ2UX/8V+by9OwOcX/I2uoV4bXODQgIEuP/RaXd
Jv/TtZJH+EvXYTVz/UXLRbrXni8Ik0MiAbdMq49qSmsI0qBmrlw36EUjsKYHYT/9dbwB0bw0F7Sn
PMtoLFDzbmXD4Cco3FGtoQMzGSb5VLBVxdFyJCzifuW9HkW2k0iF3pLzKMfDFByCN84gchxRLQli
ddgUz1iQYIfS9AQBCs9t5MyYWq5LSv4qyrX2mWz6HtOOGecthDVFYQccnd0Ha8/Cy/UokY2WqtGF
OdUgfi1JsTgJsQkqc5e9S18w/jDsW8x/cGoQD3WJ9v5GKU5sXGwO/BnPpKkJ7Gye/yet6Ez4jgvR
CNdTfXEjwAznjZ2lsdUywyba3FWLYLngVGaze7q39t01JPzeH+Z1CN2OMdOc+WtLr+DXmb/xM67N
0H3j8Rhit9p67eRi0czl/Uy9DlZ2IxvwrMhwOTtzm97BHDJIP/HEzy8OKX/CDIlhsfPh1RGsDrBX
kiOphqtKKnrvAPko+GuSw66fT0X6PvgEDB7c4D9iXSHH1YuwaLioo8Yc5VMMcs5zg6AW9roEq1Js
B6yLTFTYElR3TDoaydEJewF+S+C1hlWpMRhmkjVMc5wJPylCweABu2y0h6FN0EgKhJlLK4lFR7U7
zSV0QMmhUlgHP49s9+vFPbV4/MyNqpphOQ/mHBmX+Or5h5gpnVSI71TuCgp5Nb8EncaTmgdD6dbm
8PWda1xXRmuHt1+Iextq1P49xldlWnUrGIlos9b7Ju0UHMDk/vGg5Rg/yejJQKxcN/52Nz2i8HBS
ySYluF9nmbO585HRFy86CsS8+kf/ZBul9Lft+KWucoNNgyx4aXm3usoG6QTv3BmnsLVoU8TXhLpC
oPW4fhy2064oDqbcpQ5LK7Q7b/K5nKcEQzDHDMmS/CkRdPLnV6acZ12p2n+UaZbeHIAeNW1zBZ3r
mZ6XIRobCzExqpDcr9y0JD0AdWd2TaMziSrsFwVpzVArcFVqehRal2w744BlFBjhw1mg+1SEbaM6
DuGW7QxMhNH9vbgigsPena7NGn6UCn7uMzo4sbpF2DxJBkEjx50nT1Uv7WBBuwWF9uibZy8KMHuS
NStgZo2rxx1GQnNiErH3FeLo0Hm7NBv9tUDZ0GrmI2Uib5knUDTsOnD5bEnqeRa/lODiL9+anguJ
m/YYixbNaKhLta7yEJaHRBAk99pK6VqC646UvBuOT4gs/MSzFke2C1wKICUEnT4dcrpW9/LhilRk
HNu94mNfyKwAmlvKTDJT77PZTgJZHC81dB9qajVKLuzG9VNa1ZXLlrPQgypiJxm1mgoYYJ15pqLW
NKUBNOA5T4nvtp+WGoNjXbiSE4BQyg+wDxu5vZ4rmhSd3Jyv69KWn/n27S+n9WMSeME4JA5opQup
TY77ut2RiUyX3l+MFjGyuO/ntx8I56MQyb0fRkuItrVQGZ0ItMJaJtcA7A7PO/XH2QYkJTZHBKtI
qn9ChBNMre2jBSPK044AWGNr+w8jiGO9NYEgamAZxnGjXlp4ePxVlVEpNzvJ0VO7ep3tMRdNddDk
fn8vpRWonNd8qju5dJS5mf1NuHPpT7L87OrE3KIm0u1BZ6HU7s+c9gzzdkG1qAng6gMn6ACEBjC5
ADsOvGyaBX28wn5W3HLMFiN8J8u7ZRHl8B/55FMAp7lWAks697i8modJgGeYkzmZGTrXTWdJrQ8Y
oYXuUekHotYTC13CvhQjy+4iG52113C6FwRSZ1tmYchZn/+Zxq+1AlX2R4hXIbFB/o5VYfUIoG6D
cierzMWkFRAxzUE4nj/9kpj8p66+2XLrLAKLf8VmAvIKM0wqSay5P1mjeS4+LIE2thBAj9kM/VBa
D23IeKqBxSutX9ZHDa54wEIPBgLz4P8i9t52yN3eKOa1YyZrylvBDtHOVpXRIv3vshFoAPPPnIub
K6wm4C6Lja4b2ociqY3XSQbQr03QUBiFA19F6aqy+QDjnNI2svf/VSo//XRqw/VHUlGMGBeejw8s
U1qf2+pWnM9rcww0/dHr57J+nu1L7zo5711EaIlD0cnMIkb4Efewgm1JCOORQ293ibdKenagMyzX
BxazVTe7MONmzrLrp1QKRlEQYhLcfTK9JOab+9VMaU9jwSej5X5oiiywS6+zR+yfIzayNSZBx0nu
BvshUsnaWLfW4s/uIXJ+inzgMwDFTHxt5lCpLGWHjKM8cua0DWpXjp3lEOI54yG1Z8vpOTy3vxo0
0abVx2CMsnDybbWKGNJH++mE5xvpErD7vwVU67Lh0kVRET2/VE2uP2i9Vd0FlTc5htaf42qNYLnK
x0ETtrUVp6PFLzN0LHPcZ9nyvXaAqXU+tc3+xACsKGExDx/1shDRMa4x2wqAN/3xY5lssggEtZFs
Qv8faLX3keU7MPKR1Z9IKiPvm6dhHR35DWAgrOz0BP1r5Wj1pVYVqydtFnbTTivO1cBVrKbOG73R
9uL2xksFIb1L9REXt7cNmlS0w3m9eUaazmXsSGaHRHxfPOP4ucUkwDFAxKk3SIn0jiMOs8ifTbjx
dSgYD9o9PJGQxb3lj2LN1ERSSpQDBZLXR9KB1TtrQUf+UaByHbfrZfVDyTvCPFe9jH1nAHXc7kqc
cqZ1nVV/AC+S096IfOnFuuT5vJIgwWqU/wG9BE59b46IVWBA0Ir7SqYHE5fIKKcp9UpivYJkQsrA
Iig+Fo332foQGjl55cj61N7s8ThXUmOQthd+Ed4cw8Sd8ABBYbmP0NHWaMNaVPKsPXa7fyuSdGka
hH0FLcFn1fS6Oi920ltC/9h1K4YotNilqfS5y8T/2SNJMNZ6kh4AMdyqbHaus9jspzM3943+kuUX
xi6AF86cJg5iC6CKee8HZkHoCkuHPWdSIOX4HCY1tl3y9zLakBKvejcmu1BMEJCRPvDwbPuJJwlO
+3UVj0J8bk3apy36/Ka9P2En1h4NLF372WQh9lQooAYQEHnQe2vyd2dM65mwhVmVeLjcWa4S52sw
gg2/vtADF86nyx/LQwTou/mh2AUv8XM9XhVmTbBFjCi1YsZQSMX1C2apdjSGis0Uhs9dy6W3QxM7
qnzSd0ln6/5bgn5gtafur66TZwAkCzps8UfgJsH4zHoMOwzBFLBEZUQv6NHGqRlYEZlc0bl03ZXd
0gaAlJfExDjnTnDMB0zRiHk5MrA+A0IkjxM09P+JHS2Og743MAkKAEtjEuankyiPQRu2FOUN3SMu
mO9WB3VPeW+tNmwFNIAmuSM407hAaatTqv+818zpnV2Wx/p2ZsCpOJXjDoY5+kLapjDVqVyLCmGV
2bOp7R5AU6DVIudB8wcidwIV1iP15WXs+YLgj+xhI4TS1tHRDYEwXgC9TtgHUoTpK27eoUEaj5JH
DOMgYgK1iNBe8CSlcWi3tbO8YuUG4CXh+hgkyy8qYZY79/dhVY8LytxofyUaKsTaxYazboT0EUfB
qbPuGAC+EZtUHa1H6nMapUFUcz2mwFTH007MnDwkuXjsWaDMETY3baMuFBGbcZccTEAFnlhX4xB3
CIK+MZWZhkh4akRx8C44j0L72B+ltLeW0F/ZFz8rat/Dy9kTXBiYKJEAIt9n05fo3GlvnsXEvC82
PkrPj6B3EWJSI+bYoPC4C653tMzWDD9hh6cxfynVkA9jz9MygTdTpgLscEpe1fYo01bpOML9XKAZ
QgYH5KirQTtzc7Vo/UPuh1IxXyRnDEdZLiSETkm4JH0pAW+geREBOj92lFxJy1zFYE0UPzUebF0X
LzlIuxEIKXCUA3y8DgAseDVtQHmMeF11yVD+aHDXinjOvIx3KcJka/mCaufsoAydTRVHjmmv9M0D
MWMDOawDl6iHW2lxRTJcAmyHTxGfRmk/Bpwi9e661k8q20Fh+xwdMh0KbBeJuisj2eKoMmkCBajf
PGyzlJyhX5trZO+ziahpm2jR/WpvMAIFshAi6klQEbEyvTEs2ghpaiKuTIkTJEqBOH6udSv1/eKE
r/3R8LWoehqWQCN9jNjngmTkpxSKyR+oATXx9ngBi0zu2FfBOtiU0Ss5FFXxs7XJhwNOHakDprFU
uybZ9Bn3to0ORa1UDl9vDYwTuDiUy7MLTEpo7bLPCU1Tgn0HrWVtju2zZrl2mjG7asBl+qX8vanj
/0CgqYWPSUn2bR071s0EWZ2yJcS4RUfpTZMuKBR2fFdtinWkPn/WRN7ZNrk/ArZSFp8XWMvscE5r
MxlPVGxJPo9DPIvS+H+vO98Kvp3T3arAja2AZH8Y9yIznMYMuBdp2yXzv0vFmScmUIXtjquvq2eN
VtieUgse8KTrIlB19aKkt0kWhU7Q2PVjdjIHQLKRBF1fQD3r3pDfPtGQ42HkKeuU6trqaA7Sftv1
aXD2sp77JinECN18Y4BqmwOWbUWtZlDdpWDq7FrBlhXIym52v512TwFPsgVbt03552xnlJmOEpYK
6YHYdT203rYZA9BQRi9J0VeLKyUju53+BN8onBDsBsdc/Klxbi7C8XOwksSbYURBYv4Oklcj1MU2
6j0jnZrmTHmGSJiSV0XCFzgpPO+Od1BKvQTg+Xq5d7CdAiJdLnWn3AfeoB7OFO95ve9higjCppRq
ykHROwFDga+DGdySHvLDoL9SCIszknyz+rowad4ZAnlTW3Tbt5CI91+vtzC9nN+qIe1HwVcn/sHj
DahxUqS5qpUwTH1oph4qhI+1d0+IT+35d6UbnnrCVOn5nUH0GFHO9tTSUsWqRmSVG9BMBYPHILBl
RUvgH/W1mONWmE2ebcXymeOtyDlkQOwsF1GN/loUd04dRHXY93HbxKp59FVZ/IdvArqfzXtv/15L
CrPQtpO8eY8TGjqlBk+7S6Jf8OptXYAHAJ+Vi27HQY9IOhnoo+y+BddD5HKHUlAxcNkqqEMCBzhJ
jZGjWusD9WXbTC/itzujAnDB3IvxTsJVfbHbOOislrmp/++9OSyDG0RkcQqutrv7lCcNh5wtppHv
HTqc8eFgIy3u62w19/TZIdYX8XkAYBFynif44r2dSkQPAM+PRfVoGpBkVWGygNgX27klanZhWbcb
PyRHVgE9GqFr32MMaVSiqief6Z3pzhVwpHzSpJMOm9mn+ialMczDmtg7koSpmed/1u11cNKRLlV6
tELIA7NSsMIey9JWNi9qwH7A7KsxVQcsyLePL7i1CbhAs1VZw+2USlEBkDaKMWnSZSQRz+DoaoDV
wcSgZXf+gT6cygHvXnyzUvyrcH+kVzkeEHD2ge7s0+otZRlhtVjV4AhFt9Dsk5mX5HF2aQ9urzVo
SYWbC3j2URyB1//YuCZRca9SS+rteHaW6N+tGUPkjfo5uGQSQZUNXdkSPK4l++GzHDVtuSZGLHRX
TAZBwjESryB2tOeigFRNt3QwRw8Q/lx964mM6PqNrNUGrf71lqY4OP2KAy1gkqr49PHBCiLM+4Sn
R+qYf758RraMJhrMpYy2ev6EKd1KmxfTbw9GwOfY6Kfbp+jO8gfGUipODpWyb2wT2eb4ZzvChpfQ
lK0JoVpkJRb81fMHXGDjjVeRLGU6L70M9NOGmLlo3GB1zKeFnT+rk1NMw4vm84uU+iyTFtleyf8w
ydDgYT2cjvw5ClLyfPC8z0GPGs3Dr/6arq0sRmsLf2dHr9mMms3Gtnd1243jP0pFLn8qPPGCjFuA
jlehQzcbYepjUtzcLBa71Me6uskzAygkxyOGDJd4dPbZ8zFykWNVzP5z95YEQBFK675xoDQ3iKQF
Soi5qt02o6RwbNCa0Dyovn7EJlavsNBgL/5H+l8m0vHCbbl1GB2+zLO+wG7y15C/1KHCqkje3IKJ
HpJR7BicBOD1EfrmPzJo53XBprXUYXsMhpEg3r7YvSLdQByBLA9VreVl2zNZIfLLyiVz1bAcJb2+
XXvStxVL12VNzNag7Btq1jmyu0lFMLGMIwh3fuVtLE+zH8Xel9o+Xi2OZ8e/SdSKxONcAiTxf1Nz
ogBTyfm4MQuV5eOIZAKkC5ZkNhD1apWqsuZDdEsCj7LTmJ8YBvW1h6K6fj4EKliDK0Jt4gDiXuFA
dU2WrX9gKj3wFZ05A4ydFC0BAqSzExAZPpdun2nqF+Vi1mXxlPJ4rdwctgkljzNLrEND+9BzYown
KscumqmkjnLLtF+/uaWnpzqmIJn2CWrFgl5Ptoqy8vmEMKYzyVwIk8noaAs5Dxan6+6LfphOmw2m
CCr70PrQ//Q/A54VicBnWyhkIaSf3D9T4BLn/f9gnIQbdBVXaXwKlaZxseZgDmYQinv2IC8GIH0D
jsMkltJHhJRVNOyZuObgfPQX9zRQjTHUjQKPsrzpwbkYEtYSRtJ9jgIgTuXkpet6FUB/pTbF/CT8
KLhzlpg0tMHczoT8ZmfjCRWGP5iH3bUTVriJ3skU15CFA62OmXv57Ha2CZxl6tSSJsuuX8ny6pdV
AyZFsgKK+t7A7nZmgr9GbVbxdcMsfLXfrAfcuZTJjbCql4vB+wQ/d03SM0G7ZT53mwL3I0NKZnvd
DB5RikIFflUaqwSPXWeNOnceAT7LVTB5SNpIaxKEYtSnJ03SPw7HUKtW/cjMaoLupMdJ8U5yIaVI
DG9nbpVLc4VYa+ZI9QLCbAGSo5K9xiL/DRzmMWx08LWN0TA4Mb27cHj4CrWAl42XASF1wJ6cYMk1
1cX03FgKe1EKkRtp3twzlam+und0N/x5l2Uh+ufpGPVX7rhXqTh6yxeQam0BUJfQlc3KsSXESq1I
SanNrbbJYIJiki3RlyrF+4k3wcwjzbX7+utIucbJPo4M7c4CekmOQJGNaLp8VNL6GnDzcH3kBxyP
bkNo8bsPhWEE6T8d1pXO1K75yGXHlG+KpO0cjCKHLcpVolVywtn+E3l66L4TeO7UsQvjDJ21IbIN
uy6RPpqFAKuUsaxXk/z68+QW8JfRcdVyB90Pjtp2dmBiV2Lyf+rRGsoJbdAgvhegvTPpiH1PHqHI
BcNTMO/lE1bAGRincmz2w/NtwNio8krUyWcCZb20YksuT0eEq9GkLczs5j1XllujbAwIaZDgs7kf
2C7dIGOKy9UTTHE4sUABlwO46ES/7/c7DzSrJDQt0s7tqSvEyLtY6k6wq1nMTig0GWHKw9d/nuV8
M+b7JjaCmgSOEyR03bUmfjY9j49K8uD3z+AEs5NUEclIFAiNqnz4PTQo7O+vnRyrj+IuD03Xm/3g
ObxvHkPB88UFB2eTyF6is8/LRpIcT8okQRuejaBRA+E8ZYQqp2Qh8A8MUIpE0+2NZxeQvgdZs8IA
paeNBYIAy9JHaWrrbI95ZWXrK5nCTgLpo4uVwuSJD+zYE1YK3C1UQGN+gNfq/A0XcUC10ZYSPbE8
9DJNDqR6YT/G7n+XM//sqfKjwwXNXAKZ0O47O5st86rMvztjeLirg7Ndp6oqTSI314ihk4h67p6v
nUEfhK66Jl1JYEytU29Y6HpmVmU11oOe5Ow8nb0aQlmoqQ3Kj0DUe/en6oY7hMwt/AealV4f+aex
VgnbjO4Qbyd1R0gJXcu2my3MKjJ0yWoIZytH/cllXALoqbE0szHdB+HCpM+uy0Cb4uh/3pxr91ia
Vk/g0EDf0iglV0NtQxBwcCJmaMo0Usutkyewe+ri1SlvIwIUGWZ4+geefx2n0TSnQIBA/Jw4K0Qm
TeVB7wjyZNt+5+gU6vpH9VRmpUo8z+VSDAweqekAbzy5nGr2kbskvyhTPFBWpT/Ncmx48wh7PRF4
1CDktDxW4DMYiRbUUuFYu5Upurwd82lGZhAMhh6mlj89N0D8LHaJRSfsqj14ba9CCfcm4RYffpqK
NH6k7HMdw/+vvJR65CbsiN8UhYv3ccwIGAU7HFDO9E+KUwJ8VSkfEpSQ1ltOZfGox49UcJg0KwYW
1tZiWg7ecPRJ4JGw5l8beJQTNhdDxYwDdFqzkHS0wct4m778GRQV/5RX7b1Oe/tbmpJydSjKQiOK
g5Ld9gLECjzrsqZKCijEbK5H1v43UvwqerFZW4Fo4qjs/Fy3dafto3pDb34tiesBGTA124yYasCi
e5yzRi8UnkDEis1jqrYK9UfmODmzdfApcjSKDXvgVQO2ZyoCHWCne0pr0cObA2E44FDXpRQFCFpw
lFnFhsdX0iBVMwegy13v9cHDVfss83yTsN4/6FIyj0PL9ihInqKmBgN5RnGJobIp48xDipc7xZsT
UPLk6SmJ4KlMkO1cptsxkN2g0ufWLawwUzhCsMzYe1ky+NzN8iNIoQCFBtK5ge6J6cb8xyslbIyM
tiuBW69lu30Hid1PEvNW+ZNzB6lzegoXGGKUcgNwWTxrxXxpBRqUy3Jqsv6mnRmRftT6X3k6ryho
U7tnJD4gsZHDmA1iYajyJZ1tWjT8eiaNDoDMWtFuCTq1G9sUhpJd6aD3/QnTAQwIqbf24gA0d8+Q
y2umbGEbIjrILnGg91SW34szWSZmj7sNrv9xDKEB1Dt0KTr2tHMY4JVWuUDBccLaZ0630YfJcJRF
F//2r5iGNb+03Ph2ufCu/g6lKIXFdQ9/EjUptCmkEP/vtu3ZlgYJ86C/9x1UObQtFLlVKsHhLPlN
hG7VU5ubh00xqyryD9eimMhKc8bFWaYiq9x5bIFpBvRQzTvqkMJGA6i2SzhyS3+gIUQWJNv8sFh+
kZY5NS5KNT+NGH0BJ7WoiS8LnmI52p54UG/aD2dZYBgTtG2RPkIUOI15kUVt/MAzuOXQkZP83z/Y
gvyMLZ1fCFDbhq7mfN/xuoTfmCsMbUM9JRfHffz9Y42pn+T7VJmmLLtAuy4yosp+uQqsaZrAyrHr
a+vlrn2qFzwodQf6BCjGsMoDDitDIaodH4RfVTAugbQK4fzbcY8v/g7PU7F61oJ19WkNDknAQO8X
vDRlBLlRZXt00QNDwtkrUF0QUhtmZMtFmzdLR4rn5BY2IHevAUNHyvRsfhfG1SzqG7nbZbk5V5Dh
uzQV+FTVK9ds1fHkkX8sGXvmoEIazkiT0NGegjrtF96SCef/mYbait7KaBtU73FAYSxBozZEhrEA
g0ZcxxmMyap+DmGcA3zrBnlgIDcIrghnQsaZ9QwnKU1WuemKVR3lpw9HXDF7wvWm0Uzooda1SsmA
PnMM+jxoj6nsuLQin4MRWSeOjqHMzlgbjmbe70KfNVAk9NhrsRRPQt9bRrR75+W/y4TuZaVUOd8Q
no6hsMWKTfmaamQdP4OYa9IBnUlXglWJfBVsQy00MQ/1tt5k1jwPoQXFfZKObjDfsBhpU6s5IE8n
10BmaUmYNwW9chKmEfWxSp5ww3Z1GodH6WnLvVyTuZr2vzorudnpPpWh8R0CnJ74ExVObAqu8apq
45Wz6tmMgDpiddHRnLyPYbYguddF8NSCAuBLs0TfAbnxVAp2qjEf9Q529DB0s81Q4jynX6T2ODQq
THQolOp4x8PTo5YzH9Fd74DnE2kd8IQthoCX8QkzmCCknJug6KOd+a6//B76CfiqLbzcUy62hQOE
kxDCuooeBZpdXZsVCJVaU9Dl/0p73O+T/6AuVNLxh38lsL+8HnMeGjqrNkeIh2Dob7O4FKzqjv0l
c6xzRToocEhSsJmlTQU7Us2VJFY6ydIxaWFSPo689nnVeH4Z6OQKPG9+CkFagZxmrizf17TuSVuG
vbS71hcYWCkREgrR7hgnrPSBQ4h2WRl9ZJAgqz+gKNf+dizzNMj0kt35g53t7jN4pm7moeGkM/Sg
45UpIyA25m3/VALbFRI8k6kdT+2QX8w4Va3hyw5WJnF3cNpZZDzbgVaHJOHtxiQFs2X0Mh4Avmg2
1QvOpyvTz1ympzyYUe30FKa0c721rwCZzc1QlOyvA1t8rE2VfCw28QkxCebWjcAdfjPIpjwMQabt
bq6EV1WgmLwcu7pLxVceKE/dKYMW4OjNmUU2EhxKe9K74NOG5i3MIff1x1plnpCMgt9tJmuEk9ld
js1i/JAd+Q2n8Okq9kGFroJ7X1XUTuyNxn6/cf8lc4LC2goQV7/Fj66tG+1ItOybcQuuQvik4yiw
UR4niL1ckv0Qtkji8FZqds498NOsrUsX3Ei4dCC+/er6kPP3iJm9rGoj1CNGo2C9+nSF6IqTeKVN
W/KxwqfDQMVXxLTjyAI4w6aFhF4EB4K9mHYQxpqdzweqlg0T+Pcxd15JO9BP4JPZ2VKijCjhQnr6
XV7BJycIVXPLVZhExRFSdrDjCumNsuBktbNt/u1Ks0vjYiOGQ8OX69svJbg305PnGc8usg0yb9A8
qHInPkfq22nLlZ0xpVVws+Qm/435UnTwYskrcwCAA9aPjVRVPelj2doJ+z9e5uOBez7jqgtZjFWB
1w1qvFnFbJ5fYBpdwMqzKo93s81+JbEcvEbEu9reAKS02uczMTHf+0miqDXfWLKm5VkUYRGHHfiJ
2I2ik9OiOEyv49oNHRDuoeACUrcQ6sURjIZFQQVD/ml0vqU1HHveC7DCGfhXKRtpa6XLFeOKoSRF
Jrm86SvyjkwOINs17+h6lgS2jNCqglSTgDZCYk7fxlJqiYP4AhGVzTyU2eRQ++HO72W5LDh2k9rP
K0knuZG7U4iFwQiXqnoz/32w4/rKy+4ApZT8gC3aQET5xY8iY890mCflHXzdcg48kURYyPs4JbAL
LjEHI8K2VltAV+U8x08Iq3rYZ+xuf+qFONSapo+AW8iToWgxR7pLO2l0rxKr5zm/r2sGw78BQfeH
KNHbYw2UPtANQ/d4O9Le0MdqpSwVtAIYtLQSrvDj/M3jnB0H3OrDKC6MMQplgkzbgoWKWDQdsfD0
YBbCJe8M7suiZxzyZ2CLcv5rgma/+796V9mzBMVNe7xHgSZYYicHq1GcmE1ur2eoRKtX5c61iTWl
m0ZQlbFbyGYTjjNwY32BqRzTUO9P6VKJE0PGhszU6mTZGADYTD8fNyuroIQBbo+L3vv1uVCZogC7
Lvbj8klU0S8bCD58oRUdAW7JoijZVJZuaDUhoPPCaBFfvZR+9p99tAzsUEdmoNzMOJ/8ZtrwskfP
AX2D3c4p8VvKs6coYf2TW+5YY0OL5AOeS/zOzStx/tvgOhNvvb2Gx/be++qREqWYv8RJKGBBHPvm
z03fwpyElBZtwvGaRHIgHQPYMRm/E6I4T+Ko7LJMYO1d5gXaicgBSf6JTe/6urBeN54Zi8pCekii
RTehBwAR4KazacgCAQwn52ujUPUsm6RLCy6jLaUYEJzzwOTVKGlDT7qQV4vObpclZz16QqMmmeuU
TMMA3v4kqZlS7Ax4RFvhlhQUvA8qOjDJMX+tegOZtk7GnJbqZME3fU4cILLQPbBmO6MyUy9Wsc+u
ITgXryxEIC+S7FeGdVzOA+8KLGOKhU5VpLsLTRzKuYAonIBtArWgITvAnSu9kdcEmvx0eeY+LjSU
C2HAygLqPRC1/IPLKN1ou5q+ISj49C7u6+KppplKhT+JD+nMip+3ePqp4Ae2kfz3QB+m7mQoq2vN
VtzeT4Yx8bvXZflj7HGdxBY9Nq1+UqTYWDfqRK7WNyg/rpsUmVPREb3eVVSn90nLnfQSVJjsxdlM
HrNTBGehz0zoaiNhsAqFHdQLEnGk5eIr3+5VJStWjqh4ZPo+kMQk35BpAx+b3vHCNpFsU/dh6QFH
xNms+P+kwViMWZgsGnBTDnDOVf0sn8owGHAysWcxF8OJUTR0mrteSVcbu5pvQgkfwVfFnAF2Bytg
CntqEEL77SiUDFkeeH8gMZjDTglZRrYpECveXo8yjiSX44OJxOmnt4twbJyA2fgFGJ7Uiss1Nliw
OJSCcZ3SBMVe0r4np31f4IvUqs/kGWa4pnNyYPNw08ysVy6WOVufBiqwU++W5C70NSQJJgZXc9Xd
QFrnN0cpSklVdoLj2wNyK4HWVWAbfjjLO2Q3+/9FtTTNbEaQEiYc5eb+2HpCb4qjUBEK0ASmyAe+
E5P8t3h1zk7RaWXr6S/0g1DXp0KQiSUvmWDsTbnkNbpV0UTpLNynRW+yBefTRGfyLihuVlNvxhcK
tmtmXXT3Jv1xKUiBe98/mvDwBlNxgIKy5bf3EutSXnJOiJIgBmGQlYDnvofsvlMrfle8Q2I4EUou
2Wc6xDMICAdqsdC96503msK96aCjGUACb79Ghq2YjpCYr1EMqa86n0Qj70F+ozmMF0q2kQ6lTObZ
a3Xv0KoqxDkqofGMj81T8HPfNiDuSHCeVexVS2YP8EwlyWaOewnxcPqT4Nfm6SKuLNV07GHe30aq
KExodNPt/nkbwAQIS0MsZ2Ld4WWMaOVhNzfP1lXgKunoOY3oec5wnoGT/S23agT01YDjZ8WfCxk8
PlygI2pdT7cpJk7ggw0sLH2D7+Rb+reVnb2mt/NGFcSPvaNvhY3nuAxO9WKpA0pHi/9zl1lHMxLi
B1CxcyVg8A3xZqK1G/3l+D4kaVQMolBATUxNGp9qS93tGGtycPE6pf6orFMo09UguYBnsafT664I
2S0eE2xVddIuu9EsMAPZ9eGZ64RNZHBFOrP1u3L7D9med5i19aQgw9XyRkYKTBP6ASuMkxxOIwrn
rcm/iQeh0HRPEYRBZOepDDUf+LU2U52uBV8ZnRIGtbZEXnXchJV6zNuIxw0y4qUMXg6W+yXBnmZR
ONnzGC4HoG0lpgpc7ezJ8FZJF8B+ZoqlPjkZpGUF1Ad7p36Mrjix7YBhSk4rBLCa9WFPZyy7vE+L
L0GhF86K3ONQqrzuNkv8WSc73bPClMw89kCLuDI/BbHuX6yNbYDFr1oaRxRzw155jZYkJ9t1urRE
qRrkyDkp+vW5kpKnj/yZv9G/XYGjNL787BRqXJCQTOlMnJjfBHrY+facr0slmR3Fa7ES1pxglK/H
cqlCnVy4CsZmMKZIGRhEUSrEJUG52HeRFQV1+XZOd9TSPjAxaTwMwkKkk3PAGnw5swuyAxa/9QWD
81CY2puTkNjtXlp0+2g3ojiymXcdHf7EnS1HMADRt83vuoCbqmsKiFifm1xah9QgxsqfnsdB4YkM
BqxdRd98RV2zDrxmBUz1s6SWaFRfHGbjhRkToOt+mCSv4qz1d85d7srw5gf7T3h33yXOvVGfqtf2
T0oNbXPfJurccx25VQYT/3abaE4uTnM50vEA21sTF0LJJFQ6gcfU030p1ueLJSGjNQ91P0ADa0W7
2peabcXMn+zPO8RWXyISVK/LRAJeRUfm2Xd9r3tCICIG2DSywfzm4v51RC9mAu77WrXKuRCyuZJ+
q8SoLyVMV3onogTF/fmiAOy8X/ctOK0j+H/wxolVriOzQjPjnZvztaUkrJ6uVvKmzIvfpyME4QKX
mpCk6lEnLUzvc3uyRNXcGDQw33SLvdUiYPHAWLkjYsgI469jTT/Dw7730RVj7KRwiws5z0k/GM4T
rvT/QumXKvNuxlqBD1Wcu5cNPFJNhI5BaozzCjz67dPBvXbb0/gEMpr/OOZGd3bKxRtiz+bcHQnm
zLlukOE7bQp5r5/GrlAkhgwrlTuqXC2t5dbcpK0Wvlhjv64gXGNu/25X+p/+lldk5FvzJNHVeygb
5PKA0FSC8i6tvTYrk7Asn24MuavPSeVVQRqxh20uH2jeYntdBWz4vqm+rKBSCGH2cHwFCGBQRcNy
xyV2mASoCQB6pLMpxyhtwksD2F0eaG7tFPvmIecVNSCs4hpE2xXEkEdIfWugdXoOFCGnutRqjoIN
jkSgmeM86JdpG+Uzf8Pa1DLDtpnjmtdt8NldfcsIRggrVlAT2aTR6IkaboC0II6OLgyebEC1I35N
10OHHOt5TPylIcMFqHAyDKJc/m0pppDQt49IljKKNgerVMSEHmoBhVpyQxWMOTHZhGrtTwc0TVzu
lTk8Lt38U1QO7aFeHWDfrEilBOYMAd6n1ANVjIVrRPTC6k4BoRBydGKtqP33Rvvqpa/IItA2XKmc
KJnCRQUjt+Q/qLbYmOZ/1Dfvjrak2krt3sykgd7sTIMBggfR0DEF86XHzIkVBvp5TpGcPieApvjL
5fJ2Bonm+kPpkkGyweHxLZvsYXICbcxKvoYycmqNpziZi3MN1Jf6f6QQDOSKKeZ5GUA9z4kkECCZ
xbjVfHv0K2T1fIpcUF7hUV0em4lVD2ZOxLmeM22S9Rj1uzlTpCjEJukWD1y1X7zJlv6khtT01VoF
yfBzQzFRbLt8Jzxx4tyjKxg5mEEPC4y87G7L4YQ44EEfw06xuz6Mzsu6usjM4r3mv7glyvDx1LM6
MAJ31FThAAjm6AwLk5+UinOho8/fgwvWbRJRA0+7wf3QKg3i0n4CSUhgiRk/dzrn5PD3R7im1nqW
PnGprM+KReJTyTRg/DtoDp7wS1C7ENTlR4CwBt0Ya8T4hCFMpchACX/QslT9sCiTkuYwLPmNjKJq
mTbbx7ENiSyam/V+ernFu08vtubZLoHTJqDgqx8sHrpKHVuHt5F9BUpZWFUexMmA/CmYbgWseeWn
CV1BBQZ/wWc0NruXNxgBi9nOsklGKnwEkmxIZ5f1+Y33mYJ7+eMpvRC7CMbRtvLjxqJu9/B3KhWy
X0gBvm2m2fEipVDJQZfPDjh0oVEjRpZNC1Gd4tJWajEJQHDZSG1vDVLfEZsAzglJI8ASseCqnZU3
ouZ/Dz9NFa4K5RKLcu0ArGZjSlNFWwtA5HhR/NlnZvmWTtnpCzu+mETF3VfQYvfGB8Q4Gh8z1jdU
H3KHFesjx8J+wlnDdspSnMxvzyVAHzqe8YbBi/R5tvc2vxFgs9xAZEI/fJbrGC/KXa2Es6vkji9E
u3lnv8llHGKjS5dbZdOAmXjG+1uryB4lxw7sV/VEShqMt79ddI/dRIkEut3oxuRU/+yOUdD0hK+B
Ac/t1krVILCUJwnlIcdtE013OuepbIGLFj3psC9C+V2QSkWzUEw4u6a+7XPpgdEiWOOljaHAypNn
9pvIDp+WwDuqQgwa2EIG9SryvqEfwsLKWfhBfDbfNT0z6q9JKPbTUpndn3rmLBDk8ICcux0nHvKE
HYU2Xi24EkV3zOAd8CxiggKyo7LTlWAndbVhIrPEuBDywcpsiUtjl06xn7Az6OMbtieYuNUGG32i
gA+Oi8m0kjM/YcH5uymkFTnPFZk1gzfv/z3sNkGsouwRjdBjb/kiyTo/S0KtfI88V3KT/LfIDRZb
09U9adlWA1XYC5442zXRt8xrVgo3L6frzIj7cqKCLKtS17s9hTAExv/sYpvLx3cN2BD/M2oi8AJm
KZPYsS/caw36cBVn6VrS09bFSR4PyDVM9r8qSl0o/Hjn0dgauwupA6LlV1vNlczTvKXcwBHsBda9
MZEbTQVIGNalfGEN07bctlvZuBwgXCrNCOtrJcvg2B/QfqMx8hINI15vuByavrglOLIsg2Dn7E5W
jkW8U3Q1P9BrLe3oMjAGk6aa9EB3X61iaedBOUzRSIJ2tERzizSmFEtoR6mjLrQTELGYT5VzqsnF
ldmIuyV0xSNnMqTOwWnTmm4XYpXZ+s5gH51SOmfPcM+B3JwYnHxjMWi2cJ6p9BmhfOW4jB0EpMY9
v50tmACPl7S6wm7e51YXXbuASfV15/UOMeLL8Yzj5cXDr7ogosVqtM9muL6rE3jLyguPq455eXpX
Hx4NAF1yJH9crufbQ6//TMT+dHeU5VQgHlz58IojL/yDIo/Q+G9Zva0MwZ7ZvdcIbRUXwWpefzHs
eiY0vurZE3hB04QoJdlW9BxkJD6oNIaRCo6rPmEch0Var5esrE4ybIGj4WCBemth0NbSRqzoBmcB
RzU6aIVTG8kzcNA4BavrTCsIMdn4yKHtXFCWjE0sFiVbTlH6p0XkjXFU3J7VtHcCn2GjxoQWp+6U
QJ/G5Nhn+obCELKsL1kYiKBbLhDRsAV/Ijs5g89If4fAFY9UrnnsauJdqNICcL7GXcBjBVTiKBjq
X90avi8PiqSDkmFOheUem2gZyxrXldr/p8eipZ8eJHQlBtdF9gDlQzzd/TycnWu94NfR4SK3TfsA
rAQei7CVmg3h3CNtWIwkfgqtHIN0f88uKtSpA/E7aGbaqP37tW0t5zyNKOrPQvUNkSAgwPfZ+AsX
QVWSwcbQ+nEE/9i+TJRwqKleoHek2iar3hAYkSvFgacSUA+jHNmrT7pdYyeaMnRDVigR0yazsKrk
IEh95yVLelRHvJ8sWMyYL4h4Jxm3xQ/+swZ/aDu0RAyL7F5fe3zGXVZeLqqwlnZvI9xlFGsIW0O3
Lv6mf/o9/Khynkvl9MVUrdzdwmmFmtRsin/P5YsZruIfyVYlXDuDqZUYCy1TQ4VwNbe/B24Gacft
elAWofRnATG6iuhbCD9scUsP5JVAUVjp7HsAL7izLPO+uIZmT7N12xjc+bakGhG9q/hHSthCOglW
HcwnA/WCEFNMLfnuqK6wL6iH0MJO589JSE0eq3ZnmBhyfJVLBX8yqGPBkdYkAM6U7tbuyWYx7OR+
aMNtwMraOW4O5v402MRiXZ1TsCLDIIETOJjOiGxowe42yAuX27utSK5zysO4AvmJIjhSxa75Ilf1
HIH44hoaCaNnOwmK17w2ui4ukc4oC40ddgdav63ao+Ty17OFYQN/3UVN/qLc45LY67IHZHUTxorU
nYzOWcA6h/KFJPNaAmG51HnjwlvyrbSGOOotKvPSj/6nsn9lE/AN0VI3Zd3weGpjLaJ8ztBhpZQX
S0WWy0r7t+jF8qUam35O7VAV7Ns4ZtTqoEmS9KKs/i6VViMeDS2L4gWmZFjsrqBgB12umLuyF4H/
tqKVVtIzM4Jpcwr5mgjAEXTXJz7ITqp9wCt+fzT6vgsD8KxohfW7zG9tEKreyvsE9b+skIsbOIQ9
Ws3eoRs3QzevRAJyDgNb31gZ5eTO8c0vUqx9CM6ePGFnVQrsCD1B6bWhRb3mPVBJY6RwbKUaNwfC
WQ9prISmREW4eF99i10XVBD5y/fg91sbIoJy9/df4fVBDjnh1kncKxJGZCt/fCnjJ9m3Lq3BOTNa
BZuuLWnz2Capd4Ffx1wCxsC4FG2JUdzJRpDx62qMMNCHTybLiyutbbfl6paNtm0o1ngzqHAOIOfZ
Hp4tRNII1J98SYXSbKmD9neznmCvv52vHvrQnFkm8UstiEqA+sKb9Q2sBZNB+En8pkZdoIDucjUK
3JGfiLlSJfcHDMD8Y3l9UEnE5UvaYSLBOaDO7Z3K1HGtLPdPHfiI7+ZAJEl7lU/hyJQTT42e8opO
48/pcCTz9k58J7XoD/qk2F5Ihw88xeW5U8wuCL8pJTz1XyIJ5XulWhmvsdeyg1cFqWVlGMOr9Dgm
OkS8prCx7DivC8OzEpM+9ernNy3yziFTvj1JtLAC8X8fm5SZ3yNHw9K0gUbtWZeocXy2lAUM6rAv
+qvgkWAHqh6JG6Ubigy+U563m/5EjvZQLXgaLgHG/isslmC0IOBVQ28uVmDyYunXc9qQXwFBAWbw
+90QrYTSrBzz23W6dz6nKEUhnV/wVJPsdI+EgqnZmmYkG20rSkdbeW1oRY/d+U/EuhlgGTJ109uH
Dm1r7CuHESu4ZPGR4ZAFur/SiDSEfFH9OgvEEypARVmUJm7K9ilmMHfBe4XDW3iD5mkDSqdXMkTj
++dWbCbMSZCeY8MHICu1zb8XBHgDons6N59A994m5J2D+RDceYFLAuxc9PEH7tJVw0evE2N5RNOI
xPUxSk1ua1hzTam2Dy3Z6eGvyCQT3LH9gEL3BVYTMUya/J5FCJbq0cQ/smTRbQoZRj+WJHPfI3V2
+JK+hXLu3K/Ef2jMQLD4BCj7cE1w5C/mMj25RriCJe2Pm440RpyWXP2yfuf26K+U9l5deVqUwDxe
zbHGazx8NdvpFNzz504wbSjN+PDaR10SIIjgD0m0ivflzx57YDN0P+fWMVAutbsOJoGLM4zaT1PS
XHrf04g/Icb3Zd8VqrkZg1cvwD+xGkReR8D2k1GC4YrevJvmy6lb/TeTfdIOWQ6Zxyw9E8uJMsTd
TykOrIgmHyK/IeLx5vywxy1wZFqLvJ3pdD+kaeK4T4wyXrjHT/jP5YNwxIHB47KMF9hhIPGQcyQA
LHR9IAkfL0+WeMWDkdJxqSlCAhdglyvkoa06MUP4hwvME+87c7CWlc9pey+HDOJ0mAwSfrWFjd5v
ceBNLmLsPveS/454U2oL64qXDY9Asw3S9sCPoAimM4rTfKdzxdyLHOcCz+CMKumeqOlhYDqYtCQM
DJ1I3YeJnBESOJPGDTWeNB7UM9dU1+kW/DVRd0KbavBSTS6AZitt46AXsZINtPFvekA4KaeQO5Ry
JC5hpoCSuqb0vhfmZnAJVB8p1uZV45uGtjN2wYSi51UDOIAEXQIinCCmp8lbx7Sxc2HZkcsI11hA
uQQ2R42hdFgbaszCw3O1lE943AlQTR4wSViDRTiTapi58mtNDgm786l3OYeW80k5N0UcoU2r0Cxf
oWZt4e4sSEVkguH1/pTZnryKD8WP5gcedfgQW0f/sMcPsdJ965Q3+ARWailSIY6no1KYraSEjtvv
lcibGV2ScHxP3wpxM6fuDXiWjgq9VuOUc+203CZhwIMEqcAem61RDcb/mZNhDgy6Wl2hqXYFf+19
Hp3tMKMJW+6xrM/B4O7K1FE80m8I60IHf6ATgXXev+uFaqtS2SXkfUTqfHcYRpIvHhryLNI1IV/k
RRdbyaOY77EvfuX09ZN5SVbPiE/slyVu3abMcyArvG1eWL+L6WovCeN6bLHk66hPRhYxj/1Ji8Ym
QDPWNWfZE9MShFc6QoetMR8wX1SjlKLam5PfqXj6Vq3PgTzsmnfRUK2a2RszQwbrZOqsDyD32Jtd
vMh6X0RGcHjOcTYfFysF/auPWtg2G2w/p71piDxl4mp3PO4HPHUeA6Wpng4WEVXu5LLzH7QuDkBC
Xyqk6rI6z6nO9pH0ANghRLqid6XXwScG4ryrM9eotnibRxu1ugCKZGs3NbaQ2eSvrrXKf1h5KX2K
WUfckx+7tm+epxOtqnChtKhUlo8jAefnybfUPUYY5FaIuIidQ1viLCy3Z15VE2LD4SPmTjq+ohOA
btxBrK844fe+0kVuKUD42/tOBHjEt4L3wl4XFBpW4xL0T0o7qRhND63vzHN0toc81GbakynGJDmd
3xz8O338UsxwUahoxtOOapkuKBywB38QARVsab//wB7sulg72EcFd92pwVXP4V2F/rDYJmwXGxew
o9WkPH0t8V7LDmhM6IFNRYPVCSSQuXK23zLIIOkGqAXIfcmriYKFV8CsX4oUYx5yr4PY2qxsFrLi
nWCVY7A4Vwpq8SxxPQFRmNp4wpYbSWjUo5wfO0XJ0WYKBjQvlPaU3zH9LudWM2zxEg9VnuIIj/ql
1vjzYzZF4pj1+irAfQ06MqyzlwhZFwsQjHkgo5wunjrXIGjRpYzTmeX+78CWAd1CfP30oV6AXNl4
7L9OO5fZeFoBG38ED6FLU49uh+H2V96wQ37wGmGmevVme6vLuzwjgkaobljm4wLHKC+O0nNyR+F6
0wAcigz8mKiv9ytJ8g9YBSGfIhpmXTrqcx9f45gxNtUeimof8Ie+w5+MxwBE1yOlE/Hh1sQQIjpV
AHhkogIf1BN+mZV49Fy0EKj8VEPf9prq9XiLuWZvtAQMf/WRryTxt5UBFdRfnZZlU+a8RSWczg8D
2Awkbx7onDl4i3s5j110mfxyvTGpVIbQ0MSvWVnVgOuGQuRNcZvVaf3mMBvlSpA9877L1TEVYGGB
XGMR+P9pqqgb+0msEyNPqnHo1cglpm6x4xEdj/2KyNwB13E20CuR83934t2laCplVW8hnKaUEKLX
z1gJ0FBLhnK9Y4Jszb1e0NGAR5rTNqzp8iGHVMKtcIyT1lynde+RqP4yoxAU3WaGD8rZmahBj/E6
pcUbHYHW2hyyCkNPxeI0Dp04Zbn0IqfCI8zqmCbm2bIX2bdO8Hky33RSi7UdeP+I8/wNJMLhUxlF
/skaz7X9enBcnU3r8pCm40LHFUJOYhUhaY03OMpmBJSKeDtNRX7+L6Znmn99FhfR4Uj6EVvFVsuA
Z5kimRr2I7A0sdbRwcPIE7DiHzxNRldUzUJuaClT3yENuPzepox8jPX0p/yFW7/I7U6rkwzZ3HfF
1ZfIOJjpSi0e2zjtPi53ZYaImAB7YyBIQNrOOfoJxgrajy3lgFL6oQNBa5GJ63xfTrM+1DL2nzBS
wU3P4noRSo0Br2I5ukjmCJ+jsDKVkfihB3lOWuYyd0TJFU0WTUyGSN2CMyYkukU0yftQXxmMF/Yz
h0pmXA+TVndDitzPrGyaZOdl05jausYrYT9dCj1teKNoHMwQKAnecvLIk89ns2dJO/CtWTnqaRgv
cvwmqy1TKFFfkTpPTYKkf1JUnyBUMFkV/1fg4D2trKvd1cznNmkh3xzxluWWl9dBVEM7g7GWrY/S
dsaXCn4NgCfEpwuMGUjoZg0lcduyENDsbhRnMEMoQc6ktCuerhki785Hd0EigfKd9U3A9aQSVj7J
x/E3/0+Crc4U4F2YyyJwxGevOkiBPyj5E96dSmIMjV5mmtugBLpqdSnpWGt5MH0otBogw6Ex/OiA
rfSMczEKu566V1QQiHac1/SFV2Iyx3wOBVU6Ql0SnPG5bnYghM2qWkbDObd+JGARMmrdkStiffNR
AqSCdToGwW6PYgsmwMClsELzhVg7O7xNr9E2zhXhQkM4/pwAYEg1l7B3SCPTbo24f/RFi6NHOrid
Tt0x8MlKlN/lkMfJFbRKn5dBDl24j3daeokM05TspcrMlup5nY/kPZ/MgcDjPvweNibZOwZqQCxP
eu0+dzBC6bVOGeNJNSo1pB4d6gDduL+vLAxVDNE6oLavLZ0kkAIHKBgjs9YoETRyPboiDzdB1oKd
DQovng4zObVdXbvxxwILBIarcAnlPVa2g2+rOwA2BgWs+GEJlXVS9wHzN8r35/Yvw2LJQWQMz2JC
dtEe/XctrI6CkCwJ9fqOoHQc9A2jyb5tKHGZzXKUOjNUq/RUKIQWq5h1+DrAPuDLkH6EbyQwcCSP
puoOfAVSptgy6x1pGM+OGSytxeUboGvV97PDr6jqX8G+oALvHh+BkXLR2NfHDCjdN/SoUlIM1H2y
5Rd8LFT6e40t8p6F2ULpW1+aS2C1T4QSQ7qH2RJcebt+TW44cEg47d+Sd2TMEDxTpIw8n1LciymM
Gm3hDPZLrnBnKXQq2ZuAJDvNpxV+37wHW9VbFV+DslsehxSg1EviUNrbWg+eLvRikDgvkOiwejYB
BnIgZVRi/fJzG/ce7VDyiQj7Wsg3lurnviW3lnVvopibNPhnTcHfBFC5yXOKBgDdfUZzUbUfcjRN
YmJUAQbav1tcIGrdpupKnQ/LnvAnVVyRhc0Ebqc/jxIQwtwAjKiOEp/8cu9S6KlMP+b4WLItKBw/
VN2SbnVRn7guPG+sxd8MIpS7QgxYGvBefpLUaFWUNzLgMxaVMCl5hJ4/PBh4xQHVlI9oZaBxGHYE
kLANEtD7gHd3E67H4PI9qXH2UxRj3A8RqHQjSmB+pUPld5n10I1OcUiRzFCkb3NK7wl2JnxYTgWQ
PonoEmc+zHavlyeRYioFzNcDhtoB9LDM6hzLxpirguvO6X7Yh4i3PM884XzikwkykcUpNFAx7+Ko
049AVQN7bx/Huv7TxtNNh8eq7LO7afR4wIkCzhVqZmnAK7xoVX5NGRxbIEvlXggJWbdfRuzu/iBF
F/4MobyFRfmRNUVAt3ukgOlm0Err+m50Q9P/eZTlULEbqM0jv0Vs1cAsTagAFeszIDkFPEisMPv1
P3WvZftYpltFCiytk/O1OoRqG3MTYstySbqce7twaWIO0GzI4vmhg1TmmZU94cUFpSXh45uFO7X1
JbISqaoKKYHCeP5Gz1TkII/H/9fQcAV1+5AHa1/20+Kn9hEXgh38jNDu+BekffSi+TJLt2JOIFeB
JW1rR9DL7hLMXbFpjtpaL/KlAL3lmdc91PmBfEl8VvfaUsafO7rMZJyQV6uqwM6Ag87eB7oUG7gL
DrRauss/mbH9KgjzgraBH8GvIWTiVOvtVDeoBOLigg2zQMQDpXk1nraa42g3UgqIo91NbNICgOMi
AhFEWLGBvgVRmmxO/mTi/LS5T94rxyfycv0VTYW9QFnDkmTyQARi31aCsFzFWORovhpPXA7ACaL9
PtvH87+GG4HaFhcZCjf4AoL4jPysX/57No2jU7wWnYWYJSCki2cqPtFW5o/gC7kKtb8hC1V+Hc4T
Iyk3sLxqdZxNqZe86cM3OkC7ECAxS6f4trAvyD3/MZEQ/CSnGgEpHHir/BanMt/n1cKz2hwIzNnS
OjNi0o3TjZf2IwnZWdxFi7k1bqpac/++q3OEu3720Z9qst0jN210HGkWHBROQV3MkzTX6wA5lhyZ
lzqF7YEF+C8iPJu57difw65zRAzOfMUFrzMIOK7fu/kBstzfvofmqAw706pgm8cPCKvechvwT7KT
G/KMGa63++f1dJyn2IsqfG/ae950Wp/fzxbghlGfXRCPBhK/NcMJzJARtu7MDzQPbfcaKc4Z+uvW
tck+ATGCu/MJ3S7m+wuY6wzOasABJHadj/ifa8uMKtKiHBcUuh2w2D+u6PcMUeY8/+SU01NIrgOI
0pyG77E6+FgfLwkW/z47umPo4wnHFUj1DyA0zGrJPxTs1MsF28H+W2WjGITDt4FEPe7jcDNWi+LR
qmL+2eOrE3DVXyPXh8pVsCSXyDiZcZT0EbmQTLaM9sv0NndxGg64yKw4I7SA/InjUBQ37Xe4AnEt
O3Iq+0sFw60KpT5BOsH05fzgzRbK8K1rCnBFgubz6v9YBpN2ar6U9a7YAaknoATMy1wjGOngnWZg
380DRwxolhvfxggUyh3Ac7fXp62rxdjetAH1NnBjFscg8S02Z7iOi54MhGAo2wc8Ybum6iB/R0/P
YJB9/xrCUa3nCH/AFzpklWgdQJCQPpmoEsxz/NEe2vtkfQ0BU6ke+iZE1L3B1A3pak/GrJrE65Su
U4ATdN3EiCl/cQwgDOi4zN2OFFk888uucsZMIvyjgS0DI3Ix/Y0n8tZ/Y2uO4gu0zdoK10EpkwJA
Fi4cgv1KFJ7SmL1dEzlv8h2ihpAHB2JYWfs8Vi4jlDQSyLV9pLs2B+MGsIFkOZZmdiEIiyMjKv06
s51+t8Xp+K/qChH1W3kF1ViFlTZBFdnK/3CMQWhBMmN57k7sy9q6TYDjnI6R/SarhcZnbH6Jfj2w
ouowK2dLmdIShzaB7Us7rpqHLq1HJEkJlxcaLCzk1GzyZVXXSgc0ZdYYUvlWGSYceJZXO6frsZhb
SrCRSiADKjeD5ANqisPhOhAKBCc09P2ACbFsuhnleQIFkjdCd86Dp4kbQyIxva0QkDObY/5iUqC7
rQybPJY6pa+deDDWfahH0FN9kQpbgZxREVcuxhtM1tSleL3qLtcX+jScrFXYQ0Y3FHf91Fszeb5V
NlrqHx7Xl/wXAHhg36EVnSyN56d+EAsMHTJCDReFMZMRG/ZXLWaEcxb7NfwKNQM7IlFOaGj7zzeN
LIl0yyMmiLqN8pga8qKnlYr0R//mHDk83BLBYmCFjP0XCFYp+kubH5rauAV8Ag3c7CHxxT3nT8gu
j4FEFiQ4+9PuyUwoHJM1RQuxhxAvzGwHqWogCLHkckUQRUxztGCLiffOIrCRqSAdYGw9pUCqpcNH
6nwF5nMhYV3o33nYweoir96xbpArF3meQGqxLjkau/C99IJxzsFW9yVoLuPU44EeV8DvcYtmXEqL
akojhe00PYYNFpnCfAG8y9elZVilTw3ImuZ8Ns+StSn8MoEod+z6CyXZ1uExqyQKebOPSYJfgpuI
9aRGUtFZYBI8G5iFke1+j9AZG+9KcXDGpLSOgl3OhJyOkTLe9U9Kw9iJZDaLefScB65o3+AW9BU+
ilpA/z8ni4ThXHlUEUmiLQ9QXIYIgJpVJud5fkNhfDwOILSTasT26pGEKkLwJw1du5p7Zp9ImxA8
0yvfx6vvSBVwNqPHEUuHvUnqcpFCPX22qPinnIufWleJo446YuankJ4AIzAeT3054tKI0jhrk7E2
BC+71jgjUePdGyW4qJ9PpmFtBkHIKCpdOa4NClrIwdFsFlG7giFOVI87PWx3ipQoROVN3byur2Ve
ntuWfiuSD8oIdESRl7qgxloPSZ/z7QKp9RA6mRIxv67A0TLS+k5MUiEWerGwfQow2KlfqAsZnSE5
lOPRjubRWsuKxh9KD/VEVX2F+W/FdJl09MPul8ipkvfqfeCcyClL6xaybfRYzMbWsXA/Po4yXWcD
/y+a4OSUERLOQEFibzcgrdun3kguWBVMTAZD1aC+pIoKxRv7r+BXBW5IzN2HNqzwssUeOZ5WxLrc
VTQ9FztBguam2jAwfpYqm1CMMFbFI+s+LyHq/BgHdDo2QlrScmc6oaja5ueaEILmM5eb5nYNLkj5
O4Y8cmNqcAKW4i8BYNnM3QI0fiCwqqfunVSURlhNSeCdMBMrXXcMbgCV8e8Ks8sQIcr2V7S6cyyz
imsu/iczg9njGIguCMusHMzV1ZBylOYDD9OQqDVkaDzQWq3nBViH3yqSNqxlQNkQdwxuw6AlPzaR
sX6C9l3NHOquzqiJVQS4VDnTb3L+MBdmMwHQbvw0QrRFlm7hH2HoLywBk8pcBZz9nWwOfhPQRLHg
v6FgQND5MizlGHyuQV+9pGfEPci76oObABSVAiifnOUbsM0E+jVuhuif25gHJexfbTwQfmqLX+OC
qoUBWx4bIZBhnvVzf0ZW3iJzGeThkQ7D8CYja6190Z9pt1NXqX0zfFiq43lfqH88JaK11LxsWVkQ
hsAuZJR1wc1Nchs4nTlJa/ZTDfBYgWbF0CNdslBBzA67i8BW9FPo+MIDzIOlECjYVWYVu0+MoV3U
V4ZDyj1cwWVHsvB7qpDtUbc7DrgLAvm3HsfcizuudUWRP+3tu0sFiBFsLLJG2M9bfUjJBwskmYK/
P1OOaNU11eF+0JAzhrDILzt/F5TR5bD/Y6HeMp9R/mhXKkAtiSzw6EufMYfvDBVLMHRMt7G7r9ty
p58NuS+yieMIJ5/8JcOItEsGmVE7cheHhz90cE57A20caXNJo45tbRwscrViI4PPbNNilSUX2cgs
In5S3627etZnQrn+9R1hiiS9awQX+7vmS2prRC0br6g6F8DPsj0Skpkhge+oy/GgzJE0tZ2Y91lF
VgiLnQ/xS/t9nI5uoyZ2dJdCItD+G2rkniJ3obVb3Jwr6n+MJScA4mOy5ayTWKpPha8rMxbvbd4r
sRqSboksEA7YFaF0UQAvv6XsMCc/u7+/iLFA66z4ZmFxltqfLvshrrtQ6vJb0/FR+9HdHNX9d+Wk
CS4iPxX3rfkLabOqx9I959+Mmvf2n3OzbrDpq+Jb9B7ClIx577V5mwWjw61A43PHZQ/yMnQ3pOhR
grry8UYzx4v+YsoftCKLJkmgDq4oRSJiHA8J/1YZ+3Uj2w41gganL3ZYplMhQDXmwiC9Gw9GDKVx
L6JGUzHrsOlPpCSQKkMnv0WP5xhL1fTEt8twN3/zHksUR+9kWdCilDEos5LGe1T/Y82FOySkdOwe
f27n+6wkFpb6JN2buejA+L0jNw8yLqlfuuFRKR1JapEr9Aol+kcg53532Jq+i3GMovV6vkTlV6Y6
fgVOyntivKGFyZRMUeQTUYaM2zEw9NdkmcwvVEnxCHYhbpIXfhxxPhFDsCsh9qHDF0DzHwdVqHur
FuyNfQGz8spDLDH9h6hiFiFSe+8NHj8ffkh3R8T0YhCzVu6CvdyGoJstHqWsBUk8qYsBgRjLNexw
ytg6U1Jv0b0bb1MfXWsH5lXoTnb3pE84WSb8FRO7cOrYG1m3+MkbbNEbKN5ZKx2V2fvnGKg/GOh/
o5lTIx/tO1fEk1xoqc86q/oRWrnWcG2pwWgkzKTjdxhg5RBjUua5ai+uv+ie8eEIsD/ue7mwI96r
tR+I3T7lJLAVGmlPAyAykvW3X1wqjtiANh0udO4zjB2mTIgryJJJsWhmZ4L/8prigo38x1CNrwgo
NidZ1IwDjXGvopPw0SqYLDRMNMfQvM5yIqCcnV5KgWB1SbDlqwB/n6zyD6dgH6m+NYxGBjuMQsxc
8eiZCfz9BvUGqnv7QPrKUq/dk3OxMVrAP0RRMAYxNx6SFYtnDkfJJUneFdS8nCqGaYCja/tehgXX
bAjCgbn/ka9995CIhqgAMs3fxnpJniY0oKK2/aro39FYCZspwp16g0z4f7sIghe6CHdXgKmFHiz2
3rAHCDRA4WiizJR/Nzkz06DsFXKVpvBJU+T1bJUST+wWvsSfsDe3Gza5KkkzA0HW3MZnL6Wta7P2
gh07DEEpiS4I4ErKhhZKN/UQ2IJY3udejun0NHNfGBtSmInONA2gPqNHXEhN8ddjKmm/vuuu0wH8
qU4cYnTsq4rpJmOQDNWkNFpKlnih+1JpyYilOilo/QTBRyBSknCqTxR1eAbSwjfxo89cCuBWhPrf
9cWro77SNDBevnUoCDM2EnRsuB3obZCDOF8T1AGxzP5ONw2kAB8XoUr29eY+kl5UkL8GYmQi5sMH
Nbxy8T7VAXkuE+jbcsJoLwq8Tx5mvhfOa5eXlwcHZrjDx8t6mldO8/4CzqA1O/UiYsqbeSQwTXVl
HPRF5zl+f1gKD4XCSRYssJNP+JMefk0HHbmC24Bh6lsYolOUJPMzKC3VYpAmtkkMqvls/m8A1jdP
gCm3EWtUG4Xq+Ge5mYe3iIuXsfAEBL+H6ChOwEGaUK4zjRYNWnnaD7srhOheTfbokUlY6Yqqgiww
PbwJSCi0YLX1sB40H1cH8jQPIGXzIPxdNbRkSLIQ5JvuPuG02gVMzWpWJdu0P12vCIPoOi7KwbqR
cwviK7J8zOWnVJ/N1QaJy6JvxtSUPiuRZ9bZXd28wVtWPbZGBq9KFyEjOjD+fSWLLTOujsT0u7m6
5YpJJD3x89gAkApJVeIPI1B+KfmCOl02/BaYQQ2QsMS87PPsYdvcQ2Y8WIpvnv7pj8/c9TZRC9BO
6LK9M47US+zq+xop8pxT/KBf+5MLOHRBDsoyL02hWb1Kb0UR5SgzLXKMbjlz/jlDZTr+eFc9ZnQ7
mE6v8mt0K0yQ99PSOfSRtStvvlV2nGVU8MdY20s2BHAJdTUEy2por9NMZxZPj6df/7+bczOwEQyx
bYG06p4zBRA/GSnmDDJSOa0sS+k9YlmWGZ5GGRWIqm1OgugwGGMqNt0wD1gCAVsUnzJQOJIMeCwr
r8K9QQKpAl2/nQ9b3XOqEz0J6JjbBIxqiCbsNkf4+RT2ih/uq/XLDHCVL4lOd2Fu+gvm8kFnPikb
VGryHDopocwf/io/x+m0S5eQ1sajgbuvXv7o1ska2eRNml5VdpZqmnQrT6pLimg0E+WTLdNoUQg0
GeChqkrI/H1+Z7Di8B50C7S+tLj3AMXcgXr10bpBJQtolj+yz65wWILOSQlpGnOnf+5BpTxwl1Ph
kNYL2B4GrXJ8V4Cq76QacjgSpwwNDZrA0dk48r+NZgpsDrUKQHILVy85BEXscIrDCD3O7qXl3X46
cNTsl1LX/mga+hFv8DAh+59HDQm4m+x1vShx3zZwYYAeqQNROLhZlnGhSYrbD/uurTlyDl+vUiVc
gDA02NcZSWzgvyElXItesUnWXrxGtNH3YvyoMtMa8TWDo2z/tdwNaBiKCQjxoWbOTvi9i6tXoqIY
5/cedClfMM/nD/seKzzoE3L9zEToaO13kXhF2vGJ8/NkL01x1xE1vUmAipOJSw00h8BcMe8RHwRa
NCbU8WIMBtqUg2wwX/H5R092/NVcOa1vVC0rNCmJDV+N/lORj98HSYstImIoLLvL857u8wJrkcNn
3Oc7Aatg1VoAiclpxD8DT0Z9F5BnpdFfKz0H/McBMnobwGt91I/yPV93Az/PnuhQj+uukKAkHAGU
m8JQpmLiNGkbCJFfqe4lA+AAnxSrJ2bdTmP2Es5ErcI2FU0CTaaAKR2VpXuRpSWJJst9yY2jM1Yn
7KV2v9y8WdvTQKXrf8l1rj4vlR6O1xBEwws7KLB+tWtTGxfR7t202eHN/rwvl4rKlefVmnLe1Kgl
pFzn85ob/es1dNWj2l2fce/DesqBZ872fC2Uz8WTobSCASaZ7YIXdxHfhk6/rYIhj4Rk1STFb9Aq
h0O0fXDAAWd+EE0HKD3F/l+N+T64rydA8N7aJJSmzEBZAVJJoz+djXMq5DeUoqmyEcxYSZ9vNpuL
GPHEOjLaMV6Oymn+i5ADP+8QEd6E/qN16FNQeO8zTph2em8jXUsSR5r5MYOCMYISj7VUsrgQCDTw
G2Byq0/P73Sbjh7X8RudipI21fd6yDAE8VLqv7QYfyOpcvaQqXnrmm7vwRv3ixh4DCDiZpG4EELA
i8gnoNUaZLF4Y2YLjvZoO+sZWipjFS1erAs7TjxqDFf6dZX8LIBT6MfQ1MPE7wdPIx6S6lAfG13V
ZPTC9ZN2eyLQkv4iTELp2kvM6iFph8ak42+DVUxfarTyjusUgsEGaB1S4W2k0S+15n+0S6FqFEvT
pM0r5zYg2CBkCPrKxCd/g8Us1rq6T1NIns9Mxc4mmuNUMS0BKMIF1vJSAZXgUtwMzs9iQMx2gKX7
bbVOkvi4dKDOJKFYFxqPvS3vA9gjp9YAvHySB6I19OgOswv54lPFUie/JIL/I2sAJ+o1iWtDq6Xe
DnKZJU5kUIKtLC9DtO1J3cipO9h/VVYuTGP9+x9n3OKY25O/8EOvo2T1gQHo01LydZlCPvNUGloD
/Ry/ZOrQbO8oBFw/uaPMYMT9sQ5bDxk5nIKobmj3frPk9ZyU5t9ADgnSwAWEp8JTqYUCA9dGyFdq
qUx9Qiz7hSecwYKGhAbA/PeK2Hl6tquAWcVzrDT7q+5Iq88UdSn1rbrQGCW9Ko1M/toZ71FeOPor
VnddacdrPYlBtB5/7/jxDdfc4O0tBxbTzjIEfFaFMp1VUWB+PxEQXDLwSEULzfJg885PwW5jVwJW
cP2SEiKhP2RUzFVp3cwcFoqoj5U5c8DH1ma22dgHaFhmQXreepjn1r02hejHShTReOLuPGOVrWz8
MSaXmGAkJJYT3PY9BZmiy/jW7uTreFq/JzFyd8Wijez13VmasvRAEv2lAGaeed+jl1eNz/sNhPMV
j20ybWr27ALazuhbSf/c4bt/fCBAPWTWrPwix3oByemzN+3lcy78rpsBF6MYjTazbZnd/gBRKvTI
DTEWxPz/WjvYxs2BX3FSohYclJwcGmXHarOLxf0WTjRt236atGpYMaLnbzRuBRXLgHqmqdjz0NRV
CEk0iW3/iCJtNiEgR1SPHgTMHLokrwtty5CjifetdSTia3PkM+DzDiXMkT2TwhU34JviTwyj0F5T
xLcGz9VTdnE8z65EieNnpdMjGV/Fz8PQAposusfdP9fKxlL7coE7gjdrbDhbrQMRVm0JpVDQKEuF
SzVF+bFNeY0xPcj2f6MHCN0FPXklwMFZFxZZ28yt1vhWR6aPHFmIsge+twcE5yWLLJ569c2z1nLn
rJ7ujmatQDu4Fr96HDkjJp0R1Zi9gqJX5jX9BJ3/r4BeqCJssjJ8mBvGbegpXj+diYxbHhX5HdSz
OyuvWqE6L0+yH9Wx4167EyAQIa7tTog4icYyLB4rhtUPhV92BrBg2QmiuOKlHEJ8/LDCQF6fjQPy
IEKXtycFEGAJTs8+1sG0TDtSreGnnA7lVGcOjxMs/lrdS20TutcplmYLJbldSFv3JNZMFg45Cn3K
dJRf68qGy+kfvmhqT+yBJlKw+hDZSU82rFixNrPtwTJ9WRJsbNLu/+QWHNOmVuoVNE3V/Y6w+3wm
ynqYOG4mJN+X8m72HwTu0nhWJpoprbhZqnuxsFJXH94B/p3pMyqmegki8sPBCIycm4xFkcwyssXx
32MgjiZU/C59m5mQ4zpr+O15J4mYAsdiAIvQz5AvgLoTKWqw5FCqP0mzfn8tbqhaAqX3kQ/Sk4ZA
Ueytbq88Btt7c5/EF9iXetSozP88CMkIxM/73gWLoBjbktQOz1U07VfX7uxdA1MSIXVMEjlTD9pq
3rPL0YyBDPeXBVCkEqBxhg1snO/GRKDPzAYWNcnsz489/sCs2i2eC6nEf4GzXcf69tnSlB/UjJIj
BctmZT/nJXxH5Zhe8kNg6Xv/Uen6Wv433X19qjZKsrp/8g+Jkb06F06CWqNU+JDQcyA7txUYWy9y
/lD8p8uOOezC1Q3SO32fsqLCZ226g/pkewqkz4lr/IZYgj+Xk4Tg24+Zgp3cuzBSkjtj6CkU/FZK
psGZo61NJqd8nuptRDWq99vM6W+/xfbkX3G2hJn8Yu6iygn79Qly0toR0cK3ite/LWwhTumdq5qN
2G5D+4VcnIfvMz2UIudS9wfexaeClov4Cf5UAUhRo/NmzAMsWkWn9k7zdL6AwOzQkMt8513u8wAx
hietdhvuDtTpiNhutHV2SYTcaESj8+gJk45wU/eWoQN4hQjI5x+v2z0oLkHE+yLr9knqUV08qj3o
1IYc7habsVLLqqRF+7bKsxCKq4UFlveKLN7vDvMeQ/TtoDCS4iWEfFRKPsrhgUjQCiinas4DTKXu
DYoPdF3sSJcWWLlX2EcAn3xIAF5GV0qh7WrD39pjSt9NJrXVh2zY8ZdLpI8P+y9WAXuC/zAIIb+L
xm6eT4DuypA3uwETaxCpACHcvDYZBH48PivysnWw6yMTae3Z8IRlDVbInIRHzpnyiCgUGeAVgoon
C5ISAPXcfKaT5VxQ6hWdQP4fG50VHPzGz4k8AeKzoC6lChnkH/9xvNghFT4DPoKsB/62KiAbZza0
+5+3ZmnvPsg+rlV5rRCY0FHMMmoeYR8xKz21cXpnU90ikXjysi/gDDCMcjvM9iO2UVl6xvRpXPfl
xNF8dZSv3MN7mlyBPdZG+jyrxE6og1nTyBNSr8i+tWdgxd4PMkAWza/HoRu4u4uElNvgXTlgfH4m
hVCz4AUPxxLwj/vPZHeeD6fyh0LVGNAe4VoHRmYFT7XMn2QhNEOUMs5KP4kfpJ8FK6sATi2VtiHA
7s6WFB7BhEuTbRBJvJKdN7h8MvMBoCNGVlqFuPpjgZPX31aBd4yt4HnBFPquCxkAHDcWUEb2AgOf
a03v6oKVYmPp7Wn7AiDwx+5FopYzK9OYSQJjvaDMomYVHU+DiFsfowMw7VN2792NSN0ufuSme2kL
hk8wvOLlytdC/U1RW1KLI6s4pP+EZaKYgc9+zamhkO7KbqEpxa7ogHlTDR2NkhvBeKYnA+ahMj0X
N2XLKf3xM+F9ZmFFZpS6wLyQzVaRfG7QE3CM2E4YW0vp3wElZb7+ZGVxLd9rKaUvegQGDmLBJTYR
EpBzTImBd3D1kKz7knuPvHlHoXXZ1/qXd2OkeRvRcHg3xEtlcxY5I4sVspjrOdOZGQtdT0Dt7Jzi
HCt13v9M4/rcaB1lZjIBMfHF8Lu3N6wOlvgufiItVcTEIVGNn7OPMCKdGh62sNYphXOLuEMVhXeC
FOq+gwwCkgdfqwIrjeBdR7SC2teA++wbIwENmbIncqR7ozeCc5XBxvOcMcKUAf+qEz3z6eOrO+fx
wsQYSvlCcMov5Bpr6Rvw+Xsd41tQ9l4Mq6HQKwLCUKA/jUXriBYGX8ECCVPNJYFZbzX+8MZfWBaG
5NjSA4ayh1gNaCKgXdKPGXC4+nsGb7h75fzhk/rwX5ppiQ5GW7N4xjeaJWOlRVBThqGl3hIDg9Rb
jegSXCK2szRIepdVWu5YeP57ZUEqoRu2hrOLvTUgNcDLZUUq1qjOseWO6YliNme6iXO2TylDw7Op
JLH4t5G9QgFxGBBB+xbtjPg4BZbAPjjGmFDaItQ8xVNB61lADQUfICVAEnHsvzfuxeZAUnghAm6D
U7ax5un3MOSeRKV8dgbyxnFXgytcEc87G9fFn5jBkeHxmg77cwEQpUD6YKD2B9UBIhHJq1IZSIq5
flMoJ1Yzishhrv/yIA+i+chlsxWj5kkfgLaVI1a/Ht4RJ6cT8hPvTwcaGwceeBr74+BHa9UEuYI/
vhmbTiR36NhMP5nvftAlR3yROb5V1cKP7ifY6Fr4v8pGWW+YQhuIZeaVhWXiYKEeYk4bypDzkZc4
OUp2iEn2drkyELDc9OB0YEj8VHhXk8PPGNFrSJ7u+ybjY8/pb3iIqovU/k73MTpJWfrV8TZr9QbO
EwBqGutBirNWesQCu1e0yHPUiB1tUnDIVzzMxsrDJ9HOxvz2poniPZesuY0X/gy7razThvgsc9sW
bZqDhTPRTDI3BB/ceAiqRkfjiDH0EIR/8tCxj+61AQ6EGtX/TshT9+jWe2JelxZjNNOLOzzK2cFt
FXREcrKa2EnLc0/zgtSae2EuVLZQhz/mLboIs7COAXdN6BFr0Ry1j4ACMQkg9BXs+LyrtPOftGsa
YV/y3t6LMnO4SWmLo0J0iuBPWxfPj9X8XsLjTgW81A4uhwT98J+rjHsgtCuT4DoL9kgzFUSKzfJU
KP9YGq2ukBqO1q0/yJ3pMROnvBYzX0yHJH5ZwNh3khWhqvyah+ONKhksBT/BFhO4M4k4NLdaaUM9
sHVfKt0GqGRif8A5seBlzYC8OggXBovY5SgPbhto8SR0vxepHXyIM8eCeSQ7SKn23bi11hEkTRRP
Qd/KClCEKvUFlofRdOIXCWg7T6atDpm862QgVOzFu/SdDxVJv886VmwlmzzVJbVqvLir733J/1Px
GdJWE+A+ppQzwOz+tuXSuNRThGSe+8axoMxxUE0tZ1L1Y0jmPWSQrdD0pmzJ7vhuF0hliKd6oyJG
yppWOqMgRIDINczb1JpvrCegbhfMSzVljbjw2rwqVEkj3Lal6UWQj6HmYtsoj/1Ouiuya+0OmQUY
IJZHVNcSy0BN2eahaMtGp37xRIAkuZJiwLn+g8USUM7XYIQTa1VEE0jGTiiOjdrP1NpL58UyoR+C
nz7fuSU4cjIECI1xnTKITNc2V42EFCjyD8QtUL28j1SyvtD0RdMmE01K5GF1XdYF3DaiR0bnXPE8
D8gv18VwhGDuQGYlPRySr5f3PZ9ArbBzZ4nUYRpQwGYkQ8iQ+Yz0yaS36b65oaQGrRd9FzfKW+eZ
C5f2+AIITUOcIwKwa+/qDVSJ9Dxoqk1EDK4SPYXJwyzWYAzaSHSJvkq47+CAoZwUByfqqknmdske
jGO16BWdTG9HsBaR3gZ/wKvLuNJF+Kve8zZyhc+9ww8cCDdm+GX/7uy32Xdxak47sFav+yJbbIJZ
N+9uwzl4qIOknhJOpRGIwQa7PvO5A92xnxfTIEf7qnf0uQD9FPPTK1V7QZz6eGKsOwn78nCwOXkS
324bJ7l6/1cvYqwSYFC3GqsT3KeHWc5e7V0k7gMV3RGxGrZGgZM8bu0dfbKuvb73MSRzhAgGo5cV
gBp3xv3vsGWRmOxjAoDOuxbNw3kF+CC1MLwWBje/TrWqNHPQrEq7lsUfN5NFBcr5sRdzcf9O+eZV
383wQmvUCeMWCZX2aDSZKZZuz987TZenOf6kL8Xmn/5u1Xu0dOO/S1CkpJNtnDc0ctr6FtEZN+4A
IoweIdqblOIWlOSeaZ/quouNZ+6BE/OnVu1+nevs/7PnC8nf5w8Z2+gwm5S+ElyAcWDSSZwGgz6W
qGWZhDjk4XNoOe4G14/XPjrdevU/4SZmjxOka/CNNd3Klr4vizfs1rer83qPyQliVqzJdPVd3OIw
GlpgWNaPTVXj75aBJaiQPIlBAA7ALS4EvMVzaOEZi9YKuJUn9ecTpqcXvVHOnQpRLifU3zk40jYz
ClVOqqcTCMUJwdSX8idn5hXv4tr9FSpngoegV5/IMz6YdWkwD7AmqKIo8kzOok4Dg31TyCtw5P49
JxBi7te044ZFsOF216kNqoI7bmimahDoWRcIjnNifbuPCyGmurXfkZWc/4M1MwmVNsNcKIZf/zie
3GCuDdqphRMYEsWlTZFyV2S8CKlwNiketDONauaW4f6POi/gtFAxNjs3DUBjCraCLyofpWVbE7Gc
xhuht4H/VlIfUsGX2kzb7Al/OmOsMQR5IWtijFhprY3hKIvIsJDDHECFWqg7JGOVBPDAouicNOOq
OkgPXdgofm+1pgKDT8lL94qr47BtuMVJv2WKb5cf5Dm3y5qQGY7tyIKtg02j4IY+/ZD3OiBgKety
Y4AXMayltdNnpJphtP5uKEkMLQkYJgpSq9KL2tgFRjfbHhvSNbokbNdDzHVzrM6yV10RtJnelxsI
bYFnC5RX9O8mGZgfjAWFHFG0hej6yvnd81bAdgfYd+xsBZgp+ruvpzUiKAaT3StIwHClg4ZypsO5
5Pzkwsa6CWGK5vHD8EpJhwogtr+b2nkErnCk5kNA+w4ynQRS6RPBYP+kXBKw4l3lYN+AAqIGH26Q
5eWPTc3g7nyL7fg2R9XL2jSyrSGlDLHoXDyXuI7h5fQ6OHAHntJ1KliInwbxYvflgpS+J0lMB2DB
WjmlAiMPkZ0WC7aYPAwuIPnCqG9AI5tc0gM311bJcpJ+SGz8uDyMvObVUvZcGHa6bwEZgLU8JhoF
chi9U8VNW8ScmgW0AXvBGziKxIVVwKel5TAHV5mp4+IqRB2ZXfE/Kew//+teyxPfsnc0a48AfgAC
9RsoQi3xPNDCuUT3oxIei8lAw6nazFgRJAACtMEzUsZ5QND0cghlxBvpVLYPCSkKImmi/sB1OuQf
FXwiSCi0C0km+ktDXiX9WQJB5ky6ulb/0ZqlNUXiopTLLBsACws4n1YPuv7ohfhIkOJ3rabptSGX
BH5QIMgge+lSTkeauE87UxhREGsuvpT1yR3kEpQGh1R0gFcOC4ZPZxaP3kSaYye3A0XQKBjQU3TX
c036r36eMKmqsZIMXsoJdDuwKDrD6agSCs5YGQlLttobUrJRHexpuQk5UKPLX7jWefJsc6N3sHgz
7k3IIcDZqnISQfpBwRrjaWeZiMpAm5SZ1Hz9iS1fhR8iEI2EgcY/T6DmMcuXxHy/pEa9LtmYbckB
uF6gnaFiZJLibTDFB4MGoDpAe9aIIodxtArvEt7CRWLkWbB8wnF/7KBGhUEQbAqS42kylSK5DoyJ
YUEmG5OAaBg+G59lZTqru37a1CyI9dmAn3mag9aTBT7XtWe1xVRDUB+xegGXvQjqFF3eLLJqj5EM
CqIAbohrgp4twDQIvvoe64f7L8L6KYFydhShgwk30dOujrnLXj8jINNdgaoCi3362PCGqeUOIaEx
lpMDLY6MoeHmFuJFuBsDFl7JuYc0OrzOv05T7/lV+aJZcyKtvTnp6kVEaDuFBsGew6mvWXqhiLkw
b7n5T1wLe3+DLGrGBa6S6XlDg5zPSuYmVi8I/RRCxC1YD3WShUWy0aSy6aFX/HaeM+GJ0X5suoKz
CHvne2pCV5v/Aw3/B6rBDQDYQvFwq6PiFFW2tfyPtoM1Q4VyefwCChlKPGPwycmmPNjyKgtoE05Y
tYyXURHTLci/+C6Q5I3fhWCoicrW4GPhNWXdKO8YZ8cpJ+QHaKboEK7CMKnqks3HSA9lPKrNLChb
zn+lfs3sRnhKgDkUQouWQl11eNxZNBXncFvuXdUN9wnzZ2T0mIvWUL7o0xn9JT1d9KpbURbzTxYo
/ixTLrw2PgnjDTnFLGs+o1ceZ5k4KceI0aawZt2MYnRbZUTbZbyey/K1a2BClm1h+pjwyIby5O/7
hLntlPgRRCbxxkAiFS2baSKHS61XAKdB+x+alWjDt0WP+QSsmuJBJxVoFFEWNJyz+b1I5I1AeJs2
mlUCjzL6AppVDyB1GWmZqqtlG5aBxQXinHae8/qVSi4y24yQwmf8spywfyuqF7XxcwYDW6DP0VgC
pl/jHK8HkW26uti3DG4sOmhMUTPSTgsZJX3zZxIDPc4XSHh2b6hBn+iMaRN3jHAB3CzaOBB3pIZ4
vvk/HMAmWZeiba0Egaz/Z6vCukucHKCtV/52m0IDXwSPOfQJV1eSHnyoT61A7tGP2C6cY6Zv/YSV
ie2QosFkt3+VC5BipX9nehIaAXsfMu4yqE4kYt4f/KEcMVsYOmAFUlJ3GO929BiTFIiZ6lt44+cE
pI56c+3LZwNRDqDlw6zHhAfPcdg7XjCWSGvOAPndCm+FfVS3C/yJtINAC4oVLWD+pYoZGDtuoCXK
Oxr2vLLpODady9Na6BAB5MWvruV1lfHgMEJOJAJ6sj0l4YLY+6tynbRrJKLv7PQu2i+kmjIvCjYU
4ShOxyE4bOIoReex3n+pdW8Dty/EILbvgFIARCW6I9mGuw8NQ9SAJA/73r/JnKJU3l0DExVp8yW1
ivVZrWHZJbWuRxRmrDbIbO68afpqn2WY3mczOn3pY8w7MO572d6n9kfQWYdu5x0EWZkNSTDQyVOH
i81tR4M13dNexsNi8/x4aMHhmhhnx8KgqzwWSDEz2Ew6RzTc5tFpYCjBLzbDu5X+zT8G9DGTlKgR
JmfxT+6p9Nh7H5a4k6JFAMxSkBu2sH919OeElUYZe556OMS2K9LtFQGJIP3JfokPXUhuqz7IVw7y
P6egUmmzjAdTtE2+q1vULn3RSHzw7+7itzJQzan6ECd6QDcAU/L8BTjOPC0l01EvSlVaudUTu+Rf
ADzH6vIdMRZqKbXGSipVF/9xepioSubn7Ypg+YoOQY5D4MQ1pNNvbnzII6rvfD8OWKgxZ/GCT5mV
C0Ow+ovOMQvDKBF74h4LrSSmFPzJJKIfnnBSuMK6DiLe4V5Jpltrr+O/7m0Vc9+Oo0l6moV3zP+A
qXU+qiD2Z849PPggGhZQR5jtdUFZFcbyhKWOqoyMlv8G0wDoZcIJVb6rqWhJei0jlyfDwfSUa52j
W7RAei40PwZ2ZWDkqPrNTDwfPpWLJQ40FeZpK25WpD/reLvXHnr4JULi5t1m2XwiDbG4E0aIbK3F
B42FZwn4GI/FhDdoZHQ9I4mpjvacTjyUOxHFW7dBx33cJc1jJGDu1kieyf7A4aOGBS/8wkX1Wk0k
jcClhTaS/vQbIVm797FusF4ZXJzt0RBw3E+igDhEpIcVnLN6h7rxsi9jLKLrO3AJLM38RPxfBrp4
maAzh1she2kgTJfFFxhJr8eEQyM8In966vgNqK9uZVhFwSF56SlNIPK8zmThQteJsCs+GW6PyuEN
dbannSWuBFWpjCQwGQFwAqnrwK1yHX7S6vCNKgkCGfZqEpf/ezGLZ1V0NV9yBTHA3pC1zYTYQY8h
BGD8bcMIqw/t9FeEVTt5ECAG9wbXwNGtkqEvgK6Wje3TanJjAdnpCjlPzj6+/spem643amZb587d
S5dOj/IYNwTkPD/ySQQcgyoCwudNKxTIE1QAxm3Z2wrzhYjWuhDixQPi9oMH6w97cO7omfw/6CY4
UILS1G6PVZfJL6ViYgoD6suKkQRerE5O4rz2pPw2iI7jJasIAGPPnqu+qCpFZFO4XHhlUL1bV6g/
JhcxvNvYQt30920lNjSxoJ/UYNSqaM1CLk2yekm3IPVm+s76kNWxto7AvlSdrLKsgVofCG8fZYjx
Qe1AhKXqSmTwjwMBZn5nOOxs2Z4izlHBqB6/pqRfAChQb8+f/SwJs1RwqWPDhLHV4Ifl7cdnveBb
I5xzOssTLxkj/P33Mk24d254dZzsqFeChZmDG1dL/tW6a1Bdi73phBvifk1jTn8h707EXO0NB3yM
i4N8OrW+J3QP3imez+/WH1HRXB6InaZAvWkSwqlS7PBVDw92Yo+DpQygUnJrlnlbfeLG1RvfRWDB
NqC2aiuLS50wnn+ZEGMqmvqKB96jekD6uiEC18rcjrRIZZcuCS28ipF1i3GorxIOXMBv/EtCpvE9
ASI7lZj0ipQXjN3fXqjBN0euePZc0nqzutxJe0CEv5K/PWJoDzQtWXh9Ur9ZQK+2E+MVj1NuB5u3
h5nwGEKv/bAWyiM6Saa5n4Ic9VCslLAIQX5EUzV5Uu9JkWzi8qERsPGqzZ/bss2eKhafQdvHSnsc
p/qsS4Yv4aSZJ2xsCGg1GEb8z/Ex1OQlkiLnDofD6r9md353mKRBZX/L01Tu/53piSHhXaqegtlG
BX3TRIUNQEc6MxtBuTO9Y23MmK0gMV2nCBrHzfD9gIJsBbflQpJC966r0WyRu1jGGPhV2E3BBPz0
FN3FwtUJCPLWqYkzc4jZlYTmIgaeHPpN40j1adxnIb1HqQEEKOwyA67T0ApTsuDssfeGA7Y05hUn
sg1Xb9mu3n3iFZzvi0ZhA2DwSP0YD4/dibFfs11tsS5r4w+KnjFVyT/9hl9v5anoW2t/ci1SADSX
YlFuVdd981VIhRDS/cgQVqffdAuk4d1QKtkaUlm5UceZCgxWNsGw7xXqhA9CvnwEbS8EoYql2Ceh
Uur7cRxVETS0Hdh/6mhHsDgheLXVFw11GKeAS+Pk7uuv5Iv+Agux4CdHQxYwKDj+hOkY1Cn1aaGb
KXmKOwuZYWQbwlkGBc7hAy5j+GGyEfLZwUbNgbWrowkEROyCUwK4ZMts9+3DRtTKAc1YzHkSiV+q
ANzntJG+9rrDueR/DlkxZSKUOGN2yDeir9XNfqZulO8TWz+HeQ==
`pragma protect end_protected

// 
