/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
CaihNQWwu+qKJWjcmdIgzgKIXQ8l3vMImmWHnChjYqoa51yMcErBScyiE64YZSDih9WCUqsVfjEZ
HfdPZ9ljuyASaDAJWOBnJBbhrePBDPO5jKkFmPbv80QoBXSWaNMFc5sW0Ulg3lCiE5qq9SVr7IMd
vkFVewJkI9IJKPXIqEiYLMio527A7EkzJrjUXC11BQnTYghbA5n7/6q2WIDOwjQ+BdLZXxGdIUKi
ihIieqBZEgdd6vwETSGv3sSorIwnUPSueC94L800xEEoFQmghwgPGvLA3IEIqt1YNZfrY4rcuvTH
rxE5ve/ar6tMYP0QdSitAf/UOVre3EWtsP+Jcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="IxINXwVvXQ/n7KwTaYrPoEaEACBK27oPy3cRIdl/LOI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 321232)
`pragma protect data_block
EiGu1ShDtOnFp1/lwt6VhcKuJNvanJd3l3384Am3vLqGekTz+PFAyPnq/uY5HV4vwlfXBzCzWEdZ
4CNQMW7/D3ePhWiA9RP/R5iY1QVPFh7UXz10Z1SzmF0jR2v0EmA1lE7UQd1L7b9WPsVhW+uwEx2p
ljsiFvkGY5AJ08rlrLFxyL10wlSZ0RUZ+gRr5el6aBCQ0EY+FpPg6HC2VBjm4puEEIG1P/NvqsQD
BqkX2Bt05oiEnPOybst5l85DAUsJDnqsNKcEMtc1WQoUfBcRAHT5cLdPsiMrmYKc7Oy5bEiZQdqS
PJKJdHK7mrKXjOt080P0wFaIqlTM8ZVCN+v9nVQEOiktLkvS6AgwUqRZv9KX3ugbu91nsL87YgNq
3kYkOafebEfvfOJQEKIT2UmMFmVwuoNUli55NJhPPAEdfZOfnJRhLa9AydiH89dKSPSuxADMmcDz
1GeqnF9ZP8jaIKe8Y7NG5jcIiQ1zbn5OdBzowrGDDIELZbK37VjtMGeBUv4LKqaGPRfilwC0xfo8
T5unQ564BD17DspIuFPZh/Qm5ELbq9nziXeMjy1FzkBc+0avtsZhKGQRFVPv8iu7qCkgxQkrEaVH
NA4NlwBg4RQR6V0DNvdcUZ/nzDRc1S1d+gGo7JJxyt8B9DcG65Z6GU45hRnJbL2/O4KCf3C5SxB1
bbIy/5DnOmmzib3iWtMDc/Up4dAwoGnJMz10n2ihQIMv0AajfqZBXB/yXtvWAxOLf0Nc39RmwGxO
VDnccPbFaIvm/CZyi2jNP41U/I3e/KIKUZymWmenrP40fAlVxj5vTnR2V+kGWlfZdQEaI0xO/i/I
kuzsfaNRWibUU6YMRCJiYuHyF62avf9UDUFUXF7cuf0mkxmZoEfHKdo+MzQlyzwTw8cj+Aj3IyZx
hIOEYAJ52lH2NIHvAQ6Xeuq4L5jIQTWwZk/DN+qQ7yPQzFMYSs5pxDv4tHaJq+rN/nsDushElrdB
E93GXekZT3Wu5kuf/zQMqkq5rNipCcFT3h4JgZ42DJN2826q5aWJqjnQl7+ND63m/k5evmxcitv4
9aJmcYIkATJtjhx9q7NZorN357CCMABEwuprnl0Kj4bO33O6xjIPTJ9MsmmC1VI7lYKcEf8Mgi4Y
zWZLQPF9m3juxSubQog0NBAhGJpqOEgDt8vcPaFimSPSOwtDNFyCdqC9XtKviXFBMaQ636vcok2S
8tpHZaoPSiaYjGINN8bffJXPiZ7PWV8aspYlEFJGqkJRKKguuRD8kT+4Xr5lw6lgLsua3Ny6uVRi
D7xdqytggz3sZ1NuXFUFGbh+E3olvLxYRySI8W7do0dPJZYef1F+XCLcS/+iUxvKkldTZZ6Yufu4
XQNhnPDf5AOhO6ovG2dQa0mxnb8mDhqP5fcN1cI3ZCs32SjC0h9Hd7nSVwa8biKKxqvhoTNmuvjm
pwHNtDgHre1l9ExuZvM8MyfiYrFGhWqOTJmGKmdJgEZ4I9k7nsO7bNwa31Wfv9mXMs+OunMCDAa8
JiplFthxTEhn3P3c2fKJ86s586UdCo0JrQOG8LwOiWZ3FIpnQQWlawGuOhaaM3fJsCbb4BJFujy3
wYqTrZncEao2mmO9vxyHJcTq+4wUzTpyYAZCnJ2uqZV/NY8yTcAqgmouDIBwi4DzOLKA6bb10bnU
r0H61AL8U0fSDCsu7CAsGPaEdRf40MYndhETrHsC4dZfwRRH9W/L6jA3NvIvI5hJvxmap2FRtrBf
gDA+EqQHCf9CNQ6GpdyFX/zaR1XEUnRpif+IfhClh8Pzu2icEAhCq6q6ZHkzmyI1hVQNH2wo7XC2
P6Zc+xLbK32gZOVh0cKYvKLxNuuRWlWyeWzYBXgB5RbB95lDwj41wPPUL6jBk5KVb/7xdDxlHbZC
ljuQ6OPoW5mUkGxOT/5OhK8GF9keFIMiBWAZPzlhcTGx+az8h24pgvmBA1O1v4pLbhicJEASl/io
RZdfl6bgUat43JFO9GxbiaRnYtuYFdlteb7/OMzIm3i6HqwzvJJPf4ieNyaZ9boJo5jXsVIhG+ZL
6LcDkYpT3BWIsq1FoijtlCcgOQ27E5Id11Uk99TOG6jWAfKBlwydehyGKec7HNdSOFFPizr3ZirT
MSIZd+cnA7Xbafy+xPvBLZOt8FAmVm/mrNBpsXFfHxXe+7HjsJq9EKZgBpFMbIFRbZBN3JRDQcb+
WZrqLP/TOgdYoMzbF/AKI1po1sgzJFPDrlokb5jy9ImaXhcvs0xEEpb57rzbUcmeW4e1ZVakH4eM
fYb8h+gczDyrX7QbSv3YVuuegsBIl6gckGpMPOGPg7HTn8hu6J106EkoQa9p/pR2EQFZZ7rWGj10
K4D+9S/G7tEbFpH0TO3ljVMmO45uebIAcx6a6NlAvWASi3Mviu8AH+GQr8J5i7CkqEslAeTCbJgV
GrMFK1F/sdAg11wpnjfM9tEunkEtFMllTqQ+/uPrFf7KK6UnUWOBmUJaiW/nX6mK0oO/AcaMLHpu
okF0jR8r0fbNyZm7+wbW9L/rqAdw42SN/eHaZ3Uo53N+AWkvfrbhReZ6She0bDN+ywDDxbVHP1XX
vtPFtGLgeedWC3VENt3CC0UaL7TZo8atWzvNVqZW2Y2S9n6GPkkje6i1hZ+54dgR1wq0pMU+nsnZ
hLEey67hHcNqbaJxEWTEtho1W6B9wHMKDqLpvZ/WU8kDv/VWmK7ethGq2wfUjV8ax9cz5gMrOpuB
d2hbA/vraZMXliaFxDyUPFVuU9pcNlkeBb3svfaNNxES3fX5tNpFanxRNaMIve38c9eWUHVsrcNQ
see4umE4LMJgXphfQ0jChsWp8374RKCXc6fr0Uu4qUvfkUIlisAlmVtyEnzaCWM3Z+hw7vxERnC9
gpEO3LADayXFGpcvCCnft5wXV1d38LXk4+V2pELRwj/QKkJOUf/K7L+FdzLU4T4WKhKmK+yX2dgg
Zk3jgo1bVqT8cI81uSkuphgo762Xt3WvlA7GDSh9pz6DpO0ZWteDxw8RDsZqmO9JiGdvbaJ9jgu9
xole9Zp01y9nw1sCbyyou93s/+NrkVMvjz3e7y4Ep1NrtGayuOebv2dpxfj6Xi9lfXVUaAaJFidn
9vYY+jE4k1SsUeilQQJihQkBBJPZNbY9izgLVu9Fl8Gwnuz4N2yxc2aDP+ztL/x51UtFPRPpx3qj
HsFCoNGJuTp7VPb2JSyjqOTAqH7TDuwklZVcUyw48Z81P+ccZt84qgJc3u8DzVsBROE5Gua5LaH7
O7qG5ZphFGx1g1/SB+0aGcPyBiz/R5rhRe8Ra9gfBBsEb2HNXW2zL4gsZF81gk/UJ/9b3hLhnQtG
0YQuZHwgm92y+hWZgjPCD6ggyT758xkbRU8ZtXYx0lZ8zYa0RwBKi0VQxeijl2a8ewsa+pa7ZpmB
Ig/Krkq18L2sWdRJKNITMl4Cq80eLk3EtOfxTofVCZ+y4NTerBjlQJd3Omlct2JIAvqVHhAnNHkD
OjYHq7fjuzDAiopxYooifMK7kWCG4VDDippKksQoOou94roqMGm9ax/3KQ60+q1Yh0niQheDpIN3
ZF1xSdSSc4hlkgRbu/JFAoOa56A5Ox6wO5WQX+AcqQpsolPzxxuCFA3fLnZHieye2B0DetbYi4Bb
HQjw9CYghWQEdZn7+oxUxtrXQpE7IL88u+oZPSG4mL4mpfUOxYYblG7/02K4wxSh0+suFPq+UW8B
Ks5vueCT11iBbcyezpTIaFCG1jPx5xDbSiqFK/ai6o53jpVy4fkzaRvz+NPWswI/7FiFa4oujPbV
GchPVZr4PPC7/MGgsl3eyfo64YjIjXqLq0u9wOgByum12b8pA6FW3/qoWnOKST8wsujdrxvDLbgN
CsmE6nq1gX6No2iNp0Ryr+cLF5Si91PlFFVhFsk5D41tCGmSDTf+58bernJ6LjW5jiYh393nxg3K
se3exDfbj512CWoBlFhdT3Wj6BU+dpN0UUiK2xNEB8hFT1cWLMH67lZeJHgDyb01lLUberHXA25s
wDBO0KpyUNHvH+yshVtoIpGxlUYUTUoMa8fD3phmbWJjalDHEWq5QCx/8tvNJ3XE3Z83oD3fi/qs
AsrW6QOQNyni+uuidZrmAcR+WEd0usQ3Hy9i4e9D0CAYx18t9tkKD4bAjPuCT5V2ptR9uEkm8tRW
CehvxksMTt94w8Qe67PN9+H4A3acWQAaR4uUYROVbkdWyrY3AHhzrbzjv5D0zV+BDH+hudB0z+kI
EkCt9VLYsRm9HgPfbeBEr82dGiMzWG29poRgOnzjgLLp9867kMCwYVYIUZUGE3j8FmqykePSFsi8
zMNGn5f1+VPTAy6FWIBx4YXdma6ofa6tAgG4RJyAHqVBXSzXBi778vcL9Ylapf/iHW2XWM8TQs+S
Rs1ZUllGiFaSZBOFcQBtpQgJ8rYrisPn6JSw4/5WomdChaVfI1i/VXjsFptKWarOaiZkGX9Gsbk+
nci6FK9wZOKVi6851qSE/eYUyl2YDbJQyfin69I5CtHn+FxxGATEN9aCIqU0mJP0bektbrCVOf9V
1xl4E2aIOpy4soldra9JJeG1B3S/48Zgug2dez7dLN2+T95oq1DsyfH5JUzcNOLwdR6LEUv/k7gu
sHgsb+90pTZKYOUULGBsoTx7rv5Uq/GS62tuFHDFjDcm4lzVYg/8w37TBdPhGDU3CSgMpf3Il+L8
w9e9WyZoM1gnR0BIuw82FMqaSfMJrbLFhWT6veai1RCBgl+NMuhwmr02EeDWYq4Je3BjjnrKoegM
ZQ6kl+ITHgq+rhabVhMmqizvykMCRhiaxv0E2Q+r4a54IO3LwHQ3O0BOJWoNpEMiZvnpGqgbUl+e
F2nx7LFE2VDSgUd7RLF8dT1AamXgLJskjj7YAupdZVO7Ehk91nPHnymrL/e1f9UmjEIQhjPW08BD
NxqfHN5fBZHv4iYSX2FfaYt2/mMSOysy8/8fg1mM2gaOwZb0gWYcuDSwWfzpFrnKdQEFM2L01Rkf
UuEKekZEohFOP7YJYbkqaWaBzbeUTUrdj4Ag7iqPLWeoo1BPkeomgco7J01RKgq8gisVavlOHLM+
fY8Uuf7/jGLbixvPLTvCrFCYlWPD0Gq2Ako1JgCbRJd5X6HorW9PwTMzf+qTpKOqmuJyIQu93LNc
DOriPV/Y134oqsd+nltXdtMGmIgmDF90seu59Ym6zOkdKuKVwBaeVYvRVWjAFTrPswvRXn8mT15g
K5OqdBVJHiZe0InzWVyHO2E5vN8VxgDNd2C8dEWjj+vODXpDVtrIrN/gfjlrvFT20uonyUIog+Wo
mTPtAsZPCbuKSjkhhpXsaLRoJO9617LumkkGFXyZxl3Banvlfe3NhK6eAaw3E67EnpRi/URvocNr
aq9gcrK0m4CiZOIflOJDHKFseIue0ndNAB98yWTW+4fitLKlzPPXE5NtI41SNOBOFGrtrqZsJmrX
kMME13XLRTbuvasST3JV58VxIHPthvdY5CnJw4KX57Hhkdk5JZyYQx6uCmbTYEOujqSmK7Bf4gCT
EYHnN7ts3q1VFcM3dG2oiF84zrVzpJYJpPRalET7vqCkXH/pgGPsjx8zoXpsWtxCi5P2j7H90kjD
DViuMaoxo6aunDkMSINeAHY4A0WDnioBH7JAkOPZhki4Jk0IKwICG7B6+BdJev0Gjm1jKzbypLER
T41mrmi19uJHoDRS6loUct/YZR/pjWumYztIh3Z2OhnAGQ14G9S6A8RebueeHPEoHtet1NU9kk+m
4novNUxNCR6lAW8TxfHKJ2b5a4ypiU4WTPG9OMSwijsaLglM6n/a3N3Esxbzk/DNDL0S6wyDhm2j
7Ovz+bS39VPInAJnEh0g6X2i5B3prUpYSOOgux2MuuvYzbOcRNScKCO35jOB8ow8bAxvmmVeN2b1
LJuQ7/UzJ7t9ohPigEldt0Hyou99borSVR4wAdHtNsSNmKZqkGfr7RHyOZ1grF5Oy04bfSF5Djzk
Y0R7X5F3h9Y+1UfmIqCIP7Y+T2Hygy4KjZYXZeSdnf/KYuWZd0BvdF5Bcwsz0EKXiPGI1eE5uMz0
9o4NMGsYhkO0uCU/DTKGiu7s+8+2y+zm6FvFkShMVPdO6HILnRDgvI1TXmsHrHGKotQABtHjMbQJ
5KcRJvwFY/On0Pyy1rXPZSkNer14vX/fDMY3VnZCUzh4xXDuTtwX5g0L/5VdpsaM9+FgiCu1smz5
6924HTenQ/U6l7v0Qy3cfHK7kMx33hePsYEtdjU7vd7zFPLS/46QaMPwOXwdguzcuVG/MeqPUky7
vucFlVi2WNUpFhn2iobmb7KTQlBykvcfHJnDEcK8yWhTafzdHNuyS0ialcGGXqeqTZDs2twRNkvK
Kzwa6wnYXUyhVlJV1t3BjAeg0ADz3hjSQ3wnEBHeqHdR9piTwqmy4fL8NT5UikIwfdpytmbFkqrV
DTnQdroxZ8QsMzCgwutIYylGsdWFpqqcNZpOWg8v8F+c64FHEqnDOctTUYsit9AXk8iwvdtoQKlr
d76PgcMjjZFas/24fOQ5xR/8KOBJEKR+raKK48Vk8zvL25YNt9vmgG/6RwG0u/LChxmSmsEo09kE
38foskkZ9Hs2TZ3n+kDX434HBB1wTHvT+d18x6SfmqS7aqwIg1giBVU8nVkGm4NoCJLjQ1HuRKzI
XZj4mqmUX6UitaFmUlarxp6DWVl1wH6LQPDItD9rAaM1d8KCNLni/GaBwRZIsi+gT93Yan35aA1f
Kz+PuIGMXG2sLlYXt5mugKJA/eTpMFj4XFbMIHThEvwr58COy9nSwrxh+4To3HjIZCCpLfmFASvm
LdTpG7X/mW82ZinmitI1xl1Ie3mV9J2tjeJqtVWl3e7au5eJvYtmjJPxYd2n7c6QsB8UiL11nhIm
CbGtBhIiRcynm8N5xxd6VMfKR18Vy9CacBdEsADXrpsVpOGaQimBnVD8/53fnHEPS2zfGLxXj0Yi
FWN5Ishy7emzxNnigYCsLSbBpuC0y4G+Kk55aLi8z7gSTvMapIl/nzMvIIQbePwQgwVDff48ehYx
6Gg84LnOqYBXms5xm96pbG7R0fK1/x68uo8JTYuvb0X++ATjZmyn1dsZ8ExTpfTkexH7vjvNvy+T
WF/tkLDW0nr7Eawl8yTYzU/7Oj7pERBmta96onONr9okhyhehRjyWkGlXFo1bDMQGvRTp6X+dSmw
cldGaleRDIIfG+yBUoD0hTC+sn/E6dOxhkosZKGxLK8de8JjRKa+bdUifEUi+798z/1R7cS5wPsY
4t/3/P/235XzUQlEVtMzzBu/Blio4p6UO0yOqa9osSTKFj40wgYEjdUtCMasxQwKdLE24zEQpApi
LsOSXbVyw7zrToJeI2ZRCsCgNi5h8QtCqJBDesFOYDaIixKpoD36v2cVthW+n3s++KhKqJcnjEYT
2jSVCYI9b65MiyJVogvan6E8zhMnr7WD/yDrQZJNJJvbu88TYvsljiwofFjCm3g3IjZov76afVlM
VDdu4/nPWpXPhUq3p2/dIZnUWnEIHxbrNKCLrrso72VzMoJsWUxu40qx3m+SyeqINljmm1+X3t8d
v9vHaaoGfaFKdgqdMj+SLVZycTKdPvbvlXvnZa+RKVEW9NTB1MD4rkyg8EPEq2Sng2D0iAgrpTBa
4edq99NfouWBInJeSZCWDuzVAqbbcYplVlfT7pSRRe5Gva2XfWHM46V3vRwE/clhhNIepdCnoSiw
U82qkIHwHnY2erHro1DMx3ii47tBgwD2Bg9DpC5mYOUOem7QNGuWJk2HkilSh65b+2zY9WdjaZz2
L2eX8ZDHCw1EzPNf7++DEnYEe9EsLB5lVAiG/oSX1nGRTfDThRPTcr25rsmNxMBMSvvr/bjefqrO
qquv+meExv44sByNBcN2Wb4Ega/ZdeNbNqEX8DJwWilN5bmzSf8aasU197+M4oYFjsLay+DTZD3x
TX5VJbVO3eYdCn+0lnxD/6tJ0UppC4EgvzONXXD7wFWiYig8iVXTPOv8c91P0bphyLEufdY4wiW1
oRcnw/WEG8YkrAWlgGgw4JgPcDuUKoaoQpnvr/8Q4tgn6xhAlI6ohXYwgijXe9YdxG9w/LwFW7SI
1JeL9AHrSVpH4civOw5t7oLu2ofPmDm+QcvmMu086kSWVCJSz5xbnePJ8Lhmi6CBwn1obUPp4BRB
7CBaCWZ+iHme9hnsyHeaI6EWcksVtDj5+N9OqwnfkIEf3xV+B6FR2/N/inV3Wfx5u4SaJdbW5Abx
x1hJvGFgbHLF+rpx0w8wjKI2S+UI0/dGWFcOYjkU2FSrKUhZNrdfdXrLqiV/x9kFo6RZHp2nnWdu
SlToq2X/9PjhdclxGgJ8fh9/SGOcNNLpx63cecDdwLLJV1x/V+N03NV1Rx0c2EWiA8VM/Y7S7D9A
7shVIR0FjZMcl7R9zaYq+JoNmKO1xkBSfV3ms37/FoPLViEZLrDQXMMJEZpJAvgZipLXX7JRttok
3sEODT7nm8Udk4XpTu10U2jvedKhdS8tUFDbZeS3zNKtYRkaU4xH0L5xEvpd0IPQEQuSZ4U8cVUb
8U9t1IKrvQG1tB4Xs9+30Tdg2OvEmS4hOPs7QBc3cnqEijqvunbK2bZ0Hvg2knEKycyt/kGoDyCS
gB6LCAVu7K6frQKGFbyWEMK8NQMJbWVg5oFqXCejs5JR40mwri0t7/4MlmgbNHPkGFg20x2DRYP/
6pkacOIKfMw3amjVKSSxQMC13Ozs3+TSmmVaqXrnyrUGhAuYLXSAIRh4DxAo7SWJ5JnWTT08SLye
Z1qXQWMH0vXt/1A96qk9sfE9z6wuZ+SFpv+Jw8ic0tZRv8wyMTI0FrOqIn4i3WX2z0p77wFFBGQs
LosgIOmoU/dF09tkgupMyEo3xpabkZ42sE38BAfJpRuS9iHpGuf0t5jVl78q9KNd2DGmugLJTRL5
bZ9q0YGDOkqAZs5QD5J6kV5f33woyJiLD071hfzKOWH84zy7PWnJjIuarcXxCT85ASCnEyl9rsG1
A0i4l8qhV5mT4UdKfiUwLg+YQTsImAGNu03z+0xnDgAofgFYcOrQzbkBPJXxADQIz+HFRvGz4x0Q
RZy/eJ0pOiRe45evHIRgjuWz11DWIFMD8Xg1GoRpExTDQn/Elskvy/33qTrpCavAy83uZ+77UtPq
09dHIQkD3iCb5JHwUStsX5zJHYPfvX+ltfsPtLim3VHcJhyD9SY0s54U+njQJZMs8iN1uNM97Fds
5F1zPYHs0MKWhpMlrrc9yVhJPVzCyC9lYf9dtLKDxKsPDsaRLcG8QMb+b6Xk3qgSz45Rfp9VOD74
8S9Hk8ATkckjXa/F+FsCx9o2oYZkeSQn20nCxXmXM1jnIbx5FhObAKvTbwFE5DE0pZCXUeCADTKY
riHBZYzy7vIZOahIjYSlRa9jHzdCy44gfrNdSrBy5P5Foqavt8KBZgvtgiwTkDgfH+tLK6ta/A9G
7XRGtPzr2ntZI2bPvJToSUTH4GE+itTxOWmNFi50dSj3niU/ILk1Wo2SpE3r0bzri+s3NdoZ9vd8
KGJSH9tJIxgfRCCLDJDK9tBu5QWzjbCDOgnS4CXwMqxhmMDhwyQZ/BIt3thJ+bCEHrydjX9BGYXf
JBuFOVkzVwD404/zgKID3losQTc+kMy+SuFdmiQBkpar54Yj8zTCsiY0qrasQqo51cipW236OcyP
rP4xwISkuJ9ooey0uIfFAI00ZwH9F59FPzOizoVEPqg7PBNDhYktjzSkWwwd3NLFkuIfJeJV3ihO
0RAVguorzHxANBfW324VQRprVVa5CvtR0vCMxWE7yVhGSxEmGwJXWAwO0ZQMUOcpj727ZCx9kYoG
0UiS83ZjAdavOugPDOOM6LzGUiqkVRLBEXmwi9AKhAkVDFlms66HBuhnheE9UttIyUkyxLMIXPNR
bZ9G5XPct8BvP6dOqqzsZP/tdbW7r1koEGjcexS13WUpkf7zSDRGlO9xvtGdXIBnqqnXDiBljVfP
CdqCzYheeRXnjXOEAt89EQM/vCrud2kScfhsknYC1drfBpD63fsD/NBQsOenMdH/cz5nn7XYUZgO
ESOpP7Htk3D3TWs7ZyOyRw6DVUdAv2unMbgS9dNEK5ELeNO766+7uqqYSY5RHT9LrA+T9VI2Q083
u6vZpH/CR8jy/QiWKePyLHQxGugZdFjgyyAEDoiV+hHquZK5z5oQOI2o7ISqZVPxUU9YeLbNwt9i
o4xzsryPg4cHvsHbbBknHdY54/MNgvWm/dnwSWqx+EhZGdLU4NswPNmvXJHuD+iN6SP6NiWigPVd
ixUM+KR8y/HdPAiZ+dX5Cbm4dbKvkUV7QzPQQnQRKsMEGNfDGmrGt/jWjqvpigdJdv/YrmkX1p/q
tBboXdR55CLCKMUuVx4vPpwLJS/Sjn/6R37UybGSCFx5tj1B+G+UblXGq8m+ahMSfWw/3BHqVB8r
tM7mwgPbEyHe12tlPbBVJDH1oojTQyzQAhkKYFSvBgr1xTn+uNtvAHTLXUIfvRXmeYpFiDnhDxNk
ev8cZLQDIlE69BN+2Bs29HFH0r2hvNDrxcu0sviCAf46KtSWzoq61zdRM9BJFxeZbc75nHouovi8
7BpyAEyguvyLn8a9b5jG2lT64B4oGNbs4LzUQ3YedBtuGEobISyIYHkCobtSKUZfaId2saNOanMR
GKkiMHQl+0UrfXlxqid+kLwBD7tAlu5yMeKke5bGShg1n2ziEowPDyAujnSJ0MWPST26WtJeXweD
hoSveMAaz/KvKVEeUy8UEBwdfpszNOkSI9P/4fIlJgbumYzEIXTvNmkIFcIYqkYtY7Kl4IdKPudR
mCvGzKHQCkww+s1Gl4pza3rrbbJ0pPZI9XBcpK9kNK27r/bFmM9JSRZCHWRiB6ESFsLA1M9LZBXe
yQozSz1FSgl3RK3JqYS/q7F74rIBcwM5Xbiav9zW8La2bfW9YTD8cLdp8zBhRCoR8WkkWH8cDvJx
ZnScSfNj5FXGdlV8S/5+5ZuPmYEgV/lzdczWMSeUB9y09MEmVT2Ek5MRiwwUw/90slvdQBq5cwc3
DMED97D2zk1b0LDf1UaeOMZSa4eYGWmrekUgoWpwneWOiSVyJmuUkpHpsHbTIeUN6ARHFRPLDFus
mvhvowAd1rNJdgwNK+UFJYI5NL3hWd+58mDUORZda9QW5jzngT/YgXRzrcRqX7Pj2BAx2TmMWOmN
4WdoY+8Pq4eQJ9g7JVGwCehC/j04vfr1PDurxiRfkODodUlVgJu5AKZPtfyOQV5byf/lZr9nGujG
H884hyAshhtgjAW+bWlrwNwurjU49rbaopsgYbo8TQUChn3vdNtJiKbgBTVhycyOWQtYyZ305EZI
Gsa9F8IfLQEer1Mx5rHcrQuZ13nlDBFJeyN/02wEQAib5Ix0wcTZKOfTM+a0dEr3AZ1NWfWJW8PN
BDZ5AcCxk1poQ3L+0dIwwQFW+k1zIDpoem0rIl8UUejbTtnDkW+XSlM3PYSHWyLHwTAltm5CAIwd
Tv61N69KrXNSg/WKhV+V3iWfQ68gQOh3+TutEtBiKdlknXzbk4WDYwmWxbTkwYAu7BPAYszBH6KU
tc1XONsLz7oZhFQaVc8+/IWIm3DBxsWaZ9etNz0qLRoObfR8tRjncV0T5ktcx+XBeKFU4f8fDxKF
BZIxQes/Ihmm7YfRuQRpZ3hSQgh5iKSmmRDAGlb7OOxrRmKCkJI1v+biqk7TVKw5zoEVVJ6Psje0
bZJ8j6axS7f+5Typnb/SQxO5rQWad3bIIRnXxp9b6ChM+i9Dbarkumu20uM8WIzH4Y/XZ29M729S
LywKxhzLa5f3Tv01aizkDVNINZ6EHNSHTuPitzpx+bOr6ScqpqEqOpgzzvg6haAgNKhCU1Z6n+zH
1nE70mzwXYGI8H5uGa/2zpq+FFpeBoXsY+ydPdfojjZzA4pKiiphLEFJ3RckW6WEHqJg3bjpETsp
P7rb1tT0dAKnNZ+cSDRlJzdmIkUnWDGpaznZHmpdNOKouyLLXrJr8HSb91vt9VOu4ZJmVajjcEwI
SGil9VmCYzkmboFt9J5/Cy0oW33XPddSiNu7LlpjfybeV5zhQb2wxUsRF35UCfU0DyOAXL5eBHQc
SjBxrGw/0xzA4CNKIPZKUm/mggy51Conbnu+PyweIoBmDgGyBIh29Zt5Q88fMpnjcixuEeU5psaq
R7VSVFVTmIbTrQ+KMi1kxSW1d2IJRQ1ock3mDbP75EDZLn9I3+O9VBBpEBLl5OihkBqTvKMgZNqw
a5QF0ahj4IPv+XiMrcYx8HXrxlSAd6hLhh0Zbjlp8gL73ADstF2+W8eRdtrUxVNMA4WV2uafixmK
HckBctoQm+GH6gHLZdXiR3u5nXnq5hmq/6EfYgc3tyJxl6XXnPWHWBRpKZeOhnIBTpEDJCNgy3To
VmwsaTR1Hp57MItQ3iYmcMSfaQWNTA8j4DCGKccChiRhY8Eze0QSWXreI972ZRwj5wC2a5bHYsmp
Pbhz84/LVI4/F5/1yZAt8f2USCL5KTeD8iXrouRgYqpGvQ+6Vy5ZLZb2RXG/hAhbvg1bGNL+LnIM
tgYSYVAuyPdgV8tpHJvAxMZn4GkluNx6ciJQ6p2a2NGls+yar+vEx3zVuB3groox0e2BWDMEYOE4
Bl1+YjLZz/ftSNQ5nrA5pm8emnyQb9wgMjG6jC8XGhTXq0pBfSn4XlYphbDv97f2wC61Flfm6r0E
MIvxbHK9TkJc1A5aZd0mrmVs5JonlFRTh1eIdkTpud8gg2qTaAfRcy1NyaCgYmf3sXjptwEXUXUB
Xv3PyAaVmYImrC8MA8ZKKMOr+PqolCeCOdgnnAD+YpnW4uRTKsSwicLhUT5MN+M34NzipYdnxKJu
0rNb5dqVzY4jQXDuQMIWiTl2VKLmEwnHxNmQpoLc8vb/5abu+7xeNUiHjdhX4q0nhOlTWtMBPEGp
8bkwVymg7Lwo8iwpyiu2P3Knkma5j3bgl5zLSX2Y9D3q7Gm4vgYbMHG/kcGyyaaoZVhiUPSasxhM
T/xqu+kr/7sHTAWbzRq4RWjhFXLmeUQvsCj+Lvwaez8jqYguh7oKGxOmXFY0wHb3u0xTHCO0kL0B
ktnaLRs4Dh/IsxNxWnygHRIRIIAusaADtox0fEf8QCY6CR3ao/9ZR8U9Wrf+SbdNB1vxDXq5xHYI
bjupXnaj9zMY+5zA1k7EqmMWLGrhuC+nmfDkmvviL+w7YrqPEPJNKHLfce4DVSmFj9Ml2zEH9CFG
48RoRdYIbMGmwdy9gCOoDHQfyDxTeddOnf1hiPO6KCano8sCWalZv3lH+aYvQ97cm2FLnqmrqHNc
h6OcwNbC/15VPIkozAM1JaytnonFREm06B8FjZ7o/q5qzCzcOVlm5b/3KoLHFdSOmuhEYTo9+Y28
P463p0nS6AYMmyoiYPMVcaPi4qqr3ZEETVg3h5lqO/8jfHkKXuDBEoAu6V7eyMENL/OSzCvJWtId
cdEU+0yIprNLfbJ0GSwIYcvdjUnJoNRhBr/M4iT1h/IXZnXQopnXOSY8/HCfurqTTj0yqIhZdi1o
+X3ee70fri2yVRSNymXfaVlWjgvhQcb7nZH4oMi/JDGr5YynVFOB4P3s6zTRaC8+noIwKKPxMtYY
0RO0zSKC4PXT/TBQJsbdl/DpQpkxla7X+RAmfA8jCvoWqCAZhGUMtTqei51t3Ie44GM+wRPesfg6
YuBjqN0QN8gjjt3Vb4G27dpnCTDblI+9gwMDPGrUMgDNnJrSODtDpiqvt4uj06Nc45P6mA+prroK
1lccVjl7xiODT3qXfQkjbWIEZWoP2FWKqBYF9ADcu/9MDyubbytxOWKxa/sSnUcNSV6U21Ccz8vD
QnJEg+LtZXvt9fJNyx0pme3RPndvqy4OCPAkymON0pF0SarCbRdaPJidiSYtAPG3Y/h03j+S2z28
wy+PcTQU1PjDDW+FxIrExEG8Bgm8nb9XrbMQHi0yPu9ngkMViNOm6yM5pq2FY5dmrSit+jRSppiu
1bW+Ni2k2P4Ph6+NSVtkpYlVgoQGnCQuS0Od1SaAIo9GX81wK8buvUluOpl23BqUpDZKdV0ZbtTy
LZmF9BMyY3jOGP+mw5/ydwtvxEgfcjo0geeu9iyikKgvQdpTBLmGRBgPFotsh2etmJinQO4eWEZi
ajUntBoAAQFkcg8D5/bvc3JmYlbNPZGecKMlik0b8LceJp3EEW9GkZ0m78sEAFWHvoqslHDRds/E
V/ne1dYRdTf0MF6XeUWIJpfZ2T1iAotOzF0g34fYncxu7Og3jfIPf/h/LcQN50/94lutNM/wTrUM
h7SWcNHd7+1MO3mC0izvD1dX367FuqPou4Jcdp2LoTDj5ROYQ1GZSVkZJUfq/0ivno9lk1ERJuYj
XLDPB87JTtYclMlnZ7/EunKbKmFG3VEeyhY2SFgxbjJMa0oM+WBvcx6LZCeIeZtQ8e+wd9tKUn3z
Fo9E1x0FWK42kezoEYLuNrJumruT9x2DmZXK0YvumrKUFSzo6ecwD8gQj0TsRZ+Iclu4Y21kXkhA
B5wE7YDAkIawJPoZDCzwWFbDf184VgeLh0kmsithz0QmkvjOo9teQXBu7DTUhvX2rCjXKdnOryUf
GYNWyNh2nCxutgzQvGVGC2H4SajFToraIr/HJ+z8Ort5n5/hPfDA60QaK4UNO7acKBbsVyqWyqTw
0osMmgcCRh7KEaWhlDM0183AJYAfeXhfvj1apSh69gb+yJGF2VywQOHOM1ycJgN2EN3mqzMFh+v5
E23cm1/IGBuKUuD/8R6F7Xwm+f5VxQ5GZQORcgt6rqOIyGXjwhgpunkypyxbKEWOCngYjm8OPNXh
RBoOlL0aMkE0O/nsXkNisP3oIHafhp9qSYPxLl/G6b32BbJWzNm3LRQSxvkBkW9Mp/HFT+UXvoDw
lGZZ7PKicwSqs3gC5cTXjks7nc83NVYXZI17NrvEVaoVpgbyeZvjnRhTmgACqBcGhPoKraJURQxK
2e2uE0JvADJCJ44ekdRFajYhaCBNw9EMWJ1VFjZJ22aVmULeAdnVskmo2cRy/E66iiyQdRvpmUoS
j/ng1S7NQPCGIOBvlyBoU1XNTq1R2spd8+DaqChxOW1NSIvgwsxkKvPFwOwGM/9gYVeVOKLGLQkZ
s70ELsEdh0r52FH32tQnNqzBGlIbAGigFbcn0FR2fKgCfR7EAt5z1fNdfm/tHfunDNsapXXjPoSS
mofgk894VUjKovZUTQXZKKHLK5po5wyYQCt+yac1roKsOyXP1YinzQGviENXtl1kExUog9O5UTc1
ZFYeb+yc/QYPh9O3guT1l/VJklObvk049eAfWPi1lWyn8mtUdrMwbDJ3clMo7WSDU+Kl583bC+mI
DlTxTAdPWo3nUnBFcXFqs5uUCcBPgm/Uy9tp5Qcr9maVCYroOHu+1WXfNjXWQHEIIMBMkKeQxYyW
g9soeM4khRopjmgGvgbEvGBfaggY73nKlxurbPXamK5qexA/KOalb+O1kqhLBiPQDWbTMj9rpDG6
M+RLV9kEunlJRPnF3LmkRNBG+iumjmRO7qwocLelPyY+3TM/S4pgrAs7zjIsbCqEoJy6qOiwQEtl
vrRv3qvex6kp2+i7NVeXlw73rC/idGRegp8jIiUhBg0wYv0hKDhx0xqScQ3W4oiFli+hBYulPPsf
GmbdQn5LP/amMHnAhH9Maaht0aKAZS1zs+pGWknP6mUeHwK/PDt5zcp9wp73jrwK9fujlpaVZZbD
6ny31Gm6RAuQIGHSQdGrsxvI6QCEMps1DEqx8ZnW0728+6y3da1mchGuoQ9cqE4yE6VoNonGZ0o9
VFLwtteWvd40D+/d8dPLHfIMuAPBBXSZtrWNThqenPWIXatsgXo7ib5MzEI2eiUiq+NeDy7u1lWX
PPqJTV7rS3fhHBHohi5tWQggpwxxtpHKLyPmQv0L5GLUBOM4lurva4ViBdYBAXYZ2K68Ux9jcywx
HRCgGZu1+u+1OV52NidaY8tbEbNaBkAJJxRZmrDFPi8lziHfn5NB27aRqFY5ZJBObt3V8bKgbVGT
+wgfmn+bx5b/2EudvRhKiutg2vVeWtPaYZ37xniyMS8+DIa+UVkR6dIKrhAUbXcdMrz0pWNpGkKm
czKsQLsEVK4ZkzmGli4+YSIcaScDTRLdmmT3h0PGxbztINmEBAo3AEyZ1q50qFCGDZglfsnAzIfP
em2JOHFT7Jdr35n4lWg2k89GyY5d3RkDOycMnfKrobIY8Hhstfi+z8m1bdbNvjhsi0/eX3b3s/HI
TkEBnQFWMqqBwX+FAKM4HBDS8/YS/N41a9d6ktTlMjQ/SdOnHzxhg+XPiaN1PIHaUfSk7G/w0MqT
UAEdsqpqP2QnVZSjEYUS257KIVKyHL3fhbWAWEQdxBdXOd+y6fseB3vqo6WoTUPOWaknMFbXMhs4
Bi8x50bh91tSlEKjgM0nOL+PPqyMyweyOuH90b/XFubTCtTo4mgBz3l1QSYpT+v7Zym9jgwqzAaE
Ap88UMnc4xX4NGFd5e6O5piwrgOeRepVbfU3FYIabWV3VbcMEdXMZZVLryl2tFr8e3jOqTHH5qN8
ASrlQgRxtUodjbqMqM9VT0bZddIBYNGFm579j0F04tAMI4pu+EYz+zBE9T2yk7kUdrzGV/0+prh0
Z5e5FfybfbmiOlRVYThi4WXN65h6Grk0maxUBw1VzjMi5HaoS2tBmAOJ9f+28aGUQxCEIPBL5xsT
TzIp/CpF1MfoX0nX1VMn/rXMF4k9wb0cGaDV7kaUAqZINN2ykbDAk9lmPNBAtmjIu5VJ++uJfnl4
mwmcZZWZM7xb02Pq8+XFKyo0QMJxH9AbMdm+dmcT+Fc6ZEe4rwhtvzvXqbJ+V4vnBwPtjyLqUl9s
8GDotho08oZobrJOgtflXiwxx8lxGxhaNlut6FQ0boCAC1diJrfo7WzHz14K7gP3afDWsdEDYEOX
hdbpIqQ3EuxMX2bH8Bk7m9bjkDanODnX8OUtvnueAQuYmfb2vS54NiCSPE2qZ8yM1BELpjAI3lvy
vmGMIXJwGStyWN6lAkHs9Vb3WwWRgurfjKb87aIJtUPx9NPZYE+p0LJJppH7pTbCpVb/BXFiDPFm
lM/58MN/HnjGSasMtrjIDoVtwGR1+a2BHR5jZ0p4i8vpOfA+u6xP1pJL7+I9iyG9KHELnuNE72lq
TeauixgBIJ8956bkCv0w2rI5bL4pGPfNKFs836nS/6MwZmZI+z+SET2w43JLJA3162ajs9BDcxS0
+JaRmbruXkBXQLPF4LiII8Kuep22JzZsRq+zetwZWU80BIe0rUxZvyC8ahQ4uBK2uqvHAu0v0NKW
R53ciVBO5eSMIDSi4DhZeeWjVVWhXh/sTUX4GV30un14wuGcsWGD+mr8ftfa77OSUfx/cD3fsg19
SAydSIFdu/GPQXYR0j6pR1yUyJRBauCm8MHkLIc+xMozoJdW5VrRsNa0GNy50kwqazDvam0Rwpo1
/6agpU2q20iQA7zdSvwiStuM3g7H0gkS+inFEHSlcfSx9mwA6Lxwwrke60V78qr6tWyn+VGalueF
FWAz5SpBgZiv8HnJvng3rGh3TzZc/dciQjxfs8hacql96u3Oi0eP9wBQX9BQquvkyOSrSGWJa0HC
oh8ZU5a1PEZecYGxcT7BKPuFPHVzR4KJgvFRURM3a5snYZtAEJ3PMzS96Pk7HeK+Wup4Jcvyixsd
hb/2f5cTr2WezU2BZ4Sncz8AV4Q9iEmYCWDgePATLdJuEJWkoOE+AWi0woZO8Y9fH3dfZ8Go8nZf
vJIH/btLXqKeXZ06GnWXqjDdg2lO/Utlz0r0aG4W1ClegRu5k09NtgW1OuBKbw0LgYMxBNmc+opA
v6Ayq+5NJC0b+zx1d6bBl33RNpXOrSEF/KcSqh7EFwu85rbloUTSJeW32DjGBB23mpqPC0UfoYHn
qBaJVOVSF4ZuKbHbYzAp180NTEiw3LKWzBoUtqCu16HrE9ZQwdcmeub4vH371p55xruTpYP/CHl2
n4y2Z+y3oGtvZ8RwPKj1U9bPr4letshpv202z6eGdmc4LSD+zsbJWgKzlogVYh/k7+gVdTiAbxG9
jSu5cZpVTuqkRAu1tHWHCaKwFmwObqIBkRKwBTbghCKxpIRNmBPpyg0OhiPqUKNATaNOTxvGAmmM
ouJIoIAlEJdleY17nR0TO0IvJXEqu5fPWR4NYpfGyArqfwh/vYVVm91Bk7AozeMn0eofVsHGgkOQ
3MSRxFhNMM9ezvFZWhMYkBlBF/LMBZnCaij6X2AThoHzzEEJ7d62ZFS/WqOKNMD/inarTLD2aXY4
AdZalgdXwRRD6Q2t2LDwBjNQDhQQjFqY8D/LCgqbLGF7/579VudGhnjEMa4/YfMWRACVywYntWry
kC/M4Aa3HVZW+D96Isf3WdUWVnxggEx0z7yDwkAXnAxKDxTmLrbPZ+gwYAghk2+m6Rg8sCWT3ODR
qlhncbFIV1wPYRui+6bhqofz2hYa6ZzTCmPz6Bb7FDRqXUmDGPgybsB8aFk9cPEK+PTypShMq+ll
JxrlfWh4FiPtMrEohYWM5gunczkuz3/ZmEziR9jzo28yo/mdirdVGG5ikB5leRPLZNFaPa01TG2Y
J4JB0zNFYWJsVOcFTk3ntaFq8spgqF5ahM7exD1VAnI6qk1sYzB+8WVyXUczmTtkUk2iV2zd/xtN
GJnwzeTJzq4iEq2fswhoem1PX/4P2PpIF+DaDum7n5+uX2Lkm9Htf/eVVhukPlAxEWwS30KikIhe
229LdzwZEPr4GdhfiXbFdUM2RTg3Vvd0n5JfaJQuIfyjeEeWYPs7fowlGdF5ig+HgQCkTLVi7uKS
JUyv2FRrnuu146AF8ArpUW5Zc5m1d9YSmy9Nm1FF2+aMmEt1T0wynCXcyp0rZ7AAgHshr+zCi9sF
71xEbwZ7RMtyi6pvzqKd5mO3xYgYkvj1rtKqY7B9HmyDq/jxsFEBUwdL5WOt/snNzMFRIjXT5+/8
4f2Uot73wNhwdIrZcWierBiMXyb7cmgbc8I9HlkFnb/qV1gNHMActOXEPtSEN0OcpvQgDIlwJrg/
RJEfKw8eF/G44jINOISSzRLc7LqU0sV2Aw/gnRzvHr8A6qUjyeoZk6K9F6uyaJ0aWZgEB0S5MYSj
3ajp75Mgcfvi5McUo8gdcpDmUP06qLCT2g+Sgrqes74YIKFFHMR6wb8scz/uuI92mK78iJrJdNej
SW6MhGGHpPEB36Nw9gO6FWfR4qUlTx4peLS9hskwYO5uriv+Cj8s7Uw7C/F+vEYaR67e8yx6yzlI
em6+gNMkedXC/zLUvbGM00QO0OVknYbA/rpdDywzgTap61FBrS6dNP3onnLobDiFkyTvofviSNW/
s12nhw1tP9CcH3wk1cKK+is1fO859O1Rq9rfdONedjXSTyVEjeAxD3xAdGlPJHecFMQv0cdfXpNk
1NgoceGRRWjCnESBU9O9MdU+w8NdlT9kqa+uzpsEilSWC/5v9JFNLsGPBRLHJk5xxUNr5bWQtCdF
PWja2+qwTxMnxiqjLhRft+nW2wss7qK4GzqtYNkI95o6VGmqVhJ67w2KLhR5SwKCQTeoLt5BKZEU
XiZToBhV5aaT7oz/0s75+dIoYuST1+wjhig23HM9FLu2ZUKQwoOUeLP6ur11HPMuyu3u+KBSQ7Fw
OMCAkMVYVkZbqwq3LKMYePckJHgIhYOwbOOphHUAX5y1807IgmoxYQxnyzaXsvdwgtXMtb2Tjk1T
NKE8WQVSKJq1jQP/iyWaW5gVuyovE0E6lbTYersCPRgxjmKRFPnSt5EvkakMl4gABjQT9lbJmnRw
1+sE1a/9QKRXEGYfEvzVHMGyxQAwh7qSNDNOOUgC/tSmF97eir6sd/GXrgoHyYIP1IKUJJ/LfEqB
3/zoP1EhRyum0lh3keZAb68gHhJInrVxeLVPXttwslKwIUsgKb8np3cfegJ+GCKB20fqaPxdjWdp
3/L2X8uAQNAmwgo8crRmxpvrlPtvfs1I1HuO4ysAN67P5GCZVGEpn7QxgmcGp+d7PNjlR4Vf9zbm
ETmBswOFGNh3P2Wq15SAkRDlyFLyQcs927LY64Mn4/IeJ7ROAZaqTsu64yrviO3aXpA5CzDkEKC0
XzrpIWdPk1jSUURuplxsoFq8UDUEbndtgKyGP2xuW9J0LYPxQUpIy6oW3CKuSohQEb6puR4/nXka
ROzP2A3sz7EXulTNrKX7tKXB6iSrX+XsqHB2JqnZZszTW7YeupKQ9/GLiBzdRpQ2q01zWNOCKYs0
6nt//ucFYEYv+YzTVeFamZXpZmktmNIBGoq4EVTRBhTmm0pwr1nBp+6mjv2s5RxCoSBqrZqc3Whg
7tUlrYwF9EpPwMnR5jPyXedGWhb3wYV9CkrbDrLRFYkUE505UMehN3AJ05y09l65pUy2Yl46LSkK
RujNkRB1K8xnLtYlQSNgVc4hfbu302cui4HuVB+5oumQW2K1pRirMl2/RoOFKU7/xyZiW0wPrALt
kJvIWIp8MPLsqkSq09dJ96vEQ+XZuW4VjwKrGKgQ5E1GeMRSmHNe9z/Q9INU8p4Q3HN/Wd+lK1tb
40Bwo6HaI4WcC27cfQAYsDoiRxo3VlYPNe8491RBAZZgUXf1Ket0BVgcJ7jFaluXQlqou/A3ybMR
V6KVQf7Zpixl7t/Y5HIWLcPLwxdkfJjnPeBpIS7grkLhQ99krCr8QeSitHfvCNw5i9hRVIR2lFWb
eVVDgO3tgx4uh8MjC0F7gCkuc7cAM6oJaSrs8yzPdD1d+7Vs/gw517AVvA2tiWvor0EiZv12yn8z
rQOBVNkSntUxnxPL2X69Kn5CoxdEMXmoU1NEgIjAzIvgfGbALbz1dk9SWREPnVfvfMDxBhXYfMTY
0MC1E8EmXvNxg322DHSHSt8F8w1Hocmdewxy3SaYEcgm6BA9+huY5e2lUv4JdE8Ne0/ktuFa/qfn
jBGWJF1s8vOWzfTiv+Ymo6DMu9G6Qv0aUo6ybxqj84QjFK8cVpXyacnqYWbn4j2y0qI+qI913Jj+
P1tsrDARFA0G3MTWNvUSdT1TPOgwnHCMUSS9lwMO/+KFxEeRHjC3xDYRnil4kRG56qTW+fShVCuR
1FJRjc2GZ6rwq3b8z0gocGRTmDVl8gWK/oVgnAGgWOwMARSVgiM/vKM1acu3PigNt+H20lIJVZmP
1PrMZuBjBNtFQjgYYLtw/C/D7x1expehyAtNpH/m7eqRBeQ4gO9JidBtIhFZ0DPztIJL60hcnITc
f4aCS38SXu7QGT7IesfeTV+hhvrpCnDTBidczKY3CAxqrE7MvKcZnIyPIo2r+GFfjH+eP/rjHesj
sXRTVMlMnXd2Mw+KwTAO1ZdFS3cnBQzjKdESO9Y58No/unh5AZqoDVC9il0XXsqETjPaKj5xfNy+
QOjzvLwZlVdSgn9wTKnEmykxi1m0H4Y0+cNjvajltSFnFr/aOvY4abltiHCbUxvhC6LP17Tyw4vR
VS+w8oQEmM8Z6L+IphwYIwlyuBA0JaWNsbqF5g83KUABcxVkRXqIcUea2udoVTTpgfZqxBlDWNej
duREhYgmAWCNNAbyakIAtFjwUKXpyHUq9Jlf9E+9h6bcICG3ZNEIfAU6VdKqzhqBjJXz/GxVPdWG
3aQgDvBUETacIXCiJ9lnefLhzNhem5xpTqmLwHPXbUdSRm7GTHl1i92inTJppVBqlBe0CW6Zv5j8
cLpkmmpH5ZYiLHPER8mxcqQPwu4gcxdZDC4hlTauQoOXSAD/R387qax2d5h6HQ6vm0/hUgmxrshj
CG5UoyRgxCP3jBYAge+IvyE7OunG+jZRFdxY3L6rIcdg00BXKJ0C0xO3ufd03uPPtbAPQxTZyIt5
2Dc4VZoNu7td8eRmEnDAFK3D4ysNuZxFdlrea6fImVlcThrq7crDPQDKR9hl+KN9YYYMFhExt8nU
0DsNdrVZcgIUik84U81oeL4xeH/3HumOPgojHNVOt84Uqwh1W5xOKSeI+9IyGv2SwZH23KkqXcZJ
JMYXTMkXS3vaAg8e4bZ71alU8bELHwA3H33l5sOr1fLbnruclYlAtK6Hje1MYeiC4mfLO7UNpxm1
O3/QhYwFuQ+7AUXDIKRJoQuYP5w6HuiCC/HoYTsx4RYezFRkBhHO3Q03A9NsDGzGYLx+4T1wjp3q
o4y2HcS1Ity7//1sPj4C+8bpvB0UELjAvPgoahC2E97CoCpNTr3uHPnFLwyuqJeUbNpEjyxuTqn7
x4QGJ07/eTIYigcO4Za7p8PcjMVqOmIkAGwczzVS3CXk2/oiuPHvicdpnwcSw9Cf8wvbN9pY4Mwh
5WCJ/uhRqVb70l3hDTUaQVZtp/jyS2+/ELXjYV7753BL5Lgl3H4tq2qCTFnCTx+wxkRNAP3ix53L
k9A4vLAewCjXI4x8MBreFceTARU0sYds8NwIVsnygKdKmc8ECQJr4nirTN02MThHyB0r/hKNPO9g
9ZQ8TG/OSZofPrr47jc1sqTz8IHHpvWz+R9EnDUJiWkK9wKWUZdva4NaXxj3U1e6ZKCvVSXT72MX
4W1cLSO+hD+GXj+Qa4RvHe6VbMl9fVDpR+ZZCDwygASE5vC5CAFirH0DY9Ye6PtMdgJeQTmoFJsN
SY2PVMm3EmfCBrJAzoPbgs4fO1jpTjcMLx+YTlwYZ07GVNeUCErqd95TZnytLi9NeaPYCRzJU8ZN
zrioJprUb1wb5Bs3/SJUo/eCjy2miJObve9zUCTRsRGOEtcV+gA+hXfzSoo0fOkGctdOHdtqQeC5
LT8Wh2fzYJ2uSshbkroRcyQP0v17k6sXTEU19zgO3VNv1wuOKLHgwVXik+p2KnrguFg5YCpgV6Wu
Goz8Tp2BY1hQzmIsAd8RMsNEPzSk7GKVAIDadaYkB5Q3ekCqOkkqwP5lE6RO57qEiUmxS0zxX4H7
lG9iaxwuWWP6g+Xlp1t5t4oniyqnQmsOh2GBHYFPDO7M6K9AvFvuRGmJDlijG8NJnhjedLT4hyOF
TOWzZNzURVMtuXcMg265Uncbp074IqZ5Mi5Q2F4CgwVPIQv51+Uz0br0m2Rk9JISvd/4Tsi5sQbc
hIBfr33kwoPbo9Qwe2+qB3Pbl9jnzw4seIwBRO8Ff9detPTK9s37dh9ez6/TabxtuCgIioCUFN7V
MXsBKgP9u3BqMr82tiL9Q1/AduQE2PcwJ45cC1ssDpppB43nYWvkspy0VlSSdhfcCdvWd22cG1RV
suv2GDUM+J+dC7K54TgenCkixWKK9CJgPuJCuqbC1pBE1U1M41LJOwxzxFxVYdz16RI2HD7iSndJ
Axj4pkZ1p9sc527a/XTCRxjJWR6oIz9O8P4iZM400xp2k6FhL7nq1vo8NQtrEzYewEIMgS+a/AJM
7B7R92a3/qoZRAhq++Zvd3c2Eh1a4EuyRDfgE+Q1b7XoHu8C/qxIdZrZavUVdzXAfrP4y65ejn4s
nnPK0SMza1vKmedKQubOqgB9DkOQaWc8TLMUXbblq3OCZcHBPfV7CHCQejW6KFOpcCDyCpHk379L
DdQ5FZpsGvxhgr42+AYQDpqYeHQAFGzR3NLu4lXkaqPNxp0O+YlMWExDf9jbNb00oxtwkQJ2GD3n
9eClC9cYD/fcaxJKDPHY91FFSXIBbaQOSnF8YUoMx+anBF9+VQB3ABid++DKAAeBeCoTuNx8jBBS
S3PcUATH+7v/bS/ts0XyAhjuDzKwQDeczSrpHCcIWrzI56tcA5jPOE9FMpjR+zA9Bql0YX9vDfR6
D0CyM/bDSOYs1anz9SbsGSLEvFPL/Qz2cyvp7U1wFj3xW0q1mWwY2ZXfMMVYBR7F1vTbqf5DN7dn
dzuqQ+hpePqAijvXJ4wcwnJYRUGRprWrc2Hnw/uFaZ6UcJlsyQYygt0U+clrLotkbRuLLXHdnhKV
yuCiOeRjb6VI+HnipI7NwpKAMtuNDfW+rcdUh+DnfAKglqfm+RQFZcPq8m6ZuMV3F44fG+esWA+Y
tD6aCKnuB8fTZMZyLxdVCHzE+8Bh8tQ5QbfxVUX6jUUyodfT7p4wmYQ9WLULqNdc1wY08eszCI2g
PwRYEbQ8Md+vXxnuN91JEs6WguUT4Aaimr1q4WqqYeaNYp/zGH8d/f/kwFNrAOJt/VzmCXrlD2kA
RopMZ2DWm3kKnVpf1ujjHcr39TwDnvJljjWB3teEkj0UZVJzRtsRaVZrlq3qztMWjORKgGPeESQa
ZkqrGkjugqRzc61K8Ie54HUSkSlvDv6LyoOp4iPo1b/Wz7Whe240umvXMllgewUDXnUmbqaXc/in
frZf7JjHOqT+7MCzBc2T2ZlP8/iE9XOfsZiKXNXeOq99XjxiQY1AxYctP7giBSNCUCM6JJKSVKvf
elIvUCIokxVtyRSZb0tM1vdkmxefavC8YpJuSI0BafqfWxqlBdIbe6oVzqfYwejJz8jnNqWoXT9S
SghhhJEh0HszDlO9PSQcTsr3z891fUatySFi+Qm/ac8TIJZGOSWb6XCij1L4yum1J6nrhNGbOOSB
vI1ma9L4Jl9/xEoa2k0xlAAjkTLnf4xYBY8RtEEfF6U8V+ykNxqvDGtnR9LnvLxNNJ8AIBJceBIE
groTdllsEBrLcyTyi7VLPqsXaEXQxPjQShxYLB6D4jzrj26gVtbcXejgQDzrZl7koGrgik8J5QZA
Aci6xhvNJGl3sTMEu91nmvpUdToxxVqpFKMCS8n3ciJul6c8EQxFpN/C5uEVWhXKI5kfJ8MaNePV
3sxWK6Wc5eg7uKjkj81DmJhk/PHCydPyiQ1r3FeE7mDqetzArvZF6KHlPuATIQBz3Y/1mGWtqGjx
G6KJjo6D+Q5uR0f5ri97ycSKl3NdzLRoYIaADeXI8EEl+mhnaGUNJ5yIeVpJ2rNHFmeOKskfLrie
Q5Ww0Hzd4C9H8OMVn+YcjVRdvqf8QxQB2LGdwX+J+ddIbmgbAKkFYgrbpzPBMURv1qMwRw6xkgdd
/VtlgGsGcp5M5obfKndf4RAQ5piVL/cz+w3wH4j5m2v/+Ochvqko3CbL9zGgGH5Obu7er/NgJx9h
ynZm4/ZUY1S2FebZ52lhAShFy/n+/Te+93DBLLyV17bOA9N3ixNt7G5HgUvn8dCAC1rbYYFfvHtt
Sc8a1qCQqdQl++JN+N9vc1bnifOY0RasZns8yFdvBTTYE2tQG4iNu+CU4/3Gz16dCa84y4oDk47v
aKIN8EgmjwJwCPs57yjjcaUvRbFpitGLFffnW76yoWByX+MBqLASc918v1pYrgxgBZdQJ7zPfiVL
vCmARNPgDaH+Tt53uD9TvGDlJbaq2AWgJd2XsDHwm+ge2HeVB2yoFSGNiGCPH6uHFWdUmU9ZUhe/
ScEJf9Okdt6/6Rt/wBpoSVxcxrULkMr/g3qAa0tXBQq8/yzJCmHU63mdk8XrHdycDvtUgvH7Jmoj
HEggG2YFo3uIuOYryMaE6y4Zg+Me3+fKfZypT2PS/XBxFutvrgQDwKaDgF26n/zLQt3MvOh3Bkge
FSAXHW0vReikB9le9p1aGn5tRrJJe+q3EOGBsQce4m4SP/bReX6HZzO5ToIz5G9OgTWUe4swkJKt
AW/VZ7cO7wlpp8vrszZZvVMbMvSnVMmQHTa07xz1u7phXZWx+G6NIsQLlH/B1G12nyHx7efHdKjd
Cvt73TyqYRWfhOcgTUVgytojGN+DonrjnGL1Zq8MtSeMXhs0tir/AoogrG4pO5Rw+7eFxtPzz5b5
s18x4/sr/P0l88fCE/Ac44ESlqk5Tzlsj7YikVgPwo6FKAHx77kzopazPTACvr2MSyZhbk4xrJfP
3HB+8UdFnIkXP1lyWec3S6fZxThqn62qSLBLTsY8bkBQuoUoxOCCYLTQLdoCGuolMBqQ3YbJY3v/
6G2kKwx2L2Lz7xJ2WpcQn5xgLZt8Hq8tazGPPBU0leOsizozWZEYf3FpFbLLhbR4vdnTIHJaGKE3
8lWvpmww0N1G+69HOcalQnM08PK7JCbgcXpvuUSvJN/rhNOlCrn6PFbxGqV9i5ZSixpr9FWgWAiW
qKshuXWesv/9jzNJ0Sps7vNFWMHIaTmA2BrRbUUBpe+LK76TSQqguLgltxtSvIzwjIKrh2udhkOZ
4cyutdehoZJGH/8ZbmZgCYofVcohqbqKg9w6NCx32alFoqzglHfa5M2GDj0Z8iy66nYrGDcL+5bw
fXg/tceKxiTm0+jnObho5EtyxdMmcKWqwLmkVbZayPjNxgu3Qt+Bnl221/WykYy/h4nv0TRRMfYd
a+jLaAbEmEt3qqyuNrz2wPCx5HTLixnHhbCkBSI3vomDmF3t8VNVaYCMBu9IbNfvEMG0zhEBNMyl
cpN2eDi905lvO7LDZJgHR4cKd1+PVI/zscviB1Hno2+XBq5AA4SFyuLNmDlzn6DJFTRQ/h4IxjI6
XJrHSdhv7UJnOXB/2uroA0we417H/71Evqn5/A5pDy9e5oiSpA+nkmws+fs13NQ7IWn3elyxeKH3
skrmsUhuuUTTDca5us6lKX2iNfyVdBk4dvZIn86/WiGG05rEgr+ELY5+CVAz+jR8G9+qxUqqIfz/
PZtwYIW+eFZa6HfswMBNq/WruaytSiUUut3GzWJvhrKjg0P7n1nvcoymXIntaEjRgxjy4IDQ2RZG
pdHxmCuUA+Qy0S1kJpYFlHfisDhSMtAdFErO+sczPec4usbBaSDl98V/x+oK40qBAbLn6O5r96FS
5l0vUkahMDha8WvaB5xsH7AxXPdamZ8kOMzHAkgFm8TJUyW+2Bi3cStRBnE7UdELY45GYC3pYIMS
KJKlPWghBEF6nbPPdASjlfGueLDeuCZfTAIi58C/sbkYiSZSM70UM0Rewkskg+6bgOF36m248nyd
dboWbvCTzzkDPBtl+5ZWYp5/pq+XCgBph77bWuslcEVajzvXWYRZh4htPZKcjs1jqZO5c9IG1z1c
wmV8NknG+Jt5VMuthWktWBN/R3nwoPndJIwUrAhOhtEAlIqHUllhxYOs6L1ILd/lyFN4qOxIwkTV
7Ri3p0Tx2KzZflssZvQy0Vu5Swa9eqqKfWEutXJ/Oy2tsU+tdHQ/qfPj1U4CsMz44lZlBMCSO22B
ksleLpDF20RCy2+/f9WnmcsQvYkeeVs2gF7a6yAlG5CjX2+zDLarmwiRsI1MlTZ3hONaZK74kMc7
6O0Bl8exZKn7O5CoUT7Wuw2IkOnjEaQfzT2UgMOQDuAL2iZUyaBJ1pin2SoU5dMvf94oFy5NVKjK
sGRvTQNWKCW22vKFVw6Sit/XuzpkE02jXGbSPMRW6zjuwoUpYI3XN3l6aatSy7is8K+7ggWRDro/
2Vqrm8cbUWn2aOMn+tY0ZcleEgH75kQm7zyPHUPGqA09NXucHUtjVObct8acYGdqcvKDYCWlwXhi
0rPcw0dloQgFvzfLuul3VBtBxWV67i4c9ZBU8/JCgg+Q1BD+fyeY+2EqFXDml+2RqgL5K49Arhln
JJR3QXcqFjpp3SkP8l7vu3yWUllmzinv3fe4eIeDihGuWIfpeVQCu9OHXPqnCCtzfStmrMCq2flV
moylywE2hbnd7TyFQSC9ST0uIOQyYQYb1J+y0iXrnW7al4qvtpTI2+5Hb8MPjiELwHXdddRIp3T5
dqsFd0jqbPgNetRcqUyEd8xr9iVsWpsgB75rON9DgFlkNTjaWYfltaRBLbMMBZwhQYSqMd1Iji6q
jytO8B5xsV3Mg39TeViwywpTIlVpbbhRCij0E4uBAYW5HM18y4Gm/gzi10lGaEr87cGUdoTWhdwf
zSx58cFpGaAfmsYO6h3+bOw0srCjNxDD9NKUw48nnV3V7tor1RdYLOhMDLVmnq/NCzVbtw9Xbfif
SgpSPJj+Kh+F0Nxj2nehzHemw+D7GbWge8NCOYKzEJQCGVdW2+eUg8AGnK4RFaNv4VwKAq2scVgm
mdzqu/FSzAGnPqrejJJkSETI1xu26cYRzVXRmaqoFiGGPTXofN9PzVKpyH1qTOs7z9680538pmGJ
MZ7EysB1U+e6Xp2L6qxofv8+bSa5xVTh0dEHSJupYGzw4L42nn3QUrHLTKdkv4Ea9Pgh+VJGy2xe
dBIFT8CxNfxj1Dbb07PvTOKkiEKU/EzDVNUGcJXDSo6DyPCLHyNman4usfQKmiMWwdT2ZD+K93/i
bL2ik3tyBzNnCJLoAQYNlwdaL07fSxTEjQG7Ybqd/QZ8q4Nk8X1DMibbIw4H+tmWGPOgXHkQsFSU
JPf20a4Mx8jGNj/ru9RlJdsssCa3ykyWMN9UF01jrNNYI7tb9HK8MgAFbfUMT9TGlxNCDxv2lh2q
JQNQ4/hVE0zfreRjvJK9wKekw8K2/ysyf8uJOM7Rsmc18gC2rHM4fRlD5tOV0qfwJKo1zDoVOFZZ
OvemvPmOZ6uUbt7egQe6FenPoZUYg1Rb3APhBb7rx0YVXtKMytoCBxl8fyR3RLPeez6RA3ezg+kx
FhRxZ3R4lcnPZVih6u9si0n2mVqifqMbJamcuGkKHpNXW6EuXsfvCIbK/dVJP9vUQeDLDGzwlz/o
yt/+Z4dB7RkUnq+6yQcU/EkcqsIgTRWN0ksXdzCc2T8exYAY40StIP610N3K1dSQVRJliNcIFBoy
6/A915atp3sMqq0ekna0zjXnICKLlM7W8aJaCfybME5p+q8B+oZLGQhCL7fpRw6zNuuEuzgoFXF9
EU9vOOcfpqhpPmmzLKqxy1E8ig/yxKBrtnn3qub6F3frmgfrlQ2UF3TgC83Pia/Ptz6xPTZIZu7q
ACU/wHTjB+a3HMg4Hp9bBeGkOxszsi0e3pDm9cF0fg51PWsl3nSmVzL+BoZau6VE0uXtFIGpt/GA
/OR5QlWnJ6o2DLQJRCEvldkGL85hQM0DpnHV011+9osdj76kWZHJ/Kx7s4ZDYziDrZj16fNhiX3u
mlABL0N3dhx+ofeyRTA1oOAPkallIJfYIF8/icsPphFdwJD1RH87YADVtuKHBW2Eva87TZMwS7Ax
U28oPTGNdmUlWvsCa8TiWqNfilT0vxU0sF/dtCzqtcNqRxD8rWRUJFu30zDtwNbaLDzq8NlF77wv
yzml1dAC3ioUcGSI6d0iqTPtvrd2nwkQsV1nGqPqWDrpvznef5afgRQQmJIv4remBfMkNmWotjeE
S/4LYwxZwJRxILiwNaBYYovVh0f1TgYHGA+Zg0kUyKX0/MXTAdPrgKfFJafzQ+exJ5s0KqxQAnrT
6ljqoeEVASGXY7yZqyYrRhpNrwFvDrYauwtX6KW1b6EGGLJMjqGXMVkS55gOp9Hvzi/5QpQh50B0
f+btLUPAfTMwMHnraF2mupnI0nyKIF3GOA7PZ7V/qy5uv5v3d3VYhAnzrYhrXJKZWzHZL4PAcLJC
f/Lpi+LDxmpBDWCgU4MZYTBMzK6aKF7vfhQieZXO1tPk7F0rflYKtVwzZGL9S43XYCzd8Rl7ucvp
HDPd5UNy8gQRQ1w7ALDsVhbjXnpo28HZV2SQCIca0fIw+/13yleMv6j+d/rjC6MGOTMZcidxCMug
q92bhPa83uH+n10TetcmRfeY8BK1wk+DqO7Hp8Vf61lBVYZJ46I5J7CsiXXn6VTTbazGFiO+5OE0
d5/3Y1MuDFSH6NJJTlrk7jESLsYFpcIz9oBM6+kscVq78PhrtXhUL0I877td2vScJvixX6ktbT64
IVoFLxwijWyQIxQP8n0xckQbyvsdf+0mTFTs844XQgBleirnIp6Ty+JjxNRT82fl+5BGQkWuhqlR
gItjIpHXxBIEXbm9o+j5v+9+0ys+EaZEdbWITK+v3MfSEiAlNdkavmOTVkGl0PaYkk35AIDoK3Eh
zWwPJEpMeKbybeMfylZIpkTbWhgvWEG44lireJ7WQS5iMf6L4HmsPstXeG+xIqkYjibYkTwdX+eT
fPa9Pu8YA4Hm2JwFphtbQDBGi/I+8oFHp40X3CPM6BbgfjiyBht4/KKoNvGvLKo3JMTlf4JB9RAQ
Y52plx2UInZehBB5PPgjIV6sTYnzf9TmQdqjbVncwqAsuIJvqQpKExiZvlCjrrMLONo62/kq3KCa
fYkPFYMph9CjPJxLLqo+KaGxuEdXblOSFAoGKWONg8X/ogSCsAPLYJG5xGYYgmYFPIUzpwFpZHw5
qAP3Xm+8ZT3d93WKI+qTukcy0e7+kiqsjEa5Kxvy7GVdNnB1mA4lpVRy8FxpRD1+PnUlLF1G2ibu
Exqq51nVz0fvGBmuKwQ87aAtxa9D8Ir5TOovI9/UmlhgXnFlx/XAd+ku1IaIE44xl2vz1QKlcSVf
ZB/gUZj8uKZpeU+YUhaRuLU8Faef7L0ADd1bjTBb3E12H8pbB6za61mUZCgL4+q+7er3DbNhzgI4
64nhcWJVacBhK1UM/hR3njcUiIgLfA2LP8Ed863pbCF6KeSb/0UJUjoY1Pywd+wDhxImwCsV3hYr
Rl9wl5T8JTFy+85GxjeIyT6GTay+hgcE2pdCx+WqZQ64VvuNuJrxmTd34j9/ulyvT3hg7VbfM55t
BUQZgjZYI0AiBgLy0wd7OK866tzG781rUhL0vqoMY8Iw16RIbgbn4+48qZ+ey/fvWUKyTjUamhDu
xFzZyUs5yo0RmLKfFncCD9/rWi1Yhpys1FYAz9m99iCGuZ+ehhFRlJzZxn6dzYQhQDxhKiUUe2qh
vEmPORitZcD8e+n1/CooBqoCyZ5FvFa9hWmAJvXlhjAWeuLwxBe1RY/Bj7X0XgAfO8DOiCDR+njg
c1DmwuNuCLsWHwFe+D9rx598ayibcxT163T9Mn96KCMNFY1lgAha0vSlBd1LquqOzojKf+gaDAoT
HAc8lZeWj8LGU6CItzpYDAgio//BwRI1cWDDVbpGmzf317nvQEQTDB8y+oZNqPMVFcPvjhOnrcbT
g0kIArovyiXYcaaXXU7/9sk0MHOnQ4ebReymB7vg5an+QMQRWoh+0wjCJepa9fvAN5QeXrBJZG7H
h63rFyhbHdBiK1srpnXHKyB17ZZppRr1vFC/0TPSPkWuBeFJmwlZ0hnj3dK/ePSsIAB4QI5W7Gke
H2kLXRGIu11aWAKxe2YfLnCEzLxHidVw3DVtWSWIY8D8H+NtwsBAuq9n4rIRQCJY0Qw7IviFmibb
Qvr6YdD0BuNQTB05GiLAUkZScLdgRFCK1/F/UybnCTsXNKzeH3nLL2moTY8KatPwBJNZUcgWBt6m
D8a4hTF8aDiJ/E1bcJpeK+E8M2nyRcn3q6zN63m5D3WPRT/7aZqaQrvqAch45yeVgBQuGHLZQ/uN
/wIkcSJOxQGnd6jS8OLg9MIKuHXz2iibE/6+8FxyA/2woGR6qOh+D5Q4eiRToLuW169NLLHNhuRm
QKTzQSJYAZfsj/WXXOI6W1NKYTRa9q8+9XUFrKJQFmHkHBczTixuCIr7fY9oOIqcBtcvdKwIjsN1
/nc9MGAMmX2Jw3G1VJ2PZDPCNiSkbB3+AGe/vK4Dw6F9OS6LdobJOepx8CjFCLcqzH52ii7k/y4l
N0MrrMtMz1HV6l7oYjFcDlzQMuw34BjGZgKOzIN89qDOHMeM++35PpR+qTs5awnKD83f8+dV/eZZ
9L8FNQ7lmtl1MuaZFpB39zYOQXiHvQYWK+CEmwwqKzyCij/47Q6B7PK8rDyJ5TQXQ1OCv4ttodhT
YPSw/j6rhuMM7nmXuMnquFNWxmiOTLXE75uf+CsjeC7ZcTKdoxQvZaKxkuOrzZr102MpHDvUqOPE
rUDdJTc6BicQcUR7ADWz7Qpa0r7+d+sXmEIil61bTbPWH7eT6bxeFGp1cKV9SuY82ktveXeddTWb
4SqFcHF8yru8hFjr/edIznKWaEJH2HgKs86ldrXVmDMkeyc18V2xcYjgGw8dGWUlyc4oUTq5Qoii
gl1z+qGkPhD3IBg6G9JstN+6YaSqNv64xg4gnBznUkE7tyIXineMy0EDJ0DWELfXfdJSmLC9p+n5
iKhMzvsVRvD66sWEnWp9xsUrzmR7C2g5+VDeB+Q3v4JTRY+qHZWgiIn2Py5J2mvCpTg4i5YJZr7I
MbXaUwJmkZrHwjf/3Z/JaiuH7cXS+k+W5fh/uO4oK6FpmaXcsNayQWZRNSAw1z4jG127Q7qP9+m5
4HPisKQTPLRf9upBPFoYpFu1toaGKiVde6yl1/+AvKeQNJ789FyuzsSEUY+RBDhjX+Q+GuSDcuLY
0yQGsjvYa+gKe2rV5UPQvp6L6VQ5ogcO21EnxOVeyHDVWn9FnGCTRjaqaUp9YW5VoXSWsjG7TIWs
BcJ7kCL16yjaw8NCvByWIQzQzB32oILbSMJLF4f3h9B9E8QwHFZvDRIy8SDqsOa6pDlW3CbIv9kf
7ubbMIhuMIxFTroG0WzZyn42OMQSQj0BAQlFkH9Kuxk2UezAbNih0ajb9IH6TFvInorVYNlkT9XW
PJ3nyyN7FKxr/3avyQOIGVxQ+7rgu8VceAqYaJ51MFHsQfmP6N7xl2SIFgCfjJxWAxN7l28eo/cA
bn2BQxE2AnfTdvvH3z6yikYPBWkKCAD8luu5zXfsLwsKHk6KFcG0/aPg2TIXsFC62tARBg2K/AR/
7EjVM0//VnkU6NhRIhNSIU1a0dT5oGDNhDbKMg6oFHzTbwUhm9Ibqh1ek+fMuas+KIvYJJA4PgI+
3aWR5xjqC/eofJez5TRzFMUE5QQ/A1QCBLI+69Lo5dSP7AFudOqsCb9iBJ5GZzPbvdESKlKjktU5
BORL0OJgsPqFD1IKncxi/vptlOGVX6T74cp2FnPR9Zq5OECKsAaQoAZDCSWN3WX0uH7oIWhEtn2O
vcMBKhUSN/UG8lVYq/JB7++Xtro/WOCz2C+sbPR0PeFa9TRf3/7+iJtCULE74634XNUPWQlLW/9l
iXBuXS+O6yUAA7KOWLvxJaa0smleLk7ABleLPNjfLgZ+4YNRf1mWvCxgp1AhI2Ctoy4CSu99aqSU
LOqL2ouGXdHB74jKd8hDiW4QMQJg5UKLg3KAWIuX0wDlggI/+lFYf4vs0iC6+T7uqkZA4KjJ6Pd+
vobEOHCRepIHMLCAvwkbe7OqSSAYO0ohZFcJXyBc4bY+uFbz4hF2dWvwY6Nh2MeoTmIol6Rp9pz7
Nbo57gd485tnDPi8N+GrRMTLPxXZoHj4pC+J0tR7hBevja0Kapu1/3iaVUJrCXhFaBgXj+1A7o6z
aXr68iYnuywZdiRSdVKzeS++exGfmJ5ueFxemDEM+AT2NjEr5n/En4TkqEz+5Upw4Cm6hwQoruRd
QvarXYWGkRMgsQjysT2W8aMGbaE4AIvOLImfDinlPKaWhIneoJa5EB0Y6LUfODg991rotnWFXt/O
tCjlnXYQA6IXWLB8SplLEVte+c9PSvAGCgdlv4rx4QfW5/QSxV1qypD9hFarVyBu0ieQrjouyTyI
B4LFVe2O0QvFQX74s0ZWtkRBTtDDyztUW4oFRHNKiuW90r9kwPQwD6RH4WQM4l5hcpk/J2EogLB+
gnWQAfd1jMJTdQJB3s8eZoGF4qFh2sTQiyp0eCXXaQv/R1t4CqvwSZkssisGGwuRTBIJ4otieIY1
/ERr3C7/mqV9+8ArFBK9kBtmHx6fuwr7W9PrFwYwn6aKJeS1i0Espy2nXGu1N4DiDmepRs2O00/o
LdqJeCeYXgCiCv17X5x9246ZbHmIeMq42Seo7ivxdu2pno20o1bJBMgRJW3aLwi3BaSDqPYl54JG
ieV6IKu2q9OKpk+LDNf8HDRIl+6OwPu/vysoJh1v0pnE6za7PayizpF4JdE8wuBQSoQ2/Aol3Oox
5AKgpOwiFKq/mY1oi0ai5FMQIw0GGTvDJK1JBKUlYFbNMMN0BSof20WUbwl5MVAUF0bUQCx3XAfg
yz9XNdMndxGAbM4t6s1/M9h7CEDhde1pbIvg/n5uIKnoOXB4gzU4bu1GVsvVi1QPNv+REiPfzDi7
RtgfbV2dqIz0d+pNX3nqY9AeuGcpvpzshnXItPGT2A4mPy/eq+SteSTo4FrF3jPdQQu9G2nsFL74
PZFyQTsPiQP4F/F+3mLeIPIgRQwZYKNHVBVjFV7P38MdiQvc/s1azu+wLRbgrnKREXKXg+ABKlRp
BUf9k3poYOeUqdjrGmeUwRI/ABhN1PxvDHr2LfxgjU56VWa5SgYCNLUd2H6n287KTMdgRD/y3ctw
rhFsiwwiCLqJv+cVX6h/LLlTkj4clzPdFR84QprefUdS6N3roxqBrlGa12MsVoA+8d4CifkAyQAq
9uujSC+uPyGYhR79BXRhBGLt7kndyoWLf4lejsCOIEzUXVQMXMJ9HPwLZHHmHC0kMSoZZHLyoRZT
SL71IEBExi+75Nk/+2drhqgov9bDH8wbL7dS4qvrDOm6i9ZlwB3fsAxMocYmIruL7uFjXKt9zGe/
ULQe7S18O/r6FZHJShQcx6GsDy47xjdU3giyUcucLzar83+rzYAQil6F3WNDbngjdBGq5Ys4K8EJ
4obH04VYaldCmaWf3HEjoyzO/9/KYlUFeYZAQi3njUts5X98n3HU9OsbOi0Ri+LBGSfWX+pQsRY5
Pv72UrIWZNGHWxg7ZNFp4wCMq6k3TF6HOntsTvbuYCJgx1RNn2PZ1+0tLuRkXxpRKhUdhD+WKztZ
qyrGsRYLoMtFWRVrZjqhQyF8CuaDhmJxgDym8wLVRnhsRveF3mSrHD0AwGgWqLGii5044toEyxAk
sCdL05HtpmMzCCqaTPSTp3hfyz0Uv+Ouy3760oo+DX8UrPFbzdP71JwQg7wr6y26jG3GY/uaCIo0
EfVxTyOPBnmINzAu1TBOi7aapRNaReNcdJX0ghtS1+pLSREiQxUS6qzzavnj8oLQkgDqqRQL8JBE
G81IGZpVc8Nm3S+0ovk0ha7clavA0P1bAL3ZK2mv/k7n4OpSGQT7CZE36wSLc2sog0l8xopoMoRY
/lfqFYiKrp/JU6jP9LZMT1iPvRBf2hZJgUiafRbHGElmthO6Hq++CA30nJ8e3RJjfNskEWq2p7EJ
9ebc4zwn89l8KQRWhrmXcB/frUrgJKV84AU8F6lKIfbIPp5kOuuA+Xy3ORTKL5/1+V8iQ3RmeKKd
r0Z39AILsQh/N+v/+XAva5KyEF5A/Kz3Vtz9YKJ3Bsu0FTZyih+T/IDVRXx2pBLiwL3IK+ueifJs
WFjpf6s5WEFW58BVLoEYqPxuIQP/+6kc6FChOMaajpaXiU+s9iotoi0GwO0hBskha3+aAs1tA6y/
4GhoNERzgWOMCqdU+cUf/IFbNxHRvFes26+TE+TuRVfSyziuR+e7LERmnLY335TIsQT6LukPDxNE
PLSVxkofr/0Ww502DRdvvFwEXbhSylAFIBO208TbqheF9H+r793WBGrzJyddEen20VBCWQQpR19U
PKo1l8cix99n9Qa4Gyt48N02KKFYe4I8nXaQDChqv/Aq/jAqw33Pkk5ZWqdMsXSJzp53EAIxZsaH
SBJei2fxh7owU3TDOt5v3n9kSdYBzZRmU0E8ND3xLJL7qaf2zEXKiLme+wuLIx32UoEjGfQKS98g
e9BgadzNMMSnNNo9WeZAANXBYJEyOp3HGnWjnrZ8GdESGoeixhgGTMqAGmFvzcNKzqmeK8nkWMbP
AHmK9pxa3lRAQH1vaCzvaOTPoztQGD9TBi1Kkh3gAxLlGRmeqENl8F4Gbo/yMSUvQBo6XXQpsbKi
ExEMuNHxfRAW2QJ2jSGCOmg0K35kYAPriNLWa19xNRdyx35jr7/2lwuAF039WzGJUrbOaSg6R+wO
cKqr2ZJcANueB9d+jWyPOjiQybwE1X/I9+Bj25L6OIxvZg1SjBAANCvTUIgXQ09AtgNAc7S/WGV8
SkXqYRA5E2QOOlJrutomAXobj52EKFzNIjL2Xs1zJniCO32wLT3b0yR/G4gFjCc49IfVoipjaB/b
3/mqGWw4AR+UiNa0rkF9xj7ayu+dYbPwbCxL6qhaAuY/HpBcbLf0dzg1gzyR+8KIF+rf6Z0t02P0
9Yat5kY7YUYGSl6Fc+Pjx/SWtFQyMOcVda27slQyXsodMNDveXWw24buMwrTGnnDJBzi8QC7y0xI
x5rdbi5pM0BV5eE8Ul4AyM8+E4G8OkG4A50N7aEpC5cRCO4LTHGuCh6r2437IEvB4AnaKSb4YzCz
7kXiMglYDCxgmexwIOtYpHQ/lAQislY313wmnLvOOlMSE/aVFV/5a7Th5dhmPtHk4Sw/vSbZsXmX
OZyUxEOoXMVQ8cdMdjA1xMQGMP7nAcP0HqiYp1XjP8v7S1V2GGosio2ma6NyhWpJhHQRycxrPhP1
PgIBmMcx/dkTecllxcDrOhssF7MnTYCiE04IE7xialCohtVZXcgcc5kYdW/Ff0tlOyBdHlw9LKyS
7ldvl7IvNfl+I4fc/tM2UrbTagMcyYN1+5tumPbRGK82PqDKygb8LiwEQV8xZjYgq9XbyjvYCppV
88TUw5Y86UMX7qIKyPb84YE/5AvseJqHNNSKwGaBx7HyYExVvg0fTPOhlgt85iRGq7tSIAtxg5mv
uKpUHJK7L1nIL4kYd/QoSr2YEBE/YS0az8Clf/ONUdPaHVIa6vqwBoAybQeQ8webQ1qLc9xeXrDr
5aftQirq3AHwR4P9Ewk2evB+RMUnodoBY5fSfQszla23QvBwXN3nFcSIDhGam+SJWf7aNP8qGCdi
Uog0sikDPt7EJUegJHMQM6XHk6gs2UhBwm/UtAXYuTy3lYVWqY0VKvCgxA116JuTUVGT3+YmvRfj
FRnN/jeETlJ5sc3WaSnMLZTZRfzRaPjktkaRhCqelkoGsDWHKapd0AhGx3chdTJ6lj3e2WHA2dYx
CueHnXth78fllsZHpKjcMoINqrLWmGrEHM8NAuzj00znKXwJA9tduwjSZraii/ArebAtNdZ5YAKy
X52uT/MGcJ/Qo+RDayYfLCE0ZQTojZYUdR+C5zqfM3buzb46Pe6TEF87cHF6wHZJ8KXdxxXqBqK6
h/wTjGjwJC/V/E9XoT/1UZ1mdlpDXZH0rwDjjt4DMRz8oGl9wCBSg9+MnOdN4PWcFQPRM3UQyErt
f6+RNfw85TRqiSf6MHZyJ4Mc91ePaFoN6QqgQM5F1tum5BbteSgf5J6JYPCka04vVPz5UzX1r5hF
G2FmWbUb8TDUmBj22oIbfTF4f65wbI6kAbIVi6Y9jDy5MwQwvEEPsUO5rRxciZK0zWGyGtwktreE
lGOYjhe+OcOsT/tpqCr2fLkalE+Ej/av/dTQqlTYY7Z376Zu+YDunB6a/uBpUslKCQuxZVdTApqm
vhJtp/HbEzX5xBXwyCHp6gW7Ib6RuOngZ6v2QvISe8Dh19MmvJaN6P0GC4xLQ8JjJ9574U0lizzl
Lq0iNLWNHRUYhnciQgUj0OSV78aaAa91OdYiuivvFsJTnkbxlcMoiWhyp4lYyg8ZWs0SYN6AaGrK
8slwH7ufIxBcyPrMOl8A11Wa/3jfKsz+qZ/WlTFKTPo5bpU/zmc5diu0W0d3m1/Yj5759uqbQStU
LdoGYcyOIkkS8ouGXIMt8gA0AOlANLxBtGUCkJmd6MOCMiKDADE1Xdc7HhgmEcQmYkumCapI431u
e0SdbRS73bi9c77/9TXT6NtSgjyPszhkf3pPQK8lhZknDHz85M/Bb3XQmc0HCwGAMmaUSiy1dr4h
jUmXOu7qpybGBNwBuIu27mCEltRDjMl0o7QzJdx6EXRZ3SRXVCnFgTN5CJwkMuJAKIa28BYUMeDI
m07c5duSe1EpLFzQWxGjJEOrNxYHBGWCa1YSRgPm6o9t8YCSH+yh98RxGB99vXbdR0RHHrxMi+YG
WgSDYohUbG0UsvsJhMtHzeXWWL00zw3pSdQERimMu9P2jHt7h/evnhCN5vY+c7UibUYQDmdIcObU
FGfqQXTYkud5O4Ec0MQaXJWB3px2RQS/fLHE0Z7ITbJGiljfsXARcPV/6Zcrel3FLb8wPmY15J/U
GnF3dBORTcuS9u1GKGClbaHGOUuBQrkKsJ7SAIfM6dSyzEYwaVcuih+9YSwFGTUK/r3NJsHIn2UC
9OZIZMtTW8ul9b525Nzause6Q6gIoEfV/fTIJsg6J+pC0Kq30bdh1tXFLH/uL49aXfHusAJgDEoM
abZmrYdKQHfEE1N0U33zEuQzL2IizHOEeYe5clOSUPcjKerp34oA91ga+LHIsAk2R01CKCrw5TNG
CHokmxLV2pRBjSg+TMV2wx+YZH4UDJ5kT0mw7yBEiHFHou7RzTCYcCWFAAQScLtMTccuzxW7t8Vz
hh25Yx45E9+Zy6WezjMVLMY8r0sDzHx7JrYAOZB4K+ViUJKqGMO1rVflIn7zt1puEBWVdE0U+1a3
YswIMasmA1/IxDgoJXJbKqEkBS2+rqtfHbonnVrOf7PEjc/rxmDdwBNUcfFuPQIRR+YsFF5Y92Ye
C9XYs/2MO+XnjorI/Vzvn45s3D8JvHOVO0el76QYyeOGC9beHSSxTFB6Ww/X0brwqzqJtNLwMuJ5
Ab0wH5n0DsVLWaBsC6GytjA4rcqnTEdRdGiJJaggaj3lOPtSn/e8K8q5sRFsz/oEQHGMuJ9/lNlZ
q4nY0FqqrXsKB6Gjt9Lfjx1/sGcJEORnEC/EhcCmUJ+3a+rC+CchRLHnzSVuwGk2qBahmCb/KxYL
8IchIwl/r7fUbyuSnjCXnVrFtR0LI0NJdY6M0Flkxsa0D+tAQGljIZoPtEbRHR9zgLhYboBqJoA7
1S9gocK9XNbTZW2ZkPHDbEGHlS1OANSzLyCMXdu8SG1a6HdRuDHomkmrHaVal0D/67/8mh8blosL
k8cRF100hsevodcuqe079MjB1Lsrk02KI1/Owe+ai2eTp+xGT3xICA4V0gCzBIFIXaGIKLkEVoGb
R2D110o9YLEMiE8OqWO96tKqIkrZ+xVxKHCeJGi91MoAgZgMq6ciqnZBjalxiTFAwBDHublLazRJ
bQZdjn1bTRSXnJpZl9W0u1ZmwD28w7g7An/7cUOChE0I9A3uZvx/FOqwB/+CU7/Rh7o85/SCi9ho
QQHKaC5oqoLyCPBcP7MR4amPM86QwfVEupdaGafy/jqPW9SYX4iHJnkXspG1PbR1ejxXFcqNnYLn
tt0yYgt1pWlD8K1kNkS1b4PrQdbGpp6RWhP8xZ6RezdxeRCxMpVoGTWeS98x3ummrjjIbLM4IhoL
V6jsq6nNjztYw6voGq3ImvPSCdUwld1dVpClBcxO0xmB2e95chv39eEsOuSWECZJvE1HHtceVgKk
3ZiQO8s494BlaOJQKye4kYutdS3mxjrbBokOB17qT1QnFe6Sa9zdahgzZNax8gyjoNvg50DyYq57
IINn19UtaUxiaIK5+AaHrkfjva4N96BUYzuiWM5pLSU3hsMFLRizwBkIvgrlV4vHiRWOmVRPjYyw
QPeES9pnUrEX7M6pVxpu7JYRS1J7hFwkwB78FXeXn9SGCKQb7+pvmpc/bvcpRNSs6B/hARK37aM9
aL3kje8lagpfgtYkxfqFNkijz73cnLatPg91ii9XNvH17cnAmMqCgwBLJpCvtc+7bfLjWso3Dulx
kQnMtdXTfmTT4lxbP9ob/E644SxhrVB263YmeFgWEOYGNKkFoOvGAIoQ2lczYWwc9m9VDwutWuvU
rg7nPxaLkDq6ZuRtfSc2gJdmvT9Fro9e9h9p3d4rK4Tklp+v+EfhyyCzhtrB8j7WllrLFI3tIpvo
L3H/g2F/dV3VfrufFZujeC7+aGxBjLwstzZK/uXddNM93BQ1c/88Uq1zEBqFe/rBP7cwVGDcM//S
4h6XInbev5QcRkp2pUnFU5ix/wXzJukRUmepVb1+qzmEcg5vtv+15/fhAlblSW0ehvDj4hMbij/Z
M2fI6nEd0EHgbIUr3C+if9YuQPZZN+StGCzvaOeypG56/TXs70qqG8/6HQtzy3n83JWqhZpI0M6o
cDtwSe8cAWqu1944nZbY1aZon6jYeZjd9sigenNn/fxI8qu1E6F3BsZmsxIWjVdy7jIFcvjsEUQe
WoqfpaU3oKKXyGORQhV4gwHDI16hXl7htnRQnAF+4c+y5q/76AJ/74zRdhC/M4NVCjh2kRWK5PZJ
hFboI8E4V5vV/Bnt22JDVsPLNWJL2kg/cUs6+9y5xaTt39qHdS97wVWqQHlUWFl4s2S0gkeESzhs
35WRp+mdF2M9ZgQ8fJ/9inFp9q6ed/7DXlV+DNhLdwvqFHhTSvldvN8Pdi3KRxqGBJWV13lARk/k
KgMefZn4HLR9+LB/wOf/uNAmfoTDEmETOPGO84VLXepbl/OyGuPAsCwQrnRX6ekvpTwTrJ7pfmNY
Sd1LSPDrsG1W8q/IHXZKRIAEpEvmROqnPS9e/xQGOq1fSUyqKE25YwiUa4LgXDBmGeyIemayHOmY
h+W7wiUOTiwTnXd5Liyoz/ZI8eWdm4gkfMVVRvotoJWcOgmArwrCvsQE3xkYWkmeaGxiF1dKsaRo
6oKZcDv7j4rtnlHYSxt/OwzgSoTf1RC9yZ9Z3S6yOE1mZ5x0fIZIVtm5JNdKUHtjA8mc7+iF+BAI
4uWvmjhM/g0xwB7MTKH6mb9pqhAqzNA6icnYw+TQys13zEu7cwXVumBRIr9aDesZhp6GcX7CgJP/
L3DsAuaaNAMnA3WipOgGTpE8z8ibS+02XdX/N8UQTNm5Mq7TWbjCojGIkcs0Vp/nlWHIhmtWbV7K
olGS99/JeYn8A6nlqEZDYAw2jfaFKc04rehWU/uw0mQKq263y4kJ6wBwzMfGFY1bVd5C8nWFnFTV
gb8Gb+TVgrsbTD3Jkk/Pyu0DzNsjyxK2l6j2DEG0LZ9jfGpP/O9KStDTflKwhx8wosrvCF0fkO1k
Z0GVa/ZuopmqPBpeWv/N0C42Pj4PRm3phTSspf8snmTLFOk5ayA6c5we7f7Eu9+u9DYVObI+8ltJ
in8ABDvrcnleq0pqEwwPAhjEl3oTOATsQf4pPzARK7F9F+OSd23Cgg+VL39O7mHJVUi6kSrKOG/b
0S9eOnLafnJF715eTlwdhJciWZqaT8pqx2EEIbDqk2Jq964gmFYlD2WrqS9r28rx86CIydIli6ur
ZttyIV2poeJK+BwrEJHb8UvJsf2yAkKtUmYIeiRGkmRc5gQTuTLGU5bNL234uXQ7COeRChH5uca5
ueRnLnOT7x1FSXep3ljycUEdRdB3etOiFCVTqG3uP7aRMcHsOUGxCNTHGco7gBk/u92qEEcIKWAt
Rl6bns+UASaSXHdc4vQXEdjHRWbT8jvDuc5+6MVSwb6SttthHzfYCgUv02Uit0MUvLHHlVYcK53r
2qyxGpI0kBnNPYUVGOANMF0H0D+buUiyYof0A2SYKJsujiCrauH/1Vl6Qvcx7J04tW4MvVsxPCxg
aPizZV2nT5P8K7oQwi++dlysS+5YNDyx9FDZj1Qf0NgQw3OuaK+b/HFi8Hgn5nCVvS4h1um7XzkO
pU4Cjf0VUH61hNeALy97TY2RaR4BJEpEdjaYMuw0E0a33wFO3uosaGXuk8f1AT4014YsJazqgX0c
P2GjEDm0Lk0RVBSUrljExZ0iNTHwbeWC+id2Vg92aoBBrMJ9ptAlTKkw8kLxBi0b2T6z6LkNHC1N
WORf67j6wRrV8h9lV4CLpOXXAUtoqt2VHN69eK2QBTJ2EZnDR7/oprH0AfbtDOfJCCV+kCQt2Rnb
emPHHhbq6W7G+pVn/NipDHhNYkFsY4ALipfHqEOpDYIdgWWO9KzkpprGgsE07t6fIT0Jl5dbxUpD
UaQTMWedlLNCu76XF5t1YFAo5768sIrFQ1+RsutUveGdsgAtV4Qck7RgF4NhpZsFTBhZcM1YfSnB
sotrEmJVBf3Y6035TAgpCwbJC2BzsHbeJZII8vxMtKMNSU/0ALKjTb8v6PExpy3fYLNelF6dtLXf
n+tUcqxBzhwZXXXg5dOEY4jg5D7c0+xFovPIE1Z5rbOB4ZqYnT5XOU2OA8ycEgnP/wMuXewioQDy
OvHzhmoXrk2UstNlc8u5tr+cMTT43UecaBT9Y8OOfjGKhE6Wbbq1Mv4EHCEZL/efZ60peT2nYJew
i4n4yvOd9jS0AGgWKAyeh0uZOC7BClsMzr6xLGrkUYQh1tWQepvOGJmcNEexnPmZNuaLShqTZXjj
fvqcyLhYU8gaCMHm9ZFgCqIHvpW6gPOMyl6/jREZdudHHxSUuEB2iRNyRPZhlqMSe5CddnEWYxkf
3FSX6EJgumJ73sIOlC8cxn1mCm1J3SHT9b3SJgOXD3DhuPEEWua2qbtpVbLNR2iA66If+Zt5qEkS
pLZLGY43Gssk9Yo3tYdmafN/VOdgk8tjTVK/oqn7tWM75W4hNnWeeYUDhcS32UyI3tXjq5Q4rlZk
LGtRYawPW+pHP9GGnMCqLcRv1MOsq+xbh1rN5r790U1vpSetvTYFZ3LtShBbFhykMY7B/ItWDl21
QVsMKnWqU7RYB2qUxIM1S6QZBUs5eRHTMPw+UC34Q1Vkr65eyHwfGVc+Ag+gCM7GF28iD77RzbNa
+Ny9Ku+d8MguIgbWKt+AS2q1Q1nVbb++ALrKgf3Jg3g58vw6DTzOHjzpys44FIU2rGScF1onns/+
T5Ht7SCW+bNJpm3b26F5doLxhKseMM+8ASsF729fE9GjkJPjSmBZLahO3sZ1fd/qasCIWRVjbQE6
hMNZ4d4WZdz1yg+VQSmd4YgXiKHpFshZojpiy2u/GuKb4Kri+hE9jYWQzO5YLQpLdaShH2YsmA9M
NeSWvBcnb1Jc1mHl9nT5GV0U89Nh9vXg4ikej9W2/d399zYG++Tr9hTQ0Z3B6yGn8QybHtfriC6u
4kmByDy+oU62NqSVS/2AeQPTy94vzZJAOaV6SAZ8FxTSQXrcgd3dmpCe56e2lQCJCgYyg58bkm3e
73z85GIweWIM37vxBkGMT9JpKmjIubUcXa/CNrwU6M75Wj7lRm4/6Wjhak7FXbF0xEPdgk6ZHHTU
4ia2XjLkZGdQNxC0/hWjYjlVwRLDTiV3K8xDxOt0Zc7ZDrm+cBLC2n5aKeKOZGNXrmPrJN2xS3+F
Vdj6/fqYcbY4Ohp8gbxYlj8H3o+y8iEb/uoeUg8cokYfGSAAp93e2nR/H2h32RRyEUjzCwoMA3RZ
d7g6I5VnzTkist+C+Vr2RVI1z3W5xXMYh+lN3Va7aur/VRfOY9XbPvM7KsRFJK6NrgXZp0aYH1ES
HOVtxXvYGmD6Is3A4eWx2PTjo0XeO3b0G4Cf6a1TLjZ25NB9i9QFBzlF3nppR6ap3L9kj32dS/S0
slTlE0V8Epq/tZZ3iTnMZ2rp0a8x/PlLiaQqMHfjtaFls+r2x/EcsoYZZdwq6CBSbniVIg6AAPoC
71qtHMup/p/WnV8ypL+aWg+zqZew+ub2Zcrrhpy7nz34SO1ICI11xbuOTWkCTRMt/iuBATYl6IJ2
PkiEegMObSokHvw30are/wxiUC9Yz3KOzolQriOaFPpd2Z4W/CmqErTgKfS6N6eB0Oezklf+tIDN
gQLW1oDbPoWdKQM3Es9mD88FMoYdS/gkOo4P+U6+ii+oKqildDQwI3txv932Be14TFmVuUJMl5YZ
HGFkcNA/KI0IFafNOVub0JaivjDyQ6mIjq0g2f/mj5g3/AD2WCuuqRILLGK107cVfGkod5oV7q4P
NaJ5ZkD6IW8Gl7BDuyBeAkjyYNSZb2nhV8eKHpxCASGm/F6Vt94DzjpyFN6t4R6wsVU4aw41T3Az
DtxCG1gJg9m9ophJqOdRg2C+U+yNWwnY580tH3/0gOK0lMN5cEUHmkOfcN249NmNp6rmRbZ/EXfp
xC2l8wzGiDfx/Bil+ejOerkIKLLMbHAkUm8r+shf3crjOhi6I2834Z4FhZwhA6stc6/WzUiJhZSQ
RrYjhMv1TABN6P4GQdQe5r6rRMcveSyzFQ5Yv9sd4p7avTGNPm8FjmI4rQI8ryDfBFVHtpzxIhms
XtxKniY6VoVNWaRoZiknSKRI2nn1u+TKt/aeR8tXIhh8eobZPySyiox6hhzzbP9ll00IKp+NGsa1
RrFk8d6DWrJSuPc6F4AS73rpMri0JdQQvwuTUsmFj5C5KFZigJqmLHSU0rdxm3B3LpO808zNBKD2
MEHosOUZ8saXoFbpft4xkVoS3V/2nqHvT7Esj1wUO3PdJ2bu7Qh94MKnMjIxr+szItpHSqn7UgMs
teICLEMnpIV0WHTCJwVmvT5pXd9d6PW52B1STQSu5YbL0fNSc6x/McZam8R7/4yT+918ziViogJF
cwoQ2DnS92CtJ1ExhKkdXcaTBxc5XYHJcx7qZjnIeSzF0pCyTt8eOyZh+z4KqKDlsH1hgTKyRQJg
dAvtG0UoH6Nqyx36Y94zI2cL3ZRwss6iRsBl0KEKgU9DhXwb/YJORVCKqm+rNs8ry9V9dXP8Qj1l
YiU1M+tMsKh4bHFZk3OAKbqu1QrW7nEBWayTkZYdtL+kfuufIKkT+a3yzY6+etqGnWkTs8n5VfAR
N/KMNZCJkfs0oZ8UDxM+zPXyKfX8l/BwcRaLUq6eoLQcqKzGn6SZPMLbj22jarrXKAXct2UfZttk
zdwURNfvHLLUA176gcB5PS+ZPINVsGU7+4OqW85QM2PWHaSMCqkebhkIy6v76B41Tb3TKTgHjEmz
tCRwTQgoiJIueJ3jeiYJDpFGX/G4S5w+v5Kthkk1zY0Pd38recFLsJPOhzAl6PCOEPSwTcpCfgg5
0lFa12rAbnYkJ2FHRK07w9A4lsyBVqRGJuMZwJQxtuURJyi9p7cHYiwEApkTZUyplIW2idkb1QjU
JGLvPb7FRvNSzqzBHnADScBqgxUoJi0hW9qcg4QR3eMPo3KFPcbQMydJSrDjW/xeB+RaZmGkjKzA
Yuuk2KamCLiEu/JdQVtGbL/3OnKbvJ11f7FUBEum1eFt1iw9sZDC3k2yjppZ7kupkCTF3z7WkEJE
9ytfmgQH2PMr6Wq7d2cY0s3zU0Q342/SXVu+hr7DPuTjvXZC71ElXcJmcNjpJPy45WiHS6VJvZfO
oJ78kpk4wsW9lC3aLeC+LHlaBnFv68iRkiDeG/MtlfDcUq7Z1sy1TNfm34cRwvssSAHJEB7XJIxI
VM9lJrPoBHRJMIZFKOn0cSkpKC5cQP1jw8Rv5/1Q2uEpmX3zZzxYdUw0lK6WZSQBk+38+4BCvPmU
tSHelhU2x0U2si+j2qKh/Qe65O3i1dCDd+UCpL3/76pYdHvyd0ntwsqW35cHvCPjGdwAWf27kNj9
joadPGu7+iCyuuNmGxb5Zv8cO/4nkFtCVs7jktreaG0cJykdDs6nXktDce8Ff05IS54KrA/w/+/d
zss1M9w1lu1O5todqxtmKbHdTGL5wNqkJbfAGMvpwgRuKiLfli06aDhM+bJqrsCFE/y8Ljave9Ch
LCBc004BAbfuijkImFa2skkKTFND6cMgyznWqZVbTE7i/hyWtpXQXj/XIaWjD7s20LRP6/psdKHc
S/J4olWBD2bY5rbkaIURb9YM5yhA+R3Bwog6xQqTklmklnGGv6KHPVsrJrb8ZJQXPmePeQLM38UL
lwsCdlpp0qLTjKxbIgssQnNg5ia9/fA1f4xPmJ8eoESVWTAtu8U99cpcoV8yv+l/GJ2350JHlceK
xdZIuTCTSmj4aOc8Xo5gxi9fMVDwJ8KiAEiA98bQGUNak+LGjHxPOBvBFX6tpjOOT2XHA60hVuAN
ufKyaHcrUEIijoacWB7bYH4jeeZs8bgiRyRYVHwg0KXDgV0SoS8bIukV9PHtc6gYBFpUxW+DECIF
vWUPBaedWis3ZaP4XVxZp3DVAH+nPI72H2MvriZb8uQgoS3OMqFt6OULDNmW1rtbVkz4tC7GkgeZ
tEdXgpzadqNK1J2T7nQ/HMC2BmxqNJSksMcam9vNOags5TThM6b78lJLIawyqlxq3cdhjwn+klOA
FR4kkdNRZGfN3QYkE76pMXO5IAM0D7h+WLCxTx1bFMc78jlE9HF5XySpDYK1sCjM4UR7ZExPrh+N
DkeYIKkpVL6LgOMT4CR+cOeR+zEmcW7LEoSIG7Mptzz9M7ANDVi8XZbKeAQRHPna+GGmvG3YEUwV
51Oowf8gCprEYMzQi3KgjGJ0e3+4q8UirFfoWG/+pWZc2wtzMpYYQUUqIA+Dc+IBhtt+dBYX3Jp4
TPdywyhAaHrBCM27un7YKup9nxZgkeckMWTiShjVYq71UsZ5oxXeK7XSGn0FRmL2HQvfwRKZv+hV
SOD9NdF1i7aRN/MRNa1CWG9yKR7EKbZciry9NiEo3GeaeP37OEi/yGjxHr2GiMgWFVBsU34Qh3lf
NBdZOvHETahBpjKJ1C5tNCmlFYQyjHT/aQCyn6fdGfj14cbp5WYMK/XO1tfalftVkIwBHtTpjkHT
fxiTpzGR68EpbijjkF0mnotLKz+h+Zrgg98RddZ90zlBYhmz9cRPlCSNh3KHeleRo56/KakHNY6y
kZdfSTvOvsrEcs145u66h+WswAjAscQ3g1aCRucbm1SseA8uBTPXA0hrWjt7VidqLPc8nye1nWXB
BOjRIVZnWqvDKOQqW4Ajt9XPwhOB1RQnvRvg87ItodKunuqr5urTlDR+QEiNEdFwuTxzqGyzjp3l
XV92hxaDSidmXgyiBGjgi8trFNr5eTp0dViBsDx7ZSsJxbzl6CMGigfeXGWVHX1uV77aA0VIo9iS
oEDXEVpF7mxG22vTh3Ie6yNGv9vczzGBmTyiwiYBBfAYoX+m3EcB7o7D45Ff9amPjugGkylNZPrl
V1KJGQro3N35Arw1JLHOoKi1LcUzhTCAuxhQj3vHjI+ctwWl99AmMApcRS8pArWDthlK6KeXgK8T
rWGxHbcR2mrZEp7YyWZ4aPKj5sGA6IN1cIz3gfOJrI30+wJbaT6RoylkOjKOEGpia+q5OymvObmj
B2b954YgR9KCoZeoF6pYHfmjUX/NbFrjMMfcp/bVtUjj3bIJQNb+FBezyW+PpxjBSBw/NMEalkF9
9Edj095MtKtheRLKaDTtsi60O19Wi9foEvzMrZXlqPFa24O3/2jv9LtYlSG2PanjzkiQbkzNN3ee
2V1ImYXdgUq9iKH/eiIn/vPYusZUQsls1rM2HB9fznF8+rw/ZBwPMUujnkiNT1W7rodGBP25K5iA
XGeh6WRxaQYiO0adVQ6s9+Y7thmjXXoNoCUY2bkj826kVnT4rfb5/s48stp7nSYoKLKwlETLwH6X
VZeo7XIAe61HlAgUinrmu5exoN2876ZuKYiuYMskXhHckzi93aiiU+pnhg/yVqYH4pDa2pDtRHIG
WYCvd/cSCUBSyRZ5KqhyLzoM5my98Rio/RKDBzGp6BsZEcOi9JGROv+1jWZ53bC4N9MnUm6i/ajE
ydZJ7PFqTSwfXO1AaHZDNo+KQw44OZ8VhJuVTx09JHlGrRvSc5JGZ20Omju6uOUxKU9xKLzm5hVD
8iilMKwVAqyXmaG061OiAcqtaw0Ogtel080crgO/hIv4mXeY0prjNZIOsE1o8qYBaVl2deTtW+2l
co4BHtzW9uaBDeB1ADA2w9hOGCO078MGgKu1jJKl7yW3JU1d43SC8R/YcaVmomOIvM8IZC0MVMj5
rzrKpzGxoRvvSbxnPm44y/uN9overqT29T8shxuQjIxQdAd9eUnxUvmhII4ZevFN8OXrMAVnarKl
cqrZpxpFI/iD+bbOCjTiYRuuo2pmdXEemhyfsdWmMdASX3/7wWpP9XZT+9uJejVv2iMCWaPKZKr/
TG4c7R439sYH98sTWEmoVC5RXjVxFb0KM1B4pCoThc6qyd7oUPGOfe61J5itY9PtXEpGguWFIdnq
b/070bNr5p4d/cV4sE1yz6qL8lbVQnQ2LuW9T8BKPzqWTKnyiX5R15X5z82mLpdwd8pJXi8mk0Sr
bxwxH5nZ/xa3rGN9p1ma68SzdzpdSiA2ztMV16N7sw/baHJqnuqK63H0kKbxN5Zl4ZzmIZwajuWe
bNIPbevlgoxMvh7U4S3AVGklgRouzJncaFKqNgCxQjhEXGFu8wVluMk6SBglZnVd1d+b1Rf0sAiv
/PZgOjQt2s6dMYObxRRTSh3dA6854UBRokQrQQrM5uoPQM0RXUBGV791qZk6c7RO90qKNnsaBgVI
C3sOPPdFcRfEXKInkTfxuxBgpDDF4DOe3Dm0kc7kw0a3sczxP5MkoLtJ0xnsfH7WccdgzsCKUrmK
oeo//SzOJAzLri5OEn5HyZ/rQP4VUeWoIxSRcoxiJ1c6ud9y0zUoVhW1kIbvyq1fpsoLDSLnbetA
FRv0xG5lnvnJiCb/61mGttBv7xPlMGytLqFeeWq/hQ0C6O1L9jQSbyzKHiQpm9MZxmYMct41KeWk
FGO8n9cKEx4T/4U0etz51Yidmwu3FI4IyALtOOvZB6sJj5YKo8CbSisSXj8pEs+upwL97KfFwhtI
DOwX7kBvXoN6fep3P+IWWjMTG+JiXg5Gaa+xMyc4FIlhCAGRi1Sf2q2qUpH4fCYEVw28fjmTEMdu
8xZWgvC95VWJTub1lDqiAP/H+ruZ8dWnDSFQPpy09t3QshpkF484JkDzocpSJz9Bxj1frNUqSnYc
14xq03uPzLqaX8y0zWxbdeYb7bT2agq0Dg5sTiSndUTrq8G6anspgAXMGv0/WD0Jjov3Y8DqTo7m
tWBS6oM4ttv3+Vc81HFe+OFxItbT2zNH9IS4OW3ZZgIiDocEaOoXrRJoEfp/KLBJYT9o1KhPlitX
hPzT4KtEmK+Be0BBCm0R62WiS2amAagiz4X+kNSWc5bGFgkUd9D7LXl4183b7KxPArr6vX4JYTjT
plPzi98XRyfwVKd2FNKPeLVs4oiuVpo3bO+F0RgkdZEfQBVG5N/bYsCniQvSRAKS8RsLNjVbyrli
DoI+vnLYVGa6gO1xgbLg2eo/10NxlcXQ2swLiXOmqoEephjc7JYE0BUAMiDEhjkO1iuqMbn0srmk
yTEnthfX3uL+pU/NndHOgYVQAem1SQtyUA4oPFfrbwRI1q/OSPzYoNhvk9nSs50EpeMg/37wCOBf
2IRlOPiZ/RwwRasOP5EqGehWwDP1mZMLdsKYGdrUqAn6Zea2DhQow5SlWgzNgKFQ3VZvWWmIfRjj
KFnAfadC06gHjjE4oL6dkVu/kvNzLizyZDDP+wtVZQHlERAtOHYEgsZFd7pvTdrFQvreaIsrl9DY
/vIip3+UrVw5VQUiBFcjkAkYEIwBgPYqD36vioPfXyjtnYL5yy1VQrRS2u9ZrLZxeOG271c8rk5q
y2FxWrwr6OJwG/J04LCMVVik14+AKovLkCeEKYjJR7g4+cOCKM7SVkeBUz+F+0aiRnlxUSP+LNiV
s+CZW7ICaXB2XQaYYH3eUueuaeZKz9g3g3CzPQi8yfAj9tXXumFvxFiOmFhbkwoxBKSbUSWc5rJ0
Vq7JgratMhfASpQ2LJ49UlwU5L+Aobxw1+p/ox497JUy2qz4C+IwWZFwOK8024y2p1fh8lqWSaG4
+2aQztxwHyXDZgSgUPnlKdDdfLrmEYC9UVH+2mY+N0rl56YJkFWpIs5AUJ+/0gMvLwWj2voZAGVL
qCebBhjW3Dxaz8qeBB0CqvKXsUSIachRJryYERUe99t7L3C/P0rsRqQ2+1eMLLLpA0SlMUQre/ce
YXxSewHuRMevc3LKMvBuHA09BZ7dpUBRCqDZQP3xZevZeiRJJo6Kn4NXFNHzyZrAwJBkXuhb7CVV
/Y+sEGuwJ8EQIWOytI1nJdwXFZDm55xy7MZKqnoxBkRTSIrcMwKdPk9dwIrNA5qNyBj8D9RIND5g
KdB0a13Glhb1QNt02tID+8EZYiSSZVMQuxwYOoLeodPRFG9IzNuhCEkRB1f9Di5v+M3h1ldFqNxa
VyLya/QDRv/cziD3Ji77H6u1OQL9UhxzHHbj4aWHpSkhApI7sRF28WPObBtgGNi5n6cA4+bRhEca
alr1gdUYs6uv33aqm+TXJ53SCgB6jYDGiczvZIU7dNTG43etziAbkc645EdntvBxxFXTHjSgZQI0
TOwWTnDs85zUABO5nGJisBIyQt32S6KixaNLhbqRvlqKQeAyGxxSerF0OfymZ34DbYWTkO8BLE+h
96/nqn/SoSwHVKG9smKrSEYlqMLjnjx71Yr9Lq4EigNigK56c4s+GH3BLF3ZeYE2eVKwbnOlMmWO
AciKTHuhKu6f0yTVUxEoMHJZBBAvHQaHm8k0bv0gO/uoIGtnfwPpYD0FmysA3WNYk/ref91ARLdo
3O9P+hToyYtuCfVFsZb6vTZe9Ppn5Pn/SjTcTTJchgAlwXTFejfi7qZY3KYyXWB5XYHk3TLxPXyT
9DGoucgQl5FlEuvtKmTb4wCk1fhCp/f+xMoMty5qGJVGCTGjNczU03H0szSujIV2Kj9ASq7HUNQJ
q9WjQ8t4wY4mQgRa6INBv5i2yv8zAwfRE4lai11MguPaFzwGjuPmFvTiscZwNwCa6kKTHFpR0RjA
2RZggXA9nRELM+Qmfn0njrxg5U76owbf2TNeoCGCnLW7kJxaJeXBo2WDBYEuQa2Jghx9D5r+L82Q
xA1oBlzvDbryLcO5wVSH0eh64BVMo+dKpkD7yZA78Bd1ZBnotOCuSieMPEswNgGEPXTqJu3/rx1z
g9+43vT3mwDLa1Uh8s7gNC86zF9e74jah03V6ONmQ52TgvFf05Rfx1WuI5ipRln5YqNCmCkCwsrZ
vuKqmvMsZHpcjXFn3cePu6OdauzDXpblP1y+Jefw2lP2HhnBPFX5a9xjBNnxeiemFg19g4ocSlCU
X3K4Xh9I2e+J8mivhBq+5DvnL6WhLcKFdI5746PklYGojadt8tNhtds6SjkQSig8ofbCoIIVuRoN
i05eAN84Wq2xnHCuBUhgE2SA+kTkJ1U8u/t2hv56PdDgwVCQ0uUhqPaPxRULNyJoaMK0rDzS2kLe
O9M8QAqWVfxwqdbSGTdzTfoStHfsI6ZW1o9HCuXNxcReif25XY70VxcbBQ6MqkZwNsSeIkeQ2bvr
HPxJl6Tegz7wMXFYq/G0T8ADm0DJEyvfSPGJGngSkFVNPSq6Em0qLmTijQyr0Zx7Zd3/X1XNXtwz
FndvkrLN3/b3bIBZIswpgDK2RZ5dxRCvav/eTUb3unG6e5f8mwOkTj026SuVCx/cIToRVKO055fq
Kn1udiGNx7PSQD4v2oej+Y5t2wRosg3K9+moyNYUWBT5YX9gHNUDzkLtV/C2eri2v26apsqXuSXX
pswRhImXmyBgMUUe5pW3aJALwe0n+2odwWkSpnXr8vtW75KrwJeGa0pN+Y5w9Nes3p1DQcp1aHei
yUcPKvldpYqdymbpcQp5rkbrYSIsaZdnCSYAxw2ZezE/uzy445hm1aYXt8DQfLuR+beiHIk56k5k
T2Y74Jd8Br6Ja9Oo/P+Z2PCmW6j590isnRIEPcAk2IS+EFbnpG4AzDsotwoTD3iOUiT8gDmGaJKW
nZSnoqwqeewiudwat8neKDVjroWbhx8DzUUEDxZJJJqXRx4fnyKNIAcyAsTJ3qpSh5MFHfKioMww
7ax4ddgpEFiNkUTOuTMv+PtCUOeXbsLrQkEmOGbPVORuXoLAkUJceQ239L7XKqGpSTc6NgcySHW8
7dB345BhcKBGwMZ2+gJDxvmIvqhTlA3kUd4qB8FaEMC0zkwXYkO0BobALqeJTapHKliHOCUH5DJm
tmNY47SuRGz/sPO0JgkCX8jpFIf3G7nDKk6s0X8+KdRBwtY2iIQqqhQkaRJ8FLyEYWE24sw+gu0t
ElPiILXKxTBYb4Ft1Qdeqawvn/s0FCpyCdLOZdxL1WWwU5numQ1jHxOXW0elzaSkwKpsuqHip5js
KikjaF8nKrIb4+YQGJrn1S8PFXxf66hA4LfzTM6o/OUlT5pmItHNnLGbRkWAPyHN0nslop8WuLYG
3Z0ki7ZuWgehTqbX2eXKAuXsAAnBopTTcdpg+OPRRWQ/KNmgR9XmKTiLgMIK7Rf+4nPeRpMBOZ+z
dCQx79uz5/ryyKgs1dVISWxcbjezrf2japAX4raSF+syQeQzYvDYhf0zr8kkccDmVs2X1pjkmCz7
y8lGFZ6y09kaDh+orwPJb86i67m26XoPOqUAKubOeIxLCZDmggzCYX7Rx2MY7muFcH/U+sgf65h7
ax2BxOoajap3uMFrVRAt7VLh1oJGxBQM7PBLOfEW+STkUmm0aLdd+R4uNJjzEHpRcRn3xTWtVrjs
XdQPKSfPmqZhjCYfpSDzCxru4GczAAbrzu/5r1znCLLTUHwLusyDMfNxjorYst8/aW4qfPg1GYP0
V/v9qfbtRq9EI1bfCZGqMnHJ+PpcODB3D/UhhQbSCHkPPGeQNaHEiulPufFj8RI5Uf7FBnukdu51
YJQ0x97D3n/hHH03nGyLm2Yx6C9B77INUWJ6qZT9fIAIHPm6RrZQhv6uVzWDMLR/LvWtxcEk/ptm
43zME6PxHnTShwr7LrsdOoNqg2ixfSZk9AbLm6Q+OJk2pX7OGxB81pnWbjYFEIcUQpM55PBvceuj
9GVJLgtCJlbriiy9hPiKJ7cMrGQ4YfETmOFPtTGH3MOjN1s4yNof4EFq89cUue0tCdRRSVaIDtMc
yGPzD7OIkVLRqx40rgg+dmu7haoYCAdBLFpaJELIgI3UWBJ3HhpTNFH56Oecu017vZQ1P0PNqaJp
sp8aI14r01EdsFAdRYBytOPSazFcZi966SstX7bAHQmgKD0KFfD5nyz9kzEceQfO617mCeOXOu0t
6IqS2UXAKYANKswTKmozWDCOdC5Hd9l6PSH/WDKHux+1yXn6PoM8rOn0M4DaJk7qZmOGPY+91Bkv
1I3qbKQZAkEG8ahy4WiP2kfTqjjNd/dHkEv8sAHlFdsyHBYRYYra0SRnoceHVwlAmG9Zhdt+RWOA
+4bZfCwaPEYRBlTU3ckGYkaeIiFNftvlKTAyzSX6u2nUgP7lQuyd/OmQdPo2EW4uHd7tLGFOAXYi
ko7QuckmWGSLdWsMqdnMELA8x6smUcpp+u1t+lxhzST4nrIlbnvcOJUtc3BmK3yGSnGYVYDGZHcd
0eEi5Xh4gOD7IzIK4hOSLOoxUZuy/yQ9isueP9hY3V+PMRtQZORKTki+9dvJuZyZAeD+/V310ZW1
M0iP3E078zKBxC4KxdCHyOsGJ+cYVd7XhBUNht/l/MveS+Y9FRc9rnfg8X6ob5NlADg4ffPlYn+R
W7Gm0cjr+ilGogBjFMpw/HOT1R1SPqwnD9FrrzZrUekbaHB7y+01DvRnESDBPAsoUKj6yI5CY2n6
ey8zgLjZoQtN4V2mp/ZDWBQ/FswcfjkPikj04xQL8t1HXLABfvIwzsumSyJEiyHe0kaL1V3G51Ru
NKR+zoXT/E/XY4RSouANMXPQ++dG0MkUlqFRLSDh+ewZN2AoPJVZkDARgfPfegSHD8odFPvIxMIu
cTaOCRyfQGe9w6LHmUTlzvilJJTagtfzpnbAei2d3teCo7UGey2FU5k3hSC9qlFV6t0zdDJyFZMO
8o1J9P4mA1+Ews05o7/K4b1ZigrITgTtKXiPHavYZvgtp2rIHnPcc0qtO0KGKpG7aHg9C16UYLQg
nBzV70rMpUZLz3vW+77mkHMeyqR8G00fgvwjU6c99vAyBSo8dJeG/XWRQl1zHxygACNZLHCgBetl
OXnQ9cYCskDnxtxi8qIsgRL2W0tp78Q3CLbELqM/cjnGYpp0645zmnAzyZgAS5I0+TVbKFxG7M2n
tTspuzpyR2iMWk4+hTAPVEfci8Hzw2NEkqgnTlR+E3fzfxp+v8VAOHVkWddJ0OSryMVoWeQdlV1s
Rbe2Jwz819mnUs/xaAuYXrjQeD1Q+N8g8HP5aaLdUFL8v1ckvwoJ/w0nB9AwjtDqAVXmRpgrUFdW
nlMrpynM89a31Ho2brI1emX4RGI/urKaxNwFUNExq6S26P/BvdL1rlBca2CHPh+PrbVbU7fSOEcb
jidwO3JSmxwzMnVaJ9LPI5DMrq7PHO50NqLtjxPAvgI1jiVwtHOaZbBho5r/klKzV5yKFTxxPftI
dT+QctfY9y8FZ6cqmbx4LTEsshXG6eelLKXxPMav16uLzYWGSE+G7AhDNHVe/rrfxhp8eQ6N4XuZ
6utUZjyVXQzSmq4TYx2xOEHL9y+Qz4L+Wy8u+L+Yk533HOTzifheiWSGqF3cxAUbyIUGzYiKLic6
u7MYjE39lut2flZ6Hfo+YrA02putWscas/EGMZsXLJMXLRuxSxgYSVvJ8ZkG9SmzNIfAmuoYv+uS
9QX0fNsB/t8G4zjSWWkYQBgUy6aBpIHlgcTMZ1K/eTsSfun4ZvhF01CIRRNyJdU8YtAW7zUUwPok
skT8Aa77spqXMFSEW0tzQ8P8pCwYL5MX1E7VQxDF/ITfO6GI6vwAEtVg5CmDg+LgvcnHd8Y+FZUn
nAOijExF5zv4AzfZc3JeUEEicE9ZYsXyd5fVqAwHOHhzZw2008Y2w+YZbIy80WTPmica15t3DsvX
Ot4FFAtzqbSF8tSt5mUsg+RVgg1BzU8sieNJ740dWg/+i0a4p39exSosA90H7AHf3KWo5E5WDBg6
BD+/h1mf6kuOLa+6XMEnu2+Apa49JCiGhU90tKYilJEmJTNnwOLr15nVNYprQlQ4jm7/2UkCw11K
lX7NO1NleS+swxleNcFjksg2Z9BF5hMHF97w/cO2YdnMRI4NqXWYBoWTVRxJew+4wXleWc7bRFI6
jaAZ5bIYV4hEWtWPutVbSQCO2h45/pDQ+sPi+97+8z7gy0/hjHhk4SRQi0NNhyqozf04djx5nzUI
Pz2FwaqhQPZ2TU/YFU7y1hYkxfYG2Tm5UM7pZbIS3yiCRr8dT3IyXIi7l/m9wIhHPfgEwa60SJtq
Hyy9cA3Xx9D3tnep9rQblmnb+JOJ3zYqTpLZyDPuYJ88vgayMGj2VUE0f/tCa3ROlpqrAlH5ReEC
67Qey9DiCp4z6l/4Wj2wXj9gKjnJd6QAGlhGBfncHPKa1opfUXGeMN0ZusVntaAwBWf/j8zdd9Td
ZeBMJrw4NHFrrqcvi2pmAuvJUP5RXw/fmag7ZC3cpBRDfeGgAjr/TPOvsW14qxQ/jTxasso673Au
IqtqZqFP9sAQ3uku/cbkxHbyiMzMXpaBy8p9CExZWr9PN6YJMXk3bAlLNoOSliwpBICmIjnyIiRU
YYG4Byj8lh+Le/b4M2KMl7TB6on4jqUrHBcaBQXIKCFn6Ov2sqp8GKdDozVTY9b0sM2TEugoSKXD
n/Hrr1oJPDpaIZ47fJyC8iYda2C7B68/7/4fZNFcyP8G2nyXS8v/asI3vhoujaZApAdaHRv/8+0m
YoKyS+PZVnQMJHIFRMgL3Pqe5t76i7LukG6P8Ls/QwaQ8/G9qBWDPJrzoi3YXJ2wsQwKAuUqlRTC
WihuZesmVyCJOU/oLuif+Nwm+zrWAC5VCaLwqlHsODI59TPb45PoWsb2EESlnfBBQpTvxjso/zWm
t1s31RwkglbjNVBzmzyXtfnvc8F8oeQF2deff5fmgLFrqLUC/m1MmBDR/jRVGNGuOdmFYy7YTov8
xgywanPKh6an8u41TZvE/BdA9wKyqM7e7bwpYYfaLvD0pjqtmzRUx3BY9bFwwfcZUpGQKg1lZ2oX
P+Ky73FN2x8cpCHuNsmRyk1slOnECgNGojpzX/FZedRvq0MqevESkzLllDqqeKKBgvGkb/j/PRFY
I+2bCcorcd+B1H02JjNlES7cxwyz3IDMvB0WyK32Dpw1GBl/Q/e5372+nlFd9fs+YDScPvWcXQXu
Dibkd0ZRctdfm+z/NtKvfPbINeQhXI78MBfPY/p02HZZS/7X2TAh4oGqB8N+l8IX8R0ZBZU33M8E
jfJTOZvhp+PuTgv1+Ux5a/9Jc7K9iq5gyZi/QME3CfFdXKz+SBp8yGjzZijys+SNEURXYLmGgSRF
IBp2kNBltTkggExla3SMSqVTwjt2fQ3CJIsQp3pF2+zZaz6ihA3uMVuBlDYmWnbY0sFbclBkbsmR
CwKs7eM1HTblbPDYRCbDwTnxnYQ0LQnPVZ7C+mFuod7cVF9HOC1s9aJaDpRI8nW1rKoO8G1dqAkC
gizI9d87OExejcLSXRqFVYVmfqeaHVD0C1rULMiAYT7KTzITrss8RwNC4kREb4EDdJcMRsERiNs/
IWmiOOr3ZfaYjgR15UJFwvZmZOrIn45mCWCPpTpwbTJ8B6/nxCo3luvYnvkZbbnvTTTnFY+xzl2L
EWLvS2lAFyNraHhWBoNaPzy6TNew8CU4vB/MafORpXgIde/6uq6ivDpArz+h+FdFp5Wt4Fir4EVf
C/10xW/VuXcHOqsSYsBlgUSaYIxmD2EKmw/MOTvPiHj4fHGRq77tQrlzFzWD4V+i5fA0srlwgekp
wLrKJHkMlmWxfyeN0yD8B4v8hUV7DSJpES05dlBzMCOGhg2WAfDbrx0hFe8MlEBfzuETe5HC+C8M
bP4Ui3tPzypOWjIivnQP65p6D7tL1DlVVb6qjMqyk5rdH8xXRkY3+gHbXHPZLD7CI08AVEqD/Det
MqRVMFZGc/sAU2W0FjEXIoYHk/D5yZ5hx3M6K/qH1dj3nkUvJQuVABmtXSK9hYvBguUmwhd2cbLq
IWc78K8YD7j6iu9OWUQHIbN4BvjhovJURqnh6o4V705VKBzhjea9DqT9gYYnJcMdBNFgv8CMH54w
IiLIiX9MFKnTo6BD99bFhgv8F52wUVdGCK4hrcK6S5RxHSNzjnbgTs/bFhmZ67B2iWuWJcwTnwAJ
AbED0j4DFKeiM3uHSH+5maBal8Qjasa8JAqjIGV7G/bmif5OkFCz1OYjRrufABTI/+naXyHbuqbE
a7yT9WZV7bPCDlT1v0JFL47h2ONLFNJS434MzSZ1/mZd4kGtzBZAHrfk1yfvGoOUZLUJyWWllp2a
O6HYa80OmOQTb3mTWQF4fSWhhELAGEqgVeHnOvpWA6XON+Pq2+iWblzBEwbt720WgWdSNxoLz7eM
CWHU90Ywf6EcAW5A8XLz/l2M1+9X8t8lWtTqJAA1XLDADLrQ1jSOmx8Q1s7UW0s6gKMiWmjYt2ZM
GE4fjAn4C04Myvdj6xHD5u9BBx4lxahEiYXO1oPWqRlyvSsV3dRnDAE9/MBF1Aaaa3OGClYYqaZp
kO6k3w+dKAPGL25E77kBxiQ9nRIe5eBORxS6pW0o3WxfN3GY0yPN3lBwU4JmfDoxC67BTegeI+7o
MGAArck0BI+FYQpJ9z6zAOCzegPsEKMA/928dSG83GugRbUlwiS6viRiV/DW+3q3/urbjRdEqY6u
Zkvh7qyjRuKS7JZePetT3SOMMsQPMImDnJEZqO+GnSmWPmN+EuyWM7Rp7+kKrmKX9fcsOJbs9e9E
VlGLz/fXwidpMO+cRZi3UBnldkhincfTSMMATOmj4/t97c8rTk88dtCuGDDCt/99i57BfkAvxbaL
Zp/PciE1bVkbTHjc53WMQVMx+cKp0HrXn5lbrdQf1ULj9KwzsHl0EYAQ0U1elMcFO6twlh+6MRy7
KVB/jpEJoJs4z50CqRSrPBk7//OgQtoYMA2z9X7sQPmyrhSYcT9Qx5v8hahZF8cwCda8fQ9DR0/w
W/rWAHU7UOm/GOSgeTrLzcZjipfVJdT5xuA8WcALRo3VrjIVEKRz/25jozFqvP1z8J43pt8POhkf
vetF6ILmn6iwlLJ3laoczThVuGG5JSIzQS313bRfvbRhEl2Nv6/v+24VSsb7kZXhHJ0VXmhs2ywm
fVpdJJul9r/Op7xlSAWeDK1Xcaqfi5CzBZ6zh6TkPHXTOrdwnk6++I4D27XkldheDKYWRzZD/vsp
IKL2ERGBuIHHzV7VCEdQeZ7GtPY7FBVNtpRfQ9WE8gTRs9uZ3GLYTgvXzR1vKdUdbvHjwc6BCtyY
ooM4ySRnphV/9OD+7fmuzT4fgOj9sXixj2dvu/OgIfURWXx/XCWEhRe16uDDDdV6voUNkTEm32eE
JytyjXu5uJLaFGGGqFP2BXKnKTZC2sgHf9gxwhkC6jYg9wLno8Sh5Pyf6E0h3ha/K59UZcEDyGhC
nCeUvVk0JUeYeoPBSk1QMQrGGMKiwf7XkZfKLhqPAvlCasZM7tvd5JAzUbp0J0SsBfQofdQmDVKQ
58p/85tAeUhlpPoTNcOAkorsbZSmzsOPox+Q96cz/Jsyd9W0+ad6WtEgH3OjbOftx/5LQ7X085Fn
uTkVvBZsDPat/TFbsZgtXCD2AdOz1tJMQuZ8360hoI+DG1roYA0bRxM6IvGRvMROqZmqrl390e5l
Je/iBzz5lzzsyIeGkp6zwcQkx8Mj2UEXXf6QrbO7TtIKE2wTDnkWHannqdhEYYA5DbFPPpHfp/Sj
QrpSVUnzHh6fFbMWH/UegxYqkqWtnkRSkg1Vr1l1BKXPygw6iFaqvlf2ydo1yLVHPsCy9YVjkmSJ
0XWIryz5wnJ1UEU+CcjmIMHfJZ2JmRioFAykZUmtPbqCh1PDgih7TRzvtEZNVXQm3lTV7wGC7lcg
nWTVg/3PXMseNyJsy7ChrREBVKHpmucS+fskOOKcmt1I9NkaosNZOHl9j3YyEWy6BfBDgQL5NPDB
Y1g5s8WfVzflkOuL1eoSzxdKdg8ETi24w5DYmyBYP/HzBT8YHFjPt0Zq7ndyIFl7LQ2fnaM64bUH
r18N4iD8pQHuf2+HA9o/PE5PYm8ZnOSjSG979qwgHvHF8YMH1T1vjICtFlSMGFY+Q7uYso1GyyIz
FVCadQxzLGDZY/NdwVFDN8hfN0pDXzYxhd61dDcUZRCwlVPZHJW78dyerZn3rfiVSjsYqWY0ity3
v1DsmvT8ipPnKroFEOeiw2WdkWE0/lVX6uh2v1H8Gq+SFi/MqbcH4AO2Sbxii/malfDH0y6T+wXN
W9f673UgXFMz9CuJfKp6rMArE9sBAc8sriJssWJE92m82vpWp3Er7+1flu0GQaM/vsHBjjHg5GGe
UPTKy3WyUeCH4HiAs3sFlxV8kZal6sNGL7hmrCTd/gTQG3B2ohJEnF+FOIq1Upu1mycd21fWcIWi
UC7duwO5FCnOeDpj/QObTYb9+C3Gn0nPo0b4WOGIMllrYYEVgGPqJwtse6ZSMcHLvhmaH/bGg2lm
Ge31rIOWq+z6dq5FHMsEFBFnBQd3SvuGJsFTvZzz7tGsGcPj3Ch3+/6HBr4pG3LyfHhX4iY2wj0r
pSazf+mwoKiLLvs/ChE5bC9+qODM81c5pl7QW5y4RSBqO4jtLArepniRqKzVsk8BuVUqi+GJDwVp
WiV2jp24IN3kOi5ne5NHB6a6h+Nc+A93Nq8Ev4hqIFYNV1g0EFuCwJovGbv+wjHDumznj4LghVoo
HlwCKJtNqQv3ss3oMot6EmwMHV/4OqqWULr98COJxmBgMb0k8Fq3s8QDtFEaULFZJs3EWMTr1yDy
zN1dDKsSSVcPd4PySBPwckt3eg/h9B2QQyQEKsmpXI3IOscsZc9jTplyP7Hz50IJNK/E5SlYNyMP
Z//xgHWERx1bFGsQuLAeY8JFiGBpyuvLIVtwlVpumcrtMKN17NZVYXOTTTAa4Ly1rO8REE57ajCe
Am709/DYbtzbf2PdEPelw7SoqWJ7v7A/gHNnPm+uDVXISW22C2+bmEGeSr29JgYTF6ibJ5+KDxVJ
jvmcyQGkg6GS/k8oA2PBWa+8kUb6A1u9yhcIhlysgtki1yFcxyyQoKyaeihUXyH29jsG5FTljE0R
T1fZ/qndA6nxKpHEPtN2Z2PUb9IzU8g7O/PLER50QZ0IBX1orzGVEc6q7i9SR3WY2z4mKMeK4dxL
/oEGrsPubdcIchMEU0u42QnDr4HBVVinRazSBkg/Wgia+7l/xItfTbUbw6An1dDdiW0xl5BW1rVF
RKsXYbJYGXeoaGSkMhjRnqPUQVv6yWifv2h9EjfX/JnqJsz62wG6GZdzYB74/U6pCH1uWrribMqY
ZisqP2IwLWrCbqV7ZCOxdPnILtgdF6RidnJR2mOk9GzZJ4uP7sP5geLujkn5cgRisdXCw7lu2DrV
ySDQ8nLk7L5T9kNue8kacM9O+QsS76SLoH49EXnxnAMESTEaeSt7JSvm/q0cIZU/DRgmsVK0Af4R
q0Wbp79mqujyOLt5U7UCdjmUwvVpitA4uMaYiLfQzIA9fGKik6MKKsC+HdXDcrnRkwTNvqLkFq0O
YZx3icSDB1t/j7DWw9Kbe6fQc5AC202JD6zffY9VpcvDr++GnG+Lg2+Y4+eHb8ECOL09KMYmxG/M
jtVTs60M8CM1s5NAsP9Qa90kZAE9/9nXV1Nok3jd9T21SMgq2SxH+rEV31KP66V4nJXEVVKJSjhR
Z11AV9G4QBBZWDXs0en/vLGxOHNEPzxXhoEpdxrsSTcsdP9hGYbsXQqvpsdvESg7PXmpauVoXqfb
2w+WC1Bf7q1zWuBpWD/E0MlaKpr1o/5ZDHDM9y6XiVEO8UjVgV5i/uA68vFIMu+vUgFLXViqztBF
bF7axWIdg17D8gVZY0m0a+qZ9UciVS8wjysEgd6RATSg+7mtQFHxYH7vBOJNQt5HOPFbBb8McPDc
+uhITC5UUhIt3XiijRGS+XWhL88yGdzjdcsgffenjd89Ws0Gf6RKQwM69Ygteu1Gws3tOxeTcu1w
T44tjJxBO7gBN/OXyQNodHmf1mhQp4K5GyDsNyZC08SZ9ZKmwnCQ+mgqqTCfyNxkRFke7KHDH6LD
Onggy47rZbIeG0cSCtlEw3RC5RrNetAWuOL7BC0s+j5HitzYEP3B8IcFJq4zNmXXAfSRQUZaeuYI
xirjBwZLEJ+HgCRKQE+kzs6aDDgvn4fBRNKiXe6UwEk6BhUoEVsp4PYJUVAE3V3jbnNkRxZIgK7b
xwTueKQicGZ2M18bU3Ji3/ndx7oyB2tyTGuQ6wMcRQ9iqwvx7ak6TkMXnaTszEDUYptV/4zRTyID
gx4IoppDq0dFe1xOLe2cDMonSxevDizeBD3e4pCSfEkCuX+QpCtEbaelpnwuxI4cQyc88z+/XNNQ
s1PGsM7WLdrZAnDo8qC+mMyZg5aRMv685ZqmeGOXKM+pMjqTDAcYQrUwKVxhabsPIKWajCxki6Mp
mSGwb/xxGdmaDRSgmpRgM+WK5wTV6VMdHHRWuSWhAj15oMuKVnF3yR8S7vGGIFyZFC+gzxX79JgM
JOqdMAcaWLk5MaZ1v9Sqt0lXPagkA8KBCSvixzg6gd6b0cjP5nk7xypKs+b6xAceFZ/l0P6F8eUu
TFbqHAcohhOihE4S3qqGgmp5qyguA33t+6S6U5kPYs1G14ZW9uCOUlskPPhs3xKqfEHjwjrFJ98j
9MsIsybe5bJPCslVoaP44qvKSk43Py+Z+q/k9I4ecv1YSKcLE8kFAWA7buvHQw0r5FB3M+Ph9c/E
fSBXa0hN97YSON+LQINxmyTAix/pEnTxcIpZPFgO3LVOOE0AW55futGQAXEjEinX73+ARdPFngyv
MtwdKPD5hbUkBwtDZts2L8ZXBolYknEvpRvph4pzSjs+4XRTWZgKQ3mz+30bjWBTw/XLO2DcuERv
nJrP+FknKI7H4dzhweLTILrTbgU4H50JJGT3cs1nvIQnj4u+yeppwxkNrv5+Ka/Ueg093gAKydW5
AyWgTw033xs23aE9uXJO+w76mue/wchfLl6tfzXKl7+v+AvnuXmCNjO054bBqZ74jluZUcMkRz7P
ity7E2UYpccHHPtbW2z8glA9aafPoWIJFmKE2kpM3MLfEqYisBN6nV8yK8njMLfaG12TTNm23gze
FBBnGF9T3Rr8QqmbpH7giU9kXO0dpG8W9yjgWaQnK6xG5Jq3lAVfgoEJtnUJTBV84gtO6sv2epm6
iM3ozD7NjW3GM2A9L4o7Wne74NjLrQ0sW2ykTTKoSaOzhZrqMxjydjZBed6a21XbaPivxIzElZBS
jy4jVvnvqB/VpYcobdygF2Gr2la4L9rlGyQXCVEJ9dEUoY0SGsGLCco7j0DVzBqaBQFBZYEE6ClE
GPctRmH4QYMcgL/MAzMsF31n4n0iClJUL/ltou84CaAc2tMjAUQ6XhOY/+KeTM3nVEQ9+mIHNlxC
96jCUZJnou8o8t6OYU0qniVvkwqeOCKLBVn6suAkd7UOQUVrJb5lhynzsUfDzvZpNb8wqwvtJJoU
e92jACB0IXUyU9X1J2Gvoh1FPgjnR9Bp88pzl8Eas0IUMNT5p+OaNv/VQyGivPRgRzcl8nYkN9wB
0/C/Ro+PHg0NmhJ3G+eoU1TpIdZ+M16P71/TrYq0k+GJWnGt7jlH8Wj1KnijimRcQ2uaFhvxaO3+
dIQcyoeET0VGYyT8Xw0PPUg87wOpJav9JKHCI0F/3F6DLhMpEIymN7bpq66ZpaoZTM2w5ChHHLx8
meK1ABNQ5rT3IxMiN7qWw9PwNriStqDsBOHl64F7aFNercF14T7kXmgbSnRDOxxoMZR6FoCNygG7
FWqCvCwwdVCVGk+Srj6OdoDSEEZvPQ+mHeuGIpKYAzfqHuqr5SWEZ0HkHNh/WDAdKmDNVEz6pJ+3
BDkrTnajU6UQnMmGvXNutPqWqCEScbIgG+G3xgropnmlbPB7cWFOonoS2U66DhjWQcSKhIlfbstQ
m+eRBuTpZDjDskL8P2JpJ7ryW07Q5OmHDU6dIS+7fi91O31e1H3BO5yUkLa0wTgD7m7Lglq/7LR7
BkkCbtdRe83GNuam+mZqAjh7lIlVOwxbtM/eE4Hu6kV742nLLpAsY61++QBjGYn7VKvAlGRBhCFy
6kZk8xwKhMOkB7PCeQzC03zfIx0dcZt5JHmSiSMMnkJ3bWYIZsujAqWwnfIFc/2NIS/WWgOTKuQJ
vPBYGHCyzpSEzW7F+gg8YWDag2hx1iKCew1yzYWDzr3mYUV1CzL4IBbE2Bumtn3xzZ7dcJfgt5cW
q0s4pupDIFT7MyaIR4WN03fpPCQ8t+FWmzplFGQxo7V7qAm8slpMCaQpDUekizqHVv/8P736CGPo
SCfJCBKLOgCtpOCw5hv46pgorAbwK5Mr7fOIRA2FNUH+wJ6qhs7tWg0uTpR9CfNuX1BpOjXsQ5rj
JQFAU8QNfwmenqd2H9Z3E6kVPfaOCDl6C3GJqasS+jGqcGEZRDLTeiTowaZvigWO4h4sNojmQFgE
pQgwqEgmPLRSek10PA8W0wZWGTNkIoQFwk/6a52GOHGya7uSTNUz1htEfU6hyB37dWmTpCYHVCep
40yXDDx+6mVkNHd8u1wUuPfTJmo0oj/DVyByhxgDTsMZxRJ6RXXoed3wInmprtdzxwZPyMFPYL/o
LKSSZ1RB55ysDa6cxE5c879aAHiEh8QGnKdaFo5RJCCiB68YB/4gt9vue9lNNZnbkG3y3yj4uNqk
baByQ4ZnfzTWn5aAJs5iYb2gv3JnIcl+r8zZNUE9n9YgJuSLAwY/iFlH5ZtgcVJlu1hfta3Mxmmd
ou7qMr3QkQq0WIBcrsqo3q8Qtuv9vtBXkUN773R6sLEinAd24rCWa8KKYygQr+QMlsaCXSxwpwEr
8oHCqWxIfhhaChkNOEuPTh451b0TmVzMjM8r2Ic0iOmWGqhxF4mnLsln+wemCfQPZ/V/3YlbTdUW
D6Va+od0xNzmBrLrRSxwH5Io4qr5ZOiMZi6ueLJUMhEClIeqHFv7vBYKJAWmD/nVbEBJyRe4vUxi
jVASSMHVAO6R2e1/zKSY0g74qZCrBr+85nd9Y8Emua313GNEvMUwzkbeIRQFfJ5jV3jjxV8zo/FY
7EHGPPwyofZglNbCbBWrhq9GKdsUKhrmYeJXu6TiZv9pvbefAzrYDlcfOYmjTzQNwSyyoB48SV0t
/3FhA6w1z3OGooJL2yELNnS8PF3aZLE4A9LYhb+yuoVB3EWvZwIAIxv2TUdX2MRWCBvvysun6Z3F
fQsDRpel/SAmDd9hJFDEOZVIgnghNk8HeiV4Z70DL7lzbt4Bpi+pvj5YGElFl4LVhcEWms6WT1J5
nqXnMsfp7aQDFYQtKLc2sFaoA0cNqi9857f5LpDPL1FXSe5W0scArcnBH39UJ9kHHAXNzZsEg5WA
Uv4SdF5YNUyvhSmBVoRgeBb41w2XUv8Nmdfqf+SVkKWEgvjeAMqodYMzLZoDXmPyHjGfHVYmyf4A
2Wed83GHT/dnkQuB+u699Z2W++HWSbZdkwa0Uh6cFZ7E20y3K5NUYaoB7mi0RgvElqcvb8QwrkwS
LpoVAwX3OrPfWPDN8WfQy8HSrURUFnXktFRSqH8jD24JWRSdRk+aP6ftAfQHdbx4lsl5t0nwb90C
0/Q4ODmyWX9TJCXYAwlqN9PfR8x9/VycbGYW98Jm0muB33yXJLQ53ovlZS5z1Gnj+xui00FWjBpl
SPzYxSWgCmnZJe2dJ9Ilq1LDMHD4DcRMew4v47oRY4DZqmlTJ3+nRKXrtNi42Ir7dAT4XTw2klad
YIhaFR/TOsM9bH5DIAVuOgN7cV1tSQZhBpd1MvqwLWBegxdB+s0F1qnyCtpIV7lGGAF+UheNh+9Y
CGn/9yTrK9yJv/iNyFNi6AgThGKDU+Dd+juYgsEMk1Rt2o8gQ519mZ/IFCO8cRxeZaZClTgFswO/
2cg/nhz65m7cT4V3g6cOsuAd+KU/LuoNvGAdeKkzMUEXhBnKGw5x+GQ73sKVhZz3r/dIVJYJ5a2M
nmVwmOLI0tOfuhYWq7rTs4omGBxJzCgLUmlnQEikbQJRUCjF1DUxPSizPw9UCUDHNu8y4HOL74lt
2Wh+X7rXf0vhHh8674YieAQdXf5AQF2pxgHdZBzMa8yfVRO9CHY1MzUyIq/dCgAt+ry0zKSiDbaY
Vo1aaONjwypdGsseGaSey3DEPE0C+M0ffVtTgcetgTbf6O+t/AiVDc5u+ZgYxDKllNB0RI4tTnwy
bTnfLF09OdMKHfZSjcYQHASy/tqTFsfrX4CyGMdfxdNT5zM8WxtAmEMVhb+sglG4KuBS2/P92n3V
pkYp9NA3eG75xNR2wRe7g63RsRDCmJiSl0jwZ5ov19yaD1qijA2/fRwoTUl3AnYROpTSCk5m3F7l
xbkPvSD8O7LF231JQKJp7ItxvcJSKDQ+C/SBuEqMCq3w0eefHYBdfntIQusOqk98lnA3SoWj+YAQ
iyWk6TGmQl16vpBFUQcSy1eGLr1qoEdwxlkLTqOXlwFMbnH3JG2kxoP6mPDecJipshEDYCKh9S7O
NsavgcyM0Pqp0DZN1kRYXnVeZMwS4oAPwirUJBDaHp6LaLs6nmZKqOgrT4IZtKYnMRQ2EtDTljFy
20mJdaI+m6+5Hb1bNNjaaMcVQ1eMTxAf20gKVmB22h+g4XXtlSC3tF3dvO9OoqerL0GLEG5cjiFw
f7cMrjGG3ZLPtcS2sluxUVas8pANbBhAwlPQhL12nLYPT/hA5iGJACr94M9H1GRGTBRKYOmVIiom
ChDjply9HTj6azx/VBh2UC0ODUuhxLbHlPjudoTnZtORk+Kp1MA0+SQyjSqa5gYKZxh0fwLNQQ7V
psa0B1dxwYyTHcS56CMk39iJvuoIbCxKSxrC9AchyD9EsVLFJ1aNhheB7kug7KDOX30eNqr46Nth
QdLkDgxdqSIjDKaqE94u4SLX2z1R31fFxMyGwH6HE+44tYm275QiueC3yglxib3hWc8k0UfLz+Y3
gxko6rFlUD3WOTsWCRetdfGH2PKg9OL9GWQ2kQLt979F2DxXzPCLXhsulF3TLnoYC7mXfA08zrQK
hTGY7ZjVBuZXFYOb/XBqOL7227QXvE9IbyOwuFPF3tHORs/T5uzZoC9xuEcFL2xsaaGTGY9QC2C+
BHUYbiMZjdaHP9xMHRtF3YlOyDuqjcfK49YrRf2d5aw3vjFkdvcz7SNJUfZs9LcB35CwIZDb3lCp
Urug3g8PJ9GVrrBNLtZo2tGf/lgewVK6/KjZBJkw2ZkPeBwK34yoz64c1MX5K2cQOQjYjQCHmowe
JYIaE2sWQ+A3YojuE//G5n/nS7mGwvZowAwnhhw8foiCiBzJtCXN27rHIH0+7rYt/ZIx3wxrAwB9
kWOhlWYmz8BufPCPZI9+4oHlVM1+MO7yCdhvHvqTX7tsvu+toKnCBWBP3ofgEfAFNf+S89ygImFu
modHJbGMYA0Z+3KZbyNZPyXS4VsAVSC6BpLLD0uoEyDWZwdLEJORPT2Ng4yISN0eqqbLu3WON43t
riiqfIchXNimsVbpsc3n5Yhd8YRM4e0KrYcgcnTBvpjNXxbhUwm9mGk9gtqg2i/bkHTiG3M5jy4f
Yd1UfjeyTOk+IbQhSpqbyLR4B5NMmj/KUY0f4LCGbgrpaLk63tZ2wJYLKK7NF1JFiwsjcwTBbunb
gCSrgnaIeog9oOply3biW2IlI4YYaYZwTQIj3YadKmPo5420zG0R0HmTmnZxcydDURf0DjoW34Ss
pVou6d2HKWkSeJCx2IGmJFKbTfrFkyvIp+RZSFSV/ZMFkACphOtjtHJRNv5ehH31gHmws3B12jou
h/NVik6DEdoLRxlHznlwmsaGvaT/2C+g11dbrCLnOhxsLGZWSsW7SNNtlwxVb+136J0+b2h9uYyH
wQ9+KadVCjaj0iwr2/RfSjaW2+K79swm7Hiw77RyGWyumMOjy48EfTHYruGzRDB22ne0RjsjBPPI
CoS1J36wUsjz2dZqOq0QW9ZZwYu02rsdsv0Bl9PLSwmKf8x/lw1ya0f4jtVh6AbAdPDnKSkvDx+6
AHn8UFAvnmt6Cgu6VrHBn61BtLcwlNVhLG9FmiEYrecgL5llI5K9yP5iRkgmKtB/PC1moSCtLkIZ
dJyomCH39o1kA9bPGKa3juY+9XfK6h+m5gBEK7PPC8uxk/z2iCdD4aRN42LtYJInQgIAqVKaA7Tl
BdfZJ2Jd0p0aX/uvj4OsTIn77tj1AGHmrKDrbQBGLOKS0brDhiNbLoeBZnu65ALmRCc8w5ROdJlI
0cE50c70j52SWLf3jOsYsQx8SpiGvDnafv0fqjUb9m6VcpXRjd2dal/D+Nty8YbIkNvf7zykh0nE
n/XJmJg2V7Wn4BXdXQFYNP/g1cifBUbC6lc6PPuS5eYJN4bLEc9+b4+Mld+fwP3iAkDmxXD6eTVn
lYDqQQ6K9CVRb6yEEeMwSGVC43X0iiwDZXCa3FfL1+ssfU9XnXDCoB0wzwBNK2hxBugX6luP3YaU
abXgSwDKw0Ntjd6KPSX3NRppyOH2rWbbcE5Vbb9eDHZaG8d4lIXYeKj8qJ1C2GzmxPVlSKJG93PW
6XXoIrpZTDtLCeU45MojDE+nMblCFwtTuerSUBAez/6EzY9RqOk08jJGePacHIaoOlfCQAqqXNJ7
M4QwnafLYQQLQ+0Gx5sXQq3WAIWLVa6HtAe4OhiO1N0x401u0L3QS4JFbGxe6hjoXIR4F60snkuy
qK01owz8pe9rYctYvfdMXsZvAlyVSOo8IENzcqxrsMkOhpBitikZnhvwm3mUaxSowJ1JtQhlYcnC
lo44SnJr3Qe8tv7e6KULeXc2xzOpZrfNY5rkmM9P2XiE+CkddAslX2xaa4D/t5C14ZyHFuoQgNui
wQdP2P40tPqbxA8Ln6Pc60nuaXIiOtHXaiuD1lnCZkfyJ1d5Vwu1qSXirJWdkHdia74j20vyjid9
0V+0Q9qVp+8TuSVpjvSMtp+Vva3Sp4LSCtfrLVr8JHO0/thlaYXW1RIPIoRrmT/CbCbdangqmIss
2GN3ukc1M2QzBF99709AIuMNJUIiUMfED4TFiXxhmrvF4ZcjLHVudfKXUANGeKRKyAeDAEsAVxxZ
S784qC4G+jLEfMJlanqTVURSHEf1KQgotgu6mQfl8J2pQ4QKYbqp1q4pTp+oMYVXSfl7/oPeOOCn
rssNrDHjTMfPVaJ782LawxmGNKSqFJO0ZxXBZ06tYn+3GcDEZ1rjug/90bn3bcTOUBZ8xJUOUx+y
Z3eXKtGbYd+Pjij9nQT+/NiAyRAQKvHYkxLcBz1iWnc643Z8qVfG4aCKyrpn13/8qvGoBN/buRzn
sqmI9wgxgKNtk6jWDc8+fmgsO1ohaIPlk31wFNsy4keCm9zuKEnQCC9kZAOYRQWLTYR/vvfFnazd
AEqXkGvNQCVV6HxqsR3bHQutHuPujMkPqb7FYaa9WvDq35Ju8cmFd7XTm4RGFrCBWdmBj9AfQWg+
9AwyiofmI+Iv0LPQt1VcCzRmjIwWLS2QrTaWKRyTCf695AMOmkxRJkC5cDZEWY3+RF1fnz+BvPCJ
MhdcNqJD7WYxg4gTYTQQ5MYbH7ti5n74KyyqLtlUKYwSxcKJ7SlWfhfOww/RrMHjVPupY1a04b9B
3RAynM5xHiudJPWlvafwSZeQLwRUAv7zmbZpwySnXN0tWrWofqBZyoVswZJ4MFax86+pV10fFUId
L9IOiqVcd1cIe3Fw9hJHaZdi5DLuqtLGwjzcw4K3gnRTeK7F1Mc+9lK1tOiOUezDJJTKWJ88P9Ty
sWETK9mQegDwOQSF/eSGj9cEEPU1jnSctV3bsAPqbywfvVF+S6ZcNoTwYMzqhhS8OYw7f4OVSLPl
TsDgTAxVB6/HNtwI5kf1yJlxxm3u5k6Zw4xWqbX7atjh5kVz84F/bFvrvjxCZJc2FiiDA6OhszW2
6sp2mMvatoRyd1rOX4mTj02a6MeAVSTyre5HyPo326Vq1LUKKplvtcnx5QVTxp7mMuPUh8bo+Bxu
+6B/WmJeTqkTZ6q2eiSdJRxOdWiSiB8RiSAgLI9qWJgy6mbeYsPP0XQlTP8H7/CKiYmOL+ysTYov
RspckH+1wr+G8PRG2Wph4BG2mqjeZyT/jFkiBUrULnOaEHK69CKQKXAso4yyh9BQHyEfs0CdCe4g
LZrpW9BsUdzo/l3z+IKBaLk5gxx/nRibJnCBTF08iXNQV4XH0PnADJZZkdhYP75/mICXezbosjrq
CkJ6w9ZFAINNM1XfJik7VpsrijYCtoSeV7zkGeXk0jcQ2SbY/Zr7B4wP/ucl9wifkZGo38DYk/9Q
mK6ZN/QLVrcnGNgxt5cd3Op1Mp6b77EAvOa5RPCubEFXkgC6sGfzD2sD8HJk+l6SEiDj9afn95Rb
51oz/LyyXMxAO5HjXiWcLl5cFoiwXmLkfqElCXcmD0keCf1a9DiPNkaUrCi2zTTF4ojdyWpXOL8E
r15BQ6CWA4KILdejLWm3U9mn//ELqSz/lUzQ8durs3X3DeTs2FaprAjIbjuPHtefdnvj7CbHf0yP
3gtlhLSI0i+VJ3CJttxzUFQrczuzUtrXD1tJ3MmaRbf5Sn0fSIXQLPSHrK0+7idVzV9nRP3bjHv6
34ZZ28K79S9xg3l9aNl79yyb+o7GBhLwZOSgNlebvbSm/XAob8TDdsZb5k59WWgYZZbAZUfBpGEP
CjVWuha8W1cAiqbn1kFFpJ/f3FoctXz9Psi8fYF73sGnuLXO4WVC4S/9WLU8YxP3DBd4xbx3SWXP
lwFiP+nJTFqVks+Eoubh54+A+ubYIbnznuCUEyPR5LKlQCD+nVSg0WLJlFbMkszUXq1obU3zQqqN
fCNbJx80mAb9EkYh7MXWNW7bdAiRh2pKLb8QXUihhpxSrtnlbCR5oW9Z3Xo58PVe0HOIHcBuAgQY
RyWRVoLia3kQflCMu5Cd0hJu/AW/l/1oOcy5KCvcGglcmPeUOIoqICfkvRSnsW7tiPUXmD6XDN3+
vIp5h9kmJFrHnnmPmWSsE8NtLhBQR4LLXvXFoFMPblHH+2gPrf1h4a7zimtcIzESXMHMSeGKOabb
abO0tTopisdkMImbMpfJLhf7CYPk4GIzOdKuYV995h0XSxXfHUO9H/H3kBGG+m4ZiXPVezcj3JL+
AE8jgEj7RuIVZtkxXSRbt06Gj+h6BZWZ3UMU6cpS5PW3GOyHfRd78izXnYrSVBjTSowAkmKMcIwi
e4VnWzyB0QMA62c5ulclWbwmas1VEdmwhTitJY4f/8RMScIksetJPhadoxpR0UPxWW+S5F7+nsEh
mmhOlAZf3LuMjcx1VuS2puL9vkdGcTHm9MuUn9bQnQtRegzsbovgKrEL5OLnPJ5veExO+VIHTrxd
EstyfzQiPjhMcl9g9C9w2R1hnkk+JrkpBBzWSBJ6IVjNSNU1oXM65cuoAsJIc838jDsAvcZhX+Yd
HJ1ZKl1MqpUfgjk296ILq0pWaHmrsXJPVcsTsn89ZaWQqaFLjUhg6zslKYRYTvxK9xuJdSju/O3y
zrtIE8Rmw48TOePoj8EkCHerOOdR2p/lhQPVdNmLrnl0nVHKQXAAq3+3wJDYBivaBcVaDuLBawKV
IPkyrXGPnfL8Xr8TD+qUb17q4rIPLrAMJKTgR5famDGhXIdcGVDEjZvmIgY2Bc6/maDiXT8/rlJo
DAwPIMWACwuE0eUkrt07BICThTdMRO5wQKaYRT0VIuEfvYqCgKwVCaYgiSKGxNm2kA9zvcsslldn
uOVl2dHEI++FzmrKNZgtziIaLLD31YHeOA6Xo/T/ySnvgaf5Hyf+VjZPmWaI31bZhdbx8SHuZkNI
SHurH7qdB1fTwTJmleCxLcJnW7SW+AhjefZihk31j/7pHob0zd5wZqWeiFVyvuQmOxVZE/cO09t0
vfpzF7fEBdgElt5nro5+MQ7eyNEPkj880Qa9gWaUxdBXZ2ul29SHaiUBdfUrmXamfAv7Y+iE6lVM
C0Rfg19KNRiA98oluTW7p2uTtE2J0Qu0x/PNBMF8CqoOXGMf2yNBRv0v5d8IijMpu67gHSkxoRcI
lT2EUP1OCwlgmu54iPmC/4o/eMiQZgraRFji0fmjOsDqaSZPstvRzDDnp0ky2qcMeEuMEzarM+b4
BO11TWFRXbWhwqRTTTeXbdBn/hgz2SIYEQYQgp2vcITFB0xODgUEaVj9o+/21Kgg10WBJ4EeqIQg
mq1lf1J0eiwU1v7qOlRbeFvVxXOmNfveTxc+rPaJBbf07ZE+MBqmoSgNu5rmL+Cw0TQh1tMwimsW
SJUa5ilb27OIZRDuAJuSI7zok5rcUzrR+jml5Cb1dsynKbEMpCX7shgIaIci6h52NCSzjfhsAQ3y
x1cGNbaLaeG74jwVNJQ3/1U3rqG7kBKam6UA0TALw52L9k0yDDHKfUH7AMFukHlHNvHnUlnrdX2Z
9/Wxs7GcoG1CAi9/jPQB3yStlzDqFXjuKdSqFGEknwzimVaR4TPKjrtGXwRp0yV2i+8XfAFqYesj
wSrr1dH0lfNpAI8J2X7Be7GzHcAZ/Mf2horiTmisWnRfwSUgTEim3Vr4IXYIq7UrdkZvixQruFee
bKPoXj0lBg8uQKZOzcD8Pi01rQiBzlg7HnOuKybkZo38lPevIeBtJXR6cZShg0m0CO4+wXi3JMwa
hdB8EYYcqIsmY3372zpIw7BTOjFX0fY7dn7t51irvcPWaX6NeBMrxpj/TAjKdEJtA5kD03S/QNI0
qUv4LmxmLVCvCftDKlB46MbJz5kuJ7ONCsyV8eeuiL3NYiE+akkh9wN1P4+pLc1kJsi3gjsEcSPN
mB6EhgyUm4pEhliDM951esy0v3mQagt8B+DXOQ0Y9CrncOhEF9ormHfWx99Xeptiaau+yJ6AgSjA
sKuKMCItXEFLqXGSBcrHKtWA7lfAqnXDfSh077X1McVyB/gbN8oBhFKGfyUTzNplQ7Av2sCDWju6
99pQZOx2o0EAJAXWSfUW56XNC3pHydHNZ09WDS3UNPOhCguvFnA5I/GTqEu5ve24fJlh4h0itNpi
7/1utnLzrUKoU/041tHdci1C3b6QkbxtJqbFSyz1i5wm/1XM2/XGLTYHCmPe9e9WWPa3TPgLh7eO
h5XZf7C0Nbph5uw/CvBzefhIUiQ/vBCuJ+ejA/TghAmK+Sri2BDZjdp5VcGwXSBI44ckTXulA0fM
/qYr9FEBmJ5Ww+cCpRNo6i7LVQ2QfuM6Mhqr7v9KZhgEM6ZY6y7DcQenNuUyceMQnk/QQjVWZN64
al6KxJ6Dhlwld3l1dobsnS1UXrimSkavkD0OIqlWD2I3/FfWbOhBKWq9Sk0XFxEAK7Hb6myz3YNa
nFPvezX85AaXMGn9C+hAH/9wSAD5eE1YOgaXMrr+A2JSHj1vv/8nQSLT8Ds9idp/g8dddnITBglD
p29cRkyNu1pw2nkN1kEgBdQMBBccCtRpq5tYJO63viFffSS+nst07KrG9im+uOxMAVCBmaTonxAS
boRrPRKMRCWdAQRFPBwMe/CRHnTn8+D579yIy3RAJwXVE9R6s/59uWuy9xVmvoaPnWI05mWFZINP
Ur45UNxM+3C5wruLgzg6jIvhlF7SyzXkoPfWpDSWKBkyP9Uw+Jbs+LBfPqbynoWt8AxSDm+JAfcM
LnssGcnyh4SEx0KWVqpsQ2Hrhkv3lkJgMgYMXl1rJRGhlt1VEPAB29R6qLFBP9mUUv0GklFVyrG/
aWomYmRrRjKu3cXOBKXSUiQxB8C34UDQEsvR/1GEdBh7khTT9T/3uAWY7CBe/dwMnhTNFwoAZ+78
k/VFgHM4ImiPxfijy9RtrYmm0IRZWRFFd0QylwZFjX2HCDJ7U/ViOe2PXE9EVUTgmd1dkLSWeMGi
qV57Qm078bQn8mJoI/L1FVRTyaP9ZuAMhgfb0/ydb1Ly7UG4LWDJrMw91FAOX0xdOcq8CIUHdOnM
bVC+kpzQ21fwDwAtEucFSwRIId81GloP+2WB0YG95PxNa33VBuhCy91ppySOIglYR0DcOKPDaScE
/YPftCVwyfSvYKxpTWiYSBjssvRX6flun7eavzXT1siGzHeTX8GmMmxzvxtKZmi2IwhqljewC/eO
wQ6sqK7YlY2d+0nYLNz5jwiJnSkOYsIUdfH/6OpJGWspFrgkfLubgldk3jYaU8yQf6IFbOCfMIb1
bq3vtMq6CNV6nQr/irqzFvny0H8CFwh8vZtFRrrGvzI90CAm38LhYmtIB3Na9X4bdIZgrOYZSE4r
FX4QvG3TCX24/0Izj074CWFEo+hCkFuvuO40a39djmFzSB6PQ1ZUcmZflayqNspkPklbxM6Xcpu0
Lqo2Go6a65s8YWL3LSJRtcqq40Nkfm/WMZaTVwxh0cvNp+DHJnoczJHyk6NaIi995yALy0nHevi8
aD+grzb4JtfiAy8XgY5SEqshlB8y7FCiXG2KVDtoLxKC5Kz1pevXmV50pMRxI9SJN9NC0aoQ5jTQ
qGapaQnRw4k67sCUjmYveGoJWpSaT3FMhn4jPN6r/u7BdatNX5fl63ciD+TWrwK+kBOIgmVxjvCI
Hwb+aM4NeJw4ot+fZ3c6iF6XgDT9uX4W6YoI340fnIj/NV5z+99GFg/qbdZp+7yRwE2qhJ0E6NiB
Absfyn+8YAz765S5Max1+HE/QG58n4sHcE2gEDbf9A4TkYpc4jZTQ9CiQmx076Fe4L2dGZkNOQRz
TKDIi6VETM+x+kH4TcNg2jcCcaHyhpW169ywD9wEH9mtN0vmOL/CG8DUu+uH3E119JMAjw4iQCZg
lWUwWxu9N8R32K548LMok3hbJyqATU/ydkRKNQ57GV9cOeH1YJpLuXsvx8tTRTYm+sQLK8LwBu/N
BlfM2+zaYZBQ4sWRhMaaCUfoHoClUWQDSQ5lXUKQg0G7s2qkHrQGRKPp6yEgfeekNSTOn3lfGG+H
vCYaROUaQzdTQLKBmiL2TsR2Td+0VBtEAWixlScBkCuYxRoQJ8JdtL/Sy98l0scmMyhQhHRBmSJV
A+IOuPqnE70b/WJ25we5DRdWjwshuvx5eVVcasolC54oCzw9wCZD5FMAy2DsR6+fgIAymkXPlxnF
tE0pHepKNe5aRvvWtC4QoeLuEgrxOcgm/NxCSvmdOKpAO3/q9mUHJDu5rddlJBuglgqTKwBXQO6A
m/DocfjPT2I64XP0QnGF7SxqAbpRY3bweC3KkLKeWt9eBZA3w79/tpol0dZ/pzex8Xfx8pfYDvNG
RrF/QXHDr0E8VwKp/OVERR27/vI4Rtr9tlF1zgFMnPNnKgP+ZqnPog/UfB6IFo/P/GxWJI6N2Y2i
xWLMuPkGExFT4Tnie1IbDYx4gQ0LznFrG5wHGeic1/Fv03sPsuEbOpWtRT6zxNeu91qmlT0bd9qP
5Qk1TYG38bNhExTy5jS0e2kiz94rvGfYf2kPnHbC9KQt56b6JFwhAGX+88JayZwW2HnGs71b6KOh
/xAqUlPT5JbqZYnlpX0Pg3xKKArd+whiO3e0/7WkUbAY72X3fSEin9DOQmOuYCemyr6dVZX6OL0A
sJePBCymX+F2lvkiqybWRtAYX57LTFHnVL80Ql/dtFkEXzrlHSeVdS6U7bm3G3UInoerTJnYZ6Wa
TKlqzR2lvsUuNz3u6w0D1oHmshLRLyTYcx6/4ugY9+v8EyK+dRUaW+casMMFf86gYHD0XPJQqM46
PY1y0ZjlL9YF6hWGDY87HwJo6o2V78PerwrFwKtUOtMWTXI9UdqwfyJ2MDRDvJZlGUxtu7LotFCq
P1l8i6JbADDNoRvsggEv/4EbG2/cDWWpyMzp7z0Oet2//qN82wuFJohmZgshMUJchMhVFbPab8Q+
U4tM7Qnt6z4QWLZA5fy0mUFEx8bwltNfT9/fR10a0QtIgCf0R6ewRfMCOe+TjKzMLb50fBAIP+E7
H6vVIS4tzA5nkZy3F2o8Pt+OKyZSo4AMX+bh9OwFP+agtbsW8srBQW/nmSTxUXH5I8CWGela5U1u
NCu9q8LCM0RGGH3Ut29VfK50LFVr6Op8yRMBwePvBs2sJAURLSB2h3yFio/VGyUTSyDNCgHDmzWi
p3NDcqN9PYRN1ejzVJfZFQB5LGU5NE/tzciOE/uVwO/Zff6PybU4y54PG2rtogAbilTv9QItNt2L
FlxUrS8kOOdqlmGpcFKO7vceWfWVDIoLCCp9Oglj/57MlzwwZQkg3lDRzNx3Ap7+kEcZjWyibUkr
wxDqVUibSb8Ar+/pI+EkP2af/dMiUQfuUDSk0ICtr5vT2qI/M8uPJxgzgVIHipSv68Z1CKHXw6N9
8sKyGk2gEknUGlKMDWtHYuveS5jZiTi7hKqmNbD3/7Pkta23PFioY2zV7KTkrFL+jSHFMbl4CqwH
/RL7PaABQY+ZlvXikgyOGIveCXt8zdPUhXuJ3ROQ8aG+cLvaQecXcBUDxpzxJFr88I1iaY4HEs2b
W8e1ouqZn1Vvn9W6L5D7qHVOMIbiUBvQIrgeK/3RY81LBrdYVSze4S4FL/8vSiAUi/x9MiBez2js
CyDzaVt6qV+pSRdbT5ezZ1cCssAB9it1Mw9R90TAo393GXMWL+eh00kMnPmSaCYDUB3aJCU3P3HB
UTpYPc6ctCRx3Eim6UPAAquUng75G3m6jRuw5hPZ9tRkRqMSJPPscTaY2/82+uQKEFCboj+5CgS5
USyOYhI9nUQrLfnfZ3UuCoCX5mXVat/GZPLqytWZHHlTC5lhr45Brc9m5KDHdEz/dUFPknws4Hvq
lyTpBb0K5UCxl638fGKDqILAb8gZIi+Skg0HftWO8DNaG+9QTLx9hqE+BoDJyIngdVgeQhcDdbd6
MmtVuHyl/ZR7JLfmi8+0mzC8QObYyFAoLRKE2BiCQOQe+jcNCvehT43H7Y+kl0hiGDyybIF30xGe
jUZAmapTuzBhugPZboX6jixwbUOrVMwNRP6arcDenBCiIT3x5XtGbkK6XFoOe+qsW4emxInGqANB
gJn2Hlt6uiD+4/htSLsUXSawgF0ccFKzho2dkdfM7apHwttvk63YQ/xfRMLoXP4+rp5nObYSL1zU
GdW50MS04HCASIwcuLe55EUiuyio5TEzvBzNWk8CvTjWLtFDAo9ScpWCm8Po2HNPiB2fYBQPmt5U
PdEwmYKVRwZXDq+k4vjVezatYvlnBAeK0XuKX4M3A/mLKiTeI8GgJbgoMH7xtQrtxZMZRKIpew+X
16oSS+vjPIFyAoYTYC2a7t4R0OgNRzabYfAiK+yoLKL8CW+eX96nwZY8YlOi45w3J46I3ISLDux5
SsO0tuU6r2DMuZvLhLvab5k2WNXiGeCep/mg3nKFbl9GEfV/BEG2JV39Cd1fJfKhGJBPVbOVKhqf
0lwWTnywZdvPJi9SzMvsvHFqfHtvf32UZ+43TdOeXU/BLWh3MyIz5gEVeU/UIFJCQMLrvJxWkscF
ZBvMQB9dw3gxDBiV164GcUEriIqL81HJe4Y71uTpmqzBlQsHMbbBO9Xol8pJIIBJ9Wu9AHcnBH0V
mEra+BvoPpS+f6ED0/9neIP676sio5KHpmfltgGwkblzgwGkWLcII/fwLgEVjJjGyaa58CywHjUn
wbFb6g2YjEjBiO4ZdEgGrKqYAT/csHmo34XdJrB6Y3S0CRt9S8IVfvuIN4Z3A48GJn51+61DvAOl
/n+IHhUVuzJZQew6U13i18qiUuEoCfo9+tgeqNCqUsiJAnTpqV/ye/Ui0z6ygsewj/JSWQq2R0w0
mmdS2DMbbHrSF+AClL5yOxoOYspEseAMYAgeXyULxToQLo+O2gjAHbALgsRG+LDs0g0mgc9ei3NJ
pqWTVBVhUfRj/1NIJFxhvN65yRmC4cG7TYQGzRbwGTmYOs2/cdUlyeqW13VtZTCPVGU3RTVQsGVc
Jj0y6x/9iUac5FJ2zdQV0oqa/SrqkbuviBOUu3oX5iuURXcngKtylIaZX8DuYP3TjIKYZL/HQ13t
tw7ZxAMUnDvPtIknCPvufA2+6qK3BXW+l9yFrbFo9vaJjC8yZVFHvu9NOP29UnGmhoNHua48WEj2
Ys/K6YiDjP/GckG5zyu2+8ReiMCwputZXncKxi7RqEY6edUUXAOgwbf7RK2f612Jf4+uM3UeTgag
56BiHju4klNuH2DMh80x8uRLAN4Mm5YN3xM5BD60aFuu8AG55C8ZDdOJEMzho1xYvbe5EPQR4Fw+
guN620fsiYPCP0qo4+Xj4Phn+eOpHU4Lt1TZ4XJwq0XMFl0cp+DIiwKTL00ZN6KmvMBRYkn3/mR3
LQ7EKB61c1qQj3TFx2on2+DSa5CAIRIuJSQqCvrAmxdt3EdS6mWbLgLHM7FLYCMp/Xi6R7Sb2qXz
wnJAhagbQT+XGPr9jgTRVVdhih9/XfSoOZuDWK3nYMLUPAD70TnCN8/v1YEIecyxFfuFun5r/NDT
lQNAwj52k7xN/OoumsGMqFYqJwfO7QyzJ/1ieebdIRLx2vO5/lvMEP1aXPUYefEOj8e4Zp3SI/9/
2rn8VXXv45L3WHKAIUFv8IOjC57rZm9xqKQIXkKVPdw4NRnSvMYYacqdUdloPXShMsV0s9XsFcw+
9EKPITO1v3BqK39DG+9LlBQxgQF4hqzCri3bCAr69UG1BfZgEiLX+f0essHFeCbXq/y5MqlzRAax
ON8MkNZjs9k4HgOTDOwszdYgRm4cwLO40Bpddnr6w45OWVI8p/t1oIloHMATapKvk+1uaFvaDNjq
yeLNJION17zXutvGmgMAtyV3Ewd07ltmsSgoimJJf2qN2dIkL7gLVYqR9kdFAlNlxLZ1ETVyj6Fg
tAaJWmPEvhLSv8RL9kiGD7UuK31tKPOU+EZftPurcUvbOxWyZdG/T5jHuScflOBe4LoxdfhMV5e6
EgOyuRof4jEJ3NNaviuZA9G1Z7beU2kWHHkKL+6QB73510i0fujLJhqVr8ZvYGy8sRrb6PJHt/2i
dqawgu7NBK/2owYsEERbIwerKM3avRKOOhzWWlHzJFRZow6TP1ek9YOJxvBko4+PgrjT/NF9swsm
ZdsrAg0Kn39hn1pCKOrTF5t7ZefQcGli/nO0L7tgHHvR9sBfKbmGPgYH5EvNUrk0BNRa9lEhsVza
/te3XUPuWmmS8ngh9Jrsy6Z0vpQ781ABKGPPp+rUCUCwZM5HwaUP1vA2uki5MGABILSwK4noqifV
0vhTyZCudnbgkSL3K0M4Djzr4zKeyEYz7PGfPVaqbJ1tKNZvqSf8w/1KuMaaLrFU6Ugx4dKIZUPx
Skbx984EXAdDqmrpJBawEUfe6NvIWnghxhG+oBWJs355746sTrbMMDmsw1VAUyKF0ocq5Q0GUGjx
4IKflEhky3dZm/6Ip6SvoWuCeAcw8yYZRLgBzjwSA/Yr8WAJMB3NYmFaZL/zTkF8E1vmdVtzD87X
rd4zwUOhuHmEti4w+/oZlwCp5+/svst65DfONZ9J/ux4fVH0zSBBzlqIs5R8HLh0YZiksh9Pu62k
twyitjyrHEZ9gR1H9MInjDKlJfpaUBxe6OLceAQ2yG7IQN8rIWxqkQOXihsSjwqz4ZYTik0k9vXE
1PcvTyTyw4iZpCJC3kFLDPj3PH+Dq6vZ+IwpbuYDeE1tQqpuJBgaqC72Rvwl+4wFS4m53I7mo9zI
tG+XQFjd5bzegSgQJAe4GupdkfctBknrZWtu2nJZ2ctcQahDco5rxz1sbpFnQnsCCK92uiJOamCv
lrkm9/9ENjA/uPFnF7b/i1eL1wz7nBTWecDWvVX+tHM+QGBS5xq/UWtHOyRwbTwxHBSjQmcDtyyo
L3WJYEFK/RtMKDl8DHk3iwOybYJCom5DABfkSxr6jYj/793jSZaW1nwCyAxorKroJMHIMv/0iNbV
i7xdfYcUwYcgOYzF7zfogWPnK73I/oHeshXofpFEWCy/7B9kzUjWzHhZZEhYMh+tbyHeFQn8+bgd
s4QLb6KyGKPHMvinJ2fQE8t5nr5OphAaUT1Trx74+73bg82Zm6g6NeqmfrPLgB8po2ol94nwZDIX
wQOy9z+ILRahhKwl8+CuCvCFto9D/0CBK5HrEB94nnrkQ+zp1Od7QVNJfSXsedIjecBeDRObEz2J
7/oYYFMjsNpgnSfm4RC5WHpciM0W0hx9dQgFKwORh8soydERoqaBHarcxWWEoDg4u/j2+eNjLkCZ
8lT64UWRnndLh27LbHwloFYWlY+vtE8oFfRaQ4mnGvH3/Lw1kWRix82wmO71OEERdETo4lvZU7kl
g8PfguuyynQX24Btkn/RasldB20/xaCma9j8DRgjVy0x/Q0iJ8DOFmkhqIEbSdqpqENmYQNpb7tf
QoS/wNuGPyLg77bXhLzQW3NFgH0+UVNosQ+3602nYFMs5C58nymqtjI33oB4LUz5mwcMFHz5rybX
fyI337ZIAEDd65kxrQp6cJPs9aFickCPVI7FRvHmYWyq7l1d8bsxEi4PfOoMzmZs/q1NTRF1zUvH
6aEHhmPaosFZq0t3ptEyzaamhvrn/PHAZu+qqKZBZafj9sYm0RUpWW24IOfPfeOSOA4T1s+Gcy6G
udJ3VYdJ4G6Ufdd9ucpEbFefnTe36lS0lyf91wZpBsn+3TNCp+133m8B17lg4LlFkeSi+GTMWOSR
tbKCmnBFRqT4Q7zcFa6ey8jhTNY2pifE4Pb/f9EQOIzQ2171Mq8tI8pbsK6MQQ122EL8O4Mn6n9K
RF5ZMDSmHLjaYBHLBxzUwtjI07ilN8saOvTnUWEdhBenmST6N3FRFb+JCIBu/gvQ9/pNhS+qevKD
CTVVCfdmTLsDBeOldBpdMI5ZyB/CvEi0k60P2wzGDXtc/xRBD4zsJ7PP5bW+eYJ67/uV4uzJl9Df
m/yUA/n62dZjuEn1/0gJyWvaZwswHOjKOGe+ZFnBrux5vB5vhN1ceDrhh2fL051egZ+FFyB8be9z
pyJO+aNzlvcZtbcN8H4SOYR2dSa3pxWiP7v5e61TOPXzsa5t3qXsl4p5oZuhSADn9PGBjFPBJgSt
djNq9pSh1z6qwnMvMhnp3KTfB2DVkhtuaNKuJW0cMfnbhO2hcEv+o29cABYFxXTOzYswxoTNAVBv
ZMq4NnU50AgKkcZ3x5kMvoaNDAPnO7BeojxOCKkB5UEJAZPpBx54d7D1CdJt4vB9nMe6Z5TQoQDx
IRlHl+4PYw+5gmzZ0aeZUpnOVjo3XR5rju4wWdx2y606qzkNdbUGt6NRlCRryAi27M4Z/NQCMaRd
rGQZc3M6p8koBjUr4Px2Oejv5JagSP939Vo0J60+kw5/lrHYNu+c/FJdPK/5lv53im2M4WGODitk
4Y4zBxIABUPna9C56GyN5vGSIIDW8x71JwBbJHx4Ij8WmuEp6ETmdzcfFPGHmIHAataKlqHqzKCW
Ioe4dY0sDVpVoBW5Rd0FPHIWxdZgMDib4kbo5fazc3+CElwkXea1ItYn1Dl9Y+ynT/HHJmDE9/yK
xH2XSNLNMBgpTEBFrAI2O6EJ7oMwppoTOxsOFHg02cgDWS9VJXal+umvdiFoX4AJYqMGTDJzgtpr
NZOuEQE8BgcwHPOZzzAq9CJVA84ng1Tm1m7HeUd9klfDRb1pr1ZCX7w9oSR/snGouFzZuo+yhruB
JNLrhAzrr/g3+tlnWxpbGtHEAVH+SDK4F1pv+isQsrfstePJ9Nj4JaXksjOiUiRpDXUwLUSD5Y5Q
0zr71x4C8TqFujctjm3RxEDpWZqDjosS7ONeB+NSqJvUq3Tc5mNwVghNKdIWbfeDMWBbmEMpHqBo
zJy/1WIJwbXNuDrQ8zOJ63mUlagQ34y9hBLY6L1N+ulpF+GCMd7fzzpDtkpkWLdaa+OZoqjt4dnk
lCiRnod8H4iCRHurEbTCOEmu/+dCSZJv98E9RhcJiiLYHsF8SdmIE39VTl+o8E8kZgz/00DjN+Ag
t1/pjc3hj/PMmxMQ49mMVvhKA5xs+Pn1OnrTq0olIdqRgx1W+q/tkNFCQRpuqeJnxM+PSTFkhXHV
qDNk+oazmRJaoDavwJlF/yUSPP0unsGb79+AgL+TSzV2Tf7pEUVINA+Q+YUit4st0Lmgm/yfW0qH
OaXndrI+VkBamdG6Qg6zjInulAW/h+ZrCjfZqqxKRQeJGULvaTJZ8p16sq8T/MMBEBLSc+13Fl34
lUZ/eQghfHylZwKvKn21jOJ91ZDP5gdAciHUm5Q1Ki/opHyC7HXbsbYw70pRcgZdVCxgGoAE3A2w
9/+xGRvlH3gjmYzqx+ESiX76SmK5xDNWsJu+XYgtuMLo8JyV895vk7Yh+FzbpbARtEDAXuTCwP9d
QODkeo4xGExNTjj5vxpuWbVgafFYOnqi5uuRnOVdb/4bsKTZv1m2HsGY75kmdY9BwJtNjRObMc/B
MXUEbLO5gGJlOPiXVhn0wWu4QwBnbEeDQ7tE8PM5OXsdxOEw65oryTq6BpIpLLLBskGphQY6tTe+
B7/bJ7avj9SYPJ34w8HTXW02dsGkXenkHB9dASNP+12G7QEaKvIxT3gA5NJokrgbPVvuDembPa/J
W/FGdbZQfQeXj7Kzckp37AEF0bzTVyV2ggYKXCb6jZJ1SysxxEsz8WoVYzSPd0llANXM/OxY4Efc
RMjBSzosMka+IZ3l12VXVGWgRz7L5pSKheHDeXv37ialrz4aKTTx920vtO2C9wSQFkxCKanfiFAh
TNqfg9aiRgzlqhhzshBAktxT001kjrcb5e2y2nJVH1XCP6WVaLOxQn8SiUUTSQu2/g6z5fg6r/pO
7Klnjvi7fF0MT4x8b9e+GZFsUTwCNdAjDoB8FdXkwKNGRGbIe0EJzsmlOWhvPODpJYHCGnqH86NM
2IGc7DXzqa0TpjU6ZQGM2Rvtwe3IUhN2WSphc33cMwzYUQrqrxUqUk5S9VvW+X9PlZpq7HLHALFj
fyE4E9rcWsFmJL0JaBvXHicmmDENLR932yf86qaTyVjQxxhHJt5fYcywOWnqp7XmDO2kzk16gDtF
iwEwa7R7N0GgtYnHIPrtV1NWeaxnqunU4wYByF9XQ4WYeCcyBstg0NrstqFTDmAyJFbG9NQPRhoh
dzMPZMFrhLUCfz2gs0ks9og+Spf3n98Nkve5UBg6DrWzeFgi4RC97ODry/xdX79Ee8CZlYerSlsF
gYiFdWSZ43SiMDlgv/kXDLMTkRF4KpJgoIvb4LzHx0k5GA5eX9wvldhSoO2x9MsVZcJWnKnpPXzK
+S7siGuLcwHK6jqsKXOZdbY9UHKuJC1n8v7+sFjtbICPXSTyLHkGbxPfnlyBh7GQhY4ROCeic8uC
uRqql74eMIJJ7j5Rofp+g6qbnus534vtgUNfPOybMDlotp8shaqJHNjx+dKTDxR6ZP5Xt50qHaaC
XyKgP/3DW+M7gZG89nFps0uGANOWsa89QBrMM2DBUH5lICMU20zXYJQP56vvvuBXYiA479VidmYK
JxUSwh37o93cvAwj2npwlGAhbNTX0KOqAd7WiRFMSDX2ftd74ONxuInQ50lL43W4GkXzQM8BK57E
Ex+NvYZg/a0ALRi72pWVWw1t+ZmI5meXAopORpetPzmsZ4qq79X8dB6ZRYrZFWgHtSvBk6MPNAYM
35eiVMUSwVozfe6znvB4cyvbbp7iov0IU7wuUPXX7hUe2eb90Tc14yMkLjzPL+x7Hwd2utCTsASP
0SPHGRMhQ29f5ndDmfO8IVg5DC0MaYI5OYktFYa7Il4crU/mNiFhFCuiP2Yv3M1NFwF2jcEOEwgo
l3nz2Kti2E2OD/j7SnW9U9Kima5M/yWy7LZapSNCIJiLzG7Os5jPN7UGRDMzQRnLHqxXjKu1T0IG
gT/72m9/5O1u718ah0eW3fGeJ/qhk/k7CqyjmgRQG8IFSi1w/R2CjijqalMovrphDSGGFB+2nbgo
nYpU5NESjlBlqVvtVbqklf3y/mN7+tr0v8S1fsIF/mWzFdoXhxF2eKkzpbadVwNjJjEwxIh3YuVT
HNjF0Y6gO90R0U4ERdxtOkpOp9VAUbqH8QWpXEgcJmKINhY4i42PpN9HnKFpxpHmLE54c9QFuGi+
lhbzwQqyZrCrIblVHEYkaM1fBTAN38ic1IcYjdokqAhPC9Vr0vrAIj0GQLWRLe0K21wU8kK+23yz
qKfZ5BTW6AVaMriysQsb4VNqpyboAo1nB7zLA6wEnn6ALPWMydiFfCbxz9YAvn2tsoV+gZkb5M2B
Oc5pcdZgDvvQIh8VfboPSOCj5W3W9r0jLU6JgaSLpWvBn2zsL8tksDUiecS9sxthPrMlVb/4suS/
azorkEh3hMN42mipofK8O9OYeKSe1WpyaNVbk/NcievL6zOXnyu6FllLhsNpXyE1RzhTOcg4rfQQ
2snC8FLHFTq/tdrO1RP6Hx2ypDa2qhFwyrEaPjMIqRICXX2W4Ox6ep7L5r4lgGbX/D+cCYwj5lul
rbJ437xkjERGtFcAd41yhHrZ3iVvCTqIXp/xxCvWyk0Lq1qeUkFAwSWEGRVwOYlHQZKnlRucdW0n
rbe9I0u61NFbw9bVVKOHroRzSFTCMHziFbyrGM9PpAt3+IiSBRNsCkJvKAejwG6AFIbzSVFNEYds
fQMBFVzflIS62GQkp1XvJL1ALWDo/stoKSMp1YiCGuqtT5MWuzTOxSuTfV3xQYpDf7L0TMyiORDL
9YdP9ZNLE7x2YnspfLHioHV/tQeffVPyxazM5js8fMH2anzQ0FZuSrhJTurhcEQfFh5+/EE/bLdP
qXXiOplsTubiJJ5mb3ynvGWWNmDnpLr16yoNcjInQ0sSjIkYyuvxYt6qMp/Hd7hVCnIlCHU2bwyj
wQJrxUNwfn+RbYmpaXOOySXJ0bfh9T9OGQK8zf8VkZce6wOX8GQjM1bdZOibnbFJuYVAGx8bcun1
U+Unqj+XPkiaXUTWV42pvwkbN8UtMqMXYmvl/lTI27VdPoT+D45KzkzB2YulMcPHDs394spYLEaM
S9cJG8gM7V5+MEmZaCgSwZsL/BP/o3VZvX4IaiSZekVRdCwDczb/JGzjXry93UNhtiiB/Sz2CRQ4
OIlFoVvdSXkYlHv2eNk7JEEJaD5zzUioqlqGQgCw03H8EqP4yjxYckwx9OJROY9xFPtsV0lpUPfN
5hGIwFs21YzDwe2YIMfa5MsV78+B8+358BVS3F+N5V8O3UyAn2VDkF1GMUiTmuvLkVs419or14jj
JHmdutRgSoOnK+T15GoWUDWCCb6Q9OpeIKKglMKpc7kq5eXccLzO8pEgNkn3aAMmiWIQ5YkE+3c1
do4d3H8qd5QyvFsYXWc/GuLe/iOGkx7L2PyczGeBid8EPJlKrG9wqcoKi/CIY9cQM/MmRYSyUsJ7
71lsyizRd5UDacglIgjbqZgDjBi7wo0PSdANg/5O2IE221MSXUSL4GkbhVApvaCRVvSqlVyF16xK
Q406TzG3S1dL++lACC3wGRL6YDjB1mSzh3JpumDNht27pXQ9NmbB/7yZuvSHX5Anc+tPeZrS6SgZ
JNbGDJNF7o+KshQBUkeeXixzwOoVofJVgcmokFa/k6xDIo0ZZzJiE+T9WSQtMDanTGD3Cd4QnmeU
MuURnxTwz5AY87ZVkSmzBjoWkl7aNX6VKR9LV4Y4LiKLJnJLiUTZkjo4co/Qf2kz/Ab5RuKh6rsV
0W3n+kpc6wILD4SwVf2o47otiuOnoGrZUXgkvKBI1jjiWtVmbqeAA4RLgcQ7NExeU/e7jZkLj4yg
HbraUrbW6pGiJ0lIYQe0UtBrPB90uM3YDN12ztxYxcQflt+/uNAO2VMB8hfyfFLtcLJ3gXUnraVF
pD1Hn0sqJqOuCdZsK5ZkzDzPccvZUjy3oI4wK1DuQAQIS29y5N+dlybKfqzjF401qrt4vxcqjVFA
U5q256rHa3z21XBHAv/wt/MuCYLnX1987ZrJdvcFweVIFPTZA7UmQWghwjr6uMF4P6p1m9+Ldcut
rpBc4eJNSFSusOJRN1FSGIJrSlflolJTnsnWAL8vtbKdaudcILyLspPBOhOG/fYFSihy7f4B5Jhp
a4nkahJFo7j4/wyHSh8IxvdFCEHWkE3L+0sdZhQ0ddJrpDmaPzHDvfCx9reSq6AWep0XzgulU6OM
kfouNfacBXYfTY2G3UJXfifHqSWQXsJdlRaTNhwUJ29lXoBmqQe15nU1EAh5dHytV9FJBwbE1JRk
5osCHpGYhMDDlbBTdViz9HUlsq47wNy/CMC3Lrk3Y6dqkpO6ziydBOWz23srOE84Q5AyT1OGkKxy
px/ygjDtAr+irMQajGYSz4tiTITIr9XPvOzSALrdnvMPZeXEvRnCZbmWBu45tkv+6WD6OfMipN2a
TB9xtpIB2TxVVKNQ/FPMpFeL0G8m7Y1xTHzajAz6rERXGdlPaZdpWk/SDJzUBF7dQECUJq9Hdd5z
wv5bUn5Fk6lkX418m8Ba3rYju1/+C9OXq7l9bvMFR0kPf92hL0frop5CBeD1mZOaCe0ldydm59OT
mHzgNgYs1rt5eVYj+Jn1VDl3lJU3REsHqZpCI/Ui71WVfj5VHO0LhFnsbEl5+Lq00NynUf8u1mIY
YhvbPbv7w6/Kk+4GEhkCv4MWvQsLpzFyoYgJLCX+K5+jFms1W+cYKk5PO+DVcQkirZRAvZQyZF38
EWR4LJd8VO2oP/u0tNr87m3RfxToKmGVb/doIJCBuqRg+zho60J3gUOG/K6wXKvtLI0XM9z9R+yW
5pI8HZb4WpnnJ3ioJhjJ+om1L+ZucScWuMWyAzh541lPuEQh81MyxGNx6tmVqoHUkErvu7yJY3wS
pnWhLhc+LDf1JLVHwGR9mX32qMXOwP56SVLzjbPS3TwEnyPrfkPEwSZL7Qcu/M6tLDSKcxigHPsI
KK9HxHa07YA2FJ4T9V67yqD5cBck+lKdMERvTGmyAJg8QL1TnZw5eyhTSeDlFLZhSVp+uBDoWzm5
JANWWb0m52Fyv4NuYY2YMiOoCciWfCzPiVlgnRa5GziuHTKc2r4YLtu+f+dSvJqxYIcCqqt7cnR8
O1bMl22BSNcc8Na8gV9dko1ykDw2TSxw4votBwOL+yRqzibAseIrCShCHMUJjV8nhdEiprWFKu9T
XKFKMgj5j+sTckdtEGlKOYqITGzkQ22MbWM04prVDGw4pDLIKkDVyk0yz7CbrOB3k0l/0jkIO4Kv
63xpvuz5KVH5Zu/MS5TlJh2ejLAH3r4yfgQmghODS5E0obg+IJ5SZbooqigAnm+P0hjlOX2DJqVG
MFGeOfkC8lfT8fV/ISch/sptMZhGSzFye9DuS1sgHdp/kMir8DamcSU8QFSZVxZsjCITlyXPPCAm
r72TY0QW5cGvu2u/YaStb3p8NTaDVPL8XtGJPVYkK0dO0o8kjMIyyof/3y7pGfbUuUWKQ0ADBApE
uYJp17m7uw1FBAJc5eU0dNy7k0uBI//deAYLuhpR1s2X679pF5mgIi7FRZNYkPn1Wab77TEa6Y4I
ANRNyXdsBZRLEkjfUwkj7+4/HRjN+6IxISnCDsxWdQnqg5qplQGAt09uhB8b2/7d9+70rxu5p7kM
6A7BQLWGGNEzgSXg5z6rg+PB761gwEy7MSc1AQgI4sEeEL0KaNxH0+jhhmfukewNjl8Qk2OjPW62
atd0o77NNaQGSAUaSQUNFBLOn0+qpp5qxjmrLujL/8dWvcpCkcc4UWCCHRypCD3hpUxbMiqbNvAh
pdgdA0mVA4mRVezI4LkAqa1pViHxtx42Y+twAC7XSv56fJPI7ePCbwzYg4pngvl7rXYe7YDGMV3R
Q0//iSkMtMPevBCsp4/mbrY5Hg4UVhZZNWYcxBOUNzu3sdtbc3gIBV7E+IzYqHuAk47BuZPZYwaQ
/4E8dd2FFwgS4H0CnIMPRWt1Sv6mUvaiKai5fIuqiLKSMqELpkGdZe5s/6WtX5Y6uLqV4xVyykVs
4tfYv3FUbEB360raPcYIlAlibe4aSDP6ZFaXRw67cJq+iCY0kdUwohpwKCvvts1Cuv015/E40xqu
C8aXFwJ8VMLvqJ9jqcq9ZekYba5kAxJMQApWwclP1Ke5kXxwC1BiWOyhBSmV49mjmsVc+EXVHUMy
t8jIs6VnS60CLqz9fG3ZLxNHMUJLLTcfM4jlFlMDB11hPqrioFDTlUeTCnZwLkCWqXmHu5er3nHa
yoTmqC6bDjREO/7+7npGIkgRfR2/RFgcfpftAvHiYQBw9sJ4Ewc3NYVl4USHkePag1FoXVBBr3gC
0CYTNtzUseyetEi4XdLC8vLXPZDW49aTKkinBYlIqLTVXxhZ2F7urvpVumZ2+8Yjg29VZVsZ4v7U
z2pdYE1a6S81rjtRZcNrO/gVgujvd8aJtHNiX+I1XCvtXyIHROGPKX7txXu6nQpIcTDTFyYYHO7t
FnncitL+ZBVp/AMUHvhY/SOrE8TS7MBYoZhkHMw2Bqso1fHhBgs5BZwpIhI6Gsm/upXaZmVan+/Y
3dv/yZJ7UnwWfD9nQ0oiMqiG4iBiJ91RFfb6s6qI0k9rnHvZhMWTKQhR5m5vWWjzYRsAxRKi1i/j
XB0dV+oPqSULVCpPKWmuje7r9O93ziEeq7h2adB563U/VSBk+tdTq/ouV4BPdi/222FY8tFsxv6G
T4JWQSupYeg+0dnZcfVxFstfMcgTCKUl0YBZWFZ17Apw00mKmsxDh+/aejEQNdSU4wynHsoUbH5y
ED8x3fiGktubUrTfXKlDqQfC3k0CZ8uYVo4v96TiLPkmzJZ/t/K2VMESUrMSCd4oMYd+jxPLnRWn
89AmJ0YNAh4L3FsN81U0uw0kaXcDXAbSjSM5+R53mIjZlEns+ATK7xPJ7J1JvlGDYO/L29xtlFHA
lBatpX2wc4NTy8MNCltvizExBTwTmfdqvv3VKiU8rdfaev1RFTS94mBwqiHoDaORDCYQITH79Nx2
SDS6C6VQqSWqquksVe1dGuKKklcg3TbNULpSmikkyAXll5VHbeZIzAx2Yt7Xepy2R8AEME4HyIGR
R+yp6a54k2JjCophv4YTFEcfVN+uAn60wuoJBuLUoXrJ6ETUYzLT/26vi4pWihBW8ma0+KeynOCx
o9B6uyUiRUOUsMytv4cjDQgqkzTBYVhQT8BkpJ0A2RWt7z8siOD+GcxTRX8cCJArdXmLx+f35uI+
kghUZEA3ZclE7i0x6AEFCZgmT0YARiUsUEic5G5MKGiP02M4/D3nEN8WBFqcXiC8L1veKfxAGraj
LsMpIp7mmFvbRSQ70BmL/DXarIfn50P9lqzrG1zjnBITnGETq3EiuPi0rTM674zrW8gSNzINB+Ba
7ujdicpxOiA8Py9a4hMb7+rGsU1xMU0S21unw1oI55Id6WI2AXQgh17BCwY42uOoyFmb+Ua8F81F
NWDmVddQ85EqpKiX7DuUF+TK4j3W/KOAleMazZy7Xzmo/XUj7KPJJGXf/zwy1H7XiOUDGCffsr69
a7LovzYM4VZf5fy/SNBPI07LBg6Q3gYqiz/qRCfPgGH73ziymxLqllPbLi3WYYw0NZcLPyoObt+j
XQSx0sBQ8VCqpWuGigb1Ki5Y64L4cRkk6Wdbc8RC5XrU3cKiF/ZWjAkgIgtFC/rF4umU3enEnlXi
JpnO0dE04fkN1xucFwpBjw/94dc/lRN/n2xeYtdfpHZgL69CSAqfSQXoQ3EPK2c42zSxaJV5NzpB
a6tQX+guNyQV/NV1nyOvX3yKSXBBJD++u4pBsSyS4SKDCFNWK+ILpjF7RcBYxGFAk5qzJpC2ZVJF
xzDYIAWxSFTNipEPdq6EgsXzwio/cUh5fWFcFzcnQfLWSPfF96ZMlZnKRvnJlxNY0R0FrWspC0bA
H5GZxyQq+CKCOSEm49v89TBQQDc+O2Zeu918LdFDi5oQbXfwUN8BST1FaMNsGuuunWNaDHlSyA/W
geIopjL94apz8BNpUOK/4XnBRXVBWJ+laW5BYLnOaPIWNQv2HP4/3ca4rGchDumgEF7uotqpuocQ
LWRPJz8eWgyHVF7CWpNcPBIOIwIZsXUtpFJOr4NrX/ZXKqnIQjxVpkY++RL1vriQZ+jlGLp3JBLB
pOFG4wmz12f2a5zAfSbEzbYgUc4Ak8MkkGkZf2gq3Zs64NBBkoPo7Pz42Tpov/RiuRKzL5M69ul1
UYqX/ORgItc2FY88wRb8h6VxuxSROVG87t48hrw5qhctlg9yJQWiTRoivaYYRmEwlDxNeswrypYc
EMychlfSNVNdFq4oCmgRhWr1iawEOblx4YWCKA81q329CtFGWNA1WgmE6rpfl6h7OfTZ2NLDhInZ
dWj4pC4S2SWOSUHKAoFYxX7L0OWpWqZ+ehQ9BqHGFhptAKDZCnj5KKyxmGlztXpQueeUZEAA8thB
+6PSs8lraL/85gry0sJDT2PPAIH1jil8SldwWltou4pKAGviIwI6S0vRwGG6CtJ3LvhqQ29+FcXj
pNPdSuCKzKhU6uP6sIIpss5gC3be9jOZhRO2DakH1ooQ5zhAlqFJNoVgonTCevfxm8KV2CldYvzM
KewZFrcyvm/hPWWaUJnFfan27Cvy38eLSmAbJRd9LNqnsTe3pBg86TdUrP0ZHd7nth7flqEl1YL+
kt94iysTe5EWr54OeHzXlQ90alaK9sK3C9Cso5qvmxRtxiGZto90eGxIh/IRJJAoO1WgYxSUWBuN
i4/3OT1M+1FrF92eOnIz6zCDquEr7mamizjxERoKEiLPfCaRNT6Fs62hqzwDXwn2JAY8Oe5NWrto
epEBUhS5ago4XoapBVlcK/m+nSr7q5yKW3qS/xWeWTYCX5l9hezgqW7eRZREbnAIND1mjpwXBh+B
L7qi7TtD0qkXrEdEBs25YhMn0Fb8KREAXwHOhkOp74va9IG+54aTbi6o1Keki19m+RUuyHPPCrIG
0n3O4og8BICH5mb5alb4aYWIQgu3lHEwujlzvuDRunGjG5QXYPGsx0KvBoft8lYjoKdkqJDk2FRC
qsW0awuggAlKzgF8K1/UNBR1zSMY/jqQahs504Zj9gazNk36W7tRAfN1Ffujok1TYPUXnTnMWLVa
2YhRzHf2pPigV/C8DvE8/3NgxwLl42J8kBVsQlEasiCWrkAdPV7IlayjsT7zZqjyCePnZ9H+jap0
106FrI2D8STUCREsrkzv1zq4rOMZDr4EDEG7Q7vHOJ4q/PZ4/fkJcwMDqvljaqQFjuOyd/UguZkh
KT1TD0HguKPK1SGlP8BiOGMD0l5M2RxPtHoUeQlgmLdNYuLnjUTBcrr8jlrH/NUyZoGKlwy5qBol
PplcMlAhYgSRvYbhd8nkdvnGELCZNfrLzBWklum7NC5nxRno4zINOouLIly7TfGPua7HusboBzm5
F0Dbkq3gbdx6aPGes7hQFneFvDrgN2GA3ZVv86WdD1Ps+pCknu9g0Zz+/TfspnsHe0xlqPwOpXQx
8QNsGcg7OExmZ54iDqzPbM7YcqCYjhgp28mPVZcefd51RzXO4WSW6+MQarkaD+gDcWg0SOxUPKZM
8kims9SbZwKDJiESJ0ezXAT4Y9G2Sgtkz1ekVQvXrteMCnZj0FcBu8Yl2/0Mx8FzTGslngelpOkq
mqD0rAp5VwgjG/VLmNLNmEg2njWTA2RNe4j1Ta9aVKxfJWj/ycRL0b+0XY1fEGraujZ8x691gFWJ
u7N8zNLVMczRKkJoIsX22aRbmb6GGyK5KH+nO6VkmQXBXx1AvYgOLw9Rs6vIVl1U7l9OzVgJEpic
2GV2j24uNJ3h1ciCeN1RUJJnGHACRemfJf0A8R6TZMLIDhH9TUGWYhEoWYsMsMxIH9D5VxIzsxKe
lG02fQfoqly5GhMy/kGACMQKnGofdx5j7uL+pQ7RyBLjRv29bAXn/dkOz6ubZAv+yvcR9BMaDd5g
0jVTGjrSHl0/Fls/TPc69jQZkyWR/gd9rui4JXF1AFfrphwgjBDXk1yKF+f/TQjH2ZHjSdHizZnt
bP8Ba7rEFrPfbg/kf9zHC3Soh5dPguIxg7b5eP1SDjr3pk0In9SeWtIYm17PVarNalAr1f5rU80O
v7rYnlBj9kzRU62ndgipe8FWjlHb2hYK3krb6q/IP7f7ehkf/2vv3+sLv6G53Gfkjq+GAItW0Y/A
FPeCIAJCdzMoyOzQgF2mYR8U8htAd+6t5AgIaQ7kAnxLikF9q+hm1l0xb5MefLGjstVZMVb1WW7u
7NshU3f0sYNYYKkSv7V4QzccYNpE1SntexhfxLlyvR6iq6sFwLA0Vs5b/j1H7o4pAgMuZ7fOFwYj
uIYR51UHpi7enNXWfoj0c/0pQMnN50BjCqNLibYDIOCAZmM8VYu5b/fQaOX+PpsBckW45/S/yJZh
XEVIpXYPgOWpIdRsGOLj3BuRLtonEjBC1vgJ1+jhWe6NYJXQw7TVaiiGFssyBmrv8SYu/kcLE12z
lq2fd7OJfmYmziNd4vRooYAecpGErtXPfk3VFFaAxCUUMGVjDezfY/3b9s0MLjkP/bn0eeDYwyeW
VyBJoNkJkD9bvG6Dm7dMqlt48pJJEuXxzr/X4w4OOx1F3Ydt1bSbaDGPuAWBcHqjVWRPzEL7Vt7P
uHFkPNB4ADZsHlkqlLkk1tLOFKPnNuULkMvM85/CZGKAMi+ljXT/QhgavDhqAl5VJT/BHAUFPtNu
NtiGVGfQCnFapTI3cUoMX1slpBhjFw8wsVFaK75/7eVeO8YyntMu54brlMvlCt5jqKLHzY4Jentj
4nUNqSuNtuLb7vQ5CiZMSw1EieaX2bHC+Gfr9LUPpfXLnGVSsPt+Z1oYEpJ9B1umRo/DUHazWUbD
cWw9xgTmnhHyOLALOCvjCUYfqIzA/7kHmnIx5lt8dLPZ18cbt+3FrrHwOVkX9wZpTnQObO9KQJT/
iEA+ywiVoiqSegxKhWjcCs0I27SZNSeFo7E01wDPaJDsb79fw83oDE5rdWIXS4cX17K2+DFpy/VV
tvTN8W3ncYI3mKkJfsuFLK3oudkqrDxtRmwMXTJokkLEzoU1v4tZT3T7uIKpqZc+95dMWw1fw7TD
zwjcxLEfQr+dRGT2SpNefjj49lh92N0TMai+z7HZ/N9+t0JSt3Fy32zRUyAeCWsJQU6VGGCCyLTc
sB0ebzhHoNsondbf/yG0ueuLBLiJ9TvrRv6+noQww2P8nvmS17EiDBQFBUaXsJkZrdPGZcxa+TL6
9o66W/OQFnNb6MGbTamR5QL8lGHtSns2qyYKrbQWL6TBt3wpgIQdRQcA4JrqvX7Z8oavDLOBcpgC
yjyJpyUNw7Hi9QKWEjLIISUQ12ezaeZnJ0RKka+acUehL5LNm7mwZgELViqCTqz5fDVCdg5XHURd
xid8pgiD1TGfkfdWhR4dPgvi0IUIpleNL/bFMFSqi6NXCi0pBpcVwzdcYS6D0q7KDrlZTwrGK+Br
DEfr4+uBWDtyRthf6o6b//sLWg4X+4mwx+GrcwNns4QT+jb258L9WIvMe5S0AOK2wi8YHcC/4KWI
W6Z+9UYvD4Pd0cL662MiWm+BPOHZ8uIhkyS3GU+o59uz6Ytfv5NbXUXZhunPQP2AqzzhmAdZ76vk
VfulKsol8c3aRA9X1UKGTht3o6o2xXeV9mngtKVyLBpsBO6N/FFsHKsgzDgOuXL8Q7xp0HOtMzNz
mhbpRY1bXkydkc5NTX26ykCrIWR8JZe0fnUepwFmm0+hVihQCl7qwt0ZBfU55CEg2ND6yXmcwl8d
5x9DtFYsrd/kn+9OEB/Dbgo9nHEZvTxUL6zya61maaBCgipKst7+FMTyOzU6ryuT9WSBmXXUmT/L
xfn1nEQdDiLfhmySYbfsUOnnSV++X5kFL+nckaoeuKckkim5/7zGbcil0ALgkZ4PTYAeQFObGKIb
w+D+l6NeSPUbEYi3ha+uVckIvuSnKalfXid1p2t8X0C08fz5YVsrx8swmjVVhKL3STz0AakvC/7E
3f7lr2/AiSVLEQ528iGGw/shwzpoI71bt7ipa+lBxcKSS+A499LH145qtSnFt31d/6o248sbr/8D
BHk+wbbejLyod4NN5JXY8WQgIwsP6oOLouiPd2Vs1i58Q/+45tI2lpNR8iz+1AOH94RN4rPbQ2pC
3VxCTa2TjKWIdn9eGlVL8ozxJ07EKYpOcLL37PDbkKXDOJf2mcohKFQc7PALod4LEOqeS/j2USKf
ErenhtPNIXfmcswF/0DFbRgE/xGp9DxU2k9x15J5bhzv0k7Jxlx0s37f1kYbrGnlRJGCzUlznbgq
+w/r0Afr50+iH3z3Jnyn5Iy0qzVp5gsznnS4+XZJl1D/0AGQvfJK40JoaTAOAWam2VMaTltGl5u+
LBI715cPNg0HmP3L9f9e+lUqLK2U9W7K6aytjGMCjS1ZA+jaaK4+/fr+EYAM5inxh0pJ3MMpl1Qn
pvziG6av4++QSN+ewFHFXcdoqsun73LAK4+47iu0vvn3fQQnNxFX9TDjpR7yvDUq0u2uqpZ/PeSF
+yy5X88HbzsJJUjmOG0ubIY7yK7UiF+uRs+0OYeEOOljt/VazxXulqUowK07pf3l1xhmjr6soxSy
/7Z0L1I7Evb/Ei3UQwUk3vzbKvv3ONA04+Q7Q01SqAYL7wHlTK//uPY/m6FDoqVynbXTZmM2Mimf
YRjK6MwydlaOdkLdKaobCtI/U14hnMeXKRPU0v9oD6fEPSK/wt+mdITAHrYiDpfwfaiDdqBXiJ6l
vHjzGNy7dP1GmFokCPitnFtJFx7+IvRVon8z0cmCD+6EQSYl2FPfrNSFOrAu8wnWcOGCoMXiKENF
KbTDgsN7J/Wm1npPwiPEH2gEt6LRx1wPC+PTT3HCncqISI7yhghE+6oeYQ/Q61HzsgFSsgHVqZqK
5WtHMb5clX75ZFmgFgq1RJ8RBaGcXvgnSyo2JXczo2DmLH/fPM1mFvdInF+y3ehljITHYheU5y9V
+8H6HISJtQGdGNyqgjkDrOTGv8tVSfl2cM6QPfVIcvl+RxwTZOpfUxTifsnz2eJeMR/fEWiyeYeh
AqC91lmWIt4M+4WmaCIaxvpoEWUv3XDZbMybykTI1p5WYYNx5/9aFrG5eLQYZtdVg8P93ZW5/Zub
o5sCVXJqpuFmubrQWivrWxxe8ERvYnHrpav8+5fdUqCb9GbPjl1l/VRaLux4xmR80P0m9QT3y+rN
oPbl1NDPOdRbvOCmnupyAlmvMXFZNE6r3y2FRpwLnIu/NZPFn+s5uhIfiS+bVpFFMDvciFYmT0aG
b+OfmbNAUSmN3K3y7toJxJCJ7xjOA/MFZT4fg7nRDlgooglkkDMqiv1DUS9vOwwb/D5frUPlLLCP
NkaXj6k913tfGqRCP6bkdKcj1/ew859A1vMzUaN4nZNatD91WbKHVm+8jd/dH5uh2xP31m0PWFMo
XkXHklrwKdfB9HUp5SMiabmcR8tWsUF5h+gwHqJxYAOg1BsTiF7aygPYAaNji1agXCliD6GUVujv
30KyhralNz4cZs5Rw5kRxbcNri0HT9hvp45NbSbUpCt4zljqMOVgf7L3rKaWX/T34+wDDgYtU74X
BjH6sI4aQC+fQ0jWZmE6nAwkWKf/yXoF1gSxsn7g/DlR2KML4Ihe0NWKTXKkp+5IBsAeS6WJQrt9
vZzxmw7bfpwSMDv5/8A9zITBzdPkZ5WWDXDQox8JQ1okyklsAxslM9z0NRZsOb1ISvd0ygnbgI5s
RLUP10JZcQLMyXjuYqJ3hJolxYbQgx+dji89mSTW2XjZa8CPgQGstsKHYPCwc/uhk+ASil+azy+n
7e+yV1jnE3SAdLPuahd5Y++mLwM6zcy4o1oof7uQdnDgUXTSMB9sjHvqHLm6p8M3MwsVWDfPGIo3
zI/LxhtYJhYtNJoSKaCkG9r6ybidwW+TSyZSrel0d+ZfKY9xvcalecNL9A0loTnGVudX5q02oTE/
ksRatHCKiNWQECG7NZIkxt3UaQKaWi2ie5mzUq5XlSzJ52OfWAPkawAQOR/0smzhWAHQ0b4EPVXi
CEw0K+9KFTJB/V+n1qZ1YqvoIuaF7bXHEUWNNKsr/btixr1dxwTz71IJd1OpRN646G7ir4K8JUgd
eFWeFdXNQIxpEN6pa6+O59Tn7rvFkOwNill/8peAiuZiKDHS+9tlSVnceUKxbiag7AsksAX3CNCn
ovQj7RMCPlFbUYSKxurwF5yd6/Ya/jSCSRHASfqFqqQNv/7QMCXAytBrlECEQD+6UxJKLIIHyJuG
ipK1vREoFnNySPUMyx2jtKzVd3ApRWTCesL53rpD+Z7gfXDopSdSLFZr7YGbi3rHNxCCUzR5XvjJ
2QLyFmwsrRdcQEB0+dYkGQMPaT/ITpJiIyl6KkvxsQIVzFE+aI6uoTwULt9jUXMpxP15Q1HgJ+jo
T+a49VBhoCB2N/un9cRomYO1Ie3VsXXkiwvFinFic2mRc/a+GsOlaNuIAJ1+XRKDjhrdNqIlncRt
D2slhe2dAQm+fRYUT2WPQLDQF4aoSxcAVyyraR6rELiFugpTR28vxuLdSppUCuSC0s2ej30jDMrT
Hvqpn/5SpD41T4LKnSH/RX1AmhnR7pmUGldnMYDIfBJ2XkiZifEZTEpt5pEARNjiXQhaVxWCvUFH
r0wsyNW2ph81HaMj3D550APdy9vgrvwputv0a9XhbR62FIx/I650Y+2JP97re7e7UEE0VMJxORwS
0wxJ9pLAAipKdsDvfnl3T6q6sMFOLPY2+wIX7rtAPv6/G875tqPGMmKkkG1/4vxJbX4oN9u2y6Bj
u5r7/hhJIqCD1Vjig8+xugQ0thQ/7P2wm+QzwVBa4WHu96ITU8TcJzgW+6neDrN0Dzi4FbKWrINN
D+K3chKkGf35wzZF7SJc7YtT7/6JPwY4A9fSw+xXO0OvAO8zB4Yts4ufRqpCdhjnBleAEm6ntHcR
m8GzvLtF7GgT9+cYgSnuYndsgmJquAS7HHkSWudYKNRQESN1F0aQNPM27rdhqYQJz5lnuJj3N1su
ezySL+49ovPP87gkv6BlgBmlCDT8QzeBT2v8lEBwfMW8rWZlD7kBP+urH7UwjrNAZGhhEG9ooyEj
5nEpYyn5d+/dx16FXZ7/XLz7lVFQXb50lEy+SOpHrekFwlzkGFmI3WpvcrmZ7qdNPbVNi0HNKkMb
W01Gnhc8RewE22E5hICASUtXLF1V+07E70snhT9Vd8nVeAjfoMAiZ9j2+X1VyfuCI4N6RBnYrn3g
ZrZpV8IDpghX/DTDys3YP/ggnrm7vft/aRfmEmvhmGqI+KvEeOuEQAh3h5COCQYJWKekEzVIPAq3
+dcDlUKdpQ4nwRzZI0ZPrPJqvcwrcrcI0E4+JXq4FloHAUbOQkwmKnjSMPgWE/sP50HUS6vFacCV
a2dK4V6miGxKLhV5FMccBugR5LcaAFqRRwYgayjvJPFH/XqvIlYcZirG6+ov/eFAuQGKg/8eVFAe
qabfA9JY/CVtwa4+1LEPbzmHusEVMh/nnHkwq5Ej8QX9LMvlG8VzbRVP+xUzKPmyTVK/z/JLfsQ6
KfYdPZ5sETxunZ6mk6yxTWRC3ewSm6dXc50JcaeGB7H1FLNp8B5PjgZcz/p+fqRuvt4jys2yeIUt
qLrsRptp5w7SDv2ZVOx1VApzXUVuVG9UnYUfeKb6zA5xflxp5bti7CFB/swx9aD+yHDmhJXQUtV1
Emb6ewGNUTeOdoi5W3xMFC45ZWRL8YWD/MiFpUdJGY3PcrtO80owUHdlY4pclXPamalkodxQ3pG+
up5OybrAAeAdqKDAWw8bNCLZ3ZqigHqij1KkVcDD02BSzx6hQbZan5CXRa+AVSMGH+KND0XWux+B
TwHG7FR8FeLw8qflDb2dPKomQZ+TJwCxay6M7bIv9rmGY6J8oQlnSfdvRLd2wYXhnshn+M9G4bY1
mHW95Hvzmsga8cDXaJDNqSbpHiuDiLZdg7dsPKa78Uk8gSdbju7KidVOPqPt3hiEb9ktj38VarEW
eKBGLiCg/m2N81s14thXVrea6X5vYpl/muXniDqupEVOvibOuWucESHt9Ai3CO9KUZbMBvcElems
anluZgz4orwnLOs6v/CQXtTYMf2jmb2iSWlzZue7ngS1uYKEv/JJ9iBEBfdQ22798QPPoOxrbDDX
hxE/8Uo4aD4VTVEANLHjQ9gMnN98oOr4UDSEa4Cxd+ZMwJuFOeZeMHTNVrSkoMCrwIS7pI3v+m7/
Zu39L0SEnW7adF64HOf1hSjsa9z0BPe2TWMnxQvk8thsg+df+glWFq9vzvzEJt5DZzWCDSktjJEs
XXmQA5YgFVIwE/geI/QNE2dIVkoIYWNBk1b0BrVgsGBGJO1GxsHVYUXbyvEB8RwU2xZv3g0lsMwB
Ct3AohKJRnqvYYA5CQqVCd5qhQPI6dZ+3P7OwAM9Kh/cfNwHQsEWYf+IKlqaa7umW4wHpuec28rV
B6svIPThWBwMpa2Z22yiB/jTUuveET80iIcFIDsNRPXTgAep5UG2QP+awnYqRRqYE/p/ZzkjbXKR
wsKUeVPUnoXeQO7vg4iOFlcuVZ0tsI01jwpjlgX4lhQ5nog09+3Cb3/zmDoMCq+C07V7VIBjfYqv
6CafLoRwOh53MI7RmDcWDdxpJfiIT0Sw9b5eyDvHW0Vtr74j9rbEYfSFDWEAwzu6B8h5t4AQCllI
EJA02XP7iG9HQqjIJd/UG+lnSFxCXCXgSuHdINwgRoY0O5i7B4oYsfLsd50CT9rXP87ApeK+9nX9
kcSk8WcIRmRAJulibKsJKATbBXq70qU74gLsg7iemPgAx8IrQlDF6uLn8tCVqTLmaiFzbVT6mt55
lBzp6957fjZpLbCgPaZcCtHUhZhDtNdkyhAtDVwqfAtv+mEGkpX8cHxvKZWn7VMl5iOdvkNpcTs2
PZdvl4Qf0wQR4r90nHWrVc3I49smQjvyoBqvAKY7l2xiB9Poenl+SiGUkGHJuFOenKNEiV+W9stG
iCk85E7ET+VxGYoJ40n4xMP824hPD3Kp1awcLa33Mh7tFukmIEbdimfwvGbUr/6UFQfn51/wrIeL
R1/6nIK+IvYTmdHt4vmxQ9Rtu+s8O1Wq60+FGv89K+sOVIpqpJ4BXHsOFcqvsUuHwg395sDHdvg4
6hQXpg2/qHKtTwA4A6BUl6fCfnBN6rRH2xHEtGLOb82Oa38T3LzDNzA0Ihw6e5FQVUJig2PuyApG
HYBpUZjCBiqAztFgDiSknBJXOO4g6RYo2/bcbp7Dbhu38o7RXtuWKENfwf/CYnK5FlSE0ZMIViHl
Tyx+0UZL8QUibXkStRb5Iay2w0v53QL2q8UKJuLUdkJu9Cl4ocU5RdlRIlHETpIZ0CkvuGQ3/bD7
fWGIN4r8f+gRmmgHEMJ008VmjTkaeiwvPNdt3gBksJe2/Ue4Emd5U6FHK2P91IpS2dDLWLpdKAEV
Z2rc/vuQFQSh6IBz6O5n5h1T20gZaEi65Y+yFqEPOhhRbBGXSkRqGtmO93vzV/22lWzyei8gmYAf
XP+dAZ4xfdzrc9HzW9UAmThJcQ8IQSgemgESIPgxZxmndHRYO9HklouRM1rrRWv3qqeu14Fy4ldv
6YcRY1iCeE8gRdcAi8uNmDRiuc9RKlbSY2gfOO0pbXwURE5W5gQWJVIGF4hhYyuy6h4xxIo6MJKb
jZfH1eO6iCqYTZ8TRyQVc5BZUp6DWlptA/j/wpGvb1ra8bpBXuof3hzNlpvXS99E9YGDXObvk5eb
e0v69bTk4KBRjMQZHjJwFFJ4gqy2FoKJUu9DTsK2KBBjVIYp+JKnVFzuzNYdOlzIsfxYNbhBgdzs
l7kcwAgVkQK/oby1yTHndMklihpxdXOWfJo4WcDwQZZpEK2SaeoZCobiBeSiYNyGxd/0oOYo+h6M
x/OMZ5FH56qIxXPTouwe6+J+pz+xlgIMItRhdD4J3tN9hGYT97NCvzyTmY/3mNcWKKklVNKVVSr9
naZVjx7gDkpD1chUhgdHBdJu0QAbhB0Ht/GpJCGjvsNKA208TKU/Wf2jxNxgWKanX/IcxP+rG3Yk
Zc4/KoYRMI1y4KM8XDghG+myAflEjQrtlnddAyJZlv+bbzurq79+iY4yxb1BBc+4fMUpGGqqkYdW
8ABuLdsgOQEmQpoLPvuoTrNHEIbfF6rLKsQ1spHMbEh6bdDDhwdwXUeanR1LM4U6aMVd7LQPjMCT
lyE7zU6ZK+GI/3T7TLWIJWASZpcIDrw9vbe1On1NoPB0jvo/vOGQzWLbeTiMz4zvGdrxC3Eg1Jjp
Mk7rvSSMK+0rXlXx3H8I7noE9wyh3EvWneleV24Knb8VQ8qCrLWopQkCYdYJ47PCIRGAU73kOgl0
ZYNzuIREz4kPyH994+h7w3z6/a/qNmli02hinTTe6CcPz/t/OFSAv2xnFmqMwBQgDAX8Jk0I66ub
9viQ6saVyBL0o0a0XOPRNeb59LNxWauru1mqeb7C3zExcoVQOzsCT5FZ5c+AChlQRIojlf0AX8WF
qNrLVH73FSkeJk55+ZMkjZySTxRwaFmG2IRwmUvtN18KBpn+XpydxLK3gSBF/x7dlTpTBX2vJ153
yl9hCTyHCq0fYywa4lnHyVy5DK7hhz+Ymgrwag5DNaokqxsXfu0EV+q3WoywTnq1tf6CKlGNbF4c
woRrG1Ew7gtq28IUdWHH/feRbTypKUJ/szY6FW6pekvWUrbon5A2zz7goUk+LTGMZbVULpw8OkLR
2+aciiQgyFTakOpwQfFsuHrURsUrZIejAoNOLpQQ88+1+xJaYR+a/2MhC1Q+PlidaVaUIXPnVsSJ
AYVn+twvegPLwxov3UHKoM2BNInS7vmoCXkKPbVG2PRbgzS9yFFysOvPc5FZm1mX7+kcL42dgRZU
uK5X8l7BFfVj4Fdo3hJJaxh/eCFHXvie+HNz45DKMrKcuPnLT3RwbW5rYZzfhLY4P4unij0NqOKI
vNOFcMcT98b8ynqthA04W0fFK4VGgeQTY6tiXGPxmNQ3qe4YrA7wFqrbT5VlxQPlepLY9Czykafu
aTetLWQp9C1giS1hvUqZIfyfQSH4hkeLf3c0ARPXIV2GBIWI97ayxDy4IRT6Fx27ERRmWJePXbnh
JWTlnhTYhIiBSJeIDuRJ9xRTwzAP1j9+fvp+iSsdzbOp0voGt7BmntFUFtDcstd3hfgaevGXEDN1
bFqzOmWnoyN6mUrvQcVN4zrxC6VV+uKvVDzhBnfk0Fkjha+Zcwce1z9pjgnEGUh4FRVil08SAz4o
0muwOZY+ASP8YECTh3+w7Kafz7zD+yL5oJCo3ujvHhqsFz/NQB/Ogg1P62D5RAZPzMfjRPllCXwY
dDaVTwUCpVgg27foV+Hf44Gj8XKMLAs6g49TRinRBXcwrR7dLrB2URJfnKQy1+fxIc0wJFuYXjl2
eQX1Be+QruAK2BDjRK2PNlTugUrUu69BHx4wTyvPAgaFdNzkRJ3ON0lGjyws4/RTYI1z1t0F4EzS
Mft5isKd9TwBdmm0VFdRYjQGtttP8f17vgP48qbFJnzKkWF4nUQMH8zvp4uEKotXWwUxuklfdtC7
BHZFM9FpFm5E7SxGysruouHu02eP8MxQth3KnMpCv77mx9XojKpJDeJaKPhoXPFogt67hn0ZMtKh
PWuXNT7w2UJ+Q6FZKbu5G0c10Gez6UIvfdfNYtUwT9Sn1tf24qpkPP4bErFYOmUzeiiOZ3ZWD9SN
6ZUY/LIx9iX09lyCHTiVa2Ip958wO/w2zOmtsB8G5BpHrkj85bmSVH72iJk8MG51kqIaHY7stwty
cP3cLN+ordBwpY1IbC732w1Cq+5WDCuT5Ubd65aQ1/4UE+Q6+T+4vQPbQSVHnbtYad33x3t0+1N/
9DjBZhmbh9aE/MpNwxCriUHy9shrm4VD35jXVkyFmyPuU3EL2J96lW2C70SF/b1FBBUtl9t1Quh1
GsvtXMpd5SpM/Yqb878SziNi7va0NjvbHvMMGSiL17Vp84zOZhqvFACBXQayeDA07ILfr+5cSlzv
i9tlAYge88rqcRMke7SdH8Q8oViTAYf2F7xHXX3gz+aTTjgQvTG4co7s/P5Tet8CKLsNoSt0/AED
8H3JriKA67Zj3BuqIB/t8JlTsSxtSuSubKQ/3ADDCCVoC70pKIX3MB7qQ6pBivJ81WWEINnWteE/
nOgrKTYOEmvq9AatA3Q57s1PVV26AHfqpMbg8mxV3jJZngEC6c0k8Zvm9IvSzA5d+DirHqTZti8X
Ar3Vesu8FWSPQIac4bw9d3R7CbuWfhaLbDulu102jMXzKtxmN14bqbT90Dih5C/lFFPKKKG/ANM7
98HBg4gPx+H96Dy7N+3KWzcyLtI4YZCjj9oh1mUBcvgHyW/ZvDxFZVupLj0N6/4ayBo7HM/4jdCn
/cKSVLk37IwYrbLAklOFvjsw9sUWq47f09kFufQnBZ1qh46VmkyQ9JBA8m2Ls8pN50dAsO9Meozl
nVdIDwXJYHqnkoOKExaKKWRLiPng9uwbCYJexNPNiHPkykVi9Zf6jrREWPQRnqZOjsi2r6dpCH9H
YwIaLjA5TWVFUCmJ1sHDMavUJvVu9IiWxwMbJg0Mibscq/lVcU5gno9ejXpj1tppRfi1oXLvODIX
t2r77heKHjBtl/BVpdMEAylyEWpShBsK82AoX/b/v5mj1vIeD8pteg3Ah4fEoAXlxVU2Q7WP391C
csGPnoXeudVh7WzQmy/E+9M68fVpbpiB9zrUc8qJGYS4n7BxsSpaVMlxo391OiayZD3f7Umzsnfd
y48xArPOUPWl+ca7bJHzHnnzcfWGlisCUb/Kg4qXsUsfJXpAHghIZ+j9+NBYVsf1o4rlOavPE7Um
tO6JB/0aTmV2CbHCvjZ75F4u2x2hU7PQ7FrN9IrfNk6Ch7wTXXOj7Mfnvgek9PUxbKsow1/37za4
vhQdYUXdt7kvkLuHNPb544f5tNYTnEHF/bWjHdflnPUVB6trN/7ADBlKnHUOSpnZQ5bhtnRVMJkl
lxIyhL0I0240I707SHBjDlIElykZhxNTuUrdCKOQ66NYl3swM4wtLEGv4v5RN8TyyxXgRjKQXoqz
Cp7zLuLmWWjv2OajgLCh0jllSX5UTyv5G/jBZxJ3KB5lgoy3NWkycU1j0l9ullHL6LWvxXjt4RkP
FeSr460htDKWDOgsMlDjVy6pxraBYKYnNUTMh8mnKnv7DkaiEHMdJXSVH7qYox162Vf1XG5G+QJO
aNPuB4s3CJMfPtITDwKLcnhpXqQfYATGsm2LZBnsUBwG3vk85XRHM2e3yKG7r9Vy8+NHQA+1M4Q/
Agy8xjbQiKOmaMXXiINDV3OpBGVEg5GOJF1UMITe7W3vNwyqB6iEaF0nXa0LSDB65Y2KvEj53ts/
3QAJ6HB0iDUbx8NIcAKbGtUs7P0uYgx7ClIVwNJJNEjprgHeySv0D0I2Mb9iVqnTC32GzUIuS7Rm
dx1blTRadpFo/D4km1mBV9kkMXehOcdmZPFDloRKq2jI8vGidmcQVVDuEK1bZiU/TAzSerpoJcyl
oz5oe71JUuozhJ6wYyrBJPpUJUyXHn/fueox3YoMBX9doEhWBjsjm/c6ezoG5ThtKLkC5IFKPXGb
UIqhdwtackTnc4g2/bsbKYS62yXSGio62ImFOm6U5Dk0bp4XZQDtV0oe0ZmjBH728ZGXxipZPqk9
+0seAa3aaoMsjTDz4qjhmc5Y6yWxeGpdVcwIkAgGPqV1HsgUdzGpBtFLIrNpJ0hOp2FXMqw31V7U
n0En6Fh+GxCKMgFRlei/nVzqzorCIqKDH+7wTMcH7UW76H4sVPG2sAwB5SYrvA2QbzNavDIQc8dc
ueQCuanVkT5m9dl7yaBrF33qTmaIlfGSI/LJ3vbDnpPDRtpcnkFQsMzA4rZmyU1gKoMWf5RBhuzk
hPJkExDO0EkZc5dDyB71U6iden7PxJb4y3cBIYZ1OogVPUf/HPaTO473YfMs53b1iZBtuOjgaESI
rbHdUWMTwOm2l5J0Jd4XT7YA/gdw1ae9c5Lu0Yj8Mlg7j5n/JrKUiP16f0dzoACBonFwgco4QnXP
zwWJC/gE5ZxZfOLdC6TxCn8wsg2W2MnW4ZZ2eC5ylieZb2paF0ZBZP06YqDt2OA6xPcEvJECUsmg
F+tyd6LQ+h9B04RikSydLNitWID9HtnnidNZbYFTPMOXpe4hLUj4TZrAEu1Bx1LEnOYtKFLtu3cs
ZloW3ZM+LjQIFK6w5jtPmxH3WK30b8HiglK/WAV0SXDh/o+UIjE8OJ9w6fdD915unIHUpYwpzmBy
G5QWJ5r/Js1ck+xWZk+DfA+MnGjCA9Z3jxlkOPxevFnYDKWjgbdRViIqvT5/oDYhzNTKu0KDD+b+
R0Xbdc4Kl312FXomB1AWHlM8gauoxnptNxW/4m6CtcTHzO0z74XtQXl01ngxmnR7VxgD2xHTGiNl
IJY7/lMITzkxS2gxDy45lv/KNs249zbTOtcLxnpNUXJcSEEynpLKypnRA1c5DkBSaIq1pJx5QO4X
YmUHT87hcFxnXvmcHvVNSWa7qPd6yEoN3udIIEweg1D2boWOUWDbMczDgW1RNGftd2CAFK8yoLvR
u3nKrJTdXosabstC6LeTO9yfnpfRYmHIzcl7d77Yz2b0zeXzhdrfhrRaJGrUSztXD7uUsDoHy5AK
wXqqtdJeOjEtlXX33bV/w1eiLWBu/yAU+Ot3KtVh4MWsgT2hHn9DhJ4VFvzVit35ZQNnJpyP8hUU
8d8+mr0CN489+iyy6MKblmTQWalthwHpseJREulAFeFWtJkVlRZH1vFTGekFbJQdXyVX/IoVvie3
0ni8GU33zFebXyurix3/CtwzurlECfZivZSZJaCSl//8DLPjgt8EhA7Uv14UACS/0Puuj1rVk+tR
/ej3Wue7GV6NVOuJRYgPHfohZCx2ckQ6NL62b99SwJXYBqI05aD5B7+KIPKNft1Lsm5Wy3Ed0bkr
ksLvWspMpmjciHluUwIutlFkCPMLgiIzzEt/nZNT+EjjC1QuG2wiIqH8uZG945MmgZNdjqagjaM/
z9qkqcqelNDmioMLqcD01LitDshHO+gxOjywqOEGo1ggN8GAXwu++mXaXJiG0EmAZY4Wlw6tGJTt
wbcC+jao2PpjO161kFca5HyQCFlTTLGZbsejWHzpXgfswlEGTHs9EwO2G+MBdOz43CBOK2JFOPeZ
Ojr+sgNdXvnK2nYw7TYY32OBvjvPgtBFDRqIjnIMefH7d8NkhuPOzBXqoRdV80UNkNzvMoIQ8g7j
wjIua4Y1NFyPq57gA5VUi+/U+hJ89JsKZpqTa2Kgj+BA1FhqBA4gPwzpUf08hzM52E/FEgS9Bt+6
4o/fqcvUFg/OvUDIJ/RrpabvR8hY3ER487Mv4Vy7XK4p2vH4sES45bBj+S+0WyAwHSp4Q9PuVrrq
cvD7iKzges0KLCYAAegTyrHiODqZFkqrrCm4+ULdqYjy2W9ns3D/rXTvzUxi4c6KPnZ83xUsUYN3
LwsL/i2kjE/GHtoS1pFNF7LTMvctV60c5G+dhRPKfW5+nJ/AK0+ITdOlKUSGCCr/Gltex5pWg4g8
BVUG99gIibIT0h1NAqAUw3TDvw0VlRc5K0B4omPiQhjvEf5nBdX5remZ+kLA+7IaijcCh/EIXSuO
fSg2W0kjlQg+D+bxl47ay8ppDRAnPys42lOdICSmfXcVK94ummpt6hSSdL+WwWDPxb9RGHZtzxJl
qN+eGQ53WK76oJ6Z82Z68U/asNQi4qoIz9chM5jr+DjzHb8k941Ga3n6h69VLA5AOKywI8o63nXF
/B97Iecw+PtAZ+6hxHwDbMFF1auWnUAtc4WjM9VRRYBzJkqIqDpaaCfOijatzSbzdJCyLgG3jHTi
ITZmGg0KlmvAD2XHyzs8feovg882W/Q2EOZ8IARvC7ol32fhA8MIZUtlH0s3URCaXIfjtEotTD+k
iHtIkvnX+WDaI2cV+ZiSXg70rWXXj1XwqyvOO+1EvrrHV0TGI/QxO0Meue/Hs5ytzBHZZLKnUDS0
GVlRmrqb2LvCMwIXWkTW9s2dymz3b3cnTc4/fa1x+qFeKZsxJAqzUBV45TY70gqbXGrIicSd54Om
7XSabaJLCnVvvFY8Z9ueDu0xn7g30QDAHQ1n3NGwgTjiWVRPnpD53dkVTQH7jnBavgL1Fk50xmam
gH1pc2YBtZmb+6lU62lf75sFTsKOOMf9C4NnsJq89fik2pF+SziebRYuTOYOAAnre1N7N4yXvyzp
Nnz8+xKwNUtbBbRr3zhg6yjm4tdQFGvh3iXgQAp3mYzi4gDxMr/4EuaT+AhZ3pMpfT6qBEHBEJaS
QBGaXFbMkQKx/rEAzloapq3xLnLJzAXPght4e0ejztDDknLHjvelHZnB7QzBq9Y15UeH/f17goo8
m18xxqyx/uwkPJ+7wkZQGz9k7R/8egH881ZD7BK8Oh+CvYZXjMjl71ycRfyVDt2uhrTNW4EPUenm
HjOGXL/Jh3g5xt4d9MP7l1fkDV3FXzbwMUIQMOroMWDLJK7rgyP10tP4EtSUe0TNSZ9uecfqN7+T
s1KX2Eu90fOA3VoMXerHwTnurwHSqRArpPZ0JnbCyssAOdhUZwI3PaIbAIxLQzRnff6RHmuY8W2X
o8s67UlOPgrYE52nL4/nm/zbaMed+6VIVsrur52OtU8Db7mhXIJ5rIIUFDYDBGpX/P33TYiQXbx6
z5PbnU25/QioJDp+nlKanl7KEGEGc2BlPyDdefQ9NJf1+yPC3Rm3vx5Re5rHUVTtZHbE8a7AfhXB
ndMYaq/ktW/sCvFdF1wJqsWQx3QibB0UWLhQoDMwQ+57Od98fHllBQdRncnFKb1iiTXQUQkzcnm6
UlERShOQOwAXtBZB5O0XTfZjIzkDriv5BMFW+wwkCnZ/8VebWWvJtJl1PP9ppHkhkcU0HK3JKx43
l60JPu+VZSf2ndpZ9mEodXCOZreUjEPO7YoyQ5pCXKdHsu2P3gXlt9mcua7FiV9nzjpxEd8JB/eO
oFjpS5BGKdXW9HCgRqDVcCQ+pdAxPpHPwojhpNnnrxsuiymBhy5tZMZb7sXzWE9W/rzdENIVLPyL
zbs0eNrSBooRmJii7cW4Vy/xUiknuZvPEctuSspTsrMQxrfC53FFOh9yq6aTCXsFBiiIXkpHSCLc
AsEZUdwbpUM6lAa4pF4dskzoIUZwpZ2CIIIY3o/tQbqyjwAihj0AP45kgUU7Cf1xpAcyoWPhjNOh
ki/qyK90pXRns9vn+dlXDC461qTq127OryaGKXeBYoofzR/aDFSVNchsEqlBILv5uVaOojLH/JuB
n7ny51b3Ny3B4ZJ2OMJnQhxu/K2KcI4eCAq0ZD6AhidCvJToFHsXN8O+T237QIwhFHQ6kr17IVfX
byM5oS4L9fHUS8daLT4NNf+AcMdrvOIs81MMXcXiNv4Hj7Jp8mMpBk2xFxxLAc8Xbz4CfS9Jua5g
8JwixRJNHNmWxRcBgB2Uu1pchAOXO76BNKrSI2f/syQUsYSVzJkZTUQlWpu9czgi4u6DVlFULTYF
bab1PwJROhEtth2z/37G9z795YVORqrXdNp9hGMjVDB+CxEMSN8B/vwUb5zJXqsrpE9LPyLmHRd2
TArMteDRZbDN8AdFdj+9H4FjIuC5JjEWukGuWhMFwnUiCrIMD2xvmWiVQCnsFNNmEW+P1QfkDbj9
YBo476gcAtAMDeEXNwG9i/EgStqhHDMB2aPklQjscaJXrxCa/EhKJoirAKnr9mMYZ0wUYDWoS3dB
7JE8lbLE7CibED9v1OIkHpNgeevgYmCCmz4kL6U+VW4fLJWexZ261t1QVjISUjjFk1yoEtk2KQyW
zGnebG+jdB3TG3oze7toc2W4l6WacWtnY601RqL2oRwGXVNDOBSdrfSn4wpWE3n0sJb2uZmbWGdN
srQ8GqdFGwqtKbbeFgsFtRr5v38CtuLZ3SPOB8xfr7c9jSLQn7ZjtSXPL2w4x53F1ZUp8nDuHeLA
XCBVyiPZFptzdlhCKC0+gtU3LB1+ljj8A3mqOTNM/GhNpXjnQqjfY9EaKqcIEOZsy702eiEyvlwG
Ai6ycIggkrS7bpu0XWt3Xf6PPmHorWrLfi0WytU1arM19Ac9xbPSttjdd2yew/UG3Y1GNmHJoB9/
0P7OxVm2qpl32llR/01Kvh8KP72AnATrzk0QDhywb3Lg1pH5al9Wc+A3JQJ9HMONPQ4HgwMuGWSr
gxpIw8H9gmR+vew1NZ8Fi1apuUuzf4nLW1R8I8qmV2TsBqdDYh7+Vv+EAR1eC+m4kuuWztKSXEqG
KoKi3I8JzCC3TrctkViZrMKbIvIYmF6CS8myIVKXMM5mOJS3aopBf2Wp7QIwnxDfUvqcrbVwjGcD
P2hJQKJZI3bU0S2D0+UV8ytRxDASxfAgukWRoSztbxZlqOT7aOBpzeDemmwwXe88HwQCXEuSFFb4
AsFKUq0YqOn5VS5/d4rlxQD7hR4boE9gXVsxEnbKvMwsmQP31+E9atrG1bpBgXynSb+M5LdRNo80
5he82cVTbVm5UqbiHV6uV3j5Cj7e7UpGSJftIVmDg+3DqSJeVhDjlZ1mpTEz6kvIF4otzc2mcqbu
JLLkxIjqoYNQnXdIQF9FVCyMDwDfMgqMzbxphPngKt444mEJ+2qbvKTccpN409kKkm6MGiUcGWFD
1EEKCnVCHd17ZP9uPc2QXMcqwi7xOnnODpN7xfJa6KVLvhsebbXcp478GxpROR9HolG8tTjfOCtO
6gc0tHTahEsA9Wj785xuPbwOxDHGJ8/FTQvkWjYQXOfeTqklYMLd17SFComMVtjVDeYHOq9Rio3U
rQFhV0HP/f6+5J8We89NmER/pJdR1+fD4a3UNdYT81dLS21rkc4Z/+qjManJwnrIkjtcZ01+hXhp
csP2dkguYPQRc8jGFdd09CZ/u4uB/VKtHGYlL0i8v04cjNT7itZgvzLTsv+a43i8dMDqGZUtMQvL
NQYuXAlDZuKfbgyLmWgSl+7mc0WHELlK9+7OObPtHwoSs4/kZQz098iTyS7yZPVxGnfP9NbK2La8
pisjVLHTKP4UXaTmTNWNDKiqcIMS+BTz2Kw2Vuom8meqym99IcAlskgtxtk1a5GvHG6W0Ca+09mB
t+xUGCm4yvaqIGudJ4yZZHrFjkMg6CcHY9+AjW6d6NIZEtJ3oV1jBYOp5JY15aA1z/9v9zFte7Jg
ug+sYHVxFdJlSXUy4794owpo1LiTcJ+q0zUM6IqNofmCeU0lLnDqhOiaVTQm4iJ/4MQ/0r6f4ci+
GBvIRDvTDKH92bIN+D8g9itw+Fet6mDBWjUFRBipCDB1ySiFSiZSC4B/HyuDBMHU+tDrUtA9fBa5
D2s1rFeN3ZAh0BSaBWF07kgQTUJszvYqlOAmRB3BlZORxc2KLrK1C3xRI4mjSDVdKlOLkjQjK9/L
1lk84g7Fr2kIwdtJbrrs3ad8O1IrPQdtCkPyel7Ur175bINQOpEKd3Y1aK7qy79WNkKqNnOUnapL
5E5z0HpIqDsxgIKkWWF3ysXwsrw3kvUARh5y1UhOZms/OtAadQq790Z83lBLG/FPvtzgbnJbXLA6
j4/Sw9/PhGpoBRmMQ5x4HN6JyNVqxGxBzZuZNfMrV+M7uCmkzC7H0kl487WL6bpCYNuMcxsOQFtP
dKZEXou3RM+ISkI60v3RJEcQ5csICGmbsvvDP4x8m/pVaaTi6y/pmKTFrI4dfQBdvG4nNvONR3YC
YGj9XE+FUsFjJRBQMH/nOVXg4HGroLHTQK+UdmVI1INefGRud3EZQKGHQoWSCN0wJ+J3Iu1X7K40
2hkCN4Fo87noUinbmTNfgfozo1CIY3lCdinkgJNGG9nBVY+2eiBQXxm8F5ihHFWUI9dQx2kOqGcf
fEfY8qlc0zHYfw2uZoHZRp131x5NDGeoTY+OUgQnk5VXvxyOUO1nE9esoHdnR2tC+btTQTOSS9X6
O1tPK9g6AdAiemfurSHLNPQCmfw1CE6NP3+3Lmbgi2NDTv6INZSQisMZoO/M2NDvqFhs3E/+nQQc
LcS0uRc2kWJA1YkJSzbXSNDvKf1aR1Yn7+kEdWeUguQeQSsJ4epcITunl11SrEb+jfgMvWBLkr9e
4CaHX8+i7c3aPVo6OcUc0RqgM4NfFLX9lqVM17uPHkZARB2tryq4mjWyn7yeHxkDapUfrGuUosw4
0RspEpBaeEDx0Cam3oZdRlOPuql2fuBKSSa26v7MnPVXZ4snVIM6Onqj3macdajzfIJEcG0w4nUJ
OqaQea1Z+WY2cgRqDCCJ4P4e3r19A05k1W2DVmp8Fa37IXz08qi0vN/Jxbz9Mtuw3qS8TkakM+lh
S+/PkFuH7CDMAC+BVEQv3IFoTCTdxS8z0+f5m6mPAqJnQv0X5c7tzcfPUNkRs9P+nzjz8Auv1LSF
gaY4RjY2++HnQm/l4we91/UwKQk/K62SQuJlubE++RRuwv5cRVl21GSZaC0HspMXm6aGBzbiGZWR
+bqvuTAbTfmpX83I0Sj+rdQsGejgv2igYTsw+oedPArkuoVCv7sELoA9qd02zuPxoFl8g3P0BBM7
5F3a72uVRgNL7UIH+5orPRB5OOy2o3yugNdjWeH2MrvA5eWe6upEfmP97BJOyN+Ad3jYCulT+/OE
4bA+Qn/Er6dgmROo9m9vX1oTGtuAsN84WinZcw0Q3O7K7poCU/ciSkbWIv5RMwNpnS85hUZScC2I
UkCsb1vh04yZkbWrVADRc6LWhblxR5M4PVEpl1E37D8nYL67aftaRzVksfusShZF6tKvWzXp29ml
8xCPlIjvFE+jiPC1KUgZPmTfg8dLmpFGagbQ0eFGCrjpABN666T7O32Nznrbz1/wRAPQWbfs+Jh7
6JeuLwd6NY5QwOyPgYzHc2WVorpRNzhVdjXrHzLzO7nCBI7L77sbuT+CVyKlnf0BgE4rskzIiKfI
DDZ0ez5x50LWF02Y1aUwYZhPhqElyy12hQ+rsmNkCDlzthkJAaO996VhDkiZvj2lCIGtBXrFwIhD
RZzLfmlbanXxR89d6wYAoZE9h/8YPzKqmVVczOv+Xl8Com+gwtLP/c1Lmp52IHhlXryNP3v03VU4
i5XncpafSnJKkIwRDsdvtsCmWPNCkuML1YkTpQO6CEGRmo576uvKyMZRXxHG2ZILqZKc3W4F/+m+
4YQb0KfAxZcye1/GSG4lLa9ePBk6DayV1nHK5eNIJd3/pjJxzv8FfQL5Bd+HuPs3sktJiyhCVq3v
jht0FBfuo9zRgr3RLNtuj6c6h0VW2I8RAg7Wg9mKYZQKZH+t6f9ao2gaRy0g/aWIfUI9dC4IgeNl
EBWm6DvVxtPNIOqIV6jjk8fBFykZTH5V8ie7Xy6q1Ap670KFVwW+nQ7KhizMt2xaXXmxJWDggStD
bkZnXX4S3CTNUa4oMd4dbyMJmhE3kRnANphkx8DVQnCHQ8ARIEVB1C+puSgOcFqiJt3T19gFYDUh
DxFn4JD36S7q+4vsMLOon+rSkbCbCK4FipU0goyygwScjVeudOiA7suWOoBF/ykBULYzD400s3mr
A8l494gzN3ojiJZ6lBT86Ug5J+7GJT0Dp69JyrtmfdD/Fnd0VHoEP/t1JSelKqCXWNB9NPAGqlIw
hxYAuJtmqvP+30lSIvKlqU0JqMRDP2vGcrp7Ys3j1/zX5yTdmjtoKrjw4R2Bgi9ffUxl3XataIwr
/SBYX3BzoQxIm/dC6kZBsMn89tevJ1lCtd552RX8OwZZ5SeCCEhllNV4vTkUZ+ow4TewPDhNnz5d
x+6QvIH4wrYrVi0LCz/jQr89uNnN8x72qq0OPs1UPm8uLZxWRivqGYtEWG4yS2NgF6nQMH40mTPv
GkzuVKMFlr7XSRWjQ1T7+1xx1L25fWmwwRDXQWbVqaixPUr0Rr03OJ4AXwJ9lUwyfvPtVTMYfNvk
j50X1EFw10L2mF2uwpV0VIgnAy5z992MCxpEYjolf4WeBobAFzIk3ri5mmwcdXyk/PQ5QrYlNTVn
3MydMgyln4wW+FKL2l3mSugo8UTINFLg+4WNT6HN12hEd4AdPxlhOqKcQRkz55m3HZC17VBQTrS2
qLwdy9bOA+bMuTPpUhU06oDhjne7Jpkyay2kt+nFfGxvLENYZcLFHMiN/Tal6R4dYRSQ+e+t7i/N
xnaqW/pjB4hynVBId5S5G2IzmRY/a9v9EwAUHKbRfXgKGosEYeGUAftErfSCjYXFgNkyLKfM1JxQ
LzE+OBWsxAso/vrxs1rqGd9KakXxyp1JjGZeinkupMPV5KTDt9Y+O/UdXyKg3VwjxKy6f/+ZyzWO
nLq0iqo+T/Y+HlEsnWSNpUUK9LKCv7v2R0dm2b/SK5UYI2iKKJ1iRPYj06RzOaxzjtdPz7gno8sM
btbJLSHnLG/O5nWkORlHzotoKb7SOX6SeFL/Q7BmfvEJvTw3UXwt6eNq1GeuzSY5LXDatV3MIIaU
gTzAJ0YAV3qXvDhmFfwwslsbOUbyc8jdVVTFfUidcvFIANMnvyTPPpSn8HLNY5egmwGZ7dKkexdO
0o9b3pOH3aIhf9ej62dcLODOH/Zd2hYFPB3eoj1wpWWvBoNndzxLE/ZS8tWmuQCbZPfyzY3UVcCx
PVbiaks7QGI//AWonKr8qY/SXpSd2bEWBmQ7bMk/9TxiA30+mKRkn3yNAnezZwbfnE2RsEpked2v
ybY94usTS7c5Pe4ElTXZFEoL4a81NK6QMaVQ8qFCl8ztk+sz6xE9uxHn8tmRQTn5gnRnZFzk/GQ+
MCtRxoN/aEA/QmAAs3An/gEEVYW7LgZEbr3bbANhlm+366Y0hoc8ixuH6btiA203AFAabWvsCeXp
5EIfLQGitKDDimrMSrHczLVPHrHETOz4C3MZbygLGx506vYfY9QxoHqaVTyY0hiC3MOJQTt+39SB
PArOrSmE6hIsOgTJJwOKVykQwejJrr29gH+QZ/f6JjcmYIfhHmcS0vvy1aGd7BkmYSXPaBxNEVO1
kTt59dh4NoF3X9UH+xdVOQFGk0LijeCL0CFqpDy8l6DjKChJdFacoLVzcpeR624dtEpwkoHiCn6w
7jJsHMru+HGrck+0olkLoFrkWjhb+4RTPejFMutY44YR2AjLEF8z/xgUnfjWTo3PVjT4pAZBX1A3
cujK9SHR0qxTkXLaxTX/XiUVT+o6MRm/hD5732LnPbEZRl2K7lCLBZiaNf7aY2YlmtVn0FOdSRMp
ZBnE6E8IRKj4dflEwWZ/y63f0ZsE8oLPyeP5OCAbo5cs6U8Y47zFp6bW9jihFcNLxf05sStJgr9v
Qg+xaEVW/UewQ3xpeHqT1DbT7mulmcovEVydzE2drQQNEo1ev2GjoIcJ5gM0cgb4EsHfBnj5RyJJ
TyK9XYs0ACTZgzjQ3fnEkUrdI6dHlO8pXVt6wFHxXhiAc+IKITkpHj95y2emyJtcnzuwT0JFzcLk
rmblsmLTlOUiyaYsABYiT+mHzftCO7kwzFSPz+ZSVDOjYPETmcwx4jVnEMKwdQ1uak5sY0FMCoqi
f37l/Xq3l+rS9GHlXZ1OCudYxqmPOPOysXht678mJ4LhXoa7eqMaB8gkOSwAHYYTO8j+K301h90M
bF42+kNnTojKEo4W+hC6QL56sMVcpEKGnYqrFVMMZwqVOa7NFkEBCMw/lZ3kTO3Wjd82u66tPO/W
yXFHO9ttN4Qd3QhxiTO8BRjb6nTnl7MSVYeC8tWWospeWNovOkaNPzqY3eL7TkV/QCWPfZjuNKdk
dta9467yPRZLH5w4x9XlbNarFoai0vIcCdnZIy5b+ZLNE0vFqC7AFvbJ8snPPPtrW7E6Q6dyo7JM
uXd4yyRikeQap8pbIWgL1PwQoH06ph5uetISxiGh1mJLTb+pMN9p1bl9ToJfeVfrGNz4q/evsL1c
cEMVQxnIncxePv3/XLXEZbC1TNe7/s/MYz72892j86QIlx06eZZXhTyXUyvPjpWZ6mPMRoTe6g0d
hgO/DVBreNx5U4Bpxc04RomN8CEaXIsUtSW3b3U/nH13vPPpdtHau1lsy9JkyD8O07V39CsmetH7
9FGRAITxo9hQe5oiOCCOmcfaCofdbiegfzb8Qf+wpD/85vdZEZgAAlo/cDgem+Pa1JvsSV8pZtT6
XxtmILVt0fDRcMTA3GKcwNuHbEx1EIY9vx7d6y6KR1Pi4HBDlmda7mIYjpxEKF2Fy5DEoESDeYLL
wNcY322hiQ27knC28/08CiKpSWP8RSnDGmvQLjIbjFNMCQlhFNeqefSQeR3kCRnMz8IVgzxyS8cl
dj6XDDVe0ls8XQK86HslXoh6nXAqvrFtORLcpBXxPi1mX9j+j6xD+AKRQFMc9zIUj6YLNjuChibc
DH7EhUq7xWnQtDKUMMUqEKLZuIMUpfdNQ0Gz6JDvGycLUtbtUhgtgX0sdzSBgPAFnffQRZTOim29
DYWuoq5+zGrdZYs+nMLY+9JPcFiVlhQvpHXhX2XKf+uRGF0yRDyNvunT9YmiiAF+oB2nFedyBeP3
wXXShh6rBFBSC3Byj/9a2jsMxRluD4LDXjEse8E3WGCyEB/tW9hKSLYw4LJhDq8tgLvUWbrHhXkS
MgrJLqC9edGzJwlib3HkBIutfcsWOEi1TyD1ou+xPmUMrGJMWznTjwBg4GPjCuLeBJi6No6f2Tv/
e2RahWb8KLbyhxsNp1ddv3Ovg5btJ/VgmMCNsqmaOzgM+4pcVqhJyx2D12QWsEVyILulWnqA88nt
WtdepkqltfWVTzulYPDqqc2sUQt+GR7Cs6tRMVvdQL89DA3uLhaWO+MY6Zxe9JMO8DrF9lLbX6yo
p5abpEjrtrCJkcLZPGcPffQxooqeVEdXdLKkqzv1bnCq25AB7s4yuVWrhOowoSTNYSKRJUk8+i4C
GvExI2JupbCZi+p/DP+w1empzULJOJKxS/dQV2+UroQgH/aSWJ0xX2OgRSwkB9oDyjIESwf1G+xq
SXHtj0RWiZLSivLwSgFNCQDpRdHRNN0zBcEq1ZgoS3bfAz0548wCYdMPgUB9zX4dAoQDeLnRg4Yy
C0fwrnWzo/oT0m1NNlB2o5MEeYIZ7iIR91tT8kp5Kjea9XxHkP3xlssE9DYY47DtWjor4fdGiNXE
KFMFefsNR3p4fdl25PF9uVn60jbxw83YUBiZnRs5PPMKX3/9AA1O+y+BXG37ivgKlX2ZN9h21Wkx
qVHBKCf/EH20A2JmLyMHRNGGhePBDC+aituHDxGf0wvKEG7dl8sHW9FMYupvs67WbO31VUZEcFEj
2Xpxti7GR5sb9cVLCU6h8OL/FDmokLuaVRJUFmJx9MfTfXAMdgqsjvoWzjoJzBzDUO/ykvv8hNfk
T9FfZYdJeTDzDMLLt49VTqtbwEzipGEJxnpyZSuCavvtRxA0T54X53ffgynwGwCo+nqg6pLVk4CY
Fx7uVtHfAogurUJ/smAHrlCHjP6gkbavtSFfBKREWv8qq35VdItlYI1ga7ND/nMWIKt+MUJDClEx
TWw/pNP1EV0pGp0fD/KfZWOAvVbOfNgQ1MCqIxWvSaqZPpao+bClBpRnBZ2rqh4KcZFBwU/mZh5I
xEXGBx82vA4mBqNCAzJqmErkAqiWe2sh7zQQiCQZTtpgvdXIyUvcd8WVe2Q33LoBLPzy+Uk6I4DN
+q8CCIqHsz0ACnchaQXQh46Y7eE1GBgQX6/agVJXEU+wmdElhp+BEZniWLdMWGLln6NGohlFUntT
03WvZp/21dZJSysja3WO6y4o4ku1vrkh4KPCi+IV6d+UFrctdQVKEQBTRiBeJrNTjdkAUVcTU8Ns
RoEWQbFm8GWoIm8wq0Nc8/RN9PksMEDJOiEjLU6+9sWGXvwSTxbLEpVgOLQj53TOKLHoblozuRUV
JKPkVm9eq725ike7L3tOzqoJHk8Fs5ZMaPG2gqy5oBjut7ZYVtI0IQ6rOIAazblMwVhmw72Q8oR/
G8f7+8R8CzMyApq0ftYrg/QwbOoDpGJkhQo89pMGGDzbUhYP8VPiOXU8pffx1omi2MB0HxLIC767
rsLYIkDa8guoXUvHkzp62RInUc7tLLOSV5GeTj+Mx+OhgsWUeHEU0PMcCOpz0iPOAbnfn3WI3hMR
YnBnifLPnHScnyDMg5SfImgSuQOkASPCd9/l2CAXAIa7ufN9YvtOBVzFutFSmiiD0+bY6ML9AsU7
qaRKVFYTnPupVci2rx2snt9Rwna6gSzPwPGUcnaJiE38HfjDFJhzfPmhOWfIqrI/L5Jl+ZOg3P09
jzH0I8Gs9ldrxi7Sjo/zZrypwzfMnMQ/9u3m2hB7IY1D5fo28NDC8HTkqy34CZKbIGi5f2BHpDPq
CkMXL/fz5PxMubELePPSJz3WmE7dEKYdk9S3eKEkiMJoEK7ImENA/CdT5trgB/HXMnPFBbwy9Nvx
xAgbovl+kqUKWNh95JcJIofNewjAIpLpnkH4Pcl8DQgppjnawIBxGvmMmWPQYVZcnYYggpDMqs+X
BtwVHvmwNDrg0ov50XX4HAT5e6Bap+tzDVolgdCuYm+CHIqaCitZE4lKVmIU8mpYXxTcQQFfQIt1
BdJWTuRgyhaoaqosMeBWeha/wo5aQWE+PWafD4qpPqDv4XPPDoruiR5OcFSAQtGRuoxZpTPf1GQf
QRaGfPSdogOMFFMba7ECcjP0jUVO0K4y5qrgV+7goGRQ4r7tP00h5AAony9N/2GMcpI3FG++ThQ0
UPHgtTV8K9F+4Quh0TNpTQDxucCzh4ktRYl9gAWrm2XgQeEoo4MWqxsOsND/DVFt8Nknj3KZ3kG7
PSzZWGYgfjFrCv7uFESb7bhe3biN1GMSR2bZnfVqNx4ubqjwFPNYJ4cnBtmkdumxwSYwCilUv+Kj
x7pbAtvnaKesnScrrG1ZgftbrMEtjI0mw/BmW43fblZ9JXgAKOsHs2hDAMFP3qTkBCp+jDMKLKCh
yUvCGmF1VkNj/ONUMNDt3MyKYubV1Io/5kj+3+A3IOzqQ44JQtRiL2Wj1ptNbvJDbT2/UTVPdK4S
Wor4lO4BrmBLgBbsi5thbBfNZlxsSznUpl610OFOLu/T+kNquCI5sgN2mJJ6Xt4PxWxeQovAKnoM
fsKuuGxFZhWX5eQb9p3MJ1RAhq/ByUwlNlytAp/4UO8OIUVDViE27lyEprFAqufjsrShlUjevOE4
RK1FI7x2xjByD92P1iuJDhzmla3pOkMWE9E4THm292+kxZeeHgxy5RHRAByEa+wDtIy5+T8rSo6H
Z+b09W/L9IPIiUlyPfRxhZjdrFmp4wiQJkWW91OW88KPUp0KyKGpfsr9nmx0/wCzkDTm8Vhf/vFV
4vzbgUkQbGrznuOwupQgExOA1Bp2JCQtjrHTJIdDWADDBIfA82X8xREnF2SVkAP8HsgjEZPCVrqm
zVbTRPCU51XZKY/9PvXtscJkUAyvptdM6emRIGyMQvw4bQryDBmMlsh5cL1KLouBKIwL7nlG5OuN
aG7hK/+ku1itoQhhleJtXgiDTHKGXf3wXNnSRn/xNgeqP9uitNxdlbxol+orym4Ma8ppvtVbY0GM
8hM/Clkpy7pkB2ieJHwTARmCCM62Q6gHvNBiP54gv/nhXOhRXsGqCwruxLkJwzpZuqBcLJk9VXlg
ER3BZWBAN4pYX9mVc9G0Y3L2MwIF4K9G6XJF5j4Us5LOaOUCgWbW0OLu3tTceXkpai2oiEpZN+iV
na92EDCANIDvAIHDkX1VaPdZRQQcH72akGj6io8XiVf/PuKM0z7DF02fuxE0wIkT2PybTuhPY8TU
oEOEZXYxvlEFOAEyJhfEMi4Hn43NdMpTTEhq+cNpwTHkJLmt15jElxzEZXbqIMufbpim+Wh1bp6E
3DGBE37X/NtHJV5SmXCJoIUEmWYLWeZ776yW6IWXgghz8Bd8ilL5CPUZNMGpsHWM74GmLRu1B+OU
TnO8CNuFcMW83cFg/IEvPbI0s9n7gba8JEfyjLorUvQfxbPWJEuj9vORRn0Uwhqn/TltHFH11/8g
3AeDCqMAGQ1KkxEFICgGkhtmUGaVnr3DK8shznRxB8CNpWCMyZuAGdkkOp75BINO9HqDPE8iZhsV
pUwlCYQD+ebpwH1G8gopEtn9AklXCm/arllVLJEDADGhPZ1YrsLB53SDqVBse6r67dHXzSHvJ27m
OJp4+oyeP2/mJtV2LD+SlZUgmLcD9Q36XphmmiPelCIxYKyqoxSCpPWfHnkGbhuvgD2z36E+va+T
onlv9nsiOJd4GSMEhD9NZfizSSSl35w4hoQtuX1W4aJMBe4IAnCH7i5F4YBGG0uIXBSveIY2BaVN
ikNMCet0ZisGNIZX4mHh9PeVifwGFfRUJvPSp2CPdOgNEZzCC9reMO/RepnYn1K4eIAkti7WpEJS
9cdpguRFk2uLX2kNO1iR6anxHWci/bsO9VLtMYxmA7aRJggDnbjhSaFUOMsUgVWzD1KQay1Mhbd2
z9Fh9l5GFeOze84Amiy8uD9tkeTduh2wa+t4wGNHDSUAfc3ZfLoK/lUlp5bwZFd51dsUah+vKYpL
8T2+wJW2dkzDGcN0BVcQpV066JYVZvfFE0HFiyiAevh5E3HuwJLWl8m50cdon7btbD5tqjP00hVN
auImeYh/baJg6EHhWKmVS4bkQ7qn+IG4ktJc7ylDMPlJqWyJwRmY13SQCPPXS3EqheW2AkgoWaX4
TAdeEluB0KLX0tHJbF+2v0eirCXSRAWqze3CPltF5pmvSO1uvl9b09rykpqWYa+0j6h+0Tac+CSN
fEpoejjHBiuMj1WiaRUEYl9Qn/LFiZfFAYJphyWgbmbdTwZwus3fpUmO7MebO4wy3RldXECeufjt
xYMNLPj8jGbXbdaBnkzEs482HoCNRZ24goa/di4RR87oy+P0ZGVA8DxDck7RoW0cnEI38bEGkCwp
OUVj0A1tkEX/ji+w5aEzBUcIxts0n6GL2S7apuf3uDzb6XQuGUhYUU1086L4jjLXFPXCv4aeXGS/
0r/eSIRcJ2e+DHdbDc/svJWNesd45lYFVYNfGhs0nHmOngDDS04Zx/Q0/nYuoUYrnasmvGsJC7DS
W190i04sNz1afwL7WiuIfPnX45+sSKas0dPt6lpStZ3IlBGiaf9D13UYTIrOx5UL7bmaeXyaC3tM
bMLQwZvAZtsVoJc/HlemCE9zZJOGewfSfzM6WmfWO3847mglOh/+E48EUgomdKH5skEpbUtUQMAV
S4nMxhA8y9L/aVDw9u6lqnDjO5cBLIWHKhZ5DAbVbeKjegBMhbwMFx4OSviX736jNwsAFznwRQ4G
Ymzv4qpeIPBjb9jUCTIYWnhOAXJJwBAZYTcWULgfnW45YsmrsSd8EOkrH93G62ZCA5+IW7jYHHf8
idcnOa11gSRSlkdoMPgSZJUJo2cNx+TY6GVo+cLGU+ci9+TVlKQV8uJJzqT2YB57dQQ8qKGTDkLi
Wns15vFwnfXDoE8cvssT7CLWItL9xmz2SQQZdw4pyj51f6kkL/jK0lCWqmwaeJdwi3BeVASXzfag
6KXUYdIvMAtjxkAlYy6uo2DQn7rMyvVumIkRgRquK5O8u/2AHVR0zzZovh4OARo76/o6YqUMa/qc
PnZ6RyLCzCqz9ALhMw9b3G0Dmx8dGCRr+NzLS+cbu12Wv7ej75ak2wTabFbZ+JCuTe2POxeyrfSD
Q9/4ig8JEvcoPU1hXLHUqgZrIlQBa1G1B/O+R+MZ23xdIrfWB84t6FL5REu/Lhz0kTxFvyTjaMot
Lq/NTST254IjCZaTcRiUrfK9BUR7SYxRwOV6dPWU9v0oYB+3OqIMYoyEiSC2ABzoqnLidjnoNjT3
qUujRx1BQqoQNIaYR85Vg7F1wsLRZ32/dyM0HfuIM/bY4qca2Q2qJTzrZodscU6pN1rfasJB7NXE
z+gPBYZs+QDFRm10JqHmafS28GUFJfWYk8CHwMOMfKG6Q9g8IKww2qJyvP0Qw77sW5V+it5Mnti9
LK17j2yM8zKhJN36oe+g7EmgqbSFy2461xBvPJBHNSq9lQFAvgMrksDXT2AYDJ/13N/ov6ivcmWa
P9jprHl1ezZ4OwkRnIP6mWRmeClSNHgYeCWG1pftU4Px/ugG4Yecb51b9u+fP1V8tE9iaDT2tAJ/
BVpf1vX3zydUPduEPWQ8Ipd2F+oE4ZYYWkex1AQuStjq6asTlmTW0qmwpFXpHRVMJvJ46gbVo1rr
Xsnpb20vdHdHERE9t/ysD3HKqA/PKIB3Vshp08Kz77H/rE8ICROlUVNCpZu9gu3xLTVy3jck/Nf+
/LhN2d2/Dyrhp/EqAqviF5b3ayO0AxyoXO/3fSO72WV5Ik+uodb/Kdhpe7na1IUGEhd8rA1RW5eM
NBiqNeypYQ4SMshLnVN+mF+H6S4PBelqlqBs4TdZ5k1j0Ityl3hETuXn82ugRdxXoynNqYIMVNbi
4yLCUXVVEEUUd9pPgv2ZAdjh5ZwWMJgPnBnqzVA+M13TkWl0nj2YkfbLuqHbltjFlWPz3GkTB1Ev
446cVBaqcqKNqxlvTG9xTiIvBjR8LZG4bxruGYbNDB8yK+AMOAe2f8xSd+IywxH1g7r3iMIQDyVL
pRXIurM95D8Bwpt4XF/zInCCzctiyRSiKaGIWOOtUwdngU6Y53eUappwVUqGJaYYFFaYTMj1fxUM
zSFvK8/3Kcfz6lUv+qkrmuo7o924pvTJqtH17QS03FFuKnkzXEZN7BUlRNl7rMWXC/wQLEmdM3Ve
pj2wOdg5bDcc1lF+cXi1a3XXJflzXP2sQtg6zn65TVWSfIKbjC91xGofxY5xpJle+77QP1VVW8Py
zOGLIu61f/nWq7bn/gBCQ1mZw7Eno53gbTBjL/A/CC3JW9mzSDgkjvOBuENoiHBtDQp0I65uvoAj
vBDki+mzTlI90/1eEcNx9PCsaB0JhjeJQdf64p8SmfU4pa9f14VXDqLNTOKAISEBYWzjAjFnj3Xe
c0cJfF12rZvgqijd/XPVOA5kdmwXF0zJYIcOmP+m5agiHfVhz2gruAV0vywka3lA5ZK2UksxqQ3v
KEVIF3U2Cj8vgo38cHCo0rSG4oKztp5vqv7hajWbqe5tlXfqmnf1QTaTP0THubpFVwWLcLAL6DKd
zS/zrEV+0uR4k8zZi7pmAaJ8Fj+xK1KMaQQIvEx8TO87DhJ39DLS1B6Su5YV3Ps9WXA0kAqN41+2
HLPIVq7ED2h0bTaUSjnujN0WsvI0aJ/hgcCyk3YAkia1SCrZX/8ZBKvhj58PxXUvKbb0SDjttbEm
F4oXFnyIrNCIM44zgjo8cLQFKs2K7sdl/Pu41RNwqqBGBWrbzmplX8kO8s2irRnIN64d3N80Mfi/
I2s8aKv6VA5OtgtA6koS71RvxLS5ReGWC0NpmH3a6uG0Ea44oTzM6xfV6zzUhyS/S/P7lU9wTRP2
uR21EK7PGC7t1bn1VrmcDxPR5NKjXR1sEu8DzWBSsoC7BCcPGc44gXilEH/XJ3qRBbxjkATJyu1p
gCeGPelHQcQal6ok0/NGWMIJoXJEAprVsQUrbR5BQfLmS6h7SNWlEoxx5TaDTw/26rkEvPYzMxMK
Z3xhrQr2ed1cpSbcVQg1cAgiVzYs3omyIKryMXgmrG9rOCpdWw9KbIyHuw6QBejkD3MY4GZQ5THU
raBMTQbbeW+BKOcDI3II97+DXdn6QSLXsrt8Q6wyK35YjlDpzV/mn2yvYzhXoEW3SatauIUTDVwH
GJxPzlVFcel2edvpyjlWbE9lsJUsNF8d7P7uCKJmWonFbwLHRMzuECe/Oco2QxiMD0IcBXYHDajE
HfG8qKKO+WPJcEVREyngnEIKglBIY/mk6OtQmtXe2PwPozpugqQifJavBybQ1pX90lp2zWFjbiE6
H7B1Vb+Wqv0yO8POLzLA0H4usAmaED76uIRIKAWu2scWH45I9wrYBHahpFIFK6217LzvGnv+8Inw
9EfdzSXaLASub4b+FAaeGOMEkzlRiTXaqGcgBWeu2pyw0hI1JGQ95htjEWeCZ+Mjl+glSWUkr8Pl
EO5Wa88koAYsgxsuGNDFb1G4AwUkm2glhAtbQvYdsmIz4IaPJgzITLgLy/NT6wiESqKjBk1oinvS
oMp3ZDMt6wfk2RSpyFel8VC4iAgNlx+JLxTOj7XtClx5u8YHuLnnrMRBWtSN0A6ZnB744lJkw7jf
VCxHYN3qp9W4HDN3Pq4m7H86GkoCwr3T3SKDqyz/bAOvd4HjKMMMo0jbmaJzvHGRcfVlR5cClTet
R54Sg4gA0ZDlDCxWtOoenk6v8psmOdp2GoFV/zIUqF4PvFosaFdWBI3pjCdg1OJbvza5bIcwm/tv
BsmGIi/Ot7pFf9yrmjCfHctwGW1pxsIcCMn2E9vP5FC/i4X75qqLpdF3Kd1Ui6M28wXzIbT4Hcct
PSiCElslqW3nO/3DwAA05pLFQ/CAuB4tAeBS6dU2DOt5XLrSemzImJwaSYgsTpt8TbH0CwesXvSd
LDhA67EBUUUhvfFZM2DqPyo0x4BCW6FzexBR0CjTpWRtDYrg5oR/0D70zcQCRk6aTMDEvxByAB73
VY90/ppFFTrGmOUFLjn2ACIfcR/kDph4WMq5jDVSrXop0fTN3WY6j4kQBI1DhVdA573ew+6rmLG6
TAegpB7FLuT6CENAeYaNK1m13MF+/Y4qDIGKkSjZpGUHqP8ppcIBteUsAErXBlLwnxFYHLduX8IX
9Okyut+66MHuxEocaa/gR/01nQjdB5CWu7YprQXLLr/UqawmjBHXttjE1ko/UNgGl2n0uiVVZCZZ
W8pm4JRntZoHMDiWsIz9GtUYCtJuw59zsYDo/sKV1EOhUdwNscVyXkNBlx638Y2RjwXqOARDGj6Y
i6CzlB3VsX84KWng8CWSNMnNoqTUcNTtbZCj8yx65L6mfz41Cqyr274znLZYxCFXxT3t4fYp1jvV
afsvJSlA4deUV3/I1qbnTkPgOqgzoVhechHoA0Jk3YgwbmkVSVKME/zy31Ljir0iM2D3mUz1V57a
Y5fjzYoe+nBIBrMKH9PPBwzq1d2XqzzWql1fjj14EgGivGRAw+HKFatMTOcruYai/TpWj6cfPmVw
X1vdqXTDDI1Tg2YRxr9LW67y6tNuVtr4raytzKKQ//ubG6Tmki1SshrPgUrmme7I5TCeVHlDnZ4q
uD4dZRuG/xMiLqHGC3shMCf1sHKl3UYVeqFTufcnYHVQMxvlJ6pS07lIPZPKO9QNCP5gV304FIg1
RKcVs3MaRDZ5eFjy3A0/iqXl2rDBhGnCPt25BPhl+BZNltLGoyKWPnlS0JGZWgSWP+x9WBMixULF
nttpbaojK7/GoSE4NdEzU54L7nKMRSEOhM3yL1f2J2lFUFA5c82IpHFi8EfH40/BS5lHHJP2zC8k
dRvpAboWJ7qvBDWI1nZMApduAN19w8ZYuchRL3QhESvRal+T7lHdrRBIr8B5xtOjkVSCGkuFXT13
VPMGT7ykDZc39g73cR3VgOnT6rErLymcUm4GUDDoQ/yIOYTRT0gCPdXfM2qcIaTSeY+lVHy18YT3
Nw2k6uvQiAxiivnGczECEE9xM7cK+zY8lokSYLrOgrbj8wfptgBH3xFZU1s5iJTJdSNJUn4mbV8J
ewsMjfNXNA/6YLBKyGDQWF42LPYj3hMxZaQV75gPyoU+uqGq9Mnb59pZcNo408MaqKkd4C+uBtgo
q6m2YTkEgbaUL9qmwFbGmf/U5zwxqdrNcEDbo0Ag8qTcIMtivj9VTqLCuOemJZAN85pW0vpeH5AN
jgUSenu/LFaRFvb+nemiw0eNqCWVzhhDrwa6oZu1b3YKxUIT1PYDwtB6hj8TnXiznpWNY/qnZbPh
KxLpDPO1Z4VsDFt0+ZDxTJvfrmv3vOH+CI5IB+93PEPCxrORhD7zHfCn/xhjuFb19WDR76uR7xF/
7QXTpNSbUBeLbR+uAf45CKmaM0mAM1i7x/DyTMpVL1NgszfIeeJfguBMLCP9vIY1no5dfz/UgXXc
1lqz8G8+yhVsn5VvBVh6g0hWmnE+hFmankowXc4XSnK01MrkyBwd+V0zQn89uJlQoe6cLUkr7S1y
25JVtf/kS0GNh6dvslmbGsOtoOjsu9yC2tHPB1HeprwytzRyMFqaF5eJVEQbN9JN74GyrF0f7ih7
mcYdBHVjmZK+fe4bxl/vuG8UvN/3DGmM0qgbJZ7VBrA7ASPuHaX/IrllI0dJoQ0NkORtX0dwQz/C
vlm7gBPNDQPCGOdwb3fwS0f8b2bsLooVHnwFBZrZFQsqWoJDSg3vPdf8s7/TvBXBNV5F/sp9duDu
46sw0fVUDh2otv7cAjakV9po48dEpJiw9qDJLbfPeDOUn7+KbuC6BgeC4kZ0fr+mAAd9ethImac7
dVgj4sjmGPe+Era0XtUlcmqoMTaS2jnX0YL0pkqLF9fjYb1n2HYxWJ+iabbVJf21Kfh5UZ34VLiG
m8skX4b7DnaW1Nl3ZBv2tdZ1kRssefvYFFJRg9aFeUvokSizVcZeZz1aBjERfQs3ocpqihrOLOsy
Kt/63oYiT6+Q10YQsjRRCMuQpJuxACIqMBwKy7WJz4lf64C1GmQcMYnCC7VlgF9MQbV0YSaYXPFp
CHAU665G/hGp4HaXdvHPN1BL+mnbNpCdor4fplPEY8Zlk+oh+ZiqEd6mz44wJLpnvZDS8ozdj+3+
Yvp/Yfaq8ThI7oKQHY/y3ngBGfTzcJLPLb1yriC/ejPWb8be0Qxh3zbnuAe4ObDIz3cr4uvq/7ts
Fj6cgObgf+qjGZcZyUiRU9u9vAU0HZc0oOFnnBucmJjBueffw4YgFzbKEQKGxTqpw7iRdb0u4Yur
tAt+h72PTqDwTDtHQHHzdyGEjX5z3tvOoXsNpWi4EdoNkKSpsBI32khUgfaJRrbHwxTMeJA0vk+t
RxI2eXIrIwdDvfaTfboKarDv0kVPcz1Ifvudigs3VfU630+AimsCRxLfUersswcN4XbXiEWRn5x0
y68ezi2QMHXsm06kFHqHtFbNpGxUV64JJsbZk3XBIZCycwOIy0dmFdb3P5kHCin37LScTzvKx4VR
tItoN2CQUFGIK62pKinETozzufglfZlfAhCST2srIf2qjjdQDKg/edlXBbrj36a/ixhS8n1ZGuM1
sLG7O0ua1E7hFa75fgD1VOVw3jMYqdKNNrGTCmvG4uZMLjs1gC+G2Kpyx1eroMsTmcbIJ0DXrOJn
OHH+/W8ZpyRE2CbHexUWqupA3Yi7GIrefIzQFfpBZMiHnXLo4fPjEH1peYS8+Pl3P9Cuk1P24n9P
Ix5rjkVYm35e0pcUmdnFWC46rk96FG7OnuX9mx9GinboPvhyi/IVuaCnteIZXvmUi7d9gCS3vTfP
F/+Fke1gm5Mnbf5509zEtO2xs3DFwRjv2CQYKQivkhfaPLtOw6WHcwvv/hDdjwHPwanB5G0q4tGw
7ICvQn664iIFiYjkG8bI3pro89h/dWsKcFZ3+MiUEI1qpkQYN5OdE1X2iNLEv41RPPtvEURswh5z
EqDo1IeIgapRqBoQZpRdUM3AYhMcGNOlk42ZAvjvlTfKKiXr17iydU5GyQtdW/QdXNS7QMZEamcF
N2YJADjYpONTVQBgkp7QZrNMs1r0N1b2XKYnV9mh9hNbeHw0jVJngB52Wk5eK8usM4AS8P47caVu
GifZCdAI1LGZblI3Oim88FFp9mqE/SaO6SLkreCYLYJP1lwkWRRuVCgDGqWyS89H7XWapSTb1CzE
Z5OK4Ig3Ad94LI7ZPkLnxyfEYajjQ0x+NSIhUFFs3PTc1r6L+iKC1k8JpW7gaszXvIz54P6ZIGOf
QMF3er2oBbPc7z+VzG/K54zXi6+ml1+5ymAwHKTw2A0FCbv5uCZJI4JaZJYRHMyhm02t/AMZ0Qg8
/RgMx1ME7YSsOgUyMBhRL6fEnsT48BQPmHpKCFHrLn4EnQ9Kbpkbw/rhp9i3bd3SNzsqgFR2G2Ui
m4/NuT6KU3tACn9cSmmjwSBsVSPzKdhmqaoaKy1hhry8V9iW3uk1Ner8e/gRyKf+9ezWajNXn7BP
pHQyCrOSUqCWJiPJal85K2SD2kBuSgHQ6ZauHvaleMAlQe43t9Np4BCtYuKWeKS7AqwnrMeq60d+
YoM2ADaZVT+LdbQZNmrhIirHOIt6Tw90sjAJXG+oajzzBJN0UGxB4cbYD23RlHA9JJSY6eNH6PCa
WMLTBsK9zh49IQgnKdKW+0DYSg+ydi+kgC3NwpncCE5fypBouxe9TLErr8TRM8MJMMLRTfRXgrBI
mPP5VhYATmyg7ItM5PlruU/ZYDUOzhjvApqPlPclSVvSnNHOkOjHLYM+5eGArkere+ffkESsupDn
HvCPnmQOcHrEuQfSmJSansY53SbsfXP/6JRfgnBbv3dRMEKfmbcrOjl4W9Ui3z/7jALEaI/3G3Xo
v1vUecxM3e1CyNb2YJBIx66O8O40u06HGChyrhOKW6D9g7MagDuiixT2xSSFyKlWKA1owEOeygS3
yN7kxQKlTaT1ZznzcfMm6VArL8c87MryY1zuGatm9yQd872RhA2Jp0++j14aQl229EIhdpJ/oY2g
Aolm+PqJiVlZvyrlA0PGKfFbYgv77opZnUIDNG2eJYdpf2QWxiCST4+yqN4idqKU4hiDeFnHc+G6
ox4fV56WXO69vGnI5au2le3DtRQWOll+rnyNBnU45TqbKHH92qP8SjAwD7MREpWO7BflIvoMNehT
o4pEPUUCClw445gLViiRqwwO/vV7jJ7OF0Z/+4771s2/yHYywXIX658SPcNfollTkNshVjlbDdDx
K4R39OxQVwIwb9/yRuQW8pW5Zss3SpRFYvl8pORZeiXAITngp0pG0yTZiE64tcA1rUgGTRzSAE5S
4TmF+rDjEin4nidcSPsRzVPGwE6nAXsKdnz0FDhRleJEfyYfRFqzOPhhk4DLov5GsMZBQg2z9K22
u6v24H1vKSRe3ZhFW6cg0blg64MVOQDfW9JJPF78PulqNc2Soxx79zV5rrq9gS+BQr//uSh3EKEf
2ope6n8XxQ0pg0Ue+t+jR4bjsbK/dhsS2AKiW7oanCxwcMxtbYHWwVLKBdXCX6VnQmyF6Msom3oj
AA9Rq/tJVCm+k4jaUDLEBQWfiwLMdjb14jBq9XzYOu9wxIcArsWzzLtVfMzItKm4T43I66IzL64c
XlaLHm1ON8V/fr0N5Nbw9/cvshyLyffRy+GFV9dLAtFhie6BFLDNTCpwUTa0sBQvhKYGVJT/8alb
1NrmS9W/AebUSXWC74tmgaLKV+/jst53tCFbYl0FjItXPgDgqnPU3hhavOsU16X8HMwKQvK+4uPN
GegGwLkYYG76b7mI5+49AmSykHI/5Xeg/Uw9mp+1emIBNUmnL5IY1MYZp6OvBu1ERUIeaZG+62HZ
jmiE5kM6+hRJxbt28aeDrVCUiQWfJVSskdSu1OyNvrYaeYXdmmhL++sPbUtss2obvS0q5OOU/t4e
P32dLYOnDWUJq+TDvqqUHlgvGBRHGsTVWkPSOdIJ6dzkEfBX3UNDJwCZYxqj2Q5WAGzKeWuL20rA
qIWqUeFMqdge4JVLYxNUhXnvM3Qg/uMjrQbz7dapWz6PaH+gh5Jag6/PqiP8AkCF4HxjNCH8xEkZ
2KybqB7AnyIKWE9p12G7OeVD6dnoYYObTz6SB+tphipgmzOMuqklXe+se1MsBqW9vj3U6pXvstUx
mzz9gS3AD69UJiSpnYjmFyI1rDY/eH4vAR1F2DL6FSsxyhm32vbSmzciqAn7n7VeF0SPUQLHH5h7
6zTWwWI0UqoMGioe0eqmkZ6j4ICuHl/WlI+lBQsPYJknMM9D9Tg01m+cwI2Y8YWdZjlQNp8+Jwv0
ObW+LpDsQMMJr9ozvOBBTT0VjNJGtaMJmdrUKys7LW5HILEaPO6J80zfwBlezPaxFdpGfiqmuGYb
k9iofoUTXzeONP09YUz16tGbqMjZAf9pqFu4xhHRoYEuUWRvysn/fYxfMR2p/cAdsdr4M4JmQAe5
qpfKD0u8rj6atJ+Xu8re64NVgjtDTGJh0xd0s3+LHIwwUKQQmRAo+f7E7pkWeZVD5U+RyobpVsxx
iCXYP0LhRTYlnmidXgO5d34k3tojaZsuuAmibAoh2Y5XY75Lwy8aZgGtHY+PuhsoAofIHOHDPPGd
JluiVsnHqqB7avmDSm5OoOfEbC1FGlVBZyysdjN9CUbQ/52NhM2xZygatjdNhlixfLH9dID2nExV
1gvUhrC4Eb2DTvElXcxsk3PUufRC5RhS2l74vQctgj5FRR2ytPMqNHiFfBqX2qEg7KfENrESysJv
TbsnyxE/Hjkn+Wb9wWhe+5Lid0gJZ/w6kBRvcd6cmlIrZ+JEA1DPSr2SJVzd1FCWlC+UAX6ZVA3m
SSjgxeSBrvHPe2b/ChskPJ5UoME6WYSNkB27LNBDUP6qmD9qyI42VHwyzx7lwI947fJhWxelcqV0
zwtV0//iGqAHHjNz4SxvOsiRvKwZTEcns13xtE/xsAgsuxp4abHSXAcBo2uUr6MG2Xe1gTFPCxd+
HyoluxubsR9ykgam2CJeXSC5X7F/UUgZ8rXLDy4FcWrGoMDlF0rrUR0y3OuCXNwb7ZyevJuQm51o
KHPZ3IsfxdKFEQw9hUv8y76WanJojOpAfJQ5ikYRsT1qHyJbFA026bZ3E2v2wdb3DoYO5V369D9m
JoDf+HbiUukOGMLC3DiDf2Jz9ndcoXHKlFpjNY/q3wTcqhEUbvKLiSHU1FRqBURqMmetr/PcXCu5
zyZQhbJGTpxP5GguJ6M+HvRaJ5VsU4pL+Y2P74hiB0TypAZRpiPLT4QOpsL9q22oE0BU/+WKGlPy
wo2vcIIuwVBNGWA2QeiLptI2Qj8m209HtS6H4qMs42+K/y8/vjlddhbCJz4zirGJ4E6Kc/ssP8Fx
V17IvoxoSNB+QsdxNMS4PM2jRID0vYGE9PAhV46iJbUC/r2K2JHZWzSySY2NiGadqzq7OiGU1raj
wfb8JBFl7CeWdZXV0YQ9JnOZVQTMjZBbmPHs+nBcBUdD1wacAU7yYhpbYkM/8rTQfLtWUsrkQHys
68eFFP600COL2KsuYbBTSt3oGJWQ5f1LMaIgCGjVaLRNXGV0HX0lMbwns84wH6b2dElM6Z6p50QR
Dlr7Gob5LiAsqvfngRrjgd5TBMTDv1kW0lbx+p2NfbYre31cW4xXk2lrpA/TnDT3PQgRe+nm5kdo
fo/FguJ9zzW0hbvwLRsCSfIdE547Ozz+9wtKxhtkiwSIyEWTYBd8KNt4xMWbPxDyHjDSFSHbvYQh
XoZSwWJLyw8HXPmrgI8PshnvzIayRX0VinDN8gLUQqyz29OtY69yCx5hiQs8LP4fAM5OaP+TMQGp
wtbdwzhKifwU9tTUx1wjOqjWXNQ6s3f3c7tf793DqW9gHB0d9Xzd10wJjX58m3Gs3rmfT6So1prf
kw2eCQnCiSzuLB+PbgKBRZte1PtjQLp5+NcWPQW1CD7rQRyHuPAek3SJAPN6pbVVh1XUMW4A9wnG
Uv4LdhKlQJIFVrwAAg+cmJ0xGL5/AmuzUmcDP3J3oS3TAso20UU7u2+rAGQrkNYNFs1l+d/etLe0
RBVSry9tNddVMwVR4S0D2qF7GaxiC7R51frzOSGpGN712QVxCHGFadjjYBWJ3r1ckgYHHaIrDe7G
eGsXmmAHQQ09ZX0lbHEFLARQRooBpkV1G6RX7/CYVhOLgJykCZbBxvN7rcL7wbN0YuZH9wOBtSu1
y1TAdsiz0iBBvq9OXQQml6BHfJcmPnMMsKwOUNekTB1TeyPk/ij48ulT0CTfjfWpxX0YENuCvUMh
ZP3vWIKw45D7vcXbeSNZtN6njYtL1hffM6BQvlivgf9RTJhR2YwAbXX+hkg/+2iY51ybjZRzDMy2
GA+NDL+8auOTRt7jLxiWhtgwomFoCVtbTzI4n2+SSJfKfS5Au/Kk7/DynrOvUZIXe4pckrYb92KH
WM03Afw4smS594C2tey/Krw1al5uuMAzSQ2WB2XgahkXrxNDSeHeH1RAvQlRzYHkOi7S/udPpxV+
ggaRE/nvrLsfBv0c4Ra2bh9t9D81KoKjweIxZWTi3YcJHM+/JH3u5koPR7R38Ve1r8v3kJSCNYmu
nZZeEwC/94KpYCbomALW4ON6JUZf6/uQl1c0QeGQ3EnCxi/jDam8sgpu0/qgsLCDXAwfXnGZQ+S3
cyz/PAUOkc5ciSMkuFpuxt7OUcqrULhgMTjD/LV3LE99HOyQHXVzWkF3RhEVvhXb/ggN8mKbD7Gh
ThnHuvPTbA6yCKG0Iox6X2tLTooPr3ApAn18K5mbsacUVyEN7RLaIPI+O8EvaPGtsZ4tRCXjcLqX
7p/HSFGKaN6rTWm4HuFeTrpqBm4Iq8dxaMfoRS7Rhd26tB2I38BtC0IDjYUSoj+GnOAOaq7y00Nj
zWfz9PfnDjKyK3vWihnhbCxIPuNABdiM5v2GK39v/dg7laf731g+1KtuoFn2+cMyzh0l1/H2VZkQ
iT5UERR6uKKwTi33sTEJOnzcyVk2se/EucdhPhsPgYd0VkATtfH/JC9FBLTI2zEbF1AeXPX6Kc1t
vlAn3wapVv5LsDpOfUq5HsBSd4lTpmu5Cy06CCpT+b0GD9Z7A7TYqx+3mcry7GaN3gDhypa7xUxl
9qke4TeIZf2IRzINKGPJ1jKFluls2ZhE0zcrla7Z9tpNW2+nPbzvXQNmq7aS1IC+Cwz0GZ64it9x
GVf9bunqB6wyiENG1UCgy3Gn6+eKLhGhqlBy5rxvISYlsI4B8I7x0CBtcs+4DraP6x5m1edQ7DBk
a2P/RQ+WaKMm5hCfH71sOEVtLBktS8rhxsgRsu6ZSox1eTQNJSTR2lP2KDItp1fBbHiq2ylX09kU
fSuFSaRJsJHYbgblmk/pmCoSBHh6zvlr4JFdpotINKyL6nUWRjEVpec7P7JcSCqTUOKWR1kYMO5v
3RhsOKC2izcCQG0UcUAiHgKHGiWHfKA6U7Il2wtpNR16XlumuJYeKX+rhvRXPT3oGly9kBCdaI0T
WUOoRqtewRQukAlkBIs37BwB7cycfedf4c+nxoqYszsSxl6TDAori+R8XoGIEsQ48ye514IEvU7B
CVkeflBBYB5OOobxBOeKrY2pmnmYwrplLNirYrnEqvuCbPCkTVJSy9qNihyfHZ+S5MMoqX/2aCmf
ssVWox08O+Fm0tTkqOD1ZKzJkXAv/X61A88ncvJlZrbYbb3VQPe7xL3ydaV46hLhH1ksNugmlblM
2PPs47XD1gaD8RrMjPIKHssf2dvy7v2mi90JuaJTF3I2v58BiY0RwSuhzCVqdJKV95ynB7i82NNE
Sica2oPDJ+RcKc22I19djdtl7KmquXDi79A1wadc5bkQS0IMlgqc+xomWlauk6d+QJUu80lFya1y
C5Nww0S0N6Tldu72M2/XwZ5mvXnhme0LJF3sFB9NgspyMFw82u4yN6PwZ5meYCJLI9vfAmLjYnMI
+P+EOPkixNiaP7F1Qabaxdc2TAPh+jDEruiwpbPb8tFFynsK+hYAuUiDhHHUxdBdGybDYDf84XOX
F7LbHDadZeE6nuf5lSgcFjm3mDVEdLWYnNwtO22bv9YYdYAPPRZ2zVqlW1MR+r5fXYCxdKlhx3HC
za+VKHjfjkXPd0X/YGikmN2zHGmErRRGGJISSKZvaKFDosOYbaXPiH2b6nWXJ+oV09vU0jkZM7iR
TYdyHaXWJ0iRle92uSBY/nCSDywBEujkBNqXm1CidGPEJg9MugdGrb2M+tUOGAGy7+JHK3X7KM5S
jbXkSwRShi2Dk10yiryCJB/hm7xFhExL0ulMU1QlZXkI+E6HX6K7kKT15VYUj4qQXkYvTymGLral
a4aegkCkgs+7myDtyDcIpOqJ0w5HX+8b0tU/PCaQr/O3MioZqPNCT/ECi1vBO5GhJhQKdoTvzAii
Hdk3BtoNIyBhY3nzKlJwwe1+4dCZZWPhny391jMLAlQ+YUbC60/PsRQQkPecZqHYQbneONquR9il
6JR3tFRRRSA+wk/ShK9O374csIlX9/QsS6u6lKRdw8Kl/RiWrax7bICEAXL6pbCqjM5EGNMjh2oY
kcNwTEJDJ0L/L2j7p4Y+XvHH0rttjd4vgtkJ5q71uxoekWTzX8OPVPPN+tXTWYg+W8dE7FLVvqNS
KUYq4dZvj5LdZwH8QAdAyOrO4X0N3r+myOh5MXYk6btZk2PUK+bhXp9Qj/IlFV0Y4h58XFxp/qXa
JZn+jZdBMX3xkAf0bi8ZoMStu71fwO8mx7adrGkfbrwzuGtbgsf3dEa4UngZ/9ArkF3/1pxuDpKh
d6udRT8LLXmbrKVLR+/XJHzefKZGZZRgqwvNCM/SeSaxy+ncghTpFgT2I3MViYOCf0DYfqE19Uu8
3DyIldkysT4fcAZKyYVbxTWNZg30pEBT0swsY/2tnwZTXecwp80F35PLpurjQwVZngydDVOSnIEV
ENUxs8HacAJtEvjXiedhvivtggfZGlT8rLdcDMBXGqiVlZ9QNQZePieJmJgO9xpPOjPD8FBU2fGO
Z8V8F9FD6a8H89BK+oFXm5pIzRa/MG7SVBtgaJVHKhkGesDBI3nE+fo9JzoCd3WW9LvMlo3HUlZb
0h2r+jeEi/hFQGl9w6ohldIl7Hm7h3RGHgjWD1y20PQsNPdBat72yOxXpOyxJ/20OlBlfqGZ00i+
4QdLqRr8l74mzGOch5Q1B4TsMRACayt2pA1ijnsA1+ybVr5rDyK6PgxJhglxj3RznOX2ZNMkD4YP
C5mEqk70vY5o3be1oq1fu7dl9TmTUIhjNDKZibjZ6+gNsBU7co4XqsVYSoo2sYvDdylA2jWlOnMK
i7REHA91eg9NmdpZOkXK1TkY+Fp+cv6ZfxFzX9DE69LUCzDfIMn+DrXziYKbbzZ+iJorQEKMpklJ
ixCc4/0x8X5dhFGmmgsKsDAdk4BobqmTpYQeLVtPj9O40wBHOyq8HYWXbb8bq8df4RYggZqfl+W5
HnkTB4YTu8OzVQ8hykuliKTTlMiHxpP9tKl8x+MsXh4Ug/j7u3oMjUx2//78jT4QPEw3VkWfmAHN
WiMrAkK2LF7GS9mqIrae0zRRBn97ZQDmAzl2mQe9G/aDncGmzAYivsnQJBsGM4H0XToEEOyYGier
0k2spJYHk/VC/WNKs/+9GsVg+P0yccK3SdHPk2+9tfv0zrBJqYpv5OUxN+/l1tZSSfkwBXXOA4m0
MDmYnDmt7wTk4h/yLEAce8OhJozXiWhBIgDn+RqJs5aQ2+Cihe3hoTb6ak/7jsFzUxG47NjcYcwG
dixpMl3FwUAUu0CmrPV8wbDfToMMvYcJjn2IyhwfAe4xJCxWX1XlC4coyaUnV8bQbpBfIfYDvPuL
mWYm4OqBMmYy6CVVD/b/3GpjAgof2evteXG2D/6pJCm1FG7bi0mmrNC7iBeYDDU8Jf4yH5GAAKpO
n/OLyHaH4YgUtz2ugbTPswl7ipTd6QJLLAUT94jIXWpdoPPso5YqM5CCQ4gV16S9iAJI58v+HoCf
tZ6bYeWkCcCxPfNoVyNcu08T5n7y54121KetTv2IiJme/BHGajCTmvtFTLMEvscAmnHomtDHxfil
UxTEagQyQO1K4WfTi8Quv3BLtso+x+85GqXPFOrWTVhhLDO+U5x/D/A4KsxS5NQcd6zoDTgK5fla
pQvnd7JocFNPlYebjGGfd4rsN1lUlGX6bDxjcZxZaVlNstRQmaTRDBRDynSwb+4QXDw07SVGeHrf
sjBpRZAjlWHFywcIrNBpb6awatLSzvHh//0vUxPks+oZWAFJK8kgvKLD5c8uBrO3bpgNcZaeMwDL
QiJHSzXAyGyyuN42nTu6fZqWZ7orAChyj75S9XjZg4dASfEJzheDXhJV696sI6GarBHFApyJYgCi
yQ6JqVeDEBPFHxC+g7XKrXbGUuCecVMlBtPy/Zn9gsIOf+2B1K+vLBp6H4TevYwBCKWNqRYSamjs
YkbK5T1mTagdaQJ3/A6SLaB2m8K2s7phJU0G7d3B9RGxUZFmCaM/xOhup7K6QPRli3cRYQXwXjyA
7yJ+hFWY8H8YHlRp06xb5TBOFtLzyRReZ7slJ//Ng7z018hZcNUximcD2t2Ohff1fWK3GvQ4gc9Y
rYC/GmXBEaxVKur81gHTU4+FMnrx2cVLQ0eFiZEbpIz0lx0rZQO6ab+SC+WODne1Zfr+O1e4Nivl
w7L92Dz4kpAES/rCG7sWyZJPyhz+og1XyHn0mHYv3IQmunV4//813eaIWFMLJ/Eyj7WaEjKEveIk
Cx/m9k6Ev58clzg0q/6Cg2MDxrRMhvICXn/nJT9hkLiyC5m6IQs1a3/cWMKiz8kgRScRIGHWSBjc
+EK0GPy62uOzVxyBCha9GCJxOUc4oY9x2NhZ8XNG6njsAlFOat+8bL+T6uqi1Dh5htaTLNn3/zC8
6zIvL9KEWVWZr+LXR7EJOqtLh1Dq++qY6tZu4MXf6zH+Sl96eYqsu/YF8KJdlmUhgKXvBu53n7Ob
eZ/Jo53NU+fxbhlWCRiF61R2mRpU9KTVEvqml0SuDthOcifzJmjEd7t3QKM++QMzQIM6EUynmVPA
4P38Eaiu89ohcfX7d/b20qn8tFAbVwWpSvgvOYMHwPvYMWf5rx4CWRSqNk0VYeRh9JOfy5Txmrv0
SaRpNz1EOcFTDqRjPgnCaBsJrQkdNBN+l+7RZf4DYdGL88gYGyuRSI+gfISJsrcZvL72gUnpEuL2
zWiXNo/5h2CtQQD5D3eMXIYPGaT8nBbVCqCY1a8/cuYT56VORC2bYGlN/5vm3LO10TO6yBqk4Nj8
pzjUx2rq2zNQ4tZAOZbqaOAmi4Pp26i7l4XGLarZoik8jXPehzJtbQKzFh1CeZhEt+Ynpzqz+Tu4
4Q4ETybYbYcLMYkhEXw+EyUO0U5TYG2l4zy4ofrql+/fQ7SJEWPAI8QtrXVqNKpmktPBqKBQcuau
uYEISph3l46hGpwY4UBdhWXtjBmxXj7HmvnJ3Xj9BN033kdFv1joWWJqMvJHoHKqqiOBRcaGVIaT
Z+xToEJ8hUNjzRkyCOVdICgC8uNMYyzVE5jP5qfXCrThksCX5XJ2kpz7ASQQK7BWXY5lEFsNGkpX
dpNR6ay79rFClGRA2r1iUPPbZeOadMYwd1X+DUn5m+vpcyTpGm95mki7JyCK1LfOVq//KcxWk6kB
FIpkQuAr5N+vEFQnljD8Q1zUgX+By0Q6qihhl4DRIIaLyesOR46i/+xEor5ynPn6qBlPaj8v11Bc
Aiyk5GYxxQSkkbd2fKOU9oTjxcwB6i2l3UkGGQcF5dgo+PTQjmxL/tMps7vjkEutXqiEs0Etgds2
NCis1X9LWJvaiF7c6oNPN2EpQ8aNhAhG/vnrzzXHpnqD7314m6ZcbWhaXY5+IBVjbQmBdqqs5e+B
HhD3EmjHjCS3szyrJKzNP0HFLiG5LzeSTzeQ1C0oSmY2xCnR6WMZbWW2TgHm9fTNj4oMkgTjzcT6
rcfGPq/3c4mMlTlNZkHsHMqg4Af6GiZhbRyf9abVI/apxTJtU3SF5AEYPEjJFA+JqtzJ9TWwW+py
owfk5OD/OnrpTW+go5Kz6nGk9f4ZU4VtellzX8j2RI3jNzSbRxZzDG0BOAszzFnTgZkF4I6YsP2+
Hxa3Mj53ubB8CEPCUUNNXUj77YwBWCtC27vCT/ICBk6kk/a6EFBEtglmCS2jerKd+jOKQIqT4lpL
r2UAJuO61DSIuWzoenJl8u9guauKbuEJdgoJjCkxlwgBYDkA9PNfWra5x0rOHvVpH9SiGRLa2gY4
5qrll6F8wk/2zN4Le8BG555hmDewwERG7rFYf5I8dXdns6VYDZ7P+y+Zquvd5ieYJNrp2J6+qNzK
AAhkHKmrIknMJnncUrM6cCXAPytJVxMDDkfl0B6QvV/8sTxrRDA4+TQeEgnPfZUPKuDnbfwHyNbF
7KiZ3bAc0vkg+1OP2IfhfAen9BqJ4PanX1eVRyQ7P/5vvx7z4CyhJe+mgZ0VIwS9nD6BO2r/CjWe
zfJOtjkC8JjyYSiH165EP5iFDA5ZKwPqDc7okXGH9XynqWqB++UxprWCR6A3cquUW0aIQ2LKAqdb
KZhKlGEStbT/o4qubh0W2zWwtgG1ZdAlqDNuuCNpLYfu3ztHtDLbHqPmlUxm0bA5LffK1hyecWcC
AL5N5o2HUdZWoSXSPkUWjmUEjqlCyVxmSK0btX0UkZ6aq3uEsxLVpwtzPiFzRuAdUTdwmXE2f53t
awExlIrK31d1ww9IepZffQjWnU43dpDlYFmymE9lASgdow85QHBwcD4i7D0BN3akwjuZFGkoUzhA
k1CL20p8hDvD1fUNpfefmje8BPIrRhmjrQN2d2LxYPBd8PsPLgCR9DUpJdBxm7b8pG2zm8kjuo65
MjPF4h+uMXLEa7GmkNHVIJ+qCfH9ZTkGiWvF+yyXMA+dcII2u3UItwarfkme/7RnCQAVxljmRLAo
Df/jKqq39oiD+E2r/W+O4ZCySTgcdd52NTMHvQoiED/6UCcrrQlve7rkUCekvhpDnQlpp46KECbP
TOVqZW7KTcaRh0g0xGTBrz4enCvhKNSrpb0BN2PMv1z/68AXAwoJybpLZSccG06xCcjLaz1l0gpb
C70GmnjO60azOsONSkoF91fDbZ43VSnScHxLXpSdlEX2Au9mKMohi03MYN2M46As981RERSNL7Co
GTNda3C7zbkDPGcvS/FMIMLi231CX/fyXmhjRIRRwAo3B0erHcQGWWRIVJaKbXOp25CbZLwVt6qa
Xqp3+87rzdUzF4pze0dLgA7D7ntw8y13dJgFqt47Rsxq99LHPMUjRfdEPNBxTgNM0gMZe95cti9d
eb3IAwt7U+ZiZ9HCyU92JMpR2KUBqdMUlCs5LBEOs/zBeg5BtYDcmd6UXxZJ1y0dhsGAmQR9rssc
B/KlKtbbt9qZVYbSZ4Y8VsE6pr7gWdYsknYwCSeCSBd+XOVjGTS/NPqffEdnZ/HT3kZ0vVHOG1OM
uI13jBp3w/fJP2eiaVokEtRGFOXOm0v9LzuFX6Qi2bSn7tecHzkvXkwcSZlmis5zRCSAhvjAoZ0D
CUS7sIkDX53R8+WUIAjqeRLlmrG9xIEnkb6fbulrckmzEIb1qxR+lffmaflQoXVRnaQGR8qhnIqf
7jkm1X3GuxEJUvzJev76mGmuguvb0BSdYB+0pAVDieLok938dvzi6+2rK/DgKXOEjbwvET4FG1ic
ivrcMyYFC5WqijUtaRj3N98NwEZO7AGnjCZohHIlLgTCfpPXM0JLEQO57WWviZrfL51+MYjoRXxc
5j9rj2jEZH3w+vYYan6vT4fRgeRJXhbv6S1ntQbFzMoFr3BtrQq9zYUnpCn+Ldrd3fa42umknDAV
LS8WRGDW4OkFrtK64RDBIsGTOPF3yxjwXn8D+5xtVgkEnY6bLZflnlcgr2jnqkq197u0kDhyd0ry
gOJuVGRNBajlTy6iYcQycWN50woIXwMFfMm2YmzifuomqFe1XMlj/cfyFd1cgIEGyO3P+b+v3UsA
op+qxWTXHX2O68c5jP5hj8Eo2qs4tK8ZbRJyZH9WPs4HhI3Qh6zstFDkUQNfF2dLkM1tmAj4/TTA
wSVnwJHdsuc0frzP4SAnclBVjnwLC2BX/urWTc2bECUgJ5eRIDhDM2gvy92ke48kpEVg24Ei2fPs
E2A1k6ILrJ5R4quKAymmWg/QE+sWC8+ojmuVi8QkOWEo5ceeUldsuS0xp6iw07AATKw2ESxi6wsW
f0AcsFWCX3OzUBqwGjZ5ldqnprX+jnaYq1avbgqJCDzn4uJBi7B06DSTasJlq5zUW8FbV+YdRgOW
Zh2dIF6kbM7MDtg33LvD3HVUAucs+HNVXuyecXsIC4goXGSLir9zkJ2HifECuYyE7FHzNAMl3BLL
CrSzETr2zDrEDJFUqzadXKKLnWXmbttI1RH5+q45rZt9U/K13WNB6BqclgT5Q4BWXOetJCWY1vqP
1uV7eUNsUjjcok84O2zzczM9CbP7vzX6pQfY60DRxIz0q2sXjs/Mw0FPuqJHB63O6XBC5TrrFUZ/
bgmRIg71ZtCmpXjNlaB5qF/O07h8gklrSe0tC0UuppZlo7CzzmQiLCd0qRy1g3byWt5QOrxrp+/u
MEGuFFI6DltTdpv3nGtWpRvN/N1PEV1lH8fz++EpxRGj8UKsM18x3EB8snMEtXThssg1OEmh0arR
In7nEfAOXDbWHV7cXLztvI/naRWh4U0pNSMNy9YKzxtgEQICNOZJgeRiBRnISLRRtr/pAi3oS7dw
dZ7vqB2wzI3+JQi1NbucRF7rf7S35uyJ53kT3QAxz/nWYKkqGMOAiZC8yECelxpHWxKcwkNi30/7
3HsGzs76t+M/KJ2qxG7EVILejcHgNg9PJaApx2AKCJy6fc0ErbC8KLE7RsYuZqq3qF0zrx9qBedB
2iiRzimTTH2EA9i2TDNCQHdU1HJkqi7qxhlEf2R7JWdOV4+LdQIIZ04046FbxBYt1Pj/I7Y6oeT7
w1zlOkYaKj0WpsPMUJAZwsBRlSwUkX9HgCp7nsKtz7mAkQtJhJKuiREcIl5F2nJH7H6YZJSzGYb7
hA8pBR3f6wYaI6qKho2GIuRi1chbsIIW7C1ATm1tTaTrXgPVTqmrSTef1tIAyrf0t1+MDAE9t7vV
Hb7cc2Ce2H1oTSnPa+Lq7iRZuEzG2cGXN3TAx+LkXt/8o5cTtti9H8kt3RXURZ2q7FRry0/js9Np
NJgjbJrdgfV9I+kj5x0l52mV0+LEKPalwqqk3fqd8bwr5m3C+2h6R2cO9y1CzFOOXzD5LBszJbyB
UvadJI4tpjk6y0j2KiF5/7Nwc+VAVZknmX7YyLqAr1aFv/1K8fdNryXMBpXsWZsyEvT9NpdTfkwR
72oEWEssvfJ3yERhctRP7RRroyM6VyWdhIshp6KMrItmtGAczx0duGzjjexMf7tB+afNWpOOzjpq
8ek1cILPHr8CEuc9/0vU+ck7R/hvFUc86XWHwJsfLDynLF/eBZZHux42/ijVP4aWHPYKPw9huXdO
gER0a4syXqgew/De4nxSVABUrtZl6ALBGlCNhYTch9f4PGGjJjZqkE5j7B5TuAjE5al2sZuvXe7c
ofKCOwNeewWM6VCV2nsF3aqiwMnVdQ9Q3F+enJWHe19dGxqO8wtMwwquiR+ZQiMsuL2TuMC+C6sN
vT1aw0X4PqW3pE/beeDcv8yN8YCvf6X2Z2mfHugoRpoS7ZnCRIpuMiu51pUCe+jJDSjOviod9Rnb
hACyjfbtur7/79qCL9GvfmDarLM55Eih+chuPmM6aU3aqr1kK9Kc8ITmTSF6DDl9CNg/nhedXc+Z
nstGm4wsYuLRXdyxqJSL8Mp7OR3F0rm6ytWGvVqM1m+NQ2nHHeq06X7trX/S0Vmtm1v1HpA5wBj/
5bHtfg2rknzzCkHo2ipx9tyJrjG+OI9p/lxF4yTZUdw9qX7MViEys9zRPrH77uPvKqlFtT+U4Tsb
fil9OmFRElr/L03oc4YxjokG2+QEo7Igg6YIpiGEoZMgVL3otyuDE6+nTB7epi9BiIkRt8Zv0rET
i3+VgU41IPWj9+57rthPVsx5jJnsLvCyvO9hbvmLL7KbkZQ/DudlNq19E3n/j3X+oi4HQXbZkPJ4
wJDI3EGs177O13IWHy9l3BoE2mLijk+xhr48r9oSfBLFCzCciNKcXtFCAiPto3B30GMcqeGXfW6n
UOPhCTDMiJSdBujGiNhzcyBKIYwTw247At0g0ZPR6DPRjALDxxCakWAuoy8cV4IDuZ0F8iUXFdzz
S8H+DZbvG2ijrHArZEAleBQpIqpRnCebymtdwv3Esb+c4dDkyMXw4zN4c2HzojM/RKiZWyJap6YU
Ag0BVbJwZg+EQonQBSR9dhJsiSDegQg9pX44/84mO18tgc8TvURWcxQLEF6iapUJxyWaRA4NHgIf
D35d6DlHbKlhmtTaXpQHiI9PpsBrjR0xijBAU1MtScfZ+w1aMZth+TgtuZ85KQcQkgWCsbyddp/1
1NAtqwGPiPRbQrQ6f6x8FdrmbiAoRKMuOVI0oP8u2Go4MArGvOO06exFvqsn1qTAIxcqEQdmrJBY
3N3I0vfBViEgq1iBWNKm5DtN/Ydg3Kc67LS/xS4KULjrKSci5wRuuEJ7Le+ERSRyd/tbZ853n1TJ
9G0yQUqyB8v70okjGE+muJ1JFXif1mLyNGio7ZiDUmo+L2mec8GOXtEGIkBmvrse13Dt/KZAsLD+
Zpr5AZoqwwbZg/2vc1lqMqfnAJcWKLl3Z96t7RNwDxFwumWLJEVfZbfQUZw0m8PcdknLgiqzWDoF
dgWfRSH5NoZ/s0m3t7nIfWuI/cr6pxSzWHaO7Kvu+OFSTVbhgMi40LMUUyqKgpTGn6/psY0jKW7m
RlLfT9QUmgZElTNBUqnnGSRz/IaE5snYdP4nSy6IX/z+tqj7oC59GpIvYG6cieVSrc/nlyJElEZn
G/uWY2uKxLGOReLESUkLdA9Dv4PfikXLZxLBOfKvSf+toP90vi9xjjTh4CSXy0WN3EtxSC5cEmk6
MLIVvw0FpyVnmehlfYQH7YQjQCpPUAazAI5A4iZaCybV0iYm+HnYimcI/0hZx/ar/IndsGbrolQN
f6HdO2yfo8pFB3ernDCKxNwWJ0RVKsojKvfpnURbkM/QTgxv9DMHsfQek60YzGZjA4oD9eVAZXyO
Y9rPPZzMpM3wmJHDcLUfRLAXwdamWCPoq0kMcDFrIpSq98Gw4KP75ybycpHc2bldqhJC9AoqhnMk
lkKH8VHuY8HvlExlMAB5Je6AdFcBnLspTcJBocrk3M0F4SJRnUuiCK9MkSLYPrNYlreHmUX/Re9w
rVOWsbalM4W1/Ez9V2Eip9/N1+rs2ezaf7PDzEpxhiIgqaHVlGSDTbkoWrprBscPTrT+VvjsXnBy
mhYH73R8vdi+vHimRvMvlRDfkU8csjby35SG4Z/I+m1O7UPci1TfTWmFUbmVHZPdlao5Hn3K15FT
TyVojRktC+oeJxAoGt4IZu+8HZWkH+AnSRWtgugo52pWVMo04xx5whHWaoxqvCNG670zTJ71cFPy
oPzAess8eepMnGSD8yQDQI3USlmWzedXmRwU4a+oqK5I7LaGBV0d/t6Ojl8lTvsMrmJsno0NAyYa
b86hZRqf8YMf7VPJmehvEVobIqoAovah+KK11irdc0OW+1PbJ+rvZB639rdRO5fAmivH7+LQBaF+
5/OJK3RmB+7xoSxrGeEWUf/KHg10ijKTBcDiI5SyR87MZfBDhiqdj7bSfUZ8glZvEWhq4siwIxjL
SvBgm7yqoPc8oXxWpGw8yU5zUtgUWrA41ofMvv173dIHzFmGDU3n6Ix4vMAc0cxrlrRR92ErTnDT
JiCFhtLzCl1yYv1BRliKnqfAp/Bz9EL81nWQe7w1Bl1lP326ZUM1WZ40bwwHvKAxIojm2zIVXn2t
9LQ8XD8DynWoLTvQa8zIZ18ims2uzeI8nmU6Cj681XA5KI3L+nZegkeXsC4ic2/vVUolCvlrtowL
OO0Xa5nVYXpMYlBZqEaETCukERs5j8jdhM+tkybN/1jLHls3oe9FIw4P/NJQ+UWhQZWDVKzE11oM
PSQxW/PBhgYlbq/Armxx2sSiK3Lo+TFussIaOMVxL40UFCitm3V+gR3rUWJAgIXw2vMjwxfl84xf
n/7bIKFlbeDYG67UiDingAVdcHR27E/0dapl/uI4TxB+kBiZO0Dg3t+YEimuoxlb0e7+MtSIsJ+k
a21VsJ+IkfUqHKQYLi/tmnA522I4ojyzY5N9BX+x86nlQrQPIxMUn17owr94bGB38wx+M4S/Wr/m
dhjVrTIY4UZK4Fi2Rjw0L0FbDC8VmADX8P7kY9nfeUHFqH5+Pn8QgPBy+m4zPOTkBIbUHCuE2+vI
txdwSiL3wMgWMHaodrSaPz7up8ehFz3fgaA91W5xEsBK5xdHmZTyIYtwIZ5Nm/rZ97WA2j7vhgi8
QzN3Dc/NM15O+COYmkj0XmxquKPWIFftIjaitvJrxP0UG8hRYjSoWAkkGtQ1zYbOreOGikG+Hm0g
QhMHayh/044GRmdIz1aFr6/2RxSqEEWGc/mhlRri2gGYkG3NKwD4+PtAUSOdMubG7lCNRABCQyW3
8jnn6TQQpu2akADSXyzNMABOf7aXrm0sR3WVGQ4AqIcNUbdX5AtfWt08e1ino1/sMRFH5wjgJkvb
WYjZFdVdJCi9gnbXU+KMWlPodvhp7Tqc+10SqyrY9qVBcQOyDPd/nK/cMfS7ZXDnS6xHetKu/e1S
hXT+dzyZZdwQ8B2l8L1FlHo5vDSRdQyTM5KBb1H/V/v1k27EWxVwlH3+yT6YKIo1ZLlSseUeAnts
YlPdR+IQnFmdyY0umP4rixme8XvUdmtXcPUaP6/0QKYLUSNPpWT8hEkYrV03Mw7rHqu4adPWxaEl
cQz88wWf82thMH/dAeq6JYQVd46dHYgHtKvU11fdypojV4R/dZDObTK7vNVX3g/ZC0oCCzLoj0Am
erUKxLMLqNDQjnn4BcBA5sqpCEor5T5DG5ypxMsJon6qo5m88QvyM06CgeSnnW55k5cYhVDin0Pm
lw/foRmnxiv3N+h498lYMo1Cky5JD1s0ggNYxwoUVW6NzH8vWYwBDk+CFHYRThg5uREO+EDrze24
Q2t6OU+1W/+oTE+OpVant414IxJF1rMAAOWR+8sLQjv8mkC6CA4h8vm0o4a74MZ8H3UueOb6nwVr
0cQH770zBGrJL1MN5ycOj5tl43KlMoSGj5dvK9vrodlZJGgywsW71I34UMaNkTNt+tNmhUNCGcvI
nxHYWPHAYYSUBq1kH2uXJH2PXoJin1JBFx5y1+YIFBlWCjH2r5z6IlwKp4NGdqxfMtkOC7N23lCm
xyrySTj8pHAG6l3+lkMc8yMfeg6rr8Ze5up8Vza7lHYbU7J007dTc/wZV/+kbX1Ykq3doIEnvHFq
o1yLZbaEGLKgvV/NFbEn+r9v6GcYgIdWN/dOqRxmE0ahfOa+XLxBqW3Xfmk6k3sY7TMniMsRPolP
7YCFOJzIizOf+4A3SOs6slMnjprEaQ9sgsM9eoCXcq2miWHxFy2/IBGN0tMmBuZ4ePJU5T43domC
rQOHBjURgG4VZGMHncj3PygASRJVvaBvGM/vEa0n8W9wFkLOj897QnBUDHvDZVTmKFWtz+1jF+TL
kd3WTMg0nN2pToN6bAJO8Bh8RebO+O6e0oQFl/tF1ItGab3gdlHVYURUWJd5thtyVl2PAFivYskU
EwrSVlNLYtNjRDROx4OfY8r0JGkmWzG+zde7DxeVmZqdmnyVznRGqQMwmlXIde9LhMW3Q1r6Zlal
ne+D1wpBeiTwDmjDGxuQXAQIceZaxtw25UCuqbfSMlCc2IHSkL7HzjWwelI6anzW+F28sJ1JCwSy
wEbaQ/H7GuiPvpYdLMYvrJN1D8xOEEqUZVBxnud4V8/71fdOeEK0Mr2KHdCgmRMyPXCsLXHs4jIu
arTBiSDhzhco4V6HuNWaatFjR82bF0uojt51Cl4JTKUcQdqpbyhETuKaLgxoN07A9g4APPsY8+ro
IbmrAdYqx5J5x5U68sq2Rj0ikNYJfHaCEMFPKY31ZAiO69yfdKmXbcTRdw7kiJj7HRz8M+ufUQRs
+QheKATxyTqenvqVncj8ttGOwBzkaNgRlc6hyAFRbCt741bLquwKgcK1ZZIHi1yQ6BF0ApLK+SN5
QxKBrwwH0YXozkNHiXKElAhHAyBu93xvz90Gsd51RQEGmEwt8NAoAuuxMtUMmn+ku2ArDwg/Ahex
bw33BzsR9AePrvRYJlTRBzqWUEn38e+/UHc+rAzQYX9Vhh9YYSNPWHbnf/zAlemYxg8yvvAI6a9D
/WMB93STGkOqVTNPDcAfFl7Slize4ymJ9CEryObRhYIobuBT+oYNzTbFMFoC8YIJwdbM979BvSPI
J92/j7KoWLZIDYwrUwlADEcOnKO0xjwwi2pzDx9ClxlQpsTfr+EcT/ySVN0oSZgb7VPLeyxu3XBU
1d8WWz3uQl+AX4FhPAArjCMDIeAbioo9vrte+u4O75ILZCH6u7QIYEDt7sDbRSi5XZtTAtDfS0Lo
CMSIcfoEUCEQQYsMk/VJOtEE/2/61Yrqkso5KFurCYUnbVX4Dyyw+LUuf5Fis3/KPDWubf4yuaQ/
SD8zOO7ENKv8Jo50PsK8a9u3GQwpNaVMAYepeZEmKrzKc2u5MRUUpCZiicVL0QZPM0ZZeWRN8yFX
vzz04z11clDy9NQku6msOZO4j8NuWimlaQ8CmvszIsRwxuNH3+spHN1Ai8ufB9fqFBkG8quy+jNE
Y/lXQmBgbAHB6Jdo/anC2HEW4ODyIzqDiOh9gB2/j83MMe0ww2gXtWnBGIE+AlzmeUlycuFaEFnQ
1K7IZm7tAPOV6K104QpmRo3v50Y3DgKIVI0Dzsunnazhpc9mPQZSszM3gQPVOXqQ6WhyVac+wuVq
b6D+Uko4myWJTXmvTianWSjkJ53Y7esfbgeKDZr2iy2kujyuPiljCUzuQzyRUf/FORTrkHNrc1cK
Q5PbMLxAI6HGFwU9Eh2NRf2+GBvVKvlAknXslOLKngSqI1PKC2B/bEtOyclUmdgVPAMrcZcVseXr
DCeeZ6yCSlrawuEj1LE4nMEcGINNM2S1OG5MxmNM7C3HRbjomvi6fTuWTE6awZkt51DcAGiAxFAo
/yUT3Dul/PJiHOKkBOoYAPu4oaCfTvF+ucUKH6p5NqCf89XT1MmUGvN0eOTeFb5plJZeHuQnUYVk
S0ad3u3p5oLXsbkNZpO3xHW0cTVAboMtRY4GjvT9f+5EQIqQA65cfr1Eq7HXSLPqct/Epc/lvcQh
wRKQjsX8Vjl921J7ZNkoyyfRMNBAC11m0nY7mGHN34FzL3IwOTj/eLYkhkEQrr1ndqI0C28zjZ/s
iaXA9BlCnN4mEWDQI5IZboVWeNh83vrhgSbyYQDu0ltfeqfO8Pe6YUvNC3FdlycWsObc06iDLTRb
N4XMCY4zcDxrSip/i77vCM9QcjaCreVaEhmwtNRE4B6S8N9ovItQYhubu+slPpoFYro5l7h1+0LA
gn+GrNBwRox/OAwmwouXLtA8kT4QEUjabr75XHnU1EwnF5GKZvNpI7stWG68c/VGsyvW720wfUTy
bHjxl3mazTeAvy7LxYT8GEHFfatcDXaXk18QGLRyV208+ILDl7EvDqxJs4z1UUo7kMp2J8QNmz5x
BWbbyqpzqyt2qW8PWwEz/9pRNBB4lLDn2OiLsZD6E496/hswyZeJwkLxc+Mgxnd7xKe7wDtiU2mD
vPLj/cSqMVf7dl8tEwn9xPURB/B4q+61JXbbHASkBc9vvgNk2V/uNuwt0jJIbHAQerbYQynMRZnK
dW+x3Fw1dP0Uvp0OYcSrhWZgKPhXFMpFBzBvsRtpgvLvFddWDtc4oIwNWZkkg/j+f4a3cCZxgGxy
Mox3Sw0ZaywdTtDxruUjsf1OgEU0AqXFAPuw6gWMiBq+TS7Gkjq/HHn74A4fQcW1IEXBYdFRSUBM
YKVItcHZslaAUGF+l1v9HspM5Nc8nKt1mx/tjNJcljLodI5rQRBJoekWGl3NepxgEIMQ78MMRvfU
khdfyoqP/dh6qeat55pXMrUoO49abAc/KFJSVyxziMcRf8r8arNJioEaigaisP0tSKqPNG8w1q21
Z1wWjzhzJQD3mvkDwEpuCQtukenNJrwaP+C95n08yOxBTCn2k9ZpN443/38+z9k7lEIA9/DPaA6D
EgjiHP4XTuYi/hUoZtkr7dbBJGI81gEekEdhMomFs3e9V4vTODnA2b13x0zyHBaa64PCWfMgbmi4
LIh/+OG+gmbSiUFjGONAXaOQunWmgOModBE/3mU/M7lA4pct/z6MhrjLGH93GHttSKn9lHsy2+zk
rQmforOR8rprcjtWR8F6Vo0eN5GdaylSTY4U5t4+ua6+LOPAZUBdS2Q5nAjhq/UGI2y6+OGrpbxa
+NtsW0WViNpHZcLAaqynT23+OxuGhDgPpL+yowuZyB0q/2VMvjsGzJfDE8bjwQSk8Lwzh/UBeeOM
KeI0X9Lw08IC5j/1ds7GCrasMjjnbvb+w+QjxtaF+p7rWA+Zhp5tmURHXL6SZYcwbS9wjZuHneq8
b64lurOmCvfThMLoujkf5kuucXp+u6zAbQSiAot2YCVV8hJ2ySKOCy24Ba0rrR2lRjcBSCSaqf0F
7vGLggwkamS26EDrUBxTK3ic0l+N/TYyMtzp7vuHBHLEGxjrXtMsMuLpNd1J4VacQemVYmA0mDfd
LAMr+AoqlTl7E+GqH1f4BjSLzoCkbZtiioZfYxSaT2I0E1m+x49IoRQPjgfwaP8MAD5JCi5J+efl
kjEqQVlLBZE6CUQUufKi6ZKXQkPgXdJ1n+wo7vzBQunXBaBDRTPbgbnzn7ESxxEKztosoLaYPksO
Ko3cuE+cgvXgm4aobmSM1Qd/22aOG87gwPhoyFV6CKgLlbtrrQefzWOhDVdaCOodbS/eZ2POIuv4
ELmaiegvmXmj9eVSuJrYAfjCAc0Y7mS1znHjRRos29Zr4UZLQnLU7unJ+SYVEk6bQBIJcXS3VLKs
ImyaN/3gT+CKnDgWpNy65GWmh/8VRYNli9rZA+r+7LYV20NrMI9A8Flf72ESY7DfNnsaUFBgvxu4
30o848JBvCtqrslCYd+WywG7YMKD6mMZweSGSKQqFA7P0lWUcx+eAH1LIYTafYmZs6zASMvqWNIG
dhCFBflJbQoAViaVeqCAwJNruW9RFVcUuMysDi0h9C8spZdqzwh0fxnQvTwFOBsVXqncgH3C05lu
O2qaLnbn9QDf/JO7B47zQz/UqKVCtFflwn5Ef/wsTyxS59oE/xLxgo2hxo/A8yJG4+wBbwh+kWy1
G1WE6IXTexVHGpwxVtrJQTubLgXBPqfJvNBKroJrG1dJuIEPozU+ku/ktjAl7GzwoliUdFgBToRD
QK3sX4KU9nIA/Z7ihYLyRooijfrwtu13MQ5gopH8uosabUpYdoIJA1pSjOKqeGHrdV4atG5F7CBc
82MStv3la0I0ry6XbcIeD3wuTCaUONhgHU9O1zZwPQwkuSRmeypSztatHqYKHBC1CY5B7VDO5QP+
AjG2poF3h+oXxPZxt7CyEyV5CFCt3OS7qibQipW4hglRef+kVL5RompBfB13GLsvORyFesA7ujW+
SpAolYYtFbiHn6JNWX+ZvWWDVNIV5r49FqtrUeTpkt0jx0dD9JkpxvV2k5qFmK592LrpgHivZ9Dn
CIo4KljMZszI81XehT5Oh1Dlapjue0M9fzGkJds+UPTbVpVMiW6OHeTG24Y3ugMbaiC79AY1FoNb
B6lrJW8Mi9HV5GewJ/aSeEXyt7376SgTinFuOzlDJ5f4d4HtopZBLDhxhthKTZRiXcFVQJPjH19V
e4bj1vyNrtpkeG8BUy5N6BDsv8ZXp19QNOvAcW67r4lwLr39kuZO7YuWlXDGzDDzoqGySYTgThMI
ryxDgWzuTtcftWOvO1KMc7g7ykEbDSF8TLulxeoSUFhF+onB+8q8btrTRcpkvEwfp9lmHfxoXgBI
3lRljLf0dDAzeEVe29PMRRuy/Mnk2mIdcHZatDylPvw3yu+DGQp86S6P64Y9apmWWTAbWX3Dpvuw
8FS0r7/5tIv3Hj4YCxCyclCZeiabvJc1K4d1brhNqPyYdw3YjE/kaa5X0yxhEdsR+0e7sXvYwyfj
qeOoGH9YbJNCiqMi8m4G/BiQsY8U2husOHTXaDIN+vS8tB8RQ/PALFXg0yZPx3fNTOvtckYuBMij
phR6zusxbGUasLInYR77K8p4h98So6+21OyCbhaNd5gTV+REZFM5IffqklvZ3zkvb5IPe3dA+8CJ
7+PAhYQocj39hhwtkvJSB3aOjDUgrH+G9VS+lr5rkjkaR09IV7gbgcQc94J75HmduKpj0Uigkk95
ElviguDhs1snAfBCnDe3AyLtvjSfng28XjM7pP7w3pORI0kRBni1uSP8Eq+XI+Zo0Y72Mtyzdzjy
PE48SAvqdXcpc7M5LSY27/QeKyPtJZUv+g1aD4VYIEomCsnELMdZ7RtV1c66PfzkPsTV/slMImhd
j3eD0xEgj27gnA7N9brdFK5AS/AMJjRUFu93OGtXi1qVfblzJgx7WBVb4jspvv5lJEgmHQ6fwbea
X8IJziPo+W0pQjLjiFsVHBasQ3KPmSdzA67d1rk6K7i04oTTawYD438jPgVPWB5RfFzSadWptKnZ
w66mAHVptZh7bUxrLU/J6fste+B1QFVS4iEyho+YYqsBrPgiopkdvyPqH7ovqPR3LtEVM3UqqDc1
FJM900ivx5kN76PQr8ko5u3a2kaNyZIEQx3gDgOaL3/HSOhV/KRmIYO6sncR6wJkZyQqK+RQvecD
w65JhXSCg06zhEBGCptHgNouA27n9EzcVwXTnx9iRh+F2SQXdz9GD19AkwuCVa22bAQyUE4ufnuE
Kd2+A45KMUGbFJgrRa0tEK6aMFkINg3muaKkNIbQ/mhdEXGnRWGpyLvoe7JHNCFZnP/A+gopHMGR
M1ZM5sd9ZyGcyN/JbN2iJTOXrn8JxXd33YQvq9TPcB6qFruaEvY0HItHyYu3XeIe3Sa0Vms8Dc0Y
q34eLa4Vi3DEsgViravRY/1R9o+SqzrSkJiej/IzcVnsIZ95I+LFxFzyBngFWalxQRZIt8MqOcii
C4tMzxO3L2eO9+QS4zET9sxOWwlPim28nM8wjXkmeflq6TZzrXl5SqoRTlJnnuKv3ACiqrVI8zq/
1cwke3YwfGdp4b2VvnnxAInZm8pPJcWCSMuXYKHnPp8DERqNHVSQfDzYtZLxGoRUoz+a/QJs2eYG
9w8sjzOPskavM6Z50rirUj9cOqyDNItRwkfgAmJ+16VN0mkfjX0I+bv9tQd4qWqF4aCE4nnS+//1
E1Q+Jh2Rx41XW/7i386etQJengFhSwvHyrBBMPWAbD0Nkd+y5o7m3D/BoTE0MxzWb0uYp1oCvTDN
gjCZUCjcLvk7Kj84aOQqJJ6nZFiDebeSTBKkkhzdKNYK6czTATMZXw2PtcsVGRor6g9YbEWyX69r
RbLySsAfkcaikMTWdi8Jov+pesYKhfwCw7SmTrO8cjc7zJhEy+zFDKJXUD3wvf8tBeTW7NuH1uJR
XVPDmrR/JU7vSoCVFLrKJkRf2g3Y3Nd4C1N2iOSZZALRKe8YJIeXrwP8V9SzFQcrHwW/TdLB6vCh
H5DUX7Pi4R4FwqrLMyulx562zi1QGJD4SqFHhcVzc7aHPbhMRPyWDF+TZcMNHPXuI53wlxzmBMWR
/teKMmbVr8TLNvefH67zIOmYT2m9uHYF13OmX+y0lAAcobwba6h1ndFUIFlsq47xq+GXfJT7uQhH
jZkb//NVMWr7LOEsbZIx+sxbuLfEa4iEFqDPnzPB9pdUVMCLCz5LnhJJTl0RTXjn1VUY/XtXXzxD
63niEOu5bN7xA77aC1iGn5wLp4UQESKY1fwqdKb5FHVJhnFHXuNT09gC1uGC0WVEuRs2bMzEYvNU
r3pt5Ah8rD7+5n+n2iRvb+1oenF3qMYOVtJJ3h6v76yj5VF7wCXt4drcNjtXNDpq32tyYWZKVwrj
YgkyI5nQp0IKmM8ol5yO7l/jVJ+QdpmuvmSPgH8vY7OxgfsN+Bezd7oo8QNuDcaqrzgGlGmuHxUG
Ny8s3L95nU4l1C3Lr+zJFq26TUfDz2RJiaBqsf2tb8qujzD9Nskliuc+8nJxZkmt4bjy2AVnizY7
FRkWd80dETVCI3MMaW9FxMpA+rZxgdlgQ3MpKvMhNTdWOtMyiJDVl68hWE6EvGKuXLKhskhOC2js
+HhqV4iMR7oHdAWVbKK7UR1t/5feEr9Gk79zkBBJT6XrVK/mV5qIPn4OwnhctTsgKAgyG62QbWnH
pkcDdiCvIUF6PPY9Oa0DpPTbsfMZ/7SeE8kg+FqN9GZPWb7d662zLH+PaMbrZmee83Wt8/FDbSXz
LEO0GLL5r55ZnPVS4ivFvlb/w/wPSlmgolF9AwbKSG0wiir3oaySV9iG6BuJzjjVVD71ajy55f8R
aztK7Cc9i8rGUdWKI+ITW+Veor2BTVRrx0Mk/3+++hZvz9uXsaRMuO3fazykp9lRbtmHVOPCJLAj
cpghwUEDG4VpsNLlGWIAU0Sa6MFBc9e9ssR9dbtPF/3Zq4AM90dFZnatd7Qa7Cmb1qY6BIV6Dut2
v7vVQKYu5UQZDQLWTpw9GRyaIsTBfSOV/mZOHusEQsajfeXL5sRGKThHUly4fGj3ZuBBfdqyw3fh
GkTUV0YN9wfO/P4o2y6N3Zx3uuIbTYxhuPFATdQBdGAWo7SO/6Wm6ML/La/PmxaaDgLc+8H6Krof
I11A2bmgADzRtqjp/AIBGpL89Cd6AivqNB186ggDukEdW2Fd7XwFyRpRHFAkT/GWRKafSc3VO5QA
MooxlaDWfE9u+/qxM40xHvWrXrppLh2ZajSu4M4TfgTXH4FATJSttX8YuI3TsnIIJ/Q1x2oOTG2d
Hj/IDB7G+WP8dUgPXXhtpGnu2Hxsd4B5xEcc0x+2gb0w62iGVXn+34XfYDj+SXYBhNkvakicpyHi
UGCdusWc67834ggCn6TdADq1XwSJiijoBEFXdQ1ts+wFAwcWfDvBeYjgacRANmCIFevnis8yN1D2
18fM8OqZ6xeETp7YUXpfqF2cN91+MCtq14jhxHTCSEmzds3PZcJkTwnuddLi2VdsMdDeUdUoBGlX
sqXsOPqJmiLNdixHrlXviB+T6c7pfeuaNVGA7wECDngkLSyB/B4OqpE0kVOfv1ZhmNcpz/PxuvZT
HweyOS8y+JZF3X5RHhk4XToh4PJeJqEYGJ0IkBo7gAWIN8BMROOjpAvX4q5/feMf7KJ8lHHCnccG
mLYYM4/TXeeKo7iDA2Z5xAcxBaJ9p6RQjEFtc69MVJk+cOM8z1ZjdP0XGCQ4sjQWLxzwU4B1zLgh
TSRlzbIx5tvj2M03DfqxXI8YWo5EeBwZDLtZzLWUFXm4F8BbL6e355AhBQJOxMWLhjRW9+nWdqvq
X2pEdUSfUO+Sy/hkESoZIdzJq5o+PrZReKd1z2F90UpHkuenAQPD4VUl4EgmriWMoAtF8szSTGTA
GT7ohSjd8cqRhvYmwDjUVGDznYECbU4O6vObNu2kSuHG0KEkjRRZ29wf1dxmFFpHKya/QLmvgTS/
6c/SPBsuW6LEdaMHVjWsoaqqpS2Hbta+Yp3rW7QhHbMc3uuDL4x2zvZQcgO+/cFNyfBRAzd/lSZ4
hJE110mefmzmtXNRk+h6SMMTWRe5DTeAKP7EHdqHp5wLGLkfvO0iP/2ynOYjO+kPVX4JDNgaGi2R
wqpmROI34QAW88BWXaNUQGHi2PBlTDf+pEQaGAXZjZRKPiATEjp+JB/vCS6J+gH3aNjuOcItStZO
8Kd3Y5SN7PTnJqNJtUKMJubefp8Xhvjfmf0PaRP4SXXMB0BxwUYyG0t0Ij76nP6bpwlLiVrMGi1A
y/NiLIT0TTGV3f/LH4c4Uq2dx2UKWGYNbgmWGZM2AETJs5QeX3k6+Ln8VXZiPfAeh+Cc6s4VX/6x
s5M6HbvBB0BQdtzjrZ08TOtfMAMor1JBpbui5B64smXnA88Z8wbbTaIL9+uvPcHuokY4MlCgG5Sy
0aIHLB0mNZz9UBAxDIUCfsjrQnThwfaphoVta2tWQsc2D6w7o130NOJsCBtwD3VtY/tL44Ku6pCW
h8YVVTyzuxIiBq6EsN9aLds2o/xGDEkiv6FO9EZa9dBRPc7KP3XRvO5SRph1i3v5jNCKEWPATMNT
+Vt26L84N23ogYFWS5/qmuncOo4kg5/3tkZUilT6GaIofBLO6Xoy6hj3xon5+eKJt/83luPh/Y7O
jbu0bRQUpQgZH+xYBt5SHnHo28DOP+oDkujvx61loS9B3BotHXaZdIxejdUHz8IVZqCF48ESIKIk
mwckTVmMyUwhj5djTz4XU/B0YEzCAjMF2+Cb0t16sdwi6/hpBntB1aIx+kCwC+uUdBJ6ovu0eZm9
AHFpA/NZii1OyYAbFP/pyaKB7xCaIEXlVBnRQBUKljSTckzjHHEy/CamBUpSPcGTrHypaAUCfvOZ
OjjGWcvZtxYvCt9Aa8ccwARTRe0T9f+mlqymz28WboSGYuoHE34WIsY/AwcjfjCgOwvLr+d6Gtr3
gaH+8mrDT9ZD4plXnLMgEY8ZLHCWoWCXalnAOJLVtVb0ldhzsYdhDzEAUaPB3/rVJNr5+rj20gQC
EP0udbo2Ar2XVHLpt+pZdQbu0U3S0knLjthnUqg1B4hVtlA6qRXt/fBTILrsQrdhTQb2wc/+bmCT
gEMikqWgnT9Ml1316FB0/8bG4NxS4XYFo6/MYmQZgUed+HwwnDlEG2UvyOD6ltML0uUthsJy7eWP
BhmZIG77BPsxc3WGgb5Ov0jn1APzYzjC9mPN4YL6H8H8FlP0VIpkwsnDSqtcODGOD2h0hOxckFqA
TM6Vxci5/ZxXlVOzs9EfaX3zxMVPUumP77h4Wa53GZp+QpYk0VLQ3t1Y/YENhRENZUmvsd2wBTXU
dfxj/3TeYhuQJYazinYN/vc4TzvkM65eFBHtWhqqQu2ygrmtC80AxOiwhXbqn0bQ0Rz2yZHQ/OJk
smR5afKkPS71QQefLvMAYgqYf8UpbLN0jOG4eQSUYSVkQ8OKPaueMW/qBuY8LDc5cyBQiG5E9fao
JJDfTKCisCTb1XoOOnbiAqZ1fgz2DLoaonajrecZVA46c2blScv+ggp+WPJDfaCabQys8HKHbq/P
e3U63zlFWELSeyJl6/uFS2+jCZHs3PMLn55l1iWLxLJ+KwV/80R1+ADPlZYaC28nA0eK4i+Xoerd
aGRRyV71C6M6UHk0+CGXIPM87y3wMLQSyIkJ5kttCJLPEiAZNN14dgcEL5yn99LS2qFeJ04YVGYx
/EAcSybF/ib6DzmqSGVu5enoDLuR8vkeeSxjbjHlesc4oSZllFbP0VhWdxfkfn/h5OkqjP3Qt1Rc
FR/xFADaPNK2sAfIA0TdVdDBoKJLRR9JWyEGZLDgO3M3+yT6VGfepsT8Xtr0f7J6uh04Dx53+cvT
/Jaaos/ZkqtkzSf6ABSMdqyeTJlBotrpcuxoL8lxj4YXzy8+Jo0Y+Cz3wO+gWYwgwiyjamcjwaov
VsHupRUceCqdAAYeNKSeNF/9+sN2j9wT7pwtxj0rW1BvhJ/yxTJt1wGztTOQbz1A5ERDCJK0beBy
PUWOQayTBgjnFuxz9ad49YFqg9OiznerRMLQRY/3CrKYOfOm5BEEDudP0pAz1pMw6HdYaM/WbBTl
7reos+GB3IAPeBRudDo9tHlO9OnGhJsMWD3i9xDaQGLfLr6uh/VedjZHqmeh5QCZlEyupKwK+YPj
9uicynJQuewX8pfZqECej23DGFcSkk0R3n+gKTn5TNIKqUYontcFKfOT6F1XQ+whzeL/onU92rUj
PSpPH54tIivUF+2I5Cap6FN7BM0Y0YeGmVT3hck1BG60Hm12kngwuBDUPpSkCIWEes0XUnwKDJ6G
zzUCp6esemNz5FReZSO6/e2AhKKPr6bDt7s4oycGjZb54+mx7mHDqTOOlAgu/fGi45asxJBsCSIW
ExWo2Jv2UDmXeCuubMbneavcRHBKFF88FX8d4iAC6nw7k57icFNuOMjXJVArryUIgu6sVsyrSBiq
XRC41GdrBE1JiosuxBhHLrXh9Vxuu0EUcFEhUUuYLxRpV05BvBLv8OsBPg4Rg2vl9TA5/mzsE7vn
rMoNc2OE4V4PhzC5rAzdHj1Hape3DWq879VZ0QI3cL+ncfuPFw5BfqVjOkNNcQkUhjR9nC1XMyB/
Ki4qMubwkCSH4+SNRviQ3U6DvwcAaw4wK7mjRLDtex5HBA1Lh/FYqDD4mLHvx531XuWdtP0gbttg
Ts5toClDMdK9m5QkxWFMCoQmkcIpeTAZ6smnhDcA/tvOMODNvsolWlYjuep61A3GCTzmfVhQ5nYS
mv0yZXWoKpD+mMbZvaEfW1zSogboB/AuYhjedtsggU83pgTpHDyYe5VtF+o/J0CXmXYGdHrC8ahm
bBiW3tTDK64yS618CPfY5lF4JvVhPo0V4gTkcUANOfmhQmWKyL7NfsXIPqBna/QuKKl4T4Hewbo5
zMG5d0hUwzthpbM1c4a1d73wuNZuKqRZCqAbJqJSGRkuk6DTcTOxuDz+EC6VDnLchVF7eQq0U+qS
IA5ZA3fqev9PiZuXhIwyd95U/LYga0RJA6qIcZOAY1k5j5bORor06IuaY8KgmyCShsLvVm1Aj5oE
PUBF4YvHiPHaup32Reot32cRZINn6YOYJ3RYFUBeNRvarnIg42v78k/XR3PbXHyrr25Ghjk0VIoG
HRZQ+nO+GBcvb7GMkO9OxcJzws3sRXdyRC7MW/ZekkuzOiMDE7+0nHOk6IBXw67bXVxu9GCRfCGH
NQCZHbPpKEW9elV/LoKa5SNoJ9/0Bjz2X4E3DioKvSYkXul4pIo8fi9l/9lE5hql3Y6c7vld+jOR
IRKvt7cb/uKqR6x2OXHgGBAgHBhH7xiCF8xriRxdUg695kiz9zKc93vOJgSQwNrkQp0rK4uU6O3M
hy3Qn/SK6bk+wj0Q4okfDo0Mch4p66X2vL1nhSwd7ZQj8/ZZfQxtQS1A7xWcE6S5q9OxtDt98xnc
9Wfz2MxtQ/rswtLq5lAJcrcUikM2ieuu9uYRe7YM2PZCFQ8SLGq/UWJ/lmJyKd+x8GLzrzfPXYNp
aXEJ+1GdcnW5mIS+UETy3TH3XSWEidNNAiAOjkAMp2HDb6sQoL1FeFzhVDm2+PRPeyZVsm/WOX3X
YOEPKaBP0cf/HiD57aUJbcSQ1llgFIL7G4raZA661+3Zj2GVoXM4feEklwXeZU3EHYDfM449wT44
LQqrDwIYlC5eesKsSxmNUr3GFFf1E8hXpPJuKpJhonC+1+QEaycPC5sx8hAmz+PYjy9KCt2h6fsn
UY4ch4igNQKDBEl0Rygpeb5HzwjDzmAesCSI5pO2qXydfImvwxbd9MSfEXUDhXR6irEfxii9PCap
vRNRjXZvHRDgw+rsPmGY0Mu1GNfFmdcWcCsMwxFMr/9wKTe3NCgQKtJxEHh/rHHuROT69ZrunLbV
AbPlo8MOb4jRRNI9tpC8TlDQmmne6ejJXwC3STYZnxD9gYwJUX0Ju0MoOSSDTsonkdLnz2MHuERO
Q5j8Z+m1A18pSJbHtMNR5owKQoinp+y01HvAvB/mLfIXN7lZfk33MW6lmNTRFrJlkFZuwoFSOCCi
4bw/4Hqb7/U8y67fsN0xrDXHkYwqYHbxs0Kpnl+k7VoKm7yFQAeVbUbbCbtnfV3h0nJVMdnQFD+7
g5lCVMHanW3waNq2sr6fjIyym8ok9d0kapg2jeupuk8CVoM4LiYbj1PvamgqRb9s9Dm9imDsz/yX
hVkekthvITMgNw4V0VFTwAVoUYCj7fisKUhh/AG+6GcD0l7zZ8iYntTDgPVvu1ZGn2OSwbH8X5CZ
P7nf/Z+agLKeCeqJ3/SPb9VspdR0tHJYPNfkJPlKmMam5YzxY5P1YAJ4NYU5orvu8I20ERt29R1B
I5fWo6DRIckDw+82ZGX51z+dsXU53Vs8RGUBhQxCFBDyCQsbdmrWcHXSwB6YIPvYr7flaR/xxY/l
V3mugdTunaILeOQOCUmYEwco1PtS9QLFoAtyZMWoJxHKM3d3eLIX5xLiRm+VOcLRddrDY4BLh2d+
FKMBZThtI2qEgSy6qOnQx7rkO/9yy5orc43u2eJrQTLci7ZeM4kNDaW/ZUqTsNZwE3QlaCXHSXK/
4MaOiD+tbx9S2PeP34142+MyJxf4igZ/00xSKHGv55qfTtZwrfWzQhNJMijdFhRURVtImyPR29CW
Su3SIwEI4kGL0+qItj4gM8vngZnAl7WdjXIJFFAZj0J+hLkudvdmpx4PXF9/jMMPP9qUAVOr4vT9
80nB+qXkkSC+MxaMSQU6qYOms6g5WIVccZMBjujQm7NfPoKoGMR+y/A/p9FlN86KYXoNmkzFsmXu
rR8AV+3in3FBrJyChVJppmbeU/b56zCb8gxOIRVyja3QAutC2gbtqy2c+SASvJOJ0H9603X/mz6V
8thaWz2E9/LJzyK4LGT+TeY9z9uZ3hnXEaU9jBoFmJmQIrA1Ix0zRy/7KqIDkRcZqjJ3dc7EKB29
LglmUQagDjCiuhsbXy/gOdir/F9KTB5A+D/KcqnRlK1GVBhPRoH0OaX3bFQ2quGaM0jZwbsd3JlW
+bSjyqWprPPtSIfx8E4tGXK2oqq1ThuvGQGGWou41hhFJ9zuxYzAR6/REsC2u2whGnRUIABlMPu5
Oemxo0iNMo6DNStZKbWB2D8URfPJkEldQiUmdZQsgcuSR+Sh+mN8Qxe2BjiLiHOgAPeEB/DNJT+l
skYnJZ8Qd778QMUbWM8KWCwKOVvbXaojVXP5Ji9CfQT4ipQqwJjPYUMGQK8EArdVb5nd5+5klZlC
du3DGAtv53ONpUsXls5W9p83VJwJ7zTbrpJWC5uSTUrbwunPOx7xxifEJJem0o6UNAP6kNVUiurt
uA5mJiOZiYbQug7bNam3MnkQfoOjwY3nIC2/PwXyhnuXsCyb34ffE7ozL8PiShBuCE1Kj4q3Ak3E
AxQ0AYqQ6lP77dLAy4aXZLanDJKU/13bk3PtqDzAct3alYnOk72r5dNw39fxejevMElCbqHTi8Lq
1852XmQjE4DLbpmGf2Houkua528gbjBYXqOyf3CFbD6WIPIR5BWkvYO8NIGPHxf5I0pfLoU7YWte
fWSuUPDsyEh3Ve+TximqUtpRRzjqCnjTBwNMGLLCscV+XiITFrBnnnRyzNI5LmZgZDYseyRLCMp7
4y2+6UVLg/VUiQcjnplBLYQsnm7UonMhURMPG1q2B8OFag/AaL2ud11IvzecMaijmdfZYSEioIiM
jFbeWTS5UcfbsPZPPh4cdnR6Jgw26jx9gUtLXW3TNN6NF/RKhZt5TxFQiqCEGRNizy6VFvpe+bdg
JhjBO932NsEmqnFjjOtKz3Rq0+0gCH8LvK3SXWpl2z03uEkSErDzpoU1tWG2UyTNM5IXTr2/s+NX
h5BF0hW6FJaM56Kz3qylUllkaQ6aCWf230z9BxF6gX0OGiIpjccg00DkGBZ7AVp/W0l90U+l+6rg
yjelOU3D0Ga/ziwJ61H+dvFpOJUI0QqZCt6KgNNku7LJ+ZGz48yUEuyJvcte0heEC1+WJcOdOWI9
JZ4yJ8zgeCgNY9jImBIplJ5G4m810WKyM9JEYeVFK6O4lVN+Q56cvGlFzzSleFd40KX76V6HNru/
l8FXcxEudPtKkB14kFYQNweHvbBs2N8U94ikGWgL91eUzOwi+cSHY3b/szWlDllAhOT2iG/4YeWh
hT88+TU7eBHnX3wMb61Vpd4Eq6jurFydSutEBIBO0lGNcpyMqC+9I7fZHt7o66naya0z/K23quDW
CY/cQPK9F/P0Ra1TsHgpA2Rbx4dSPY4g7DCCF4vpNrjU8z/wlgvSxfyctrGF6yDQFS/9AIeWZtut
sBgWwy0mWlN6MQ59Jg2Y/5Cz4OmKt4cbgt9JeHYU8JNnc2Sef+eivAaJwBA47Fycd6IheRsP7c45
sgnDWGeg9KAlHZ5odsP2S1+k+3j5TEKn5ey5bSrqU3xpXGPLEh9fufth94ONWN4Ftm6YKM/sGxzi
Sls66KbI4bkqw3xTq9y6mQVMShpD9QI3XmZRg9D3ZaK91SD0XsNMp8ngSaDrMTxx7IXFug6y6KBx
Iutx8MzhbUFaTcUeZYggiJTKNbJuwS5IWMnG1/fC4Wu4L1YC0KKC8VGGAEz+2JD7VY2ZpyJo4IeT
tiIJpoHONnxNPFimK3cNLu0LqMGMCj5j0hTtXsQ/TLnQoc2WpnSi3VdfwpfMwXcWeDTTdjr6K8rj
VKdSbtB2BqaKNEiYk/85dYhvZ7TcIyO5r7SjnURlBiNDblh3qfUBO4LPIDS10sfNq8QUUEUCv7Cl
Qdsool/eScq3A+vrxv5jUBM8VjID8+KtThvD7IGDoKIQGxIfwMCHOszZvXibuome4OeRP5lWoZyF
l+eZlL9kYlGwoIADTasxiKPZVUYAnyOGWAOMkS+C6vou+s0wt4JojtVO0mg0iptHg6f8sbf3+HJw
exmezHnBOFm288bM+zIY/khcQmRqcApI0KPflZbUk3Zajew0gszEqQrnbvm5mIgKDkhf34/CRMAL
2Cte3uR6w3A+SI/lfZbzA04mXkxSB8chufaaRNdELfsjFQ27NlIBpg60eMICeJVVnz7qUd83FZ5x
Q1gHbUHVtMsMdl5jbXlglWBzoXbZr+HFuGZiNoVr2HruhbqOXH3YYoD/bQgxVcdBTotqOTs2l2IB
cxCQoSrAUq3nAY23TccBmuIJ7mfkRM4IrUa3mb9QFKD1bmchRrFKbT7Hqys+UMo3WZOEuz2zeoOS
nL8x2KZtGo1W8bWqwwLCGivwO3lbbzWWPNZ+u0ZB3Gr5eJLfdA6oPaufqcHRCcskPuwLy47643X3
ff3SRRl9sPGHUe3iTrjQPqIQ4UcXjuxqh4iDUkcTWeR2PCzt/zXofCcrFz1nQ8IEye3W0xoo5em7
4ajjNZbFfn798BkfRBFcZN47pzXt+WqEJTtsRaO/SNhQoXUk0uBCSuqlwUQrFlWNjLGfkrzANaKN
KxGqu0NsuXNx1emCFc8i6oc04t1Mx0DkEFTJ4IWgobD+4zb58p1ErD1kuAK4H0v6pXVs0P6L05Ng
xUdmUVNGN4VskIGAs9qw+1XVJ9M7hZ65dNsDZn9DqzEK6imcbqGzgc3qUFltlYVLF4i2sx9qyg2r
7wpY1T+Lea/tiviHGOVvqOW40xVVjhP8EE5xUGZmJP3GvhU7/IbRoezu+1eT6ESVACYEl4hwIj7K
F+ZDQLuJcsnjuLWuVvxNZ1SFL8UUP1/YTFqTYv0/ID3aCztp1Fht9Sk13kNQE+omT7Cttf2ikNaf
ZpyaVABk3wWmbk4mWKVl6wR67qTditUCiiSbH/jUi0SXEmtQmC6Am1iTGgzPTZaP9/0aLtYHejar
CbJUX208iwBV4ri5RslS8Y+CPLXrtNo8GnXGne7ELTQyIwciUtYoY4vWvHOrdWJ1+i3eunaTmb8l
wcIuMzgCv/pTYsNjGSHjEJ1FkTJiLueItiOAVewZJmuA0IL+UR6syqPAT5IXBX1Szn3bNOOrc/ss
fS0rPOInupdMZSm3pdqYWp5CssZCOBW3/TUbCE/d92iLxoBkTbcxJ+inJ3syfygNndPvoUp4jm9l
cdIlYIK+9NaiyJXqsyhsEEWxOex8f/OhxOuYDVcxJbG/W1eKGuqfFDEkRsn/Hnp0vRi46rI8/Au5
I4owpn+ovmsFTHc2b4sUfTxKGZe1YZZuSUBDRpkGhjjh26rqJxfDwbWwXm4CpDHBkEzwLUNKWjae
lds3RdPqjltpO19HSh6xfVDGLrGW8EcdaRfxEgvt+E5gQN8ZswAAhXJ153zJxxZ74byCPiSB/3lI
E8kUNYzoWyQ2S9G250JDMZj0O5iArXAIRIrukLbMR/0ReMu92aHL8qg7JeJy1zjAPCihJBuKkgeU
ILrbV0UD7LC/E8mXPk0izty61FoL/hNcjfLKZyHuNlC76SV/PPO4ZWeE0uVr1vyTpsNwP8aTN2Xt
mcgArjMkujhPuRT2Oe/t+mjkxGUV2pDn3eu2kgFdRvCJUC87zV8YSBTdr66XjGDoLWwOMIWWsH6Y
zWcSB5BETsCw8SXhdFFxltm9Zf17XBsebDPXRTr+W7aQWk/veGxF+/+a9nzO9KHAJqgcliHU0Q9u
N0J0mzgQUjjPj5KkMWsVHP0qEJv+bwxxyX+wbonZSZu8k94DkK0qN805sMgcRx7B8NjKDW0QNpoA
ezYsZfBAg9RWdQ2tsB5Ffzo6Ooux6CL0SbYUyDkKwgGszbsg5EIgZWJQut3rL692hJOHXtVjBhtT
ou3LkDUc0hS/WYcN8MYn7gssZKXfn4FzWHa54VUdlVSvZpOHgEH1rymqf1W6PHhUCXH3sxpit6KH
8BNdFUWJH0uJf1RZOkPJ7bsMINasNdlk7silu2TKcuoll1P9FEAJd03H7OBiufBp7eQ1pNkTddnb
riBLuCEPIHXdmRe/CAlI92UBsxTVOLBg6+FLFohsxKMHJc18PWBFKs/cpx4jb0e/n4hJNSRv5k4k
UcdfPRSUxWoA1aeCHZfXi2SKA5g9NBUFdcJFUjnoiC8TG9EqH+AKmrBJvO0pFeJ4u4hXtmFJGlc8
UMyf5PX3AT2BJaOaaeKTPjtF+JockbqgsXGEgfyDFQuVKc7X0azPGD7jq+ZMXQHDhNNflBeHc64F
8hneB/zaxqWYeTPZY9m0xk99/0e5e3fmVXjhzwPKtEIWFKfdksfAPAPki/GTkrvruSZili/LQPPU
PelbzKV+B9zVb3TwPdoYI6OLuur9TDbYRxWFZBPdo/I5FxBa7qYESTt9M4g0p3FOfv0YqMUtBROt
IEry+d0ko64NZdHVMJ9Vh8/m6QRCPlNCufAo9tLl4Shs9PqsegWODOOHcXdFrZ77eq1r7qYGJEni
BGV3rLxZZy3nE41pF+0NXbYLc/s5OlnDqXdUwuvWzqFVv3mNu/N1ZRzN4DMauZiRXKcW35s3gfTm
hSpmR5RHsQUXLlZqAoUFObdor+K66PqtbV5ztIvGWnTUSTUovqSoqWjcoLgQTKHUl7ylPBNQvC6O
ZLMt4EbnFLrswrN2qtH5b3GsQNdt0Ruy2coVLSKhQmEt4C3xEuj373MuDkwk2pSgVlDpyaLybBnq
J+0r+/iBmRpBx0fOq7aK94jYhOXtOA7piG59u3iL1C4pV4wYh2cPWeAspf9mUiKJ6tHPtpvlNHDm
TK3lzotWaUYNPfoS5zZcbNeP3dQDV9qK16IjA0T7YpMpsroU9BCOMlmkoiBHOQR3DiN8OvrkGCQ5
jIJ7KOSpyVuA7z6dr5/Lhj1V+/yHqKyeGlQm4oJEDXO1aHCv+s+Le3tM4QGgMSz+L/DiV18RJVNY
4GY5606vPJP/cUiX38Y/loL0ZXb6vBtzeP/d6m3RUy2yKPj2BsvTGz0estWI8zrCCc/IYJnyM1IS
b2i2h2AXA695PtHLjW0dni4zf89oGFHrsGfhDWHbPedgcPeJ+sbnglneWENySRWGHf8W5seWIoPu
7JJIBPl3bqlJCB9RVtnkUk3Afdi8cwAaT9timAJC3xictbHKsWOoPi3DHChhd0iBMjYNVAn1ezUt
QL4gLFoXVi1+4YK3c3zFTJbH6NKj2nF/u36hUVQPVoBydL6/BxSlOfM8ufVP26li07rBEXl3bn5+
ErfrJI6zzY6ul247pHJR1TWilkQwqtOJ0w8lX6uuHB1FrxBAYWFfe380+EC0Z4oEwkJu+/n02JeK
PgMe2t7PQiT+3Wv09rnMQAp23HWtLukAvYmaiQzTDHpFF9c5o2J02+a7C6yGW/3bDscTRQ/RFlbc
DIXsHZ4FnfykrBAVsx+9nQR03/24ujwJ6FHQcSAKOo6hUTca0FWcGZy/0ASvfb4P52Tab1jDo9QO
uPXfJhvFdi7zMdfkvEnZPPVusbT7WLxKlj1QyI2CNGBF77ZUtCu82rwSamEIDmv4Dden1FLDyK30
W7Csnna5YCbYrvYzq23QkOb/gX9jq6zXixLYQkPl0/iRrkJxORFGwvWYlOqiI8MnEFGDauzxM2zi
lu4TZOpfA5JxojB1Y2teG9qGwUb2SwS4Lg7ghZ0dRM4G+rzcB/S0JgmbjFvOWd9vj7Ge50qQO44U
Y6rzzdn4hjTFxRCu6ghbEsxYtaZ0y3X/EX2KGlvhVB5gLkojENPrPpZ+BVxwr2I51sWsbts1ksqJ
n2LNJo2gZQKNDkGudH8LBN0x1aQ8MvhyP6ZK7dSk5YFUOALIa3SWiuN6ILV6sifBmAgHeVA7W7vZ
/PGewQlWzW77HXtLtMnmlxxwdKeHaFJ1gjC4kMM1DetE7+J/L7rklCFqt9mHKHyd+4Ely/GPoCnO
1KdmnHfQGXWjzxU59YGzB/V9BdkX4PbuDARy6Go7KkOkwUsIvhIW59b5g05b5qinge0mi7E/4nK/
IsX3oAKYGtrOFvErTD6mBdmvJ81412nbLOHThGnjsu0eflslKosWt7obwq7/eva2vUcV/V3qBjRw
/e8d1mqEAzNPTEAmBCrbPhtgOKK73rXgOh9hPqE15xCvQig5vnACQ3XfNQNavlR1lWB+w3yWQ1nY
0I+2zlkn30QW14lmbs4f3dIguinIPREWRM4f9rP5kUKbUEgWQ27n2E1MtE40tM86qB/U5/laSLvl
TwvzSFatWTBgASf6LYlhYcsrAV57y9ReuSkEl2c8KRfT+Y4avmbKX0LRAAfScOpsT7n3+ZmBWv+/
WmHadfpJ8o8HBOKEWD6r2krC6DxEVf62aTi/olm5cUyIyrgCXcz5WlxYuH/plscAVgK2VSg/gokh
SSjyeljDjn4LiezLPAvD4qqwJrZkzsmOjtQHhWfD9gadUsLFJOcebvvD+irR1Csv6S4wjcKstBJ1
hybRCaYxVG6iX7b50PvTLgEiVJrEPU9mtxlRrlqK2oE4Cxy8I2Q3b8zMjV2hKd0G8b/NjpKXOULI
XIJdcuRf7/3Rr5eAKerpYdPE9pmmEZTXSyKdx8s/CRvj1qGw8ImISokBkhDXLyg+04NcqgVe9tud
lm8uvdX6YHqjjVwazp1+N0xCUsGiXQDZEFa/QacN4wk/0K7DUb9TFwY9KtPL4WhQnZ+LAA96llsg
jbD65AFrblyREiNbVsv1Fj38GtSWLr0XBRas7JvYDA2K72FFFTTDDzEaTOWtufL2ETvu3EPKNF6U
VN38MnEaRqGfjQJ7WOKYc071uBZ+B0uL/w3GHMPAj4juotEenEXqvMIOFNGRIOc16gMbSJWzgg+Z
mfl4LIz0ysVLo9NK7eJVYGUkYj0PlSgywU8/9NsmIvRHJqL2vZgg+17SXI2I1MhBM0CzHbmAgb0d
N7fojBeR98NmrdEkuDJ3ApUJ+OezE6wQrdWeassKQFWiBjiEnksnyTiFwMbGFHozTHN3h4ImCJdE
uDHsWAOPdYSMs2+YYFZPWLjTtCcywWcuz6PE5wiYEZyL9a3Z3xlhY5IxEF0GXsnv9kMLIa+GwPi6
ZxYTmiGF3vDzlCt5W3YeXuJmWJrfoCp7gcz34fUyMpwZyhK+7nDi8By+z3ZvfZseANil8WbXx+Qx
VneFFTQVtvgiHQbaHUndGKrkYOF9khXjfSmRFslZTwNUMHbOq7M8xhZzJ4oIi7kLmujG4TGm0zmS
JHm8/xFGQEVmimVv8IIHqaAM2W6D/INm/IXbZWisCIlrnkXmPy7tEJVo5sUHPJ2UK2t5Dk3aF9ro
1bV2IrsoT9XqXxVYQwHJ/6Z+eRWNuaZw3S/EiQphCSOswhZT/FjEkoMHCtPVz7v19KL3j/GHL+mc
yZZ8z2zSGd68i964/9WfaP9TItLpikuyjK3Ac30WLEcXr6vWqlM2O2wimyWgburdAef/jC1Y8xba
62ata7MVpZ7CJKP+BRPkaUk+egM5NL5sDV3woT7lh3nNUubiqy5P0u8rlDQDqpSkPIq9odwTl4Fi
oHGNzRDxPu3D2ijLXWzoGqF1k7WHJM1vU7I14F+8n50hc59ZWj1cFjPHtgdbjEJxbYpcHkSg17IT
zQRNISHH8Wmifggyri9TPm9yQLvt36GtplLNxRh+txsguiPjp//io+57abH/Hh+3zclRCHP501su
a0fUXErM4qfKSswZHRtIdViTC9ZlWKl5hgZFJCpeg94M+MN4KfJbnMihoFyJ+bTdzksbsP/MQOZT
FQiEL5SIerpf+WaJWIDCNvQfP7RRzCuFQnC9XxICr0lPGtCsvtr6DJIYbvgaAdGdHZUYvQVnBZZq
/0qJm844tw0lkX5DrBhi3OsGhCQlBsjJgO14OhZ7BHS99vjsXgZ5j0b7iZj8QsVD87Lin/CGq4q8
iNzZxKpbGtvCtagvupBgmSzQLIXWfGM4nj4omBo7h1s3e3WNtU2CG5h5euGMPiNVqluBfcrjeq44
OKrgsPHdcb2W5JswMuRHHfU0kJAQdPRJfUoAPRY2lyFdqA0qOulMqruxdWYftLNdjjQpKMnCyKmB
yeY9A1jDyX2CbwMqlV5AL2N41+U6ylsw64RkuJsZf7POIqCG0Y9Z6lTSqwUuRHGOtGdGCabHcnSW
JUqK7y4clyMe7AQFqLJW0p6ewMhw0+I5zayeQxJWjzsP1QU2qIdMS5ByCObFHMfhpVjdZqFEgH16
qAYcXuj0yKaOvcmoDLcykmOSrDoKRrb6HpaIE+g4PTCPUIHHhzXNeVBwos2gwNWniYQjpzzt6vt3
QePG5i3dSz3FQRKNedSvi+hKMt64coqAl01cJZ9sexG/zy+mvgxxIO15Ah1SzK2EB8iicV84HBs6
NkEEOcAYRuTU3afBxHnEj4FA/4ySnxjji6lo9c8zQVNPiRHQOGzQRM/3WaPvWsXQRYdLMU8gq23y
qFEWzBokRWJD2cwsUiiiBM81VRMk4sb5rC9UoWQAFamtbb2aSrmef3uB/yM4rv1e+dyBaSjeIv1e
hXrKeOIu6hSkw5ot9MpVpG5o+HYt8hLWMcHzYq0Dl17OvBXv5QgptZmbhuEm+IiON/mVJZjCIRxf
UEnHakLQuFDiMmxyHTrMCl6CiN6jmDnQybuX1ENSJcMnHOxZ8eF7qx2alB4AE2l3aYdeImm5FdQd
pc6LhbitYWL7ji0QyjiYnJ6LZN86Abuz9lBYEKRR8IAYhLaHKknW/zZ6L6GxVuYWiVMT40+6qIHm
6jbtfVIMbx91gS/y3DsS5coGdOCpkQmOXsc7HoJVSHy0QvQsJBRjFm4vgimF1xIB8/E5a0JvjH+k
BL+nt9xtKvH808m/w++fqWnAkeDQmc0trYvdtPnYaYY0Rs+pzLIZ0Tu3oteyj68p3jPjP6QSRZ/A
Xrmqf9+Hr/cKCSQijG0P+4uKeCW1hQx/oAY45n9DCRF1JFwZA2yihBfTCsJZrsb9FRiJR7Lh7k7d
LNXUfvm88IWJksChe+qHgGdMpRnIKQYH4izfSfVKsS8/P1uFeoWYEf7gvpdjqWZbbfW5SBf6sySL
TD+yQKqirWIJ1SSEQfuSm5l3A5/PVywHCxH+bS8rqzcWRM8V9eqsmZZeGGbob2tjjekPuhUBJ+8W
QKZxsrZZpAJI1Xqg+5fP2sUKIqvzxPoKLo6AbzHLGN8oLokyJhwu3Kkk6UhIF9KhI2wglr4nr6tP
phv9qsD9uBtBDYOPMEeOGDbajvbd7OtW4WlgxXKbiY8Bq8Lx+7JyOsicFUhGO45js4rfv63bXANW
ly8oKiOhjCCNFbH5ti+/+qWXRVUvZeMgEU1qAXwPPGXAEwey4XyBvMYllouI7FyHYC7CqyQj0WxY
HPbHFTa7gl2RTYbe8P5lZRhVllOSv3szVmr9gP1fcfLD41P/0Ol9S434JHgS07erz8fVlku710OW
zbiK2m2bFL6wVfSrxsHMYu8b/gob08oJ0Dj11ZVv9tjIe2flKQo7+4sQKVs+0vyvNfE+cOIp2yaT
kXJbNSA+Tp39oD7UON1JQGjMWlnDxzRQkYYRucZnfOMi5ysw4vCzITu1puWR+2sJNRX1c1kMZPQ6
4JjQcHTi/xZNVK3esOJk4W2BQnVs0frbq5/yGdchpV67oPmrY+djM9EYFZGTeGDX6cQFrRo95rPI
ngSVjRd34312HbMN6WK8o4/yABM1ISQN/SNRBioA18vXvRGJxCIoaE09mLqjxq6EYTNcNwLes/YT
tHBXClClF45l0+GCGLPSIexqac7WhEUzTPTTbgWXdqX7LtSHgwTYdjTt7cKjSca0YQHLbZVJCRAi
rTb1jnN2ahjZTt6jW5/umkeu3vW3oTPd0MmOfjobeB2m6IQJQiLoBU334VBtn1Fu+PjejXW1Eh52
4smhjmotCaYxq3iiMI5ahJd4pFguiy1s6W/+X8U3ugW9js5+M3sBgtO7XnL0YTnMoqs5guaHbkEU
yZCBnJtjWolDNDxbndoO3M8JrCRkuly9mHqT5hgCOMbeZRlNtm9+jXY+qeZ9TT9qInSSjtyVObLI
JY4lL5jfnE6Z74iLIv7pUc//eYx7wPu8foUMNMpBArjm5K3T7YPUUwr2EpPx7jEh6RGDeZML52SO
kiBDLJ0O+PVeRRCAmCDbgRiXHW6fONRPFuTXRdgYKp9IdUehxe5p6bDT717HN8dFIMKQrhEtCXu0
v0nls2af8L67VOheSQy0ElDgrtsGwMaV6wgoT5QxGeGpV2e3Rl/QCcp7Va2JLXPyimyS8hERSIja
6PjjbR190SjN6N6yrqJk51p2449TfKAdzQeY3CDr2mjMxdlsGohNPYTt+/v7y2TYSm8nQ1hHt7J5
1OVbZybs39+ZLoNZMqtT7jES4JaWF/Kyac4qn5jyv4B3UPCrNqy3JvAzdGdBRofxHSJCYqtQYyK6
A14ts4pqSqbn/AJpI8reVs6Lc6XVLntUsXcpYTaQJLMrDePy65g3Wjq+xr4NMzoDkPAS1lTEwI6M
mWik4Pl+Il9FOqQyKvONGOrUOCkGxQuahLG2Oly22dkQ4SxmVDW1KLP24kpHErm3ETAFTCaOSI9G
48gVXX0ayr6I2t7IBqtbEJl8gwk2Nrctpi1Eee0GwoOS9H5KB4OFCqgfqcDYUs+WIRBshprBOfKP
ut6wbYuXydcfak/bVm43SlYRTL7wMfTyav/XlYLwZAEFApz7m/m7Pe8j87t4vQXZfr1z8z1yOcdA
T7R876ws9axFMC9twmN3kMXTvcmVaxuT2Wjfe4Lju7YMjwInUzQ5FTLAH/ZTa++TCvvTHjHHw8/w
/4IFuQALELeU1Fy3Q4+20xhWpRsdLm2huOGUTH0f0ivmdAlQ5Jmk2bgnknpZnJSg9vhqon+mdqE6
dvlTAxyKAPFfmMMMP0fmn2azF+AAqpSidLVvPfuVgRMmcQF36bLUPgKYRhNx+0iEdEPATwEOR0gz
KPXCSI7vIkwBQ8WHj2Ts8ipScN78JtxQy2JpQeXUwa+c9+F5y9CDHhAIObEfF+D5V1qaagxtxhwT
mMj1lleBEttoKayHaYjHYgkqUlxe4AKka+NDelEosttNvUGBHpl91JPUcIz5fOIp4ADe+NL5kRF3
4HZFecXMDp//GhidlY+Astrf3ogQ5fum/zvC4ctsqivJQ/mPPaLi8dTCeOI+fFYhgKnFZvBAIk2G
qB9lrWcfFMS7SQyVRQzP7RYxn4UUvqz9mapsVvs+bPTlJbmzKJhk/bRcDNonLlnlyredfRhW+dUm
vsy2TPFR7AfpLVbWwUNqOQgMpUxJNhhDymSMYHdb80rUW2eWe+R0TvObWsStTqekT544wSnwW8O0
9gL0CMy9cYF6WP9slXjn8NzqdjtQZL76pOUzoO0tQ4HQLNmfVDVemteRvw3YKItZPNJWUOWsHDgE
eAO4IcyEZpvj3lcCF5VsyJKsFXEcfH062TlePkwAzpCSFtBBFveHg+1T1+qGw1jwTH+NdYgdddyo
jG47y5+FG+VsnZFfSOpDS7xg1BwCR1+D1qwuBPAJuOeJ89Hbqg2QNsXpsoNW4DGr6/OAjOEpf6sk
WEylxwxkNw5LxDI/RAtMULBqtsgHMCOE05U78fgdbA28ydxAFP5UblP6eg44+u0I3f5HN7u7nZbI
pq3AYlZv6M1i07OskJYGX1VZzQ/73H5zHCYZkuKrqgTBcE2hqyUBpyzE6nQetsZnZG1g+L2cXSnx
4+YAVCWlOJ2768G9WxPS6+hisgMjAYcBtALbQgyAP+5gnVZGfn1xmmvoaLljOLX/L98ROnfceGjs
4JP3hKDCRxOAcvQiLxalmONAHT1+lIp0x27DMVw8mXHhPKivE8HhmNmLPAgXNnL22V/RJvYAvLdf
pZFYVdPgf4Fbd1rCxi9jC35bqGpl2NQ+wyXfKxqiB/yRebGDkp5GgAdq/9qZP+l5hu+RZbJCxseN
6ILGJFgWhNoc8luF8hMwzcfQTIGZp5hjESTdaxUpxWsC+Pfj8QjvbjwHnEZ4JplnTDFIBAU9tq8B
vcNFm0/bisocf/qOB0qhF6z8K7S+Y7h+fhW/tAxke1MJjNS9qNb3h2vKTGPCdAqktB1l0kMJoUAM
6FEhYzF+QQUI601oNyt7bTBeUY/Ow1IuHqQ5m6vB2nBzkdbApxLU/sFm9TfBbmSq6dUegyFgvy4I
ZSTUMeekqCX1YzbjN/2vkYthf2TS562m8IXqJ6L8Sx/s6rJQP8+c+JB1ewOZ5FkQjjyCukHuyceo
igERORPe1KeqOYC4HeqXQXttMsSyLtyIUKbkCidHFu1/0IAM0n1E/zK8qmaN+k2yqXeX7M9Q+vHy
qU9F84pxL5jbnHFPp706h8Os1mG2kVgMVy1cfFooHDVPZfNrE53d1s9LDDxioUHJYu++4JGLfFzP
UWcf9riD5Cfwo5CKfXEbGKpYhI0TPZu4VMxWO8zflH18VUj8wJOm+Eb6W6IeTXfqL5rO/70PauED
SCiS5yKzL8iLOiFBNip4gTuqaH32w9ikZ0hd104Mh2DnYZpPR3qr7g/YcNPR+OXSIDPNdNVWxrmM
ha2Uvcgsmeu68yP/UAm5yv8TR/UCpPxyywKBOYbdP5jdoC3fV4tzvQyn5M01CUGuOKNzAQw7pN/R
XHsqq384wurVE5DVER6XV+XVwGfxy7NH0987dhCq7NOwk/sANNhXB5qUzFfvM0OuTmnt4pPYPYs6
4S/GwL8ZNIIy1x+NZvQc5UO7LSt2hvU1P3BGliM9ZEELxP74UD1wZJCtidPDeH5wK9Y1t1qAVTAq
JDfTfDiV18YZKgGfV+c/jgu5oUc3E9P0ljHQXXrrXBGK8KiM/Q42nJyw6oadwM8hYV+bV13JwyFK
TdRqBqXwneDyjpZL/BONjDAzB/4tJ/vo7C1qd9Wdd2/cvongkds9Y9xHA5IwC4ut8aS5F4slBfeN
dmSWYS7b9n04e1V39LHR14V6YjVLzqaviMGdL38Y2HF+8UWpwexNu+LqZXGZuuQyHlktm9zys7jB
0XacyRMzY305vdlPHtAP8b1jxQV/07XqBYCe7MRAw6oUTpFBmRobazJznRA0WyvLxDP9RMKOoUzG
1Kza+vMjgNaj5+IwV0S82vPvtXDtf2WTfGxpxkP3lAX31JkyaEHpjo0c2eiT49d0mxNij6bbtTk6
1xRfQgwc3ZsA4tc49RxZkTBm/3ZLFnFzbEkeFbCoKneXE/NAmGH/bUF2iSBiSGNJqZHQXL7G122u
Kg+76G647e/hy1rXQJIOpa0dqZ4gI45IOpBLQ9fGRv8JOaNACUuAjWsoXGDnUrCJfUCBzvoG9DhL
q/PCr35B/qeIQQHDUXACY/et59djBWmxEMzGB9BdAYAmwsTIawmgkKjT4LYVUIKaCdWPohadVUeo
ZRrJcBDFy5GIkApN68wf3LdTA3DNazjJ4klsAdTnzOluP5h+oGLho8aP0/DJg+bJVNglMxYyqywB
o1ETrozLxclzkzMnra0ohwRRZNIKgC+Vf/r0Yz7mOQGWjVhqX7uhNw6N2PxEfRqe5x1ebhPAeMe/
xJWCuBzJICh19k3Q1f/59qhLLbAxJR2CLGHIkytsRn/qeQFJx4QSmsOiVlYmA4jlNNW9fHz8aHKn
B+VY02Tu6nGZwzPeb/kpuOOq+weS64a8OgCsUz87pzmsM9Nf/HEJ/y4YIzG8da9oNP+gtB0A0f4s
xGHlRHK/ggXq71AZm16AN+zC2S9LZGkPbqyloARIy5Ynxqzdor7NlebP3rCv25++xIZ8e7nySVmM
17bo0jU95/DtsujvP/CQaTAdXl33DSvQIkzuMmHBKHxTSzHYF3xP5p/X1gYupaRk/ITfGz/bXkIV
4xHyBmC8/05NTA51eY6Twsbm3jwsT1LJJOOsKLFVkjSp2W7FMP4G7L5mL79X68kz4tpReMhZ6Rqm
uT+npXLU1/nF8DQkGywXTlgkSwmyxdpwDhiEX7mbYMBUoXkVPsoz1WN9r5Z8QkIG8EgsX70KHswE
Du/OuhFtTe78ApCVMlzNCZv9clbZDLPd/rtnLm2wWSY8H3OiFj7P1JyiVHgnsw8b5MfMJEXl93vt
62nnht0cPyrSJKSbjLjfy3fWJKwqpigfuM7zrnJT5BWGSm4EJeQiKqjzkbjpnImRquqKPsp1VLqM
3OPZx28QSdtsNTX0UROLuRjn+HZhUnnFpU7PAopd114c8wDS9R+m+L9kVoSlG04Dx70pElNW2NJx
bJf4x6BEeOQbSiNkOPTRRzoZXghm4G5g7Id8zkfVrdyzpe5GS7PPH+7mPKBbhOb3knMZY617JPKD
K3fd3Srwg9J0kB/RjrMdc78laLPBRtGKFk5LAZ6nzlFrpfUXrIb3bUJNt6bXNJsKQMxkwMXSUYiH
z3oOUnWymzU5KLZnmHmO4L/u0Ya0CDLc3gf+9yMhWrJjDG39UoRrogN+Nu1BdFJr8ANvsLAcZy8y
X6jo3WCtwC2ZPSKmywbnwjObabYzhiMoTJ89UUW5DqqzukY2rbd/BbJfQ/O0ul4yDgXHon3eNz5j
U+SiwjvuTgFEq0E5E2TNPB6FDJd/ioOQhqirgMabDVsznv/0HBMrndxyDNjjkNxjZkH5GMo/0u0B
tSFujVPteruRAQQf8kepmi9tsRuLfOnbjnZMEdMfGRiFpEOTn+Z+JXI+1lfpNqDpsxuOpc9Lt1ry
3wiFfWYjahb5e5rknElEX9hTbqRn4VX7UHqaW7+WkBQoHabsAkageZbnWbDhxp4yrqeg+8OmZ+BO
/ACoVfu+nc+5a3UhF4vAgKJYSFHvh31Z+Inwncy6462NvVnYYzuY9JdP2b2TE+ufsg8CxNRARnqy
YTC6XRP/h96xndEPgurjVYIJwbc6VAP1/7C81GI+fgEXnd+7MqnPz0kxpBV9ldV0dDwV7iiRpeEM
3w/Td/uvCU6LheDYSycPHZhOyDTh0CxNfByd2Csd4NuGvnM+2s/tqIxnc8jaPLtLlIkCGjPzhH9z
DC6P5O/ZlvvwI+0VbZPFnOoXX6nr9S7gV5CIj07AhYsqO17XmMylAN7H+Fc5J2ppsuIC5WpLaYP7
58k9cVYS1jrxlN8FDNGCe+RgJJwS8BsGJdlePTBUej43NMWWxW97MKn0q9Whz7EWCLBX4lUu3uA1
NnOHE35p50/FXGILbqc/mk7tpr/mpA7JC3olkXaI4sW4XawqdnHxYRHZyLHMpbGtHfZvGUldTqn6
+HmuQRUGGxI+MY5dUOY5XOGhmOtKa6zrPIFzzkrop2+PiM0nUbm6t3vzJQzRZZg0xWm3W71vpjqw
ILeMd96DAv/sLTs07vUchwOuJ/AIj3xStcA7uuX8O+/di3pSC29JuaSYWA252NJZ9oUfnTPoH2e7
BpTqRT++heD3ID1M6TQLJ4yBe2fB3ImRPyPgqLA0p/Bf9k1B6UsSQKqocI+dcbaeetMXj/D/z9Ky
/hgcDjRRdsd8p0szWfUCBoAT3caE851fVjqLVKk2kSC363NqNdjQtT7yCaonKq9YXlQT7SCjWGcM
RZ1wrjYWkRnwf7KKaJynKp6puCNoqnYsDxYGoTv4tJvYn8Noxd5t04NNFcqgjskJnsAcjK3/Ynw6
zJuLF0nQqU8jK5DtIckkYrJAr6uLaWwo4uUpbNNJqCfHSXf+kYmO0WYPKUQFCBssdLMcYXLd+OPp
j2VIGrEd+ksxzuOsIsUR9KbAQ42qhNx8y7ryKAv+MtWf6CAgUMxrS9TjwxtQG6RWPIOZSKw73Zgk
8x362b42FN3onYrWxq9/COuiqYtkxUAUV33j3iBHpYJMP4j0ipVJDXTkiDJzVFlKIDSpE6yb18qA
7ReFgamuMUXWOYIeK9e0MBvCRq3E4cmCvN7Yfk3OWE6Q+JiBUvtpa5uE1UA7yXWDWDV/7DOez5ws
Ta3VleImam7PwC9QtIpQeGWHPaRunsKtQfn3smEacUn061lZJerLWK0j8ej5VMspBROOBqAjv0jd
m4Ec7IrShcqBve0ZDWKT+xu2ygYAt+jZQDpvIJbYiyT83JkWyxDBp6g72eP/fIEWj5+4RH8OSrdt
oSSLbrmwgKJixl41q/2PvBsKCbRq7C8CDNyyrjCNPGY/ecxXfeJ8RtNRBEb3TTZRv5fyLiujdFc7
ERy0Y8DK2GbkevsFDX9ErFb2meAYJZmKKiRi+PhhjYjtYR2GZE6XlrCnXECKAUYWXtUNFT7W31/X
CvAgILFNMu/fGk4GW5B17T/rkM2xWIpAv/GIf5Eyap0efoPobnw6fyYwwnLlxD5mK9Cay/5QFgDz
SnLJ3V0lnnRfXtEAQ32HmUM56nbvKoQjdypMgebW7v5DO8xqStcLkuehkhv7zGJtoUtGAaFyMVtM
/dDjQLAWNxN6Q/vrTYABXU4e74pQJs2N6D9KJFed/vYoIvpzn+v77cv2RaV0dyYPH0NjW6YN+ui6
voJWMumaD4cUymPUkOGsLmStWJFxoSpO1s7Oml5Yu2dZSxfQpuoSdHdpULLncJ+2veGADwREcSgM
FaZwg9ibvgdN/mS5TmkjjB5jF+On6kG28WG1So2urj55rKBjqmWOtZvw2ut2xTYYtgFGXut9S+VM
0ZTehndda8Zboe4vWSnKdJePVI2mKUPY2DkJvaAMQzHfcvp3odwTAnroYBeDorWZSx6vt9s5ZZEf
RcYwjahosM9ZJTVVG7hFIekYmDZFbkFk1XqsTT7fX+Smdajf6ViT+ExtCHXG0RCchom6XdxxUyxQ
BrIgC3ibo2p5xTRJ+lGl8plnHY1qeLlwNQFtUA6jycS3JocxUBqUKAa+XJQE6ryM+y9wALiSwvtZ
XMCxl10ffKkgzZpOdcKcY2fqSmZ73XZ7SsFVyqqRBE2XZrckKAZ7RaCUevcgaELD2Ejyclir5q10
hmjIaxnf9jlPMm3+ZXMRbJPReP0XxAFjiLmHbQSu2/aLAVtNLsjF5alH28HrpM9IkD+LggBTOj6/
ZcYCuJdnruyvLK/9xfV9zL2SXSmpVaJtsQwftQ/tdMK8BKKTBvn4uQkSc8ZE7csTPdGmKADJ1oxx
UijxQoBLm8GTjf8X+3uyJVUTvPhLkT5jHqveQ/8lPCBC+Oz1hAbcxMXKwH3lWT4pB3/5JFJM0RJw
gH4/gn5TdhUaxnWoCYSMPiR4tZqdwqElHdRHm1uIONkYlL5ic5+/+Z6soC7DoebTM+T+x2N2/aai
/6HvQo7HYTwf/jj64ytCKqOz1yLZJb/3YdDOR6R5N9nVjVkBhaIh2+o/UIDnEjecXbQmaMuTaqyX
G823zq1wCdnpynmUKYQhwhpJ9m21BuPWq9NKngt4czRCALNwdSbFGmto/9QBjldfnJ/b7Jl7Mdub
DKqIhbp68FXDDtH3LVwuYTIQmpifVTOw7i44rw4ohQ3y+EkynDlcElmLih27PvA+HDTHL8J2bN8k
fMy2ygvgHH2y2MkKMu8+Mx7tSlRYsYOr/7pV70DoozGqFbS3jxhAMLlbVTC0LSQl/Ea4L2tT+tMU
SBhz8OWkdb+d+9mmM+WqZK98S01dIAGHHPG65r1e442dBk0Yny5F0a/j72+wIvPCiXM8/vQEwo+H
czUdyV+DxV4Tdt//9SwQ0lkcQsu/ukVWH6h+FPp7FyDQJ/6gIoatDgsF+TxtS8SYKReNcZLXugkM
efB3udkHbf/gNTXkJ2ak+gdHkwpo1b3IcJXmlkRlU+bb5hYwyyT8pWzHqEZDghG32FvYL+G7VwCN
dGZL465tRiCe1x88txQbQLFirVlozeA5AGMY0iEIqVTdZbOAxVrc5QZpFYS2VAXYS/Da/nKt8qNN
6MEC4w2IZVydRfJJwsHJAGtraV2RwRJDmsAHYOTSELO4EFcdyl5sybJSPrsZCxtCQI0d0ERLqZEH
RpsWSxZa3Im9DJlHFv9Buf+UrVSv4pMECp6n+yiZL+0IPNC1gqgxYFL5RAuKX3eAsoQnVaz4pk7/
FdtJfBIKm1OmXSLhu08+fV24yqqucnU5WPRHRtlgU7UKFC7oTTQLSTkYDW7m+ETdzyohmJ2LKU8K
4aq5GlL2MvXxPTxkrG0RcIQ/4S4u3IQa4LF5aMrQ4jHw2YraeOWDikP+PXp8LVaVrTj8driaJHR9
AokbAdgTQu0r8wSranBxjvGqsptySbvc4PAWjhGJR4zW6coN3MoRGIfqR8aJITFxjxxjYOVLgvCI
gU055F1+dCgR+NuGnRp28K17nL9gwZhghXKCpqpCAlzbwhU/qrLCYZZbrNJ4GfhlZ89q9DGkb80U
rQmch2Y5JltMopKjhUd1uuuRUrPMnv9a4O6yZvRRLnouddDAgBz4sSrwy5kh8Vx3AMVMPQyHSmfb
AAOSc5q6KgNPbnluU+LJVZ4EhFbHF5M6Zv2lh1eltZYljjsjyvGpWod8UtiC8NA6/yXE+msllp+J
dA8ZAZIZl7MaRZE8snLzpPR0OlBAUyI/p157G0ycjD6KFJ63qnyy/T9dB6iOqcM3R4DBxRvZ/PJX
8OhclnKf7bff4NL2UB+v1sUAz/9XbYPuyqE+uGJc7OS/cVHua9GuOiKsNNIy6ufXVXK1ARqDGWiJ
61B3j5EVflrkLDA67Adw58BL41SFRD6kOj5IyKhJJ4ANiViiG7lmTmimiNX5RFMduROGzbG8Tc9/
nE5qN5rS8BbW5y08NC6Eo/ILEp3N4bV/T+ADdMWanyANQ7KmknQQPwInycvxnOpyBN/Na//hDeNk
oA7eTFzVtGs2ant2ZUziPinyUhs4G5lOR6Cp952clxo0YVlvs4GVxAvikmISnjChk0ElWwjIEnbF
pBACmkcmQYzjo/PvOJeqT3nAeHpIHhbxNS5Z5uMqanSx4JBTMRipAgZfgbfwIe2tCiF2+kymIXK2
Wr5SfwdMkCt1FDldhcOGDmnzZ6wjEZv96dwdJAb8S97ITBPxViULFKjkQQdX7CgGtUKlQ1VIyecC
MgoHgir2wm23s88boDDchQjnafVjjed4iN4oNi5/skJDb5Ad0fb+01Tt2+QFAhZnkjIIQmNsTvqJ
WGce7x8+Oh2z0JXY4S9IRmasMj66phPjYi8XeRbx/2P84dOBGikVaFv1G4agdI8Sx6nwjMSydiLR
jycrFGlFfwaY23xHVbqxgRKd0SWssRqM6v6BU/LVmDVMXEX1WNwrwiHFviyAJ1KBAmOy/6VR+PKP
R7OmzhPZNOppB4WoainQ6o5MosK1KGmD1u7yQzV9DqUQRL6mWuGEz5el/QuU+qPn91AqTGmvGB4W
Ts/rdRYFuh3K+BkKRLBecvH3ch1l9FDSIpoH0Cyg3tfsX31u+b7XHWxCF0IzOZFLsSrUpT9TDKie
OUB7xG8id6TZY7DOMES67rd0ErQfZCib1k1svRsru2jccl93qshrsRg8U6gzamTd2hx/Hk9txYrb
2KTf4JNZNx9gumIci4O1KWe7D2vUEEWHuHuLwQzgFakfCS1HhAgTa7ZiCQVdCPOPThGF5MdB4X8p
UlLSd8nMFa5JAFSdiNd+hy1xdVYozCY/dNVja8k/hFkLi/SKYbzrOQPYEMvxK68KFYLxBcvWLIri
85zMIC1kXPAttLR/3rea/B9ZGCdigydDjXIftcge3sUBSK8zPiQSGwvaJ6c6xozLhpVvMLuuVgz8
Ci+LGMn5xprHifwjjyBsXhNMvWG8Ei1IpHK+/xOirvodSRANTmqCpapj8iZZy0leoTOfF+4HF3a9
LL/w6aukSKCXJki2jaQKaPiw2VUT+TgPfD4Yb3i26VynI5kHqQ68Y3QTSu4Qm/i1upD1+d1kNfZF
oIMQJZkrv+9KhYq1DsU8vvxM17EubOflW01QdW/TahOrWYAEItO7GVj5WkXUbWCxbtO6BO7CS4AO
Pmj6InwdpCvhlnajhGKMaq7DFI5vW3eDt5g11u7GIy0B80P1eqfcMuF4PvvBMrSrkt+vzWwh+Jkn
INf0cXU3EiKNKvwOn1/5VXhPA2iwxXXjQd37E9LCV9o0UVmWLbJRIoXrRhpsA9hf5aOy5yOMOqEm
HOB3HaoBcbgiyhXVtcrv94cv0J/yidhJhjRbpzdjWpNB7WbixlJI6YwLQngOqhBVBV4EXwZRoLA9
0nVk4H2wAmRo9Ng1IthO5eh0oaC7zFzpUCJLV4ppnm7FEogCTclnD7UHJsmz9X0VTPfLTHOTMRT3
eRfaSLSr39gWi/C+xST6faTAFzaDVtV2H5dIIMGoFOVWkC7WTO6HH2L9eCsRS9TgvO+LAWJ1yWa4
+2jXEptxt1olgPaROJtkG7HVIhfU0DUnhywdcrI2AfocsWCuP9qwFGxARyWAWebXkD9oLI4mC31+
t+xgVs2zHhYKVpFApc6FqaNJiFzm/dhq/NxNK02z8ZjosVyLWGlycvumHdkpngvta762ngkADRrO
Lelbv6aXKXYsmWlK5PMWi1k6koJTDY/F2n9/w+NMQgd0k1aM2xXFvh1Etee5OeTTjL6xVLoIrCxs
Rjwk7CLTWR0pmXPW3ouek2SRl+5K7RTNhEc/EaJFRaxivqxrTqSvt64XdaNraYcXnnLSVc0m1UsL
VtDc6+oCLXQztCzkumax/WjgTbb7YQjVnj1OSFoNl0cH1CHU2o0+ckZQYvg2ew/ax2y/WkED59BU
sAk1t8WNcM5vlhoXdcqnm0pIvAHwbEj1HbxYp1ttdwPMIi2zzhZkpp3JF1ceoWpvG2SPBwH+7UKP
BJwXNjHprYQOyfd4bjSlK0SpAFEl1J/6E5fyHMWADApkd8qvxWGNfNcR1+9utWmbBK4ro1cK7PBA
5XIiLcF4/jIfYuEfUBpLMwWIi+An01W56Hl8/1xK+VWIeTtMH1TSpIBOZiHLjFnS4+pejPmF2wta
wGQ+vUOWxPvHqrJ/rEb5Wr2gjKC3pYf9Temu8ehDmF9RwODxG9XZpNVp9gyo4+KD+nlCx1Flmrt+
bk3WFrVhAYUScjDtcKCrcdghjsqVB1uzSntPIaxypJu3YnMlWbpLQfdWCq+fVcszmnnqfOB6pp8z
nJksBr9DxMWyMTW/6bMB7hx+8Yop0y7gvST4FzdTr+RQ+oDm6VdpUj/ngrDtLI+cTv7a1sPYUa6X
YVbKU4qmXxPo/Z7lEwdXE5WNrSTnsB6EjZNZhCGt1UbobJjVWhgUf/D8SNEzFTRvsRME5f19xL42
jKtaNZD1qiDwkokPxBrKpEW2h8KTcjYcz+zHR+YK9iF5Q90QbadtjSdU7buS4CjlO51fFV22X/Xv
yw+9DpCp67RT/5f99ka9RA6F3uqa8RqZcrMrP8Dkggke3NKxztmnonDcAtqHePWlYnF50UTzVRlo
LnQsHGVzzG1yShnwHA4NX2u0SMUXhZttiEF6TY4kUWo72TQ7CsGzWQIakppv8oEp9FckU+s7fWQ8
mFQzC/ztKTQihhXJNuFmqM3e8meWBoaDqLRJ0zqLjQ60whWpuIdesKxvBGdpyxItuP3qx8/RlChD
ZPKYA5fqVBImTogBJNIon0/mO1TqguVCBgoT2BAb8oYraraZmyT6NI0+zJn3xio0k1yqUcIObBsF
3seTlyjp4ieZklwePsmpB3apkX82MyE63duOirPIqGw/fG/5Expc+ba8f5E5sYK72IDL+tskOe8d
2VAbB5+x8nERRdFWmD34Oo0j8HiWonWy3/LQe3yWbzXgKgDTSXr9ZzZpOBilZtclqH+EXcc7+Jzf
/Ck0LL1HaUGDwBEZK0V7WNUzRxV0hU4zUWbD5cH5Ld0HrdjOThvZpqTU9sGC6LZx+PUd/HWaTaev
Amb2IkfbD08zkBTD2Q3sEFTv2ZyBjBVkytzCCHx1EZ6I7uC5dLBNGzMVkXtqnxBFWwWvYZxmYT/5
Z0iy0C6CWyn0dEjIqlJS3RXigs+BB0c7OKaLJBLKyUPvk/hV2I7xRzsC7mV4+WSfPEkeiNNySgPY
bbcEfc3O1wfdqBhmFoF9vlkZPOcUD80GFZnIhlLswIxk6fLy7c8avLGjQLcjL/cVvF3umvF058xm
Gh4Nm8szb7r4gT6ww3CqwF85NiDWYDbnDki+1+5RzCfFg7WJx9Qb/eYmkBmBh4D27KhcFa3AKj0O
sattkxZZIZyO2Zb2pk8n9gzFWj7VSk4R4wAvgNkSctwjYizY0v2lHoVeOQBrZ7IoaEON71ubpiKI
Bp5n8pU/xM670ulIyuQciYo9UaPDv7oX+tIxWr6+IhgjxefSKt92AuOl4hjSk3j4JOR8UZ9uZ5Dj
Q8QDucIVSMjpYYqq8MfKKVUTmC6kiFDcY0xPUnOFj6nbwddVEfeHbOjxoVtOnR6HcyM5nVMUifyI
ZRklepw/i2xl3fDj+e3gmVvEYxSwcTrtle2N34QuMIfmY1vLQkKaqkAne/Wads+Y0Ob6FOCyAYrD
nS0XEerM2uxohOPKN90jJi2FjLckLAOu1LE7fQ9eI+zXOQNa8dKCKfoCBfVArkXzd4LWS5A3eyhZ
dPcYbWu15ahCGngR3kejSJ6ys7ChEKwXiHNZd4VdWufsMrUFuWgVsivxTc2q8DtgRHKRckBHnwQW
wGGAqTsZ51jILrb7veKqM3G+Gz06AxEa5kCdLN9MaU4I7kW5Yl0p0deJE39lGvfdTKX3Ev6vq9M5
2WhrswV/+teUw/VRREmUZzgNX2M1HdKZ23ptCiDQakji+IFqef+VSD6d4LIUGxfbrUGWVwkxE6uD
eBgs4bIuMDi7KrtjCiVIHiT6f3CXELEeo44liJ81kuxdl23kWiEfmRJbpqMxO7r84oFfcwGlOPAY
yDd8VLEq0Kk1h0F6+mBQqxrzi/iokzsQBOzHBf/cM7hseyN28X1rio0P1nshY2DE7v6HL+d7DJw/
XJLc0k1RrgAXTNZ5hCmfjSt9dFLLRktmPmeFkea2OQs0hwp8dRAv0g80DX+J4DE/4gOlDtmFapzc
IVSC+OLA9xXLdaMbjKRXT14pEJfZiAd04xGOXytK89TYBmiIOTSSHsbrEe67WnM9pqyKayAsTDPH
mcL/rbJY4bgJyf4N++hflbmcUOdb9w2AqPyKcnwylD3zXPgdYGNM52FcbmTbEEBaNcT3q/QJWkw5
M37n3V69jutbmO2yVO4Z6OIJWSE2htcy9buvgnFMi5C4IT9VNjO4O0xg8e87xUvFowHU8xJnlMLd
plK6IKnTQs8DqMKmuqUWLEul0bvZ0xnVYPGYf2YSlcSAFgVxfXprkgwSo8taa1owQAsTCGIAGVN+
VirwBeVIiQHIggbWuubeuraa8a5wtMllOz2JgcS2rvpCx0pMjwSWFtIqEk42z83bFVwhBQxoKveg
neLk6kMlorMHURRWzwl7jAqlTiYdc1rgGdmhn6GVOMpg3foqqHIzpdLNyx26O3J2Ck+DK/fbEVgq
aMCY7Q1Z4vpMh6NzQS/69acVwQmGlLPugHgui1eYsLrlcIxgjSpbR6sHUfqQTZvGfEo/omIvhyyZ
rIOISa08cUNmEnoroLVsS0aVYrKE8yxyPwRFbKFttp373xZ8dW9ccwVTuwbl00d8nkaoJWMwbZYt
a480hEP59oObeDs783P0xA99lPUIjOSuBgQhNymYdNgxjMXkGx1VXeovgddtsAUCZk4OMJv6Cv7I
S6InvwEfoRi1vWrUN1Qv4bnmRGS1d62rng9TYkCemUmg7V+jFZuDVmZ94ZjKsKdqdrVgIHv7kksk
pUdDIKvVyfPXlhWcXFJJhmPknoxjnqc62hzVIIqbIWgSjVnR2+RQDVW3g5TYtSXD3ZMGtjiwC+am
nyks4+BIew0PEZE2Th/QEweljplpLqyec4s9P2DpvWWmf1SVy0sKqUVxEIcd/zrIqmTH/Fk8gkpU
2CkZLE+NIA78bAJ6rGXwqmLNm//07T5pr4hqonovPIkv28nYbLneluGjH7PnNxPA4I4btbVGVuWl
f6jQN3OXycTUykhwcLxWJQ9Yc5eFKr6HcF+915mXaZ3W81hnPzU3+4C1ipjnUqbVyHmmnsROua5e
X0euOk79v0d43qG4SxbU8+kruKYa2GOVz9JJn2PNTodqokWr531ZOgwIoYyIsORTSuOL3I50pIHA
xcAx1fnig7XqsdjrD94nHC7PNS838pugLf1hNeaJhrBnRZB0MOTKFQCvKCJaNUmKtgedk94KkzFo
CQzNNkg+CM2L/EkW/F+a7qYio7ohbXKh5gdeJIt4hnLfO3uznJp3VodZ32LuRnTN+FdnWTMppnXC
Au1c//eE6Dj0u9QzwywGj4t5UTpbLC/ZMbJL9+Rh4U5n0NLp3nIOY+s1UamRkPlgWjm9qTfkzsLD
O6F4CBZ/kxrHFxvfDj6SauUirerwkFBsfqIXb2P3EMaLvCY2GbwpDBk0suaorZIM3HLDGEhx58v0
S9WDTqrXrHwirVlIScc4DKUo3X4TOh7xay2Fo8/MU1wZmchRdgYbXYcyMTX9Uk/UCbgro8nvUVq6
dNDxOII2dkk3B0G0/XdYT7DgQidffxp52QV5kJee8KtxlyJkeAtLLvrnBryMl9PPmGro75pyfX78
lkB/rbMbPrslJwnRFooXcjPxxczJll1QNglHyVn1iSR/wpjEzCubOQXnUVNpUvJ5gqFMqqlL977U
HKp7xvivxo7l1hUcvCFiJM6a7VsA6ospjgQKomwqQwC/tcSq7GI3YytI5tQF8MVJ6dW0NqYWFOj4
ILjKKBKNjHUTW18h9uXk0hb5MBbmve01Ki95UmwXtfHR15w32HSqHNrxU1OcgPL7sty4mjIhM6fC
WYhD2O/OstNYr5zDkjksoB52ZsfObMLf2fIteD8itsulgDoAJGdYdfTiJ3jbZOgySJfxJl/iIKoN
i0+JalX+XdtgmPvg5geAS9A1gFuj/vuFG/v+8awa34o2XYO5PaZRBKK73fBbrSWK+m7CKpoDeOTJ
1kG/axGyME++09OLGwJrxqqgdoWlGCVdIGiBrqtXJWFeXAj1EYBL24Xh/S0z904seodSpQRn3Uxa
QjaufOyNMO/LuOhxW2AggVTodJl+iEDoPIARJ0AL1UBKRwFXJVCAU865LoFKR/lY+0di2oHkSYkE
L+/DCku2HMf+zNPiTCIwFl5wxAp+brt9GPuQxV+rK1Qd3GtVPLubisdcU+IX3Sl7V+1hXorcGZQ8
2eNkRmJ52/ySYiFCXwu/MKXLdo8ASs95firBqGwTPeTU2IY7I8HjGi8FZHEoUfWeDVS6JwBbdiuJ
GUbAVPvp9sqIIB0UpM4msuDOzUZoLs4d6dB5nP9CtrV8LDcMCeN5QQfH+MnbCShvwcs8Dg10299N
mnt3P7LuSWDMYw7QwDmtl5EOvAQY8VyCz6VOjCRuMNs41zkmw+F8usQ8RH2lsAfgxiCtGkTDYF2t
6SreRdR7AT1SFTY8CQ2rCl6oO3o9k1EJL2NRDRh8aFbAJOFNTO7neuwxK6SO10Q9LHeZweuO/vDO
C8c9pUkC0HaH9t5twmy12sRFTZfRSAZW0gylzwZ90TrQQVAjR14Q4CkB+85hXLjJHb3a0anKtsat
KD0cYpqH4Y3EKHrM20oB0tO9PSsqSIWqnna9JbgaZkuPRDiBdxpV3qzSpZit0QqGrXR8Z1nrT5L3
ujqPJ/x3REjL2pmzOOAijRxZWW9bQCiLrz1LLbc+pShIwkGaxGlzZhRE5Zr4nJhfNFiokUfeUS1o
DpFrOMGSdmQ46JuE8yNhzWTTIsIwCs4dkacYjlkNM82uesWysonO2m1/EBtdE2IZtk5z51+llBw9
R/4AjdnS2uYiv/eqrXQftMrw1/z0KE4d+j96ajFic+HJDz+8Z5nGj0bfmda46YDTsJ+OwrWp4JoW
VuVR22ruN/UGSlVSTRYjpIEvZhAb+f9DEcg/WtGoUIYR+kUj4Sk4pItOKt9pvLY2lNhZpDFL/gs5
qjov3UzAmGkzzHOXMdP0NEeKsJL0Kiy4wbu1eGySizyOJZk57NlGVrvNha7+VuEA4p5FTi/JWhqr
1j9K0oY8q9D8TCfIL3jKFMUzkAd6Gac1cYE2qRUdjjZkGGV7DObkF+pWg58C30PV3+6Kx6nL9w7b
nXgNn1wNwHTVYN/3UQ90XhWHxG4jJKiYpDUJPw4i/tAHGs3tmvAg1HA5O2as+quDNiEFqVNGqpQz
wnH84AxaZw49EqML6QLKp887UX1T8Aots2MhYK/iX8iIpTgflHtJUBuQGYkSUpoN1joKB7l5m7TH
i6I4v5Xki71VUsM9C6GtLmcXRLRqBsxkE1cVEZryqdDsVDggVYDKjEHEOOBMaL7+PfF04EY9cUrU
jzoctHIpvyRIa45Q6iHU2IbPbUZbhuDT58u30kFOe3Cgy0Rwq0M05MOM1KcNB0wiBHGV3NHpJxb+
/Xxt3PgA6asCGXGwHHlpJdP80hRmwFUP/rOsNGvXyiPn/AxvFXUYR1KuCRlB+375zfQ7jXOJGLcc
MLxcvAc7Qjidm8OUffaAJDDEz3F2ZGAHqzw3nnRp9FEPf80e0b1lFxHCrvb+OV/jXVwNsfg9nAsA
UrDBZueF2fFr/zyqU9/BvM+W7TQdaHb9elpSUKws5v4/cqLGfzktDJB1oRe+JXK4xl/JkSWCWmQy
F7ATM3t+abkXvqJCynN7eMoQOG4O+rjCJTL3d9Wdc9ZvG4xucDevv29BhwnU2zxgNSPs+ufjqfGX
RS9vMQQoqS9Wnzy+rw1xytuR9dKIA0ixyxTPd9UcIl7/pmRI1CdLCo2EPTW/17IOOTybCfJ25TIZ
bXV/S9DeVugisaf3F6GAAuY6XKfifl5MIOYKSGb0364EXKGeSNKAy/ETnU2RRXJ7Y/bFG8bis5z0
7a4D7zid7E9unNRP+rTvMV02sYTqJA96kvytKBWPwme/9/LMncjXuEkaK7p1M1qqE1t/mz1Nrfme
kIX7/5v+fOA+xUse3S3yqwzgdegSYJmfgwnyJ4t074pbfDSdLx2WHsfpqqb71Ot4+ecTbVdx1KpA
wrqLoIN5/c9lZKttiKVZh415KVOIIEradD2e+b6BrjGE0WrVAQozCvu4l0+UTxyJcWIGMWx6iX/m
VvYpTYZTEkGJPNIoRYSxUX4UDqZtKHPGL7kVBrcX9iZfxAa0ba/15L6QcH7AV1icBzJInKORy4kt
40EZmZcd4nEmI0XS+9nbC+iy7vKbUiPkO1F1sevMSA9ylmWMZdKjQ7QO4S8QeUp76w0bTqhmHQrw
Sn345/I1plN1XCKx1FlzfKJBDG6+KHb2AZyHV2LmmFGs4tKawHd0NrWWoUlqgqfq3FNUJ9j7PfEo
iQxy9dgdYPJQEwrLgEzugeWc6CK6m5LSW56/UmKn6sUqUcTxBvQWyL9rLITiS46MvRP/H9MYBsGX
mHIOYLzILkChsA9IvrTYBDoVrCxy77diqIPEXRAyVU6YzZ3MjVOY8Iq8EfJY0XsZfbnzHVo2vXtf
9cw7EuZbwZg9nb6ZlxNOY8vo+8Y5jn9tiBGl0DzJeio4pMbHeWUcZwaIYGIUe192EcUM1RdzCAAs
DHkhNaOc7M1/KQJbDl3L4PSe5tN0YszfCuE5tJqtvbGWH/aLz3Th6p4BMmShp8h5krHckhDVw1S+
Pev6v9PiImcycUk+74YQMroiqEDulP4JDRQZNRtjC3YssvR/M47vSoOmTtNcJyvmVj1MpgOaOUh4
IFJO7IsLpXzq2RYmHAyifc53jL/mTCdPoo8IdtRkXJ9Pwo9SlHobeKcR+S/ei05VnfHMkm6FTs4B
/PDD8AlqWiRNMVTgel49acGvRTxag//2Bm/RafwM4C1EvaKTPKmKw7VgNR8x9WO8GJJ29cTs+W40
pGaJWa+5M8q6yjrQ+PRvVhn7164w7/gchCSkp/z69WZXZCgTc+WJ1VW2nDnB/CWQNchdtUM2BHVQ
9hhk0HxaXD6ooOkN35/x1pwHfGSCX1FK6Be6TPja9PFRkLlyZlaSOn9/Z/GWYafMthsfXc+gYRMm
fGJ7XUVLdYRkdcYPag+Ed3hdUHCbqnfX9K+jTdtMLYaSGcDxzzsSV+4SvYU3THvtf5jTWFiV8gT0
YR4m+bbOujaxgaDsO9z8CPPJx1gDp0CkRCMdFLnzxQizpggI9lEZ3IbKztw8mxlMSC/pDk7Eq6Da
/rCv2DTc9nvlYA1l0/vSfRnkPCA490StBuj2P7vzg2Kk5rNCNyHS3jEUu+sIqiZV7da4AzR+ytJr
KIw1nNqkxR1QI7hXEHcDIZI/lVC0VwenFStksrV9p1SauHPJ2L7msmRDxoJX+i+Cg8FPKCOLMjUn
70eQHzN3U8T2RH0gQTSSgd2/ib06WU5MnAOY5Ow+nTZC5LXXoty01s+GquVbq93x70W2fU3AtplJ
lUPOjxg3zccRSS+jWdbJ1yGLzgIQL17wcFTuy6W6FrxgBsGtvNeIX1gRP71STidZ7lUrk6697akj
p4cpBDDKsbgc8Julztfwkb8IZH4Y+eqq7kaAVnxLlZG9xd3btfPsD0ucFJ75zhRr1mZAdkKcPhCj
XAchKFPaSz0IrVsfn8enDzLPC46aAFN7dlcx9J5ABctjuRb2wUmuQ7G7luX1JgOmkHEx5JJ7i6uG
5tIiDFkEYKh3Il6vKIOk25ShhWIeCm537MOIOVUdbbpXtDKMNAry17DjQ3rYDu1n5JFlekbxMwY0
Fb684l6xg8MStjpsExyS+IbkjqMsFMydHo2S4KKZk3JuKhl0+ZV70+J8G6by2FNfBZ8aLnizDoNd
o+XkZ+Wu+soabBhRdRSDCsNjbLnlwM1xNz469meORS5i66FMmCRrwy4qXmMs3ga7CqmhTBuHaYpo
TOo1C4ZitXcDE5CFCsrWkHxK3E7vGQob//l3n2ZMdvubOfHlj5WubQjEZlmlm2UlbVfN3ce98Ce0
rmFx2E82O3dYlbpeJewPZ9C1pUcHng9LGRkKnEVbTCckMvYUQ+5IZX+rsm/5ujyOT1NsrACS1pH8
U6DddVWrcZfmhyN8i0pJJSbnTHc6GVP13nBw4wRxGC2p31rEfw5X8GOpUBTEmiowKVzP3sps2e5A
FL5tpEFPhrjz2BofZjbI2pz0hWMgmytLN9rpH5vu0/9subN0YuiSegGcEGF0HnPwFkLl9p6B/b2b
yAkVgEcBtPp+6MMQipiDwk4PbP7ziO3Ych2TWZb7u9DVsFfKc8+1oFFnRtn5azqOewSO9kH367ip
g9EpzY7cz1wi5Xb7/zK7eY4kpE95ZBMXJxSiVyfl5PadYh8HYkLhfSiclFqDr8jjpws0ikX+Qmkx
zMSIGP8jgX/+lY8mgreLG8gmOaJ6Ca33u/loDSp8sbC7duIi/BLQHskEqAqphZhW5IwZeR0U+tYN
3GobKpF2hOi0TezASzvSgRTQLuuw7uRNE4/Artp//K8P5VFhHM725MJD29vL1laYnhXikHHDGU8K
zNaLXS5Wz4aqotL57xB/zWwGdLgRV9lVf5dcGexDUIJ/0mB01o3RWk2Kcjj2SiewWDDqWR0JU74L
5GFKsjhzU7SUSumXig9sIl0KqOHVi+ld4lb8nHSMRNmgkGA8fI7PpTwPe37Rt6Q2T/xbvQcRgQzk
Q48MzXtz0gW5MalECwxvw1AvWpaqvnDYmAhyur50aA14PzAbL1hBp1KWWiY62Vrc1eMcESrCKatZ
/RJzGEMAhsJVxkGE2ZgoAaTNqR9tK9J+dWdLyIOQw3RBclYrrX2XC8MX5J9jJ4tQfeea28QfW1lG
HULGd5B6Q1cjCbY/kz5dsdC1LR9DoJYJTe8e7ya23Xi5244rsi4pBmjhsC/ht4edSf2K2AbD1iFV
j7S3heODkGFUNRmH28mXKPab7bBvlgQ9ewwSDS5sORMSNCIc7f9U63Q8Lj3Jf/4NSKZgFDnPBcl9
BiXliUp06md9n6rfn7rCWdBJQU8Q1tlROCBYWU3HSxeLPM65KGM2rBsNhfUCWXp0dD54oA7Razjt
H6yTXjiCnL5EPU2iViofBu4Ssb93JNbifdHuGYg8GK+QZer6DMCJrQIKaK5znF3Xj1wuAd7nJvSk
72DOhsiYLuKzJzGG2AEblaiFgu0Lpx5UTOSbjYLu9wmmXhAwqwBEW7R5l/a10ZHyUluJ8jqfP+hT
wY6f+Xxye8wi+2k951KKdFbaXDaZGJbsS5FmTLs3XQAWhrr9MkKMAG00jDqBouFAZLwUIAl9sTri
1I0Bx9QIk7mIqS0xJwWTbg+YaXDkIjnuy7EzGPtMh9wzO0VZDILJdukSIPQ4YE/TKUgVqD6CZeYf
vMK/+PRbx7yHI0TX8e4M+q0J6kGBy075fUw+Ga0IwuinFiGmxpjHA6TiK7VhduEQBT1Jx4UCsdYB
f5Qz1GS5Ak2oRg01eT9/9XKGBRHGNz8esHPCaZno6OJT+EMk8PXc3+sCmIOCr9Nj6xiDoiUChe7i
YQ6a4ADsBnJUKMwbkCPxULh5nzwz9NrgAUvqffIyjzM/esLy+0H/wUcxlCgiL0eqBZ43TYA26SQ0
qLCk8uV8/1jVAC1xeYhOtGze9ikLWd0MlJB0py1xSQwLSbaDYjzGNmnszBl2Ck65YdnhgIJ/TVxF
b/9IDEB41dX2ZsEnLCW2xzxQdjbYmxglUP7C/bVpTOfG0dmOwDVetwI9my6RQO6i3bYV5ImzrGhI
CPt+nS1rueQpVtxjXn4yHxrKGwZUdF+KYz9D+gaLpCn5njPltfdBP6Y2zJSId2TM8mEE4cKq+kpz
6bqc3WcZrm4/Z1Jec1MC0M9+DTy0nG9TAfUwZO1eD7jgSitw7I/JtM8ZGx5gXi7NuAEH3TsZRJij
3h5YVk5QY32BmixHPDk5XhbMBWL2nzQtHw83WeJJ4Fq5i2RkEfKG3u81cxhu7D2bJ/eVpzTU7O9K
Kl4geTVQ92Qx7T1SsmElLFPzC0jE8pPtQ670l2Ub89L4Q7uVBlHFcagk2qI69+mOe4y8ehNEJuiu
vzK1dg3HYsXCr8QXm6SFNemNZTsHFwbS35lXIsNLBqqekctIPr7FIqcc9WyBWJXAyrse0nJJJbCT
b4jFMnwRnBiFN2sIqSxAkD8BGTEzxEt/P7oS1OXGzonq2zrNC27zJs5wzw/ryYpYMuSm2KNlliGo
xyHcZ57nq0QV9fbn2dea5LGGF+KzLqMD+eNJBaYcmVOVB1nkjJk84dm8RFAvEIk66iCT9vLCDprs
8eSDrfwArre+C8CstRcfh+f1v9UCwrCwQD5xGpRbjyJbna+YINtPI/IJbO18AeZ0lcccKAEzKLe8
xr5G4+zPlw7i0jDn9wukmnWUzghoGVREzgO7M34PnJvgoRzNKqQANlH/+PlqtY9gENzKAaEWtU9x
uPTKLVzCb5ebJKkBxn9h+tZbVFxx4FPObtDa9DAc6h2GFwLZ2Otv/gnQIXbbTAicHdlqdDeHpaKL
uuNf4tjcQXV1xXSJoJwGi9GdO3T+TQTfuODF6wtCUDRI8evCrJlYBDVHudrIuCsR2ADA3Ilp292q
epIkHO0WjX3pNWeCNN0sIuWF4u3PzRXjb3nnZBrFy3p+6g8g/QUomZolAKT5Y7j12B8L1UHfD2OL
uZFvTpDLG1igkxHwOG57IHFLLOfxl009qRljz5hn/gga6emY2kdRWUC6adirr/9IvHGFDdFDsFFs
C465JztejAWokOXtcpDQVtG4W9XvVLy/1xoodHgxO3Htohc6LuzQBW8Ih/qAF2FAZ4Y0kOdUtthZ
h8urHvOJyg5ABWmXQCDnYxpEApWlAZMEtNUeobyICoCDNCCj8VrP6gzFsjfxYQfAxNy5s+nwkrFd
DzkYmNs5rz3/IzsuJpbqSxl3r7LXDLDdGlVvOB6iK8AqPxjUSM5oKIjbBmTnz18mwf3ewCIqYo/I
fC8pNiHjAuFf9KF6XlPbZmjgtv7jC+PlHwuTZu+Rr75L0mseMSN2gp690uIMyw7Y83zrKrWfhIvs
dIO28rbaHJ4Qy4dDUS/uHPok4huh0c2Vx8wsnwtym3auWWSkjhPZE7DOu4zSrdwWYeGbioswGtMT
UxRYwcikTWsm2rcScfD9WBtlNuSfBjvw/0ogdoA9fqVf2Dh2jPfKDzEtcgdnOJYuqAokXt9vDQMX
Nbrsh7p0sYkdvZ5q/bG/qlatJ7SgGdN132EkhbVOC3YjthC5NtghwcReZQAIdTwg3mPIScT/fTlQ
22h8QL/BJKQ42UjO6bl0pHPNn0lKmZl64Lf289Irjjnj23Awb7j9oulhKjgCIQLx3aSznHU2shM7
G05ecoL2NNE/NNOy/vMFppVSAk4UEg6MGKq/Nx/5OxYMjnvev4a+LuPN4C/k8S2zzUL8D7XgTTDO
Cb22lnu8pJvsytrAcYRkBlhhXNPY9hHY0NlFA3/dkVcX0h1iD+yNg1BvCBDV0f6kFWpTyVBC+juK
MT3XCEoGQuTLApZvNjLoufMsMXSpNDWqqQDUVxebY8Ziadjl7kcjMR2Xe9aC3OfxSLErXHzm9+zu
6PcBlKCMLCmoODLEEXpJfx6wu0nSf350qPlutjoT5FRz2I+jgD6xGCdjMm+uN/2Dnw5VZ6mBSjtD
spjix3DFkrAeW4OKIkNs/3cpLOZFOdZnKubkKjJfh/IOkzfdEfxPSuF5ky1m5089sDYHmvvW2UoQ
KV2lgMV8hCZ1FstnXnWrQpLeNdGcdsM8gAFieOHH92JTydx9LJXhbcE6COa8bDkQVXZZcVLB4i0Z
Y92rxs+QJMUmfFbNRCCYx8/HX9/JjAmdCFMjo4naD7uxA5ee/LyaD/O+S5KP40H0Fw/N/rM1jVO9
F5BtqkcQ6MtwW4AnOTcutk+tseFbS91B5PwDTxove1yw4/pLkrKIGs+st4pNkb5cgSQ4854U1JGE
DQV/4GyhbDXUdPEX2wtq9/JYLFzP6Z+xPtflJRpY4AN7+dLaHcFMGg4/xfpqnGEwXLetRzVWATSt
wgufqTwLkgMB8OsGRV95zmQnDVKz4hVLGX/CZqSt/PhqzTBqPX9eIPq5z+KclhYP5O106G1m9RD9
Lrra7bFoZTji+o3YMAFcd4hyVDl6G9t4UCMkl+GZHadyO6x14+lWeBABr6r5rNX1vqoVt01jUtG+
jlHHs+6O73Hm5mUv3mUkQhVJoVwg1iVRlROjcVpHbph28/7wgSODSMP9jdPRyixuBpdiGULyHmm8
SSSqLFvyPNC6MOgt6tCy3SBsjxVPq8cAClKl9+wamp8tuvBSS+18ziI1pLYsQZHuQJzaeGlfhxis
20Ipy2yf4xto9+d2bmvXsPX94IK4lIp3RHYU/iGH4Oe+GsKWNn6MC9LW+UU3YM/A4hFcA7tIJrnu
sohgB0TV0b3Y45M7w0vM6Klqq3oBhmiJvzIp3mCbFXEdyrTrNK/5M0K4glD0losHOtlJ/2XrAJ1D
23SC6CLHwvR9ZDkrSf4lCwv36HjWqFbA5tTrMp+AVK//zPHv78YaEok3xsEbeNv/K4yDIgvIYG9t
XUu9h+hLOXZM1Zz1JHiypBtfAMFencahJC1H8fj/iCnz70VrIOOM/u2LDVFsU65VrCYd3C4v2tHI
se2dydXc5l/obQcVVNpIhhlBfnejoThnDKcJqqER3jI6b/PM5LKykjYpjcRQ4vh7cD1p+hbEdsxL
DHEGubzYrfndXFtYW+wzNXwAv5xWd0NpSC2emx0vrPiPORCOwH/la68mws6T1xesK5ezw7l2jptT
Pv7RLxpX8ToOs1QhN7ASQwwAKcXZmtatietsHCBzSHxzRDY1Jmifr6FURmJVh/oi2Jc7guimVYyn
GGVf98RkCHFf3WPtZItB77zPickNMllZfmu8AfqHTKwiNGxKoh78udmRSC1RoCqhKZyChB9XYtzl
25jX/9Pu74D6I+yE4vHqcFdU7lUL0sJLPWQK+Q3Kidz5iWK4268kj+LTnoKl8MXZeHl4S8RG2h8Z
RLb3XH+08LgXvU4jBncwEDpXA05UMSfrkwRPbOpv1LXjkWSoY9Tw1uMBSLCotC3UvdmiKN0XuISH
2ABaY6c6HC+idnDfFE9Kmn0Sr7HkXVGfwf5W/THJMtiooiW38VK2D7rJ+/SAJ+HWplzpo993wwSe
60K5PJsoGxHwpwnl2wU5JUrCuvaxWRjL9Nj5dr1kFAXcFOLgv+w3YCsJi175J7QdNEFuaSfyqBw/
WggyeHWC0ikqtwtbSqC6zkWlHWvrY+WS01lE7VJ6Pgz0j76ctixFLvwwjSflT/rBgyv32IuYqFrW
DmbeuMH2seGPspN2zmmtSP2F6UiYKO4AnIscOi+Y1Df6sO3NJy4ohQ1Ef4CMaUB502p1TCAlUejE
5enAGaVxgoGRKxpzeHUva7Vi/ClAaaQDRXhidP8JpVUx5gAVV0wJDu4Oua2nigYBkjcxdE+cMZ12
RJzxcTkbYFrgxyAS3DTqb0aWWr8gz/sYM/vk4KoHGE13x5UfyCy1/LqlCXLoWweiGdZ+0w7NHAMK
Y8XSt+sJyFqx4bU1Ygd0pxyxn4NtdIribzyspgS7cl97y+g95pRcetwmn4ozOjCNi5S7/dGzol+3
RCifopCcUKY/R2bc02bneGjD7lq+2/JhH3VKGiN1xIUuJH4aZlae6Uf+l+d4GFcr4/XWUgn9LZ7i
C8qweOYx/uZJ9L1jeBeT5F5gdJy38fXYf5JW5SVJGlK5vQI8CeMFcaOPPO66lUZHTxXVqNKA39/W
hHWarda6PkSInYWSlC8F3gk0vmbskw2TWEpsIVYdWcTtwPvRFIA0T+4abSjvk80VidFPjE5ug9KW
oRJJR2GD8wkwE/sI+4pFjE7vVvF/e/scZIsBPEUqKoADkC/mheWMWRd/hv/kbN1ZMHrNtS2qyx6K
sKuBoC15B+N8C1BQ4zxVdWFsA/Dtaqfb9JDGuprh07mtYjXRCVmFL8p54aAWCvWr/jQwDEcjauoN
/Fp8ZkDRXcwfp1ywtE3PF/OX05VzqaAb2HUtn8mqVvsfRdp0Zr3/3a8iz+ZTUW4yoFSvQemZm1f+
f7r4VrIa3Xi5ngPL+jWAGEJ8JAjPVzN6BAMbr+EDNIRAY1pThb9L/Oi3D6q4s8ZWhvzO0P4RXRaY
jHpfapklUlxNObY7ZpK/lned37xXZQK1sbE5hTW306jrtgH/cSEkSAlNR/VUuBp2Ocdry9yE8MHW
KAB6GQh4ugMObcVIoG31aX8vbLNa1p+6CialfTVHkj/XYnKJDRK4DybzhMNpx+M2jJAKJsI0uzUR
g5iHyD1HsF8QF5C9DpfIoM8KA4C87QQ/GWSCMxul55g4RJiKsw1TByJugbJMBxHzKt6rj8mTnZmB
V9keGmepgZlzOCDTOrhMK2izqh8p9GDFx/PzMleXLD63Z25IB5ki3KFnAy5i7KYIMV7iHEEC+S4S
2sQrdPxA9GCE4eJBMUAt0RBiL1mdkZYg47eIU29n+TljN0pDfRaSNSrM9/wjuwEcr9/2PS1yZbUo
iijjOAhyMbJRDjXGJV10lDh7wPUkxz1Hg4F1vVhX3aUO+VRUm9pDsK6mcx0pOLB9s3TO6EaFXdQu
IYmV/fErQAUDLTpNYe+Pn1IRufnYz8ZCV6IjKKJ8RiRE9X+9HbSnsJyykJjm2kv0CcIpr6ri3cZW
d7i9tOHONE4rUXG0GM8jANwYHSqUW2ZWU4bKZfBDdNOCJqDBpKloqy/ATxoxAp2muyddwVwTYEFy
HuJ1a1vyAH646Bauf5y8xDCcMR2jgUtqERJYVnEE883LPMvcLa9umXd+06Ux/uQica1P+Av0EAyu
ZmTYG63L2RbcGV01y8uuMHZKX3am/rC+ZmLwQohfeVyK+FKz59j/QCVuPsuaPTWKpBx0yfJsshgU
Vqo0OrIbd/DIRIPrqlI8cRlR7nOHm0gfuyksOnv4aCfA+nd+UWlq+G0UtXjv6rtLO4c4B8/1vzpS
KzMs5P7isFskOH74DGIJ99HnYU0tVdj+8LFBdp2BHlqAWZkKFZIIfNK4/4HlciyI9F3QaDxwDOSv
XgtzHv1g/KIrUTj6AUT5plze+WoPtB36fVWEwm40DhCZ9k4JuS0u0kVdPa8Z3gpSIrK0CjcdqaZD
Hh4lfC4gVFw+QGoEn6IUK+P6ajYmx5La115PdYfWA5WA8b07C+vRJu5cSb8TkjDunikQDuP9t9m4
AH6DTTP7nef0VCOxFZiDinGFaH9Pe9bx+6UpI8Gzwco0sSrYAm+40AVQefqTCseZ2+lN+HgNsZVt
axk3hxMMLZl4p40mEygaUf5poy1EWJ6jRXkZ+uJwy72CGHmalfIv4L8ajDYwdBPXCX76T7mZ5aaY
CaCnr5XxT8JSLUQCzVfUgNp1oWHzB8F6ZXEyugLRH/tA/Gi7vn7hVR/2M/t9NopbtHKmXnpHzvBb
vmbBBRFcpsx2RiGx71FZzlxtneH3je2PD0Gj2r0eFiMt2TZxSa8Ko3aAk1Ji0mbd5T1rt54BrmRS
T1VFebu/2mQBN3TVqiU0CBebaEvQv4OFS+fCSVjW/EzxI5DFpjO0wcRn5rrwQEn6DLsN4wTQyaTM
9kjxXMGfV0/SGO0YiEWVB9UjeGFsaujRINUT0ujvQQYSlp14pLt2ofCPvVfpxzGeT38OsKne8iT9
p7pXDNshYRXWH3IYxuohGhMlNMSVzuG78q3sb/kW0RKI8YXji/+9cSv3hVTt2wtLgvkbS7k13/Sy
Oisrgg+u+stXzcNzoX6hAUmaVTqkcQ3e2J8UFKtdSziKzlLExGOdP8/3+BitnsKnmzxks19nWPu6
3NTNphUH46QTFYB6qvlCpA18N0kiilEkfTOFGvFs0pIdfXfkXKczN5zK+xGnLVAHeHqS8ssa49RL
vsewG7OsV2nbsoXXSAvL52lDI8M5uLn7nJPJa20zHWvgPZRQ51z2ToD5RKdzU8+H6c0osw+lmmmb
6+5RhC5hLyKZo5YWQzKI5ci482riKZ6sUZDZs2YPaxDQNBnHj93yWptoWzcHstvjSVT+T5IeICDA
7pMNYGwYJBCzfxi5X2AD5W4QRYtVBqNFowReo42jlksX4ERKrc23iLhf3/yyma2telTqjdLqZx50
PDzfpGE7SCUWJe+rdL6wVNuqeVtKO3499teXQaYOJ+dOEqWzXZuTdyQ1aGmbM9XMzUEsiFviDC+0
CaseEJ0EAkEXpMgQSHvYHqK9uECXwavx+B37N+lUTIrBZr1BvwlR7z/vsXu6jJtHuvz/E0wb2OVK
sMOC5pX5H06tj0tZikOBGdeqcukOvWpDLROdX21qj8HPwVVgb2jflKGX69nDVHc+XkHiQ9UTQqWL
NaZ/3mlDg4YC00AHbZzZW0RTOx3qiQG2eU3UyVvXhhvICVGY/3iTtokFxD9wblGU/qh5RfklMMBU
5d9y77s1vi5B2evMLaz5zNqCIH5gByPMNH1/BIaqFFcdl9jNX8xALAQrQX1JL4ipQp5471XmKRgV
HPQ7NFoz48b2jWxXNNFgSLGali56/esdCUwFBvITuBCdP8aqt1FK8vcUvm85E2UjPXkgG7Gct1YB
/soyCZiSM1yFpHGwRpVuPm0v/1Ip/kHu51Yq9rp37DX9TnXcqPZ71dZqZ9lWj9twpyfg+W0TKKw7
gDSGVRRdQ9NGX4tVenZQ1C8sdOe3c7fANbyXu/OSjtccnn3B/Q2ouZEH71nGPi11K+qT7KiTeSsC
CC067UY6/a4rvIdOJLE3/BOoQnkCIkOurinnvdPuUJNP+cVbWVjsV51/dqeCFKrpLpLZuKwbhVWg
1WvR8fSS3J6OUVvaHNyxD06j0o4YbDKcRoHxjLEq/ktD/YoJjMhjJQUsPEq06K7sT1XnAvJ4FxZa
BPhHaFv8ZftLLSqMhPfkf/c3wk01mreH/XGLQy/tklwaDVofWcZQdlNoB22kw41xk8tnig4pCr8t
w56SQBgtuXPin35aw0V2Pg2aLeCMwi5Ru1OYqHdwKOx+qCo3xqvsK3hgRYHmZkRYC3y18+0jD+mc
9iIyy3zcWap1RV20156V0JEI9hXyGTVcdpsV5nEjnwbQDznwI6dI0OeyfmPXO6A5408g10ouucp/
n/pjHSzYFIyzm8xkDxsiR8sAzYfOwEeeM0kSw5I/KqoCMo8zmM/tmCfJIdusdCxpc4IgWDnLJzCT
m5L/8VblGBwcFsp3tcdLjCGrEm7vmPn7zui72J5O11Kg1284SmbYTk8oSq2rG4kDqBhm1rLZLBvR
VeZNalatlHgYsknHqddXUYHxWdkw0YlijmgxuKG0hsQGnJbh9ohN3OioxYs33PgQgE8j+k6f6s4D
dJfMGpFfXAY+Fnof6aIwuTJv30vgMdFSETvWuqaYHo0mewr1jfA39W0nwNavyC19ttHgjKOHXVlk
1xgr1vHYNQZymGj7ZmkTErA5mgHoWEET2kQIbQ62G7ahw7vOgKaQLmXcEH8+7OvXCgrKMEH2gTBp
knqdsqK1fn8o3deRh0oQTrOX04qCjuffGrXHjX0TztGoBzyqWHlUuLyB1FBUi73rzlkW+VCWzdz0
8gSBnPYRvpGz+G0O0d42H7lAItFUz7OQ/QRnJ9L/GNiRzOY58m4K1E4la8W+deqXjqbU2GKAvuJA
4cFHjSmAStwsbTnZA+32N9FJGL9fA4DP7J+hrGa7owxG5DnauaiI3W6WqcqCntHwc4XvSg9A6q7w
NA6gkgVooGjiQBmC8D+Myez9N9UFEusudTW5FOmGqrVag+jPEW5iJ3D2e2DcpJJTvjxJ+S1ro5Ra
AO47uvhZRvKrqCegoWAcKr9+KWc8QfuG0YHVPE3ltkcATyNWB4Zn1m8zDS91xq9YO5jQKoRSTIC7
EOW7cwoyBW1kCYSvIH4oSk77uCJ6Tr+1y5EPOvUmnGdHjBrNMe4ySa1HnLLGubLYplFlQlH3v48C
qUBIlpeXDCVWsNUo3X+j1Ao9j5rfbPmEb0yUHZopfdmNvVUXAfmcgxQ0+qEGjRfuSP3qKE7TVCrI
l4iVJAHaDOSLBFGwtGk/uQvxmJJox1UCuL+yDgl8LH1TbmxzOchuRgdaoTmxR8b4EwTzig2k1Owe
mROa61t2N2lT+x6qfQ7yhKlqKhaV4uGUh9z+h7jDx+UWKK7x7sfUtco8JB7+rt3ISF2jiTmQIaBF
wMAUqtvKOHKPNSmx7d0qS0oHWHy+9+ZgngIPAS2xlhOjHrGGVds/EUfFlyJx5DkC/pILTY0rFcg/
r1dVOXgq+bAA7KelZyd6enqJELJRfNzyJ3iB17dQ7brxu5HWv7HJMSAnntbkuBaZAbkyf3EYvmBA
a4lcIr6t3YZ/ZqC+ZHtjItfCg+8XUYlQ9yDDTvRWmtKnCGxH72S5rfES/7IR8XaY6xapedtng+0l
/Xyzfuw1o7eGYeplQAsoU+T9u8f3h4q1pfoyr39FK+2TdRnzwZGE7iELgt4BX4TMfAR2Sn1Fk9vj
JOVmwD6di2E4K8s/KDTFXIgrWrWIuavatFWwdpF9iSvBARuloocvJG+wZMu/7AHS3KxM1Tyeu2jJ
aQZS3gfzbVD9gI2X9JTrdCo3/8nVsh6DQjgE6BMi5h+0M0eP6o9idIM0gsvXbXTsJZQEc0y8EpOh
R4qbMg9ZsFJJVvs4Fj2VnNWEzJX/yYPeJucYJXl5Wdxe7CZjQaQLfLE0dWNRhLqgXe2676dSToNJ
zkh9fRJedXiGwr/VSVBcqgEPo4WFwuoOkGATxtYyqHc+TujEpVwUdH7WesELS1Vg44vgWpf90Faj
UMrU4dRxA9F3AOPxxxI0yan1t8ikhwILxjKFhK+CuF/+/xNu6txy+vXbnCABloBHPp29JRerJYIj
JBe+A1rpj3i8jO098grx/SgzgvG377Xb/euPEo1GQ3rg/PebiU9LGadnrLMNmYhZhlpUbrj9g6oY
R5x6RkvENIID4z7XYZ18CTURdXFjMoKTLH17hNbZX2Mjrxhri9M5EoJ9ffbsUYTYrTYXvfE5slKP
1EgphpOsErpenGj4S51llLjFc+8gUcDau8NjxtVTJ7kjRmK7EN+nxZmsEsSlYXITULi3rJaQAGBg
evSD2llQH6OEq7Q+rqAUiF7XNUxQBhzmkakDc9djhAR8YQyekFTww3xfgkzZ7BX4z+vKi5nwJkh2
bxzHB9hiUb2QWCezlVx/9vfV6gRGhTFC9r8+MGMy2++eV7L19apPGT7knCYSZrH99rQRADMEa+Ty
9BXTnV3qg/Cp7fJl4R7F+WdapavwdGpy7s56DKZ3AOIkGs0H2DrWfBBmAcIinU9jnKQmpgZ0QLfl
1MIcHp+3IgIXICE0JKCGO6bLYneIpH01QGabQRygD4wHFOn3dNEa3aNPjV2szZ4hQ7XJxIW6isJN
Ajg8Ws2q+OpSQFTAN4I+mladVa28FTDY4ObmEQb4KSCC788oxkavMLX+wukauvSK0IoAk4i9yWmm
D3HFTq/8DNq/FZRf7yp0qrkjig6gMrg323ECd3QksSwkYAtMFw7wrOxGV1CkooS6pDQw8ng9s0AM
M9JCgRghEGTVypJ1FHHJAZ0/QosungYqsi+xg3KrXX5SNAuZyDYAGvZL+IZkMdESqO0RGzrTPyvZ
Q2bIr+RADlNQz5c4GpLxg8QqGn0nbm53j64ixorAT9EqCuxEJlGEZMND734rqz8nBfiARLCOiU2N
rr33EOedx+TCcrJNZC60QHz1oNIhoXsQBFW/AfdfHcc6WRcdc1BVZgdOnVWBBIkem0zqmvNwRge1
qupA13DG4SLRh0dROxWSKFWLNSKL78eL2I8AaGj+Jqoa9e91dCjk7yNAVJMkbAcJw7/8r32AHW0J
DlNh7xoxGRyZNbAI3PMz5tKF/wP+6I04fJeLiykz31naO5lWmpfgjUwlsKp6qdeOxvooC5BoCSmm
VsPfgoT7/rKqaIYRWN8gJcBzCW/SsYhkoMQPt2LJbVOZocgBW6F4fnxcARwfbX/Vagnn9LeGzYDZ
DW+jWE2iDuOjufOuU6THDwp3TIZMV5RLIrtke9M0YheE80nsUU+/8bLMk3tX6+pQWt9PeJ6uOKnK
oSfS1Z0igzORuTlRMzHRG9+8W7qAcCBOHD2saj9cJGRgGK/RzzYu9kP98HDdPJPE/Hsn5ekiuUxW
g1rqSD8FHhn2dtWaula1JA2rgxfs8/Belu8PGAQPzGxwU8E3jivhHC758bPz9lHF0FeFNPT37FZ4
ydP6aovQzWbsg2U+lz4EWvoFkozhe6bEkllCfuqTg0Z+Fdy1Z1qeRner5wY1bq3PqXQA1FdIfZ28
Sra4eAG1Ee8q2svUvtNXEy+En0/RlA9LSUsz+OiGxJElzTSoPP3Ln6x/39hhpk8dvNs5X/+LEKyd
CogkAc5mWXuaETYSM8cj6Nz2+UHU6Cq9OolrXWsMa31NcAeq4yX8VwaaPG+OtbPHdVpWtPEKwn6Y
qLMGGnsk1mbheeOjbpCwqIQrVKT/ikH3xbTqGZAVl21pgg5jz2+z+kQktn5obObRLo8VYTGlWQZc
Oe1pBH9jBskgKstLo2R33v1eQ2NFW9WBj+rY0tDQubOV3fh08/rsycqM+zfSHyxKqp+SSXc1Bwo+
AMuOzvHpBsm5upsco9ihB/aY7da1Ayp+yeP5eL36jksn3BUvQqxECpjeJ/huNSuOzSifXAFII2tU
U2MQEDroN1kOC5AyM82yDiWDZXGmFWABNEvz7MFFS+qDSuu1vfsgMQ8GFBZwHnrJwdPbqkNnC4eU
gV2KWMgjTa6ZWnaS7TEG5dOnSn7EpU0WdViUJPmrc9QiFfZlnxz4IESoxvdf1atpJD003Argy+DN
Bb9h7/hiccJZPFg5yid4MqrQvugwK2W66b75ozkJd+tfGE0vlzGqCZ/Ov44o4N7i4NH2bIyy/eW4
rHS2PzNwjP5+zoge0KW0i7ixRsmgyL+WEAIdEHi85bwFCNk6sgVd9z1pVbhEeLIrce0CfJA31KEj
2JAVJilAf/JpOVxxW7pURtF4UNmXmY9QrLrvNAxGU/X1j1xG61xs1fq6kTpD/DuimkGZNsFSmsIC
sLnNRqJMBBDACoJON8wKdeNchdF8YWjKL6mOQXiOZ6N+fyP0CKFANlV/FO27skKKMoIAOTrcQxh+
kA3eOXtN2YvK7Jezjb4diS8lJjTxrelXeaTueuKI8/ciRcJ4SaG66fRBmWDHhrGpSi3hstpyxop9
u4iBBJjl1mL+B0g0n0AFHCC/WQWKnhLf4zvO4vkfs25ib97U8/n+MbBi0lSoKAusFxr8DUj5GaE7
kZcb/SrKB2ZGy19EncziV9owOaaRv6SVkKOrN48MyRXyuHbBBoivs4nUQrAQgCi5snZLdpIzSCP1
cJsPOtsKoX4JXGsOGcIP3ibwbBclM765laBoyQ7p3/GxKZrzpUyduKaMsT1i7x3lNEYvsr4LI+/g
RplakejHE+zJcwus3GRDBVv012ofHIbC6pKxAbfvKVAcV+/OtwWYtUfA2Q6LzM679yLzy4gVJ4ms
b3+eXhVPwip/eBP/AGeQHa7plLsjeMM0I7RP8dN6ENAIT1h1Qf6Z7PpdOcCN37mHnnPL3INBq1sS
21C8lQEF+ootUwgq/dzf8ynCcJq7251qs6zy7wtiGU6tGnZIjKH8aaW3rfoZljOA2bZErby9P8qp
84DLwTwHzE0T8QDvKYwhpGpnbio0dvHfdCILnQfTTI3ePEHGsvVosiJ3Q+i61j7DkfNxT0F4OOIM
D9OQ9QwBGiQpdPvgjtZFrNwf5DoWFENp4KRMmAC+BXdu05raaPq70Tc00OTfHCo6h+u0a/xhfQyw
KDUa6cQwqDZBILFnTa2g9xl29XMeL9dgGe9Ta0uurz3myxxmKwTQlZxSlptLEE0qBPZxScJRof5d
mwZs/72p21EM1aK4+wXLDEYtIkzXpniLcnghNy2MYg8/WUWjPtGfmRyJOzP5xDMvT3kcZCX4tJnq
MxDe6bWosWCkYj1XRySlf+VJV+OZZmdYL2GIj4DEddZDmi+SnzcETaPlnwRwe9RoZkLdAEs8cfxS
AUeqFUDLD3xdisoRUtOdWwi74IRJpJyF7Bt2LIcPeSUUelMxwCLGUPzwPEfITUMlu65uKz7EObm2
2TYhPB7ItlDlTUa5CHmXOiXnFljozv5lO+gtG1LRNZBvrpFYSChfkDiPJvoAjFIhG9xfoHuiclPw
IUsdxWUXaY+st6KFqtVvWfOXFdgWu/jK/V0c/Ww0lIe1Rlf3CqmyQjAz/yjT0olT8u45UZ5ECkAc
VR8sFyrsiGjoEmq35Kb5yFunvTKGWDclyBwCkEQPDex8AqEP0Uj6JmEeMmu9rW4Kpy5cVfRAMWNW
sskPbWUaMv8rRQW5GitoLup40UQiVyXsdB84pJhycmT+OLLkHOzO+Whi+Ks/C7E98npq7RL0xsfT
052Agjk6eT5A9MWCyFUM8kwbO/wkq+/Miurr8Lykk5U4xW0fXebzcONUNIhcT31by+8q62XSxo/p
BITCga0kapq6W/IAJ4KTIisZF2k/Y7rtxmd5POWbc8QlgWKuvkr/Akuka7Dy3qkyq/nqPZMtXquk
tEjoP5cglyHSKI+XeuQvBN6OiX59t2Uy99K+xzq891WQLTzjd7jc9CoR042S+mh6+XV5Vpr296bY
c1SyOLdMHw2+DoWAT5q/g6PCZ8sUcnuxCuLjHu+ROT66hW8tLcfBB9mOBNBWualc66llQ+vNOwny
2luavucRKyJyjzpDveVStyfJiVeHHtsQfBOi2uSZywm2Oi6NVSLFHKvLQ9tv3mPsAGSJ0nutPqtO
An5o0o6HFA2mAR4mguHpaWPsmjnq6k5X+/FGk4RGJQ3l1/3ts5MH81vpWJOZz1bVnqZxg5Ko4Pdy
4Xph3GAFLmNHd5QUGLS77MBQd52m94qR1v87Mk6+uykTtx9AO9YuW36DZt62xc5BadDRpJpnNf6n
EunzVjcunyR+ww7b9U7G/1Zpp9g5b11F6MP2mT4A6m4JSrKLlhwLo+VLYyuLBfORT3ZZgSSQaDpT
BNPXzvNJ0M+H07yXHpckWuumyZYWbxlKDHQufUvfAzMz9+PAPsO6THB6qVBF1cf2Yi780mTXqMH0
1MdUggtVWZGOl6jgiSWE3iQVxKyKNj3sUanVnxSKg7NcrCv2f+A+wkStUsfnz68grF8hFw1C6R9m
VWwXT75kcs1SHKlrC4SiDz/dSAEZ4RGqzXDSsB+1imFI7C7VUvFljNoeR6aVDKVsxTfOOgywTArz
ufAl5DqIKM0FSF2m7BK79b3KcWT+rvPNq/5FFqXfzJqW4PSPg8M4dwNQSsZKNhrNsZXDasOT2rKZ
IpZnCYpDxwxl/mSqmhVEtOwrZM8RyIBWWLos5oxuSKloT82Xw3TJdR4Wk+/9bbY+sOiEhlAMsmip
JaIfJ27buNlsCGh+ndgmrgZwt8mSeMXjvgzpg8VYmuc0rUZL725wAjbNaf/+VwMIMaQSGWUnIIAU
dq/wCsBEtSy7+TuSvYFxvkBhD6Abt1lUhkqwNzJfzay6TanFaNB4wpYU2meLqTZfAzpqh8vPGJsc
A+5NXT1ccV5jHIPCsep8MB9ZrjwqkYShY2EpntCbCyyI6luRj2z9fyJ/fhKL5dSDk2FhIIey55sG
AhlxEFw2UqDBId1SoVmC9Sh0QBo1wxH43peXXFg5J+dY5p6+5uxfbz86gpxlGiD0YcBzAGDebCvb
qtpwlgCwLNcSatXqslVcrvM6cWCFCfTPZHGBMB9EVaD1s+lsMoULxex7lAu+WkEkuqDhvgC3ZexO
lTqRMe8BxoueTkwEmLz+WJlM4lK5Q3ZTzu6Vg2rg6IxIUCtGb6AX4VTFS3BmST/pDLnBqzaPy7zv
knixxITkSy4u9BiPHWswICtb5imHF9Q+yVj3/7GXUuYCpQZPj6W8IQXnxb9zcqyktdr9F7mBsGR/
bpGaAfEUuwnRbj7sPtAAJaTMoLR+fwm14yr3KOvgLQQKnk85K5zVL4Ztaobmx0Yrbj2HlwRxby9G
LCPABGEIe2f2BB/7TE+2ykd8Z3EutKFD5Vibt7roLIEhdUcH/De+f9Qo/ehiTX5nwmXGLyzrDyEE
OAmTxL/hiI2XjjmwhjlVLBh9rBsy6LtU9ubogM7R9jbrYmScapVLTU4h2sG5Xs82MQ+RLLCdsTib
/4itQMM+Rr0Jd0pklJDw5SSCEBj9iX+nmoo/n9winR14WM1tambuFG1eoWZwpyWMKnGXwoYGLyJX
+1XlX2fu0z14NclYSSQQ+/YIE6q9HyUf4K20VvYALoPpOVkCk5Rafdcz49NyRg8nkjCmYokoNSYr
uOh+B4rudjRmwieHddd4LH9vR2fhgTyvUibyKP0+pHmVfMiEaTMW0KlW07wUcHZ9YhjzZN1+WBBv
wrsHVbtDR1VmDfwuLdRBEQOfS+ZPKXw/gvyuY7znhwx75Y4pr/x7/JjoWXsjTz9TwJ79dLZqX+IQ
W8P0G2Y0MLMoX5jqJJe41MfssfwU7ihaXdt7Bmns8ZmfTRRGGtEG6xaF2xLxkMb/D8BVsCWXtBCA
lUXLaiQnQs+CweiAyOcc1oNF+QxYdsUBdruwIbAt/sbG5P1PF8l6cqlqhdeq5MwpMcs0blzaNv07
3dJ8TVoNec6Vtx77Vqxp6Ey/zwvowOLFkn8faGc9lQhcWWP9kI5iUzBfCLl7FZffHSnZzIYyMS5t
o3pdW3u3xnqUr0mnAxoJbYUN5g63K1cQZSw1ropcbeCvbIYhGiT5jScFTd1fK8dmR9aJutExV8rb
bhZkNJfiNJDQKH8B0BuJ/m0SN0Da3jjZdXO8efQDKB+PNHMFtsQGCEBMCIp3ehQQ8QIZHt93oESZ
/fdXqPmklKycc0ZvUvRYucV6BIwDuys5a565LOHxksdvBcdnO7glX9ZK4eBGjsB9HB1o0IznNJTt
W9l9Rcwn7gXnpxgXwVgYsUdf9FsE5JLdezDW10kp79CBqQI3UWStf6FvV9Fn0it7QM6g2cjblEy1
qIzXGlbisyIHyEsUD31ANfiLxYa4L44JbO+T3+GGK0HA1m9TfpWwEAst8NdeJt4ZaAl/lkWbqPJd
HB74kzZFFS7ZPCMfNxTnLsX1RM1pM/ndYQn1ObsFcTM0cApZh2R2T5EUJBhEJSmSjaIKduCbaD87
8RKry0a4UJ5n15cXs/+x7zaF/SqEIS3M903y57pPLJ2nmY+bS1zK6t6mu4+qnOs3z3hLreSF5nCp
oBtMtZhPM6f5y3F1UTjp5+HDT+PT9QwVYXfncI/02oEiWlzBPf9ZiMmfwJ7hnY5cghyk+RDu7XBR
JBSaEpkNt8B2z6TtyXLdd/kuf/OlMz9Q/K5FmS8ShSV0SJ8za66ScqYO1tUf4eHMF+wot+1eMHc/
xYOBsKrzCD6DMVIf1ULM1m/JP8lnv1Io4DQpei0HtWf8I8NxW+7qfTuQebhkor/6YA4lnu63Nird
Ojy4at2OrWOvzZknGbYDSCW35UkC6layFgtu05H3OuPRaBnQ/5CkxCmZwM6zhcCipRUNdlck8SWE
pQZzvEek7doEoiLyB1EcddYscfu8EESOEWYaPexgRARJsUj5osU7XX8mxnG5xd4PTcxPwrfBptq+
vvJoNxGeWzzdDFgcXiktuumx4oKLU+38cpDHpN7+pfDFrlMxXEUSeSjDn4HR7vNkVfjgiwfeE4lA
QuDOLrNJ6qGesHCizjFlFg5NM537BOBDRxdgmdNty9eEZxTfEoj3/b4lsz1co6vBxtGSMWiii+sk
pTx3DVHHA2kZaqosj1k5YDpXn1+PtprySfGHYsArcXA2qV6mx14gBap+5nmiwjyfk0fcux9YzjbK
ozxyV6Wv3prwp7uj9kCAfZ7ogL4CpUeuoClmIXlyrl+/LioA6h/HXSjnOtFIqsH06wbPqSmsCSvV
GpNjuywH4Cg+8p7lSNDLgdesMsa8hM88cV/XvzH4CJACrsz6kzF9/7jb8XWaqqHX0FXrWdclPbu3
wz8IOPgaJNxmKbMZPqRBJgHBdi0tH95yDi/X+gl/BrnOnDMpDWNLFYYFsf/UqlBs9QQVQxHEe+tD
Gqt7/6mAuHoPdPijzqaiNSbi8NpjUeqdwnkOOAIeKl4tgBulivmzttZu0rTgZV0VCuTXlrRoauys
9wUAGLhlh369oYSFSbZH0FFAxvOmiyN2XJhHjCJ2rYGgV8Cc69jsnIQGJNr9cZQczN2bobDzPr5r
XCPYX420bXTzQQ1gBRkSGbKJdPC16gZJjeoOgPbW5tRIvv7DSu927F0/EexChqEAmYlsUUUzlU07
hFV+vP6noxceMWu+Yq6EBU8gWqIcvCZRLimXMZ1hbfE/ZfvapWu5oI62CpthTzmJgNe7t9/jklPY
9tEuXpbMyr/pfphvlhPSRDO47tpyFO4MwFux0P6AWkKHKOSXbk2Xee6SloWvlrvvxOyNOBla6Gs1
NQhttqvISkrtPAYKAnpGkCP9bQ0wd6Q0vUfwCGMuRrj/G4kMdo0fM6UHLZbiKRlXss3vW0RJvDqu
mtluAJleru/IXVVBFJnyvhma/XgNdBVrgdSPk6F74uo54I/qV0B1qBIh10wwvYFIcmfLtEVzX20v
eQHXqQYyBEFLbMuC7TAE/YogO2pnbqrv1nH2kCyT2AYZ0bQMxLAvqh4csYJxCBeugxQXD0FXKrgY
86MvS9sOy0aips9boyqwSDQAQHkn6+H8xhSP4k5raP8ldr+rJbqbNm411BVt31Bx7II4g+9Ld8h5
QyWUoP8STjU0p7hOUsLw4BQLk1V+CSBBJ7DaVqee51CUBdSOQc9qbk5GtlMDgTzoeO44Z99b6yvm
GyNpX5IJkbY8tAsYHzgPpbPvQPpiGqqB6jJzzLlgfoxZEeq9az9KrNtG+o9RWSeV/AQBhd0FUqF5
Wx3w8c1V11dCi1mlNQwnK1w3drYIiiCT5u26PCcxi0KQq0WEng32Y+y0qbuYofpoXW5a5QRtli3e
+QSV9nCd0rdF6to/H6Lnjq7WLcxCjhyuRaP4PdeOmZUDp5NXBBx/+ywM+3hKaNyWGvHAg/uXXzEk
+HvDrNFyXkHuQz9EEt76WV92PbACg+UEFDbYngD00V7HJmWJi+qSyxXIzE4IoFOm50t8zAp/wS1i
7we7Omm1gxAYfx1/9iZi6y1H79MZCUQNq3lPzQ/JAdQMMCiEyPgriBMT6KJQt/upsUQ4d9VDcpKO
DFKAeXAjiu15uEy30p77z6yhgBnrDYBd7x/VGQ1rejsvi3W0pJmQ5vTZ+noFJfu/MgsRznKcprO9
BwklXEwmeAnSMFcL+4B1PHg94sMdMIWFv11MHWw9cMSn1E+vPMQnOZrlhkeB8tbruWeaplal9BoK
Q4/yLXvjpGlE5tZzwj76R6xXOGhcsBzpUXvdBKYv/b4CZYOELzheajaDW0yJo3MkqsM29i3kvmcA
yfc1qY7u9uCPi88/eyFrfCx3FQ00A3b7BA6+HN9xIgHPqB7/aH0HedSqE44QJlLDzbBek4t1LHTC
zrgc5uOOkQeloKo2NFkp0QdsePiGkAt58BO6BaIF4I6+/59xG2N1nzIMJnEpPfsUZKCKgiV6ze6K
vSqmNDL7sR9QtGl7sWXN/ziZrhYE0X/hd6bx6yVaW4KF7RYehpwRqesCjrQMBPnnhsDUho1MCOaX
A3sRqSQ5UDdLWRhtzfbnBp/5QKsF3g57X/btqRTv9b+d396D1ElOdh1graI6SvOtsNOSdDHBmgns
7CCySTddikzjRUEvhahKy+vpuOjT1frEjZAVhomc2KfUwBiSAMvAbDKXT+yMiN0WykE6YdgBvb97
gsBapBO80vIJwA+qj9i0JS/Kcsd5r2YxDc+jge+Eh4kTNlwF8l0syG+WCJJwlVER479SLbX1VcNF
Evs4OW4lrkU0cKQEHMrTpWPcL8wYBsk8r0nxE18J+2ESE0NwcoG/2d68JgJLx4epW7MBv/XUmhIM
EpdSKnw+wB5X2vUWvtFSpvOzyj9BfazxLhY9hoVYZgQpWEdUOHAvibLmdlDZYyNzBbFYG20dX8oP
NuqSCqugr4usKv7YXKM6tqTookdPry7w45SfMe1F03OrpGTZcxQHPqIWNhgTTNKgsivhNMiyHZOq
e8MpCcSQUXKR+3Pqjd/4UiayQiLQmOAmLZYCfMGKMZ6A/Y5P022gHHs+C9iR+HB5wa9kTPDOHW7R
lPvapqNrAwpeNfOOc7oWSl2smcG5Yw9l3/OIOEV8E/TqrwUMBf+3ow6B6h5313o3PuwLYZazpuOi
9kM7Z4pLAt/uFShXub0mjV7ASFDVs0PKRnkNmzeM8RdXFnNikYQe0b7LCasP+NkcWarpxwz2ruOr
cF4Ew6LklGGYLoEf/4XiDph9BZGbEcorAGwZe0AAcnfxS8DNoV5jOQVAL81p1nVM4jZYy+dQMz3z
4hF0Sm/cyv9gL2nEsoLCrYBdLpyYbnSF1S9zmyOtHlh/kz5gdbpd3mSDuCKTqkpJwritzHH3v9pu
2kdUo0eJllEtkvniVT7x1nKvrOuu4a3w6D7KSrgXK7pos0nzR7SyQ1AhQ43sOkEYhmcZXWUnmmXT
axfOPxNfY4o3eYARwBykoz3t8vHkkj9Ykwvz0p2fZy22SF/hxFtAlDw3nWKqzmMT5CRzqc0Q6ory
JyfSpdRkqOc9oyLw7MxomSe87t33vJe75fAeTji8/VfX/jIrIyZUIY416CMlQyq7Ygg2tnDkJAB5
HVv9LZQwBSZhBlc2x5mqgEovaO6UwZfTLI5BS71IdQEb2McxxStuwrIrM9sXF6BM7Aj4+jZvZtnB
piPX4nrzgza5cJGKkWi6NsAnxMst/wOKO5ujO29jhny3SFU+O3FHm4SqkkSOCyhTfy+pW4GA0Ccc
zzPVHjHLWHQ2UyOQLjJYk3EP/Fo2LMLBAI19JQml0gPS6PNYyhVMP6LKjdhG/RFurH+5rglLkghp
IorylYb3mqR5sdLtM3kmRch9vi/ObCCf0E7LBtPiMKMCqVRM0Z4ZMlr/l26J14C/te4Sd3bqgyqK
azMed90GQJrqQ+ulE1dNqIKFxDYN++dly6jJXBno1Umiw89xe+0RrV3xaxprIKtEsS9aQE3VaFQM
7JZAU63O2OUbmytdkjl7OkPmizt1fWerrox1KBodKota9y4QnTkRbaJVfNc0Hjow7Wgtp7kLofdQ
syoA/e/Fg18snDx1zxBn1bdf5tHVTkRH4OJnFpcOLNupefclgsbf9udb9p0siMzHXdON6nudkF5z
Yb7HaU8dDW2VwX+T9LI4Qrdp04Mg4pNFldX34lc6Ht7aR1y9gBH4dQUUji1sQjFghV4aXJ6G0OCv
n10Wg5/Hw4hTwRrRnJxT5aoRG9rEjg2DssjNJNJzk9VgHDgqze0llssyx+3PHpziiPA93kefBarI
X4xfae0TYZUaeQANauZ2t3tW8ZmJq4w3PbOGL97qE9sTOGIhgF4qQP0IBRcRYktrnNekbbshfJQo
MuMyGx5CBc31/hZHf0pEpKCL8tDAr9N85/B8WFuyK35n1f4ujb0KwEu04zQpprxwbYFwj7yzxGC8
DRyYV+kr4++Ug+yjS3t8qoCwgGFWGrYb8m9zlTPo5ChOwr+0Vg0xMpOHN24AGJuRhk6CDIkAh0M8
JbY+pZdMF3vGg/io4bxslt0Nre71xSuMD4qdWSt+qYIDaWTT9cioZOeWcl6Zn4KCQOVKGyBrhejP
5i3s07IjWaD/uD8PVmFY5qCSggBTXT9fQbhDoon4IKVCQ5A6s450UkNGdEN56v1NsZG33UHU1pZU
mXyNNVjCu9zcvlk4Akt1Kx79ZU18KSjxfT2ElnUn9ALxUDpWkyHg+uF6EoNVGO7FQYjsjOeSNfxb
WjTqnGZhDm9NrM3+gEeFxkbAEghzOZuvc8tjY6O59/7+bZ0IkEkvWJYvdGrz0zJtv1AJQ6C72+cj
MqAuPUpB8skszrfLyR5PKD+5gIxZZ8kz2OxfrjUC2x1oPXc8We/cJCaSp3UliOUjV+6+fBPo7lHK
Zpitt9AZeyeWDDADTddosYRL/LqznrPW7xfOpfS80V8aEmaZelwDJk41A8NrXWNnbanrM1OEb7O4
XoFrx2czvFY/BTUcv+X3iG7RXueYgiDUCrSH9Qvz1SnQTacsms7+fO434b/DzyhB4cLlKb5QNJNc
VyHt5m+2LVkE7sG6aDchu66gVl4FywKiwxguQBnCB5PGWr4ap0VrRjCN7aSQMULAzMl89SBzZ7Ok
yMfJwp7/flZTmfhudfw15CN9sVG2c12QY9kJyVHUx3Fr7jJze/dwCC3wl3IrbJZVw+1wIWqbP+M3
8xcJysVXh6rr54szLrJ1+Nsz31pvJuv+tbe+CAemwNm3xDCmsPebNPCxk46QJPEB9qiMG27cg72T
43qu4bjvHmdv9AbVr/Cgmb6zCNpgQ3HrnkJQuoKmtxd3ACf18vPdLHFxa0Y8MNmZW1lUUsLdidmv
NtPhAR5KeUIffj4eUnBaAh88FUVHi8Hu835L/keWKhx0e0s4k2p7Batj+4D3CizriNkMf9bDf9Ts
GVT4qjJwfW5GrMVHIrhBIS5X90T0wqeiw0K9hDaVFY42wOuJW59NqUY1xOhjvSXjO+RaevQyACWr
RdogqGDf6WG224eRsjRAZ70yL82vW1APgI6/naFPW1TJu/n29khm6sYQSvBi87WbhOeMtSamfb0G
6VZwokaHTDi26PWRfdAamU4org3O0zn18B/KjKmDvlGvyrvADPMzIoCKPD2no56hnPi71+CU/VZS
EW8a8Lnz/87GAvP6WxeMw6A7hHFq9cEDAcwioydJZ7ao6O/vOX/RjvECYm51GC8OuSkAsFZOm4ba
Hvn3dN5BtlReHQ5gmqHoW4cQoLY6GHKMaiP4tjBnS/ApGsd34oveyX4hLS023UACSK0aG63vEdgK
+2IA0/lf/OO0pm76TFP4V5eFkzXr6dIvrIx3bVso6F6DHAuDQ7ng5sPBwWghwOJvlLwSuiYTRXj4
+M7bc9gDCIs8pHUsdZTzOH4Uu9EbRiwVIA7XJ4NfqlOS79GxQLSX+f4/WotTZFzt71s/84rJlZZd
wzBNjeByYG15DaPcPWe2z8bkCjBHdF/yEvZid38Yw3mFTKma2mMVmObcvUORohET8pn/TdexuSRV
9ksePe/1DaTqUZEJgzGxVfcrrbZzTpth9Rh5pg9l66B/n/uEAiqXqmSPKSsjKnXGXze5yLJpqnru
YjCiI2r6MrSOsgD7mEBxyWu1JUdLwdCV6LRdLxX9kxKROA6uBKpTUWKItqWKngdHr+tomIYQxRao
8klhyzqCyjk+dAkEOo5Swg60x80/tHftKyb1SieO/q9oqHV8e7qyfYgdq0Td7c5P2gMxb+UfL/De
y3whbUv+NbGCvSx6oWmeXL6nhQMgnYbHXYx7F6gR+WqN9B/sHqnrRrd0J8hUXK6EJNr8YFxmj/1v
VZRufWs3s+NPnwCkj1tM31qHZLdeIuOdZEO2ZGejtiqtabhj8xIEXKUrGST7Z1C13PO5LF0ctmti
QF7n6bgjuFmnQagG7uHkBAXCSOkMUiSlGC7j4OK5xkxXEvpV/mnzhefPNi0Jtcc+Sj+X4hZpFX5/
NK89OGUckh0y+o9F6myc7o3sqgrbeWLl75BCDw//SMtm3sna30S1OFWF9eFcXuHmifjp/L5+WT5l
pAIygLTgmwX7pG7aTaBD1HdxYP1r8+wmieT6gsQN+e66T2mDysWDuJAypYFp6PHLWO76tA2Tx8aA
oFRmlmB5k6lGrO+Jl6YT70fz0ZSLvckGP2sIs06e0kZkWdxGB77mjhLU/S649U8YQHEGNBxvTX1w
RE+F89Ldg0VhLdaSCkEZNATaZXOA7/0ms5o2j6EMJo+gulHf7QZJMa9J4hu0OwKlsTVsQbWzAzn/
+JQ7lrWj7THKvB8qy+UXHwJYKqv7lLlWCdqGKBNg8mHNMyM6NbxWLYiqtxRsJeb+RckRw9ECdBZs
jL/pZnTniARE+FeZh7N/WOODIp8naAhRCpCGo19/XIwPx+2kZSnQTDF/D3H3BrNViLJLODkdxoPu
nX9fJxlc0pG7kFGhER7CBu+PR8/ct98LxdHA+FKSL4tMYVELAVMZSJAU1q5LCeCbx39V0kQFdY3R
jl58AM2lhG8jj0VtLoNC5RdeC8KvY8YgMV0xSo42lgDD6gddKW8/HJ4v4sCRicKg55kpLF4Q9jX2
nR2yhUMmEU/H7PBMnPsMD8dBrPjEaZnABWv6+iEqPAaiJyIaTEr+NncP1TIZmoExOE+DhPtAGlV2
YEyzdqn/FXqjJhh2b1H5rk3n0uz2FiqCRYDWWkErhm3KbWs3Wkh43qLrWNqYwoZ9lQvvju3UA+M5
527M89ACEIfIStFCMKOIP+OmPlYIxt+vwhIJGy7UIHC7VdWYoSDfXM72rASvV0lGwJz2wsXlpgSM
iuE6jDCsjzA/+CqYZugh9PjJVAHfJShOYxRzxgq6YLq7cr9+2IKllMlHJstKSqI/nQLfwFregduQ
hBuVmq5nPaAvYJ97kJR2RPIxWbTxjvPJQt9adHYSPTObB2PKptVZMqHdJkCrAtNPZCC+c/zzj6qp
EPOL93+/8AGgmg2/mxX0WTcqS1ulQlS+l38Xcokf+pqEqtwLJZ1GkvKifxl7Lx3EMhv9jdF5Z6FF
A8IMKZLHYU84gewgXJjGgMz0kCarGZ7CvBli4lRPp4nWcP/49vm7T0Cc6bM2CfPNC725mbL3iQyz
A86kpCQFmmXw7ZTdWudVuljVM+xFa03iqVKOOenTeUNkPCQxeszHekotVR7SsM76vRg0O4lTI2Vb
Bv2gel7TOGdC9NidF+//q6PR0ma5WabBuXvHvRguN2QPv3yNS4qkGKLNN4BfZFz4ybpCjyZq1+Oz
JOVda7K8XLuybv0rrC96cbwUBz58HOI/YJGctc6isNqtVUDTEIF5S0mxQlwFjV71KE08AqkjFwAq
POrvcsqS8JA671fgyjZHu2UR577d8lmN4AIKelWpHEoa3hqx2iuCl5FO4VgU7FECbkAdjNesetrx
eeN1yA/4LPWRnKFZqpK1HVVj3xmid7bkux5pm6TojdlaXsKhpoIlWBOtrqI3fyJRklVTs80UVbFd
SNJ7lPFcsfsCGrqZmt9jqCbwL3Ul2EHeXuzscYEiDnKioqh6R6fyExcbnX8Yf42cXb3mv7qhOFnU
1TCvP0UKVwYXghZvElO1ZmXESDIRMEKWrByIm/7X/b2EhYmm3tM0AMMF1RD0iR/8CWUvyZ5rucRT
xFZ5JEC13Fl4+zvLgfdQNM6/KTMGspl/dICQuUgrXt4fT554P5ec/iVg/6F/zi1+148ysjhjAXdM
NABVZZzJWOMbuJ57lgWH6Vljra39NO5AzVfUL5L81qGfZMw3Igpx3om0KbjPtsr2GQfETxbCbBey
hVAMyehyLFdAjTYORurCv9cS0XoP+K210BlJZPWshcXyzBRwl1fLDsJYXgWtl0+P9mrVNyrpq6Tv
ZvDrHzyN6ngG2XeD1xv8pD+g+HPVWWALbgip/0dOE6ygIa+vRJS8fPnsuSG4rERi3EGG6VGhPb2w
liYCG7agp+pFwydoW/IRJZOe0erAm5O0E4YRR78IbCI/jHvQMOPeolOErOkTw8G8nRrXi++LhBzj
8XT4hEDjs7Aq5G58WMp6PSEAKwJMXOuiX2vaJQpQ+ngxR1nyD3m5hqJrkYR+sOoyHhGBN0tUE0Zq
w/7Qh6qcG16SRhSQyNZr6njLhkCaFrkLhF1LB21vC+k5BOaTGaQcEhv2Wdgjk7HD8Ry8sappXpp6
1tfLGpd8/bSyJ9r6G1+QtBLS7jD3DHFjFwuq3UmeT1ImvIuiwHBxDGQv7AmjfmiorvbGzTTj89ao
AmryM+xbBWaULtiRCBOYOm0x+AKgWNXfjW7VqxQD76F9P0Zuk9sK8riY6adS7WscShGtoAHFGyok
wQXPh6dUTXSQfDa9ZkpgpjVjrYSwA5QY1xawJteSPiUtQ4+Lb4WA6l/Q2wez+tNGjUiSoPyFS4eY
5wlvTFWZ+l9Ssgv7IX04tlhp5jLlMspgktpF0qWFk7+Vu3IbhLXLBEjHsxIzg5WCQ79TlaChb7Dk
OdRAnx3beFgyLrAipm1gCZ64sdgD7KTpmuDWBh34HSIx+cRo1NTMkNLaOeP7M0LcUE9VSfHolIXs
AQeUFySRwHRqhM0LdjBDa2reuc4a4F2Sz+hDNcGsWPQNK8fXVBTJi96iRJQVmpwqG4zqbkhTZv5s
F2TIPsIkNJRwTq5LdXyZCQ5ftPN3C9vv3PQQNv+NIxXlgGmP4gQ9Xs2tj5tg2lh52IZhjSW7AcKR
9+rvby4iEmNKZFSL0pXpvaZyOAXkiR3tbI2bZ4eaA8+YKxbi1Vv2OtLMopLwj47UXXA5kYM7t4ip
OdlhtoyCWlZ5zdx1LDKnQA8Wj4i3YCjC3NRtTlS4kDDmvfAptJ8G1qJp1aYmL9xCvb8POvjv+COR
OxH71ql5zOgZGMdlOWoLxEGmHb3zslIoU/bZXPUKvJxNrnQOzOEwYfP0ebPDtir/YJSMlnhE8bW7
XmZ2LBfqfRuR5sc+pXf/0uq8h3SexdXxLRIeH1Hm0hZpzb1leeTORXOJqqVRJ0h5jZw9YnaFWZRM
/P9RnMdbDYtgKVLyvyZLDU6vAZ+2kddE1KfNVWIxl3q47+xTe5Qsh/+gZdIcitrY7cyfI5fQxn4e
Lrj7TGlJBwcOXdhmr63j/WZvIXzmX81+/QW0hWPIqsYPjaEboZz85xHcy/Eycr9SyVmOPhqZtpYn
eNRPGvuCzm1E1Z3v86mPWfFjB9wxo4i/Nu7YuZh5acUoQTXSxiFFS5qzjvHZcvmsW27d+kbzlg16
s2Qg58ILnZMIUdsi/umuDuIfnIrC8TmepKdgTYRIClhHFjP7uZ5kULV0Xg04dXO0AOSWm6lgDiBB
L8M2WreX988/VxH5DgLgv7Rumrusso85bLgWm1ygRJ3Geo3hfK+5FdPZkviWeMIixc5wtDlJ/UM+
56Qn5pwDq0fTLjP+818ynsKan4+TO8SHzlalz6RQSt8CFtEe4lrVqb8t+rDnc+KsuO61OnO5fFnG
9P+M5/lX6O7zTfSZz61VfV3FBHSCJwZ09D2FOS0MFc8r9rXibmqfzw7kyTdvH/3c27Ue0xHR3JQZ
CxWBeRqniDv3zUIKatrYinQHyRV//3P92shpuvhq2qrHcwgFOEFfQ3/vw4IX+ZwaKaCZmBPIcSn0
8QGQt0mKf8J3yxzil1VgnwGrtboT36QgP7GvjF0ekJZvwlBcrvcLwBPdE8djK4n6N3AeY4+HDEcy
mGR5iVgv7QswQ435b6myqPmqCEeHvwB7uS9OftblVsTY2JfJDBGIxHoOYOrn5uQEHOV8NSpAsl0b
xRAvefZyWz/r6oi4/VX8k5a4mx5MF8MfpXaAeaF27z2qAV4raN8kuVEpjpmJDsD8CPnx+JJVkxrH
FrXLQs67R8OAYjzDXEWoPKqW5EEpe50/tsRe3I5blQZFOR0+UuSnTnbKHQQhikNQNqs+R6Zaz1vO
gjkuv4jUiVkVe3sLpW6EZohdYpQqaB2emKM+42Lr8hz91eIHxYQoGdsiBoGcdwY1gQXYd8d9npTG
gdS8/V223YmTimPyLawf2dYm1Ue4QFvr6+AIO0RyhO2foQKJlVOwUzPn/j8mv1tRmPmDLlNy/90U
RFjRbczJIVE7S2w90z91CcM3Px7R3FPJixnTH+B71v+W1cuoTodNud2fY6iDole9pBxVs9NI5nH7
/WBcVbhvdBDUz3nE0JOmrDADFFDJu+gqnQTjt1VqQP+Bqp0FHb2maeYRsO2faXzfyyrjuTcfKrsh
xeBLlUl86dmZvSN1E761Y/s9SA47jtgadEd1bWLB0iLhL5j3ku4F2p7NJGCjFX2sD1Y5b48w1vXz
zC28eNXrom1iPJ5IQUS0Aowjatxp4Z9SPNk1rTpnXxd4X8LyT/PPbAszmVDTWuRruDQtf3DIhx/v
Z63yNa6bDpfJlzmRk6Yga5e3fiQFLuwEOHLBB+nIQQ4EgYSsCSdFcLfiOZ7+glCDPScdcu4L7Lev
sXjjlgY7eBnHrbOJR7ma5U7iKfhAw49ExvcHgH1Uvgs6FTcY/BsPC83+MG9bpdbIEzkAWZbEajAL
jjjSqn1J/aYrBbudyMuLH8LR7el1DcMuWYfKZJvUbXJvhgWAa7tS8uyc2XadI0A6qOQKuW+Huhwn
ZKU6FsFRdRaS22k2e1m08P4fX5ITIQc5bS1l6hvk0wH+RT27hq5yuVi2h1tajYtJuzZyqFwNmPIa
/FGmBXehwG+13BSHvfyj3YxGjKY6arJxPztbrM20l8UkAn9as3Pp0ZIkprWQdHYLJov1PcIstSU1
Bc07YjEDq+Su33zz45BgvFpnM4LYdXDEknE89ecFW52TOwB29NItxFg/IMpQJ3r70J3uydRGSTlK
uw1DZNIz1fJff+K4cu5L/UaL7wcEaOypeCacxa2ywZ8hW7xL2zB7UkNuP6w4n+9Kka0XHF1/xC2k
1nWHL5+kzcJBLTLVP3y4/pysOxIx2omSv6KA7WuA8VzJABSi27POufu44iIqXx3wth4yJkf+D6zk
ULbJhWREgH0n02RYS5yPRY2r/0fEQZ/Zlvncfu4J7u2ZUc++B6R0AS4if6NX5x7O7CAOFaU+nFKz
VLIthSO4pTraf65U+ZDtK0txeI34oQSDssM6a0p220yD5pQ1BPTdNIptpvTopF8NxtMm2MblUPNq
dkMRAZRDU7ZchDETFT7VhzCLTtAXijT3tSLMOD8i1KISm6ae3P9t8ia6MJx32MedS7K22PJpkO5g
ibs507iv2R3bi/veNuZ54B07XVpuFUnfkZsf33isf8IafyWskiqBairpH7N/dnTCjHV3PrjJlnyd
M5GQ1Gk1u2oVqeEHqUrBU+MNuWojc8uOVQgDTN368LGLESX7Ad5fNsvom98GdYrB5k7aCZEB15Vf
pOnfXW7Ze1TNPL3JoImtz3Abw+iNUSmr9tPrpOg/PPYQbTQ7IltlCc06hoCKBmyeyCGJgK3T1uVc
Jkes9e3B3HBc/bDL8+R7n1GQVamXzYDtTTGrjoR+KumIoGRvnfLeKxAnf+6IP8/yOVHNk37uW2zy
ffRvcHfGJ7mpGcXNl3Y0odlHkGyYZvDC/OHoBjDXEVUgCUI50CSRZIyz7PWN6RZqcT8YjubnHMzD
OzAP23imSA3bdbgFUsG568jVpFy09uLJclZSyyuANzf4+bkLjARw4hWK6fhd4WJk4SBTdTpc3EQ1
PG50whZfPRaaOeLbUGByAk5xx+vnDfPsGJLiAGW7umLYmbdYwPZ1651AQ4V44eoPK0nhWLAFk84E
RonljSoHLfCf453PP8FdXpl+kEGa2bK4omP2YFuSBxdGTFOSZpka37TpGUygf3wlKNrCngDjFLco
abmX4+/eFqlnAoYTbkVQHk2ZXuzk1YhVG1pIs78fvb1odRl5GZT5p+lqVTtdH18SsbciAP2ktxLa
iFS7U1/PyWPTD+Hu5G41X7LusVax9IotmmFcMdhWb2KrlhWLHC9C9591wXxgwrGgkZJ9DwndrZUQ
KgYUyLVO2BxdoDS5UUB/Nlw9Lw8EKW2gmcgbnNZT2ecUjz9d4ARQiePxUWNwZY7sDgc2+mRaV+O0
lZUSS0+MH1G5UWtZml18dzzghHvT59LEZKojzkRiADvrA/8Z0xrFXgXDLk3WUuT/C2e3s7P5CX6j
DXXiBuLrUPb0kIZxBVg6LLvVrkvgGpFeBNnKsx9CguTbDHgTMuIdbpeYt3HMDLOzwrQJ5e5zlXUi
NykTnC3j9+hPF2JA1AkzpA5b2JBI6UM0euPQ+0mg7MWbuJARniyM1zwPhklIywBpTZ49RQKGDZ7t
YB5K2DfEiZvHzq6LCHWK/RXOtevgcvg0hoMu/iM3GMHYrL2ZT5LD/NxWIBuFEYK5Gx4R0Q0H0WIJ
hmONVCIvg2TuaBtyg9wYP6+YxqnXDf3k14ew/FvcKrgRTGHTfa4DfnjCR8SQ3mEKZwFzG+o6bKk/
75j6rqyvU9cWjnDkBBNxeQpkOhcb7uYKk0Fjpw0JpCN1R93AcWCYmFjsURfxkmvk9O4tT2SMWZIq
JWFktqQbM/8pP005qAuHepd7ee98cKAzEHIo+rA56TfSXl+hRLyAEhlAr1fI1ijdpqueecCYmvHB
WzxlycHl8DXw/1dzGpoId6nYeQ7OJsyPIxkcqNKfn6P6EqcYCsXf+KW3Am4qpPCRI+MqSB+uFKzo
c8WQqsVtbfg9NBKEGxOhW/dLUf4byFAUHnMos0vMaB6w/DnNSC+8+o8NjTTcHhPezUdHHEbxdReI
eQ8JXcMXaf29lYlq1f0nBd9zSljXb9j0TIvthX/3DJmXG7JUdLTKmnvjf4MiVPW3sEoNe1mF8XFw
L6ycDQdfKvK5TVvTCyGQ6anmvVfEFSr3UudM0HlRwHJ+aWCoXf0fNJLudWjKHLOuyBqNWXapx+Yz
h8f+Uu/ibzBKgrAEkTL2XwMgYpImzR30A7Sa0JJ83ut6xzK8pLq5sDqP9NC6Ki0Aacw6kZQlNoKe
YioyGO1BRv+H8eknGwHr8zcSGhisgXf/4NOiAjBdYRBfi8U+7Q1nF77lTV7r0l0n4fEX7cboJQNi
TNQxUExcufg6+mdNzpKDQiH95Jn94aeJgK0VD5acM72KoV+JfHl0zQqk7e/bIpQBmRXnkjiSx5CQ
MPHkwBu7JRu+SGrxtsYzFFAgnuOEHjx59pYV0BN+OIKFq0/An3xwkzPj+C95IXHeDrm88hgPvp0J
5b1GvV6arJgx8K0w5iaFkrD182u+3coIv00YQ7u7HwFd9v6jZxDjDBjfGlUCCy/RD1RlTwek8vOY
X5X5bHmJIRbzXGncO+OrOd04yWUgG/w06/RJE3BAKpIXMygW+hJBU6NGN59+hRWD2Xc5/2EESYOl
k1Za1Li9YgjIRstBRQpdr4sPQABz9P7abRsOXZQ35sxnp5uaPT3i6VFbMKZSSfC00Q5IWuU1aMP7
GADoT9bG9WTAxjpmyvSvEzRh5kNW++Y7siKHGxRF1j1awvk5mBMjmfEFF85lBbAHX1cH5VjfQNtE
45QZXiQrBCxxKZst8aCZBsCPb7FGv8w69pkz5YyeVnjwfHQ94dLELWfjyz286hSqjxJ6mGAa8DOR
G4vRrDYki0sw/ms1jMw+bIUs4MGh9Q9wuUMd3YdgXb0eHZRmKDOx1xfG6hQepoQI056yklgC2kX5
v55ud7g2nMubq30n8LS0WHXLQuUfOl8ZpgtSy2hqNgpYl1qjpcU9FdRypHS/tDLS9EmXuTUxdeZp
GalLl61MuCVVCpLj5yWsPUIMigdQKS70lIciVvwDbeCcZkXsBA8l5UMFU2EpE8uCHO+4XPtqRYtN
AnWPeJ11FToNakotjusdHB49hcrftvBmEc0wOlf9dcvHXG+WuzOi+YK+FIEoM3dEzg0WoOKUHpCG
Dg8xQGCKk5ZEcUk+sGSUfdtQUJVFTgr06cmuCYr8CWXABsBISZYiOyqYzLlaHA/kEA621A5TlJoV
cT9iMr6nw9jzWB04lYOmTsw6L1MX3arJ4zZF7fo4CMBh2VFWM/UWpuWPcFKxcd5ebWBaJY+Wmm3c
iuUPCmS3wiUTiraXbJnZnD74of/EA0O5/MWTYkEaeo//P6bfsCW1yGUIHxGY+oQv+4Z8Cln5ATnk
n6Xwe5S6hZyoNnsgXc7L0S8RwZUbNzSaO2UtGuBqR5NdmCbMzDEyAx29SP8QRm9kLeLSnPHr7kz6
eGFxhxflRJ165Ie5aCmhkoHYeaWuNW7gDxkGLJNCUYSNONdID0bAizM7nConofr63yxbIkYefFPM
XJGgfeAl4rxMTcEsxSg4mjpZhy1hL1XNpHPlNXP55k6p5h7Azg9wTt8AfSilcSHc8efOqRI+FT9j
iIVYFslaGKg1wmYpSQBQVSot1991v1bqwVT7PZZzHMHLgEw5flu7vL2IdwzbxE4pP+pX+3H8xX+C
o9nE/0Y0R/qzCBz2rrRll8o+NnBQkoWg4LxVjSxZRBm/rcj8zXVGoaqOddesjc6E35UubrPCBMMg
6WaDmzuvpKYSGORdY4lEGtpp8IR0K+46kNX5+sD2AbZORpObBBPxBfw7C3/dN8tIv8QTSHyAhlkp
iOmZlXP4tW7ZPZXR9Mxf2O3q4mTWhAmyQyPXZbJnGI+jVGJ12+b2txd0ccBPbm1ThU+8kpcGB5G9
7H95fQ2weeQX+/Pe3mz+3tK2SKqDNLGIa3lwJ9Tu5T2QZoQr6ZxEwq/v0rAXM3QiHJ402Reoh+45
6vSjc8ra0UWGv2tdbJ/iTW2GJaq39crjgnyCwjfxb8sjtpahAPxahF0OE7dcG49X92+HteJLCp+J
kqLR8RNqfwrj8Ja2E86xNVg8CFNvWeYT13wcGiUl2j0eZ4RzhhvM61wQ4k4QTvpe7s2FkfwPlQyz
QnuF9uh0Uo22ZIoWK5gZ8UkJDK5e4Ykq4Bl3xS5fPw5ZmDQyrvL8r9sQ8/2YXSbZuA2v7uO6MZYZ
GfLfbUoBIkkx4D3RE9Rlem77gzkELNmjjaVZLKerL7EDRAnqXuN8D/S32FO4bAr7BIm/txnP5v9p
X0xXeZxI6gieTNbe2bPeysYGQk3NgLskXlf9fpLcZkZN1/touFsv63Of1SM+WWglrl8IFbgPxd2b
IxtaIDDKz5mcxVh+UwdfyDh24WVbnpAJNYGSYIsRIXyN2WbnCJWYo/x8+IuGf6JrUpApR0onvB8W
uiSuOyELH2BUuB6P23ra0h1YnJ5b1AwazkjR8uUkt/3K+p6nDzJSko8ua5YbN2Ye02OUalmcoGpF
P8D3vUMvcFKaRO5YmmN6FocvE56msqwLWDtatJJHMPeSvGu3iOPameyjH8/c5cn4jn1el3oNClrq
te7OTsQ6vpR0TCuJX7ChYDiz3/+TTmUj+38T86NhCGBWe7c6A2ywP/9OjwCfnnOSC5SU+onE528n
kSCRq7yf0avHw2zbT05K31eQL43MOIMllbj84tjGgEktdSPCuP+3kcF4fzop+7zg/6zBbybpVofv
Il70SA1x/4NP+pePTxY3h3UGI6fOknFgqxasKgI071wVHWSaL8Kh6vRky8eASd9ordXgbPigSi1/
9MoPpbPHG2sZ+Lj0ziI43rOkKqxHiWNq953+CDGXg3ebgol/jUQ+hIzZBzyRwBgNMoeKaQ7/kKGT
AxutoI6wIfa2NIGn/vFE2PX87WtegveXjYxd0WInDGR1NAphiI7+qvM7Ct09Tbx7qH/aXJOzxJIn
BKjwzNSbelS5xOshaV3wGwdZ4NlnmQDQGeEaXI0KDhjN5/Ae1VqFWHjguBTDxAs0nZKyI26Wjage
rCgjdWOEK4glxBz3YxqC2AeZQY5sFfUjuNtYtU0rnPaYYDq9Yk2X4fa1M3eOt5kMXBUQj0AMiKE6
ksUGT+q5+z/1qZ3bKU22UTXle2LGifB8H1gNMkMs087HRZX7m9Rq0qS8TRIFOMHPyf1uo1kdStyS
MedDIrFOXpCNP5r9tUNOKdNHRIt235uNwprmAJC6epRN+PWQ0eVDq8QjfVvy1M2pbSBeRAdwVjzA
E4/ofkfkzAj1/5a74fdI4ZdEoHgCygc9tbUA5UpyNPpw7/KjCIEz+vF+Vc2wutZ6mjS5MecWnaL1
266YwGAQ4rvZ0QcbtKPFg5xwvioyQhipd/2NPmjKNfWVcYJuK26KStH1XQkxVQv3FOseF3tK1afX
gTP8CpBdkI/9SiKy+CKx6SKVfwU9/zk8cIY6ceyLqNMTKb6xnCQpLYzLcweSfHX3m02TqFwnua6m
QPewQDOU0VaT0uuqAJPs9ced6oWyjmx+kbIIU5Ygr69n8w3We0Wkyhz23jUPupf0NHNRmJuQjqIA
WpF/t/O/rmbBPIXQsEqdRUFNkLK/s+l5TJB45VsPJlXYaO/FRQccicF22y12gfPVC63k+s+fvNXe
8IvDJrg/4gyKcXSQsCzDi3pT+nkUzptMpc8YwZlSmdVlgoW4xp7RzavsQg0HfR/jd7c1DPgSEx/z
JV/vJyuBsQAmqRgHAQorFoty1ITlM9Cz35r/Neaf1VHA02N5/YbXosgAbqwqf70YgKRg/FGb2Ihi
/1v/40QWjGONcuecUmK2vwz312GuWfIIlfXLTxmzUi6Ydk15ARkYc3PxIsgG/9qUqcG8xsqtEyjK
SFzvHFp3cEg0/2PLIQ1BU67GVcIlirkU0DLk5CZ37otPRiWfjN0WBriOomk9+ipqZGXTK7BVoXlg
eMNgtC1V8ySMD9VNqullhxSQndH7dPOJSAmGRAeuKdNP+p44y/qWG9WC1K7gTE3ltof6N88AhTAn
4LUxfORc8E6qalX6+aHR5PXIybzUQMioV+riyT6DGxoea4YmMz+MIlT2xKaPne5KkfetDzWvqKlK
EQ6i4c9I7ATRplwShn986D2jhGISFnH/SjqiWzuaUgBD7I5yBWCDJrk1dFSBCAXRdxC2l6E27FHl
vhOqj+IaqMhgP1ZLErai7viVFSyiiKwHph3uraUellSIFXeOdUvk/A+f27ujKVWoE2sHEpGvbcRb
cxYsyR4wHdq7r7y16c15tgfdWnBlqes2BVKJzO2TFd7cypZkjIIE8ZIcl0Z3Wr3E23dG7N4kIz0M
ZfBqygUPQ/JmA5IdcNhftqj9wgqcWiIBxUMMcziBnawXFcq82bGa7U2kFBGla22N3QUUR6bqeqdn
iM+yNrfXloRDNd9rxfnaCidDBHXkSeIGjRzO8NTKoFIXKgky9WztWwHjjGZQ/1D9bBnFc/mMs6Sj
YvjHpqbeC0xSHWnGsYv8veZpYDj3yvDotTUxeV6v6JgcH2Xgq0zXv2xryBhtTv2In7obx6vt97Cc
UhQB3eitVwRGDYcdHaNuQx+JXSLSympD7A/Yf4sFTBqSk0TWe+4ncdXFFLAfHaiju0+i//O1c9h7
xW5pPvJdfTzwlL7SrVDLltRuHsHu8310bICGknPIQixdV5BZocA/pdKJsnKGGMzeO0nO6brk3rji
5C2BKauFNwgxcRBm18sUQ9WefAf1T1CTkKpI89txcWUUUYo20a/EoLQVhf4l1GNcwLNLstvesDN0
d3R8Nb5rdsFso8ctjHW6ImvFucFQefSM3TFbjhSilqfbKy/QqpGUydPLvL8/+4fDih0PhSIAFnCR
fN7xDg4A88eVIsX83tqUS9DaVSEeS2ObYF0PAA8oT3n1Yz6glvns8Zc5GxmPDyPEYCssPGa7kc9I
McRHvZcsJmwS2WYHDxzMBBlI3iu0CQcg62E79PKY1sRcORZKZQc1PunGXZX6DJZ3LP/mt1k21ovs
lId3JNTNr28WP69PDn2BThlYEO2ThgyG6+T2lUm/x3sTYnReYvIHDnVjtyeYibwSVVrfEfGhTWdy
8IqTIWzchj1LbDpcfz3QrY+GM2rO649zAN4Cqy0Hma5sM3wGScfEvg1bnPpZlYZ1alBS8+OrQ0bF
9CG56AZN+QUfs3bvsYzvM12J0EbTxBfFnnOpI5EzQvRWGTplSEx4UNhlhxFxdVtZPgnLI5Hl2OvU
7Xmzs17eEX7R05AC+iblH2VuaUI8XkA6OTqmi5ov4RvVtF1GUBgkWc+0YxFBWh1jHPG00Im3IESp
mdg7PisdMsAwhGp9fY4dl0UBCJBz2pOhoVKep1qpl0smB3V1yD8bDA2k56HjHoPiAkR9LuMx3904
ZcYa4vAC+JAF+csul9V5xAWlEZc+h6erkM0tIyhsEcat5oQQKu5rf4Nutd2XmVAKXc0MBe8u8RHw
2sOeTlDBwvrVDbJkcmI6A7X09r5nTMDuLzcDI0JN8cON4W2uV0Z0G6jK5FL3awS7S5GmSt1VNaoJ
5as5QHTu7JWTWq82XrEdHMuykWwn2qXgDo+7rU+nQ7pJNCj5obqUX7BhkxyWLoZczqdaBz1Uq60O
ujFeeWdtZyUtbdDTFNsahWcUEIR4qmbmyHWrdAClkFfI4PaBTBSh3aKZ0oOpJnTXdnYLwZy9BzxG
2wRT1ksaLHy1p/fUW4EwZi942t8me1qWKztwlTntTytue9Bqbrx5D2zNnFrkKCkbI7mEQpwftOeN
3qFtFQGyH9pRv9cPXt+qC+ZiaXXf9Rechf+YIoD0eTwa28lTV43EwCVk7PWSkHX8hf18xEJfSo1q
IqP4I3L7L32DhFNMU2N6m94lruPuJQOAqrKv2QoofJ13/n8KnfL80EClZyzmmYY85mfcwuzZdBye
QceNE7tJpAjjFzKHL5GnMXMxoN1qBeX7/kU7oFOfRRHCTZLm/XnVhSmsKEQ8Kq8NDOpJgvYo4yK3
umx8YSF+DY/pBD0WMg3ZFlB6yXD1qxvj13ff55ESJi6N5F6yffPJEiqK00Yu4c30WuXrnzGCILuj
gMULOaQz9UUA3C197l7yPNyEK6EBmQ8I0XLbmFb/AZKKTEpfo8/NEQPJK2uiwzDcTh3GG5bFY3rq
zHUQQ6NIQ8+0RfTuFywdvZJHYZV4sPVP977/ipdB4bLyK+YXzhgfRnEnrUXetTj8BPj0HfW4tSQT
WRD6QIshphEGp16n+TAjVMwaombsb9MhCIlMDS3+IjvvungFe1i0zOmgx9y0RDYmFYkhjSjGY4od
kgCBgEfdSh0Ss8YS07TkpaZTT5rPc4x1t93w96tAjuXP0771GVpi938NoSyaAkBgoaSO4gqM6beA
KqUpPyTkN73zXBy04mz3ht8/cpHF1vqjya8Ca7zavVrzMHobGJbZ0IGno8Dbalx4GdFQEc1bDD9h
xcn4FNtJchGfBeDp2dt9yRPh9Nnv2KBVmToDmFC1hxnYMq9Pc6nkbBMPxrCXj/QC6no69ozwUYjY
fT+qqryAjJ3z9XanuOg/uBFx48VWrrOklHBt1EDU5/rRCBaOVNi+WeMMSmBNij6azAk2VHHcW1Q/
t9emCPgnYZ4f/2l0AR1sEmUO7CRKjZdjFXQk2flGmYyaDM+WIWY/lfRKyCyd2OIQgRfdVF1UkRz7
bQdZj4ov5tIPtenLY8cv41+lkdAIg8FHaHj6h5ov+tBCgesW24M31qkp+er1h3KEd5hy3kHtQyFw
aVfpjbkS41h29fIrmIs8K4LhcESs1U0YZ0gQFgwGVrL0FdP5VOTKdysoSHjhvStEQGxt6GxgsjVr
AJP9w6FCQZPD/HASqRAPoqJIJOf8rdMOwBKZXLNIIKiAPFDRYKAYMWJ9nh0cBuNUP+sBeZ4N+nlB
Potdy+cP31ANJBRyemuZZr0kKPPRfkk8fgnhYBn3MaCHgDk752OvEYZMRSJlvd8Ucohvo8OY2/AV
tX75LvdNaOL+l92lWi13yb4MU3d44ejVA4DMjG/88AK89MBpZrKsB2irgIMYPGFUOGQFBMt+Ke2I
R6F1fE9yW4XV4bwiEN8F4ZXoQlytehkH2JzszzR6yEG5X6w3nOZgrCV2umPGo7sjimou0qBp/ZRN
bzy/Ul2aI8Yn9qyGikjTjXPV4ChbyT4ZwXQgZnlwovZEVNxE1K4uc09vrYbb7f/fVU5dfj0jsqiT
ZhN5jvZIzJ8KgmwHOhm6zcQWYNGNXH7UiK/354FRjZrgLBMPFu5tXS4A+jGavveo2L9xn6jEExRI
PrHTyYDv49nvOm8C/vsZaj7dCDJvfP9egWo18lnD2rBvsjBfGZ+/GIXC0xhmTDYgSNhx29cvUUQx
qLlL/PiAxfAdPLhVo8uj/XL7Q3mwk4en/3xIzVzxS+4JqQBJq7D47QChmtjca+NZNg3AEhfBCZvC
EFJsjr/6k68rf1UNowM68mIFUiaKY232UT3ukkhSalIqmGKthxS2b2zJdPjqdtaswlpUwU+fvp6z
8UP79Xwc2DcoIIzqSJpNULNw08eV0NraM4Pyt7MGiGg0Mcc8lx9eeKEfQvu6CUewVMTKPcJ2lXKD
WtqCfA5AAIgRYUrpO35Fac/THQWMNat/4s6m12gYoeIMsXFkr2ItFElbRihl+UfKDtZpJMAC0dia
mm4WOqXbERh+dBjgSFM4XKx3nzmXs0W8IYDnz0TqwHCfG8XJX/B+OVEJKKfWgkLgH76EDSq6wp9f
A34nZTyA87ujtULIYU/W8RfxMowx7eMHsQ2O6b9UmJp8eI7G1hZjoYtMQ05elEPbWqShZD1zisXi
zRPLNNF7D6u4hQYa/Ge8FhV/Mz45A13EJYiQv4xm6Qz10opKokIIH7GLZfeCJXzchkWYIjLb+FLV
kSoM3vHPnhKrto3x2zkdEVHvsFG0JVftuYJDBTxxW6E01wHTRSBfhzl65NNfs6PFS8/z4VP2Xvvn
l1+SmurcmuQRA5l0iOTPhaar38hjfe82U5G2opWKx3t7kk8c9+9DcvDrJ0hJtw3439BUaxy2qUNV
uk8miUTATMfoEW2mwosml79EsuV3xSRxUedMnjX/BDAjbAwVGyPvQRwUArpqMsL3HBrEF2PACVbb
FaWPQ4s2jhJXXqIZdXyBP99ExjR7FNitN9F1wOJdPohE2h9iJZ7VW2TN3iy/3IUsPg4qAykS41Py
8YXEdWh7AAM1q628nZ677L2ZrDDnZe/aBvc7nGzrJGL5cTez1ZzCc93zCQOE90myM2dpZ2h6eHLf
ZHDnTf3JVL8Jl7xQEPr6TTfiHzhCmkwwRga+sA97yHPz2IRhqmTTaphwybjqPkGGbCkrbZHPT0oy
CuctYg6/LYkVD+yMIoTC73bOfEvO+epc1nexue9Km39+7jgDQoc+iBQF6bc4behvYWQefhdRE+mA
a8kf8SR62i3R4OZfd2qjyOQy45rySs0q5oVgjC68xbTtIEWzYAO6L2i6Kma80u5Wi5hTcT8cD8pz
TP7sdw2p80m+8ZafHYeBi96cgvupLhZRgsVdUARvPY3JRT5CTv/cRUrWdJiEb6cb7+Z+OUMZBLiI
okJg+uOahnVW7lIlGdxSHpCAZEqbBW978QIcRRNiXBCTWor38BeqOfXEe8VOW1iMbtfsPChcXRjD
PEjGmoLZ+DblfZtAIq2kOxcACSBzgRtVEMhI1diefYnIZ1qP82tvEPhqrEXDXMENEHcdm5veeWk0
U2sJ07iMP88eV2g8KozdzDbHuMrD5QpCbC25R75Obu/SFpvpyZDCjHZKUEVhHagXJ3PrNNUniHbN
43dwxAEz7Z7EwjXB2ctitv5KB7FWCS2LDRnnuNAXTVdqPCLy80otQnS1STEb0q9xeYa9qHysuHuc
fz/4tAbJV2lPdeMUJLqhAZdHbpcEFYAVqdvkrrlQVXHn4bSODcVCeqR/+haPBBjuHmrJk/LUNL79
RNFK6O0qCJbWzRlmAch4d2Bi972ze9ouzpzWcVClFZdasYqq9+/qQKk3ONP0l1jx79SB2y9nVqGc
FZnyfal+u2idgxy8jyg51Y3bRmnVmT5FH/dzayd9W7PWPEjvgPyytolL5qrVxJ2MZtux6NW4h2xT
cNvD/v2nIRE4SbEEpj2ZYd7zoid3a7P41cGe5gV8gpRmwVQQsV4vcxmJX+VCikhk/sirY3cb2IWJ
pSW8/BbKtGotPQwT9nrPDmWie4H9lZwbTdoxJfF3KQdwSDuFMKA88UxBm3Ir6y4cDjFqL1goCZCY
EiwQefl5o5d61SVRvvkJdOKLXRpHnImNIM8w0DzaloaxxLV1Y78wdoogn0EZLW82bMIKnNdX9wsN
7DWcjackYyYYm98IDWdJgeTkbWHa0qclBkI/W2QDXvRR9svHJo+Qfuf9KWAydQsKuVsyYgibJRGp
IXI0KIYDFEcta+lFbfbcViOM696EQAPhANefeC5Sis9SeGupiiU8GdDWEucuUy2xP+B+rCoImpX7
aPvnOspUC9yR6A78iAMUEItHUGk1K8PkJEQhMa5O4xEEpzMYTPZiaqhmLAT736rTzjoSKZOSrFFp
9j8s4yW3e2hDMQQQ5Q7Sny0X8bJJAM6Lp1xWTDoOM01V/TMuI77cehQgs5OfU2IeswWbtzuGkvnN
jZdOAVj4QSbBaMV9Lv5Y8YPtXv5WbxYaA9ewfWESWTZfCqSMSnRlDeLmSQQeTb8L4BSE194HX4p+
aW4w5bYNXoyaV9zJ/7ZwErNI+cL8oXdrARPP8aKk9aFoNtqo2COEOs3il/XaJ8+mVxQZCOfmfY/5
VmSQ5tWaHIIESDgyXJtW+wiz0FK6QUDVaKHagELHXsPvsZ8siC6ZTmqLI1vQmYtRtmIec2RLofDP
8QIjI3btwQn8pR5ywTEmyb0l+clAu7r3p8etLhnq37eH51EDVdxDV/BbImWs3Mh6RtDh9zWuS9Ab
A03mtXCz7TQM1GFJqTHLAso1kFFVU1RSXNX5gZ+Rv2SUUI+xSwlHFdw38VZYOjxZgkSZHRMUvZJC
L9rBhsxLBuAPY7c1UmJYpBLEuoBX4WAsiXZTLkYRCm5HZHux+qGSRUWPMxjXPrCuVu0P8zQbnZNg
6R/aGEbMco0mkyATGM35y4TAiQIHogtCrlMsTZy6mFVxw08oz/6ntByez5FtkQV14FVKdg4YaDu+
bno0uL5GxwFGxwi7ZrasvlhIwLzIog1mQXXyEPvd1DvDq+Bk7NTH/g3ROW/nv9wKw7YccR9cqN/V
ur3TekV0QwViRmILUsxZ61Ra10PSCoK2lo4PlZbQ34gaeMRffYY52f/ZyN8Zs8WNCnCRmIb550gP
rxIc97pi8DzPXiP8JKUI6I0SWTVtucOJ3kPO8yEiHE9YZs0V9ZvErwCSXD7YsqGT65hnff7orn0A
K4Bf6J9yH1mP5tmSmyKna6LnDH0ffaXdAfEWKQZXi+W8bXslXIX6yBIUJttxTmI2GmanqQl4F+/6
HDGHpd5xe9u8INvAaOTbwjR3n1ByDRM8htfGJ2BKGbZ5DcBNFfl4PX9iuXL/lkfhPZc97W6Jm0QQ
1X7MRKUhIzbFmMTgenJ6tzSbZywFYcJB39UZnCb4ObArpm7yEa4YOlPzMjCR6minAXnzhBUhelKO
oty9kJjIqw3IWmrh/GMByBIRgzVzfsmVc/ZwbN+T859eOITqZG13S4614SR1fQNjZElvmiM2hfqa
gtEYLm5Wq7e7mCK+obJT6xA9KrHQSily5FWwv7XV/qJGzXxQpjDfO5jwU8tYjyRfwk1L8tlLQjgT
Nq9/oHPnV7kjhxDIUOsn1VFIcDrZQlMJcMIXCcGXkVDkZJUAC5xUDhAvXorLASTOz18ErpswXjaW
jFzew+O4s/kftI7YkiCWGB++XxXAs/Zx5TWQoBqR6XqkhxlmUtETGPF29w1RSgaRdeeHuDqH+e8b
D7iPjGYnTJb5ar4Mx1muShW4rN74n6feZpSlN9ElBebsJTzMmFzqh3LS2STtGGuNmrkDwOQ7G1mU
pAQLAeSa/O7XzQ7iiH2HOQr8pO2e+HOC1lBodkcTNUgPpPSmt1rRRJJElXCuhz5UqaLSCupBwWuP
am+1WvAN+Rjvf5iTdGD+aoFzG0cMctarIGnCnqAwP/wlQvX7yCKpeJfxM+kutrJjeEMxJx8SGcZM
0kYFtzfq1IcG+9/hUXpSLYULyrXq3JiOQV2JVIv22t2CVHFJbNY8WfyYn91URP/cz7VgiZsZN3HR
eprGcfgEN00FQCyjpLtPXDRYudpxkBsBbE+j2yZQ3k5UcBL6Q1fez2Ue0UHGPSg0pjbiwOYpaggu
/aXPVD5lfBhgVob5aNrHZ/n+DbsoTWk24sCJwT2LUh694Fgxv7KxH6bpd7MCrkR35pTqFwo9XmaU
zDSVez6w+gKDq0RWp3wCRTZ74eyIdVdsRJVAvU98miIpkIMzLjtAqDJZY+qlqNBuiGffv8LLv0X9
Sde/ij8GbqkqfV2kD/YKkJVqXoq+ZHdC4WBYzNyS+zreI5IhvTVEN+Mz9LSh740uERTzu20x5Z1u
YscLMzBNTlSg4skbnTbdZnLMnMs2lgSn352+r4fn4D5/bwM+CCevqrtJkNMws/axbbWKO8fM0jNx
ovHVjvhC6OGaEQIyiXJgy/EQWRP+tWmlGUIbr/K8yz3V+UAwQ4rsNo2Fh7LVSH88p5tp85h2IZTW
4Q7u+qn+R+6tXxWGuK4EmUFLaqz/tIQnmMqhZVo3QBHlueOaz4BdA7D0NjHmGKz2m5TbFrptENA7
F/9g4XAXa2gYxjB9QkqpvwSbQ0xZPLY877Jj1EoKu2XznoHXOYS5jsEBiqcEmKSnLj01E2ufhnmn
Uea4j5cnzYh49IjFDMFFgINy5p47U+WyhU4/OtO2SH3fZgn5LgmD4KVzclbDNabB1olqIZ2aOiTG
5Wj/FlSJaRP7jFLF5eZny08Lo2ZVFQcBd2/wf4m11VKX2EzdRepNi/TAqMITp0SnaavjV71A6Y9J
PApJskQ/QAuvpk4E7YLPs9LZr9PWIzqOiR7IlPIpDGpv70a2636o+Mx5UaVsroxDGbz6OwC6J1kO
7/04vJ+H74naKXaevHoQC8c57+MBeRNJAAWrXTqEWKbLrRgGKW/LDprAwTphsTD3ldKNCzc+Y98p
D5XBfL2Ieso0caBDC0KNDK8iKgwgN4FVZU7TAQj7ggnbKY9SuSkxxS4a3dGWZHzQg37FQ31B017U
Puu7ci8qkwxmF25xIoPYwhYTr5GmPqIUjqW3w1l8nJrggmBbtQCCr7YB5tGi7LlHGNHXkdzH8W3u
QccKDQxgwPPNINXJ4S0CWxM/STsuQcM4n7ve69ioBmTY80V59Kv000o9j4WTdqLq7KqBHlkmXLNr
Jkk/PEWFFE/xPudTiEFTauEUo1VuyPJ9hiOr+g9HbzUo0uFi4m1uNkgH4ViQcHvPg9CmW5qZH7QL
RqIh5KNjziWUf+VZnUwlLli/TQJ6jRO4Rojd5MnjQLM7WvMdWnmhnJjcX4myzbdV8BMekuqCHTOA
KF8L7uTHy+guTbuw6k8fKuUPfY8GUfJnOHg9xJgTUyprkR1zTgy8MlkSmE7lAuCSgsL2Yc1aafgq
7lQoKUsJt5tJ59pBfV9md2JtQgng6ga+DpFbgL7oUsSOtZBBSM0l5hzDoZDK9Tp2PMVLlGSJntoe
rUS52nxwN2pWDm1Y68+LjDpb6U4K3Y3zdOZZwyYCiS9VkTbKaY1O7yh0Rqwp8O1DSfZiMDPKOnck
fadILGoVcBlR9IvoCnxHMRvImULjTXv7JxgKgBN2xC8JIp8W0J5C8cy+ryWd8qe8gAb8MS8JVOjA
2FDwrKm1az442JlVT2Wq9TF1rNF2PvTDzehpKJiYv38Vg9DPvvnY+3NtBCegk6MVJQDdn/2Gw/yE
j8vHSdcAhWv/AL6wXifs/UstAVS2wP1QX8V+tQqT6mUHpxpU8dbRbmpee9x/yDaE/Rj07eWRi+Am
cWz+5FXf+z4/73YOAVlvEAiBXFl0qI4ASmXm7dzYSNym/wmiXMRihs59wKjZwIna6Ss0sHS3oXOu
HDb3+MqJUnUAIfP/LEXJb1CS3PrFk0aW+Hx0MrhxHLv9+TNx4aZ+EAnYxIstOk03DDMgJEEaS+B5
sC0iDx5dZuLORBmnMk4Y++oc84UoVuyEgR4+5JTjexu7PqZrJktmPtR2vSAX9Y2icpjDjVo/8hVb
B8r8t/IeXD02Cx/eIbhsUZfAdELOkO0CLxOTuAhFOJNrTGJwPYSyQJgBLGJCsASab1TLGZ8gotmi
GMVnyB46bn28V7W4Ueg2axtIHU96MaCPZUHD6idNtqkWw6PMMlzIQkrWBkLd28mWSlUCZN5PzLM+
10kXRIo/b5ADrcN/25c4/B0WcFxkAHyiL6Yl3Bj6pQwlFYaCEjFYO59DjZt+rKC00v0Zb7urPAlM
dNyhLspxe5DAsSmfLCR3f6N39UFTFMEQcVRn2/qiKwmJ0C1+viUd0X6s2U3gb5CdNUi6a9YVsXQ2
0jp1Q/igtTdX4EE47ZmbXUk2psko35alD6VbFRSDn7PwOIerAidd8dTMpJnbn1GrPYRfeLn0xid3
Lp0mtrTclArp2A4IFXlpFDI5GHpFFDCLo9dxrFnSjntHps0y9qPCb1hb29KbvjsOB+e28yBHfHyN
kK2lXRetmPmYjAlAONy0w7UAF8RTBcEWsVUgyvlKg89V1TbWHdQI9WTMIGqrGFomRhn/AdXGTwgp
wJb5pI4J0wyTz/tVYwEXUnQFeztQZ5rN02exfuSiHC5B2XYtyf/3GOGNh+OHsbeCEUOqDWvY+Hzw
uDqIWGyYl+ZL0cb+kTrE5uAyvRhn1opTiXvJoyoUHRJaFZSdAg6XZ7a68abmnuMMk08POuDc+vt0
KFHkpA5TkZvctAKEZyu0dajVsbler+zawEqpkYHpR1ez3aR6eGpfmkXV3ARI7kWGGGezGiF3wkAK
oqXBUzc8BtgpdBZAGQjGPVNTpoaJkQV9KcaE61ND++5//F8aCbjKTmpR7D4EqugchL2qyUurbkEO
4ApxeYt0r9sS8noLogHff6vDKw3UIWxQ1GpJVlF4sa3dRVGI3dAdE+2e1SHQdDAlsamETGpZwZDI
ASwiByj/w+buvm2o3XqeXLHoyS9uYDjcTnOIMiKcaXF9NqejfWkQozUkTQmSzdgpQIDW4y8o0Tlq
P+HSENe/rKMJq/Y8a6sJVuRMiz4DjvZtMr4TKsdPh0S90ZIUxxkLypD71B9byXBG06fwrKV6Ltpy
dRU0j0rlgoOEvfE6IitIf54cXirMBtTVdnXRMXhebqAc7+99aWNo3eXbZHBnWVqBRdsJ1l1xpUEQ
C6pQZ3H2gEH0307iSEe9ziPqDJZI7QIXX/UOPTmSMr1WUsxBDLUo8sYjsXyMGQCIaCK6ws00zg73
3HClsFhOjm2/XUwBZdix1npNN8L6adasgzE7BXNL8dLpbeP1XQ/9xsQ4l8c4XmRY7mywE0EBpgWc
uHaVOOYNiUuuEcfz+fW4a6ncuc5CyGYBhhRwRsgioVTm5BJqYacA41rPeM3+rC9yEuliGchgx2Jq
Ffd0KODNhWNGQjRUqy4p7Oicsr29bdyP/aiHh/OkcnBFX5/3Gzc+tXzG4RB47cWzMl6hQy9BVBhz
HFCZD0VLkWKo+Jifwfs8Ht5Q7cSQD8rds1vIs1qyVjh/II5wZMkKpVtSMA2GYIrkKtBeLcI1KrvJ
QDJTXVkUGjnXdEVNU1h0fn1egn+FpVSHxvHFTTjv2KOgzCda8D9fSO0weRvlAZHyX6YuYd6PqE6j
7zeM9n79KRXLneZ3hzxOuS/lz93bbIGESQl/DYe7WHfsGzXoDroXQWTSeQQWFWjFJh6RZFBGTNPc
2Fa10JUL6KZO/71CgB99qqPCdutwJEB0WI7O3GUhkMTF6hhLY0u/Ba1t68kGapBoiRGEQFNdhT1E
6rE+ZvnqyFSkJxeu+ims/a3qiOlGQZZURcJ10TllEOTlR00IwnEmEzHXwoWqBw3lo54LcMPjbeJ1
uAlEOYiX2lQDGFbSxBvNQOVV9roLHMLihRKdtwYOQCvHE1MEcqCYFcVSUo5zxuQiX8S+B1uAYqgs
Q5no9XpEl0ZKsd4H0PRFUpIEyMIiS3aHtDTWpSK0DmySxt6WLMe8LVGh8kaAKt6yJeS9epFgdWjo
TACy95w+etUAuPnd3cwsl3w4qKJLOsUD2DSpGCVCjQv873uMoMVTi80MuDKvJd8IdDBY8F1fGQws
z0ROkJ6hbymAqF5lWGcNdshAiB4MD8ZgV1f5Vy83JLonXcxr1CSrfylHE/TMAaZMIHdLTU+grMO4
q/TaJsdnENCdPfk7wDEfGc74+vqnd/1bltW5Jvk3YS8eQDkh9RGpg9IXoZtBIBiXDitgeIqpekFm
V1yKObci0Zy+QwgEmGRc53flGirvm6gpEnegXq0qX2XUt66Eu+VJOoziTdzJTCihfxgYu8B7VClS
6mhsLXypGVB58Cdk6nxmMoon6xPNZtiVqQCu38Qvkntc9IdQTyhx8xIZ9+Y6qczLB9ooWZTbnqkb
cZWBR+ahO9V5IDTWH7LD6iOIV8mpQl8BErVED5ewXqxRaJWdgy0GWvedZbt9b2mkSLnrdqB1CH8A
qLtpqMGOqNnKiXm7PbPYgiyWMDD1PjvKxf59YoCUjLgHHk3lu16NiZmnAPiP/bYnkiPSBBHHu8ZR
VdSMiQ/NjYknGoDrpjEoyi94o/z8Wq4jGwyuCeAUqVfp7ZVyXFwjEbve5QkLmtY4aqa6h52HGUtu
8jBcFpAyoJegD5eFNKAJQ5GB7tEh3ThCPc68pvqygVUjSGUyIQNpc/aP7x3nKLbpDa+abNIzc2Ed
I/zeKDAPhqQR9bn6wKFkLnsr+YAVBC0z36rVuc2uu4Yutm0dvBzQtAMX/XTEBiJ71wZDJmSPT/VX
Lafx27UiZSxEFX8n95H4TUVLUlfidFXDPwO/Z5eEGa9WjGLCm4VPX2Af0ZaIj1bFwX1sYaRBkjSA
pZCmXkWFCFZHXHlwE0BdU8Fv2NHkPjp7585mr7o9+EBPoX45zR8f55Y42vAqqTLnZVvGVo542Omh
k1sz6VbR1BqlChqFUTgTcuiBbB0s2z3Hv+lI+hdBquvY09eY2vly87mzWocVGrz+IqD1rwi9bXZl
ff6YUO+SzGIq5b56Ns9kYkajgO3hY4T84j/TCCHlbPnZlFY4BLnRV5x8kzP7M9DHvusPI/hEcf58
srGkL+/4HZqySSK3daIzrma5WEpvsS0wI4PIBAFyxzgq83NqY0srpDGrZDbNUeECc6AHeORHXHxe
NlZH/RgLMiYll60K7N3/KiN6rQgKPKVd6luUZ33jY0NPtVn8hOwsja/xxKA4eTrjFPjJMvqU7YY6
wuNDNRcCGDuOvNjj77tHAxdaFpRzRYrrxkVYYDL5rnfmKZl0LWY7KpIb2Py1Byv+bwOieniKCffh
qXw/2dI9mN1jteknxCSUV8PRX53K7iPbmqr35L5e/kuHWoDXEUl4MYPYBA10UScYkc51ocZZB+gB
kBwo7pel3PZ+fL4vtmlmVpCExgjcCK+PBizh67E+Cimh0IFUoRrkpvwVNyBXCxR/T51FEbmW1mzQ
/aIH+WvSJRvBeZSHvikm5Tx/FqFPVG/op2/szWtyPvBwformdsX/m3dVNiOs9HxYMH2ewklj7m07
/ctCGmAjq7bTqP6xQLlF6/pMHH1FPB735CPN1sJvYVcKOvXrmlMZZit72RsNMaUVqBB2RYXWFvlI
ZVBYiH3U5svHwdQ2kYbsBNBJnmTaTByPj4Trkvo0fHzZyIMyeIXh4MPweH+JYvYXtthZRowUA909
+SziuVcUD5d5hO49zSfvJ5D++BF83nJpHtyw7my6OJBoPxBl5I5tXDZDLppwDY1uDMu8kdVvIBf1
o2IdiRMmNWckdLcEOw6BTZOMZqvWCRGnOFoIBkXWKtoGjaV1QFmdciFF6BGsFulsW1i73VxU3t0+
sktcE2UXC9LRWd4bTa+oOlWxjyd9CKWpT5R00F51AFUJPtplVyHcqTGW9HSquyMEJTbxWrEaYMLH
rFYkQt3xmZe75NiGlaR8SP/OHRg2DzXXQQUk0r4U6klxrDAxstoARdFV9Z/GmPZfV1yr+uYDyhKM
AiR+AP+YJzEK+ZyukES7sxVyr82ddNGTYQgJbpiiH4eCqWfJ+fsLL86SpAJJMCbf6MFl0kcH/3xY
l8LBhp1dJu41naeng9aITiyX0lv4x9CkKeLe5BsNjmV15CiayWSrqTPOpAvfbQgJZLnJYsuA5HwD
eE57C66bPLgryFckbldQtev6wDG/hlTkysPowS8B/+5STdJapErINnr73PnyhJK7YiqzFd6cMve8
bfB5LDhAr4lAA9JwSQwdRj3ERViUW0jzfgalWeUa30N8lb1CHd0ZLijdwPcFyX+y7cD5uB1WFuyk
J4stcDUCOydZ3rGgvk580DdosCfJmmWibdYhAzm9a+lAo9aYZgk9CmHWanekbqwf4VpouEl/IxNA
H2PBJqkOWzpWmjxbDQvecgii4fp4S8xcWBPNpV99Vz9PJsZNWhP1A9mBIO7SymAWArwLCjpV0SlC
LAXzVLsMYFtFel7Uk4HbuTDb3j6e9Y934LXL8soGLxKwU7hCzu6Mut5XXfO0F/2O/1yuzMQX1tZh
c37/BnffGvpby3CELEOsuLVM8atZzCs2c4zpp3J3+c/QJiHkleG7N+ve03hSgXjNH25CnT4uBwv7
rhvvFVmIZTL4tjaclBeSpdW8p0XXDRJUbUNKh4z2nRjA+JP/unoo4SSW3Q3ODnNMwEa3Eq/nwjvV
T3vJFQRLjDs/likwc0V89XtJRGE3mS9+Vebw6bwJsG2gziQuNVK2LVw9t3QqTSiYPnSI1Xq4nEWG
a9P3qbSwGXuBPZeJBYJAoU4n7ebKLFY2nF+6m4lPM/E8HUEbBmsUARu0Yyybby7z6oBmjmdz2K1H
PPI9m0wGHuXFgfsUhKqEuMMRof/QkGtm5BzS6Lo5s/gySf1fp4FPGNDXwGBWym7I9SEazMKAYjMf
CoFEgss8tmQe0ipnyUn0iRVCJVqoZxWkG88aRQe6Pb0PoDpItahRIdM9SXAdwO9X72CirrxhaXB8
/NNppPdAibzy/Eb2Kj+sajLfI728/s9DHtIHFyqTKuFSsG9bJ/RuUG4E7BSXmVCNWkO4/CdAobAs
Appj5mLrjBUo2Rc7JlkLWGY09CferAT3xhW8T8/8tRq6sqmqGx/vvkfae3joHq3i/CSc/PO4aDUY
KMpPdciicAyFMZTdc4KSujGwrE4Dqii6Qg0jgoR/IqIrSS56z4kJg+AwFEK6CpUnHUoW9OsZZlvH
WHxskBTIy60KsJGYOXd3WojCtbHXFnOYo9UnJlR3+Sv3Hawqj1Aam5RgDKctEEgZpo9FvpgsgrKS
w8kQL3Vj4CgJiAPoGZ1RrGYz7Jua1/t5JHXCFztyRvGBs9A3AKHh3FzcYTt+PWnrKAIeCe8+waRr
EdvtlX1oK/SebSVzSgtwpO6N7wflGbYCdmwABXgQK2khFsD4+rTO/Bop/UnTbhm4hLjPHy4Sl3UI
SMgUDSERxYqiUGEr3vSqol6LWO5SYiX8oDJ3LwTKThoGgYdobVc9OnVAG683ahsq5Zk2dOAITYpT
aDr0+cYlA1QltC+XR9TrVNG9V/4CyiYCMhkjFiqWupHEnwseQ+MSQGKan6xaqtwQwwpAHG54fD8P
UR4Gs52VT0YC+I+Yy6cYceS9yI7Muzsi7OrJW6tcXTcj+QWk/Ep2gPVEdugZSYA//gSV1nSpB73s
gpBZoiH+Jf/TkGZkSQ3wWz/InangqveYQGj32AKUybDZ8AXIAL3BdHLGNERZnfriJenc/EuP4p8G
Y49cX65C/r4Y4oCzOUl2uZSavYlz/Sg0yxstJf5Xzw16F1gZq3xCg2cM2hQmIypDOuHOI6OC0M/6
wb6imVgEvfwzoV8AE4J9BeA1GzD+bJLMY3XJepqOwIptKum5SehSc00TK81SfGk79cv4/uKvdVDo
l2rbsQtGn0nkivxNDp2dLJxPBdhbyM9Q5ignK6K5o8dH5iJkDEJAL5piBTt+0RZ2wlyNqxvMHmJ/
bK0tCNxdK7LZFtZl5SzbldFOhJ8iIwciuZiMoFAP3FNE8/EvZZqBhxlgtG1dCF0TmKs4aNie7uRg
V8OrDkA1EhsEUuHqLzKvEeieRTHhO5wpxzRfvITqmxscRDctk4+JjZmUQ8fRhG7/BgL/oKn4/EK6
IE9RwQvArgquDT/mOgApqU9v3sJCK/ROlq4dn+DZ8aJA9xxL4orJVY2P+VLel1rluO1lwGf7rKK/
kpcsy7yLWaraQMYnreGC+gDdtOoOXwQHP4L10eCkUaoK6YMDyTfagzE/UdaOMs51B3MczTIn85RT
Ppq1tvPW+nuvudmt19Jc6o165AvvZBId+DY9U5gyCLfq5EUsL7ICQ8IBqEBqy0OJ29Mty3X+t/17
Ff8tHWOGWdYqiIjOic5PgEwhsY0CywsE6FkIUIc622E+pj4Ftw9YDRRwTc92WOCQEgiqyK+AuHo/
mPPXaDB50wUX9Ijt99MF/J2YaCtB6J6mFBXPxaj/cfkwV9VoEMPPzCGeaoawoYmMekSGw/adU6OG
AFzjPxLHffF8nEggX15N/g0E5rO6Yv3ugoN3gw+llwgISAIcmB0JlhvddH7VEl8HSH4BAqi8/okR
tcaYjhFnN3HoLiAPnScbcWmN88rh1E6p8mCO4R6UDJqdTsCvtWUC5A56imX7QYq2z3DTndf8mhd9
NM4cHsHj8b9z94SfVTecQgLpdra4W3eCQMh2GO1Sy0t0E4T6eImiS5NYG+CSvN/Mh7iNZe1j07LD
yt1bT2Pn/M47d1cS30KciNqxEmL8Rtx4s1f1W4d+kJnIsB2W09KIq/SvauYf2xyGPcE5e04pCKIe
zDUi+2g6642xpTBZF2BQA5l96RkpCHBhGxqC3fQVDIyoPucHxrMxzldmdAQ36GppFGs9DSx3ZdYh
1D3QURp6Aj9joyItdMsS0rMEdL144cAGRaqooTOujGlPpCFPsP8JC66JlcSF+TQppNCBJhCo0RNt
lIMlEGy9ArErq+pWfQvb2ff3cdkKDX9b7fPWQ3741KB8vIhcM9dQLC3y5zv9Dye6iQOt5XpGVEkg
hdNDHxqbCZQfsAG3Jfm6LQ7m+rVT56H5lIUWRHz17f5dIbIEd1rsr557npWRPn8sRuuIQUlKxspX
3EfzxM9D9bW6HIx538GRoVOlvhlQmsDWN0C56PKCH9qPt1IARJQiNBCtpnDzxbwXcpAp+BbDUBWc
14djKNEzsJpDxivqZq2kyRc3+eYSfbzxfnJhFcbT5SpKnrHensZr6KvxuUrmyX2jBcnW/qOZfjC5
rpQwHRBOwCt6jz7EgxB8BRRfV36Wv/gNUt0ssDqIery9HRcMgsk+dEDGE7uYHNIbqFDE75givhYo
ibnTe33Puyo7zNIKXt4bm0ciiaG4KwCXOnhxqhgY/71TvTj2SIXaDQDXgiY36wFYm07y6hgsiCtL
m40WOkzqx0Ls8TaAWsIRTokCGZexHHJ3tHHLQ7KH2F/sgvQ3SfXqSz+FWcxjYNPgvFp7XnzriiaU
sgXGNZLSBrQMBntz9LUKFac1IkANn1Cq0byXkHqwAkRa8M4HQVmlvA4uPIXNm6tt4DtBf5AxKzZ6
Nlfw6YJdvOnVjLXOwfXim1IHdCt9hLJWcWlEXzcSIlIdD2p8d6hQtAbvLrF1GYaqz4Cn7f7jfy/g
2rpZlk2pQqlKubkHodPLn+cIkaJ59uL3bxO0W2b8T+og4LkSbkweyOK8+AL0jYJ0YDdbwXNBGEhZ
umTtZUDv0ADw2yP7A2n4is4BS1cgOM0hQibWUiTTn4jy45yN6WaVyL93scry4khrGYjahN685kPa
9T9aXyy6l6CVEWYtI0PUIiaOJgSWCI0iXlKG0LKpAwhKPXWhn1tVkcVUWvHUtxDSjcFQG53V2LtP
zK1XULZFmu6vhqHf/CX7iIyprS0VzvACPHM1220qwVjOH611abVdORSu8281Rx+vXPZngITnj/Bx
ZmC/0tnwistdR0zycoZAupEybh72XPk/DDuBvp+bl4mizLKkLzaR8uPDXMnaJQqm+gATbLxHFyr9
Rk27Wi5l4PbhlQt0CpWErcl8gJ1mWZVOutGhZnQF7ESEyZuEmNCmPldT74Ko9jiUEpca56Z2Tt13
+35VaWK4sNkMxRg/Jp+W//36mj1harn1R9tbdTZa1fXt88vXP0bkMfh0/ixMNLoC8NLANmVkrOAV
X3+Zp4zg6exki/UD0RiNdY3dqGbq740MPI7twTm0bybEhXwUKUpZh6FQsoZxSPsMnnMs5DabR+bp
YxmcDm31ZoXXeMUgYbp467+uQeROpsFnQQReZtkwZFvnjlQ7jfDEUKTGKTDGwc5T0/jAl1vgll2T
h1Fze1alhPUZrESuRPmkATwJSAZ3hv5yD1pK7gRQwZpCHY/pBD0chZIO84ZiOdEkf1AXqlcxuUmY
RnvMWp1a5l1zk083oQMBs1TkOkGbXsxMTXwxBGWd4qxU23QwsLhWQv3dY6BdAXZkbOh3X+U8UzvR
QE26KYViWxPBG4cbFSmGtpMbmm0sz532IWhG3lqWQMDdPCtbAzyRF6+uUMKOXHyXmXbvi+52C3BO
lrtn5kdBgQuKsRoI3Gehi6mYV+5E3b+7gtCg2+xCASoFQaTN3fDSmJRtnNIk/ZjAsz0FwB+cTFAG
nk5xh2hV1y1VZ0I5aWfAIFN7H4PFsQbXBfVgZZIJvGEmvxxVLJDBnGE2FPouJRDmbPdgyA18YUL/
5vNmhyM2iPlxRoHwlW3zeJrc19iQpRY+0T9vB61Kq2mTihp4zhXY5iI7jYP0JNCJDQCpD9QFZQ7N
ZTlXFI+CiuWdScXdf2oBNABCx6TI2AibR/vqk/O1K++UKYYEFogIC7v7WPS1yzY6OauuaTGRPsL1
wg6iDfiXFuhN3mnhxHcxGKC14CIL18miI2VLo+AU/KZqQeAVgnIK4LCiLErJ2aimhAunowPXXSFP
1/hpHiZwwczw4wd2ALLnkCWDoMqQUFbMCdgFDIpYJl++15UHJYFAYoQW2iO0LGJhAy27iwiWHQNC
GSTnW6snpfIEWFavvKkzNBecwNP1gdLXtIPzY1bW5DpnBgbGOtsaMuPHaDYGGg1kUgotD1JJiNeW
QlYT8lb6u2Ob7TBHFBNdlMVd7ZSwuAifpooNHTMS5L6AUU6FjuZXYdKacHcTlUT3BAb1/39zks3p
mjwyz8FrBphoLCAZ9iNUb6fB7mbBss54sbm6PN8+hRV+w1jAUeGII8IsvDaFvDx/rLjLqixcQqz7
U3O4RGLvCunoRS7CyiDpSIImmdQzs/zQMpTMxxDymcolON8efJ69rys2FaBzy6xfzZQlnaHh9Tco
fE5ue5gURMs88Wqc+6ZMH24Cvj7JDpaM+9p3dBH1Kbb2L5P35ug52Zqh52oN2ibiryexM/zJQFyp
NyhgFrJlouE3d2l6a8wyAABt/0h/dgzqTp20qkATPvNmsKYOLs2I/3O3Yyn0AhTCjOlU28fpIRA0
px7hGKMpahBbde3zm17Q/hCsE7S4OokW629PiO8gaKt6uNIHdfBsZBwdJXHPSKMQz59DfXKzYwHG
AHztz+uDKZC2een8YLIbdCPTawVsiX7RfuG1H6y7B4hgMTWeQ4+pW7zVHEK1AYYHoz5zqvQLZDH1
XcKaJUjD2S3IXB4IukZeLtM4bbGDpFmvAnQhk1I8841aGLRpHpIoj6j/Z7BljpI6XG14PSXP06Zw
Ixuy1rsswQZNI/Qrs5OXxO/Az2yznyW7YLGBQ8otqlIuugkQgIUcgCsrN5EoqAgTq7Je5CCzOBL9
BuXfY8hVa5WCjP5sbnHdfJkYk4s8dKmLMRY6Nm6maNrundhQGeKrdhA4/hNE6gHOTM8fRXvLlMbi
9BN1xry8WPeLPcK901+0FWfYf3dgDU4ndysCw5VtFYR6XcEbeklTXYWDVonPBCYdiGXl05p+FRDq
VGryh4cHlZ11MrzA2/it5XblKGyi+drayzOk3anXPiBXvvElEW+BLA4zZBdpyoyLFrkeo7kyA0GV
ARz8u5eMtLk32unk4Ult73dDesTMkvRpGdhqefDqSlo1zwNswfNX8pBPbzLEld3jLKJk3n8NTzvp
6IRFXGmxCwzLawZhJ/I9gqeVP5g1wct4Ux1qjZNeErKFqDsD3+9lmWyjXPICBADNi2jJbxrBc4/h
qDhqZ3zJ4SazYp1wnJaS00ZmQ5iWrXubMJZqcqoZaZhHSNQb88rtpgMd5QsZaFayAuQ1TIfcWo/z
94vZkO6jqRQg1FIxty2CyXESjqKkvdRf6TH8sDS1kwVwsVrWpbo7UGp9yjKF9kPVkWripqCLvuS6
cecjTYIaVbAeayXa28i51ww9RLoAIj43j2LtTwZ923iZ90a0Rg9U5yau+d/PJBNEAP1B6eQvYjZs
CN5AUC1QqVTglnMLBb4tTNMw08MzQf7mHr04SMdRyAMEsCC9hqQHrW2IUCIhW74YTG8FxZzDnYmW
OFLH4F4n4sa0GYXZLZAXLa0HPZhaU0ebOwWC0Zff0/escJ+L7bWBP38Uy1n2YG8MgWfSAdgGYV5Q
S1dYnuVpelQcHvPVhSxiWRgcWdt9zrZfWDumEcBdkmH1BtGJLDBazxtKbkIJRsBOYZPjXY+uzN5f
Tj6o/Praoe2/JhIoay7vCcu3ZVMK0qw1tKCznhbsLfjvLWWtzHk6raPcYhu+GtPCJ4BUZIPEf9uU
LDRXEjzym1TwOV8vLGC7mo+BO/PpqwBH7tDeW+HAit8e2xUxhSlU976DZLuPNWtJRdajpHPptNW5
mwDOwuIx1EldEDAWejiQrS8JHdlvrK2APStkV0Ok/CyZle31P+hVxGg3EWD6y8/xryHAaJrJo7xi
WeynEj3LNw4JhA13IoOenU/ks8L9RsjnO8koNpydf8DorW3Bo/uqgviu6QRM9LB/CmGqCOPE/Her
ALUH2ISfrK1J/WnR4u4utq/ozB19CR/UEYXnEZgGovunevMI9WeTY1lNyFxc6qe30ndtYyRp4u+2
br+QQVOMuUX7Oid5kiieJ/2URANBwsIyR0uNcVLPXTW8b6bZ7ACB2tg9JYSxap2EN0XZB0gvLrqs
pSsy56tXancpNGTvDA1/YpF+4IBi3ZeiWPLIRihFD/wbnOd5d3IhNyuqagMXSdCd3tiNa6E3ycpl
APZxmnK+iP1B3Qoin/OIRM6mE7Ht0zEN9rxtXfEo+tNt3XiFEZBXH7DdrnRjrgbI/WOLpkP4A8vg
FpuxyMBDZkchvUIcvJnwZ323osdk7MUT5+3SjCveGkv89yZmMbRiv3GKokCdc9FNSYU9dhyt49Jg
5KtYe8OdR7oxO58Pr0vtNwDCYa973zY1POSYd1X5wTXzPKLy/dNz6h0O2AoeAuzegW46ggJpK6/e
FBhps2fezecELj/j6pwj2NTZeLnm8O9x+0eOR5g4yUoydDtqAp2dm4vgDSISeCPmi9QvKAL4qnFR
xqxrDV3kMy1QIdd4KdyHtotEya8o9iIYzZrx0VLpJlA9JYhHmMgMoItLk4Pj/MCnf1eGc+a79q5Z
51Pa+9RU4f3NyyFEy4fY1GazXN+3cZKXRZYzSd4U3q9gr9F6IuydstodZb/0lnsQZTQknekkUnV6
NQE1TM8cSzIa+7+BJw0fMpOZO14EMLnet2uJPDQWOCvezH0VohFCpFiy92Q6sf7yLJPqSH3dW8AN
TCnBgQ5+Z3SsR+NuYE+yeG3ZO+cGBDPn1yq83tvURIhHP+Kq9eWf9QKODBpy1mVXnArhwKvI2iIz
vDSiQFOrgTM3sB2TtbvZV3dV4c6+7HeKIVjFMs8ZVRk+v0fBUrvv+Msttmt5kd6k5iCEjxns5yId
V8RqVgeqMG5I5f4X1of508av5IEx4VXmNXzxn6Fm6JuCXiIwBfnDU0WdWcnI0HNPmh0DKV6OAt4Z
WFzv1tGA4j1ivbQcYYa8rQrdIr/0ILSwa8ALgx9GnRVnCX64efzJerDdYsPjcqGirwtgt9RbKFiw
5itSpT9n9yZhrSfzvxhEzujYXiNWrMAn756Wmz8uRqiwOXivefVLFUWMpaBITXX8j18grYCDMYAS
myVgUcmzgTbdifIUaWoNMSjPmRsUkZJVDWvJOhVlRVgLg2apAcuEdJtFALeNd7u2ONx0/B6KlTOM
jX2GH1+yE/WStiONkt59KX9ereDKysSP5CMFIzdphSlguk2dtB82udjx2R72GDvDCpqRn6/HmwtA
6lE/PSdlyprXbgOfXNS3hFm22c+vnZ70yhcEuTjYWsXnhaw3hHTtufJQZCRnqDuAMDzZB/VF6tuc
mrG1dvDcSvhG/sqSJyGk2wjtjsPAM4BvUgq3m/NVBVQlSNEpA0hWh6xgxwyKAJYzTFpXAIvzjiF6
JDz2XXK/IeVVv2cwgHcPLKeUfSpqiW3PK4Wx0yHrr5y/AZKHEkHs8b97grJcM+FR3hNtJNFOvTww
mLFqFNn6NGUFfLoQeJPQ0sfiGcDOX7BpueFWzbnHW/+tUem5F5A+jgogNgjWkKcdYwSHNKGmLltn
FVtPNrwpezFaczC0P7SBQwVN6rNxkczY1PL06wRTVBLYp1jmTG/W32qVh42A11iuR4u5ktBENfhS
OeRv/GP4u3gIyi7RU/ELh5UNZB+xaavH0x32z4jUUB3kvpMrvodugwDl1P55CfnnfQ1aG+MQcGY5
YuRssqN1kJLunmEYQfUX7Xq02E9fwYExdCEt3FM4ieHcxVtv1Bm3XjpwG+1QYNCuKqgXvLrawr2V
3Hto89ZP3qRR+p0HzV1oI9myBF3+uJnv1IB0f2q1MQGUDkFJiwKTccTQwEcQUKLEbg/jfil9zoF4
gvCHKXF/aqV87/4CHnuueTLI7YdRqI8Ajx+/ERd78AaJLNI3+ahrGSCTdxlqwlam/+863I3oxiLY
PVSedmmnGBBGf2Ug833TiwjxxlBbebselhRKvgb/wTt/JH2AMiPQqVM2hrsBAq3/fX68cF+JrrJK
nyD5Fc+4bCJ5TaqefDH+L3VTCHOuLwres7mr7M1ZeTBAhs5TTTm4E8VpLRCdDbiTTyIYwO68kRIw
PWnQDGyNZbh/8Iry2CE5D++Lt7I7SYCk5goANQ8HFXgR9ZkPldUaJHN4YkcmpCxsuRqONs6ZWeam
LsI3c7M33Z+6Xq5zaz2SKMotlD5YUJ1zM/NZ55VdxZQFl7GeU3HDsYm5mvgnDhpTIGrFdQsF20W8
Ws1aZxnikJESwk/U8zvsRqDmK38/B0Gt6Ha48YmRfkhODU8S9oENX1MUHbQlDQ5ESJDcg/fvApMI
kcixitKtm0toxl2ulJYgRXNldb08YY5V9104RdWkmzZKFYzZGdNVbIFa+O4uX3H7qm2QV8FmjF+e
uJVMH6blXuIa8LPL/+z9B5k7n05DQn7XecHipiufRajIsJb15F7B3dJjywivkxEs+GSBWZJ7rn3+
mvtk7sNv74gel38smkX2pIHfTPrSYyO5u2RPlODSY4wNgaqZl2D03bP47PHvyIiDjUNwIxVq2gO0
T6/OLYEhfYcDFT35ftf5e3N4bdAA5ZsP+PryFisRU0vwqb8mGK5gfWDuF8vVzi5Eg0sa45JtmU07
kyztJTAGAUlXfaC/eVM4gxEVLCCK5gBWIwgU00gt7Om+qnyJGCsqc4WZTf0cPvds9Pil02/pr/4O
rhF4qsNM9bKWbhMtvRHuoFoxtJCsOtHVIRjUWky37JKcEQ8ex2J1ofTOANLsntIur/3qBm5HOef1
0b+wiACTxOnMo4HG2fx8SQIhEioTHSZNoBEzCI5QnzURo9P7s/5Y5LgDtYM66Bra7zd+C9djQ0ON
AcQHLnRwV1Ak080cGtpLochGzzAeiyj0SRXqRHrEYzLb2uYc13uLjF0BRh0LOv6TeibjMV5J2Fr0
VhII9u+dbc/c21hjeb5Rm9wdk6Ua+j/WKY8S5xa6T9bKBwMyNc2GOkXI31tnEJb5ivZgeifot2qo
Kss7jNLhU0+UYMMx3KyaKnU54WyqWf10JrTnbe2dt+0LKgjEcEiVS07Nu3/+zdgBKEeKvtNbRjcE
B00uGEtMk/1e7f3Pt/D07iKMpPLrksJgbks/7RskJCeFDTWBbZG8VHMNpawRtoFnQbrgfomvOzk6
39wTaXnT5c+dLdfOKU5nQ7O/97rtij2FEF7FpDjiOfS2wRLxdbtbylAj64RbELDcginjJ0D0SpEb
f5n8QY+C0cxc0UOYEATJ0C42q7H1JWVbKwbZtWCCU/rjfzAugDntJ9TsQQvJAz7ee4UHMl/2/r0E
89bu8Q65VbT1Gg7V1ntMjCJmcX39g2zx4Xg6bftGeV4D+U2j6FzxsPHcc5NiHAPsYq6vDgTqRulr
1OIRkS2mIcM83coIduLkzzK7LYqGKNcgJK0kDgPBHBDBtaGwtQAyLBsu1erITqe28KS0mr2dlimx
21wpO0rLXShy4jHlDl9/DwvK63PvkzII32UcWRo2YvL4x+3C8B2M6Vq0hbedytrUoq5irU6PbyIQ
1g+3AxNBoq7ZIIeKokY7UtXiqYVMOiXGXEAquYDDPst1qnFDjwWJKhIuPTyTk4jVImRD8PZ4ZMSH
v3kRmAIMTSSE4C6ayvcvqwiJRDdmACDC0c4hApc6EuV3PX0gQqsXHCOvAOiJB/G59SZI9VXBaq6q
XM79Xrdb3YjS7Ewps7A2FejAaKhgxCcxdNPtLkwMjdG31vuQDBLXWDdoKdnyE4LPbJ+uhUcTJu6N
ktIzn46fRRy+DZnwiGsAHpVCAKGDX2jtBtuBuC5l/vzaiDcF3pzPNtpjCk2MnyBvx7p45fI2iLhs
s9gaCCT3k+xVRW2QSZLNV7z/dHGxQbO9kH7REFl01/eFbgevdDb/TqbxVJ6YMxpqVbUEgw2zeMIl
nKg0RuaQkKT283J/AfB7jTitmGMceNtazJC8AUt2KwLeF9UAYSWbbQ/9L4EbSIIFj1hkn9Judw26
VXS5BNM9k1aK6r1PAz8iA4HGQ+6A03knv2+jZaWRc4NC8NDNcUod374b9+zI6ROKfliEigKWumEK
xnOnlYypJRRPujpgiVZEogLb90y8GlCMo0FI3p5m2AAP/pPJkvhsPCS9vi1shUt/KyEfOGw1TtC+
+lrZsUm/vQK53LApe81FQCyjGOEO5OcmDINwAz2KoRtYm2bGPsrXX2IfWxKXhCRCK5GTcnEa2BbA
W2qV0eLaKgCLVHEk7mVPhUEUqzwQ3pufYlYYMaaG5SzuRnsT0Pcj0AT38H3jmzhuGAspDof8e129
skFb87Pq4f93pZIzryMgrIp3gPk0yNJfCyUv6gGyPU+Bq0wOF3OjHgel8H9EY2hvPIXQTqUBmpu/
weWunYgWarU7w04jkcYzFoJknTUyNJUg+RKgyEux2+SgnXySzfusOI2AzBg8SWmdsZiOJ4XOsYpF
Dqi8Wi11xXU5zn4oxaMTrVHdfsG42CZXsMVknK0xW2pQtj2eyBHr5vQMNpoEqkevFsfS3STbyPB0
xJI+h551GtG1mPfyGTaFs6ZTOUf9HntWQ6/jhyD1jvI5a5hMph/Pg3igpe9IsYvMsKysBsDgqQLO
ucpgFOdzbTeQVt840DBoQ00RXKGMdOQw3UScPzp+yCl488dAZGWZ0ITmeKJbvpKylgDvmKMEu/4Y
9E6TbFrDOKF7eIpzLwnCaantucRuXcBLGfFgCOWuY7GxxyLYeAFGE1Iv5kbyamVEwv0xJGh7F81c
7Hc9Qk767uqho1BR+de78ZUv94w5hIm46MKFKJSv7Sf1ejTh3KeMODv9bZovxQg9AxsxowB1UPJc
cdnjxvJHwMV4w9yuo/eXt/xUMQy3/cZdSgHbiXfROXWBd21VpMYtmkTUOtE8phNV4LIIXu98LTJa
Ll2pTWdog6oRKgobZet56hRORYwO8cCmCduhyxK7oJo/Lf2FoFSuDu3YaruWH6RKics4LgnBb9bj
RA6nstY28f3opnrzmaMLGhLBUBPTIjYZ947Oppn8CFPxw7GyqSVhQ3uDSXkCuVIg1/5yiLytSyJT
v1T/Hc3dMmMRmklaIF/jZ9DwCp6KxsDK2vTNhlVevQDYbY1OFz1yNPqV3l9wdozBgbkqdjT42fbr
DSAySX2JlO3xj2PkejviHKWJBOSNavxvLGAWmeMhTfdZUVUxPsYjBryTg5zoIddqEoEtfFN20VJs
fObSA5x74H3TNRGHuW8IonGFj8RjjPf6nGU8SLU+pRRBCu8tqzG268hnhvoO77p0/VW9w1EFpBZa
CkqRC6937Dk8moRZybSqffBpMKAFqXvYpcRROU2McvoGIvolAi9hQP3vbWBg/ikZ6ajPku2HuHrs
tNfd462yWV8L5MDzXFOz44vXWJmkM6kV+6cypwTZm6jhUo7Kd74+0L0qhHdJ9stuTTmalflC7Rhb
NjuXbrD7637fjzpl/d8pu8bwg2E5QSsLnUb2RGB1uANNyf98fn+mCF251Ra9a+ai4AxUwf1RfO8/
zJN8oRvBvLeqoECKbHofMqKFrE7ZwIyrhksE7Ing3MVwfi0CkZT6uE+kRGFIQhCblZqp04mZwtPx
xhYrAVS/JPrlLYEFrxdk/8fMZBfC1n+BTP4WMlyg3LL0kcv1HjKE/16XcEwndfB1hpaLP7+FpbB4
pSdSAZXe10yNVDwa/Q/+VOvjQHrCPWMMfU8jC61yZRfEQeB6sMhlUeOIfLYUoWuu4w1aVsMuWEMa
FSUv+s5yxsfG3an9SIJ75jitr1PuVhLD5d4vfhfcM9JFB8WJz1Oc9zV/Ea/IWcGOtB0PecxiS1Ua
//5QYGZBLAsVwH/Ghv4oUn2xlOllXyzYtWfs+RryTQtJpLYTbjnTc7ICYGyG0TNwQ7f941t9ebKW
xNfLwVU119g1YEfPDQBBVoBjPUAfovd8OjvNTDLop/jk3R+Nx4TEanv/uAo93+CmHTkVW3wvnaEh
8vqnPxKArI7wUemvSNALFj2kLxnKBLqOvbdBI1GOxILtrg4gjWJWbu7nSBzpANhRzlo4K9/v4FWS
C0biROjMxZewARjZGvnI4TcI4XkZcXogR93CoVkorJ9er2GQO0aDBe/GD2kbh94XDCTE2WJ2073u
8N+Yc27ZVZ/PLMSveZBDjRDHwLXL7Xk24hrlnWFvmrFmOBI3VrzXTJY3Uw20RLueYLAx2uM1Wk7F
c8tbPY94kaY/MnEkUMmUzaEYUw6OkRKXwzfff7Rvhj61NWAjoLV3ZWpXzjrm1U7FkdprBLMASWjR
ZqTOqAv+jBDPMCMEowGJ4yOwVM1eboDbXxDs26O4J3dqWqrp1Q43atRfNRR3WXDzK1XeIJjpWo50
f9faBnvf28q2prVOhBfErGjYDAVQu2nv5RMU8Pe24vQPSiXJQT4AXwc1shomKTcpIEnAQL2ZnY0y
IqDw1p7/zqmoGK2crrOU+ZiRLM5NXV78HrgTri41tMJJXfDRwV9MIViCiNxH8snqp/bz13+2oU4G
VWqJAej/s9BpPT/JCBs1pd/ht5Sh2NVNC8LD78pmj17ueEPja3fPjlUF2szh849hbcAwWzfuUeG6
vKbcZxNR//tB2YGOjr/sYm6qmwgUNvVY7CrJ1+jxOMzTy5aqxqNx+C2LEjbxRXg1PKp9k/Yb2bsn
ffUjnu5+GzuIwCSCyFmqSWW7saVFshxEoLvgmbLKwVnj9sNz8PFDCtFbesxcS2HKRzkkhnE/hmmf
k3f0dctfgAt0hGOfYwaCg9Px6QqfsDO03AjCAwYxALpGiaJQcmpHn0MzcPexVX0nu+uNatYHgKmX
2tLq5uAHF/Q/uq1RgRzt3e2//1KVBQANBH+n1r4LczamTLq6DgCm8JUVnxOhV5RQ/n78+LlZc8vV
9qLEL77da433MCO/MBJXMTHZhRGySLBhw0xgbafmB8ODwIIrXJgswV/Siv8wEelWH0Zy8kIM04eJ
Bw3LbRnSYrLA4jHbSWbUdLYtKlju2FfxtTv4xI4q26oaxi7gnLChISUESgkttWmJgCl1tOzJSFOA
kDJaAKExIOULTyw74U4uEfR103RkrY8Fpb38UxvAxOaE+XrtBK2D24MnC0UapYztvDf1pgAlwN0S
CE3KEacq8COI4gnrhB+vqyo0xsZU4wt5TairmiqP2aHXxRKLvybWBD4QjwGTk9wH4nYbarLNgbOu
49Gb5LnT7D/Q2Bg9VJtvJpu+fAbP88V5ID7pZcJZjCLbSWu8snG6GJDsf1TDJu5et7q305zUYdJW
fY+XYoOF/DnHI+Ecfloc9dpaej0vkPsj3cG+5Vbh8s4fVy9gzUeL8doTb5wn55YS7gIsEbFnUPbw
AaLIBIuax3fO2AfzNF9rBT9/Fe2NymwKM5xQpqBlRlmAyBFR2TvxwB53fiwcQjm4G90kZjgtAzzJ
mmWiT47CnIc9thfZr7B2FcG7HJlwuQKaqYCWQNTHUbxEHLKWsvZej6WmL6/khUWaFNUDObwf46Ti
1DDtWlOkkZQ+Kh7GTkTBtG6ce0ZjkgwHKPUPLiqIZDVX476d6eGwpPs8f3tm4nRwti4lkjS+Arkz
Dh4CLhV/1NX+3jFjf9bwl0GgrBd9xVwHnk+Uw2pN1ex5wr04b5zU6ris+J//3z85GZU4nf5tPBN7
ebPIYCVg/vRMQRSh39usrIZPogQHFcz7e6hThaog1nlUkpr213MAdyUHbcd5ZjEb1LUyI2nAJ4J9
LFstvU3Ov2q7KCgg5nd0AOCGzyiXueLHSkmhgBc4sWpky4OAx6nq5sVsFm3/aLytP+25ukVy70de
KQkHWRcdSaRfjOGYA9YKda2yFp65OJrpn1XjSKDWWEzalDyloQMGi3MRbV+ciGqliOp/m7j7COaF
oUU/LdNyrO4uah+p3h+Av5NlQWmYFDMUsUhG3V0XeBR5eqPE1HRicKqKRrla9zITnLvAxXHtp0W8
9o+0wDA8e6oASEuJQGqhtJFzJg75m4I3UTblD3+qAZ+h70rOf65eE1k/QfUx3UbikBdvxzemPtgT
g0kv7LBZHMejKkPjcnFhQkjQ4CuMxpoEGj6hRoz2hY4nTtdjyZJqQP1/3knf+leYW58O13/04r4H
S0QF50zUcOXVimEhE3NvX7KYAAdlaZnQp/NuTpZiFXKMHucNjtYN+YcOvwwP62WF8Ue5x8jmaXx/
Rv3KU3vHWOIdzZlJTxCBOFz2G1TzHkOX0rhYoF+A3JvZBn3Q8xlHHnYuSK+/nwen5MxQJIWSlO0O
Oqz7iq6HVBHxWGx3faCA5jlNBIeRecnu5j0Mtqy8+VcGP1r5jJduEB3qKItRCPVRKMo0ta4HdtDQ
bufZwR8m2EolQfujKD1VdZrwSvEcd7xN1lJLpXm5ErXTtvhUU4G9rbSVAcIUiBNxHmpU795I5619
Fi1G4U+QK9w9j+DPco8y5bYrNMi2AvzhmDdo8hDw5zJ7tTmAhRRSgTYvQMZCG+zvwdCWtj3cU6aL
2eBL/wxViny4lkpAJV5WXKAwU2QH/cVb7bH5M0/iMrk+Q6x/ktc8bY7bzm2hkZFJFHQSjXVS2otW
M91wvhIxUSRdqGaHTGzB+Uw37HpBZ+oBSRWRCCBytIVQ8N2mblxMl5tzn+gSdU3QQV1t07aTsu3b
jkqQ+CocmX1gTsroDkfLJXsnLegFXFNNQJXAzSNtA3sqNcA84yXfLw/s9BETscs4/uHBroRyjHHN
W38URjHkoOAJmwOgmrbIfkxmvDgTv/hjhEGXUKlQFMtHojwStmj7W4L//Ov2OcoZFsgMCwq4hLix
eVQAs2PPr77x4PgbBM1nlxfFS5W+mt0o2zDPDT7eAa/4Zym3MBh6t9AneAfmvS4pvBcSBMv3r7sW
eefggFH7xPC+Fsv8ETxqElYdfBHbI7Bpx57eqrRXcX8WGwsHmqFpVA0vLtaMpCMw5WCQ3ahshGU7
GtUaeLIXk1oe46V/8HdVBeUWjycP78cbchRHXts7eXhF555Z4ReNoGLbBqHPLZV558T6xtsZxf40
dQN7lPO+D+xMTB9tmI5Fo8FqW9XB0MEmxyhICeRdxQRqNx1WvlL+z9FER7NBeHe1tUrxUt5gy5sy
G+uVxf0Q8uo9lpdBxAnC/o0Pk5cFXzoU8C3yZv8tvRGEsUf01Bs7J5+pdYp+OQZONBn+tD0uE6u0
Na/Q1eaR3EXOBoQc6zKbeAueu3QbcYRgi6fO5YggNDRuZs8iUDb6qKWI4p1YcnJ0UDE9cNpZHrNh
u20Widks0Wlo23rQrnpt7UVh1o3TIi8AutfgijVt+8ImbNHEF+xVLzRrLBf5L8sJ1G57uy+9R1Nq
5J+ptM7ys1mJ0BEOiloiPoQ+pVxH9Xv70ncHKh3bU7KL3MtoeJVX0q/XdShsLO02loMbNW+IJ4Bu
h+/Mcs8+MKKv2HbBIBET/D0gP8LqfMeUHuSUcdJ2ZU01JZPzZLGGSMAFPWfmmP+feZpueh0uY5CC
pep9ob/INZKyknpuIUIHDXTcJQrZNIkRhjt0WLvltvomgps15wvYewgmtdhv24/xrrHrbRyFzjL1
sJwjv5PZ+/Z00xyvTMkFP/SWIc2lNPjMjRMZiuD+j4v7Q++NFn2ibijpwHIjIiRjzB7o1J5ORYiD
lnp5NziWRYbzc2bkMFGnWIdaqPw8sf29303T+3/vmkZSF7bHcr09HT2thOVMM52wklIc5swkAmRP
KOL6EzQndwJcpPkcIdHfB/7xSUi9jvWr7XOXuafHtJMQHvKhpT4/0M0ULz0OI6jzNL7Ve68VNZ/B
qf3LZ5wQOh+0DCIwoUp8BXqo3Ri+EAyT45DTymdqNi2K0PGSXlKvrnqJIdCwzeInOVUXe94qegD7
mpg4W/WkHPGuZchzA3xVfON3W5IYh2uhvAMJ+nps2A2ffCHYV/2eX6+LpLC5e2MFNHpxPbzgpois
T0DsPdgZue3temOw/YqF6stfLj1LEnLzBcRvkf0Xo85wxrHjQnzP5/Qr+E9CaHYZycWiAI7ZB53G
rayIyyS4e0n+qkIxVw5ROkZqZtr40xr/3m/Id+nFIj2SjjCl/HUSvLGKiCNkhEDFJYATm8rT/Qtg
CnQX57/VUC5Hvz5rdy5Tf4Vnis0M0YwKgK3D032PhDFfU+XYRZHwshRxDbqum4receN20GjSLPOA
Wl2KIksRQrkHAVVfW3sqStJ+NpXybf2B51r5UgblAknkcmw6/WfafQv8mgNJPIFHG6Izv6/UAGGb
NuO00wQnuyxAtcbHCLJNKb90PMCGjwNSEAViK9p1/RVTHmr8bqZo6Yh/JD2FdWnTvupoZbuha23S
+H76rjx2dQczUIyHOjboHlp/7BtLb5Bk6+SAjMvAdbwUos9Yo0zqXowhl9G05ChdT+YGcCiQ3tMC
B/08y72snsVpXAW3CTkjuRhs82VAVNbzS30rEL/ulrsbYEA7c7qffMSKwbusCkWz24GrIfkfBVsP
GZ5F+mojzgpPiLi1YwEeEWB/HcWOv87NzdoTVwl1KQOWllpT6cN5DL3daCqv5Hv49zHmibn7deFo
+MUrIQQ6JBBDMdmR4zQyj2kd2JtdwXohvWaagP+JPYdua9qV6GAWOWiEZhrZASs0SeWax21s+te1
xXrcfalN3m5rL+v3ec0UKfvlVZcyJD5XS0z2f8QQV/F5XY25szgv60qFhWETtDM0X1kYKDXnTUtO
mNo/hoi/axcZS6qe5pRm36mwrM7hoEnG5eT6nJewlH5Go59yb7L2nYh26UmD2j9oXIhdoyHCxrU8
pASIuDHNxxrGv77UO8gi6bN9QuzEQ2l+JH2daaZaZpyAjPl9pHyyU9Mi9oGMWnwo+OKMvoNAzpfV
x2l9GhYJf7bcodrikJVe/8UeCUSjwSEdJS6bQ+YbmMm5ZR4QUEO0lu/Mq/O7NQ1KZ9i3WeEMZ0Xi
d+vL6Ts4/hxD+EOx6uhhOQJcUDAjErd129FipnVVk0hRNh4Ppg5CZ+iLm9llDvh1u9nxYAhlmaR1
5bGCIZBrYPwNSVLfnLzGl/vIDlcCr5fiozW1YV+yVgq30bBbK2YPJIqHk9vaRr26fJbHbmv7e5EG
VKLNtocklVEJuQmhz5CEm8E/bSJwld8OtSqnXhByjF1nS0hNy02CJnNfnFuNMzIZHnAAj+ComvNd
pe77czt2cvXMl/gPGrAvDLgLKiN1mI6YEg5jOHyavZAtspfLDo2Ff+QM4hjMPQaAIR15K9eQuJHC
C9TFe9j8MmAFWzD0fmK/PIweQHd3kEXdbckw+3IzRVGdoxwTsiLIm//HwkkGNcKPM7ozWZK+TXFX
oSN2mh6U91Xs83dvbhDw8uhUrAlcr3LpgCsO5ei10mnKXph7Q7x4EKgtM3lxyAaY4cXmlqtQ/Gcx
Fr6FRbEux0veVqn/GZwNOpV7q5QZzuPV3V5D+kX60BKUOSg+6woFpOPu94tIglXaZSUTfsXFsFj+
SSPk6qtTVfIDA7UEurhd1qK0tjlRYESAbl+kcoEpwzGEfZJ8IXmKz0dgIo1WNzP60O7ct8uUbe6c
1kbJtXzqpXe9rSkIeH1VyXvoFGhGzhfMOktooPb+QRWihUge+aICGq7Ca5/0kAu5IcJlfSZzrWRU
w90TxEGTEi40EcGPNh5wnUaxKwaIv53NGV3wsM7bo9WbM3XoAsHnSInmlEp8b3ItGDDYiMaGYoSw
Smx5Y8Zz14R1qV1In6f2Kk4PCG/SRbJg/VTjcuSZNioRdnc0/88YiRfQxzWLRJU9Y40Bu2nbL007
9Y1pmdIcZinrahWF/3ImqWfqzMKMOKy/X/3my7cGiDroI7T3sTNdWPNtqcly16MY0aUCvAW1+W8q
2UuvqLpocbv9/qHVuvOknsm8iuBHZVZbMsQcT+7Xf/S6PDxuvAWv1tt4WsKHqcJQo2czxm0WRg/0
3T0GxjfUjNjLnilrhCWKw2zlNf3EQzoIXJnzASdWVlfHge9bBPhEYtgC3UFyzGBXopKhYtzV5+Ep
WQb9vBuyMvGfaWXJKNBbG3yn5H/VhFqBr9aDsiz+Jy+aTnbrbV9fPPFKi8ZI2ajBRawvFDMbFCnr
6Mtli/e+bGlBz5bNqRiDRhjxwYNh9uk/JYvBkKTzslh9MVbFq11a5lLG5syDVpOb8IeMWmAAUVVC
bpm55U3pel72euQMh3Ock/reT8hEr0xfI8JPjeT2Ix8+D7wJvObFjM1R54Q8zeDDbJIWm02RAyii
tXe1Y/ng10mRw2f4fRde7PPfv+m8BBPKJ50lDHGQCWWZ9hS5lZ2jgUhZuXqLr40FQOeK6Gbv1ONH
ZMTvwH0vyU0wDJCIlUZzi2RUNfl4vU+MjbN6tEYK9fPfF6105vzZn63RKvEpbRIERADLpDtDRo6C
zafteyuTp0XFXN94pAx3rSCjEyRzjDIxDK3EjP4v8zDR1wLTeeLZ37g19UfJ5eVr9r7QtCbYZXVE
MoodwVIHSXlRo7bxtnPY6Zd4c6MWOsjsQYYtP3HBhnrJVrsdhzNKSUd1eESa/yOHgb6bt6k4KCxT
tC7/hU0q9SNff7L5JhDrD/BTYpJvdB7rcloTXY70eNN6+dAjSBh+bNsLHnGTjYXxD4uUewQtk5FA
vTHHlYTa/UcUmMfcp9A7ohZ7xh+Q/HGHnOje5YOFgXDkivR4f6CwQaiKhN7TW/1JRbrQh2Mx0FOD
36e/67v5PKDVPRTVenCXDn+DjMLsPSQcBtmqwIiCPGLnBEprH5kWlVMYmBEweavXAqkA8Z1sadmW
lghTIdtMoHl/2HI6UFeID6XIEejBFM4pDkXhHVIZg/Keo87Rfp2OepAVZ3Vosfq6c6bi30q55yoL
uXdiIUynBjA0uly9HzaDc2V/Oum46iem9CQfGRgI3RbX1n38wA/XUuXx64/RV04I50bCYtDtFqlL
iKAXSh/vBFcrhUL3Z5AyJl0O0LFkmejZitZlY2FMwVg3OYdl1EnlRv7kojtPbPl/U5Oj8aCnKxXt
+e8X+Xnzxn424Y95+Ud+e4bAGETAwl0sAAKoK35DSMyhpnwjqHaOKe0x+XqGk2hyaViV3ZR4rwVJ
WxMc4qwAC6FuJF/Qid25DsWponYlg7bShwg8NqOSu2upHdujliI1KSpFVFpib3xRq8frAJkgkMnc
cRy3qfY90oYQu/bQZol2dYPTJd7XkdJlaWR14me0DPMv1oy6B6Q8zTE6t7/64CgFSIGZLTzIBuXj
mUVcKyukOs7KJ3cmR7I8Xc3YaaiQLoFoxA3EbO4yjtuN7ZYolN0dJuLfy0bEMxEE+Oon9AuKWZ2W
74lWp3+wfXSTTW3QQIZNg6caShg8aCC705oSiWqerwHurDAEeMFqh5V7oee7pQbSm2FYClP1d3ET
8DFkoOdme+ojNDWs3JOedTVPk2fYrn0HJgy/cWZR+k4BYIXV6IW46QSWp+JBux2kjwMXq0RMMJld
0hw9vvAaspdVueNz1S3Lsd7o/D+ySp1lR/uB3MvCyINTsPH/XQ0+i3x8X+/iF3z62ED/UTUVj4b/
rPRP4Hurq4ykOahEE2y0LMOs+eFUgh3CABo6B81T1uMcG9i+0O4wH8aJiY243TsjoiyN72Tz/3l1
4M78ngChuHOQJgNfEWk1V2EIrdqv+2/xjB3kJ46F4LsR9KRizo/UFJx9faMRvGo2Ar+LKTmk9SFP
J/unD/cfhZZmW35gro3FlrCPrC1ha616Nl8cs2Uplp8TRDY49OIIcA302I9PLDOvn+MQruT49eA4
ZXdbBPCYuC8fx0RVeCmN9Orv2INt52W6gLTp4OPlFgQJp+aJG7JPeJIE+1ShlD4IOqH/7YmnTIJF
spYbGdWDmknocLH53XnOyUKqVMKcPArr9kKYHJaLlwSNLu3sqhSqjIra6csZdBWB8hXI/ElcmXSK
j+fjrSZhfUV/8HuFv7fW1C9NzUIb/GM3zJe3Z4ZTBRHh3b6Ph3Hn0KAu84UiaL+uJQdFa6cVhIb8
Pi/diDoIFGuxa5Xx0XZaXJ+ciqtR1cbYPk1EbcLX1GvzcDV0rYu+9SRPkvVR/aR+nrVYvg+G6xR8
A0A+z+Z71B8E5uKLxpPBXV46cuLTXEXpIv2poZkf99FGKmnI2JIeEyRxPFlnlnqVqrdLwnj+bqgT
Lo9CxwuVu9NL+ZHwjFenxqokdY++CeedvRjeWLJuPhFVRgKhk1OtyAC2PEc5d9NkRA/pLlHYLpLC
6f40sxMWS/hpXSw3Dw4M0DeElTefyOwJxte1AAADYyHrUs7OvGQIuUWpYDtwSkh836uPKt2kAXn/
lb5ND0z5SmrHb4mp+hwJzGIbi35soaJIBywY+650JHKlxJeCFSvFutu90X1xOQfrfRWpmOiYBErG
9aGncqc7UKDIjStNHwtYgqrCg0oEvIZ+qHoBH8s/9NczXeEeeOe3kQvoXldpjX6/yoXXunwvhZdY
Mt80nWpdf6t/eMHU5tZkz6xlJuKn504EOFdy2dnRTIC9YqiZO8ai2+4ZGRYf5796CBq5HkShthb+
cdBVy1aU7qw0vVpTmSxete7kIFE71rdSIPRYsTo7sXtrZfp0xodDfSu0zZGEfEYag+VyJMIoD60E
Dz8cHB4zQlFKxt6Vc8W9xebh5OHjwWJFC+P+TYD/Ly1uwtLN3EZQlFI7nAISDfIAeAgQVTP2b0Bh
UGWYO5I2czNWQvh2ezY6fhAHH1b6Xk1Y3k2jFCGDjjwfVZXQpDY3/Ik87+aSJlSDt2hlgFDbiGwL
ajk1csmEM74cxMZ6iDYAvAMDjlCRNQkb//PQBCny8tMfdkuzJOWkyHnng8APMaFNmQstmQb+Ir28
NKMxHMQ4L+pXxHJHDxvmZd1L5ov67Y3J2Jv2UM3j0oYRYp4GX5pdMaB1aqnqDUHh22SFPr/e2D+y
YGoIvHgQL0t8KRBww3x3wgYWXNRY1IfZxXsF16xC7pUT/KfbvYpCTxRfMdnFa6MGeu3SnmxFBu74
tpTbG4YyHQ1Y4r8BTQhxcyVdyvzv2ZWhYAVmiJynFPMEUDd0m825wQIiA4X+9B7pIao/u9a4j80c
d7oA32NuCktn++G0hAjNoFQdaUkzy00U3CM3Z52dzw2oq5ADAp54di1Thog3pmhx4105fEdrOw7z
PGhF36ZIhwQxPuY4jWqRT8+K2vh0j94ez/gUxzFqjCSn97bdkyQd5Y9lWJXTUqqpc9KRWRP3TdGX
sw+XUqtESDEUyXAJjXkczK1lKX7GjUXKRTy8sYmAOjSZWePTus46dfe0fL0cGdoZ2DAoY2FEVKee
z0Q+PEdTFJTEunrjjam+/5unH5Di73Xg79ydk8zUA92DJfmdvsdjJs3jdfPBEd43opB+tyWALY3X
GszPLYGwo3LdOlBGrL5DZFPoDVfcbXwpt9ThZYMqfdxTHyYOCFpjSf1hOBdxm5hoU+gFGHgLM0Wk
Fr9rl6SnJFC+41xO6enpu+XD6Kp1U10CnTonZJxvLiZRYfEK0clhf+Ac3GUpf2rUWG7gVx5cbdXw
upr224BXdIWKqu9k2g6Y1tu7dZ7OOFE/vrIZgv3Lq9qkwTI8JOoMV1uzzK+s5+g7t/GJ7grswwL9
nRxmjZX+OYzvGW/AVS0kB9QOUWB2cm201DGRjVqt+ze9w1C4XymUF//OZ7x2v+rfo3y3a2rOY0nX
J5lcbh1JVj0FSvx8TA8CQHPpe6ni6RrIYeUaCjPGoAzEdWjAc4uFQH1xfqE40pUIkZv/6t9IE0OL
Pq2NIwUa3elW3bVkr31qrJoIx7USnAk4/F58oW03EEhcIv/F+koNLRGxNX9enkiEZO4eiOiWUzdy
HotC18K/psx71Zu4Ln7TAV5TGOr66TdUdfMhdfdiqK6fgZ7Gs7PUpGvwSVLjHIqhxTUd7GwfncaG
6AW1fpAXww1wv6NvopwP0YKW4ZYyM9OIjNuakwGM9w8t/F5Ljq5JLiqdXFcaG+RparGVtOJrn7Hf
t+1IsSL5g8w4Pc0CymCjJc8vGOflRffaOu0wC+YnJsJ2wo56qbelY6aG+cckl8ayPkDnIg9iLQok
8XrmGo/8wMW5qnC0/cM67YhMF/eMswYouwoU/CTXek4/oIMlyGs00zZE+yvHCOveGvToo7H+RaEG
Juqq1I6PxTLTR5nP+8FvobzF+YPv+XAHoZ3664/WJ9oDb5h+hSk8JU3G7XlJDHxEnLc9fWTbXE+E
UNXYGZ9/cQdTKAFmy3ZqALGRDq3IqR3DAEFluEKDovW7VuZDX12gSxpvO5xDm0+vJgDQQySLumF9
Z1lRZm9/JD11QeGxDkjBH7KDiygrwB1tRKjxuhqIz92TEY3oxGRAG4HRkmVaDNW2CYS6wdYmQXKH
D2Rtv46sxDSbCW3o2yK6XYBGJveJwBSlT85czh13TWLzlPwlf5ILS72ypiD37DESXR308J0HHUmP
hTwDL3Ka7uOi+0M6EfSfDx+Q0P0cIFZsDlYpsCT4eEmqihPzni8b8h6xkzgQZ3k4SzyqR0QATNmW
52IqSBH/vXVXwL+HIEWIlkQqn9OzLvLPYJ8csNpgHdhEp98tjlKNvEIOPb/d9+jWnHD6ZY6SCyNA
gcnRDMes1p0bR0CJ8o8fKlAU2lSeWc2na/ve+3WSEveq0/oeWFjbZI1L436hlreuLkcWlKEXEkZt
shXsKtnOpFZC/p8DkEtxMYLgXg4n1OyK2jmL2C22qZoc5VxSzHlnRKZIg085ku48T5PUZY87Kfcb
vIfi3mS9sVVzAW64mfh5h0FEyEAu2/zsPLTyzDrGNESQSdfuMP+uOoYa434ktdv74t9fPK8gkE2B
ny/1rqUXVLYbH7lhPMr30M6hsV5+MdagQ3P9VfB/GuQp4PH1WtpM3r9jPMe36aGQYCvL+8urE834
3sPo7awkO5v3RE9HkaV3ZelAqJkIIFgn/bffOpeBm0axtoh5ZOWg0R5hyeaCacAcZtczilR8/CCz
7cGrXa+nlIFsTHDnxvgTJKxRAHfC/JxxjPtdG+B08wJSmYBtkw6K1pRvucG/FDMRW4Pg+ThI/b4f
eEeB7JOMMztZ1RxHzLGVzlW5q5CMOj2W7sHmSW4tm0eWmU3Rmg1VqvHZv0E9IMW50xV/74eqZ5Fo
xHC6f10kOyX95eiM0oIv8fU8Y+FTYYNpxZAdxXIKgHm+kV4WL4nIADlbtBvvTzzzzoz8h19OExoI
2xgZWFmoUdqfWnYnziLRaU/c0b00Mvh97nWwsV/EsW2wXhxD5y+feNcD8fpn3y8qyfXBczfkLRxa
tThl66kDFWxsxhRPhdzgsHXnumCUbai/b+7oASMMbY2t6OhxPTWeLeWBsPpdwFRfoTCg/ZXRCZF+
e0NRrfk5Dlkqa+t5mgZ/HgjCdNZN4IeAiGO2SoKUMiSsG6TLUMRYv8qSyao42l1b5C5q/f1xOpJt
YwNkzdqV+rTWa16OqAEyM2SYLPjtJocwXdzPP9IxnM+XZ5AUU7H35E0p/K2rwcwi69fwdni+j1mw
XC4oOF7bG9EbzvbdgHy9pEq+J9pOWD0cnZZCKrAnwNCxf7FnVkIqcOARbM9t+8m826PSFIBIwIZq
pqseWF/sKTdNWniJyVjT/v3odONo+7FRa+2mfk0rwQwme5EM2Rik9/mhtQKRbXqNWMFKCpn2f7dK
ExchFzTJnpT5s3dOXuAxmeD4cvjgVOOspUcqTIqVrmD1EQo8l9+En7L8hwgQ5VEZHZUttFB0S6Ub
f68YxJNBZAbiZ52X78wqTtRE6zRX1xg9NyfsP1safysnvJNDirpElnRipXOdMq//Sy/9qQLUxEl8
YFKuGiPluE1mIWDEZggHy0Q5Oo+4X/+E9zcG7M5OXM9Fk+GADBRqNnuZD5hkbsnvwEPqax99ddrt
UeEd+Ma1zOnKyhJsF1fmgk7H8p3IgIhnbuGiefoqMjoLx7DulkAssrVTDKPV9LQMCxCio9HvKAN6
VQsg71LT+uGHmNNhsz4G4fb6gx52vqa/OiRkyn35xRMsorNyT798uIvqBuvG9PKSlZnz85TJCsSm
5MWh3VbJoiMOC1NHeC8xYzwkZFwshcLBRIzUpxoT0XpKw4Tiy1/760n3OmnMUXLeWzvWCfK3s/E0
tGBa/H3Etu9AotqL3FKa2JzkR2C4SEmZM0ESDe6cuW4EBDSuraOPtBBq40QkSJUZKiGQBB74qgcu
uaAJRFPl1JoVMeMddqnqXjwH8u9N2pVk56ttXVN/avUBbZ9P2YeJvaqkY0d7gubhtiNVa5sHWllG
Ayo/8eGIapNEatKtzxmDhdWg/jmqlGL9WK3FxumIGlWqieOK4RRptHmpjqsIUgwzy6swW2P/hz5d
SjybAUJEM4/66FCepKmoAid7ouS5C+MZzYEchxn6QS2avrM8E25LiruNyerkoW5qHqAzkMRF36If
oPxqr5d9VGmmbTH+p0Tj0+zq/0ZDcZIDEkC5STILfstXvoy0Alxwgmw5B9/qjoMN5w+VjZ+H6L9d
uKlRLUmIfo5htaux4NA3pFs8iW+5piaTnrX5fND/qweD0gRyrzu3//w+lLL+O8eyqd8VjoJcjgo+
yNKeEjV5hJSLSCDqBSm2YIXUBpWuktPo3frIcRjhhT11UuvcgXHCqTYFtaK+4Sp5uwuGt6YWmgIL
swVxSN8EPcIgpQfCecUdHWbbMhGzUH46JX6F6tpKFjARC6Jy3LhrbHAo0dmYg682b8p5+BDsyLG9
RbuC/9xxwCjnhBLYxJJgbH5QXHCD+jw3qLRVB6e+r5GQvp31sNKFYiwqneh+FM3AYarQyTmIC5Pk
vOp/D/fXYvb3hEru31/nRuBVLxEE6Cgk9qPgQljfpKhbiB+DUAey1cE9KrnOjnkPRgxzuQ11XTCL
YL/EhBQ6IsTyErqBlNsvHtEnE1VKoStY8HSyEL8gfIRWWsSbksku3caEwDQD+ufYq9Qzmy59iaOy
+31I0bvuTuN37hDmouR2jEZTWztzMj0w0UwvOSsed3RB3n+CBDwiAJlnq5dynfVTl2vuyzLqm7JU
3BqWlJyQT+OWa+dBXss+s4rrFqRH+bB2bZybPwYemaF2AY9coSTfEcIcY9dSoGEDb+UleMvKw4cT
c10t6zMXn0b101YFqzxjysGMfWztt9bpV4XFj3Tr/7XE7zLV75tWTJt53SRGO+CyyoWRjoAUyNCS
EQgMgfY9n0uBKG9N9UC0cKYCmTfOxf7cDhgL8RQy6NsJWjozE1daeS40Ttc5+NdMySrzGnKN1Uu8
NgQS7vTbWsMEt5o/B6AYSOnqyoVZ9sX1RSp1zCHisL3WFsolm7DPQQJHwCrDiXjDE9JQLO/i3gxC
c8YaLKQTtGDqzdQkmDzhtidHRnAm+GL0IBY/KqOGpuSoY99wiBOsbYeXimLyFl0pPGIIC60XTl7m
iAB3BLcr9BgeE4fWN1FT5X3J8O1Q8202ZG/FwPcrAXTM51aBhJ9BuwcXQH3IPi0VfPX2+29suCGs
cIUWamYLcrt7TjKup0BcDKQAV9lODbxOCKBf45GQTkq4B+EIcS+ha7GG9eC+Hd5Veiqnf6Vk+sIt
Eolbxx6+zaOePsCw+voL27wMLKjqLN0KbWf9RgMAZrKzDPKfXTkhVjAijSYphjXaEHjZtUMO6T3H
Rc7/kJqgTWJM1it9u2OP62dswskkcZMMhLY5HQQQEy/t/iMg45QsiLP7XrdRJXwYA2Vx4ssYcG2w
r9qNazKyowhRb8d11DU6TN5r+MwWfoEimmddJ9x2mNDP07qQpbb0bOdM+QJfb333FIQDrbZrh07j
HKB7iNxn8i+CndSHNOimjvyyNYip2Ns2Xs07Kj1hZcRtk6hCa9D/esjK/EIt0CIxKzLNMVa3yZS6
u1Q84HBxj2bcn1S7kTuP19ehpigWIGtt+dr8a1i/DUUFUlRhF44uGDrtIirQOp4zNFdFlDxAKNf+
NXNchfWMr9Q0n2e/FkP2r9ZMrsAjKwQkM3kfe7IAls/kgE9AYHM7a3cJGWxiB5rDXiXfbprGHpoU
XVCwcND9RhxqA5xL9cAXwKo7j4LDgzIZSMqvg0NnPgPLRr7/0YcVW57FmMWRtgpEb5v/pjWHRG9e
1vO6noITG4+joOynwAOSUpfxmcq8ze1Bce/zi8gfKCbQt06KKgCJYrccdt4RDyD9t3i4THZieDP5
6MiTRd/xDgTfJY4Yc1K9j2X/wk0DWzmSyuvElt81EMM6/A80u56U9A6T+9iZBRXnlZaIZy6MrIOs
U5eUtSzsNPhr1YVGVcBi8pWDhA2C3DvxyzAFIVRnoDAlkEN2o3RqJvJiki+vK0TiyymLDQqhZbNW
E5C0Y/8nWh4d9diHHjEhJklg5TX+Sm0rfbfxNUb3+hcXUu/tZOME8y0DTHbELaa+K4mgcLnrTOM8
31izSW3vdKYzzj+yFJfew6OOzNF9ZX/BWD0+is1+5C8lJVLGd48hwfD1gJshkWiLljJUTvGyn8uT
/1ctaOET/d96mWkIw1SoZn/qTIAFkboA3kvOVga81v1cgZtS7ZCSc5Nx3WVMOa06c/9OsvkRfHhc
pAC1jdNoWZ07mNItl0/iBzjV0yLNeetXPxmYQmVPLTGlZ4CtbXJ//tRTMsbivi+5QMb8bbKYiSfL
B7P6Rkle0ycXfrUyzqQvlKnMRiz+WF4XiI7sjtwiiG1pTzkDn02kEaHi66VLUL/zxZACDwyrAyB9
eLyNREG756wXuFGo/yB4ixqlq96JnigIhSdDOf4ZTgVelK/r7qvuHmBNKna7REnKUDH94cUnidIs
O5EX/dQnC90Prqnbak1mQKbr2EN4NT7bLYaL0zvNOB+uQelC84bWjdxIKkbUUe8qdLaO1DQI6rtg
t0mzbPerOhiVA+itsgTEhhNXmMxOTLUpL8usF2X8LOnlR5omjplj81Lejma3fp5I8B4jCm1i2Jns
5Hj9m3uds4u5c29oFHlPeHbPkXGj/gLyiT0ARiUbDgq9tZJ5lgfz33KtMzRNj2e6w1TfhuTRTrXL
olxNe19fxpL+YKQkGDvBBnoJpnj0TRmG8CH7QzOFnrs8z+PQ5zuKFMmylxgyZgHQMIdSoxYKIvYx
m0gf52qSNoshih8yUKW6N9KyFtsMTlhvxCZFAirCOkYUe1EPrMkcitklrtGFMexImWBkP3B4KBRR
uotLgqCvYUuZySpwb0sjtJeCNSoVq9qlvup7hmabUy7xHgsoKYSg25gTQIyGd/NRXK/y2P+MMA99
EeKnI1sicHckOe4+3ySe+8QnNNOJbc0c5iuHCo1s9ds9bmeSYG1JaUa74gmOw2CIWCOrExF3VFeQ
K2ha1ovcJaNJmIcibJONf9CEpjaA0M+qya0PQVEfRO+mnVa1ZwASaP14xt4+sEdsrHeTo0EPxDBd
e/MzkcFYij0pCGCQTUVMyuRs5rYgd8NKtqP3Hr7AJqz2OZUbi1a6GIw6u3vDkMJcUjcRnlwV/KFQ
l6rbPc+csZSsUnJnXjyJlii7OJHnPyHaULw7UZVzNCvPQnFg9RXMSjQ5RAjKJGRHMIanprFsfkI/
Lh4jVNBHAdWpXcwdflPZARaAfdPln8vm9ublyF66mB4vA74Ax9G6YHTcSnn+IsNfolAjqpsUY/+x
lQ7kpir91EXRxEwO9s7zywh6lkF82wjudmFfXBelyMXba1+b2+S3Mw9P+6rnfOpQLXmHzWCgkX6c
7a0TzBernlR0j4dmQrmhqsBCFDs68HKyXySzxUSF4CHTpJLnbh16aybKzR3R1c0yueu940z/euXg
f6gzmWlFDA6rPPsWiCqfYsldZSEcJyQeQno/RX1yZ28Zfw0nCruS3XJwabaCdGJhc1Cdis9wS/Gy
O3aFERpUWUV4oOwlm4NK9wQQmPuGX4Rih8csQoM7scES4sKD0KTa2mCBrd0U/iZqLX9sJhc2HDcP
e+YB0irS1WKz5yC4SFCAmzpYt6goIcuocrdD6eng87pACwmcdD4QF8fk27J3wmH9wtNkDybf9S6t
NiASNd5U1cIDLRs032L74DmetXXFrqvyvuMfWtAXl54lga54sUmTeCqVq4j2PZdTLCmvQwLR932S
SyQNKHCYlqIJcuNWcj3tdiaxDBZbdeJFFuNfoOf0UTP5i+FbtwIdXUKXuspYUnJUNnm4i7+N8gBz
pIC4ozJrzdQrtFG4ltp4p5H0mHFuF5ZWQh2aPErrfHB1xG1wq7HdmNRUVVoK3e7pxU+Y8Zo5Hacz
0XA/EeNaNyg6V8qHZWo8hFHn/KKGYLPbHWZfRe9IYZP+s6DAmEY++4j7J+ZKASvUfx40589EpZ2f
jENJNAdgoe4tt5+DCkmisEbPAwjU0UTQljktpT1AAl3weP8ihTglFxtH37sfCXE/nZ8tP15sIypW
eMv0FBHazefXvaRzfJ22LuO8bNX12ArxE4LTwUHo1fuPVPPwL4Sa8VL9e0+Jd54Ud+mlJNtUqCBb
pw4HZVx7f6zzS8nCg5prSRmDkUbkLHMbiOn3zjxFkjRQpT26d6fblzbWD/h7BzkjKm/xqmQGQyDF
+uWZ8O0Borz8q6sccCqQ7ZuE2znZ5uYhS64o/oKNKHb+MIkiZXpUgEtUGTFz2j52MHhVEw6zByFi
T3Jt53dME8RQwrOwlNZLI7vuSi8LCkLxMX4jq8Q2yDvk0e3WATRIIGlvZTabWKYyEcELlJa0bjlC
J+igGp4pEVhab0PD5if8trOhTbf20dgneCdMFPSxaPXx9dOwofuy2qjotoLMQVQQ3vwL3auijFku
DlpV+TeimjFCoFkOQv0zcI3G37n5+E9cVwsU4CMg+1QpFLVHQRajkZGERckUNFZLsLZ/r7g442t5
bfaPACb5FZ64GN77ufVnBxa5sKWpnSaXg3uTr45I6vsb+CVUFBPEB1rzZz5+AEP5u1aCnk0KqrHW
KlZisV04HBUUZd0A4wAKLLMLUtoY+6SsKkej+qCr8gLbMQOCyjOln3+vPs1goy5CFkY+uVAh/4/C
KFgLtYhJsFw8NUi3/Ila9byxCbVya44+0UM7QRLw/zn8DEpgjp2UkPDPH6EEybPvPwZXcBZZidbQ
tCED6XTy1RyUNUtkUj2AvVgHFOaHfMFi2wS9/WzcCYHy0cUuMmgqFIo88TGInb28fPl/oc1hb1RE
TFXyvDauKS2Wchp3IwYLQjK94exafYSxP8Z2gidKMLuob1w9T1YPP5SCtqQ1RSkdZhnjFsTYMiJW
u6YTGxJUkWpnXuBbr1OJuaAHPYtycAxOq+mGbah2UEK7SVc+DLBsm3gp2erghQedXsPMWnhwSU2f
3xVMhoMn3/Hs1Twst8An8GcTjMYMVJQcnHDEsNxAZe76RumPrm7l+qIMLwYcicfWYO7tOPpAOU9D
aOv86R3Teks6nHRAdYUt9RyYKwjVBquL3TXCzPG6TrPP5o1OtVy2UKcNZJQJ0wjaqBukIC2U0tTt
1lWDxYs/Q63uer0tPR3Dds/GYynBuo3oUtlw2AeblxrUKKzGTzMjzaNAfCm1yTuGGuvKPmZpPrCl
0+nDEUX1UWevPT0og7Tree75V4Hu2A+sCK9aim/j8zuMQfEz30O2EH75kWT0k1dwx97rz2WqoxwG
PYRtetbi21us4fDuxHNpCD8Fxmkt73JaF6GYR2Jx6QbaUIW1sE/4yFcy5Xi4LeCg5F70YqMuGjLl
qXG6425PlZpDeCAufqHs+b12WfQkp9EewKh6MMQ3O3lz//qgkb6ClxSQ1s7P52QelPN+Lxyp48HF
2TDxmIau066n9AXFLBGaRz+sZVjZVXbzkIE+/jLIZp+m9uYKwpnVQwtP6Ofe7SRXO2xGbPprHm0t
wIAXFnQqU3J6aTv2xgryzh7GN0apBGkvKXBXUUtOJeReMeSHcoC4EGthK6GiDDk1x0qW5r/NDMnC
U3d1uKbpV35OKTm9CUKhC6CeTgqBzfRY0x/SRgxAIfc1YK7HARluM0ImPhtUqKsZCSWTv+G7GZHU
LFz1oWAApPpQUHonpq9SxVdJz2S7EsDMmZpcpO8wxxf6OG9Sg+ADsRCke8EBgimEP64D5MY1FeeC
SjPz12kmBAg5I4UG1QDWM9bp3KeKjcqtTPAHjonzUpYKjYgfENE/2kIFnObUy7lkYM5/+ImKBtc1
S+h78GloA5rAna8vIni+70MjA0QFhmxAnl1OaXxu8JvYMFQYLRMpjNO9EN5lwAr8X5SgF0ImRfNZ
5qnq7AxgsCkSrMCDUxA2sPadXD3QGtpValpg812LgLKNi1qRA4Uxh7+gjxWgIRNzMaXaaiJsjOHh
b5fz4NTFVAjkIEt4o/b2V2Aujg+aHsBVkbV49ZMK4BPH0KZNah6wifQOCGi90gVc/dsgcJMG5tbI
1h8oDdKPNyteptSy5h/d8yaoA1fM2I7W+wZUrBZZUnB4x01OgNcWL/oqLrfHbkK3zRfzD0A9DMX/
WmobuauFpEfLtClKKS+qQfIMa7KCA+ZS17rzNT6XzyWk/ddmnSF8t2GD+iNt7nfIJ1LM9QlESa7f
jeRtI4cYySnr3qGp7JVIC+npfZ+Z/qd28z4YiTm1liiGa/yr1+WyKgtAlS57rjR3kfXrXrHip0ED
LhU6ssb/f6oB8yaXAscTMjsMBX4gUl1+cL93Wbya/c1s7SBrgfNGvrkWOhPRofvEeNpWdcfBDea9
KGjOGBWBZL1sQxjP3wzo1dxyFdikNzA6+WhhoZg0WatUlpON2N2KwF5sbp235U1JDzFqCWSe9mdz
TH8QCqFwdetdJ5RsoQ5Wu9f7gASq7DYqN0ABw9l7EvNyjn6NJ/6lyvIUAHwQT1d4Z8IwSYhFyhT3
JEvQdcGm1rGn4b4N/VEZUPZ/bTTEaTa9SAt+7Ki6WU0xMOoN/Me8KbfvE6FE+aNrTSASekEdRZ+1
s17S7dU2N8TwRaCa+KWS+zGJJ7fwcmi+EfvxesRFJrkEdg1mumZCEX3SXKAkMpncIpHFrGJ7q3EH
MYlBaj97Y40bAyIfB8X9o4FR0e5Q3zGevBRf6jiyE+1QjzE1aHjUGgizO228jjpvI4pmo552hIyv
YfHOYTWTm7FgQ436IuBKXKr2Aq/HLT5R1sGGBdT38nR+522vJdPJSVEr9t0TVr07c8URC1qKtOOF
f3G250RBNFn++7C/SrEww1PRMj9sdG3AhjysVU/Ro5xoDMosOIVkjtAOPquD3DhFXMTHA904aup/
357rM5PkijKVHiHrWkJUYZi+jLPHGmOmMI7b763dBlKMiN8kJA2o9o+hSnsZLgoP+Y2YUFyH9HnD
ZRQl5m3e3Z5b9K4J9ZoiQ+sUfDOYFpFwGH3qCsfFdrGK8eeDv4xCGwQjCjS82br6oCzGt5P9pkwQ
WWLseTtAZpsBkaxyio/AGcBc9N2Uyp1DxBN1j1BToLWzpwfYI95z8us+eiHshyIvX6oPatsNwFBk
hkxmksE7/A5E+/JqQnmE5aWsCStBqIWGMDTuIa9aSFRn/5EnNwUJvxT5nPioXarHkDUSiglJ3ajy
XKyUXGRd9dkGipRjSCWSIUDD5SefiEzgErcqdvA4N5M8Zg5Rf0h8m111+Dlm2r6dAlOMdmEtmPid
HBSdM7a/diW7mOnkvI/IqTGCBHv7BK550VD03TFjrTrVcab+kUbRbxesY/zU16m3N3hx57cdrFyu
fGcwjlBu83aWcFplOkKl1xDxdkpyjYNdf5rXjrFx4Jk4/1VPo1qpN3jDiqdlRVB0LDxgIa9A93Lw
lfJQIcxYVG1Dw2DrGZSiczG2wi3Tbg7la+5THuK7iF+mOCRNvqi/9QCI9m8NG45c5VnI7uVASGfu
80tzDlk7ucb6x4m7X6G7kIwIYE/EaVHApS+vZcbdmM8pX4CzEMu0L55TCECqCn8wjHqwA44EE+NZ
+ubfAjGQgmL1xVEvBSvtuFZgpzvuGbF+HAspBqc9ZmaRFofKkeWG333/fvtK7GpgV5vaFdsULZwN
cd4swSfCG6RwiunOuoCcxF5zCNmhZPFX4xPxkYhaSc4bV8BERVTQ0ZXT1VGVSCZv4whbqYg5T3gQ
/5uvH7JNus6ieIG3yM2YzD+e9yrbDX8h/UsY83Gvp9kbZ9EqOICTsJPjti5NBSFggb/RY0J8ks07
2fYNGVF/vbwNytqRRRyq0HsfOaexfV4T9Vs+bp/jLyC9a+aDis6qnDwYJUkP5prsnaDm4lvOlJws
EWbfSG3IlRM00/HtOmtKSAm2u9l113DG7JH7FIyL3GFDf+2g336MTSTnEARFlE4WzqlWE74jDcmJ
YS6nUl6aoXW9NaP2xYmEbQvV6r+cOqltE2gaVdL9zpJ84C1hfHfVeB1FFIajfSXBYlxtJI8Z338k
Wx6QwGZIXz0s8m4tlH9zPfDxxlPIG2cEIU9cmaQAlre7n2O11dB2ISwZUbWvidZgTsVawzKqbYl+
nBuh1TQaoQlUkkRuYGfYVgcKgcy2+QvuwXxFvPYqNaBdwGfYswhPmGhlRzApZMyBQxf4KQmlQBLz
6RKhN3J2MWCWYtCD/Ff2KYQgx1T8T/kOY/2g3fhOtK6feWsNbxB+oq24AYgoRlL1hmRCSyiqysQv
AN5KvAHXkjePi+R1z5t62GFR1nyLkXl2XLB9dDA6KazvSWaXv4rMKDz+POEyphpHhKEZPzBYfnDs
cXPhw5+3+Ygna+Yj1Xg7vE2nn8/gHd5ZHO+yQmQiknzgfW13qk2i9ljQ4/qqKtSbAtaF+K8A8CL6
PBe0/Yg99E77fe4/6SiCTL6qE2PuGJzF1C+3tXI4W4vhoxFf7I664p1J4BMjvXmSrxIJwzgeWcPg
8rKrbe3pEejqYABZk08J61MEQUYKt1OHS/yfrXKM562+/MwEIdOFnhHLUEps2qQbd5OTLDnPl5Dn
KfJ4PFBIkLwVEX1RP76inKAc5omk43bQfAJJw8wW5h9ExbzTfphWvSTbXcNio8DQqy/XrT+F/ppE
OFh11F9nrnAwWbw26GRk7DrA1QmwUsTfTdHobWNz9xVmOXyGsk/SXFv34+OpXoziR6C878PmOp3H
dOlMXl9j1Yj1BJ35Z6/cg+SC4gxpbZobplOkvjGh4AY9JiUElAVMnh4ib7JcTVRM/d11OCqpv0hz
YyCc6cgVSusDQufJf56p0xXySXQ/FJ6fEU9KQlHBIAlCaa17PUupizEbD/Xa/bp08Ld/qSBhPV2E
HrJndQsT379nTclZ7PUUu5yyJA2YxXqYHMH9cXWOiZzQ39EQ9MKZPezoy87qX6YpTqCxdzFCbdjU
WdwojCGw6bPIrnfpe6ftf8+gjlKfwQz8bSbvArhDwz4vIJhzGJ0d3AYiWsAS24oO0Qxs9dg9OHfr
XH4iQICfuofkX3WYS9t/0lBmwHkTc3xsaOAdoJRLK8rC8RB1YRn+ZqOflqvy4iQf3ehGnMAdGSwB
U2ulLJErobepJHrvMAHa2sl//G0Y2MMihDx0MBG+lYFtIy1prMMoffxmukAcWpb7qRD3A6REyEmn
0JoPNjrRFkK6B5x7pQEgGvUQYXf+c6rA0lHr2JD4WSfhIvWaYIS0Na79Oo1lDKynx24FVDAWx4XG
3L7KO/YxTCjxU7eBCwedER1J+ytRQ9O+r1Oj3AF23yCtw6/p3l98vakuD8SCT1PC3N85dqZQhfQb
cxWPmm4JMHyqR5m+nnA+NfaUgdaFtH9h5akXqDOJQcYGHhRbyiKRNFHI9qq0ZCdx0gOGhorxUl9F
eUKiu3kPWw5G5OifWqAeph7oFJs5T4VnQigAm35MFEqu19oeXOYzGdrjsxlQtEwtwyHBPYpDEsQB
M0DH4qo5h9qLyP2+8eWJogtkYfbHfsNCDu99/EvCEpzs10qq4TOH3OiXREAGg3PuxOlJVUKxe5Bi
a/i3k5bCHzMYsTVxPsN+KtJYGenN1vTEH1nrXf9eWT4AEqRb6pHX+Z+9D0dZVO+BB24QWnbdNIP4
KQY2MNhHJ7f10me1964EVCHl+XB1r5/CD/jZ3cDcTMXXuRbCE97FOlJguhLxcyklapV/LujEqOn5
yWdsYFOf1Prvx2+JtT1GFlpXepHife11WBGH++3NUiRnUNanMMHM5nD5VzpBDE/L+7AQkXjbL+FY
sqFKeFJbOOfUclRax3TqnM92txAuoP3LgnXf7ChdnKWSGxtTfnqHKHrQF5mcrSCO5N29pZYwknvc
dUCmC4NKHwRzi0NKFg2yajNs1INSBmqCkVon8+wQs6j71RQY7PPX1sebwUuLQoaVIfQr9zJK5sy+
4c6UQNDOjcz3hylI1iKf46+z3cRIdlTYLLnah1E36DdPi5XtjgVaf2EwOnyYVSVYz9T3YmZFzHz4
PllWNKbhda8+U16ch0V6sGPr7vmj4pJS05DFjafRFn+KC7d+m1hFL6xCLz5hXGQHCxdOfPUFbPBR
va8tSKozkZPoQ21wG3xh53IYPxDJDnjdfS9eZCZewnlS2lAD+UMpy3sg2FM4FWkQ5z0a9Aj9ERhs
9zbeyD++lE7xWH9r6lhZEIzxqhKHh9ecqvz2RMOlMMEXzxM223kN9Lw5t8o6/DaCYVZqSXE06+Iy
+uYvkfityqiWjxyNCyyqXuApgXlndBAdmwCtePgV4aS8LjAz87CXUpuCFSuhs4Vwx1tYuIzLn0kd
5ZnAL4jWsl993qZJrG1bKtVHQgQZwMOuCfpOd6cjyUXphQADkmhBwOQX5vZh2bCQ//B2ORBF19VB
wwLgKih7Ma36qrd4oZ/LhFbQRZND+mOkDGG0VE+GaSsXUIcYCeIA2po9A7LXsYip8d2A7TOMASUB
s4y0DDE7VL5qeY1ZYI51l7V47VMcjj8qj6S4Xja2bWwpABDbEMPYKl/nnUSp7NNvJGqmQFQJTGUc
hKeSdEUG9PP5gdH6uJs6XmUUemrDUGtCIEagwcYz8CvKDrC3hp+uwNFhE635el8aJKZ3DVJmpZkr
pM8wMgKSwWJ6o15Y03xODW2A+UY5wcOEP5eZ/4WBOhjDjwzgdH7Pu1vGiGKsniOtl/iLxddaGM6O
RA225I5FcgA24tDffU+eFqSawVxNbWwtCvZU6xCC0rYvYyAClwdVcIPuWNoYFPQMDoxTX7Jwz0QG
RjQwh52U0c5i71WBgjdLmDNDL0BLjw3pLrok+5K0YOjgPdYjbSX46LC1cUTIHJJ/m0OOwT4C0XUt
B86yf4Vxx93bZXeAGJzsvAXSc9cWLHOnoAZ5s+p0WaDl1/ReNj6sQldPQqt2D0PZYh28aFYEyuzp
KjpJetlruiNM7CrnRE8OGpvGVy+CF2BZGeLrT6LuDvYJqUaUOiPdLurCKTCFwz/TlTEYnl4ar9Lr
jWU9kdRuyi8BaKRAd3Uvo7/HJJxDHYYMwCn68cbqeu12dpxK+sPwrUI4PqpExyL0+aPCmeZS7dd5
uzC+wDwUQW1PSKlz4doQciO7QA0arLEqgFmONLPKX/9PEMsZk6pmdwzEdqf6fhLUvanoCYn4TOH7
rEQXLyNOkMmgu20iU3+Yk7An89rkv409P4er48WsKAqFe0w5HmGZW7uzE/GJI6ukfDsht8kYFjuA
inajTf5V0eIXkEvurp5rEqSimPbP9hOlz0Dnwoz+CDF1ZTgBIe3QQ5ktf9Gnrzj+KclAX2VrRdGw
VKnUQjPnOXJcaELRtdyALnNYsiqZOmsDVI5RKm5U170kQQp+gQs5OylknYCmu0UteXNeaHrQuzjs
LlvHub84qO44pUUjvM1CdihwhSktWa9rqS0CbIiaHfObkDxxLaA3713WvugdCMYr2eJastkzP2ak
OtyUpwXs1h1M1uaVi/wfRLVVSQ9xsjTmniaMQA1mtoiHjBb5gpnR89bnQ056fcPZEqVBfK1pLr3l
UR0EPEuYI7AHo5xQ0IPBY3o+VyF2T0C0Hgcmoo1kwiUD8zTclym00FfDs7BwfGvElmYzVGwgF0jq
QSjqHacSu8DyA46bp1y9sObj9nXCjKNs0JkzcPMubXDxEpH+5k9dZzTd2Fv9Mrjz6DM0I3SVg0kX
RSromR6CaqgwI7E5FT16SbnoAA4HTraSrXPZLtmBgJN6PS514N8bMycV635BEIlwZaoDOxlOxzi8
2N/s9grXpOaz4OXxUG7vYKiPhgdD73JtHpy1ss3Nc9l//GwfvrsxAEJEzMZwfAUZMojPJ1/gvJyh
PVdNMvCAUQXR3jV1wQwyKn1B577/5iktMaNG2rUrv/wKF5aJU+tyfQK6ilCy4xknw64YW1sgJK57
nDuU8h5oJmsEMn7XLKF5QBMaalk1wiR+4HSYMWU2mcuEqRwF71KXuzHRu0XrUQvTIYgSZ2maXBwt
KNDGxDhGzhLZorPSJgR6FDsP65CvTIj7YevXEUTiPZRaKJJb3+TmeiRNenh7eaxUxxUrj7okEhbV
JyT4/kN9oJaWl18LWZhY81SArVGUKP5Eo/k7TtcS+p4RiJGzCrOAZFv6Ya00LVsWF9V1r/IPTC51
t77/EVfS9gpr1cJqJvQ1PHTUvsUAYF6G6z9GH6Pfca+9P4CZ1VGrpcUXhjxYv2ik/sSWSoF+45Rd
sZnV4fYr6nyDv/WyqKNBeNbeZn1fqx4XThdG/b0aYB0JTSEMf02/NTJXtg3EQHJjwCf5BuvFha3v
7SVh+LYr2gaowBM1AnR0+2KrqYiMLoqI1rCzpeQeCyvOF8JcDKamWyvGKwctmBUGwZ/ehwDvL58O
MEIDuVYAP/N7lt3AUwgSxO8gvV3xyyUusR1aEKBhu2bVcoG4jzGT9C815CUGFDsiVDYcDCF8+9Ht
/mglrOJjnEJV5ZnYcljDOwbyzpdiE2f56NwThHp/oAhQY/TtHMrv67lSWIAdiNF2LoGpH1l1MRsk
TNNvI9tsfoqEla3UQXJsyqhQLDldHKZZsW/p+R83JY1Jb95j36/fg5LVTDYSmkLUAc8CQ2RypavN
Efl+IjCNlWCW71NenyGt98Uj448aUa5JchAy8x7kq5vVLY78tcXlROW7EXfCl5FIwNdE7rGwESaX
t6rhN2+1a+5n38W8fr6SRYtkkiiaxNr6y2Du+6mGOtsrsV/+p2c6unN+zUYrgphOEVeV1/zEAbA/
o0dn3gklA6wpY1kUiSwFTWPdjwISTQ6R1K2Vycvvjxji0pgMNPV8YVWOV7nh057WYOvOCyJhpvxs
BaqzGu7iok8W6XrFJsyfc37icSS1n+ibNVjpcYgv5tt2JLfkE4BQO9tu2JvJf8oMmxonmkNoF1n7
hL46dJWl5Bbm+P6BoxyQBjzA47q8ApGOVAt1qiqdjDHN8M/+jCSFr3vOcm4KFZRuYBveo2b3FXNw
yKMkZ8RQ9zhEzdORM8r3YgwsyoC5rfuGJJzAkCztqiEffbIijwWU7n1D+Of8BqUlhoQ9rHv5QNQ8
JdAU9PVqo+gWYqG95exHUOfNWNo6zKnkQNwfZTKofuPPcWKoJCYyImtaEhq2GDwf+2M746TpG+f0
4pX7wJaZaet6vdFXCQ2VM0eQWMJn/ldsZmSRP68Yd5zKdqXUp/floFfJKVHhiOc/YTvzkpisv8dl
hC+7OD8V3W83gGSEpq20FqR3JUnl7zWpKcD7Qsq1mrk4GrmvlDZh32NJ7OJeUG9jZx7lHTKaSx9K
dnrVv8FCkoTwVNm7wr6LJEj8COlg9dH18vLR9osyBig7DHh8vJcOHTuX1wgZAXvmJuf/F6dKnCkw
aJn48d1QmAxyH+5hQMdfH+W9wrc1kuG7c252iWvdSigcNXu67zA/2yaiU0l1rxynPxu8wI31mQBd
M0fOXCmlZUAMJWwUdNhU1Uz/IQsYxW2XJku6ksG3hc0iU5tNxOUo1vfZ9SRhWWMviU2HrlOhGl7T
3gwylazzSVB5+olh3R4TJRqAAptG/SqtjRPMqko09MksgsNECjJqNsKOq83ScIHI/GDaauFEiSDV
s1NlmCI+LoLkAjqX1lN23a8cx+Q6qZE4+bsCc9wKgVNHLHP9fsuEsykq6Q5mFxCHhd+YJHJSJHOG
PT1ec4PZKmLaXwYudlOliCs4xmRbHs8MOdYrytpzu5ZV6X9Tu+Hk5nG63Iu/4lDsGu+DZA2nXcZe
tu6VKvjX200FRABt4LkTH5ewV8qk4t3TcDSojq2RbfALuUjIqDB1rb8bGGyWcmfsYCTehxp/8NGp
Zpxrf7i8tERcJynzMEGj7gNVTGsBex9aiU9AsN/VRu7vJCNahtyRrkLpyuA458kFb/5CROirkaEM
srIXWOuYzQ+Oody3Wk54s2weRBN07NSuAM1zhwEGTqBH3sxgxN+YQfLGohBnHrSzql5Pa2gYTj9m
I6n/gzuhpymO0GgvJz1bE539OlWy/hm665QWX6U/51BC99vWzMcR8g9m0AsaaXMRGC5hX2tzg5XU
bbgae0SyP1H7Ygx9z9uQWOlIIvUyZRyx9cFxWug2UYH5DZ6FID6HQMRudo35UptFJYr7bSUDF3YK
J1Y+9pNYHCmaSXXXz742fGlkOkXog9W/sh3WH7exOS6pkr2KrMIeRcnTto6+MwVqa+Ptnfdr6uTW
WxVDVpob5KkFqu5l984ICZyevbssvQl4Ymn5t7S/UQO/BamRJfQGeqXHQAzcBHJLMIZmjbKc9sK1
DnK1lTuhYqgiNBYIakDCZEOGyjwzfG6aOEKSa5ykbubRYxp5sBTjNlk6ccdLA/Xn+nH5wldyI7A2
HxgFXVKMIgylkHTqs85FslD0TimBhNbwWtqsBCjui4E+Vp7C+4eSLruDBgcqPCsx5Q4jF7XJG0k8
P5w0NrKLGZosAhqu7r2bT/F9105183NFs7EqKROD+6tMrzZLh2F1fI8Pmja8I77jEPslbWdFZjIH
k37nDmCqwSUXEQoHhKdzEhAPc1kEwnjf/kVbt/0cniTUsKaSHOYjKtIAm9GFMiBZbwkNq6m7pMAa
tmFXkBRxBQhIzWAhDSTry1QuADn1O9TI8rcmIL2uUpXhd//QIjST0/puv/BTe6qe9rXhBqMxOeB8
qyuoxdJ49srSghKVWrSjFpriQvV7xSeJXQVhuRYFzk71FW2C//e8aV2jZY0DK4n+Eb5hoRLbNzGB
mbhZkbCqB1ZxkF5ndNyCavowsC/CUpqQAFti9O1DmMCKaK0dJEpB+z8FghgcGAFpvuUMI8hL0Lvj
qdP6rYDh/j/LD1yEsQOZo3JK1m1LY7SUK1Ku3sbQBaN83mS1Q2h08fQwNko2PFdavLg5Xy/AyQBd
WvAtQsPWYZdWFEVT2YO52oNzSTmIsgQBQSLu9cM/uz4yWKgCnzgD+rRtd+Om+oAoK0Cyw86Dz+gd
/vOA2tLL+X/Arc4Bo7FZF5DPEmPWFuQZuG/tdlhAQIqpi4nZ6qrFUSdonBDaOLgUpIeZtlZ8tFxA
h7pLV9wgbOicl1ijsMrudLMsmwNzDFhoCbKwzHVSnVo7HUnBsYd5SykvUlWRj18C5EBIMFBkCEBi
vdKaY6mylC0ZIUD7k/8mUhCDBrD7KMgKx5qXZxw9evyNgL54g4DQsQeX+uV7OmWrOmhsaLGFYTTK
6tVNtNmtOI+XNeNbbwMZbLSbbfk993Fe3rQdJU+Y73K3qXtpFGcwx+TKb1vX88N3WJ33v+iwn8DI
vfP6ENQPGICeDkpljlEUzgCb2C+w1LgoDTeBpldl8a9chzC4ygDY/sVXpJWvFgVcueQV0nlf7cM1
SmLVcMkloOhwKJp7IS51iagN1yqu9j1lqlgxByJM8FSjnbNAteyjsjhDNWq1d8MHiix4PKIvdMhm
hNhRLbSLSY7208hyfIQQMeFj0DhHZdchp/NgQD9655kUaI5x7wAMgJO83BR3lWhwMdPfPjgP0kkq
Wa3Ko1xyhGMnuXLlN9vZXfTQ+7ZsJmNBqLrxyl0WVW8NWlCNXlNmudyegqUcD6z3BCK2qCpApC8s
Dk10LyV8JcWK6pZ9wRHizW+ANHYQuv9BAxXEUPNN1qO8WzNXjYAPCN+0jE5zScfk5cIOm13+uTkl
dRPaCW+v+nI/s2XL1i0SYeYwXWoXBcEj1W0o2N/LY+Wi8z0H1MT0NqC9IZiE9RqvxNk4eH/s5vck
yKLQPx/tWPNkbvc3hextVwyOsOMRNEIOVe8MWehM+YA7t1BQQrGQ0jdEvkiRf2MUG+xeZTi9Bxtk
DCDHkO1GPIZZUUkHScd9SFpbOs5Wu69v3Ld4QoGS2iOPXshr7Y8kvl0VKaUmTZCYD6gXwbx1tQXX
Hfu6C2UYAcPmSFmCuwx4nlFNUp1GhKhn8RJKZfmXJMpUztm2zLLXm56pMbi1QSlcjE8qkcXseivv
UMTG3NuhRWSxdFqL3dNP8mgIH4RxnxC54XhsJ3OEBeVZWNcQVtgTCvEx26C3056FbNueCNrUKEOu
S9nq7RLGzFMzMkQyZqwmSqU/j2ux7FnzR2NW9Xuz/u0TrxfpSCDVeyH0mq8hlFGRz1fuPfnyfLs2
aF0H/IqwelYx9MfP3JkWuk0L8Ked0pBrL9630AHoXiVaJ71IDDOCw7Hm90oIcR8pRbpNA4RcSlKo
uLzupsBDL7e1kzSZs1BhDoC+UYQ6UxsP8A6esMpH9AUxPxBtHkyokGj6oOw69Hc2dy2n1b4wopcQ
QOzA8GyadXrYXL1/nsAUs2rWB/tQj+U9D4QrjtzwLuZWR+E1wsSR5+zHFq5hX/0fEEMmm97pGl+A
a/KieDrhD64Ss7d5IEJHD7V1Cm7qYjcRYlJxxQL+JbOOg4wze1oFH/aDfYaHEswPsbosLmRiA6eW
2GpuJZdn0ih0v++Nu1WdOHj6DZE2wY3FUrZR3eTMtA8jATCJOFI1QrYyR+H+RnEbYytNuK2GGEIE
wT97FvMCHbhhRz/vrz+8pBdKwOzgiEJgPgZl2ttri91K4i+nGGs9SGgevpoWx4Ylh9avlt8nSKNY
DFA0PGO9Z+qvUuEKTdOCk48uW0D+n8feKD8/GrGAc5pXry/qOONmU6XGTKfj9b8cU71DqMu6jSoU
PUu4fXSmpdDJxc9ZHgl6Z2YSNTQS7w//8pE4hEokuVrEcvqKDmJtM/0fay7tINdveYFK0E3urnKd
y9al9FnjLbZOgMtLwa2vKiNL6O/zPe/TXh9haeXsgEmqFdo50Y2OWwzUcRzyFV+gca4wnJbgAvFS
13gEsPtDnYic42GjsBEkDFfo2cIVyqGmMAUMF9u0pGAa0tMwIh7Q+ykF5c4JlozIqUCTMEEfN46d
RLHNdTXiiI1mO7c8/w92f78wblqC6/fzy+kpn/GxvJf9MqAHUeNk/oihsSLlMfufljPcN954NwKV
c1uz4zklk5UsLRZBouzZE8bk4ZaYn/aKQlpoOsU4vf1JmSji8s+ukpI/IUv6MwtP9eXgcZLksuuk
nAbc7/4hagR5Go7xwcHJvMSMyqlaqgxqNPgcqJG/8wzjrbu/sb6Xg7cAKqBp5CK1DfV1Ph76p64P
AtBt8e/6GCeu88WSjkRHxQhGVDW0TL6vuDnWcA06BDwaryDpO8Xti1L6UCG6hQ8ax+0MgnBXPHY5
302Rhu8SofCF4yzIarjpQ4Jiq4vOwX/Mxj7HqE3zZ/mFT+pouKucYeantUXPwF06KL8c6nc2oXF6
kCOsHyIN6KceRgy4rnoJwW3pQbIjwyBOaUUSaTD0xf7HrY8o1E4iS03+2VfABVD7akzKkUoDjf52
dhCrzza/EVYKDSzWKQX16mnh6YnAp2JblwVT6GxZB/T37Vh5XqRlMz2E+nfinbfLeE42ahzbGlHP
SdnoUcglT922Avje1CbK0roBAZzHOmhSX9QD3u4sC8Nu26tf3bvmWLZVo7erNABzh6GQ4p76BQpd
RjPflXxbowgYy050OnMfgHPzhiyJFgDfxETq9eiJCIvcSvzh6Yaq9yh0Qchmy3/jZwO3KfmDBl48
A4fmKQfc7TChGLQ5wIeFDFYqPHTWKgNte/5/5jqcg57+6K919FZqpY+anL5nb/LgDSE28749Ke+H
qNJaHONgynOLtgyUi/t50c39W6FQ+L2UX9YFn22z/FIVSNnHW2yxiXRBPv9YfVmDsN7cQoFj3Vkg
A6Pyzpq0NJ+d/6gvivDmlY0gLCPC9AELrSE4oTwGmpJLU1SUAqzQJwRdCadXgsPjO6STQNZT5fzJ
KCXrEmKSRdQAU7sn8AaVnRTLSc8VYp2yEArSity+C9ZrmqC/+px+noEs9DkpgMXC7QijWZew9lgY
jwsFAQlZhw8VJVZqNgqV/oIK/gZ/xS4aqq8oy/HcEy1nFNVxsv1R+iUomQIdNxAw31HenfXZ6VXS
swyeY0ksb76InO302GIqfpOLgSwB8EF25THCv/KoBQ9iqKS2s9ostOYp82DEyq3qPzek98mejD4O
M4YFWVsygO06HHKsyDB0vhKpnRCBYx0uKgiYrduMN7KNZWLMLeYtBJeLC3CL7/QvbSDQ6DtGeEbB
t2ztHUq1WDauVV9rZM36VS8ZtYNwLDbeup6JHW8Vnc22xiEH5/MR49TZRKpukZSA7k956leYj/em
TqMzSpJD/FcxbjQzZ0Fm/VbXRjqfYxAoM+W8EgWNF1JQ+hAybanyaBMz4eFVzcWwBbWSPECiFDVg
XWU/37JcYUE4Mo01qww29ARzFo+fNb2fMzQK4WmhZaq1y9CKS6xFnL7thnK7hKEzT30xV6zF/gGQ
IDiVspl+rYFpfcXKr7JviVSRVH0F5ekzOPMVQ/FaeURDbfsM3wScSqd26KORpuYHvcscLQcISaaC
JD1HbQGuKbaIDdNwEtTmsNfwqWOVkf+DFQTaFkRK/DO814feNTYhB/PahXCmVWbSIiDH2ugmGIWz
jVZZQTtwlFFpRXyjI3phy3rzoiyeG/b8DmlZMyOYzimw5xgFirXrfTCtkZLcGo+O6EUZ0Uk8qI8B
f8vohuDazh/BFmmZdtMyekopXSUY4N8qrpW+7lTw3z+Osl6oMSYABG7MM/PAuc1Vnjp7f56YznX8
CdzkX3sJeIeIV7SRzKWtmxjIxvKpHY+zTuyQ22bw/LUiz3gQgL5DBAqNg5JNy6Un9UilveeYl0R8
D/vsxzL4ljJelpRAY/zyl2RX2pZxsqKBZ7f5kq3fABb0WQXBW2Mh07A0WPbS8ATFqXJzbZwzm0da
JrucBC+9G78G+fTKskwTc3RY5VXGsKpLF+Mmgj7Z4D83WtvpCYW9JCdke3vZXdr2C/6FHjOP39fo
KPf8ohiZy7TwX35+vgxX/wyYBYnMo9K8ljlnvDbqSfX2bnvAzPZ5qYF5y23V0tgxX1JjLALCEg7a
KkkW8P1NTIEpwcJ3YcMy/EmZ5nqmGH3DG9AchxW50n/TlY3Mm0RL8t0elk9PpsqqhBuv4GcC9j+z
O21+CETGdVmj8OZEqmAs/MztvF9JrflOjrd6m0+rqHNJz0Uu6FINgytPQ3bdcIOwC+07xRkN8MA4
9l7idhap3RN6euvU4WJ1RDQ650Tur72u6w39nkkY1eD6ozFfdRSxXI2LZ0ITudlvaFzGMvZpSDEP
Ss2QYqfA9kRCJ8IfvMGeb3H5BKFZdg+7VveNPz955s9LJie58D15QjBoAL4wuqSKYOpW7On1M7Bz
5JPfo0g6TVFPmCuRjnYMojQHySk5HHBakQvkmbU7XXkn21fM2sMjnryCoURerFCopH91XciAkZtW
4LEAbkoQom2O4x/3cvuhbMeierFqw5AuoIYY6hMI868XFUHmNbREdd3z8k/7K2duyn6REDrJjvN9
G/ahcxNfIDn4OkwFLE/ZOVe4SiCf8mTry223pHp0Pl68Ri3lndEpmMvuzBVVO0FYbCMSTvx9Q/N8
oVNoLaJ7U4zYNcbkZ4X2FmAEJu9z678FQ72bxLGOW24wcjQ3SW7MDqwNW+rP2yhIBbrlBnI5OHpf
/3Ry9PbiMYMGwOVZWbzi32f2zjuPX4TNLhbFzFCf3y8jzS6mMVgpu6j37RjjV2eb3Nq08y+0XLeU
qU5qaO4CBPc+WnzkOLyyZlaIHfKJ/fjiFiZQ4B+byj6EgWiTJhG4Hpm7a1b8YkKHjKr/6xa56Ukt
U/vKxbDDJoUQO4/Ri/RCBQy1id2jQvhAozKudd769JhtFGjLBJk/gmF3LyqFdse686SkhwQcoS16
F9Ys1OlcOQRwwwXEv0YvKFB3w6jVMmdMkqBNonPWeZsaRmfH4bLMD1gpoZ+BfAsp5ttdKItVDEgj
gEjWsOPxOCi3Ytla70jTodmZXAv3jRHAsRgtuL3MF18Sn20I95i+Fr7pJDeomeE/s22gsVrRHG75
tQeyHA8NyFIsheiY7kfRS+PnIu4gg2mDWvF6sWzT9cKpjvqv68wL2GKFF38UKG+aDegYyN4C8i2p
5h4GoG0WPikJNexxnmb63U3T8MGCV3r+rhF2HozV283E0BkOafwACgr2gUWmXewlbnlm/V+twRmi
R3hFb6/1ytaw8pJK7w79E0p60flIyR/MQ95x4XOtr4lGh6OI9l1JvJHGfYxrZlu9hfvt3NqsLYyL
cWkLIJUt3ooaHSnjVG2lmY3wpQNXUn4nz0elqZVOn8ZVCkZq7IEdqtVhZPG2C6ye3oVEoNUK+9d9
X1tIMKk7JsIXTjv9F0EeXuU3MUkre0xnWwV2ohWmNJIb4h8CCx/kryZhVAOgZteajw6muaWp9Og/
i+ljIYvIPROAoydgRfXQHgBKeHwrqZSI7g/tcNzpN5iDWKM3FoWCU7MtvD6n58hNs0RXT+YOOoFq
KsmtbAoVl6ZzqqrDTw3gF5Av4v19mGr4ruQYNmB0jv1cjFatZyfTEnGZk2417XRix+SaUAFiTZ+T
D7Fzt4OfZ4clBtLapYgjfw9y/W3BXr8hTXCZoe7DG5Db3t9oTjMt/q/isf1kVTp6A8IVABYNo186
ymc2vSbm16arrKA1Fgs3BWKrrKTWwpO5buv8z4SNPM0Yaf7eYtYqRnBpy1gBmsogfcYQe3IWhnlt
RORJA5uVJ7UmwLvNIKCYhbHosHmAp8oKnbGxrpdfEb1GK1IYMmcgdVaw8whO1LdQrFmdx1FZn8kd
TdjiRhy/zSMBmaMZnv8sLUpqHakNCgOBnHVaybUWrJCipRkyXyWX28qpxmjUOqs7txDXlTE/v6hK
I0HAmCjJtedxvyBs3slg/0B1Ti3dnAFa2CU2W+xRwsHXuGm4iQ4NtOJP4w6Cm+9QdxSYP/wYjjB7
DSdnVZWvlGWDqg+PnIzxwhojg8i0fCrhDDgTOCW7sTlnFndnZhPr+r4ozOo4Gx0y8ZadBqszQGUb
2zNdX2sUCkf2yN5B4ybzgeOjkVSaP1zAqOBUZKmyKB3MkKeeRJ6x/QhL9+qEuD1Dpshy916ddb46
CClt+4mYusDt66FPtZm3YaBsfNrypgFJfAU5t9AljgRGEsq4hWr0tXPXh1ImqIgwN3ddQJEPZ5nf
BZjLe4WJAx4AkTrP33rhQTHmq9A5FcryQPVsUgmiNxLuD521ZLgv9Ot+mrdJGMJcdgvMonaBtx0/
khD7iEyfOm1bM2s5Ib0HyxqdKXZ0XivExca4ANN7PnLqdKJAdREchMC0e2g5U8oxBIqkrXGlN2ti
j1XIyN50v5uUampnch724YxhvSS1AYl5M92vve0S4lx9Dn7rH+CTtFs5FR2cT7mXzyOiD7zAUnNn
3u6kzlTId8vwj0ZPidDf2wnXCbysmTZrGeXhFp+VYBzwZdh3Ka1JxkZcyPqldKC5bQPEcgSS9gZj
fYLW4Qp8AuN1ojDDauOejnYxGNI6JGHNmquXHkh5DhFZPHvRykjzPvF9SKLJr2ca652kzIySZ8U4
pkUoWVNS/xBx+ziolWvY1EpuXh/nM6CtxpzOjwZ/7sNGh4uNGDwNhD0wnK58ibulqy+vHai13BLn
oA7LPYhOmSTLSEU2hTaPxAmhAWPJvh7xrg/EmYH0OIMCsi+oOdpUnHf0x+TEb6KnSzWLnpXv1E87
xGL2DIj5RG8pU2nFO9VirlZ3huWkL9Sy56q2+83gIEUn09ufeq9pgpT716Nn2jIlCl8/doEMLJyt
AyjijZELBI6UNZWdsaCoKeQXFqSiq8OsrFSdCijuMnjuq5CT9tUhDZuBppH7g+3nWqc/Yfh5Rw5p
1ZXu8pe9b4poIOhx4hg1g22lnLQ8A+sYOzytQZn0WzcqMgKl1gcFe0wGl9LOWqBtaw9fo+eZYu2F
5EHa0FEa/81dsR+PeQL7NEyj0cI0qH+EUlQAb10M+1qbUksV2ArkoUAlAXTxMglzKySNi8/obYog
cfQGFg6M8Odl5LM8OyT2zkBrIbaLere2xeXAk3oYIlslywv8NvPqRjD7Z4NWetA2A9XT3trOH/o0
nWFqKagskNgvRbuAB2IA/1iZox5xge4ZtaXYLuw7oszquJ7AwRTS3mArSt9R4obx818u3+NW2Fkz
AJvGv2itzshiVRmjwFzQAAhkLVKAd3tRQSXptdoOA1VTb3rkQyiwcB0w4nWDLxVGDK16BeRyP5/E
vnB1Q/2GAoYRQIHKjo7LRpZ5T3rJ7gNRqG1AopP4agjYxHAh9o8080BAc7PAP9R/WucRrtDH5hfp
EyXhzKByyHBBsGSN8AFxjwgKQxhQjDSnx17pyZ51l+Pbxaj1m4W5uzGWmsLt+crl7Ys8qt0CpPrz
BpjL/dhaa6lu9ug+Xz78IEjFFH8EZqAjDcQL9JaniufuJXHKJQP4/7zkxvdABq9RiFZPKL1p6mWu
H7WDf8RbUFRAJbzx4A+Di+LbCXDzFZmAKZFHsPjDZ3D0NBqFi9VKiVXdbus0qwCnrnq3KeLBeyyQ
u8jWbVFzLPfNKQKIEBxvHs0yUHAiU1CWDBwf2Fe6F6UiPSDqIgE/FKaWj6KV5bCxJnqzWmBiIvcK
9sA5rBFpOw3qU30c/6b7e/CjbaUEaVQo1Qm1nhPu7ZXgsthw4vSYpBpXVoQY7SmddPZkpD4D1tDU
f4UKDlg5AztyBUeGJQ5wyCiXzexsO+YR7SvszZgmh0kzSK/kSWFdYNyGkhqmjeRbx0SXaaH7irB/
dA8CM66KDsfuZjrBFJhNLrLo9vteOa2eielXoi5PNxXj5bZgLQNZVU64PFRhencCSjkHFOrqlqw1
bkUxfrtEr3EzPHX0ro2yR9K3IjQPyAaDS4hmc9XEK6Kwmordm7QOhgtSs+Bdh9ZctAZHAeFxEI0f
U4hv/OPZvV/sJ4U6hXtivQ7DF7LH45YYxhpPaI+yCoxRJxK5VFalzmkAc4TV5XKv62qkVoImOS8c
WpEZm7A99Lsybvmy+ADU+wGcJlt0MngR2Ge06uou0eJKbXDQ0Cq6ttlHkJFmu4bGO9utYGC5JBmi
o+oV75kW11a9d0rVXMzXo5SR3vbUqkLZHpfQ1zQ1o+YKgRmmtkSLCptHni09WLBLTVhT3X7Fsygy
MsleDBu5uZPM4FDXSx99oZzLWuvrcJf6pbvAxSK7usNfgLiPk0hlMLTrUHrrtpotuYf8iPczw80i
14B5Vl30c5ktIA26LaBXn/MQfxi5lSz+li30ZobLLzKgFds8kmjF4Yo0/GqNBDZBAX62tGjzeB0p
9p46cPK8QaYfpz0jTnCq3L72RAKqTTZt2hCsOueGbgXejig6W+I1Rs4Y2ED4aXtj73XiHY5emJHz
ZoOXLrEpH2df6GVzMhbVl6BN1q38XkBrg2zRgaT5+IZ/chf21XmSrdA/dvVIA6XUTok7ibMiZtlC
E8UmzYuTbcHIb6McJb9dcKNe8l7v+8VJ1j3sGztKoYUfKYTRKJ6c7zBFvV5xkTxRTTR5F7S5Cjbk
NtMd4AVjSKQMynIsDpuQcVhwrHCOCOLNVxLupotf2RKecb92EaNxwJPZ+9Kr7YFu3Q59IkRm83xS
YkJyF0AlpWp0+VstV8zX22nXWqE1ClbqFPv/o3RfbnZhZOaEDyV3TNNhG5QVN74lWEDnlSfxQZIG
zKueGMvpHPmYSX4wv9Mx1uLTpDCZ7qnYRvy78mETvknDe0Fq/xk66T2AcfoxkUeeCmbpl6BelUh7
eOi7dYtaeJf9V51FOZbgx72F2bUUnpjJJe0MAGEXR5B8ezXiuvJg/x0YQCPNf8ZCX8KQ4Splcndy
iaREXoBIhWfGIHdNtxzzY6wrHj0NfDPK64Ht/G+4RrV06ilyyT1C2ykQlBm6jPZzS2wuQDqv06tH
pqyexAZJb41Lk2I+jTPQeZ45GvA1SjHF2KUjCSoTg0cp71vFlLWtJFkFjFznN+ionhzgMsY9EP5b
vSUP8DHA+MTQ+kxlVAHYmnJO0WBLk2bnzUiq/hOXXrPVsXPUhQ9v8kxIZm+tgRQZBVBIANEqO9dl
XiigS2jCmi1QOeKiyOnHef3vhaTSxnVxcgnRLJz+pWu8N5itayC1Jr3Q6MJLwIaJ7zI4Gk6yzpA3
12LQUze+txDEKq7J3cQwAx8eHySkr6JH8btD8zP8HEOTgD8j29+chBaDTKq1VikVDRe2DkfCEA3N
aBXb81mA/C4dmIoJp5jPg7GD+JQpWse0sPxUE8RhRiq026kn4koVbpQ3v7TYW80klSIdqW85yIFH
ZbnBeTviDevYFV3nUdPebs4n/encrg00vkeG85OqbZrj8iCE/EfP6mydbQ/t50NoOoqxUqwz0aza
tz940pUoeySuLPWcmyVbDbycnOrfeSarpUksi5RcV/WleLHAa0R68GMulWAUDc54tDO4xssY58G4
77B3yLS3LMg0gJJTKzqIGtq7MGWvV+NTKQcOAhmbcolIKhvGON4tjIGnuhmVB1xCQc95BUQWTbmi
H3NjWfvkDbRhlL7Z/hXnSa2eZxRhyu31UTkjEWXs8iYDliP0j6ZnnstEtKQQE2Y/NGkzDU8LC5oe
keJXvhva5R8+jnfxgOisQ6VbWnQnjVIHjJ++Cm4IUOqcc3p58KR87b7PaBcf/rrX8O7rG22SXYPG
1jscC6zorXt5RfcBuZ7vIJUrBthSF2xx8/zBcWNcmKQV1TqANmYt+jkr5hAlgk1tM3MvLIXQCK59
ojZtquQJRi2lbJdaLpF6hDE5ekVBRZo4l5zkw+D0FRZzniHUZkKOzl0wOkeSkTXGOIi4jPohrIcy
QMgM83WJrdaB0krFt/OYtCxmcWgs9wsXlc7fLDojlKr7dIiP59RnTh/7gdil4Uu4b+l7t3DLoOYa
PlUqBQaomzr0LNwDHzvFiUNm0Wi3wXVIDV4ihJjUk02b9MlSW+OAVVvlqkSW2VMUcNLDcNbliD1e
qbXWsHAG1vkLrq7ATVExHhh09cfgzMkIQapew/mBhrjhIVn2kIXQH6YWiIg0JKa4IskVzeNcTai9
1gc3O6CP7jOSo4MznB9MHyOxU48aqjNCv+VjH6ugqZVxLwug6B5/Po8/rhRcW+DsNTJ4PppaIRoO
P/x7Gzx1W8KJYsgPTpsMICpA0GTp+NlYWNok5iXrV1eyaKfaQ6S43+2KJxdCYmmCp679g38QMF5N
srvA6bafz97IOVvWj73xoEDEX+XdgjbcJ+juSQ0WVjouL4TcWmL8h7JnKdmczg9SX1hn92p+8J+1
uMxqjQWNtL+c47wePMKGpM5+Ks+FODh3nrdl0Dbbjg7gMQuqwlgvBU06r/c0BRziZ+yBJSjdOVk5
jCIGZ6H2kvxc54TY4e1tAKj9Yx7yDGqkI7R1q/3ghHdr7c75P6E0DbqfAWIzOPg2sSLM5pGinUaB
wZrmncnWkRoRJqZIh93v7Hso6oCxlbTo4Zni3GsDL8XvOLB94A1DtTxNU0mQRnc5p5rF2oVZCsW8
E0yc5Zp5meWSalQZOUnVXR41PzZX2GJ5UuczUvGHNk2R4cAmYLqwIimeUPnM40TiVNqy3Df6qyyx
4KwMdbmS/fyAcaiGTuN5e+nfKCl+P4Lf96i1zRq4Ol+q3PWxdsijahfueExVEliOMUcFga+GjVgu
SZuzskHPNEiCI/6fLZuvkrOFAGDlJvETeauMbselmHLLQWu/pP6SqLRpOMpxdNDWBvV8zNoor4M2
Ffdan0h5e5rMplZyLr4PawYml0NEPAwuUIXMf0jrvVuW0VAMWN5szZwrNd73ZzreRS28g29DLRXo
GOBQm+B1SroRIzDxunHKEimWHf9gpI1G1cpxuyFG8tELbWB3XfTl6QQhnJbCzMQ+7SSYAiLboy46
VSt8uAbeoF1Ca/GGxUtwpbIjFP5xE8s4zcSmBGLU/rC9nAbmtsnLGMtJwDhLjw1zKU4fK7FRt33A
07RZigu1825W0QpRsTcWY/uts3PO2ZPkb8AyM54d5Qu+MC4YdEPzwcLJe2nnFFY/ykc0CEOnJXTf
kh1jdtDdmN3lwYfZRucx+BYhikAejm05Na6cy55i2HPz9uwWGNPbGp2RS9onCz7ffDycESmo/pnv
ioZPysugDXyqPe7gi/dXQHAqRlwPifRrbtd/1ECbClM7fGyWa/6mgQEhNqfzUzn7hZ60M9hkmws3
82w9uTmslQHJFWXm/VYcEF0sOY8zXS61/Ybtdl0UieuSD0mtv8WohBHGmRj066hGPdq9sWX6eSeH
7IlZecWuxJEXv7KhE76vsXygym3Boea3EYin8HMQwMUmawWuqOQDxFsIQEmyG8+cNKuSmxvwwwkl
23yeOMsHaA/IYbYZ1kde7IYCijZcsTsf4BZoHB6/mr4gUmmHVGsAjdc69dJaQmFFBdqZR73Lv1Di
5FxKZrld9omZIuT4xrU0FK/uptl1Fsy59S3rnWUlyvzhV97XFQWW8hlCKWvmQ+KL6BOI9zYzE2Ix
E7wVMq/CrEL8c+PCnjDvBiUtWuff4AlJMAhw+PfPRPiE0UGyVZclde4BeKwC1wa5fgYsOdSGAe93
qiPmRs3LtCEW7ierztYAAjUralqQAgDvzDS7iHUElPP9+77Yh/fSXNhhHfpqp3zZn58lojb9A1Eb
Rd8ZqvR6/tl5LUAvBllgizQtswc2tPeW1xsSxCq6t1H7GuS8caj5y3OnbpmOng/D8MdSr+azsT9k
Qi1kA7ZL9BBMVoFk5IAQ4AJXY0fu3E150Bld4fVF6PoyXN3dkrmr+uk38NaW+4BAAzSdY24x0Y5j
FrezdvZWX2xY/lw2di0ffdOSQCQPyhwfwukXDygNhHCqqULhdfbMKN820/2GBmonOpjDxcBPq+5x
ANgqIc47ufOBkomwovj2w1oq+VFeGX8Ul3gLvLcgHrfuv+tx9Bem/bCr6FLhVZNslwEybd671TWU
clu3mddi6nKK1YyczGvUJNieAbROsUC89v5KEKSU3GilJ88UB5q93xEzLKtsMZNFKd5bibhz7kWw
EFAOR2N3/wLEoCNwvNvzTq8ObJhZfwfwV/yuFemETIeANhB2iow4plH9iVF5s727dmxNTfwq0xjB
JpwUaog9F3P3wHb/4L1aAOH1AehYxzVosm8NUDo6xvGm+qeqq5THhEwhI37r6+/9CVeMzzCFXLN9
c1iiPr4OP0d/DSz9UdxjXc6gvQMp33lwxD5t/VM28Rt4RRQCfFIRwfk6AmlaYVHt0H/5rKHODczm
Pq5b+1vdkPsCA83WTgRx8clS2oBHxkbG5N5XYZ1koERuPGBBjP4jWy8/qrr/5FM3YfensGhv0JGY
sfoMrjdMFrnIDritUnGMmVnzz3r+G9uKxuYDGLYp6wtS8Gn7BPtxcVrMqYkujmf1rlYCwi3MF214
gUFAtSamsap3TWVzYDsqoB81ofbkPaUKg4oDQh+y4g67okIHQgm1jM1F/jLgeD9tM+PSpG38d6Od
hLNv7PsFWAciPaIGRvb4uJdAUerCiBbw87fYYnSxLwjTrlRLkz5of84E/Jfer8uQoEdMMWNxpvwE
NYKH38Yqfyca80m2/JxCdJQ3gfVci9EoXXP7/V1mJ/P5xmzq610wWsHZk/1Gr681Rm5S8rX/x++T
Xt4dNjjNLnfOVjIFlgt6asx04zjJCImRnLgBUuiuRkcXMCAYP7YeK9aY3/6+zvSNbfiwynwxHnvN
tLybsX2WaXxCrQe1ZfU7TsvwMKhLX8p8Jo8yGUrjBxCDCoNIHV0PZ05ij0s671GBwEGoT4tdxXjG
GzyfVWKzNFHKrMVd6ZEqbNaSzZ37OF9FfjervSVd1Un988KJplyBGYkJBoeGHqQWXD3vNBC9/dPL
qynyEf8m0BpygU4p0VPFoiNZ9f7US2XmQa32E5mEZauGIf7rZE0h9T4VhDY0yhTvD3VVoMjxQDXJ
7WJE0ekakUsa2b1+XnLEAOoL0PvLbnJKTA8VQFSoZXvIk5ADyRYV5MEm/Sy4QP3NgVwYEaai5eXJ
28SNjcwxgOd+v/lsLKqgur28lP1uctKhPF+WWxq4q0UOMktiiiJcUVtPhKqym/WBKX5WOKDfANxU
p0MrqO0CEUunL2AgDCae4r5OVJn3SSwf6rRfXJHFDM8mbvJMQsc03rV1+aOpzw9Ok9ZdHz8Bvdn8
zE8J7dMgxvPMDuwO9ClvJ/2H47ELaEBablqv570sQu+96XcjKLo9ZTG8C5T6SZFOo2UT1LM1qR/Z
bsr6qwuDjAFlYOWfxjzthZbv3rxEiUXjCsk9UBO68lTGvvDpmfsQndN699n5MFRJs/rziR+TAQdN
seLwDRBl5L1zqOFC0i2E/sYaJ7NQeZHmZEsL9pqpfcwvFgAlZXmjeoWfKVsGhPTprkKnQ/Jk60ft
xEV0EFFKa97RsfDC9/4yIj3026pV2jC82rgPg9yroKyBv51zQwrQRcNYn8qVFLvV3j6X4Vq3wUBH
OzwtgHchRZwzA4uX0NlDYxUQAF8d8kl8n984iZTNfTuDR15MqHkzbHjAN/MnJe3J87KSPNrbbyhU
BlKGCKxtTngONxdSahp9OR+0RtjIns5ek047pxolyrE6uMtE00R7A35208gpT4zjSRmNDC0NYnlY
0Ka2wMwTLtPFljdOADZoMhCDDUYXzvHIbiZJ5FL2Du62vG2oUn19fKINX5aQBgfMtyBTX7PeFmo5
Quy2S0qo0/pWxc+YeXmXBA4Yj5ZZvq6tVK37SOW69L1TNv83fsBDFjx3G7Ir/tWGJsyfuxudK8m5
3wCza7wRPHI/AGGwZAY7ajskqMlZXaU6xT3yttmmdmFY2Z+Jxx01hI1H8HoV9I1A3k3vYuNH5eu7
SHs6vSzLXNgHbi1MkNOihWk7cwJUpGH+k7BZccM7LSXrKOMbG3d+TPOIuW7lb2vXC1rTDVm2tM6b
0WiItawDRNMt33oW62PJTd3U1Qo11H6kXjx7QuKQAjSryYNVj6SR4S98GSn1ZzzP5V/+7pBAMlIq
qA7OZBs/HWb7fSf/xTFeUwSwLneUaLWD+/QEdlBwShTLevCM6pn5R8YIi1XiUc6G5GhkmyrGPRas
ZPGTGDqsC+X9ZpWHJCER8H8tKUZF6AP1qHhNTHUaw/yqmIFiAEPWWXk5dX4gllalE0cMviIAuuS6
H3/tez3dIBZoElEJlKPVTlYNOmOkKBugyYZWgl95byLeWJOGSfWPI/6563/nGyma+ipo2SY1mIGu
qOuDie3JvnAguN+vrdAyXx/ihRj6MVFpVSDd0ZDTtfaYj3lWBwYQyJnrJRalXm/uFHyVyK4FEtnf
2mWLgW9MoPefiQdmsaRuJP1cE8GnPwVJ1VDC/4H9rmETV/essJvtjYx7q6OynID+7XS6qXIb2ClD
P9150EpchjRGQLNbDAejPW6BQJKyGeysMj6QgyiSvkXa3iN0FR0Z/zsn7tbxTWVrZVicFZKQD2ho
BNGqUvw6bQ5QEBGSsiwTwOwJssChj9SP2p2PPOX7cgDfKlODwYxM6bu3AytlU99qBqn/ZubPO/zq
ci24m7D9L0vkLK9z756JbVYVrtDWbz4XKRtYpJbz9iKkFKZvVeoNgy+XwkEQCr6TEbdtPqj05KIO
OjerMIK9s9SwGAYxK2AQTpVQvO+e13xVPldIA+ayo1KSZUDk30ukTLktonYnBjqJ+KFaMnZOgHdJ
LGB/bGu3ufPjnUO2cH9am3eqLDbBw86GCFOn6bBBZwCvKhgDn7++jOcuEowgS0S/oifO/S784Ayb
obFNC6jZLsKzySbpvYYpE3mFjeY/F82bVwzWjh1fKOdjCGtfr11ciQfb2lWejwi0Tm9k2C4pCeGb
XP+/35v0MzkecNwg+W6ul9uvX4EMnQTE9wV2fDEyouEFIkq0OqhZxJ3aaVqChsIYR+IT2pvdT9Qb
49S+b/F5IVY867rcWDvGSjrU4RiMfeo08AxA5kthRgZeDuA8vNIGetMhAeB76VmxYHmsRCcde/3+
Cu8gIMw2piEr6n7ZQjqusWzvfJCWIo7qFGjHFy7pDRGzwhncY/MyFoEMXKDWb07ObzU32nrNbRAz
9PvCQugRgVo6uXB+HmAEvUv9sbw0cVfD98rUA+3NyPBea0RDKTF4UDpvLj2SweBtN5BjGjdeGXZy
riYyBnmNHpkthbAJYC7neqIThqV1ug40JrRD9Od04BXLlpqjBHxE2576KKwL+4HFcvVzZmrzCww5
DbSu1wgmVEW8+cH4zzua5IpTOucorLgPKlhLLgvYDljeRPFFq40U3Xtny7EM53eczKS8eWIDraIK
Wn21n4/V2prg1mxzeYhhUZXtb2hnrO6dmiAh7PoXFxNYonFW3gB0aFnMbMD2SeGuwf0zbf7A6e4h
8KnfErLcBhYlICPdB8/moOFPEyCIWLHjvbn5OhEqfDcHaad6dK9yAnhH6bzytU9w5LPdUX2ArC6O
sh6qhqaTj5rPf8G2f7EBILw1u61P0R+tj9DKD5SWnhM4kSMBBw8T5J7of5OkkJp7IQXRoyK2aZRI
dKbju9/fLruux5cCajSZVDXGy8q/CPauRYppt53832yfUFg2AEWqdugs9EE9Ksz+4pZDXQCYPgCY
XoPVS+b9obwx1iKqe3n13R7yS5Sl9Nsg1IERvB5u3O9i7G2zfSGIBxVsWojyjz5DmtOQUC9wcSJe
rPmPeDkVr+krLI7MhWXHpql9W1Eq46aEp8Q7TcFx3kxs/QxYmK56wI1nmQ/TigWwlVpvW8bvrrPp
02ldHNxmOOY+igf1N8kf7SsaZzRwMCW4EcSqsECSgZgZZSIVUPuB5bBQ0goFa8jxkwUsa785/Me/
Mb6zz97yjjjNQGJTPLYdtDPDdzIA9rGDIVCo+OiSgc1h8rrBAtNMtRnV9Jf83xjrjLG+YK5lwvpS
POtk/e+hcSGqAt83zVOynC+Qvm+emPRs9pb+BTUo5Lj1p1hPb4ILkdtCr3fGYJOuKb17RQh/sN4p
3dLsaG7hh1OOXdeqtwHfhyRQklPFu1NdYPJa4c/Z5RAUDNMpAumciKp+vdZg7syq1LgzmD5CLMvI
mdFa6mjqERpTjEKwyAp2jP/JVIG+SDuDWf+YK9hrXaVeLYHWk480PLMLspNprl2Bhx0IOnXZRVNj
pFf9MX9hnVdpXQE9jNfCE6mhbMwAd1FuYJUa9t0OceMmGKlq0RvIQ5NYBjGkApaD3EW2ry/g4vlV
mXfA8wh4piLOVTSHreuUFE4KeJ8eLzJk/JlqQGMujL4H3KSZXFK8hW5KkCk+3RQDqrb7uJwqzTnF
YQNEhqy+wOO8aPSy7us9VjdirrOqcot6El332mUdsqgdsR5/BtZxod0dsj+Hh3KT1UUvvUYkalUP
BzxiYODzzBi3sbBRTU6pTEIoA1CdboZcVCu705v9CS3g2NK+T9KGJuYyehH20V3rAJb100FoOTfY
gdv+/+M/JkWztIaFDi+hbCbt2pjiI/m4VbtqVl3/HK5eGJmM9Oho5e7IJ7BLdIJU3ZmvgECsLyft
v7gJGapGsniIgAFo8fk2ltpoiyPnTozByedrdh9074qktM1ptIQ3oXSPmlE5NxL+vmkX1aSh0n33
8/TlOrEsWwOTmQIEDrnVUjQ5f1kuib2Wkhfj/UmReDcQy5D3DHIthHGkcOqwgB1Vam71yGCnIe+L
tXY28gTw3vXi7GEjpktpuw39mtaeMuS/0nw3Nu7tycVR9VNtuZlSMuVjvrxoZMthh3ftxbzHAwym
7xspTzr0sGEk6KErnFRpTNs6NU+/4rhNa5tKJfTuvGfXveCGLCiYyj4jGzRd1uUZQum6sjGxvHTD
IyzdDc3lc+cmsaat4H1Emunj7tTQGHatlR5jwNn0lzhgEFiQeWoygIbFBV4fJ3CW9fhlUGVm0q6c
ePseuLvLi/obgbMlJEO8e+BHancxcvMQ3Zv4EUr6sFRIg/c6Z7U1E+4L9U/v/54QDgaRgwq+8xEb
Qw8Cr/S8rI6LbFX2hJeKupTA/qZ/CsIgMi7Tm4RzayO6qbbuUjf91CSUNPUUymAlZzMPCj1HZZZL
Ml222uyUBBVQUqRfCKfKA0UJVvjgqxT7cNyiAvGY7uz0pz767L3HX4eyi7PAMUERuyuEC25MAxzH
APPH2OJmSkmRCy7w6DBKOJmQsxv58cvqIR2YNVTOHJ8lKH+WvvMnsvj47WP3z1FEU+tgkxQ/Xzdh
enNyMQu4EZ+hJI4VlnBjQYsrGmP2URVGeyiQuv83tYOmICWfiaOiHirdXcq40hPkMIKumLERY5p3
flUsLZLYUHWGO87N3cOon2NZ2p2kDMgGK7WoLRSeJscX84CRnuVtdACWAeWb/TEscPy5j62cn1zW
ypDHflhA0klSkwCdAbLZjuiUhBCOVfBtqoE8Sq+XHVUQuaj7O7s+3O2m3TgBI3NMauk7GWKghLEa
6FpR19sFwN4bFCYHsDQC/qPOwuVJYZu6uNcKFbO757AJtlvk1KZarXaiYmoYia15MO18ZGL6CvGf
x+83EquuDDiG7ZNWroWSsb0kHF4Ri88ZrcNsTyN2uwtNvsver6N03C5PW9k+Oobn93eVGuZ0L85n
/6mXHI4QiQaV/yfyw97UbWZLnxYL+28ifC4BU8tdP3Fmmni9rYkxkVduaSbLTd3x8ZKcbprfwLVk
/VvMsA1eHcXGgpQl5rnTfm4Rb1rFqw9JvyDeExt9K/QWeyhlRhSWR+nM+tAeWjmo6Kfe1oDE11Zz
9aMrtRTDjG4F2zOotFsuAmwT1RUlwDmARn85OteIjsBvvUUl0dCCrD7dK8n4j7cOnWKgEkZsQoJt
KpHimMHwCeQ3YSZQuSplhlGjuwHEX8WjqWtSuu+0PIL8Ps/5IKQkUWndDgXVm32hcnKGFOQ2TEHB
t0br31Ovu3tNXv1HtFYsZvZhtVhZUcW2XRj/vYY6x3x36SzkaTJJxFPfswROZjEPNwyFPTc2XVnG
DhKP7gzeSvBmrkty9X5NZK69FLzsvjwV01vEbu86iWPYLm5eZKY50Pit4oiVlUPzd1Esp/54jVlU
ZQFGqd0yzZCkGhND00JbXYn68XjDpqefqyXh72g2VvdrF9aTEIPcWrkYrI6aEPfwiMRznQCdSO/p
3YRHKXDsmMEJk40wCXnRHEOJb899GwP9L1H6VsH2DyVh7s+qxqvsZihzh7r7tSPPPYlBGJQwJvx7
QLHZhUOLWCw+CwaWteFMSlbGWJZBTKsmyD/7/aNK6gVCAwJAr5TmMT99LOIvWuVE/R3UWkCu6/Sp
/0dkDlPMg3kQj76imbi5BUVdwumwP0hSAg6qy7FYQ4j4RrzRqiieDK9sOV+RxGYdB8qY0cdjvYTL
vaj49u0kzZy9dkNnMIbyeKS2SZJoMZbobjk0TF4pFJ2QmYA3eIwdHB60wsZTNDpapVkavZb9MUAX
HrQWbFDLubTTYdE3TI+EMKeFBPw+Q3+zBUA382D1Sz3ubF0KSqT35cLVe/VTmqv7K+tcjVmdH/f4
bfHGzXP2iVrvmXGmWex7pex0YdvZ/nePZ2uaJ2pb5lToqg0+YQEucMgy6vCXGBUG+yZ7yQkxVLXH
wam5m0i+w2xaiA9aQZi+hlWPFyQrGW3k/3OXO3LIDhAI/yORKeFFvnULbkm+pqIvQ59zuuTDauBY
cs+INFkqcX4Aw7NUZLBB7C4r0/pj9L7wzp1aKba5lW7+16/IcTUXv+jP9qa6rbLD+dnBxQJCMd8O
MZ0aHw6xu91QGjQD/HCxCmUqrfc9NJ4WDXVViiyj84ZpdcCN3aCHz8usTCbuaUPcNYzKfglvt0i3
5SiJryHzlHhFrb7hLzXfSTXbpAGe/M0veamA67jXIEW086Wypyn7ffT0+oyh1nf1l839OhtqRbU5
n3XiCPjZIPnhXQfn2Fgy62UyNaw4eQVu1aM99PLU0m3k2S4cd8NMNVePpuEfCxERoPetupUJHGQl
rMHxH5wzUbXOHY8bS7rQ/OEnZ1JCcQDIlz99KqGr3p3jNMd4PyhEBkjKAzrYlYa70Ps2bq+y3ngf
Ik8lsfsoV3brA/S2vUImH5+k4Y6mta2XFfL8LYUgiimMtqCD8A1Iz6TO8DE13EdOb6CGR+gUs3NG
tZVgPm9m3hE4yTaA3xAMR4cH9j/n6+kSZ1rRy/3z7le1Y0po2lOCYCdLFYcvyM+cnK04oneEMfyf
erOlQOjGMX1b1JGb7apbY25voeMmckLLRKKHy4sndR5ATRdNdS0yk5jEgh3d7yiCOvJXnW5c6xJN
rWj4fJ232Vfc+0DxcBWengfZQuc1KHiUxX/IIgYNEYgp5JHz+NHo8XhYNlZoquNOhry5yxQ2GyyF
2+wfcKeKK4y14wOvwbMceGvvnaq+5FbvqwGoBEIDFxf+VHipW9EvKLNHU8kPto7Amih8NL+sMuCI
XF7gHtH9wRhOeqmZoHsO/N4GEXnbeHlJo3ZuG9eJ7ACNjI0qkYAd1T98haVD1v/j6VSikQfJ5QfV
L09/hfbV1N7Y80pDKx8VjKfIfgyRmhHs6r8m0HHMQPc2J1Rw1Uy4G8WQVM+Tl9HDwBpqSJzxF02d
yueJI8J3+KcrksJXm8ZLF1KYDcjlsTnHXlUYli0/Go85mfHg7mZmKz07BgT0gt7zolJSSD6lTs+f
7cEsgDB1cFK3aE1gfCGeUnJb3e/1nNvvTb8kbQioGG06rktpdiHEkYlvk8gz+oIHW8uJ6tN0sUsC
bIjD3TCeef4YmhvHTyvGbQB0Qy7CK7/dMHeYyamZYkpBnWWYgU8sEtmasm61AyIwc9IElniFE/XD
e6zR21vidGUa3a56ho3f8f3JnPAZeaGeFI+co6UJNSSoMX/MTRbr46TpQ+1yJcdWFoNr5vwbjet1
aXm04Jfsj8sopP4fZKUpAkLzgMzCEA0GPXGyBWkFBvi9amjpE215bv7z/mYallbTV80TQ/dyl9I3
Y8fGmg5pGA0HOhoMeFJxZNxGa4mQNqyp3I/3mAPHEaJ4uwSbaapCWZIbkejMcKOrFks46aTo8le6
9yZjW3Oxqxxy1S/zRWps26bJLS9kxT0Q9gEvCWBfZApSfKOI5njjvEeTwpVVHJRtp97yKgkxWJP9
SyeC3El85m0sUNdWZzSXfTmiS3W6rwag/dYoEsU4IwbuPb0FP6/3ivgHywLjiRFBFTjFSHZzvTZ1
IZDfusTkmGivwWP3nCHHxRtwRqyp4jezhu1xsmQsh4sJMmZL/poMgEuj1TfulFlJuRp2Gj2MNWYr
gHJrX2dMg/Nro+7X1kRTxQv88Q5BvoIc80pi4DjogzUFVdhMjt8mtFQRO09mibqz5iqtFQtX1z90
BlAXJWaCIr1rK8CZE67YkHdUmOSqfp8hR0Ug7AQiHi1HJmlRbU8ETlCkSakOg7QOfLV/1i78MuS4
JIV1KPAHuiV7or1K1AId+xoGo1SRENNU0Z7wfAsw4pTZahrBC9r43cYza+PoVctMsEp0v+QKTJaf
3GHZH8UnwQXJMaUSR4tNlzhHOUCc+5Ua519d96FvfY63pf6xj9g6NnNm/fE7I+pg+FuweM9lz36g
uR06B1wWgos4pj5zfHu932EJT6t5va4tJpYk+/RNrP3HnfsVSKHNNjY6q6PpF67w6DZf5DLUWDP+
PaAELwtj3Oi2OWcoaAq4lSmCg4FlX4+CmysfhmRPQAbkJBkAlm4SBxiLU0xAnpZi1PIr8IdaH7l5
YGvlcINT3zR/FEEPOMn4EUHqi+ehHaKMRbp1SkT+2obhsnUz8WRadwfqcHCOEzQJqdpzdlVpSOo9
EGPgpqzlylR+PaUzLJkPG9lWp4k/RwGMJ3ca9ZnTkgkQSYkKEsaFXav0NBI6QV7fo/iQhDJCOmTE
7+sbZZUtlUVl75mjumvVmzgL+dtztRIdHR5JYgKz1nu/twlstwyne/7ZmgQg+V5A9S4hBCLF23CN
tu0/LMsKGYyJ1jsk7Zf6G1HFZutr4y628m+Le1mDXgnHSxewIN0IcYFP7V9fOECudxp+X4Gi8WKF
TvJf7Q2AykL7BSORv7WeDmz9rRkAFr4rYzwQGJsmubWY4J3rm9orM90lUTAtDhBihhWUKxL5fFtr
GeuRAIhP1k0TZPV4z72Bn5JYnRzeHEhEa9ybFnS5WTgkCehv6K61IFYbFlLR9K4wAe9oNH5j3nRY
HSUluGsu5gy/HUbewBVsGSTLvikt2imJp10+W3D071y6NQ7K46D/FmvL/fpg2jAQ4QeFLQeMfTaZ
/8BqxjP8yXHFE6Kd6+nc5NdnaaRKW+yZcaTQygglNwi0IEXIPgjyES5PlBv2vm8xiaqQngy5Umpf
BOOk06q0pQI1P+Njpx7TsGybuct6JE0vsGXhOUtaLWl8CcIHTgZ2bSFmJxauczGO2oF+B9xp+cjp
oBTX8cDfhH9s1cAdWcAjZUNEqDMXQv0Eug0A6L8jiSJ+fSq3fQQ2kkx9XHais6pztqMevaFLqsKO
HeWzKMIzC3vUwkDzKHRchWSsgNsqVz/BVnUtdJLmCnts3PBR6+tzy6N3Vwggy2JabIWOqfp3Mgdj
Z33l1EVMZCZz+57DsBLGtFGRLTVZvtn3EMxP9ROkuHF78A7dQr2o4JcXm2WiMnhrJfIKJtjFyjhK
3W6T8cPiNZ1PYVTfy0q+CqJYeRq25PWbnMt5eQAP9tIAYOJrzj4JYXeB9POgMxzIBfuOVQlNPPSw
k2hye5mp46hh/zP6OElE76cBbKk+mk4DfOlZ8YoOWtyLpLSsYIcVoRBv8BacZUVQd0/G0DwbwC4N
syrKc9LdJtoV5++ZhRjoZoHKXUExryzfCk2hcdQSoGw7RvjY5+J2ACu4I0KcbhBWz8yobcFRqrr8
nrAqCJ5EoVmWYTAbU6CyYsklbXngkbMkDt2Qz6Z3PJH63f4sRtgDuOvBfjtJcWst662LKWBAjtiX
1UK+wHMulCIhPEwSVDVUvIss2Va0q8dLTVOqrOyA0VhLVM41UF/8Gm8jmupj8xZDw5jSj/lufzoN
+lKYLzMHvSjonxIP8j1wIILiiKHJQ2E13R7G5EXFKB7eXJ5hXkarMxKCNapEnhbrvtBLfKhfGXkz
LwwYTxpnG+nlf/juN7JJIN2cwXmzyUqTTWwgXewvL1Am4imPoucKdtJ54N0IpSe0zGoiOiZzFjMW
FKtQhM4MDLwH/1Jav8weFC1mZl8mom5bO+i/RD9hcJ1Mmg7uGYi5qJ2bAnmkR5zJHjmbOEdJDlsl
2/9NjFzRz/y3jAf+cmYG37ctGOCBG5Tvp+CMgQyKp/k3i1CmbsFJHspabp8ysnVAnA73+CkUUR42
fJl+86xnccI/7PWpRAanTCvufUgqKUtoHe+nuHnbnTHJKxo7S8JXK57+qxzPxhm9uej+nuH6Pxr6
JOQMC00uIX5+w+2TLPu7oxL6N+UCSMHV0mj/0gSf0D9XIm/HMnZdXjPgFOvk4el/LaSSfw80u4kf
IRAoTYq4HX0h02NyhnkDxLHZKiCJk7pC935WcliQXKELPkasDLcZHhjQjWsNiuFJomL5dGYgsyYT
dD12Y65ABfZGA+YB9R4MdH/+mZ3VHbX00MoPl60TfAU5b8X99E2InNmYxgis+emeIFT/eon25dtk
V7tjM/H3esJ4MOqHhYnn/ib7VJsqUZVxBf1O6ReEORQxrZDryB+Y2SWXIKO1xE3op4cOSzUJHHQ3
az3kbInuPcPh3Qwg30l8kXbnf0/D1vohB4sMzXdMbWIRyOhQhhy+AejR1BzIegcIkTRadPoAz9wp
TD6xHE5zfFh3cDQFNAv1gwVAu5oenGC2PoOQvVWwg8yFVpB2L54nZ2tiY6M8MOSHmP2fZJiPg4CP
TctPNjCnblUfiozp4JfYpYGN2RcTcuCdx31X5Q7bZcUr3rrlv7DoDDGaE/ZWyBZXKJGHJp/4E7yb
1l7R4DOcERhuhxSZsbEVlE38Jy5Cqz8DRQR5Kl1l9Ikb0EMS6n4bsyDMOkWJDIPtFjPKEen+v8sY
QHD1Url+FeFuXJ9FI8SKzy11n34QiFBGhhNniOZBnYUe+OdoWkHYs7vaxqvRnjJzxafA2/tpC2D1
BDW8N8LLf/GH2mf5u94V3vVYLQEZIlZM/SR8FlwFRKflgf9iL9QT5rAMF14UjB5j5H1FpDRIOicF
lGfKeGAZXr8BOQXxxq/k9zKeRJ/AYBFV8z91HQ0j0Yt5I9KRKGnI/kHsv/31yyd+r7dWTMphWcBf
kPBdFiK4zmlAckIzicVncoOTffZZw27X3in1SxFJrsnyn/NQHyPhvHr1xYl7Q4P8WL4Ganh24rYg
frRXozCcCvxjbmIPm2MCGpKnQL5qcaD52ogkAF9sHSprjfQPxWZBbLycLcDJiQbweQkRIIYeLagC
91tDB3xGxlDqONq2xuYdJ6llADEzn3H8pdNry+5JfTITBHCl1bA35K+/epHKCiGxQncvmRwGZLKq
Vqr/1sFOsQi6w4tGr/8zOTyF5Q4nQdYCjMMcItSq2JhsZdKFMdFL1lApZy5mPVmn2Tcbpv9dMcRV
S8uILn/yKUyHq6n8uQe72t18L+Q0OSHQ5m6dNxhFhlTtMZtqC8RvEehscuv3Gtgf2m6PUODSeXeH
cqlvtgBzSTb8idKbP0FhRER1bpRd1qTrDetrJF5neoLEkHB+z5OZ8huiW65koNM74C3KHX6XJtAk
+Eb8BknM/DWPVRTUEjAtIUKyYCbCVdNeo3vU2Q7WN+QmtKpgFLCERFf0f2nDV7S3gN4Q17+tIPer
BuQHZJorUBuSI7mn81Z7zi/AQ5Yxid52Qcd3oqdRbcdfXiKWoB8vNrH0Yg+G292uc705zSYwUitp
8UW/GSYKMkFK7pi8j+1wI2gOcBd9/IzabwWLPJIrkZyvEpiLdVaOZl/YZS7TfNXZ8RIc9naWwWpm
AznXpqThsfYufUaz3xFQ544JphYjQfmlt7Bb+G97DKZmMCOnoUc2RHc8jjZmOrqsBktC1RG3Nr3N
K+Ejye8G9irLssaRbA8/SJcv1eSFee1fizhNdcbBb/ln+xPXpq6B3UzQLDJEa2vyIP3ZmxMt0RTt
gkOzw9il2wImk7qBCsO1pWHHn+m9FMfp+9zZ9Ea30bGQmJghnBJYGKrrttZAMNTkDtaklt7v1KMM
gyv159IpV9grQACa/T56gNmC4o8Ad8CvzGmk8FUjtbn42ismA7EwTmuBJDikgosbxM2eL5LLaPKB
13UQNm6v/Vrq02y/ytj+pMF+cyjal0XTY2oKpxgYgCjQnY/s9PxF2LgqT4C2UKdq7FvVr62Cocur
0RD23JKLgSFFUtrKuoQwoOM7uYMI8VeGTKTJTbnSp5fNFRKVg/z8/Nx5pokWnjHgzGTFOpQytbg0
OzKgN24tEOph9fP6qBmSxrBC6U/7W8QGb/M9DKuEGoZSYCzyD0oG3QXr0n1AUO0m/r6eFjQy+MqK
dmICoFCUPE8VDrQbl9bshmCFISgfvrP3NKzB0ofT6epsC0SjBaUBp2cW+UtneJywAtXmAjR5PAa4
UCQB2DVeJGgFveHm4HPfRgCD+DNn7qzY5tQMhM/huV9jOBCS4inPaKrsqa5niE/qisZyHQACMPH/
goOqVkxAVxnPosTjWhhQlWmFGH75RN6fCL32ENpNbeUSH8wbbTkvCFUQ3ab1r681GEiph+i+uRkT
+HOd98QeqORBIvqZDMA6cBNjxEGZ875EQfVPMoVZQcQ0AJlKy/aQUakQa+NjkFkrLzVC2CxgWABL
x/w/aK+6Km5cr7UfMh+kQcjydXRH4yS9iZ6Bh2PTKaRWYU3SDZsU9tvGO153OZ30qnDKTWwZH6R5
+acQczi4xVmJ2iFF6w8C3t5B/qn6TMNrQaxt2O7LASOpOCuEjykf6GISiOj7JxiZEB1kS+08mFTN
phDlRCGDe9Zdt0ihVm70jb17i7+5YwBgaOiD4a6u8RfBqvaeWyWTAjpG8WuRmB93i6uVAFJm22qt
7pSyZG1+qVmUOCiF4620cUwI5S9OBTf0wf8SUty0HklUU8NqZZl+4zPcmQTqkLvRdGnk9NiHzdeI
24oP0qGHk0zI41jLysKsGVNATt0hxs03yW9d8lWj7P58uuDdYRQLpXAEVj+g9wA86vek5XC3ak31
+XcNm5iGUe0xi1hZWWThUjv+nOxUWyOPS7+W6tIwmaV4QG8A1s86DDOauwqoXHytjd25A+DU4sea
3cGDB7XZBlTFLDYv97780FFJP8oCUGWwloCkg2hnUavMxv9Ynjg8ki1vQ61xWNeCJPcJqJJUDwh5
zDzVtlPS7CAmxmWeprgm6UxNdK/5wTwd6oolff0Av3tPFPEsPGH7PfYrzDqTsFvSLnacwEPewoWM
AE0nbrI1hgKDV0ves1U/1K2/MrVvL4w9MUx8z8b9198FnMVpe7iNI/FPpZbsRFTBta57r+kmq+RM
B+C2j8PnTGHPnURqy+zGJvZ3mErm9qyee1D8cqAiDl9J7cGMDNkAotAQWfh71yfLCXCH366VqbdT
0YmBOHUKDiHvoh/Ylwv0bOEFrLNLb/YHXwL/q5TnGbCyh3KRyZeYVSoo4MJiLtBrywSwumDQEdVQ
N5YmGQPwrIsj+HX3FJ/rfOQs9P+INhemWPaemT22gYuHDeJUgEo6ryJiuiKaYneRpFNlpRTp0kU6
O7AKnKJvVsKse8t7sS8XDc+zsorCMV3BWkRivtOmJu4NJsQ89Bq8usk8v/Jvs1cmcdqcp/hByASG
UahF8ZAxfd+I38MZeNMh8KtE9+kcbSLddoBxm3qVa5D0c59VO+0H0AujX24rZ3KGan+PtdEu2Hyy
3Qr78r29mJ68eozuOIUrFGUReHG7szrsjUC1kmokpVB+Y8FX+9Qqf5darq9Rzgk46j2vKVJ+O03p
cFYO3evcKV17R/S/0Y9mWhPLOcan1fJuhfruGHr7dJVyR1FAoAgIj7rVXm1W12NqkljSKSh1As/T
ON025FY2T9vR2jlUHwwOpKgyJaDwUWfsbBQXzq9arLVgIBAu7E4j9QNe1KB7/ryHghIMaummgPEZ
YHhRgn7rw/zbC8ubO1xgxDFccwK4YY4Fj3iqTJH6n2OEWTEug5uMV3R/9b/+uSqZvfQ8LcpVg37H
nXn1/VcQ07lYZc47ifbuDXv0mF3N3fft/I+WPILAwpZ3mvMDRZMOBhqHwu/FtPT/Ql3d1o6/AaNp
GCjRgphfj7J06mjB6Vhr82yeBJv4MsfWuUpS1AtQAAZmx28e4MSt5Cky7hZgwZWuXPyhlMRzaNkS
bSp1ZJm6y7bwZVa3r4KDznaU6phYjqi3zXzBPt+UgLBvrLETbuJimS5fuTX41GNYr0uUYFQzd6d/
p+VHHYrpCFKNE6/geMpgasFCQ9w2IH9iJJoniFHg1gQKomAZSSFLdW6Lro4izqQCr4HjnxEfGJdB
JuqKFmCiNADg2lSLHAU797uug02Zxq2Xw4vo7VqoNBHTceZ0FI5sHLY+kPSmes+F+pr8CKtAHaOu
WZscYku2RKKjquliQ2PwKWKBZm49V6ebvIJWz6r7fx8otXe30BFA400KpWpH3mlx6fPbWnU146VW
1hPVTRoIHZUIEnH24TXukbCBKYAjpKHLnt17XPPc9Z5IELzqzMf0fipa9qiXTM0iArlLfs7oJlGv
/w8KeTHdLuGYtaZCtJ5vecA5BBmIZmj53zAdwq5VA8pY2igckac0Vo2TeYAk3ouD8xDlfWT0IRwp
COVU3G0LHCgDCj0JuRv5xoBdR1J8ResNmsKFBIGreIvJjkeBe4k7M4ZemJ6lRwSCjKrAW3cY23t3
qaEvP98vsS/S+/RIA2OxL7Vej27k47nHNN8SdMvq8ARH/lWynxezIs/PGl6OCeLO5zH3sPbVj5E8
oIb+EHbMc+QrsRztjYQa25VgHcJb6S93tk/k8Myy9FzfJzhZa9+l/pW3N3Spdz+IAz1R7LUAM5oL
OKP0NrkXD8QwEQ8su5+pbJuIWWUwihqTy6FLIA6ITD0fWvY3Ypao+da9l2oF10A7Ammp8unbzO09
ZNgeEz7dNtz/o4h8hzVAp9pZ9g0tWJISU7e5hVvmEEUi3VjhLJJOdWlZIaMwrvEFSNMqJEO/zoRQ
fsD9l4jvwjaLXn2xFmBe5LbmAH9wJQBaHTL068eYI+cCW+5FtO1egMAcMoig0mPyqZeFQOP+dtDr
Te/6k4vQ5a6RyWmZyMwfWunIML9ZNKyJvTpP6+RIQiqm6G0D9DmXGY0dDrKowd6ylnJq/D6HDC3O
G8dDYj2MN+2OUGizUu6GXIObguglp/0d0oPF9lxC3F5o7gzqNh2BlVBGzjKXZxvyZDQ1SAE0aoFM
nUr1ufrYlRyqzz2rDHwgu3TB2IAgWJmaQ44Ppg2vb5QIG5P9IUJXuNUmSVtbiVjDhD/TxaD9tVrJ
ldpXrluAmJ/H4brIw54oWQpN+9hKn2JzYkhjjdsmlXMhxbEzECT6rB5gbz3GP+VC4xf/lQpO1ZxO
+lGp5vfTFkDw5ynxYC/DZfou2z34S+QNQvEiijpfaI0LbQJiXbIxObRe6tfGvW8DY9jLFgtcZ1oH
ralQZ/0CBNIvlfcw209pOkatBk8tTBuglIu9PybJ/+0npCH0st/t/XAFZPOnx+/hIy0Hyae8k3OQ
8VSqsEgCzTubdtilrWVZmjZ4HWXM9nj3J5YJjasA3GIFCPE+Qw3E60acTH2S1HJosacRLBHCJrNl
ZcsBFWi/TcykohT85wNl/OqIewEXGodrHMWGAYxnh1LXwCie6K1WNdJPfJQV7qoUwmnnVpEb5l7g
iWOlLSpZqc8hQQy0q9MDLHSpCo8eM3p7L4bFA71+YjbXHYOMyLbdB64oqNbELZMFEXsyBlCw5n7a
+B+xBKodHrxj0Ng+ORMmrqh/zz47JRFaUQJK8z20G253B4b5m354h1OtyXiV8+JCcedDUrAlPjyI
dko1q9xyHa6PZOsaaH+Laqe1/WUY/1dfweWvIK3lQ/FWysqbYu2Es2F6E+jHhP3Td7/gVVqMXbeI
uQhrlr3tDV6oqCnBIEV65yBO1FR9ymuA9nnRcVgsUuei4yEgxl8xEit4roFFuWJpx4TsxzzpCDMJ
2eJxDrX/NcKNmp7liB2VPgxLXR+HEus1qiPcEoheEuZcmLKlpozLHVM6re/ebTBbJZQGYhfAX26j
SNdJRMShtVBvmlW0hZHIa2+rFkU35QQI+MVtmH7E4LHF2sXodzvGcIr4RHh4xQexh46jdDSYX2uY
SVFtBk9E2uGnfMs1vC7apEEpVM/c/NGBLLyLQdX2JJbewjDwPwZoeoARGqBMRaVKFKqcbpxrGvAZ
Q3yiDFiYNHnwN9Nkk9bYRC8QMBSs4Ju6d6SyHw76QCi6V60fn56D6M2aZ8EorGLaHs8BXaGfv1gz
OEuUoDYHID+PMRg1Tu3/ZpZ7D+7lW+hxv1EKpnvHHTpCb/bXcZoHf+HC9Dm/GLz8Y1gcZ3WzHgl1
KiKr79e1YyGhGN6AMNdEICvWo+BiSZhfEs3k7D6nrOxVpILtF6i0aoNC0ZN2zKckOGu7zbVyvHXQ
gVk+tun2czgMEX7XLKQhLh8bBpg4+JBZ+oCl+X8AbUAqfpHgwq8YJZ+NNqzgGYwz7+k6T3SlWHMH
20grcgh8jx/NS4zCqysW6mF8NQ41XN3wAahBSohQANXgjtoW2K3lm63h7zEWc3MzV5yF8juA2xdw
/JXbVlxrakje3GS1qGvAMWkwaLCI8eb/MLv9WhPKpM75mRi9lKjJTockcKV8K6OBI9d7WKpE4d8U
69szTtmljOb14M2mMoSTFyXSDGOY/azJHE7lg8JpNDdJM82ePaaloOhi6dT/s5MUnx8rjMAGWGfL
jguqT9KzdCIzR/Kqttdw7yoHsZWoJ2IiB3/AcPopYS45Gorkyi9SZKJYmQZva8tVl5xtYtmHzMh8
ePBKO/xv0v/cfGs11SAa9DE2WYxrHdZUofNrdXFImbVuMWp49QMOPm8yL9vQp6zn/ybGJX3KS6zc
fc0UcBKlL+AyMUf7rxZxuPatVwiqcB+icVbPpgTWOCriO/oqBT6zbuXtFMqTLO8AnbGXIlZcpFEQ
nyOjFLbJ4dlcfpA3K6GE9DxtxqMpwtLPYJmZpba7ADmJHqRtTUPg+hRFoUGM7Ba9g3+mNFqOr9zy
u9vVBTZ78m2XVH+rPMrTWKHR2mwW+kJqxUqjIkZP1h3i9mkkMShLpncf69RLwHyUS96BIo9wuCn7
13cqh+N/EmoiG6eGQxLRAZVO7eTmSV/pXyxYUb93GYk8HR5bi/iXYlY0oF05OixARWftdoirpZVS
5DSegEO01wKKw0mrQJ/qzn79DA8Tl+uVhp3rNhda/dvFkptZDrrOI2apVXgnYckv5EVSmhFOQ3Zk
hbYXk8L+De6naJMs26t96cY2GD5ju2dfLgKhuldFxfDV1R0Joi0Vhg/Ibv81k26vJ/tevr71JtIZ
vX2oKZqsdetBQIxOW377cBZ0IOPvTMG3ZsA7NGOcFoXrvWajLmq+s7oPojZ54UZXwInjs63Tj16z
gMKRdtPACYzDDBdF0h7Gu75I9ccTzEZ136e+cJh/NVleUGtbs1Tu2qCC00iBO8LHar7A7bcm/ChZ
GqqBQFvfEduqBDnpT6jHYRUekZtNqlyJ5XbA+gbQ8UbS5gnqaDJIuuz/cwubs8MwK1KV+61oeJ7D
ZKBUbR2D1jsGzs9/1ddNndYdDf95N05IRdfTC62ylYn5R+hNuXxbP3O19JFz3mk8p5Zvu4CSLuHN
HpXyVfk2gw08iAuAjf2UriwhPavs4PzfxvsPOqgLUKSUxu/kDFacVkQVuM9+ZiM3JDzsELTxbRmH
9cBM1CG6MioWh7s3cHWeirc3zGdyrHG/fOsvktwH3yKMUkCN7pjp8indZNkeV3HRLncJEbaM8/k6
HRiiGMj0kqkWFHe9w0FpszJh5dv+AJUIJh3q/wN0fc2inp9D85SB5yMvVOR3Oraers/9r8rdZP58
Pc9apwhSGmWSwZLs1YycISsO2kdoKH2EVqCTcQcLvE8AK+k03+DdXKvPeAAI3bDAEaKE2BdKGOlZ
EVFZ8tpXydixzzIaG0vhVJdQPUsfAdDwi1sVj8Ir2ev4VezlQ5ZVKESSOfpcAbM8sPHlNBse3X1e
LNkVa6WjqcsoVUnlC9wOkV5fDLs250E6huhL//mh/cpZf0Iqpzgtf/MKR6Tcl+tP+J9IWvDnBdDe
c8LE8Im0SamJuKFKDxLDPK00CndebWhwg3n0XUaM4KBDXbV7sx+UWkwRLPVxUccnfssGPhQTUT70
6uG/w27IUrdU7j+ZFgesroJakK0ivyo5Y4RyUo6HHWnTUvgRJusz/Py6RD9gkMWQWUrZ6K985Sht
Wk+LAk1JKUEduuNIc7Q5cMntC3cbJ4VSs2ySRjdQC7HzSWGGDknHWMjgiGdnHF3bpry4rc3+K3Gr
TyDb97UHA5Li+a76fF+u5eRqddbKMFxerpYt7TXiV8RF69TWDNcL/gWapUynty2z1QD1x2W16V1s
TZiP19FdsuAh9z5e0o4w3psFeOKHlNuXDgVvDuat2nM9VvLi1t1sFoo1GagRm8K9aTKjkEjIqd57
x9D7XRvbyuSp9oEjDo/hZ47WtLZ8h1N3FkFNx38s1jMjHCUiM0OGg8cQx8ap4eNrCRQiHNR4ZOo+
GDJcFOozyjsw4NsFqbEqmDD6oSKiFyifbRAK6JpHSr+ZChiqoI5eYEKUDbY42jMjKk8nugbnOa/A
Nw5k9OrukTPSfxwehcVwlFpJkZE1Lsht0t0AGtd5v3ucfPiDKYwwinkKjLeRpLiE00NmxiiGhmIJ
yb0qLAPYeu7frQWLduxd0AC5gXFuOT3Fv5uo3eCpfBQNNqiOWWhOxGfnOutByUl/4Gjxk4IbG9F3
F79eQPz483pBWCjmYFnAPjzvcV2lSIQIjKaRHXm7gCZsK+rVqndTzLze0/hEesfSh9Xr75ZmA/wi
hxmflgybJ1gILiy/+tiJx2rlEtFLAfGkan7BQcUOMw3Wa9VqTc0K1gsZTTiwyOEmZcma9FduHAr1
q8HZZtv/cSrpXuZ6QmuW/ql4+zLPlD8UyXkPlLNEpz30DLRSJHKSawXDExk1N/GzioRmQII0FV7U
mvwZMU46LjQSBcmIGE5riQXudkOx21eZ2jrDCgJS3lZQFovkW9cTSgBuS2nYIlHf7M4Z+VeD7/U0
N0J/kYnU63gykeCtTILXzu2wVWF9XT1vAhJd9ZUvQVBzDBzbhrJ5MNFf7gkePDH2InsYNKclJcBq
c/vDlpSTCaM5cIacD3L2XpWNgevsIsU40a84V+HyKNLQE+hLkkb1QL8ZK3tNvKNord2vrme4jHJH
n7WjPAxdUD/1Kcnjl4YjXkyxQWPlpiGtZVpg+xggdP6MSOP5+3XZA00KTve3/T7EIcTVXQKHF3FZ
EjOE5q1d9TRGk6KlOcJ/L0mGqdTF4wD5fvrKgIG/HALRJ+TncKozce+1g0hhOiydFt77hQkbcjCo
VZFN75f6lGXrMazJKdpDVu92mJk5h+VQZb2Egcbl9Xg7WRzrFq07mVlUP9BCBh37gVSSpdeVjwmf
6Pe+71CaEnb1xZbYxSm/e0ifN8RbobN+yh0eRcPNI5jJDOBJwc3SUBJ+KM6x6pOi3f/ay143Qdr7
XZWqKawnwONFmGVctAQnP/jOdrc5glwPvIrzksFCf+WgRhd8ZY/qkdq39mYhcAWsNK+WVXzbpdcA
O0S9oGUr8bFOcj2AD9wgFb6hmc88XCzk5FhZtZhQqgNup5LQTDL6CI2B57MczWaedyoRXR9Vs/Rr
ltwyvgUU6d23oYLjF01unAkNnJRCdS95BN6Zy8xRov2G1IMZ030A5rhKFdd05hR3fAzUaZAU3q97
qiMCfLd374e4GaDHgYDHTVda/rIG99qfI1w7/qRL2wsCJ1n5G61VTZ98jmax4CzH2EUZspBpCxKs
A++xjkOlYi3MD4jAGrNZGxFALJLHr+yDzY4HzPpWvVN4w9T8+crfkAKvbvlhcj5BlkyrFqS0hMFA
uJyC+d2g27hMTErOFChGyhAUI18gkFUwGuOw9tYlonXQ8yo0t+WbnimHmSLSImZcBaaBNxo29V37
437bFxP5bIKlQK9n/7v/TWUpDxlQK3Pl+NC32vuszYtpMoRmdn+dKCiw4KAZlgTqO0Yqf1vwK0/b
WA3aOWTh9IIk9zK2XuwoTcZNRK6Cvf5HraL1O7lZfaYII4mWpepJwntWJUqTP5Y1e6iXFX1pmu/2
k0z2OW2V0tTWvdbbVrVtLCr4sIfTOr9ViL8WsJgqqTWFjvy66OznLD/lythkGfx3YjxyOhYpEkn8
WrTkoA+dftauemnEJbpDtZ5j7Vpl+a+waLzQdTl6+yjVTko9/MKYNNyRHL4YX9B9eB9Du8486jpY
NCYOmd8/UGi0g5Jb+wh4a8Wdar4igdok/4N9rWThfulkuN3lgBO68fS60TOvljcRnElE7Dv8A05L
W/VC4XR5g7RVX7L1lA/lzEuhpZNGltBKLTN1/YKRAWHtxbszUC1+1fO22YMSzf3tXwKR9w9pqNUg
6XhPdFJhwyDGPjuTsvjZVHu1i/X2t+HeLVL2NrHGzOa01ePtvpnI1S1Hl69Dnfi9vLehd0nag0aO
BxDrCnkAWJosD4UoewbVNDepDHnoLhlVbMKUEoGDgQCvFyF/8NpBVxGLX985/S8jPgQvAs5+0Gdl
YJHObQXeHMRwQsOG/bNa+XWDjXj05PB8in/HLEHt201FyyK0Q3pllXYJpfuGC6eDEVbJI0peI0AW
C7d096/hmsUmnblR0AHu+Owxt32uUsOhiQI1xo32VjTOXo7EkC5ly3+YTyeH4kuc5sgn+GLyd14a
u8aUKAeY72GqFFNHYA0V9OF7HIwjxrcGl8mBdD0i6Pw/oeE/5MSFkoRjO1Nb3hMMj2rXG0hpW5sl
0PUCuxOGXyjFbu11GQ138ut8jSxD1QVTqUFzPmYf0cY3ErL5zDF5P5bQZlWplWo0JLCjlpxji4pZ
hyaA2Lz//Mu0JrufEPcLKkq/b16J3V+VC2oFaJY85RCRpEfmRZuAH0amfwE3/NMXcFICJLA9+7Fu
VoqXxcFKQlBW1IYpk8BgbK0GuOWMauxxrxhlmhPZ0Td+8PJuhmJ4H/sp2yN2GfGbGT8txzF3rRY2
RsoRHpsNBTo9QRhvUffJjKKl7hNkoEiVFYeCbG3PkpavYWHkAswZbQrnz7t73YOZT+/RbwY9Ew9g
kZVQalpZnap10xrjvhfKkP0v+uM8ytw625NPCOO0EQkS9LUN+hAb+6ygvN79z/j+Wx5MMq6usEs1
RNvFiOBNwMbdhjZZ6IUaTWqLF0Dh6DMP9wPydfJ4jrGEKDfwm2asmFST80NCregfi8FSu99lIoF3
XR2bydHbVI4hfn2aphg8aOQY7QSaDip/G+ovPCCX0wG7ilWHVf2CGmEBqH1P53sVvYqHmx1EpJOq
EukTBdLKtthuUCnLuoan3jqAGpMX5oPBu7lGNpt85EYTGg8UMgUcbPWEsVvtC02cHe5maOqxENU3
Okv2Qq8zJ2WxNiBROt7db/ce29L2v1fln6Oe5HtThdyYhc768k7nbACXQ0ym4c4sjes7R9rmkiQ4
w3fT5ZCOhmfKcVoPbB2A/y1s8qqKHmReDrsuVsGYyIKxLC22SYgQJ3Vv/3zRTxcaNNjMRPXlEHPG
4DVS5R4wE5MNHaaE2p0KVLDV0gH7HyMMedj6K5Ng1fNssnRM/AkMyxGi0AvlWXGz3bOWCMwZKErA
j+UELrMHouu/TeJDNiPdgquInIjk94Tg63e3Y8m/xR3QZpg6iP/tGkh6hQg0+tnvt7y+GJXI7SdG
+E9tqlZh9NcvP1iY3Mo/D1bMh2pKUCre6D0Gq/qT/xzZayo7JbOoGpK4dFylMmM0/MECGZinCFxa
celam5+BBQ5b80R7SxtbP0WY2qa7tu3WeobNYbNCx2qI0gG7d2nMrjWuJxR5igqRoNLzfdJoK+zG
4RiuHK5rYrt16m/shdVGk1Z41cZwapDyZNFlar7KRNGuJ0CscNyRPVcsTt/aneU2Xrfl48Qhwzcg
aKnSgvm7GxgmR3hESpvl4D5OaZfANCBHRzPGQIn3JHVaX1aEekS91RtMXPuoIY2lb6/JqtXzGpzq
npJ2MXZXca5KDcBj+ELMSmlR0ZbNVVDa5Imu+iHZYZ0JD1fEdZD+4O1deZvCf6jn7G/QQ/4byH9t
nm3bu8RuWS4u3jIiU8AExcJpEyDDzgEa6xJyAcSkBsEaVac3S0zRMUiA2RyOvHAMlaUwVqnYkFoq
35SfwCPG8OYUOSEAYBXRCsx1lGBtcn0sYwufy1GUbLbGLOH1P6+djOAeUptqfyCYv7yb3En7JwrN
vZYbU5FrG4dvmYudvFFf0PvB17WPp7wWZ7gPjM7qceSyEgf/J39QlXuv9v73VDztAuKku0y2aND3
uFJFSYu/UbaaiHQCSme0mANqGg0BcOWDxTsjKB5d7NJiBkvqQMnrMzhcwH0kIKXgpOTBO5JQWE9W
812T3oWaAJnDo/+Zo2uVWBZ5VxFGy4sy6z93Zy/1OkZyjCi3wJbTX8lQEPsGgo2yR9MFQDVBniNa
eUwQ0ldUsUb4W2E3snasyVmxogeY5xpFjSNHb58ity8nrPeNkKeFlLQ4JMiH0ku/AhOp42vN8BpJ
JHYqwuIultQhEgbA7fBa5ChLtqpnp1wXZWl6d5NiBoMtfN6nKwCVhpVVqUxzpFfnGoQANX4lTWtI
Xg+LiSEjdLN9N4NBaeaayLQJH0ICyDFYp4pXcGMo80CfHoWCvyLYXjIASMNiRAFexE1Dd+xMpFty
iROSVwPJ8Xugwxdp7GrZyCBGrp6jYxw5GMvy11NPapXhdDH4ur3jWIhXHIF5+4JUO90TeYdJBSOe
bPIyI8PbQhTaDfyyj2CJNNlq/tPlAra+9Ye9WF9FP0ru4ZQwh1W+iVU09ZqMJXlubkfOmMPJWkGA
ghm3ngZGG6BjCgHAKhcrFLa7m8u6KH0/S0enzCJ7fLuI8f5WQKJ/97uvkJOg9FkwYI6mlBVwmM0J
gEtIZS01ipCsO9+s1zz25ZB7vn9bDHMpzcOw21TJxs6eIhWfLOxHo4y15Ig0yBlE5YIfZXG40MUh
zP8114ZRXIcdX7TUtY+nVQTUsETCnFawFjLM+e7bPuJGoezKEE7nTRQY+FqKAh2G9YhLpgPGM1u5
3Yfe2WzTQIGgAmNw+KqUpE/DZ6x00a69mapc2csljGjTK+jm9OsDc42/TEDNk+iddLFPD9Oo3Yg4
MAMw/X75x4aJxc7WHTYXGujIoP40ywIOajXnHh/LwIE0gLRCEa02XyiZ/NhdA8oQkNAd9+X/DENE
Mos1IQW4RgDnktTclDov+1/7W1oHxIEynhXSmg54dRST6qbddRF6HhGKzo6zKABSUcw8FgArkcWo
wxh9B0IdG3RsFfETTWLOf/YQD7TKTqUlxNK54t9hABXck8TEUYi435ZLKa0Kqh9OSbRS66VInPar
gtAHoOQ4UhEl1OQJ+lJsrj5TEIynkpTAOkbTcCVsBSbngE002nt05xRVECVs7KS8rEWYMpLhqBsZ
DnBsLOxBrijAV9s5Yk0Q4jxOFdvwf/q2vxk4kJI2O8hrRT5wLb8lZ1DslGbuIU9yhwnqpgyQamXM
ql7WUkL8fqN1LEr6FvkORZFohpfIoFyt01fveoVlO5tEL3vNdVnsks7SjZaPxlQELbnCsq1sS5wF
0eaCgQqcxDqy/Qjw7qG+iEqJzVLw0Tkq2ROH2aqMMZMlLpXiYa4IwE5vQ70WGwbH6FfTkdOUfWH0
rGuks6eRSsJE25tCyX0P4cxsG6q/6HBCvacS4mGrHNNjNRwy5HhQN51Bv1vM0OklaIt1tnp8arw+
YM7/AL7HI+RzvTMm9bbXWypiAe7bgaZ/ruvzjppoqBxWvrN+u8cEC/+v84Ijh7P0vQ8Ze5p45hOQ
id20qEo3tXletaz+00XS/4h47av32dNpYq/+oYeKIX08vFw8OByel0HugSi+S6M/O8pzKXoeXBTy
A8hIWehBr6gHoDtWBDAtMFUklkD4Uy+X7zemm2Ky3RpcWMDMcrtdOx2Y4+lr36sRNf+ykc5cAXfd
g0qZ9MhLtOIFJa51p2de+GE3y+vGwCIIR3fvHy056P4dYSBdGn2SAq7c8AE+LRnqclbPxsRcQSj6
dvUS3mHuemQkSE0x0z+X1YKpZUTP30om5uhaH+uK6qXdywbKAYw2Sf8ja6a0o9818YJYXcMdDX9k
xU9GnJLc99U4iNT/r4+9zCwjGxqZ408vHHYacXQqeoU8MrRTjuAH23C4rmdMBxafBXkUeIl+XH17
2MIcAI6nQFbciXtFEKInSw3T621B3sOwRINEqIkBjfgMw5YcfIwPiEWaSGJLz/mafP5gP8uSqYH0
NMhJa90p5MzaUtMyba8ZE9zwyhfN+qTPPsmn10nLr/8pMDzrOM/OZsp+DEjSn8XUKXIL2iU8mmcD
LppwxpASVIgwN1NAsbkp3vc4yq35JueekfneBuCyuVK+/V89g8rVc/nJ68mvNnyxb9/t37+1kZUh
kjn4/9+B6At0HNY2MH2U+RbSRwhtPk/e3kiPKjuK8U7M7bV/D0iEkm1/WtXQ3tKzJvlsAiOgFViJ
XoQ4izsx9FZZDrIGgio4PgnIu35iK/Mqw+BMbCXfUxKdrNv/DuAhbTErplkotnVQkAhnczLfx3yb
O4bzguZxLev28vG0Es+Uh0DuMTvFKb/zgfDQfVAYwrnQGaIBd5JTji6egEm8l2ZwAacJT/BnX2gH
fEa7SncYkJ7MyEV1NUHEDdmZrDnC9fqejj8C2lmZ6clHjMey2JH0JY3FEFsmD+oiVPfG50H0DufG
5RrbajV+P6de/nltkszua3oWXUlHirsp0pWmdhcqPKJuk79qw+8C7vx9FHk0LtqwsLb6PVbJDHoE
jmsY22yng4KmPMoOQXkD5dpp/IlN1JkoT5PSWY7R2R6EVpYOy+VoGz3kmkgYviKULSCZDI2ONfh3
CF40VBHeeg3k47K3R/ww6yFQC7GKhatkyhLqlACl9b1Poeg1Ey9PHI4gbcoYwU8rubhENCA8o6Tg
6MwKU9TIhsZIQlJSWaqkvL5WllyzBBX6adip/miMaQs1P+UhzXZY0l0FIRu2dMiqPXDAlPoinhdC
70c/KaJrhwjSw1y9esFdVZ1PhV8R2aWNEQ58a00dP8P+CXa2MYWBjdkrCy65Z361NMKDRuU/a41n
3pdGw+WkeQ+PRgs25iO/sR39DJmqlwhrYWAJhUsMNI5a7023n+PzL2ysET1O0sO84C/m1EM1sbHh
NLgqOV1rjboti9U8wvO8su/++1535yN6vEZmZL5P9H5JpeZpewfDCqT41hAHxrF0t15zDzbAAfvg
cFRx2gjoudy4MaI2KgO94PcO4XOzOS4zoQi2ngl4s2iHKS6Jg6Ri3qrO9XkRELJcDekg1G6QII9s
+yKZv0Om2RoFrsFhsX28jxJrasS22Ewh3zPHMbhUg629hX5FvFZT9NIMUYxA+2+lqYnVzqRPlNTo
n21zX2tXwhNgK0pq818LOLTyzCdUOGkxNRS1ISm1bK2SgBpZqAlCnqy8n59NnDt3/pdLPDPlfURa
WGjug3KfbAsWHpfjba0BCdsIE1pn6OdWQhiEHbbfDn87wlqdfiYhAkJ+mA4y+gzpG76O6mN6ieM8
tfFNdJ4gcx8kRhf+vy3VpvJbIg6tLiDtifZKZKYruMmWreUKd5pZzqgeeCnVLNh7nJzRrNZPT+PL
zzFcCopfRuSMXknGhLSQ0WUdtYlgZF+338lWtt8YSjY2QZn8dFPVmlLV2xiQd/AafIAU8stxYR2b
WI1aQaOWvsVMiIJ4iRgQwBTRza6GVbPCKFiChGPF5Y8nx+K25VBoFoYkMUYOZtYTxomByDzyz4lc
LYe+ZUGyVGUe9QGTVBrDwgaPYUuTzPzNq0QE0xdlBfCRz9NG0/Chb5bmTCYlvVR0spRpH0LL41qQ
Jnev21X536c8+hGC16ndedeFAxmVvxZbWa1ar5/3bZUID6Usz0HYMvBSRjlynKkRYuVD3j2Vxy80
dEPQ69Vc3MrR1B1nMCA4UlqZGTYf33tOhj9v/UpY3HrdnHb+f6IubmmXhlxaIRENgyq4i2a3qX4u
zuH/LfCdWGBdgyg+WTd0LQTBbn6Ti1q0cDTN8t/x1Xi3GFu0zreMSSXDkvkkOlEgjJ0TPsVBEsE0
82iOKFFG5oQm2YxhqQ4tK+BIm87obqLNMcJystmcQWJv2w1ugvvgV1Iaognt43bvHccyg3/0hLOf
+4bN6U9fJP3tTdOnS/TrksndxAcabfpNKgGvivErcloOd9iok4tZbf0kVd0QovPh6qpgQvUJe/Y8
pxtthEi+RwkdZxjlfWTlEdDDqRavXBofV56LghL+jRgScFAzzxhmtpPYxgfRh1h+nSDAl0CW+rAc
NwW2czjkucOR2n4VwAD7V5RuSEI9D0PBV7ublMQ7QrhxGJsmPnd4BKOfjDyCEhYLITGq3FUb9U/z
6UDwxWBgGZb+X69NfOZ2cGjBeSS15c3BVRnSAM0SfA6kkPVtktCN69d+ynbKHLAMa6Oj9xF2ilYU
vLb7in4XkK7dGLrbfNniqyaV9HimOIJlPoNVrICbrTo1fw+L0ekXnOmqab30+u641h2Pyrcm3jSW
nsZFsP+mtPx+b8zkSr+pyjYBePcRmzUyYcVgN5O0K5d7DIS/wOhO6p2u8dYkKWopie1Xbdih4WkY
snJpWfVwIMPV6uX4Uq5sePUoY7M3Jn9Y0M6eeh0b4CZHoyqNTuJ4MhXfNt/a1suvUoQTin1TxJtx
D/sAMpTAaapc2yyHJ67QGN5wR5ZKwMvijumO1T6VD6MCdL0H7q6/tfacSNWSdz8cb67bNAuqkK7E
DiiU4VMS7/S+T4nHkyeYoKlJ7EEtkvHCraLkAZlSej7XrvkqmeLHQhI5cY50z46Avt5ObEKyiBT+
oeLEOEu6aQWJIWTE9LecSb9NdnFge0t2wrzTzK3xW6orUNo8SgOHldX7pHC+K/2dQcumDCOWTxFy
+A3vVefe/nBmynyj+Wz/t0R/jCaSVB/UEYQmmnbx7UcLWjPRT9X95btqaw7dqLvaYQ9Hrckhs/mG
jX8zPc/BH76X5EmiTqGADyq2r9PvI+DHNIug1mn6Ia6UGNGYC2udldt3SD62CW+DpHH3Rq540lMa
9MT1wJ2Roi6+aKYgLSvJTE6MZOlCZg8y95XXgyWLiMLsMfri594B9kI8j7LzHAzczRr9ZWSj5Pxb
QDIocAocMw5aVN0R3BibRleohDZpBPuk8rwORKM+/1hfs7ByBwF4B6HahwOaQpBpHDoDRlns31aG
fHkso10o5D5cNIbpE61EZke7mnuZLGb+KNM6bhpFDA/EdKqASjX3YAGFviqQayBznaH9ZWTIUbSy
CuOl7CdTP+nAk0qFb8E33olcn/czUUxulq83QCW8Uc5HU1XbAYfiVmtsMeMmCeviUywdzl08TrQ8
opCxBvvlM88Qm3hxaItBeszq/FwTmRsnbicnkCPnZ3cURqDpttTkF7ktKNZ/qH5pQ3Kzdvuv9/Lt
PlbBzzgUdX30rW9N3CWC05mgN3tsK/5XSBGB5uXgt9mZcqN3IATRrIMnRKbt4e2c+bqC53deKywv
JMpgCmWx1N3zjRUe/pnt6Ev0E1YzXQ3e1Mq8w7cx7qKsRR99linurXIJOqy6pquyEU+pfsVLwwEo
k9SpK+aEGCeqj0yryMan6xcimOdNh6TYxOR9HW3JbLrRewO7SyET1ZhkN0il+uWyYUzRo0QYTAuV
pqxtCHfanzPg+H/bJd65m9BMzYhmQ3/aV2O80wYtihUAGQ5InBW2wnJS2uJKbQSoTCRp/IRAAAPw
pSsdNhxuSyuBwHVIQHDGz8ZQ2O4Z1xCJ8bbvntL/uCnjmtJh2G9WY/T6ORN4fhJVikxAbgQsLZv8
ahCHnqkOv9WzEsCiQW87+5GI8gXqNe4zWqbCc5yhnSrWYqc6UIm4v88whb8x5PSsMbmQm3fONaHw
mz8bnWPaRrShp0NPYrIdpSxVV+y4AzkqGU2dV7Ac7QhoAaXaw/8A+OF8tsHBGNkejvcFR885CGGJ
KH78YEjb/2s9Vug8oxfpyW39ktcxzUDc+oG1PFVnQsLbZ/YArzAK464U0iWFBiJjkTFyVlo2gQ4i
EyKZ4ohvy9sePO9gMMI+s7x794U48djkMDFjRD6FnkXSwjKaveY7PYd08jkHB9rjQcAkKR874ian
FjmOoR17ojE8hunQrXF/gV+dMnZ59KcoAcdPRDaiTT3+kjZeZHMavl0jYND26WCtp4q7JcOAZweY
cleNTs0axoPT5eDei8JvzmREfoBxLSrQE7jcyywE3f1sWrdrNcEbIjjanRnPQhx+QdgHOSa0GNrf
U5O+NmaTlgk398qmoodOl0fuN0NAgyOj2YbMGo9G2UtsmJFmy5z1saS1vDPJtg+5ZSQrDcL0rhvx
Q25iOx7gO0a1HNXe/yfYMD67VW54wCO9ntYNtkfVCz5Wkx/XpVdrE8nlA8B7Hl4fq+ihygD5QpVo
UWrO0dmLiTzuG9LPgXMJyVZwhqCUbo4CkWIyU/VDUcHnw7iRZ1NR9nApZSbf7EJ3fp/ywxDtobEg
D3HU41DAqKmDQcij0XODOSdPh7f7RA+QbI6LZhW/656DWIhlUB4Snzpwfa3fPX1RR5xKq8xoue+C
/J20kglrwrZTsn6EVGixvNF1ixi0LPj+P0guAWdKON66cdLsaIksqCWffTCc8mY5HdcAT3NOldcV
dvD2ZKx+csriHGjVTAtt26y7RcMx3iZFbqcBpZWY/HSPi2lmXg612bhY12L5t8COINeVtTFfjUsL
t8d9szXJkDuiCi0vLCsRwrp/ZjssyIZ/dkLg4Bj/FKxnImFgWQSaD8gSyIi3WgrslRZGWC2NMAdg
ow1iNml49ItWXpDVcFaEfxdq7dTdtv3UccphM9rqL9XJ1Gz5ZLCWpbJBk12TVzDTOkMD3aPGGCtW
360vN3y7SKMgEU+G5QFwlkPDVpE14yk8it9llUtHeXAkDhv00BpzwcOEaA2Jx0UNqM9KMRYKLoDj
nC3XwsenmBQE/jwUd+nngk4vkz9Whc2qO5EstGIvA7KJcpjfjQguhu/mKiBpAlE4sr0bzN4twyqD
JBQ6QEHxfW8aoJ/erOwbdyh+aVukVdMnzUe6grQv2OAEHwd2crPjroEoaE0q07VAAfupEs7vFQgY
M+CXqPsw6vx/ZYYAyA0vUsiuNECTLXY7Ubu8Ihap4Cybk7JFa3y7qJ9q9A1ZFCg4QAlZVE0hHmnw
zJV17JLy8mvks+A+BOpgna3J7HqVlkfDYcKSHBVnrXkDXk9qd7dA8NzONsCi1bnKIevkVlVZP/Yq
4uGEjt2zER1XASub8dLVke27qEyWdtRXFlhYQSgavj4MuFBakd54nZB2mIccaFNGCoxpc4uSaDY5
x60AhvOu4iKFwBiOGtyzufB3SIdWeyxU9knBhsEkFvx4hWYwM1ccRqXzNwE2eyt1HC9HNUceGPjt
AU2jWKtTfbr07/IEAoHXQaoEGyLNBlzxHa3cjtq8NoLEpfz1yVDgo1BMRK+3SBlGrxiAkIjz8IAX
RbP2NVqlaZzfa2pMg3ZB7TPTDb90xJUmsn94u+4/8xJCmWCpDzSdS2uTdK9VyUmDcfPP+hH084H2
+oF5Dszl+1TK4sHl0P1YBUJKbe9lH5lDlLp0vRfVFaB1fIKQ+LcYAgb4EPtzGssgX44AQRLJJNoY
BX6//FuNl2zUDlOiMf2JHTv7r3ivnHD4mzKVzIWnnRJzE0zX5uiqNKWzZaullnPPzFAu1BqrqIk8
GLRS0vG4UZo6833e6pL3FUvp4uVB2/iGG5tD48g+XMy21jTsW9Xn4/GJyeTAn0qpkLNQVpoIwvVN
tf07nJiRqwHZeLT1bAyicUXxjoQBM09L+4Rdb1Wc7SQYrU1szJbxhshaqke1WgdqePUWSdEkHF7G
qlQl2DEQ7TJKT+KuLdMk4IqzdfwOh4hBHoQ1k9O5KyVQIFZpyuvusgyf/gi5oIA+vZ9UnnxF/V8K
qTFHdgqv+PyPmYJTwj1zvfbn0S3yZekJh2i04D4L+VISOggxTuG3NXd3GK8ijncRJnylxNdzm+nL
y+2OilFEmQoLiZYDTBiWqCjqDlRO5mS76yRJmUKaRz/Wr/n09sOwlYBaWNnFuH1anBg91RentqAv
gcCQUnY4SRoTX7BLPrbJOQEI3kRVKXs0iLRoXBzkig6WDKm3Uv4wMjTawWTkSWDOu6tarV5Sr0D6
DSYUdpsoD3N28D3+9F7MFvOVJuyxfOmiVVYakqits1cazAwbN8Tm9+1fKr2WQXJgkB/HdkgX97hp
dffJMEDD64YD2kWfVuRgztt9B9TQ2Yh4ixiKme0kwkpKRZjFxhjA1EKlO/un1Yyqs5lOguWOLZtC
MqMFN7AHFNAwzY7sk2bHkAM3oDv889zl4AN0FJMwLmewevEy23NMUW0KtevW9LdUsw9cRmCxjMI2
9nON578l+SYMgKkf5RtxZSbz/uzhXJANXqcpPLUfqiCe7vWKnld/crgyJDY5ouRahHn6uT+GaEt1
vMaAmsC4yNmArIZRrn/eGNfb41keB7P/P21sPnV0dC67KlHI2h2aEavzEEYsZg38No66rV9ZMhkW
3K+TsRe7FLES8XR2ik88x3zXwoHFITTYnSp3b9d036Zp2mKQ4uTwyA3ovB0vhzGuCjhGiTdCRNeG
qy1FqXNhfflD6PuInyTFetrjqVbbTk3wAlop4TcNeLXzECBIwGZrtBN3ZmOzCL13EvGYsOTrppN0
8Xt3KpBHzUanan471BS5LAH3c/GeZS8s09n6Re/FW5WH13Z/V7wEcRSifqRcf8yi8qVo+amVR6qu
6NW7fEpD5c/7hUmsCQ9a6D7d32D4uLofxMfL9i/sk8r8OLIYxsdc9P+CJt/97Qn/z8C3OUZ0HmHK
Z7K+VXr/Id6LuBjwKkECP2yQRAcgvc7lYGiiV7k2uC7/koUGcdnUsAkOkc8VZBvUbDJDEXHR+2bw
95mrhhQogmDxS2kLu8953PG0oArjPZ35/+FYtAjz7BffAtnaM8ZTz+Tk4OCz2d00PKTRkK24mRfZ
tPET/cv3QB1Yr8r//0lZFcWqjwgWjQXMbx+vXWTg4UpNO3tov0sAPnsXOBQ7Ix3Dpq+BohMwomlb
t8vhOKD7VSdPoVelPwakKVpUIqkZY8yB8QCSAZ91sQhK+jbXiUce6T5yDENO3AVSMeCzgqsPvJmn
BRAc/udob12S1s0QPD3jqTaWvip3KmBYWhmVh9R2A29+qu93uRjVttDBaPRaCM+dND4Q1qXw35Y+
IaZHycoGagh7q2zol4Tp7/KCufiMNZuEYQveVTnVpB2snmX9W0dc2YqQf3+o0yUZ6gZMBwtso3/V
i2hNxhSkyb9LM8+KJ5u+BkkmLLwZNhx2A0m8QSIhIMSgsGu2BJ1neaIVo/yMAmkF+uTH2krYY1fB
kBNvzqvNtgpD+VIeSiJBthVGKmEBY33yD8PtCKPfP3pXOnDz+DcAN6zvri/PpxSDwsrc5g/hb8lY
eLloG+Z6m41uPI4h4BQ4oI9yYudAgDsSz8+bTh5oIObEnIDQhSLWw5TzlrstGSS7gkrA7py05dQS
xk9Cu8gbVdGaC/dDf8rXqAoWehV+EiDtRfNTBw2Ra4O9JC75K8mKg3E3qqmmMZ15eIirUtep5K8Q
OQ45Xe8Q3FmuX6EgWOBCW+uBbJEl32f7p4xa3jueizs4D+GjX1JbPlyn2na5Sy5IK5PxwHvfG/ZL
UVTDZFsHcAbsSR1EPEKwU6SE2wYbyqPygrXNXFBunpeYyX6LBND4QQjR1uGA6BGcg6BZ7LJdCtfG
SkH89uugCn/Yet+MYEg5CuA8iAzjZUDEdqMzJ1ukyXQPvlKyzRLUXjdZNuVmdpQpK8Nc2m+wWBJH
pVEjOa1RZPqnVP/lP5zMEpv5L3vjjbNH1a2LVTmExRCOCBkp01ZGn3IcTYpR1VUqLfAlaeXVe3UF
83+ihGdHfnIbHZh10iITd1J3tY1Gk6rezRZEEQ6T9kxN49iRBaeXVUldk9C/57WbCknrhNUr5jO9
1wL4OQXaMCDxemSOipDohUF25prrGZU3mLcoq/cyL8rcmDDU0WqvR/RniyGPDrk+5Ahmnfzdke+R
DRoRqD2SFIc5+nFKT6lsLvokPfm+b7kPTjsEcH2Qn7i7aeB2PYV2Vq2bZvc+g9zYFvoJx5fS//NH
V03TjiEUqGCPZJxLiCMSVclOm7cVxR/W6eR4x0s+0lrn1H4kBtvxau4bHjsXTxj7YaPxuyzfIIMF
H1wrk4dJUt6TdNygKqUZEjaNVEl1OaYHFLPHpJYkt7NcEaMcBT4UxYDCKLDl6WBLy3aeX9fIK94j
MbOhxVupkPCpCdbeZrPaol5L2RYNl0WgB4hsxh4AstAKre9s0+k6ZwDWT9tLX5exNveAGTdedxKx
H5pS8Yj6QNlgHDRfgKIgyP1xA7OoOzm3/fbgTnm/Hwwgu3XRc/BendEM5b6uJSFIFRn17M0ET5BB
Wodcse9R/5gU4PumnPKmpKHx0pBq8S5KfEOrsM4GXkxhot+YcoSJcbplccuReaLZ7M96vrb1+q2f
bqyrUDIMeI93hj4aDXJ8bMmeeoe+HRa/FihpIx6nFlFRkJ3d+sAA4+/o1eKz0uHRHThGvvvJvTXi
ZzIryEH/uM5kUv1vVXudyd62bMhHYOV86IKCaavo2yav8yYXhrIGchd8Gk4VqRpWff+01cp8dhqH
+vq1vs0PlxHZ75m0ReFE4Clp7qdi8uGnYcG4DhyPW9MGx5TKhuD+pBC0LWMbSv0LI7FHfRJkol2b
uVREYlXBWt7BIE3dWV6/9ss9O3D73NgzWVAtsuSsi+ml1P8KUshVxryGiC0brHKde9x6ij5OU8ex
GvJEgD7irEmMHwBrEDJXPcb4feTXgUENlH2NYfaLo17ui8kZr7iS2Wod4+16dKapP1V+aOfiBBXC
IaZOKw2DbKpvKYCOV0H+fIHYEQ7HRjWKTGJXOvwnf0bquALUhnZmTrnhgx05KWfEyRPWziIYGH45
C/OQtLP9dxupFTvzRFnAqyPAFubmKKP0c8xBAJu1pcdmINrsG/AmzuvW2vYqT0d7avSOkNDfJN+5
wFUHTJLGADkMXXktj5ZMShBJ1+sGU9Cf9MTbTAKjw0hX9iaEqpa9mu2k2xJDU8krzZAnrTxazz17
mTUNnPf2bCzfJpUfZCtPWacMmaN9UiYHo6550T7pW/O2p5Xqbw5lQo6taaucSCE1iepvj5HZChcj
KMBgEoPnCODOoQLaDCCAspchpyOqRfSieGbzzJNWqJpi9tLE6mM+IwxdDBHEi3stKw9q0V6F5vNk
vNVEmNEoh7eZb1Kau5H2i832CgZiaxFJGGvfWgIHQWwArnSbmct82Uq21y8Hw6C7qP7aw92P6rIX
btvEY9xP4PQa82CuLvPPqB41uoUjrs/yRza3mf6xknkB5nu08MN0GadTA4QKLmQ/hqTQxkqErJvc
nrvBnledLknEGvJpfWtXx/Meh79UcxrpirDCNOI+04N2//aQhESMZj3GZpI2kf1mfqOt+HPn4k0n
IJQypiMpYwxhLFGjLfrssh+1yFUFy2iqXMwz3zUMMjmXRdQneX8Ksgg0fxlLJcRx0MaYXJpkZjte
MIxuzsbV6xqonoPhPnE7OvIaA4SaFo8/++YEAAjywJR0eQcuXssbzZgfy53enVsL60VR724y0bVo
+UZGlpspV70qGdBisMy90yhKWFEA8jh6u9UlBIbeMX1DwkZaWkWZ5qfLlLDeVzsBMEQhsEVuQqRa
tgZXFIvjqnI6cA3JpFwfPHy3ecwdEugCEoF/4L3E0DhmzhyUZYwPBiAWVYpB4S9XkxqWyaCM+bUJ
EgpBiwMNgwXOu7Lzaip7np4mL/tYiUgraaQtdwGV3FIZ9OsLLimIAVMQG9uD8Lgzf0szQ5nMfExS
nH14RtD/zBH19eltdNsuz3DT7rQcwV2xYVz8Frbcch3gzrXslSgoItCGRgYbKhs8F5AOPcbUhaMb
N9WsqMnGrLMoQsqEeJPH2lIYioRC0+gB+jsTTuKUAW+9JaS8pIhkJEKjrfgzx5AsO7VDe0p7Z+nJ
Vd3365+cM7HgWv7bMeqLftraqt+W6ooiOh3KPhZmx126/q0f3CeQdv5xBRcrduXhh+v/CmT1vLBV
FWA+edI9YjcaaT1vvNYZj5+U71sAk3JQjhuzHLrv4R2tchHljA4HQozsmImfo2PA9zjQC2T7owfp
MVny5g4BwkPR4wF3MZa6Kx4VkK8yoVZpl4om1hOX49UcF4BjdiadDnL0Kf9jr261kkd3bbaZy4I6
GlYjJalmMe7yWN03XrANIO408N+gx550ijxABhKUeL9S14H8522oEB/LhCNJ36p2sq4c6nqGK15a
B0nPIiXkoRyFIZkMy4qUwyyRF80rbrptxdRrNXn376OhJNVZF7MdK/U3dJ+v/pIcV1wqI3hm4fjT
AkIqFeQL/dw2AaIWpTdHtEMtI5+QUzJ+A7Vgp4KoNuDAeWXW2Z02KfCvtcb1iG+moZUOUCG/s8cM
SMsqFUv6CVmodwkvhswA3XF4hUTqKzKdpXWaSY1rbh1g/1ROnaJG7L3E20YGPzA/HSE4nFrxq0tS
DzzknQ/jUc67cVd1YDXfpTcb48Jj2HUpI3RL8F9dVDkyPIQucpnKuGvf7bivIxADhskAHeObucoq
9h/Kn8gzjX7CRMryD+EjHo29lQa7i8QWtV3c+3SvqHmJc8Em6E7AVMUbcRlOPC+VukDNN4VSBojb
pc7UuTRHIZieMrX82OmVrFbVEb/ByzVys3e9WtNEu0bFZWt9KLUuknUnswrhEO5QNSkR5Z3PypM2
O9F0tQm8LtSyLTSBKB6TkNJABlNOh7RuUE2F0KmZwEVaudj4vk/ychqqQxBXiRZSJrQ1ZvpK7Pfb
2StrCAeEfDgQVjFiJ7HqD/gJqxPkMx5Ci4Ov/QoLKaYmHow5llQNgsm5COvIEsZC/2VOB/2yMePs
Jn7EtmPTTleJgVPgpnoX2JTYsrOeu51qUzi8/FysXATnQuGywt8shnGItr9ezDBJhhMwsBKkCDKL
rBUm3zUodKyBKRtGMAwEukVDL6T7aTzwzODyv5+C7w+bO6puaGqU17vsEmpPHfzIelegyuH1z3Ji
EUFnJ3REcPeCqzJoj9bJuB/lht+DjmAZHQXZI3zr5DpLF+bqnroR12/5BY9JfU3zNyRRbczCA/Yn
C9AfaSXcfXjR/fUFQyB6LHSIK5y9uzmNVbFsHfA0s18GrXbCYi5xezGeDNBe4kbxE+pBpA0h+3XN
0rqtcraAXMI3yD9R6H1oiyt5NvPoKmCYpWQAzJOZqWojjRzyvgGf9tl06+PRMxqc0sjr3nDrXvvP
mVLSI4LxMX3vnWfuyL7YkyEoxCUOmx8rwqIGae05CWTgtxurK23TpFG6ZvkaNyE3WBZkZ0mP1fgW
hGqcaEOyULVa1D+nxQUSSh9+ecdc41QcMy3VS8BktlU2DcGY9cUfkqAtxy7tpYKSIoucHcfzgjw2
f0fiDoQedLunN8mjIOBsZXS6nXkGgieuuHogHVzUfXRZ73y/HjfaOmtUQVkYOfd05JKWzQa5XdnE
0dkRn1RyuPy3gqqBGl1Bu+7ENFMUVZ7VNs5wBT3IQ07mco8jCtR1yDC0frFiTYtCHv7RH3MSUkhp
QZpTk161PbSK+gwSsYKHXoDQMibk4RasfOaT1fLEFausQFugMfcZWyzWOK1788hfi5ieNsJIM6hW
LPWjkhIwAXLeOTSGXK1xtukKa3N8bFKLhHKEb+xi9yke81HflY3cZ6MRuUha5FcUPH422UXm1pOs
Dd6iGNBDtB1Kl01PjyaytoyiZHRftPXMFdwQ9ZKQxHwoBrWCc7fHcfvsw51T/voZpn1CXUnMDs/f
f/CEKmiX/Gfv03vSBaPNvqYIN2leLJse3DmbjiCW7DdM1Tnrn7gPkdQNI/eKxZUOEQl9mUmF3sKg
grYJrQdDMRQjwYzatcwLbtQdEuLHw4EGwYM590a2rNkA1ccLYxlh8zEgrBMgcPkspbNzX8bxQg2A
PsFKbHZbQwNqxb1I/3zLXSB4Rom1qlstP6w7LOR7RqGTAg6XcAXz0VjVSp7u3+pFuif4HvZR3QkC
UFjlEn9az41qy1+YP+UCV/VsQ9YXWuaTOm8Yb//LZC/ApNOT99c1btz5iWSr4bIyxPN2Qych9D4G
55R+ykburUb1gAFTu+obBJhnfKlyXAaUyHLkVxmSWoCs6p0d/kbn2a1wBaqsDzm1fXqptJwVHuVY
DOEE47bkYZ+4BFISLatDGYWgZ7CAcBCxkFYy3e2Ed4H/W6KDN74fozNSiAxiFzj4zm+TXGcmy6vM
FL6pwhtznI0sHJ6aB8+ymtorJO74C0Pq2l1wYefA880kfqaxRJ1Nfam+5tUDqZRtd5HePEaPkUvK
Vuw7kb4o1Nh9IvCZF7VXB/igTJ/W/fyBQl07sfgfVa7WBDq255J43HlsBEDRHZaUJA5pvGEhkOSj
FXZ2lFzugz0VI10LcDNLreFspazsDtPLHwxXdcp0n/A98twCx1O9U6lXKS8reBRkhq+GJ8+CYrMo
WZQGwKhjmKF9wjffX3yoH4yhwUHQk8laPAmq4rr/Dq7jp9th8IKRIJJhnuih5sORWd7c628ONypV
a17KNU23UN+oszuLR2JnMRC5pWjH295MW8r74t07180iPDhFPl+w49bIYHGVfi9Ke84UWjkZA4Rk
nufMa9dkZCPmfyw45GnhLI/0/4b8lcKydpqEJvDssQdZeC1wKhBS6n9Qu8EdiNqjAf5EcG7Kqm3Q
rD6B2d3xNkihKmPiCd1sj0UjkzVdh7RASIWhslkkq1sATN9ZBxlSOKfeYpF0+JcusdpGkVtwl3Mi
W7KYiEcQT2G/vbLEN8hUeKKP4gh/eTaGYL8O5WS0TARqY9NlZKd4afBcL3s5hMo74vSYsvqMi9Hp
Gc6jAX30Gd2AE8uuM1D9jAEcHdjmDL5Ybq3ZNWTtwmDUEsVG5oTYEfguZ6O0UHiuMXphnZVPH/1s
1ETiSZP2vwE1nORwleuzDX9gqWV6t6cq6xaeU4bawx9o6mNl1JPhztW7HFHy/igfHjB7hKvhk607
H4H/6rgu9hN66ZT0BtPRt5bXs9SNSO6v90leXYxRQ39/1zlPeWa7oeR1YKhffGVC7hl36lxBzju0
mPutC9sd5WHkjrYzzBdlXaU9qgrUe/XUgnJLJnWdwXGRBRcAcS8qJDnPFLtZ6xs6Jc3vnxX6pgM+
7vJJ2VAyMDse7MU7U/ZAb2Ty5NoR/G0vknhlXjxUx5nlbXX6jRWsaaVhybrSdMWCglPvR905NKNZ
2+gNbKMbFPb/iEnrmBRglDd8D5RdYk2wBk2z2tpTnlGxdD+XGVnwbQCTPfakNySfv2bxzbC2zWi7
94qRm3vGtT94fHekrydP57jNQOA+4eNOk5/6qvushwRJxSvm1tDX6GpBlwc5ESae6TyCshpAsJVo
HaUhg0QRezf58ICOsH+HvmE7huYKn1vQ1aTWbUtrpPyE4SNWeb4sV0yboS9FDM4OVZb9qs7Np7R5
iKMdbZsdjCYOzy+dT4GhpHlTQ4rG/l7eWw7Cu9MKnDQbMxmay9wXVNqB3XaaeLIy8xCKLyU6u9Jw
HGvTvjucYALtLGDu8c/JeOLJoeXLsvlA0DvQ83YIb4go2eFlf2PaAjTHPstZbng7dzzSXUkUrTwj
Xe/ATWQE1nNEldHhJB2PDU8qRiWQXRLqTjk1kuBZRevnPHOuIJdnk4oglBiGbI6hG2Bi54VK01E2
NX8N+yKTE0HPMKaFrwkXUfLAEZaMeNCgHNSEXOtsr/ZULFeNEI4lAv/PUDSO4qhfk84LD7NZxNWN
/2Swl5t6xecMAiaRUXQZhLawCjlTmyEcznNYjNVmRygqAWvC7lPXCVDmT7LbtRDDRT5eyG1Oj8pW
QnmKdgd50G87GW/3J8OEzNaW15oNRnIDfvoxrc+yGdHuuxzOd/jkNZ+vV+u9GuGrKXSbOYmL+EYU
9zUlPfX3jtm/7Q6MRtiK8IMfARbTqgXMVvoNH7R2xNoPIL+GrcwEtKkuTlqrUAWe0IrNbxyGmtDG
g1SJ1jZoCYbH5seWZ+ZOzDzDhNdowVaa5LkvK3Cf3dLtYiVOplYUDL/QTbN3grNIbU1tqi30paQK
F4xhan2q29ScsucQIqveP2Itj0/SL5O9cWw6z5Meotwp0n8e62KDlAsJ1/cUw/Cmro29sJNi8Iez
wUefqYeqUwhtwwhQxwEIZTRB13OoyfVe5JC5NfNRqavG/TjLBsbTpL1swA5oK9Dn2VfG7NxrAJsa
Gfr/xmhwjmL/4cbvFfwyb9rtQHBeCOGl/oNepRRfMYgkFankS2RXMZbgCWNd3uucIRGfnkZa3H+z
IqSTFbNV8hIMGU0c7hKyYNFVZ8Mcn3/GH6KYk1vBrjiBz4bo5A85oZHzvxQwVUFCAMYL5OPb2Gtx
gaAb61F1AsmWUz7VXqFFTFeXt7cvFKK627TjCY7nCb1QEWKxWWJohDOAE19z8czLox4+5DjCHn1a
g6mOGVukBkkTTa9iO4B2+uzll2jIbFEdmKLv9yrthZ0vFLXuFGJxgfAiytKkDbW1E3uUS7FOidOk
3FJdL1cQ6KO0gX7u+TL3iHFKWk8GlC4EcgMuYuncq946HU65B88zpYw4+v7Zx/sF+bbZk2hFpC45
RHUINbu/SP9jlAXScYepNUwCZC1I+6BMjXdAB5cvjCrZjC+NN9OOHelMoD3qqcdLK9XsPvh7kYFZ
jQ/E1ACzJb9Mhbq5/PPc+hLBlLyTDxL304CZCGJBoI5ngP+ab0FiZpxDpWF0jMThFa+a6epw/zp2
SiPX9bOQICl1j93IvCcdoIRXi9UjzRrfs5VjkEszJss/pH9+jmL3MYNt+rU9F7fjLRVi4BDaeYbw
hUj8jamNtxSGDhC9Q+VW49FS9p/ceCGn3L2nqekCadp2x9e3mqtbaOCwhjJjt2XYtul59cOKz96m
WN5Ar3hEGSIITh7lfAnVXx22weLAzHsnR3+cPr08ZYBvlF2vmym8tPRSlv9kQqtQzClzaZUflLrW
JLjV3NE1bBzbb4L2Px6uDPR2no3Azjs9VRQaPrg/TWJKlkJVEkb7//btMIS8V9nokJmzM2RYMLN1
4LEnnumC0qPnx31AR5c2mJTe5jyMguxT49rCJcAt1ZGXyYBXJ2xh/lN0A7Wj4CHlLvsz0pM1q21p
FIOU0JHxRD4mTcu5WDW5RDfUd88L+SeP5Ggp3aYjTD+x0tMlo/rqNdnT64SWgcA3KDN+FvQhsVoN
y7MukQIayFxN4BSysa6ljdglqiQJjg5dZpou5KFlwjDe/12pwFH37UBl0J3bzCTZEF0sM7hHHbRK
tO7ry2+4Zd7e5c9Ego+taOPwdHUeSSe/WCn71UQWtTE1zvoFcrqIRrNYIXdg3sBEFKLgnjnTEdSg
avkFHApjRZzZLayhSIhhzdX3UsVKxtoPBbZHoL6oxzBNW9HufMOK5jMvzzUc4g1KwIEpJauHhc6x
Rerd3kbPaSj92YEEMeB8OsH4DVwAUBMvT5yrc01SEN1BlUq75HHqGf/dEli3y2O833L+IcfqJgjw
T/OEXxeXz0R/8/z4MZHSHtJZG7Iu0jxw/7QD8+Fz7fFyQWOm7ka21hac8FC+1ywOIama4S6Btz2Q
JPiVMZjdE3xfkAhBFb1EK8yMWFFi++b7YS97kd7X/W345NK6KOXlHAXGh/Zn/umXlyZcM4NwFFGg
hRlNnPPB5i+R6kyeWEuw2icyFttcijfqh3wenXgHXrLtG2HYTOOkmXR8wSgV2mmPaM5UcqJPljDe
SM7K2a8GCRmiFb7G21E8iwSsQzBH03p8aLM7C7bPGguRgq6fe5Pny2FNHixMt2pXhiJJD1XYu/7u
6LaMqJnQaIkB7ygkceqa4Xn272mCBV4G6a3jEh0QIyb1Foee1R43eTG6GHz9/zm+lVGCM24BjqY6
/59H7wLjs0yzxDQAWCzheGI2gz+51I9Fn+AbqzkKWjRwaRlS7dXcHh+ZWCXciz1LTqkkOfwGGBw1
78xUMOZMIAjc2guVshB2QJm49pUCYLv0ycMn/Eb98yPgQnDqCgKhOlOs/o0N8yMH8Ai4HeHS5T8u
iE4+6Q/PRU6TTz2M255Zxg+v7EbHmwt6Zva8+Ji+4cbnFhmvo62OJEIqBCteSzRVHsRy0B8ZiJxw
hzUpf9Bh+IzGcnrGdfB91C7eK7jxfyZoh3lMZ06KYWlyg/MNs0Spi4a3O0/rfDheBqzZEN/dUZQg
fi9la085+8qJETIOzaNZzBWddT/eP86oOsXOrzFsTarsJ9rNCMQBPv3RNrjD2MhIMdB0cYtBhwTF
lZzbKfKQ17yJBsAcrdjWjJhA3/Ju44EFBJj2dQGckH3kbD/y0YgDp+xpw9juXsC5G6G15rUotelh
E0FT7VYxtrhb0fzGgzKu+xpwiMUD/EoplpPmu46H3q8M5CR0Bs8TKjHclNDkkFpNstR1nttuiwv9
P1O6r1sUbnBuXEQp2aU98J0xJlHB6Wp2vGu4l9rNEWRu5+3CjOVuKvx7sYp8z/uOIapKKfKRbR9Z
EywKJZ1NASkoTRGUqCx8Agyvr6E7QmnGb+6W8kbeVk5LpUadaZgVTYmxvkCOJDIpyyhvz/8j7EQQ
G1OEAgEeU4c0nLJhMm59X1f5wrmbDHsyBYsgcaVLgd0NPcIalC1+ZJxvJzpX+C8k452LPgtZ0p2m
YpGiAe0+oC82vFEpiRiQKadDlAL3KyRfWvumrZ6Lp/QQB2RmYgRo9UKvKLydTYzS/Voowgc3Fot+
ZHe+iQZ+gkqqZzNVdU02ADgxZ6FJS8Gui6QTlOGxrje8EzVkjGRDyGEUv+5/SVgZYZOEmH8gP9V/
Dfogye2Nya5D8T2IPZDHjcXd2OqWM/g7qCUf834VioHaPrEc30yhOiWf8TDALxDlxbR4HYBrQG1k
ZaGydW0xYRxV69CzGskXRtqSd89T0YQRJh+241AmjSQhVLNW500rn+FeNkJntLIjQBgClM3I1kS9
CZSW5jwYpPJPmgVQUk/rZFZVBzTaaHyd+S42bCKLfLAd2fJU0yKr3+oG3HM1W4d2tQ0LShABctjX
dymD5S5AOGvBto4NkidL6d//jiZphT4Ke7x6JuupkFl4qm/3olg9MUBiq3ODeXCFVFzy3uP0fUK5
cGRGi/haSQGa10GR06AUN2NbPXkvBuaAJZI415ATmfZmQea3T4RPxqqNdmMe36JUrlOZsUtOjzdS
hCcYxzXCLsokgHZfGrK8N+WckCA+rr2VkhsUFsBgJgWQrb89fQ5v2lwnsyVnEsx4skwjdaUqPyPM
xH7gOGk+9g24MYhQvK7CiCMV2PpzWSARcyhcJkcsy7kyRvEF+Mw/R560T2Wu19Tj6rK70nITtFmx
BE2/RWn+SGgsXV/bF8nf4X1PywLgpXQru5Qp6cS5eG1zthh/v+g1t2HlnATAuaRjEHWz/hqtMKMw
m0h88nVS07JqIkg1nlYGsNca5O+rrv/XTWvuFdjOa0RJ5xYOawqLrONxRUcwB8hGE4FnrSkvPtSi
DAe4XoR1NwlDNKYw9yo6dreC0Oo63RfY2aFPyAjG3YFD76CfSFqrd4oz17Q96HmHqM7nkbxaDa03
Gc4r+lfbohKp1Km+mBfzD1wiEdz4FsfW3HbBQZ5Bs2ZRAJEYWxN/w9IN3iwW3/ZwK3XXffyKRGkF
JaKzsBVTg7qKsWcpua2KjvvigKHLp5qYPGYxuTzk+ASGi50lhI4Vxm/zEwqoFCNFuoh7FL9ffBzz
Uj/yHf1zeENqcUl8+O7wncQ1gm5GBG0uY3RDOrW9KUDYjxtC0teTnJIXF59FPoQkw5bFQoXi0E1e
Q+RfIykQ/2sw+4XfTYxMTfLa6a0kfKeB7AQNpXw2PXzxtGU2jGxp0xj0RTLcFj07b7Z2okmxi7+Y
Fn6+lxsDCPD1tXiBzmcRyaWYF781Q6uyc0vvS7lYoEJ/4en0dlkrKIvy+5ht9qJphmpR+MvBHzaD
5HlLN/M9zKSFGUsfPHpBfvg9sLVRy9ZaeTDz9/bt2M8CWhAS90TeSM5zfp2E9jyFEVZf9RnCuLGl
aLOVyCDanFzNeJNhj9Xq7c3JE9LJCgSwHzuz5nI9IdCEZv/eHywGt03MR4ipRX4G0R3ZVOwVB0u5
P8pkjcrIFzrFW+DWJnltQMupLlGrS5WUkF0tSnU4xy0VGE9eO9PcOBZQQHWkYIzXQKAQ6UKygcA/
aDaX7ufxi4onDsgiExRFkwBT5l+NAIltfayHlnkHJZr7t7jwmMTwvrRvR85WKn1p+g3arPEQ/Zl3
d6RevzP2cnX1ftyJ8uwBmoMRSI2s14kd8ErOen3gCTooyNiplyYU/zWC4sXhHVj0bDKyyerpbfwB
febdWMS2J4pymcvdRfAEmyTQuf9ef2qPYRRf2jk+so4380VCJgeFZ7Pb4JdKf1MW99itTnvRcMkY
CaUjIzyLEacmQChG26dUFMzjN/CD2rt8XHqPCInjrlWES4v+qlhewq93Dln72Xkz/gGI4nC4OwCW
DQ6m4zIsm6ePAksP+bXrVRZs721nJwmhkQxsdOXzaecXOCmNajmrmbyma/qOPUtntAxaNny5C3J2
U0UqIATfmDgKk17Ni+4psBRxI4Hl6VWs7bgY/uZP0lir2DRoTSjE3+Z1DrN9S+ePANE/vY2V+P4z
S0NHEW3MMWJt23dMZurG+pcsHplz6bTHLhhzHobMx1WYhGVqoKh6NFi6zkdWmK9I19oFU1+Ri2k0
OqEeVWUJNDL5M3fZGDg6Ljf9+nfBSg4gn4i6VfS03Tcmp3bNn0muXGxjrgOamT84xymc/Iknomp5
A4Fq3I1WjZPyCGSxstxMupXbBedzTZnNMgqSehVTanHag9HwjSH5QjT7ZvCfQpa7jOwqYV+r59T/
eMAKrX69nfjGDdJmIE/dZRRgh19vIiT9jYONmM2SSO6LRB1HXx25QbNQQcQko2bN9I0mX9sbzbyM
C++jvmV4y8nAsNOpwhSFHgs9nrGHQVaLBeJfyBh7UzSCjQQhCxNhd9u9otGARN+SacKlkJp4X4iA
NmAnQ7G2VPTWLgvrIFHi+UMwjQsmoTxwr3CDuQO149+SpgRhm7t3WMvUmbnLT2FXRY6+665H9XNa
Yh1Ca/bgaOUFkCAyQb3GRvEVuZjCJz4z7CBorKEGlePUOiG5wFDIT58YBRx+Lr2xcps4JQfWBAJq
g7olG7CK7OrPsZ3NNSfmqjEDtUhawuBqu3/doPjv6ZDLp7jPyvM96OLqJRqXNtRNYc3akt5p7UYJ
cpLjxNeP0XcgIeIlG5LcEkhFBL6K0s0E0ygtSPcabuJ6veQvVpwvP+2CuYgFjxhHYH391BVjnUtM
+czOEyBGlIz9md2ny1jXvSXs831R6GSviEg63PP+AxjydES6rfWgpBm+5ZkzwkypUl6cBPhlK4np
z8ZkkXthJlmjIyUsslVdZqTbq6nWDjthUKza3cCOnIbyNfM4f9qYvh7HS+KhDr+NZ4UGDHvcuqmU
5wWtUwUtlufX/yZpRL387JQ9AVaW4Eq56nIPx95el5pGT/mnMJ+QW26Xt9bpRPyq7EI8Xl/ktkyl
xbQiUQ7m/kqSVASdYK0Waz7bboa1WYiVXNRt2/Iq/ZhKvv4WP0yBKRGfCrK02955pQqriGn0YL6X
ApaFEBkVu3AwU3MtVfvkTUeYlCdawBaNiJDoxSxgNZ3ep1x/VyFbx6cNu1WsEz3BaMv8a3pU8Xl+
/gzViDyuN2iumZoubBp9JT7GmXUfyNJR6SYJ+gtyB6RvLNHJudGXtsOyPbXyEC0WdlzSvaVdK3Km
ndmFfEAT9xISTTEsSZ7AmNtOsZLyY7N4Qiwxepx9wsMK2jbIBifhqJDJhTbngTrgKjfuKMAsEuR1
asLZm4SoVh27/UGW51ykQDq4oL6xPA8Fg/kvIxi2VP+IDv+mZBypo/W04km4xxwG2QNgrulsWJ1S
vmV+R2ESJ0i84NM7OPdMv86v6AyWNRqzr8XpYssieIf17S/ITKgBSA5nJoextnpYSSt1ki42meyh
U9UNQZi9cr2ESLHMeFuCjr0LkW8Xqtt+48ca9oMVVSImHzmrxjkjQdGQgfWScVeCEd97bVYBvdsV
3xVEXB3Ml4/m/3ttInSYhrnB2kROXINM38daonTcFmAfL3Wv1345shZqhGcgFprJk5YKGSacrtjd
Ei7tBWhUpMiSA6c4dlAt3A+AnqUI6anDce4JN25ca3CFFUswUc8PRHs6dtzDaDycISibmXyl5qVV
9CYpDCxKxEt7sVdyRFjJVaAb6IMn7XaZ6GkvtjoE4uAcf8Xshl7LyzENThLJdan9GP2ny3iUTZ4t
Uu/bt6Tuu0Dvf0Q9omgBhvy1PD+rWuwmy6bK5MWlt0d870vyVZYifkjvJzmG7s9wt5Lw3+EElLXW
qWYrivFj4cttn4UlzBxieg51w0MTDnEKtHYp4w+CtMv+AMFXDf1WXFKXZolgRuJTxTagB3ov+Jqw
TVpmBG8HMrEY9EtNej8G0AScRY72HpYqSA6gRqFk/SgpJbCnfsSvOnS8vqvkznmttt6f2PSayB3G
ykWZd1ifJt69n/OMpustbhm5XS8xpEDBVsx4VwibGAtPkCxqw9nyuX8BSLNBFmzHePM+c75a2zTk
/6zcRlCyoeTiyu9opjTZWrxmHpg2pgMvjtK0VrGB94fxH7gE4er/N+vgMUyW5j7wXVdsjD8GLg7G
QqErZYQkHpGOtiCTselcOkx/j56Nvrzos4cyAIZnn2q41DFR1aj9EXgNtEG/U5ZpPKiR2NJlzge5
A043b4ltnmVeeoX8E2vzWgMszsfxXdRduWRsGfaHdnuU3wZE7otRMZjq2Ch7MUwuzU7tewA3dOKi
fRjKTqeie7fi/LQML3CDgGGnQE9tgoN3LdH1JBOG/6gKP8VDjqe/iVRcAhF52FPE9Qpu5MNAHY8z
fGJZADr1Cxkp0vq0rpVewO9314UcwES7avu99CUBSUX+oMzwXFbXKzm0HIh9MlKqQX6KBbHqUjXr
UDTdV+j6XbYzulga96D43l4rxefWssNcp9BwMkC6CrZ7FxhjBhqTYgtC1u+zvqR4Z6o0ZkVIBgSf
opEoYl4Fv5BLSlfBygPE2TUICGYaaau92UZSNW1KIKr8rm0xy5p/J1EfvXmW+xkzdvVc2Ysh0Jxj
AudWOAP3V/mrpVtiYJmkAKFyfHZSwZxWqiJUA0e2pkRaREaoeGRjP0GTAdhJIZl+t2sRjiq7ZZZp
goO3ptGjkXmOIcr7Xuafvac/tG4p2Vv/nnLz9EbkiZnuCHXXzjMnDlzvhahk4KF9ZGRn4D5kGuIL
b5YCXVNK82VXlAqrZZ0rhMnt0Z+4sNRVEAaLw+HBF5OV6fBUn/8VciqmVa6lqNTcFEgmmqitxiJJ
6K2fB+/eX6uySek8SxDGyzOG0DPd/AGZW0Av6Nr92WkcURKZLkpemFsPcI4I0Go5fFzoit3iwg3W
lcnTtmzOxKB7RGoU0By0AG0+VT1KhBiq6lwMyCOD77nta8M5CbQjJQq3FiRkwKTBxD3TF/6aPGfF
4RLUVbqKrcAZELLwpSe576ND7KNOQ83OoFT1BUgOaEDBzBjf38QGh5rDzvqKQsqurONvu31dodbQ
5whUmMcoiORUm1A1qecknzu2El40hcpS8y7pdWntEk7TOcidT9rJy4GPywI4vexJFTue30FEaPiD
WpvXeCgqsNNuixb+FbK6B47wwxoT2O5pAp20YMO2ZrS65kthfTDVP+1shXq45qfKmO8x1zVl1KCF
71AFz/cbCpP9UytzNg8QnWV8w/X/TuCWQlFFGmVLzNjxyPeEL6Fuv1wiP/pjJZryAeI3YcaATlIB
7pB/nDJ01eKTViBJ6p10erWETcTCG6F/NBZ9XNOKXCY0RdOt1AiIAbzktB15p5mlQf+q/AYJ1Fik
+IFXktz733d+EBEylS4uFwRdkHupsVabCHwj2TrwQyXowUxn2jP5tSLrSEQtK3rvcAwiobuoaVK8
3/45ndgI6oonghpx2p09XAEHWEG0KJRoaIga9cdbf/fCDvjXqtU2DS95iq6+c/5ykmxb3VSDQgVT
gmTEOLdXNmaZYw/xt317GIY/dAN4kKhujgYB53t3bNOpCI9Uay0XFehgAaF/mVIt3IjUVMl7NW7a
aGs900xmgmiOAwsdh07DwczaYuXU87R8oTWtVyM/uq2L/8Vq8yr8ftyhvNcogxDO3EXbIJLWSMb0
U4Eqg2PNVF0g/JGWBoTMYFPFmcMYaqDL81JiRnlNHoDptok5yLYAFgnUnU2QC0JNqzaafY7Fjizx
MI7FAs/NCSK1HLzLmrKcsTcjnUSdbcBlV4YaDS+W7ej1t87jfIt4cgC+L86L4o6IYh46EFk6lJf0
hOZzNwruSSbZqlxfTeoIvZmieym+jt2wO9YqbHn+Dy9stEEx67eDTOOaKHWM407/IHzbqsUsbbZm
nm4/N3tlmK1kGld0BeKGanPgrEbMmKYsxyyt8kAdkTZGLgMop9X1jVqugkj5jQXLDyGhumhbzYlQ
CKE1XZKNuwBGz8JqoFN9lqtP/HUvgxk4JBb3kS42zzgjGHlkbpGw9aQ7vbjQmr3shuQGKsadYHQ0
ICWFN3dIN92AHu/zFPsxVeZWiaCX4aSRw1A+z/iohdXTxTtalXqJEUu/m2lHqbCfDE4zGelwEMWi
J9cNw/z7xhhJS0PMSx+JsDWnGI87ywUtgHYZ/tvuiLoZa7VL1M4LrEMU50RfW5JOvk30UsIyfZuw
+PQZYCP0tmG6xDuNqlP8ECjBVvD1iORc/9cplUvG8wtJufuyfkSz/W9Gm3KfNC+gT5KYKzONABNO
bzFGz+kzcU+cSKUgJFXANTjiq/32SwCYpzaGqaQw5rXMuqT1Dr8dC1x1JDg2gpUTcYHqkyUsDCu2
Pvw5bOCN3NRoK2V03NxPNlXiB4AXfFWhnoxMDa+rChyO1P+bpWiKzLEee5/RVYrzQPd75/JKF7aa
RZbPyC60kdhUqNPeB3U9Giu06qjAmsoNb22T1qpYANXqr7hSKzVpe/1DIvQSnJIudhbGyq6xHtzj
WC+2y6Na+I0m1p+INPZ779y1s515/5ehYU+0n+CH2GY3xgzfpnmikp0XNqEjYmQY8tAp/7GHX/zh
mdE23JLpIjMHj7cG353P6/86PGlCXdZWx1vnKPpxXCnfCw+5PeQNi/Rrgdvo45lIeYz+GlLVu6i5
eNu1wKKZzwZoPEeqp8ZSy0HhUeoqhRR38v+37SO1aKVZITCKCej8IUWpZbE7x2gJxkDTT5OL9mrs
XQI+DnMrVvfgoZ/R6Gs18oXPsGAzPfdomcuJqFCGwmUPdiPsrdKss/uIkgQihyg8Ts9WwCPQz28W
D4zW66KbmCBnHsxXK3KwOFVTp7M27S2jlhh+Etd5L7yuT9Az45Bxy2fxNRdQaglKOozl3KaVO7ul
pZ9VfHwLaUwZjIz7hzoESD6pAANf0IIy6k1y/cFHjdcm1E15PHwrlsmsRvQTJc66jDAfDXZAJE7V
nRD9euTF0DIbe0LyAuvF3Oqpvk5wLJotFXV6YyNuQ28aWOOurop7uCh4EQCPcTsIt3eMbD1H/80O
LVXsuM3NH4hxijCjHF6mISY15F5LidOwjCJuJdyYYn4YaJjfhhdk9/eCwd1ffKrbrbXDXLQKyP/9
j2bewS90rZbNnTSooPyl2X5zNjp5pP1HmedBuwCwnNNhFRBOkW72j5tafVOu07FXWa/u7Uf9fZNP
hXXmvTqYC7zUkj6SPOmBPDb3/dbQvEROptQVgtBjDlSWXLo5NAHIaspkKHpo2sUWrsqR5yUCkaA+
0vkW8rg4ZKAqJJqqDi0z3HqR06yKN1zbGQ9iK8J0mCQVbf+k+nPvP5AHCDFd1LDExb6fq09+KZsJ
FXrS75bwQUWvCmLZUP09/jeCbBk3uuKEaylhTZiAhwjDLkFq58vtWLF9F+Q2eGw2ILLhAuIOQAGg
rzg9Q+B8d0qFNK69G+XFyY4mEBrXHS+Km+vv9toC4uGSG+KIkgvyaZTvSXUf65l26KSW1j6oQkH/
pBLL7eIZiZNlIbnYlGfEdr3HaXTvVK7HULd8spL7Mk2iroG7aaV3AH+LcPXJYFryEcZS2AlSRzCk
DFPhGp3aDleTHC7UumwzBJjuGyv4sFhoCbTKKGG2BWHObNPberGP85gNNmsEXWwZfMMsccg4fiJd
Cp9hVsFsMaSTEeEsfRaM0CxiRhnnmuImSYcJj/sIpF1dJLpk78+Hv0QuRHbBCvS+PlccsCag/Nhh
FVTetA3tuEdoYSm24t60jEdnHwUoPyuO/nPxqZuBgEF78+ciYemxivhr/m2co7tPwImaxRWLycbX
UmyM9G8kt2WcfTjcY78ULcuG3uWNq3oQoIWd3OUhHrBqz3CLR+uWp3H30+KUpD4JhfDMo3S5lSsA
mvRBFwjjcmUra5JNuH14ueqLK4kQstxM8ByXYYUo4jLb3bHDrzeu+VHRLoISNH3bOgHyNqHapUFc
Bp7IS3GJIuKWQ+aJte/PofVPXy+bx3momVTsyf4teIqbTJ26h52jQ2MBLDxfg/Hyj9LhT8Amr1Wt
7Yo5xAZJLpBQqYQMhoAtkCibu/i03R3+lyAzk7rXijs8EAUz9svsR87BSPqLTNwMEfhAyMW3JBqd
SybwW32lqd6OionLRwZa9RjOR+ZW9QZ/oXj4yoc0OBJCFGA9topruwgqEabcfvdAcbykYUjxODLN
y2CC4vorEsnSQADSciUg6TvyMWgXPfqZQFheo2PcCo0tJ2yXPTUlXsbKj0mEmeK882DtuZWW3P5m
i+MRnG1MmBKfJP7dUAaZEMcwAao/f6OCWQZt6uE4A0QdBCHTOSnM3BI+BfzlxvUe7ZcweBSqkZq3
CfS1ghUOw3VPvHClthstWevJfH7vI57EE5FaxEUXsLTc8sBcoeIb9ePKtBmNd+Km1ata8Q26L/Ga
1Ftr3cUDbOfm0gpdJ4zYNlYHi4ukrXkDt0TwMXhxW/Lm5k9kPfUKm0i++d697I5cKPzD2LSLcPzn
vxb4yqinzD7EeKuLWDn5lcgwan2IouFS08B3n3sC56DoEmmTGgKIkJRCvqCGzkdvaxsZnNaGf+sN
68U8Kic2AeaS0Of0Of4K1HSGr0mC88Ksjll/TCUbUFvP4z3oxNej8hNGOwJu+mNk2++XJNtJoseL
8zrVYygc/EvRWdOXyq2+R7hajLt4GpiBadIZ1EOvV2+FZ9oj1NjVP7+xaEbtWm4X3nhGFolZojZ7
AAzPKJ5g2ekSaH7cIZIQVThUWGJXAL8453R6w3L2NihWfBMfixTOggpZyHdlNxOK9L3B6dIPVU2p
zCYoi2Yay9ZDDxofNmItjxhsIn8vKu2rCJqI9MAuoqVQ7V1xxRtLWjf3cA3Qo6tePfu1xZSbHBYM
0OU9KAHZIXFZRkG6WDiT4HC5fLtXwRwBa1/rym72rtKkZ/8+hQUpb1BrXTOMASaJ08CA3cADReLD
3XUxU6dlfiSfzKyZdK4CFmApVd9T6gcuaZ3/CWTilIYAM/yLZWuI8/NI7aDcZH4V0HJ5DuwVoB6f
Sunah4dhdt4SKYgyy377Mu/aNzvhoXfcgnyLTO6BsJSpChWl8qWQQV94VQl3DbESn6PtrEpY6B9z
+pXzU8lpcgDWGAc6VN7q7XStDHBdWq4DVXA0gQEOZhNZp+WHVpP07yPh8P0xccA4VmSvHb7njZt/
r3g0/GeFyXooDGhBybjMrkjWVdQQC8tvojnTlPFgaMxkrr0bQ6Wov6mYQ8s0kGivdOFju3T9mgdb
ty4FHm5yOLDeDpYzQc27cOsIaY8RKIWykI2wKDTeTEoKz8iN27bKiYCv9Lwk0z48/d1Lvgjodd9+
2gA2dKLfnlvIj2p5SMgMCxOA2wy8pBbK3/HY5Ac2YoSWb0CwwChYaXJK5uMuLJiJig+EVoB+pF++
abI1FFnDSqzn1lNc0uuQdN4uSzdh6t9cs/fgBPu7yTJ7XkLMf6EP7sZjDfDIjMYu5YcVgpDbOl0H
eC59uuK+7dvP03Cc5sBj/uIi42slTUhHUDf/rouJXylibxewX1ngEe++XGUMIIJJb4ZhTq8f6zZe
CzMTBsDXmZSOn1V8eS5za/vpD9jS1CR/DVlDaeKKKEmnpa5nLmhFhpL8EzBpvEBPri4XA6gGXCYm
YjS0eUAVXoXzQw9sxPvyW1JZyjCAxd4Nxjj9YeNVTlgSGWnwmP/JMouAI6u8nV9SPz8DP1Md0Qqf
Ym6h+PwZMT34oqz4QQ1MuUNTMv0nEl5b7IONJ04rRgZF69UDxn7qIfHjCy/7v/FILv/y8FHE1Gvj
272wb+KUwF0i/2fOXEFas3YzYXvXaNhl2SSAAKc+/+fYYhNbOE0LWI9ewpnJvyKzQJkEckprRBrI
QpCIIMhGJ03Z530EQZeOQ9+2b8XpwtFPeMYx2Pl6sHP6C/jbhkcW+Zu/VIyAvnnEmmgQrK0R+yO4
p+lh8BKCiWAsukcrZMrvA55vEi5HQJr8f8LAePn9C+ReWTzkIw2wN/S6yqGOC51DG5lvPKBYV/j/
aMoY7TmbJq5unoxWFvi0oj3y6MnEcDPEcQ1c2Vrt2WZAfOeYIczvmCjdDcp/0qsFGss6bDdkJ37g
nxrpAcJAmcu2dJfif7Z7JXCcexVqvfieBRHNs3wV54OAP8HIDRwTMo0thpa8IfKmPR/zQHHcPrxi
r5SRAm4Nyfd5Gn3SsM6MuE3wdFUlVwoVO2S9MoAwNooxBHnqg6lMYxFAcZoFFawDx4fXQj2uurVp
9JduYlgCcRFXt03cB/L89phIiWCc6IRAwoeP/4falzg5IrVwa66XLQNMSSgU9AcR5k4ZUAN0J3pO
Xhzpfix0vwEP9bf+NjZ5rQtva5gthKDTcxpYkRxGv1wJ7mB5QJQ30E9CNjeyu0a8Ej8/D7xHXtiG
KS5Kf3L4KS7GP/QdXUadGF5CfGep7s0vcWb/W7wrkkg90NQbjJZOjOhoWPi3t1n8aFIOHaUKWtI1
Y6bV26NEGThg0tj9mbMu3OqGzmQE10vP8s2IS/ehrGX7hcJc64Cp9CBeNwI8nc+JZKbRxdJw2MW5
2GyilFpt0nvG92Ybu5jcDpvbTamimf3nuC+mvA9UuNK0ZAEC0wgcZZz1oB2dvL3t8HAoOxg+3Wk6
EPEq1Lda1HzIdb8WgFbmMDGDKaUqtCUxYMfs2THshbWks4UcPV66yGrs1xz/urrX1agh7fPsfYyy
YPSnTLno5Fv2XdPH4tCHGJbRp7qQtLDG7S9pj2WTBhUkybdccmO1LhOKhs7UFmQLeEEwKtj5IjHC
0jArH44FJqwYAJujkY7kbI8smmWTwCOXCRJ+UYi8/694mXteOryGrNv/zAeEZRhr+np9bwSO/624
BpXeuz5oFrzmCY8HELU6dAgyj7FcossrlBDce9W/zOydMFa/YR9QvO2XB9M0cUWrrHnIlsm0/44+
O7reiSS/RFP4bhOIdOvGX5nZg8sgYufywvwkiXRDNLJ3x0eW/3JRznFDh0NuHkHEsSl8LbLdV6Zj
eX/I3CH2oYZl96/QBmpdULgz5R1Cmt+0jagDpMP60GVAszRMeyylNFsP353kmQ8wDBoYzFnS1hvd
0/xIOCm0jERTISjFTutNrbPemB9f4svdE/CmMeu+h6IG1ckdc08MblnP2vdoSR5ABuB17O8pKIvT
dOmtfJXqWfz74NRqTtYZSnz+/8tSEviu1H3GFvDdDcBjF+Cqt/L2UiArIBCOhbyzVnEnvZ/lHGOV
4y9xN3r56cBex8twVcI2n5V3VrkUq8qzOWKSTWO+d89d2/kddb3firlqnTVn1+8QadIV+yxPXDMk
a32foiEo1bg8nK+wjtcOYpu+Ld9Viilba2QsTfb/dHrI5LXqsuR5ZaujasPG/OatyFDU6hNvwzXJ
lMNAL98w+LKhge0KnYHT4BNeuxp/EZhDLdnzcwvgOd2C1dcXF1Q12XI6S4KdJzU5pATsD25SJa3B
z5s/xYppJcB3ic8F1+YY6+3vrDR5A8e1DgzvVUe5O6zfU/PRdLLmVhihSNKnszCGgbB+9tT+chRJ
4HCczhkv3u/zA8Alw/YLm/HKgYR28i37cfMAZiInmYrPM5mGmEj2R31YMn3BJXoLfqjL9XVmUW+i
AdLChBThiwVCdWIq+v3HnCEwgOn2NIv50HJZawI4Q20fcvYsFJsYEFPNwtys+ZZBNI+vAVXCrY25
9w04QEYJ0TheVI4/wSfqIGRd0OtaXOl07LDZU+gaqB16vmAtiLNBGVTTIiIu5czY+v1V7KbOLKFp
9cAaPGPiPhtPSb6ZQA36r5Z/riOi+j/R+ycT82mPmHoDL1BKczcX4stBHYs8faNrRpjxzR7jvyBa
9ppuFl8MDAsicWPK3CkPlWI9YpHvnwHvizdzgHgT6Tx1IHqTUbKombOlmbDSYtAkgXjH0sJVoR2V
G/Oid6STRhr1ORNtRIQ2ZrTzJc/vy+/5/kocU0D6WEeQ1z9diFHwxB0LnA2311psyZp3Wn+hKZ27
zCOhPqHibKTzbIE28oIs6tE3VEBiu8dSApecIigv8eASNrNlxu865xqiDPK6dUgsQAmaXr5KIQ1f
FatqV0o063yKfLLJxU0TxWeRHgEfJYmwtCQ4kdd8PphfNM+3EjNDU21u7Rqp4+MZfETXYWzTVroa
QbYxB+m2m6eOU/DhRdbJ2UgMj1+GRJwBfySE9XAFzqc7NENC1pKIWenAM/gtVZ0+FeXyGeQnpP3L
9dCTzPKmYfG1TLx78tJSF+JAAGp5rAFshVROIOjhsaBFOaGRmp/Qs/bYFkTKSKCd6sn0PegBBkpO
lTf3RGmutcpfivJE9KnOAx1gA9huy/o+LhW+M/yR1Q+G9vR5iVKAMo9BgjZyVsKROT0wMGdrl0Wi
Xyg6NvoxaEZdJDkE73+TrDGSUco7NU38TzzJHs3D+cb1DGXRPDKKQzbSWIhVRSb2b1e/PS0FMxKF
1AvwGreBUqNUrpJHWN4eQbj1GCh5wHTRotlKorvvQvrmw/XsYLjC/PGW6F09iWx2sVodpXZ57boI
RHVlJ5+Prxox1dTRhR4OiCpjnUkunHoWELeDCVk0H7P1aWb3t9Ep0qVGX1REM0vfGyl/PwEpMKm2
jH2ID9GfVSXZ2iVtxWCp1dvdKkeBq27zO37sd0o5OrkAkoMBbKeE/uPaX93a885AD3V3iKtMuBUR
vJYZ2I4KKTDQxnHwO0cHK3TjyKHNHpI2Jt8HLfOVgqno/coFGUE2yP0cjJK2yjHqJPuG+VMLyahQ
OHyFsE5YWEzYjhJkTF7ne/acq8mYPeLnI08uCYZViih/Tk6Lt3d5C0GxU+K13VGyyfA9chrcAi0V
mSZl5bu3gzxvAlTL6+8G4y8xXrSIm2Jo9nhXdRboGwoAq/XNH67QNudqgmei/GecMD9oJS3b5Jw0
sHjzWcbv928JjgnlgWks/Ly+OjCUaPE/5qnbry6HnOX7x4hMdnyTMuwlT6holS5lgGaL3BfBwg7l
G+4XyFz/Pvy+iZTYfG8So7oudRugHKYprND6JRUp4TThpdzt5B3Zk1l8+1ycdKuMgSRR5GCGyX6V
lfISjCKnpRoyRacVA+aq3AUG18/06BvS4AnMVOu1xwbkqUi0aQ4Edhn6IgnItztO3DLWk1OC7gh+
YOF+SyUAwPvFIXQwKKzSgeKdoQ08PH9X/bZpUHZDKdMcund4v1q6FtdIqr7+2ov8AfXUq0mTEFpb
c5PWdaGAHHPmkox9DwXAgokex2MTx6i2IFs84aPg9+rfwdu8T5P4tr5s9noY+9+dCuThV47QuACb
Bx3xS/5Sx595xgY+dd7F9JyYC1Z0Do0L0M+doEMlAN97Cr3TReYdQt/56kd/20d2vr15WnBzjTn4
u8CLGDmQc5nRFXC3DDtmhYlMiinS/EO6xwDL/iFHJa9NgDOrWeT7RWAYyZwLgrH7Dad9OD9t/+/X
MaV0WzRGXGLaLb2U8CjqY7PBL7yDZpP+kDkcxZGGfTETpyR2eHv8GnYbDe8EbqfBemw3mgeYkEHs
1P2+mnsnIFT/qv2fkSYeTtFL9DvoGWB+Dw165scvRzCRS7JTCuSBz5SwSTm72Fe6Zkhd0ZMt1Cum
Dg4W1TDuVhooErwdlLmNSeKVUGkQ+6IkoFV6cn1atAwz9yDzxRtXtP8YhLe5z4JCKtqd4bYopmOm
4Gb5e1oBJuLv5nyIVyjh34cruhYQcCSBszkXgoMjPX6JGCqhePKKlFEsaugV/KgQsh4JhRJQ8mvu
fZ6EwCrQll07la7PBenuB9QpQOP69gV9udJHQuajVUnEJFToeU0pvQcCDOGqAnsGSkO3nJFT/vGf
VOH6jERdgCTuwHgp0tr2DZtwESHY0xJLyGpW/NYXU3VY/mOFmYA5MMAPr0/q2nZb7FBxFAwxhbwy
iNSyF5u95rc8TPnP8CTcDpCBEmStiAa0xyj+vvWviv1JFCTAXCVL2aoZL8RUkWZhGd6P6erNhBG3
Yq7AnQ4G/RRHXGzNrNarqw3QRqHGxsfoNzGo8lSyFhjlYWoOGM8fFG8QKq8oIPGmTcPh9joSlZjq
1HAlTtx/g8ocLULcOfyySBYh8SzqWAgVilPa+DypuXGZ83mZix5Qdobbo4Smlw/Kkn48HxZ/DleL
rorzndJszCfFjC3fWVpXrvI8KareosMQeUiVFYQBaURTKoua33kP3i+0ZW9u77T+Rpb1OLrzdFu9
UlVVhlBSZybyuB38E34mk8UK7WDP0hkfcIJEtpYRjtUxso1rlqEx3CKwWYSv+8ZQyUonEQq9qsTl
xREOV2LXIBdDgEWZtWYG2U7guaZGgaQOI9f9nkfcrDS9LlNmvXFiblNfxh1X3sjdwgMlFIx/avxc
VxypkEtau2kiKIz0S0DD8ucmO4JuKsB028cbIIJztC8Tr5fUzBTbws3dEZU8efGgpF06yXuVbTUf
xGLz4nDrOu6V9X5OEqh8X/1kwPGB/oT7jEEcp6RXX6y3gYfeFcly2B5JUfSdUYRQov4xmaHOhh2i
BLNc+WlmQu7u4ZfnzN0xotbfI1V/FZZVJqP4IoYkaN+2X/wt/PM9k7Nq3k6TQiMZSiLHj7RaeZ0O
0teiTGIrEzlpTb6T9RGXSSNY/oD3cKlcV/teaZIIh1rePNOTYN20oPN5Hh1/lB0YruQxBq1d6X+d
he9l/PC98S6hCs9jAZY/SSR0NYW1npbvvl0zC6dt8FCVqmTfoLHaUcNofsQF0ALEHNMFqsmD6byL
OiKzI7XWEvZmIdNjHjuV0TEts82MTz1kgno831n19trIflrSvNNOFyFSB1I+n9NmQECR3xf5K1xB
WShBUadwk+DCPrH9CciplYZdSghlgt5u/fTiuycZEI0+xVMjgKjAbp2XR0V8jQRPwq5X1VcI3WT/
5uZ2lby03Hnkcz+btAsPzgu4z+fdmLMUuT6NjjatcfuRLF9uwH2lTsW5HYJ/H9z7GeW9iTJw2Fom
0A0CBkCCc50OvjIjNZnPfSnxCDLyI64bGtHzQS93wQh4pvTHKAlGwN3+x6yzwt7upUhUJNZjDOP0
ZxFdY8HYtYnWIcUZqMVb2A5LlmTQvfFyNGb6bfIE2Dq9wRzAKb+CCq29rPsGpJXtBIcFcpaGch7Z
fSN+iTqirnb+KWPwXqVDufwZ1hYCFKVnEF3DZZxEm5CM3rFR1HoyRsQT2mGmbLgK0vU1XMR2Ru34
1VrB7rKLs1wazQTTfjRhiv8Pn8HdPOKDiJ0nh51y/jNXdgsJ1FnuoX8hih1mPWerwvfIolFdZr1Z
KqxGFdn1NIJaFqb+rTGL76TSoK4ho1+z9AoudIwLmPEDmHq9niDPKjqVgCDU1UsrbT5NrCKdiYhR
EHsk1ZkyUskaWyoqW34XZAs6bsgkNEGqwICfCMH+R0wrIxW3G2LQnvt2X3JDIPiq+axTZNNTRE50
AV8wP6h/uL9DJ04IV3/V5HciUHniTmX0FkPN73BjJScfiFbSqgT7uTAyBxrKVmZvZc99vB3jK3Kr
jp9zzljcxNG3PPzaEgmZIJYYVXPINUyNY5z05SGrs8iDUNOZC4gWAMuLfMoZiBBwiOgFzrGyQj86
fwi+YJpxJdrDK60dSEcCTb4vUsSGZXd5hkHgGTeDPWAgH6JcoaujAjFtnlNRHKOEhEyrwDRUc7aN
MqIGqC4uJv96lFJ9xy7Pm9BrzjtKEMlFHNoOrhAK7DfXH/70TpY4NGAo01bwgOerFxUhxEz+Q1+P
rWJhXd2v4LSh3KEBt87nOsgzitj9sT0KScxs5vxHJeyqmGz/D20kPJphd+5ok+X1ULoIEVal9RCX
ROjbYTaeYVtTJkBOvCJXB2QijWOE2frQ876YBO6J937LwZTKBm1TP4W8HPd1thx+xaXUuVGFfrN4
PHDg2+yb7BEA/abjAf/GjWNLtiHwhEsU4U6iJfexCwfZCbEHSXqEzp7CQNJUXdR4sLvmHwc4yEAd
qq8EJiNJcxNQ+t4ik7SjbUzxCx719c7hZEuI34o9adWRI3xkC2cIz47G8iKt7XC9wy1ErJqxM4gp
xM11yl5u/EwhjftWW4tgNykT6QkUqa07jTBPlHNda/HqUczpqw5C9HFNjcPLoSt7xzMoYly0VA+L
Vc6cKkLXuqhV351TY39O6bF430+IttztfD9CRFMsOjfNgRRi8t76l9j2p9g6WSoyrtH2lsG8YWpN
YGVD5P8QDXu2XBxJAKn2icrHLFQb42SNUofyO8ig+314BzsMjCoRzIle40VfMGkD3G6hE8Kx+npH
/Z8Og1m+W+5Xv9O8jQrlOpl0frL7dAMxtySbrg/GMBW0pi9RirvLH+eF5s2DzYMEeJ4CHvidWyOH
4cWjllhgnWBDfFJtkCr5nuSFrvDCGL4pUxWbsM1MRLSd026k6B9D23JDiwxAhv44SFWYtwg3YgxP
1+hkwc/zD1kYXW/6sKDxQs/CKRVqoFq5RGoyItpMWveoU4GfAOZY3R5J9a7opa8mgH+yQZ9W+xj1
pyLyVkAqJ6wV+kvkNDR0UC1FbM6e2oqOy/RKVF9hnMXVc5e0fCiaovu49dDIgn3lBtSh1qIJ4sna
vlo7e+V9U3Rh2Zh1AO7KPiFUPFa3XuySmUDzZrG6ix7YyAiOJrH6w+3peQeBCdEloW0sT3dNRZHF
PXI32nW6T/fv0ZuhW6W1JqnerI4wGugu9T2VHxXZE2DIyqnhFRkPkBbZ0lluu6LsBlgTs21jmwM9
v/crPkBN0MKS9Am2kxJytS/GCP7MJOtg8ouyV5DFEXK1oL/Js1LV0vSvzD0UDFYQ36m5LkSB72BS
vn4/xDXTpzyhORJrTzJRJwR1ckyvljKZB5vOCwjovkK0y+GHc42zopZk8ScYI+uLmeZM2Kkg1oJa
4L1DoCReXxJXcjmm2SYJgzviU5sXkrCuxgqXygX0rDitCu8LyHUAvFldhtj5D26ZQugCDCH9MqXq
wV1nffv8l4GrLRrUIfhV5HMh5EL2aIITUKqpXcvjDhO3X+Hy9sGr6xQpjHVFcUXRIM2geZUur1m/
V96Y08OvnV+AeJUV3tD4Pc58fBvK4mAmqi1cea+zgFL/Nxskzco/dVOOJN8k7rpxnU+krq745ZyY
7iqM+QFxHssPVEA9lfXNTns1E1qP6pHfYXbI71q0Lao0OQxVv8ZSjMbbw5UIVBl1eYpENF8M9DO3
8VQwdJytzgwOoHZ4AnGevIyCBqD26ob4s/R83Huthb+F7u6G65a4k0mDI1p/6cs5+5YpeU1wM+Nv
76qT3HrTM97h78M9lvkZo4I6LzYLDhlWrqMA4d8nSdHg92B3D49M6AqutRONgQU1ZdjL5kp2g5Ip
/vRH4NcZCO3G3yQ1aJ5gEUjLuqMLDISmKyWYXJYaNU5jHAsOEOIhX6JHj8GPJEP06Wl+B4Et1Zoj
hEAwLnj8mz6Dn9R/pIclCRYVl2pkZtqGcmBYJCEwPQ+bAeTffILTjTEEjkp0gfxOjUxI0t732u8Q
UQuX94YflTcxUrBazc+leHCknGIoZsMEhQPeKsdaZyL63k4DOX+cG+KOBygot3xWI5fTnL2FdmUB
jF2HqF+znEbrFcpsXrbl2yvYyMbIME+RaPC9IJPW6HZiyZ6M6tzLNpNlRVRFYzSQTFY2AFWSbgji
Jf1YpvpMOfuQg5G+Tynf1+hiaDqy6i4Zk19VG/jID4lGJq8RsS4y4KXo+gh9P9BsdE4FdXuVtCFX
XaT4kfeBsHGQqob8G8xcB8r0n2x+JclmGZ19D5HIRTOnIRwbT9wPwGnBzQYahiHnMnd3Wyh6L0pn
eeyRv+X+ATafD8mJIX4YuotzYmhDddIp1pxpRi8bIj3Mg7zH1A75ZW/VgN810awt3LZTeWCKlbcj
tTS47m19dTolxIH3EpFggsLfoHPBiUw4C4BprWodPWq9k4vg+RtGoBmgyidLLwEQo4Fu4nCZmkiL
ycymN1k0AMXRSgN59T/LHrvr57emjL6ZOgD2dttOn/ffvtP1VLssyiz44enWldobXoSf4NohsBah
2gaU9TSY2jlmss9br04hrIMR7JkzTj95Il8H26TPgyI4O1REdUEHt7jw/WuQ4Xe9v2i2vlNucQZo
Hy6tw3ldkL9VulViXr7S3D516VUqvKfKXgBuKi+mD37RU3H4pY7xqfGyzVv8t92DSnaUzchcnhWG
HS5Qedl06g4uEQK9e7lkBD/H2GYLjHsn69PAbnqxAX+o7xGRpn2NAQlC/tecY7yoAdyEIpNYY395
Cw4D5Pt29QAyAxYiT2/jBFCqZGQzLce4aaJR5/XFQ7s/Ur5zfGteYJPtNvm9PTiUKnlTy/oyfeXs
q4qLrbs8NCUfWqpOsv2tt4AqM/k37W6dqQI1Nw5672ELIzbHm9vUsP6Mwqk5oIVv2NfEiUdCNw0D
EI2IwBQ73pAcxWm3IzEPTKSl3GB/JvQ6YW5NCiSr69RXvCtCw08yZXtTsDOX25Q2jKEYyHXcuOS3
iyfX+oyHq09F81JoUwtJlnN4Tkinm9+JNCM/BDo4vcJ1Yb7veXJpWNaL8aQRRhzSfI5GBfxJ6Mze
eqIK18g9Lm5Lk2tSQOP8C4Jx5wmjorG80aumFkCLpcJZn71VvDZ2r/nkmk9ycH0vePJsD5xPPrun
r+SRlvHfQaX1yJY59m+6Ws02LwTmb4m0xDysB0byX1Bh8vm8vyxqAiwQcG10W3B/N+4C5xiLB9y2
0xt9QGrtIKJDdQBtD834Kq+2Qw2aLOg+r2u9ELTsmaMI8PTR3wmJ5bj0tAvKxMefTxUACVJhrusT
Wf4fIGukdMf7ONkxWW0ep1wSVW81oco5UUGca78ZRoZN9uQV9Ee7OPGKJh1CgC1yOPL5aKU6Lr2+
/WKwVqaFeFnTvQiqGO0rLA3WqH9mRD8E5ZGhAinYMMpSuB7IlWGVosVL/3/EvhhNkKAtegg00OmF
CApndm0EfylKAZepdK7KeMorvOVr6Ow/NdWsMH3XqJrNM1HcXBjciXTSTkUE+9REpbQry1dIg1uH
4WsBCscD92toZEHiYVzHwPJ+ReOV+4g8VsS/CcuzRIAV91Lses93YkbAuOzeBuMu9XwUlmE/Zqp8
a0m1jqySWbgHVOItRcLZibvDQ/Ys2cKFKeGFU7hWkdjfZocFmDOazY91PsjpY0L8CXhKVeihYvv2
0JSuESF2tLwPS2bHpHoJMxLiWa1rcjfLVk7d2GZcHgLXQ5lohK/NcvfjWUjecikvhQuZ5iH5CbhT
DvXYMIr14NNajIW8AqrQ3snKuJgOeRohrgPPRQB73g/MqWlL7KvZxuYntDwrD2QRMzwXFOFJgYnY
Mer9VmU+EMnZg75wlnaL8bwq0gizUj6tFfOjvU9RoGtf2azxtUxmzffWU6g79NM3DtyuPlIbb0TH
BUs5uNASnS6KHDUyzF3OIlrYp1dKhDV4JyclljYDL/u5m4cD32qTaMFT3qT2GqP0jt3lDkoviVZy
dCGb5FDyMpsUHGGQoG00IRFlaO6Pr2kuu1DnfmTfz2x3kU5tDIwXFVxS94rurcS940RZsETH0dMA
uFoM5k6cH13dFUMqIXk0eVMUCtz1Q7e6InduaEfUNKpOWhJLm+7mrYdNBp+6gG2gYYpsaGGfVpiS
WQGigR0+qeAyHm+DlHUgR7iM5JMILPr4iRSiwLLxuGsNAri6Xuu26vnXXafyrA/Z3WFTIqU21Zaz
u2nnlmyK/6ILRIOfadEafgi9GVzePm3Ntk4tiFWydkQnGjgtLTDWQVTFq5BWF88R2hs08x7zkmkX
8KlGAjzFg5djIuIK3gTH2qh7A8q74eSa+aqLNNEw6Q5KJ0cElBKD7HXGHZSJYifhSlRdWORL4miU
c9ZlUFOaWe/UyBuugmTOUzSuVYTZriMypcssvetRfa2hZ9AEU7l9t4d9BcIiasgYbUMZZqnHElWG
I1nRnU//PvTxs1bRVmmM4duc8T4MK/Nwj+FfpbhVgF8EUhmV/DtZTmZZ5KJ5zG8XljzGjkQ5eWtQ
uPqjRUGjnb+OnUvwd3/yaOQjwdXb/ERPSEPLmh41Tv13+zjA5ZdNaG85a5ZkJ2SR9Cr9UWfM/64/
XnjTCqNhA6IsH3fDo8FxJNBgqUSQywbQVSjSH12IFWeE3B0WCAsZjyMN+l+g/jhgnusgfCubULNG
eOUz50ssTPa1TdjFiVIV8KG+STsTUb+SLf7kgXhAfkMpojXaSZFwhRcipoKDidC10vJjYrzju0+/
fcsj77IbyaF3d3zDZf0ke4eZ3f/UEURaI83V3twOllnwRp6+qGtJNcgAycvmnSlenRXT5oyJvCXu
gTv7BZ5KQvt9as5yiaTB9lZ17ctFY65buAHzaMuGuCPF0+ghMTfUMGxYQ+kFvxflJJ6NRad/EoWK
5D9z1xTsyHILBqY3A3tnXtHH/2dVG1eAZFFQ54O74CU3D67sXI17tYa3RW0ply64SBiWWND3EzhJ
GNPXG5H/ZI4FyVULwvFJ4Mirs8P4xcw4mjJr3wqOVw63X3QT2PBHLaYEwp5jKx3wgJgiCqxMbcNF
XUdDsRij4DOOncNwkMDVSQBNTzqdcWCN/ldP752xoUiwbEh+sfrXZjGMvjboYKF1bCbNtFUcndrd
8BOY8ZFZvQV2X0TpgRvKd1Z4A8+2QZOgbQqeD/rmQoTVq631Iux45oI5dTtsoTKeqeSQPONPyHze
u5fnq+cOXWj1C5rMjrg4qz1ttM4P64hRl1nscbkHLVo7RTc4EuN6/8CabA1jIBK0DRmwhnXs+Rwe
1GVEUl7wu7ziWrNbdwf54UCZsLil+h95VaLUAeKyS/5nk33/BzhZj9OS0SBg49qgLzjlZHIir4H8
BjhgcEf0KY6fTkWOvdw91XgP+92Ee8lHMrfzHhEfPk7Amq/THemNdWzywQeJfnp8q9yz+i6iB+hf
f3BNxkNQA9KZa/j0vbPt1bHypP6LSicTw4RiWSUhGlufswrVFCNEkZycD3J1t/srk+FPij0G9+MR
jTGcrjOmfL8kc39CFF3feD14VSTftMP/9tc0DAw/UwEzoe5n4UPn+7yIJQd/nk8IXk7oNcyvfYmt
vrcNyY+G0XgzLcL94/IOejM4J1BJiDjHwsCtNH4FgawBxgtpUY9gBCE3IBaFtSSQppMUMVNMVubO
pokhnTZoIBdFiEldqxKohuvgHqQ0ggB+xSBaSXg3aPkOPJBpiYAEAQ3PT3jarrpE5MAsOO9DpPR8
foKmt9ZaXWyaRE9G1hdnKq7XD9vjRVkpWJQ66eaOlavbDnle951ytJxySAlGRc1V5azhU5nfQ5GV
FDObUwpO8taVPutOH/zzIYXJm55XBLh3pMFhun8q4LxL8uz13+5DijHY1hipNR1nsJf0vd1oSK6D
jl4KriaReUcgnX5eAE/ghB5H0jACd6LgWzDQ2mub0OEP2HxtXz67s6ZKTeALlBsdNPzLcWc+Pvce
edEu0N2WowdqjIxhZntW5kJSwuUDddlePTIBQQVGKrbiF1wIwyH/RV7O31sGcYmdaSUzbaoyKEAx
JNGx/aExAKsKSYsEYZ7DVv06pnQdC/pAZUnWeU8Jy+3WVYWug68T3t8+EDTyaxbXks82US/gQc5Z
BlE/TDORxT3o1QtcGxsS0iEaOEJ6IJT4x7N2llJ2XpnV+gMhy7lZqvSBJv709aNT5gNBWHOmwpwC
ZgfqKgXn6LjNhOZECQ/WpP2o7y31Jfln+pVh+O3gO2R3ubAXGLxGCRkkeGKbb1AJTgcZo8SEaZmi
WE3Tq9L/9t7gM3UiKvGnlY2jCWEbzzL7zbqnIHtXa8r0OQy678XLcRk7qfWpd/3CvPd+2bWi+UVy
bxxR4ufwEm1SkZZYvPYub2aiPPMdY5DWKUYxDHtC0Orzyl8mtff8qQVC3jTLFgTeV6/wYFcogXz5
KskGByuWo0p7NFCLmIHofsMn5h8fSzn3Fm6IAs6l1dLptv0ihXI8saJK0zFpv+8abnFrnSOt52JP
Urgy74Q79wdhtXXPU0VVK1C697O5uqOxA7LzuJNyK6r0kCwI5voU1tocAa+SVvNV7piYWdMvVzdF
AWmfVs8U4e6eqH2GET19pTnLwOti+oYyHTUaz5o+GoUvYwgOgM+UOze9DVrO2CQUtsp/weEPIMGk
j1jD6rvTZFeqai52HOrsuoG1HL9eDOw4Ne7xDTTbY8JVkrCc5YPoERy/NjFRiMxgiZAvPLYNYatW
2frVmieC53UQs7BDpGvsVPq9SldJpMEltNQrpmIda7f8pgKAhi3w6CS+jB34JKX1z0lQedn+F4IL
bKH91ECbWdaUdstIJoHvD1FCsN6U9n0A3wRPZ4d2Hgsq/XQHwYa0CM075gArP6vf9dnAuJFnQW1p
XdQgVL3gdU3DHHuR1KqBkruMx/YNf8FEXnD4ndOAWso5f2Im0xC83K+7cXtt5FALqocTNAz3ePA1
hnbkyFfVK1UDFoCYXWz2Ds0Ccd0FKlscwk4h+mJyyW22yX03n9YOy5md1/JEAqdbSFLN3HFGA+GY
Qz4P5CrDYhz8N73PS0Oeaht808d/ShuE5929pSQNlxhek8yq9V+6posETOMvkHA5dnoVCTk/ReYs
WwhueEjBPreYU1nmlGcDezTLZ+L9MpcXQoGmx5ptMxI0o+X4Qolp0la04hzlaqWiPTSj0dsm8xqf
SUaLsf/tuF4pcIJfb7IE0IYaYJrWTBPztbuu1PjwJeyoX24ODcLT49t9265Q5GXFweVpwW/jSt7N
CLu/GRqV+oRh7rY9S6K7rauDUOF9zTaK01Zcg/L+oGl/Cj/bpuZa+6RRwzd3+HznHno6wiUzw1NU
3NBESkEYSNQmxbco1a+VtTcQsTdRl/GoinY/0il6cU6KtRvLyS2lsxoR+nxoVjKCJoeV8v3ms4XE
qD6z3x6JArKkqr96t1lNerhnW/tAgmvbLrqlQ5teq662aOaLWCOgxuM7CSZYwxd29IaJJmXmdjsG
MAydiTtapqVcy0uIunET+GJ4toSA5SmLY1rxt35St/mEeNvW0s8yKy0s/S8Upx53C6//QTLrUtTW
i+z0bW8hMO/fISZ3EeReeZhhjEQOSlMI0lYKD7jhg7shGrPf55zroyg+J17NPq4cdrLL8p86pZcG
p8NfiVcK5oaHeLJCBTX7V+o1aXJMSt1DjVAPsCYzp0oVQwh6DzV9ZTniiYHz+7tghb240MVhI7hr
cjK78xAf64YkRlelZW5UTYsd2GkCYlQCvBkSehtLAdBlnzukmx9fjZqgUtU6yZbSiZ2D4EX1jZSP
cQu4Vrk13MpIdO/+GixQ+F033C43SZXrazbZO9Jlenp86p4EV9lP50paKRJclHqqd3GnoLzSFXWK
HH4/sXfjyTAiFqCBCGigPjgyrWjVkAj4ljTq4o3/0qE2GsT34k1Ssxr1gcY9eqZ2S9+wUjUuzJTd
FkUwV8eIzKjERc8TIxPZG9nAJTU+HWibivEtjyidYDguBMn8MeiXaiHpspCqppuSBLWdJULxLIeS
SMibGF557xAjsQ5wFr0FvG4nTyJ54CAw7yTuChQWBwBMFTxNhjK0MsmRGg7Vi8QyCPC2JTWJyNKA
IDDIkfydNUV73NUeicDxVe6joeR17Zy/LZ19+STOGwu0j8Ob1o+sVJMM8EkQCvTtR/9R21JG6OqB
ewuPgZlMxZOmOupzJSM01PKT9qXIu2yshOmOha13EDZByFzAAp/ms/fKqRhcTJU9WakDOt/hT58a
X5XVqU/zsve9VoEmnEyacDmro6VCHxdAunapTOCCSNPPJzHFa26YNSQbRf7C64TZQnjOdOUTuqpD
nmZA5KJJEuRo1ngpA0n2Ccuswy98XF/ewEJtL+brutca1eSiPB7AaIpa/Zn8rGX3XxunBxkCyBNc
UPwN3y13VBQq0vtEKfmT9JuTI7bl4F8rFZ9SXTWalCGkssNEZZuwcl/Jza1qtZdBU+Dq9butnj5o
m647F95Dqup15ex3dOoe8DR9+YxolgszkwtLFefgikyTUHzf8C6wIedm2k1RA/c5OcMsTkDngoGx
Sf9V9FfjyjfLaMkIGj7txbJHTzYPP3eGzSFRornQ0g5R153jB+Zsrjn8hfUT+S8PjgInwZkVbwIs
VdNnlS7l1xFH6Zhf8/rA45OVgD75llzao5tgfLP6QDnGYUzugbTPBsRSFIujD6El3mM9PPT9OYqk
azVdVF4N6NLsArMpSbOkL42X8w8X2m6VJzLhXjJjQHoIY/LuyByaVueCILSfZSR+mme9IooQlgtl
+pdrYBvn2+/vzZW/tMhyWrzsQ/JNPRWJQ+iw8yisGRiTm2Tf7FoUHe9dsi2glWDksnB8q8V2drW3
UNAlkVZsKrDG79/2lyKOCrt81moYtk/4O/5Zi1wUyl/bzyhbsWVFQtYWuYm617uVMw5O2AXPghE5
ar4k2XuL9L0d7dpB9fp8sSKgoJrF9zt8qmALyPnK5Ut1zuDCWnlAxJVlOik5t0vWjsuPDqtfGUSB
1boB4qL7Vf97CaLyCz96pPYjWLJNNt708soDPHjvYFpQOklsjmVPpX5G3juKXuNiOD8vzAuZWUeB
weAXbe32Sco95foBfICVgl8WE/9hS7LSXevhQe5JxBpq9tvd/qalVDgiWXbMhe5fMIDe/y5YlNTd
diHaYS6JRgAuMrL3Sbm4Wun5/Ji9KphdSvznsN58givYidpmy+oD8GrIEYu7FL7xHN7wRGRw2xn9
dscPKIpoEIfm3UvBzT0TXqUkg2W4jTHKImm/Z6vNHvfEdE7gZkjJ3uwuP43QZlWADQKYOWyG/8cj
MyfDVCWrCkC+oY2DXJV9JmvtWNtpn77X4uvsMRaepVH+8Nl7DQfCDQLsxo8krnDzTk32nbTzsTFX
5+wWcnOkbpwEQg4TTdNVIBI586eerliPUJ66ucLXrBymSzdMxwecbPwO86p/ULMWI8fV6hNZD03A
EhdTajcoUr7GUfMB7B5l7b829vgHdnLx4rMlkpgGrKKyJ8bnlnMCWKk3erxkxQDqx+m1q320Ykk2
Hyr3TynTp0h9H8Lay/0N0eG+9IeXLvVPu2oLLs6fB2Toqlh3BjB/QV8q4wLOXieuJ7cFrZMAzc6i
1ktu0c4KXRhQiJQyZeAxCShHGbHFNF0Lvu+3fSJJBu2ZAjkdAkJ80pmO6ZGMkJr1Lmz6t+x9HccN
PBPI8eC+2DIQDvTHuUru6lKyDTv9ZKluWtRDhMMr1ZTxf7bRJ1K6epJdUKgRrJ7Fx5Vlcl4Ba+QK
wcx1A3l5LJ+mbZdQMc12WzCRNlcsh1pmut8wExegMRW3mETjotfrS80+lJVlphIrO1g3hz2B459p
7Ci/0lgxvQ4x0/ouBl6JKuyZfcZusf+cRAVW04aU/S4cC24EUWvvp/yhTskqPyavM1Q5EpW3otQp
yi3Q7p+OHDwWQz8Jl4CxZs+oitjMvFZFx+rAVDEJtt9kSs0GjR9th0x/BUR5wewFSUP9O5kq+KR+
CRzlliULrW+4HPUZAD2chPuu0YXMYpitulgOLsrQFTsBxqvOVQfcg/Hqc8NznQujgtzaNTSFiXNZ
i1cn4pCBcrLsIgC0a91A0acaM5Y94jremH5NIaZRxWZ3yh3ZdymqVLTBEzrWYFjUuMnwhcD2uquE
ybPJ7VA8rjhlh+MfG79q6Qk60KWBOkBCxu8cAptk6TwKw8p/ksDkwnh1s7xyKtNOClJG5/YUKtB2
2PFA4EJpOMIGCep/BuoBtH4tDr0XpLLTTJDRzIHX7PzY90pg31VI+GNwLoi2m9lt3QTkrgLyc9Wv
eBuS6C5oP941+i0FzBhMMewFfyFdyIJy4Hpn45GLBGSK9TpG5LYszZXqJPtaskCgV7XMmaLH5i5l
hQ9F7Nr0uWNlh6zg6MS2M9Z5SgwK2orUCzd1ePfZdDQOrNlQYmCklSRgpOc1UywwyjErg1tZb7FN
lNrwf5cBIkdLSvTMHJHQ9f6l14vhoLJsxrAW/2RKFhrgKkHVh8vndf8lfaP8ksQuSAy4tX46cnKu
WJnlHW5qIqaV1k4i4+JN9+bV1y2hX5Nu06vFo2RWbku2rT4fMLl+1bUAOGpeiBFjZ09w9+yi2l+P
9lZAwa4JR0gymqwxtBiUU1fKCMpV5Sw4ZcGOzt8f1H2Je+Nd3XfEZO6PiD6lcoYC7takMZrKSPpN
NCjwI2Y7mUAP35nhseVmzZ36CnwTH2XxsmtKEBVjDsQt97a4xUUQlfpykDK7xInowb4aVG9mjDXB
kDFNRjxnrVFxgvS6ysipjIT8VsSv8St+T88CSsCmnSYmkDh1shc/xWZj1U42PjRzsHSz0HgVY4es
nZeS15Czxh7iBcxSwE8YohLJuTVJrQH8m6iJqIuF/QvxygrL2P33PDu4Db8XE5NupBDxSRL2h0kj
u8pKJEQGJ26LWCBgbBIgo1YVm1CXk9qER1KDYsL9jqKdXDbvk3aUy7Un04Wgpbo6k+cCuiPBryFe
+0+9W6jogAS0b7ybxpjGJhAEoyoeabzcgbRwVPHnZzV+7fu6rMDk00vgmllfmLubJgNG+OUEIZ4Z
8Fx/7cN9ydjILvjUy7Ez47ygDIXvU26Ib3/RI9SiX67T1pGlXSj8NGM85D5py94Cayy6vOeApCLW
b0AKKgSptQ+BdGOQp4VcdyFrMZzvy4b2eHSuEYPMkrJ6rCR6nu/Vvtifgmcvt+RpexvpXmFGCnd8
DH7x+JOF8GfKhFpS7hNdM5W0ifzU1bw4YVAAn1qprGAEd6axvtIdNCQXg8lnvzY7keHB+klc3uS4
31s6JC6zpv4jtQTnFRf1lNngc1YnJuaoHsZHmP9pAswc1MsTsH6wwVNtItAWw95KRbtBDUet0MkC
6UF3bqAcEyP2lwXGz4iJsZ5Lw4epc1oZeEaXo+FQpQs/j+0BPVpwCszbSsZJKfZfOjcu9zVBh87M
lxBFpGfOhMu5UyJZLeWlm5Q05LFiXN3G8Oz1y/RJcBgPAxBxAeon7rEeJSsjCOVivKBVlQovtzsZ
vgPAXd5OAJ6b/MH0AYZU9o+Q+l9HHssK+Dht/uZ6wy5h7YLv+P7CKGgZH6MhOaZw5PHrSM8cUqT1
sRGrPzCFiexpSQf6kcDcdOti/LlX7+n7tRFoGMQigH/i2yN9HbuQyknaP1sLxzTUNIqfrAReLAU2
47LYur+gbn85Z/9i6qnefDRXTyd0h730CY5p0TFXevfl1h6migQwOq+wwy+igvTLeqn8efZw/XP5
GT4yxzQZSgIdJy4vtRqT3N6jMU2DKzujGb7/JtJX63N/KTkzEdTaKNgocgaLezeeIYffvpyqutoe
tpSXD0RYIVzCR9GAzrNZH2oGRErRde+L6z+a+2JdGsGphwdqdQsz5zo37+DNJrLNVpQiL52iFGQv
H4TK5BkTC+lC51XXAfgukGjwbq+T02d+1+p/KsVSVgcZIrAL/yQ2daUOAShgTiHZZ53rMOm/tySi
oUhkok6+RNpi+eX5tqRtBto+8llXkHv6Wop3sJ3NRbRiHbxQ7wf0Klx0VF3B4LoUIREpD/0fFgc8
ihtNkk6PY7nMlvvWL9jLSIEOG+lYkCnshKqqp5gzHvWIIsR79jKT2aYqTIZUNtODEuccG8PBhrKf
qOtRa4CsCZgPzjT3uKC7O4gp7/CRB+tlcBEL1TKCltFZcZfogNryPBnV4SotJ72U6SZG/kkdRvwn
guDTcTy8BLzOafHf16SzLTH9KzTfh/geT6Jkavgxl9yHp9RQMgrUtoG4e1/NE6dcSxg72Sct/PHp
ZKn/jmhVXhi2/RQsE7pRbhoYuYyYAWgyfmOQdtjv1TSklSCdBGlsEy7mLoVQlwGiY4miPNgqWLa2
ij9JcExbPaqjnzIhEKHe8mZknAFkD1Di6ILToejJRE9dZe19M+1xIWeYLRqk/QTQZDUDkyBEt5Y1
+f8YLmGrytuaLJo+pun/pbtTBqCzA5mRCCmqDOm30mu4AFA2M6zx3GSS+U6h57R3ybXEsYGScYm4
xE3B/ey7wVeaNr45Cp90ODT38CteF43+MdpVkHwMVncoQ68juAdku6FfqrRNi0OeIGtm3c7+vpXX
BHsFep/rMXwxxiFqV/iP1PJ60rEBHWX0V5kkNLjFigl/Kgdn0xzwFinmAjfvNGTVEgovPf1nLR2y
34ARcPRJTG/3Qw/oV30ZxXFhbdu1GQyURpF7pjlEPh/EsDiVPl/LNurKKr6jN+9q4ktv5hCgCWVr
4b9QrrfwmizdWvjHpad8F5tqvJsrHkllmnHfFYeQvu039kuzHpfBCJeHcRsgqqI9iKQi3wfTWN3S
9w1xDKFKDHHMzMOpc7tu895Yu5PExkTClVsOQ5jdzTIuRzU5WZgbq41ZxvPfEXMZ7f6eepWiFc2A
tskZy4eMcFkBt95aHEzM7q/GotFzrce0SljUbAN5qD7PtLd7tkVKzt3eNApnUo1Er6PQyQf1GWiE
VVc3nMl1r/mco6dC+GFLrHMTIuwHIGto6+5MYnxtbFs9nhcZIKp2VnwbkCRiTdIJRULbAyTzdAG8
r/fBi5sVJS7W+BLC4bRxY+G8vulizmUDNDQYGesVt/hhY8G7/HAJkFfXoOJtEFxmAUCArFo7GaPg
DobPIXTQBHmpc/fR08w9S7X6qB/g/R/Ae6O5hid213qcg9q9otRsP2xkJaFyx/DTO/cjI6emZ7bA
SdxtdHHfGzgMIC3GgN4qIMORNW5CGsBzwxuI5Kj50/pJIl3EaDojJXB4A26v9CXQS9lT5nvmbASF
265GB6qAajbn4vtaEeJDoFJnZRbOsBbb59BKu47dzNitQgSwi0JdAO3r7CgHuLzGakL4bLbUq6Hy
f1bppLf6rxw2yyWMmb/pp061NiTlv8CGawI4OmCTWj5RpUU+Zl/gVhMbqPNHhiGvwVkboP6wuhvb
OrPVr+yAdWnX5iG621+UZZYjZ9NoeRAmidRrOE8iubN1vf5TEmgAioHhHceCGx+dJbOHYdnncALe
6S890XCnSgE0WEBvh3kkNZoeFlqVg4F988G8K6HBXkFmubVzn/L2PLGYKe2g9xrGV//bhrYi8b/X
eat9ZhcQIU87LOjuau/OpZvcbt7Ngr2YVlNzuKzelPfTGHwjmNnpL7Ywsh32fqHIkDCL8F0FmuLY
gc3E/nl469KfdciRfKnUweiCfrcTUncuxfkFQm4TyuaRFf2lK4UL7ebZCOQI0P+dnT5YlU2YPlXM
hd/J9UCZfU2S5urKapn4L3LatJIGCwU1g6qv8/ZcTX6lKdJXTCJxKKukJonNFd9jdw5fuv+WpO30
M4ozpUe/L40PKeO1TwcQa87B02c2YkY8PPDVbE0iSt5Do59oKbVBOXG9agf/1BcgSc5WLy+ePPnx
mYShK5WuRynoI1lwnQHC1zuWrUMUiRedz087tees5rRfZPSWsGnDRypDGsNkYMNRRqF03F453PZq
qL5ACyJt8BRGZFt5ubGRTSKqMSDeYiqSj+SbYUlA53iYI80s9GLi9EQAsqTEQj9+HSOi2GAejbaB
BKR4fYfQTNl5Jjs9KgILtH5AvxkoNEbwQZLK0f7NYGTl7d9AkcvfFvnPkFyv/YWw5QvcP5nRMjSD
6AaUFftNRRAYYp9DGs0TYJuxWKyjTHcCj1xhXwWrZw8mXFp3KvIC/1dGWAgb2uij53/T6RoS81Qh
DaDX96jvlNVfAN8GpZq7U6AH5eHK4wHaVRNUN44Wkis/OMedF2D75q85fSW9B+3LinYOG7UMSlo5
VQUnreD3DdYVX6alznzL6/jufWk4f+xKcBauhy7PwPEQoHwCjJxrxHMOCSFqpUnepxx6DnkjIK/d
zsjWYuhpzUGXDAcDZ1XFmpYgkuRHzLQ0VDg69mso31N8ZKR/e2ZM9hWXiUrg0L+5S/UFmn/JaFAo
YzdSymnoayoctkmF6RCTrz7impfMJ0n5OwIEo30O9jWZRrstsli8Da0pwYg9J6LlGFqtZEALGRKY
cNKwCgKRX8YsGE/fFqbecoLuZJWvKeHjoNJ/3bAXfpOI9SeU6bWth2wTyrwMmq4JTRzCwMWuxewJ
BzFny8rPWnLJsB9vk89tQfwNPoI9s/R2EVRgfNI1VhVr7U26MLkuAuFQgZzxPZUCyEqIfyac5cCw
XMO3LDus5lK07M4ys9F3j8YrHIrvpfE7JkNvwBpXHCjDlUahNtm+6FqckfieorVGX0jx4gSywXBk
4NXlpFou3n1dViChmRv32/PMijD+BMU6JVuGDD4w609I0jLIQ7w+YA7MPCumEPA7nz2ON8I03DcQ
xybxF24ZWKPsVfIcZ3KIU21yTF8j47V6EzU9r2fUQSSlF7tW2AjX4cPxFMVw4+8ZqEoc+XH/W6T0
/goSIf3LdttYwZ2CEDJ613ozghDtWwnLKA2DGmypv3xy+5HXe/6x6NjDegmJ+wYA5z86i/NFrPvL
vJeNpBVLNH99ytgik1pr9Ceqzj0XnirgGxCe3Vb/U7VCXKiUh9lAgQNLU3yxKCvKm7sNBkwVI8Lf
uooK2JJ0DK6xLcnowDI2gdtCT13ID3bx3ITEwFhcuAQ0GS6O5VlZ5gWMESr/AYlzV89KtKcE2Qrp
EYg4kL7+n4M4WlJHPdjSWkW/AmHx8BE4U0Y2dzoEI4f8Z1YrWGzgEinAYQk5Gq6qsVpFa192ZAfW
aXmyH8ziwDR5lokdW4XLj9G8dSn0vRTHmvpDtwipFGzZrWBWlGP+PYDBfMxKY0c/gnl2velbmRZO
Xr6unRGllmanTnPlfYlPYZdnnWP3hmaLpUTZkdUaBclcLh7GkR7x6KnuWD8kP85sGAAvfk3PHakz
9wzacYC8+Eeiihqnc13THIPWiPaFavh1qWelUvMy0IlXL2L8V0Y8sAtHYymzLw3wFziI2gSzqRnD
N5mqK0HOvwA1R06JDqV0sIYewerX4iQxWzKpb4a1CROnXqKy27k0VVrNwhrG6RiMzYdrilOQPAfJ
fDRkMlfPn9jfZZhveXsjf6Bh3aKZ8zKexKjp0aOTua9zNc06aF1IjniH47IH9O8C1Gj8ZzBxY1+T
yvS+incTeaKd/xY9SVGrHbubrLfcIRNVdNcvz9gzdkYY3H7ksavG+y6080RTd3aM+AyyaXrgQeN8
dKhExzhS9W5RNw3eAUsOmHDnqnJ8O4Kb13AA+NdMFMuLKJR1WlExsIXNW8lJiOlc7DsKooBDCOb3
wwq04aL5C8ZpjjdATGcH9EkxVQiyU0erzWFp0h8AHFOkDGJ9IzBd+HT3h4BtOACjqHk02IKI/TsW
HPPqXwh601Hcl1w3ZfkZtFaFe/9f8GGFdMwYUBHDx42h0ehTm9TMVo7dt+cI8YcUzx6H3USWuQzM
HpgSlhl0Ag5l2xs3SFY3ahOGAhBWqL/OdrcsbF2+HLmsl+tYLoICjWPfEOBHH5I8cBCZ9jC66xoi
Y++x8fL28xP1LipRCeQVi6kvpkBWQUUYW9j9qlNc1WuFI4XDJNXmTPCZsOco3n4RHvvFfc0Aei17
AiYlWg80eSegtYaxIqszK4Z06yXJLY8MYyNC+XZZobm4BpBw5wk97VdLo+A+USv0FyANbUog3U7r
6Nxc5k4nDwkf+IS35H6l7ew1d13e1/BPjQeFBUp0SEy2NMZDaBO6uZcAAHKhEPUNAdTyxsmNk9N2
VYTrKok5EcLlxMlpnZFI++TvTYv/nxZHIDi4Uao4DJcDMhqLDELzu9UWVKEuALXOCkK86suSo2hY
K8Jbex5XFrfoIzj3J1mNlU6Fj5nBj4+cs75BcMoRKpVPAaAhQZ6Z1n/UI3zDR5obwLD2E2fqkgwQ
RPY3W2CZDhC957BeNHl76NUovJz3XWl9RLYUWggZN1b1JcNLSJcDNAfkD0PvbnvyJVuu+BrznuSR
sED17z1kgEXkZvIE73tCTcrENKQcglIuqAn1pIcMAM44eDET1HPv6uD/BQBNURZ431b1sjwt30yV
6Dl2dBthCWqW3eFZ4WMS5G1svnGRnPd6P+iAfMxPDTXJdokb3Jy7O/9Xu2vWke64TPjq+dGxA8B4
P6rR+iPf5cyE/4s/LQ7Qigsu0r2oy8/llMnyQUdpirtmdEMdMcalcwhZUJtfTQqNdltko4euQ49r
RhfjsshskZU+ZB7cYZJNdLPU2wIl60oVyYRO8wNZBM/4zcbSgx+0gUCXbHLfmGt8770q5bx3/dxp
jaNecs8q7jhhXlfzcsEUbli9Td+x1layRZlrzfWpxr2DW5UxsivVSKhVhKqJmIF0kiWgV8hx0zgW
PxZsKr4+I4bC+anLxCpquoU3vFhixUwKpzPyPcXKGEXz4WHLftvxSQi0W8IBDmKTwLGxvF4gCi7B
Ycqh81EYCSqt5qgj3pcDNKT2viRZXF8aU/4t7FftPKHISkJZ45qcMNDZ2tn/AqxFlIIEt3YyXVkN
ArFdIWf1FP3wKnARuqWH5OFqU/9RW3s5UAWayR6DC2LDBb5d6xoGF9g9nb7gwI8nt4g28hQXRIOM
cKO3P6P/HcF4ZbTb//SV+cXHRw3s9Z1CXtHGKmuVZpy+MfNAel+gDvrsFdGKoVUJWVTeYakJKok2
jp3shONflgsCZ4/GYwqnJzSP2ZFs4diE+lyg/txWIwSUWoKje5fkqkLsgGBbuRbCeNazC8cHMQ6G
IWRBDGsHnGI3OEzbymc70ZpxPAtFVWIRyrslyIRTz2dJmTg2oHzsy6rxGVv304M36kwHmejwOtnp
2iYIXx56QL9hzxzRyCVvUDgGr1x5Vjd6qcSU25nvPUb8gu4s1RHUm8gtVP3g6s97IA9QniT3Rkf1
J6S+dCkWEboMZzI2/QJIhhZc1r0PV0jkyrY0j2aGbb5MrMFFmAYdu5yFzkOTr5fTVCgkMrEezbrs
CDeIjpFhBD565ekhV7WoZH50h+m0bIQcLPRordrFhy05olGMUAgHUCUzmV3aPpP3fFXpSkJtVFpZ
zT556g/ZeB15gv5cQ2DVwIEIsi3qUn+5qZ0hxL5nP8R1DzXtiroyDNy/ZqbzboM9UNFPNqZ1l6Gv
HRjJsftSZYRYHGLZ1UvEMtpHmGnC3AioJhCa5+U/ok3jLEVUmnWpYkqIq7HQXPDOZLHjYYlzTNBL
OqxT/ewrw6X/jEPQdd8PAjeXb10vtltri6xRsrrYowv4fWvuacm6ovDHVQbj4NmEREUAN+lhhhpe
qXBJ950+p2Se97JUI98LUg3pRZA5yp7m3NsVZbb60QPEhDpRmkaf7tOCznTQc4je+ACOfD3AE+bJ
UrAE/uA/5LveX+N/P8geT7qYNlqY2pdEbvfEeLuz/DIreufTrXZnGDA3ocoHiZqVVB+QjqLStfyx
qvBz8CIzFyyropj4OMB/TzpOdt2lQ60LtCte5yMqgaE3Ccy7Msm7krvVglpi7IIVr5bV668kyQXH
QuREI2UsD7iDWFIoiuIg8hhFM+40UcUVmz5vxLaZf1dHIP1zRpUjHm6dYb0bcmJXtNdREoJ1w/PZ
zR4lgtXJnUMo/vmnDm1SjRZ8LW8+tf+hQcN3sBdBQ9GonBXjgsaoh9as2blJBioreRyNC45UEuNT
vVT5rNwtO5nDGER6TD7iVbCz4dBtCy3DZ5beetcaMbfgyZQFSrKQdXVQOsp1UZYuxmWX4k2dGU+u
C8ycpSwrYvlbEnIFSNr/U7Cbl0nemNmfNqsQKl4dV5R6mQpylhbnveRGUF0WZvykgwo4KwlvhcEe
H/ISZlo5pVbaXp5FqwrfaWWojbFU/ApGEnr8MRfS+acDW4nSvvV8GX6QPazwxUy2Qn/cs6bcJyX5
KRG5Q15e7PAvg3wL8Y8Big1JF8K/iHCRqoiIEwJgh4TW9biPHldZOMyyWiInzuBUwBDJn4E+6LU+
CLDxa/+3vFVUGKPuI3hMdXYzmjTb0cobjYr+vp1x6maa+RdkRQqDRX4C6hgaZFKpXZgRC8cYiQx6
+i9ZkZdRfAexaxiuh4FiEAAgyK+ntzx09JiODaU0SObPvpahzDL0Mu8z/RkwCX1Kc3/n75pCEM21
uol1hDeAsE+/vT5UpSEi+Hyuf5ya0GhmLCayiPrS4Q+S0Cp+GSZelUWDWVkp+lUZ3k5l6wgzjDWw
08mc+L5djDJMpdDO52AeXBuUiXQCpYckte1OysLuy0WGH/XlLFXiFgBfeKEokDLGPbE/kcs8quHh
SgdXRl0d4LUEYW7JfoZsu3f3o9zD2MGte2utZawziumrxVO6BcQar4nA/rVF9WVSMvucLp61Gpej
6Vad2ip6NLFzzZ4+D0kRDnEhe9qLPyf1CT05KA6iypiOC5hQkCRkE1b81eQ07e4Ox7Xq2TgStvoB
1qUFmy1aW5NfJ45h0ew/h+CT64Q0ueJPt1Iw42va6XNQTnn1u6bEby7QHlhzpnlfvfD1bscbLNaG
tPr3gcLpwnWUVegttNeNAQtoNAbUDAngH1TstVnamUvhZUzFUHaagRnmBGHh/Et1IgBnoUO4E+gq
oA48OntXLu2VZkmKImBD4DlG+dYMlPoCcITlPewpW7nUyhTZsOKc793r4sFPnXj5EV4YKPDNTtik
culDzbgxPccc/3E1fpG8D1fecDqEYHjd4KbPiPXt9I1DcGuqy5ziZRwytqcrclSBX3nyLCVY0WEv
8ZPhrN+ZALvEFsokSRR3wTUhdCDyHQc3c3FSZnbJBjDk3eTdehmWo5qfUt9R7IKb8gHMlWBw3e9s
ZvrQ9wDq3Fu7mImEoM5DRhrvjFEM14XVD400z4zYDq0ki3V8WbN8dOheJ979pjG4t0tSuoLyRxmD
WhcbcokYcQxmVlz/23mL0RBDhL9n4JPeqIVR4CyUK1Nnb0m12aobvs2FuDyXYmWeHTzrqw1LCQd+
zYO7k8P/ypXuuRIxG/YBrl99qi5eogBQdKMNTwGE+HuVchK3lH4plyd0Z3laTxr+C+6BPKW5dE2d
SyQWdi94Rkasyv8yqdvpRSKl2bmjPQ086hu1oZBPMtAhn0jX6SCS4xtUM/4FR5j0tfjgTc8OfpJC
hPIhewxzniEUYmQ2s+M6YkqL3OFKgiV4Ycc2jnvdb1eLJMGlaaAbz9sRYYCV9ni3nZoTYZZjcMAk
onAu1qi3tLCKNMYALSgWSzBmRUzP8C1CDkmmaVqiEWEGleodA9PhSqulqAv0ZS/VYIDdnLLpRzLR
n8XoyiHBMccQj9/8z6qVONzfgbYxThKtmFQAuJYmFXv+iAGklk+Oo6hn4HwzXO10cZ2rEK9RTp5a
UYuSdKEeNf1cBhyeMnY5D+EeIcdDMEBOQn5eeiiLcl83SlOczWuUG0jO2h/fALWXgDLs9R2P17zy
Eh2pXvqGXvvni4tDo4BepkMNSGVW1C0An4cCtGfVS1s29z4IxzMvqOYYeqIH7egJ+zZy7Fj0Mun1
Zz6Pan+8WIGQU0mBfQc9w+NRFceTCKuZrVVPeYGMS8dAYJbhjfJcIeEOJ0Brf6BuUkB2z3uow3lj
tVTEobt06CvnZz9Wory6feHfWgH7dMPXmqwDlbUgAHaZdEXm8Ecfb1ZCCk69FlAgRWesBKgeB+4Q
zMLCdSJRopBfv0id1SRF7PENRw+LWjqOSnG0VOWVAsVH6l85S5qEJzWpDjldpU45oH7Ut6GGZP7X
xsLbadBGUVxtb4FL6DsyLCd0KWqV4iq3wuVnFC3oEpSkPHnOTRAJLD52OOhpJORmv1QayDwDDwUi
9EV3i2BcDA7k/IKM+XHCd24nwgNtuk3RU4tN+tSjV405xxcebVkTebemi28srcafUJsGg2/ij6D6
BZS7OPOpB1wyEhJrbp6hxKJs6P8URNYvO/5m4nXSx3nGKCcPRsMU5bhL/pM+ga6o97/kjTT2B8xA
cmRxQ6SdyJOn0iachwUx/TIeQH878BmYu7wyBtwd1YVhDqaAsc+GDRRi6XxUmgmmjpcA2Y0+MfOX
CpRDJqXND+DhXTW+HyVvjydAvZRoLy/0/yd65G6KsFN9VyXPF7wHOYdWMlYO21XGVrRje+YZ5/oj
6UeJ8da+uqRw7Ngd286CvfLitE3BZuQV+Psai7MB6cfgcGzqZptDjprbrR8ZaVPD2dmwHHCgMHIf
9tQ6IR3mzEymwpNvUIAAQ+9YQQld9YvxLHm5QS8DiKmWuAU3yam7mIomJxNIXbbvLXOEYVBCzOOV
uczqFwO+iJ84NGypeC9+IpDkCOMknDfCqzpM/rM3DoOytkJgQ6UCgzT32brzX9vPXmBmWYqMAD/O
GUU76vv3CLmjY4IRsOiaaenRtRV2+KaE206AK/2fgaCKiJ0w7FYRLIciRsu48GOqi2uUKSNdGgYj
TpkYrUonL0+Emc340GXiExgtvZb00Mcpn9ZrQ8tONpvWI2t+PaVORI5faWV3YYXadyoFB4YuwBwK
WbaeJyg7VyUtTzAjsP9gemJQ4HNFPVxSQBpsixoHCGplM7Hm9AHlGtcqEoexWH33eYwJaRiGD8+m
HSICWPac/vQnRIESAp+7kG4SqsG4vek4R4rUCCzObQEkMsV7+KG+0aK311c/Y8ZkaRiqXS/qxeZP
b32CgR4PGJK655OWT78+Vded//hxwy09LbhpvhTY5i4lueQk/T+ZdIKXeaUzQ50/mTILdPXI0Sgx
qG7Mlwc6/as9Ua4n4uM9/memYV5j1WYTGDTtASO2B8QTizscLFWYO+9OtHPOhdMEnRKqde2aI0D2
xmhtizpDeIbKsl2Givbpo4Sb7m5daXQTxU6iFk5DZ9LJ31y5Tuvod1l2JjbTEWltCOTEqPkL98Ee
M5Llop8NkZiryKBguIzRsSWenzTjTx7WLLdyBtR/691xdhkwBCsJOIzS7lx9uF6lv33WLkG+71Mi
1Wf1cOkFxRl1FyEADTxTlbeeaixW52JkPBciox4xThVOBcpHxNuWy7OEoqySEtMyY7QMlFPpvNWr
oQMnYp5sP7t4wSiWgw+CROJaWA0AggGJJ5fFsRfYl8GpSfOogFAphNf240ZF3RmrnGO7rhx/VPRR
2gxBOCXYr3OqHHae7kZFtxyYn2yzOIeUmRJM3Qk7ZiQAypTfPWQ/+KLdJk6/sxq3HGFqnd4CaKhS
jy5tW8tfYQGnEl9D4tJNcXPi2BP9DokNb7MkWWqju2x0kWDWdsOU8lOtHjhgRfy2CJGNgX3/BFHs
IGLH7ar9VbxRlYbIE8knulxNEifY/9zsU4Tnf2IVr5q0BOKcWmAY6j83wZ4cF3STJTaFzt/aaeT1
SP0no54BP7/2/FzuxIpQEWTytwe1LqdZ34hSrNSlRORmAVyetet/9f4UrMQdXpHmzIZNHFrvd9eg
j/tsngF3y1jvp+qJ7xKzCszcfgkYRMjfBYgl7XMrvhD0KGIBkQ0SYyMm41yNJ+KYWESC04Rg0YVW
e6hFvsaQadNSxrHL0gRG4MtWss6fiy2iYtAB5aqC+5qG9n42Ame0KLW91gzGeKGd+fhhuY+Cj3ii
gJ/IfbTIRIgN+Hk5jXCgeJwnNi2zv7jodgeYIh0Hw7WCYf32D0eF3IV0XqQtsSjWRAc8uUcjR3b0
BgDwDo9XkgU4iyl+1r5wuIP3q3gEvaRRRSyY64CsxIP+LO9Ndlr5bG9nl/UIECRBRbzm6fxY/bFf
Zp3pKXHvQxnfhFlX6HG9ntk5DAY6fWlQs1Nzq/mhfW4cvjIZ3h4nSawvICIsm7hqa04iOHCLHZM+
ni3b4Ses9aZ4fThmyCxyXMsl1kQUIZHXI9NptwiC/TJeRABfCK/+AnGtD0+zCEzLHyowsBnz92fQ
YbxABDHzVMNqNLrqF2ClxdE6Qd7quIDaaEiI81kNZ3o/EtljwuL6OwwaFRh3OPUxgj0QSRFZRTA9
6xg4Z1Dk8yDJfp+MOT4vJS7EfzsnFAxmTRToZplrghye1eYuAuYMzCoNeYlufYYXXK3a001haUVr
jiDVF0KiaSNT4bDcevbtC2Jb7e+9vIPWkapopqaKTJPR9gctKsCxa42SqkdQeuME1x0rH/OALW0c
o+ZaIe8xN2YolxIRO6k5for2/7WJmpG959xz5kGQ+c/6qprKypaHIG8bXEnpwsmeohzc8E/Wfg6b
yCtGttZOFm0O6HXNzxRnOzAOyQ1qfKrPHKS9LUsC7wfJCcM8+/MOp3/mVfDuXnVZjuJbgztxhptM
tnrRQIKhYP9jhQfIPQCDsf4JRMA5hqF7uYHFGnkAue7r7FN+20zI3sVXdHg+gZsoaTcard8mcNak
JhO+6XOZupQM89hu3FbBg4ZjzSxP8t6qqSwQLOSqoRqaJZZpzTLm6LprmcfUJFtV1qxmB4hQUxbu
a0D17ZXmhpNZQcIKakFG1ZokPof6P7x27E1Rhq0C/91zo6MsGJsucFcDLrDmgv1SFxzbmNyWmJyD
pxlzRM/vJxP+koIDsliQc4T4V4CUNA78Ksx4z9dgDe0SKtrb0NqA3jhGCb4N0KQkBuoy8rHnjS+8
/Tnvc8VBMwFYI3Qbxtfj6LtUzdy4651lRp94PfHhI2QU/+71Y2EI2b5m6OQklVtIKbe8zr4Z/r+2
jrNPSg+8HhsD8KpJ+khnpZjkDND/NTsryfRigXkHgr+/M3JAI9oqZb8ghMZv7MiUH0yIxGKE2/VB
g4scduIzujy/H75uiLh5/b8SOnrszc8WaHC0vT7ZajYCKnxULuhUfXpTNW/hCrKV8Xmc7Ti1GyR0
kEG8NeclYOzfOih+0bhtQ9L79j3eRJBYwwk0VFhyi/8PF+g87cbNd06pyIC7QPY3ajqktmaexwlN
C7T4Gf1ct5yFKCA6quxntHoS14wVz1womwL0xnFzwukDbvTvaWbqMoJmvP1bZ/xaOhf6UPCAL54J
RvUsFTwaB8BESjfTI9ST5CU84oX5dBL/slHmoWvnidl3o4Mln8xpkz86ZA3eS9SeE4jpzpoX8sQa
ReMty85DH7yljxkLuYAK0mtg//R2z0d+nD/vpdky7PI3Eow3e7eV1Gf03SKt8j1p8PkW8klIr6js
sHmO6qvQn6eDZItKt0xwUlcVs5QaIbQf9RARxKBL/VQ7mj3B+VHe2WKY1RIJbvVdxSUaK0pUb0Qc
URASYUV8skRLptGcSCN8sSlLGIe933NQJ58Jms6X2rLkvOY8BQ0cpCm9gmtjsQhjKzdLRGhfOLka
g0T/BvJonqifzVB/1H1H5FI2YpiGi6YD1CE9EZ5T0xBjM9BPqFVkl1qAoXBJnDn1vjfI6u3vj69z
BCHQ9QQrtjYul8mJ48aw/3HruYxFSw5B2zye0Rqdbfrdbhli8/qs61gYg+vjw3/rbbLlHG1sXThy
uF+9CqtSt0vH7g/OgTMQ/kh8KNtgUxwJ3GSK567NzqgdGZK0chT/GTe0ngJTJO2Q75IqxUPEzB8V
tenAFzenOcDBZlGJqrBOLPkPbp8C3e6QHQ9ivhjt16lrW3WnPfYtuPt/TJpuz2SBtFAT+fMDf2ZH
iCIx8OfzVkBH6R167RpaIuXaBCfFunkmhFTP2zf8c/ygsmud8RazQyr9nsurRGUDyLGevTEPuKnL
HtP5tgqMREu3UAwHkwx7TERh/7RTz15323iYj4Yyam9tTyDKGPYENvO9IgETwiKndsBAsYVltBiu
fBK8RdSisWQZuquR7EdkyS7ghvEOjl9r0A58pFJh6IeAKAV18Ixg73BqW9My5jE/IOiDUDvEv6/F
Ll7B/L2jR8OBT+BahibkFqmMqQf3NThHFNZN9/PUTSiRqBhZGoaLV9Kjm2Yuatvq4UATOOUMXqag
95WxuHQaaZc8XjYfZaanmxUUVa281+5RXwvsHre10nAl7CPwW6c0SaJ/aFcx62NG9c3XpcmyFYKy
/csROSYHxtE4oFQ4cUAi92xK1ccCpdObLD6AF1othXP0+jUISCQwbNpFDsy7iCQFsVuBX1slsL+Z
5B+kWuqPCIUvbsIYfiABfV4L61f8blN16BxPm/7fCsGUJ3vei6TSLHnT2MTL9NRILqh9osH3Xtkt
OQAG/MN6S08LLK+x4FXxnsEkPUnDiVENkGMRININY2avGg/O4ns7TzbCmHl+VOavSRPSmQGe1tCk
NrKZq32gi942dyVOKZPm7OPQuKC8rSeyEUieJ/VTkTTRQFxsk0XXoSzDf0O0x/WFK2JrRrpGzySg
Yd0J2OoA6w75ZBbeVceAg6gGt0hpDVHOSit5MjeSP1id6/vVG4qbG3+xs9pFkCDIDrYGl24NuZ6D
enDN2AflEs/d7HtxSz3zwBlr8HULnmH/gIci9jRcddbctGbkngDbdcPC/FV7aDKQ/cutW1D9CnoV
/+juCHXlv8nv4F+wuHzAJwPglhvZt3SDOVlbVBanl1Z1cbQiqZABkThpK0YIJULxaQjQm/4DenLg
wxv/KYTGtl7e8wHdBDKGRYD49Rn3WrAbM1undYei1C0dkGU0p5aNjCsNCOl5iy84pQq9Z8aVPqOI
qIZBViA9fBvrv2Ysr8yF1df/6SDBPA5KVdtUv+1oqSByv8rWyOnFbpksn4xSF7oBXrPe43Bbwu0O
2W6r8z/kaRdFjavCdbB09lw1ZxsMiGpagebyC2WiZ49zNiwOOg0TCKHCoEFl6SICNV+fxakchoZR
LdonC1khMgGYAkLYG4eJI5C6m2JKaDSI88s5jKBsjb4uG/d9PxEfLDfRu379dIpDLwXEcOyv9eEv
dnMKfpKsQayPCeFg7XflYRWAYCmfrIb3TD1vaOfOTMmZ6+faHvvQkWMlK+ipv6Dpdfzej7PW7/VH
eAQ99CY2TbHrtX/m3ruuvX0xMj12+J5iOBTlp4/HDQKqlkl/sFYkdyC69j3iTzLD/gH7En+WcnwH
UXo7iD+NqYTmMl9cuWUP9xV0/pP2MgE6H6FplzqCdSG6y3/jKJtecunH8Qqf6XfUW3dfUhBkSMck
Uzm/wZGrAGXKlXoZ1sh906OJOb+g5U2CwR842AQri4eKZ8VAa9RjmK1+iAz6EiL3OvnuqE9cGGhA
fMnLUvAr51XLIbBSUmX3XLhUmOCvWddW2dz8XPMgEOGu4Qr0IC+bZY1WYuQ6GZ1IeVWNS7gymygv
M5A/wRzcuagrwIl6vLfcYz1zm4WrC7tZWgQt2vkje5mTyClH50Ae0Ou3q46Fi+hNlpbhMpd8dd49
XBy5KEI269Tp/JwMTi/0wn0kr/6OwVc1z+fSDq4RgfrDHYIfiCA/dPiP8lKnVnNHnS//HnwQe7LM
4LSZNa9IPVLNvrJ4fNwCGTJBF8h4Zm91i8eYSZ7TSCQTDzhNj0EoFGAnt0+DZayL9JtTuY9RCE3T
7R+CZDwn1i3et2ty6k8G321Yds5Wqbhm4FoaV1MMNVxYtY+vSe+wqecl2wUy1d7g/SjXWdtdHfH1
L7QozyX+hd+uZR7UjL0IHxEvW2HSy6z+303xGGMiEZiajOVN3yO7HWhwx7+ul2K3Px7iyL6uUoiH
gSSvWlsZC5vuth98Fvghk/8p2b6c3+nW2JO4qPY39DgzQBl0EfqIsdvyZaOxoL5RZBLF0TTki1MU
fvF3BUyrDDoX99N5moLHu5qCNYD8T24hBdO1gzm5dV1kT4oQgE4IiBlZrECHWRshAOs6AkfDcpnI
fyNj9EuJ7J0Whs48UxX6s/unqY4Mty8qcco+kMr8lfumA6yIES5a/Ymlpda63ao8xFgcNBXVmhfo
l6Yq9NV3Nzf71Vydva4bTDFXmWFbj+CqI8WoI8wCHTcRJPg8+H+b7S9wPkXON3Su7DnA+8YfHogy
nGxyhWDQNLOaZncLaXWa20RETdsFYnrXzMNPMvaYkPAz49Mo6gvMXISRlTchQGJ9Zd4HKFs1gWed
+U2Ss4R/0mR76CA49WNue1YBQEfJK1X+TrCMPm83cTUaUYawfmNIE7i1zGSF5TQuqSO7W7cykos5
86j869YyGoHruGR+ufXjCwwJqKE/I6kJviSYLbw4cjGKYX/luo2u2mjlKJf8qV8ozeFbaB+FHzyS
iDQIEHk8JcgBYiJUdL/NySC/fNNiGqEbA94bjEv8uQw+GVUZp5hMNCDo4SjVKxMZzBthxYyWY6ep
f74uE1TotHGMj6sD1vz4cxovq4tKbqcY3vdR1gHcabMXihCvC4KP5e6Z17oJcz9itKHqe+svpWMT
CX/SzuEjgUaeC7KZXq3yeY4pXCXdjPYVHuNCGlHsMlgecpaGKqNorpsUWPGfYVBhqbQkOle4Iy3R
buv1fpsvAWKtcSUNDymCkdB/BNviUI4odDiNHoBSL+PipZaMLjEUCCg4WEyRC9W0vdoam3T2Ha99
cTV9pOJpj49eWUrGOn/Ldwt4SD/ZbCKMYUxc30JeLSPTDujUxDsHjCM6ZaAq0UOCDARweGp08Kk7
YlCaz+D3V7GYyV6Vsmhv45gfjH2L/WGMoORtfQ0aUuWS1QnhpTSh7Kc46yoNWAmqkYKraJHTXvat
op40qWIw8WkOcdodhWn4VWMGz1LRUadH7Hu/jcVQ9negn42Sodcxz25Ka9Kwukliw5SYtKQ+tRbC
rK3vXJztUe69VkhkHmuMThD4NEG9ftx90Z2dfI2sNjmvCgxCoySQRNY7GWlMCzQ50YJUcJTVhstn
o498UKEso6Ts+Xl9qXw+k8UjNcOqIQ42dH7S7qEBiWlsI+NPe76QljbEiKktzC9aA4uPWeepGEi+
KFeEznJPWnK0MKoujISX63JREoRIchxX4BLEz8v6AZH0OEohlEqCe5jDmkgCmWtJzONA+UzHFFfm
AJp/Yt+a69hAuk/VsVlYKngN8qziMK/bC4arEvX3QL5rVZRH8d+1xINnIuxwRbEnP0w5ZSWn4esb
dzTcZFIXD/ofWd3pwhEaaRq89ZtKr/KU7us+3ht8Xt/SjEsePN9J+GNDh328hmulK42hy3USmpHL
aRNUm1nB70RNboLdJb3M3roLjYdlUElCJ9Tfd3hMNo0y9dQg75/cxRngQP8KbC+sqm0glZ3bSf9Q
fxjMXNV4Fy37UIN8eCdifdMkFn+djm1gZ396S/d7UfAzl6rdWN1WywFHr5/EKDwhtiu5j/CI8IoD
W2SDqGnuMqEPpzAKf93p6BZG89UBA8ES3S6TTaaRG83Z8M7NqOwkRwgYFMTtPADzJSd3Vu8Zdesn
e8RBOOB3iWNsHqljif1AHPjIqYIJeGGSlxhQlLGjuIab5YNK7y2PP0yXynHIGRzuFGQGmdkOBLTA
Ia+m5njuyO19pOl8dQqr0t2yys/HrdyuEWUZj3SVUdgJiQz6vuIEHHKdmRm8BTFeLKUx0rDI9lWF
1i6U4TNhqBLen1DXl6INO+cHN4UZxrt7hAWXOHNScOlec1F8HdIyN/2nnkGKNshBeVTROgNWW5fz
O2Ai+zvEMEd+uDttXjhFAENUR1AooqinJH5dm06x0SNBKJL15EqlBMo+ZtN5hdRMM4vpC6K8Mdd7
r9y+uWPAKJ7NzDno84/jbRd6ySrbiKIV9RNqmKzYSNhMqvuoiB5PzPFp/UbEIXh4bVEIvHozXnPK
HtWCEwI9d1ysi68BYmpXPfImJvxv7mNcvRc8pd4gaEsbLoblV3bONOb6sq2LCvjJmz7QKe1BoJgl
kcIJ92X28Et6Pj3KG/HASN/3WSCV2/M/YNCeIYhFICrVe0qEKkWQ4s4YOehYPaEyayfIkwIj6qg+
9u45N93vvnrA/CBO9qwTYQqIlvv8SBNbW6Xz2RdTSZE7F2QyQUyUh4snA4m0G7wU/eu2VDF4cSKh
EY1jYl1OdgF9gUjfuOGzOyOUiJ2bzp48Hl+h3W+QaTdZbwLfo/NgOhuvjFWEHcJV7PySS2xsH1UN
gUg2KfxkvFgAaYtFRO5h2pejCA3OOke7owB9DBfS3bZKjQgBMCskJRSK0sUFWKvfQqNRPrL9jq/Q
LcOsBtEe1XckGlZIonA5vpT4lWHpUV8I7gF37i50BxCxoo24f1zF5v71LuMpXD6Q2LpOdAbf3Z0J
t/foOvJFzWtkWQW2HlqvFr/AYSQi/5qhzZfzxuM3ZplsB4iD9xXCIt+jaQfFNlovUw7cFrbbekip
tQ8gn7dm3aaboPpqNs9oNARjeGS3DMKMActNT5PR4OvVk+MlSCfF+4hHqWBhWstV4TEGIzAnoiWu
R7XYVVdv+t2HZy5EEwqgqJsJn3Ipta6fD67SheJZ6Kd/aIvcyyd6+GwNnIgZ/KRlSekeh8OycqDD
z5eJ84KkoejEkJbjY81197eA5fK2dZVkooisu8qjibqvt4zwEmEoN3b1k4U/FkMDzcWpz8iV7paM
e0FsfkpV8Ipv9t42LAOTkYcc/2xj2yg2qEv3HBnYdW/n95hVob5GggqdeR4uV+M7SpQgEQUyF3h6
sKLOcAG1jS8W4/Eot4lt8Tr/05tKlmeUWwMp32aAMBLCc//ZqOmOxWHfvXzDJPIpR4zCRM03PgYv
ZawWV5VqbmoEk/98laizeA/Ke/pMUh+UpoPUwwFmatFoC06nrFHnE1Doy78TzTG/PZSalbwKmaJz
pgPevoNFCeleYEKkNYZMOKiyRskfMTz+7l2bDZwdykzApOHOkSwukYaucw06wdiehs56uaSe7LCC
jOf9nT8OHBptALTgN99/rZOw00GtpVgDikhH4l8s83raqZy+OmdGQaDpNIiYfx/8GFbENww6fFfA
GPzy6HOJoknFqAIX+1R7plu//fNu5o3bkCdLbFBViXLVK/zZQUOQ8lSN+r/FoHHOdX4z+a1UFVz/
Qfw1tIU/UJARj5XtI+vBeEsIFkdSdCUHc1+c1kLRQJnJ9a46EIet8k/CphyvlhVrXcruQctAfQTV
g70MLfwrP2SRA/quSCQ3IlHBr3DkvTGS8AEU2eQ9xKCKQyAU0fwpSLkrITrcgBurKcp9ZJLQSZIs
2V8H3usPVK4JTZTFzFEibL86V3JodN1k/RsO5SDXnhpP5Bac+gP2jgEQJjl+VEpxsthUMr0EKPAu
iMJl/xOFyNMKLacHZY9po+9f3HogN7QSFgkeS20pBio2199B705dK3itKf1uID+A9fSn/8oAbUa/
m2we9k07jAqGq4ZUN34d9cjambqdf5lbTiuPBpNOlqTojoFJIxTqjMmwTHHNCV30n97koTv2YItn
AfdSmnSc+A8DP/gsbIZPLQBBFW+25QqeJLLY1Eu7xo/rK+iF4XEuRXsczzkId79TTCnk+tdJmmha
Iewf29yhrXWJcDZNQ/toJNzc+dVbYQdaUZkuM/x1Q/wsHDCZoF2taNWBZlvc7yi0q8AA5oo0MrQ+
UW5hWx08enj16jsoCXRpG4EGFniZbOegxMcsDEh0DEvk7Mqrk21OUBy9enUXlgABHMbB7csdKzsm
c8nwMu7Nr6QYZM1fi5kSCFaGZpiuQ6Nrf03888R3nN44T5BRIqlvwqFjYu/KrTPrLjzKbTqVquTS
qvmJUlGlhwA6ZEzjZfgme3RgXpjZflf5xanWnGMmvnH8hp/BvOx+/WSpiGG7I7BgF3Kw5caMTOI7
KlTJCfGKbUb3VFM7La1eeZeABPqUEpeC78ao1U45oBqohv/mfDEmgjtoFzTIkN3ED8kk6mZGHFHQ
7TfzwhrbgTJewNyUJMnuW0ZKzvn9Y+gF8cUib+1n71h92z/fMkPeTOP5ZJwkE90YY3NMIBmcDWwm
bSu0B7/9njiTO2ff6Pp/2dyvjPzEPkGRxEIQCwK0ScdoL+n/wITDQXngcEqiRLW/B2wBX/VnT2xH
qL0sEhZ6YDCyQ8VBFO+ummlgzbleNzmBmRtlgn58e/++hVox8Q5BZHucUhKuL2GkTSj+tmwROAOT
ziMP07QfhrgdjB7V7JFKohjJH+JG7jH5vkUl26YRS4MgczuXF0hmTY7gaWQsMhdxaMNLAxIm4lA1
GO19j6NK8F0GMhIxDydAoGG1ch1IqLQ8e0qmsxcLOn+KMChVJ4YDB/pPZWznxICMG34k+YRxD24Z
HeNP4fhYhQpTlO42Ee2kLw5JZrYX7buxpDuIlVPwbsnurboE456PGjlV2Tg4IoRXJrMRRiMltNZ+
T6Ex37erAQ8GiN2JEJuddzgKMdZeyqXGxzqJiNqG/77xRzcIk3xdY/VTyL8fJO7RS3gLDoX7ngTh
ud8kYSE0uOAnuoe/1lO7Q5jxO3khs1P3SFvpQZOLUcop8WXlnw3Vgfi19o6yKc8pg1o+W/fGWfh2
Bu/16RLiB5qz1B5DOxzZXORIYtqgv1pFpUXqGC2uEN/+lZNqY0NS0sJyVCesuIYbu/CQULCA8kWr
aBMX15E5Hh8ShNhOmOr5tywGIFZvWNMaKo2bjmZSoSGb8uZNyj3wiNpDuw7ZPWWm/qxnlR6qSvNF
TlrscwPG1XZIyW8t2sKTjBvvfCSCn89xWJMiOISDtJfprrM3W/btbWbJ8NsSv5NxB6LRxeRRsHMx
YXU2Mst+/tpbmfvh6i+3qgDhQXLrTGKemKZfD4i7EVgJE8p8fGFs8BLpCMhllehKh7JEGASFoSBM
aOTcvjTMq77W/fVc1ao3RFRFKqc5zinjVtPMs4Q2O7dLJA1ThwEsh2czfnAXpc2c6MDYoT+SbpZX
lAXs/hmR2wNG0IuQJyeFLjL+B9/T0tW6q7mjvsv5jtMXDu+OqJ3SsFiO2BPF16Ce53wIIBDggm+D
PdFyMYAqMQqAhBqm/KY7hjTiMyiPT75gfQvF3nyaUytugooNnB2Wx45Q0ou6E2Liu33u5RaWmQnZ
cEBjuEAxCJ0BI8XJSXWqJ2ka9O7vkcm6CLKks7Q/IbDF2x5VRgMweX9doOfcMBC3eKcOyba5C/7N
g9xvktog30HdYLBLhweIG8l6V4TvmkCfXfJutrIZY56za26pKbp1ugE+RDjb8U1Z92t9pyw4jfua
kFRMyDDWtjJdzpqJ7NIfHqhF+IWfS1iRqEOEDjNXxxv4kihLmaayrsh7ZKHaSqJbaDCCnyxBa8qd
T4FaWvrXtZNm+ZhtTP5yMxNGn/c4AgAM+5KUfVsFmT6/lykeMPROZMHXxsYhyEJYgs7uU/kGE+26
b/GwCQ197DHrcQknfen7U09WIZPKfSCkG4RWseu88J/xVQAYjhZiBdlfLcmxSm++GMyBgmbxg4W7
OhZInHZeP75/4EXkeOKbi1Tf0uLlWp3/BRx11dZapq8oAYw9IYPqdgmbytvMX4DKHLaOMxIz3Smr
tO46MNBO0euSiIPiRGe0JNe0wSb3ryPXf3WJfjrCxiVkuxH5dI2I2ckP+sj/jNCND/5Be/WPOkdB
dIukRU+ho4lTSD7C+Qim1Om0ClInr0EUOF305TmMqHelEWceUmXNJ479YSc2cmonqy7iRHv0Wd2I
DRUWIWzKTE3sSCxKxRxW45GcZxc2W8zyeOEdsC4TGcS1VcBh/0GLaR106T5wMRSJ2b2XWvntvDtZ
0IvLgi4j0PdRyb6/SvWMGXuwgZBdFxR/Lx3vvUSocQpotpN24V0MTJFFmofQ49jo/5qWjAaBfSb2
onHTRDjc8E+8VCB1LOOVlOxhTvCrHN2ml21lu48wsl32F0S6SC5v8zvzl8BjA77NAEqM1LxICKnI
eNw3P1teJoJr9BM6hVRCgJ+0KzDSimXq4ZU1/YLzytxATROs0skcS31uF6D+nB+OkUMPJygpHfKF
eKEAg5G6ELwed6EeUh3uJRq1Pl/AX7BjZb16dAxskjacVvyDpwQaDSplv71BwvaHurQtLrZF/W7Y
rDBMAn/2oNg0olNKJBKuRz56uNBxdiuSyLngn0/++qJXOl4/Dn0PaBYny0DcvXhSNLePJYfyntzN
q9JmJemLuhG6A1SyCXC4JCdv5gEKRJFyKKqFD1QoiAbXNZ9FDM/jR6/3BJj9kInpT9kwf2M1bTST
Th+W8HHvMudeTZdl/4XVp6E2zpvpkSfbcIpQu0q5AqSTtO1QnxOyiX1G3C4a2wHNmzm5srUPgv/K
FhHHzs8XQ+Se/1NOr81PHT7TtgbGWLq7U7ATLwOKDBBMFykcLK3EEUQAVspPRfJYWoiO90QMQAV+
I7XZkseifIJyxNfBzg/NpB+Bnv5S/a3BXAZlGfZivsQ6Pd48+R27pkHr/wv7Q0BUA/odlW4taklG
ddTlzBjB2HLZ9wNnwGS8rFRf4GZArCWYrvGtyrJg7ZnH32cns9N0lGE19y2fh966Xk4O0RihwJEw
QpD/jwCwcopdyaDFlURgv2gtKBFyZnCWsS0JduW1S+rtA8IrYsvXgf9WeVY+CRvAIpT4ymuYewrW
qHfmTTNPVaDoKNDxoJg84W2UZBbEWQ54HxqelQfonfmWkBogUlM7VWzDQyPXVzCStXIC9T3owyd3
K+XhHmG6Xe/Iu2jImaCyJ2331+kZDCCKt+DsY79Q3C5RJX+MBAaLYQKCsJDuSOEDIa698y+hM69V
hLrGAVLXZDhQsaEct5aumdb/rGObLhIojdBjvcZMIiuSg4dBdSek/PksFCysTzKCU/G9cn27hoAN
fFOAj6Xf9mbGRS5TI48XgiktqXooT7RGCDSC9YDNiPM33au4N791hSONdAbATn2cqzRKY6N8+8eM
amuDC9FEnk5fyFLkbqfEsv5ExNeLqCzdmrUWPLPd+Z4MOEa7UsDdLL1E/UQp+ucfPWLM6IhPyeLx
5AIb/RNKavDzQBZxDHTJvx/z7k40CN9hePDT2+bjQZSOhXTsBRlfUNAEnuJddHtu13/TP55rmwnF
YtfVWFDlTEoPDc13rHWp09VLhA8Z56rsAJwNoxJg1AW0DKvGXbuqb5KczRfmQVsN9H45WCnpM9t3
QilN+qYbYpIdpCW45eX7J7Dyie7R4n8H4aWRbe8WXaEMM3JWqTANrLncGuxE6rDcgqLF/oop0VeT
Dsk030PnFaMrc3O0RPP9Lh2Lz92pcDzW0Yhkx4xrTq5WW1hje2PbxCaTe5gvTKoCFr+d/Klx35M1
9PR9x3nE6msEWSRW5bxCGCyOyvKzW0xBIAzoolVRkcAl+44ZrgL0sLFNWeDYfDnWUjZn8QZaOwKa
G0rp7EdFxcWVg/rL4yc0p0KWx20ZO312r7/1ChWJqmURd+6D+MUSLj/fdOCdOexDyY2IO9pzZldX
TMuMMYmIs7C+w4OncUwn9JuYDdV9V1hP8gVuvlJQM7TdG47mrsIJuEX0O9lE3vS62xdv/Jv28cBN
kIDpm1qtZg2JIUkjA3bVA4Qb9iYaRfgS+sGPPw0NTJYpGmCu9BvcoBb6Kc+8aSIEreG9j9jKZCfd
Rl9oC8ooilYFprj1jPH/p6J1lDjRulk1Q8RcKiRCjsElaKdM4rBxXaci6ATMinVbJRuu8yDrF7td
OdGGZCkdEUuQ9aJvMwNIbfHEj15BnCKl0wEHezP1bok52xZaACmu+n652v4/4hxQHIiQhEjFAUcx
WYfUmR0Hs4tstynvnRsoG3LbWWltuGUVxlb05ntNzDpwJIFNVSIUBl29AH/DZx4z9aRTpAMQ/+8u
ED/oFwG8HGgWPQvwRm7fHpp1Rjzpend4C6pi2ZlVh86G8TZ6gv/huVkrOU1gOKn8Q71DaWPzy5ev
7zY++cbjijHj1L+br3Jys/nX0/DDLahbMAdRN3wnFoIvH6tHZThF6E3w1PvoDE+DiUfsxBr71Ojb
jjyDk9mtSoCiBGR7+6wTN3aKX0qqnLi57OwLZp6m/MkHsCnvnieMhynntY80tFje9Pe1AOLA1Ch9
/zBjVdVTrlPmEQ2s4lJvLorlcxyNCCnhgoK+foN3z2LxscYmByecYtVH8OxYyabPlUgNnWpSpD2t
dMjxesmL0ik0A24Ayuuu17ZKpZFiKMgrzSZyCQ3WlaYN5RNepSTDtFKIZXsEv8oPEFbTzuWNd8si
c+ttGE6+VtKjJpkNE5jZYEzY1txSMFffrpfCi2GePup5ip26jTYd8VENmhK2bQnuMCUaETsdQ9od
ltT8dcXneoghBNdcWqCNElot6GM5ITSgEaqiXx8dLfuYrZxnETHlBh8X9qsTfpYPF5Uan6/2T0F5
Vlj6Tgc4zixWHKIU2WmbbY3w+m2rEafCEsR/5zBUKXNv9sAzYqDHaF6qpbH24ebzRHeiotsxGO/E
naNyZG0Li636KjCxL1dCcNNZwM4erRgbxujWodSNSt4mWDe4K2ifEMn9Is3/FJemzip1Dr2glseE
kcHc+nR4R+ZYmWKEE6nw63q7vpzrRfDrthEkYq102cCLefnzJrfmEqruOOt7wNpeA5YPHXWF+Zk9
w/yevuDN0kWjfpmP0wVyRDPBfhIloJO49xchSOvJrRole517o9vuZc6wjFDRxxOQqJd/J5tu7+KS
hCevJOA4d5jFemdqmQGfxkHZB8NCWwtaBA5RuLl0Dx98niE/AyOzA+kYv92sJgUnzpGgDnLeTJ8g
AwGFsTVz57eN7YMmNieJhnxH0b95ePtVsOsNmdMgUWeCfs/JNDvGE9sQqDoVfGWu6jqwcD14nZE+
VheEvi6+iK9LxAeKkT2iweutQzEqVKuOhblrmFUph9pMcOEiAS0KCpV+hjDah7TkHidmuqCqJRQ2
O4xhW45qNtgTk3mtIpjXl08M41+VTV50QHI2cI0DsKjevJbJr7XbfbGEp0F3oBa2zuV4SE5L1wK1
SLh08WjlO7iEiWlpjglmuX2pDl1Z5FOb7g7ioDwaHronhkujSJCSWHhkDH0UC82MfwajMnMBhRJ5
rZo0zFippcy8NINxKnqIDGP1S/FSftiF53yAORO+l5YNizzpiX1XQjbH0JxDshU8pLGJeXKGvMvk
i8OA7DOpHDK55isxJfenyUKCJqTGz+qSGYM5zJcdcvYb61p3qgnuwvWIcngVRUAne2k5ccx6j8U/
dh5deYe8wAFRS7/hEBDleFOx/nUMSZxJoh5g1SSSn8qiG02kWHxhdVYlD//UbdCEgaQiDkiOcu/h
1j3TmI/DL95X28xqDM6oM7mIyyfHoNfTaNYgCdPZ6/Vno9j3dQMZAv/dfruUbGJAmznP30MftYR0
cGW+soaYkitvwhmJXAEyAmk388zxJizELOtf4iKmYJqA5y5IX8Kjd5mbaPmIIQIcsO2hQ1EztzE5
0z31M946T4MwzoamWMqrsV3xI/qa0z1l8Uw8lyLkBj7DnYDP8ocJ24d8Gg7h8N3ULmWepm4mnzB3
e+2AtJ4JEzIJaK1NAFmLBA2L/nqJpeYMuxxF6xBCJIIGN3oi5bjUi78BoF45hGSKnBFjI/ItoWlp
E+gT9kTPhdhbiJUm4JzpUPuetqVPhCMFTZgrP4fMTMj2re+MQMsDoht/1//CWwu1rAF65pUrroBa
Pncv/famq7WPICdvUQdTPNLMFyO7c9YXSE0hzeT0bX7Orft6WdnloGrMgBpc8Edpypgw8FE8rY5R
UM+44HtEH693UsxIupmxqU0YoAMh7NQdFsC/9i7TwbDx5BTW6H55hniUvz9BFMMuoTYus5iSux49
XW3YSp9bCS80p+WzXJz16V4LWIJkjmm5VKAc2YqqmJg23eKW8ACtnp0YwP+Znin6ZZKzTM94qrsu
W1mYE9aJhSNNEudWy6lp+2KjNTs68z0p+aj/8uK90dcA2jejRk8WFbWJjBlV76uT0jvrdo5Z34XL
MnyHb0o+TgXctbMJXztTp/FysjkWmSWg7TElOB8X9Tf7GhS4BymlD8ulqE1gwsCT1aF3Gc7h495j
cm+aQwxf/sAt3KfibwQnHul0D89JVXZgr6oAeJ8S424NAbUb32iHP36LSiIIIUuiF+nM0ATBGdJd
NVwU7LyaEjTAC7mKrcPtKUQ9/68jE/mhvDrW7YdA/if78lP7Q9tvmmV35IeCpOFC101E2FJX2RHp
Q16e7s/r/SCTmffgu/y/SsYKeDaZ7XS9wThOSI7ts74pAFSihM1ydWwlBT0RqN/gYcKVOMy7gmop
pRzq6tuQh9m7MoQhGJElWRTlUA8aa7Y2d/QkSoBlIDxjuUjzAprqFNOdOFXf3QuE+ped5Fms6oAQ
8/kTjBf0DpM5FVw44TcBYpTxvyvLhbxtWnIq3boyMa+gs7sGdRYAN3If79IpjsWrczJKigPQgGMC
lxl6TRqNUYrWxl4+jTPSj9Dc8twQHm5Z0iqRl9VfOuxyxv6O8tAtlq9G+zQRcj4VyyNrxX5jS9kl
hDQdWCshlXu97ToCcaSmXxfcxcYu7rqjXjwoZDCBRFIEClrWnp1ojpHecuhJs6rZCv0TNiRL4LsA
2J0YVxqrbx8BYhDv0SKijfqiQnSwWSq9HJEArtcs9TaHNRCoxdfdPOACN+NU0DzCG1Q1kuTblaaI
9GIW5KecNIWzdfkwq6cq34eU+Tq+5myk61oIrf16liwjcPSfQKQ1ZmLQwm17qlgRnUZCPCaskI8p
AXXUE7UcVPt6Lvltk6GW9CzILp9Eujy2nPfTAvFNmKAhfu2ouNm8Ubuf9OTyp4wHBHJWCnFL9UX4
bTxxJznLE4YNSiKrePbW8x7jvYSU9LH/pbOvCR+He2ZBxZAIaI145z09fjYxhxxsdf9ES7ekaS9l
DwqaMn0Sp0cwOE3k7i1/S4A+EyPR9LWCA40CeDcc9XUhhHfFLnIUh4Xs44+GTxyEfnSWp0XSj+Og
JDmISsE2o+2e7DNpzvQFG0yrJx2sA1L1W3Uq4nKyzphRkFOOyqPd5k+taW6NkYJSfD0fj+Uqt83a
9Foy6cWDAgiL7cNBcd2aMxNQ8gXmSGI99GHNs3KAyc3Pw+78zDnLJgv+l0Ux2hzjCraJAtgkn2cx
A5xRWCX68o6B2XqwlN2HGa3YOH6I1VFizV/Zu1lx6ge+M82vICJ3r/Xy0ek1ra/WGBsyUo3odvqD
DQlzC6l5yl4JBfb9L4OwxvrACDhvc2LZIkRovtHps89+OqwCtNlsb4/cZPM0ZjIQBc4wF1kVqAKJ
vtGRsI7lw1YaUT79PdhWyXbBDsjVx927X3ruJapUhfZqIulyU/1HD1gexKOx0lCdOQu7wvjY0O6r
AIteF2PYsvRK2RB/ONdqQcZeqrRM/az71P+r9j9CGKKHrQCxRGu3EmVYqQhOzwXOOyTl7qW1bxYd
IbIcRVdbAzXczmGHfAHLPe1UGsyegiiFoNft4NABq5uZxB8yXR5yeNRUbTarRpEK4lygv6QHPHoA
vLBAGJAaUscAYdWQZgioSWU22GbDGiyIfqn+t/IkERCbkSacjGtl/YNLC005GYXzl/hcBJUQ2tEF
1IOQ5qz85vBuXQepPpwFvmxd92joL8erJibjYbZkMQPg6QfGumSUz1IDdcstI6lhNnd5j2O5qGa8
yJf53p/pNWzXXRzCANKDcKe9WVAQTm2TBiHwXhH7/2uRUif7drxAyRV9HL2naReI1jk84gY4Rqtg
TC872a93lB7DtN9bkTZHIQ0Icqv8C3qRX1fJ65F0/7NPm19nkXIZaeatw1K2wgUxGXnYX4YM8lHp
oVrEFHH/SzLDxOx8dDdALmsq2WtBkhwUNhP8qhoOKgaZLfC56zrt2sRS7hkEqWA3AjdqF8KU+n2t
98V7Pxwa06MZj6vZRiZVOeSxeuzMQxAJNPR/PdTY/YLtTpQQ8FP1RXXBd1CceHmSay9MvZtFJ3+x
uGOOv7j4xH6VwF9FqqAhqjPceHLLQyckyGE6wa3bIdSviH7xN/4Ok52BCrwMPNCoyWNus1pJK4qC
xy+9YPS5MdJiOwum/5V8tCmGHwA5Lt46Zaq+A2eu6X8lyvuSZtUixpowcTXmcQrmhLtHpTtRA0Pg
MSw35DiiYAma43x8wLdIct6AAOc58HTe2T91cBI30geoLriX8kDvAkCOzVzIzSWdGJSUX1uvK4re
b3Q4seA197yHNYFOSbnUt8oGcShXk9RoenwE1QUnshkyswWEvcG9SwNC9yjrUrO6Xl3zs2FEGByv
jj2KzATL+wjNlSHgYxN7veYhfdVKIwu4KRBAalTQptzOiOyMGeGleJapff9HzRQQ/gXGBQ1MaXqw
arS4X7Nhb2JAZhVAnM/B8VyOCK8C4sYpp+Gb6YxwuJBCwvpLctuYIo/K4XNoXjr0CbYASiPByhk6
0p3audBz2htJoKbsfZaoWKXYZQQe5MzM610nX0p/cpGjEkDKvT4ktPxHQqN4n6tPy7CaYLN/yCeG
Fd/a9elkxYcLl+fb+lwDg9WZn9bLwCeHkT/pUF3A5m4/jx1/BIO9GIgnY2l2N8QsYuF1Z0Jvw8GM
8S+XgOfWlExxpS8VXcfS7dXYJrc1240hwAuNmPoMTefAHB4hk2C9G5gBMBjMi7WwJ6MsDSrozRRF
0gLsC+jxmU9jth4ec1Y7fjXh0RbMu9cZTTcgZavrePUstt524sy3/fijdo8beeNXgPuAkMlypCde
9mjd+ljaaNIujjqsVoIpbvuHqCudEU7QvwCMchb8yKAG8y/S+qwscST+shsgrgDCmpbcGabQN9cr
TUId/7jmioETOL1obuFlI3AEEqDw+FnY1rZUK5JvSwOxUNzFkhGThPPgChEPkIQKh5hCckhVBM1A
luQx3oCCmUMC9LIjQwNpzuo+dLjs5Oe0nU6TAakVJy8i7irClTMqPuOf76Q88fAXW20mb/D4hLDy
pZkuypiY8KZgT3o6PxHcC8BMNRCb/Hl99R5bH0mZF837yXQLvlKjPI/24vOVVAbgJL1zD4btytzA
DU3GIen1NFQEfguAypQZnJYCBCwaHOepQ4MQvHrO80M0zJoHpvF/0P8qJlNV/McVfX9d8PYnfSMK
UEQGjTLwCSYD14rDOb911GemsYkETqqPuyufjhGJa+NC2Bc2lyjKzO78ulU63lvcMxT9GzSI/T1A
q8fuvs3xv3mRwjVn2oM4ZtbRBstyrw8U2EOFXgj+zdST1mFZx2lEksYODuJmkEbZ+abkwnEGZOnY
O0UQJi3SSOC4QwTlQ7GI4dnGQgX2MgPHfHEAh1nwCXtj+vf/atcOJhPg9qpBdAOQRjj5bVxJWKP7
fSC/jXZF95UEHtVoOsoH5KxfjmQsEDoDbB0DwqSPCHFv8KbW1hrJqxkY1Y9v+bxkbKwc46Nj6hH7
jBWpankN8Y6jFU4ftBBFV95hP9nOrhnMJ0xrfuvR/ZGElRuLIeEROaD+OyMX0HQ2dWQjP2Ap7ztf
gxs1M1P9t3eB7OnXjAcZuoReI7YvF3LO5O8tpkrzkJ+eppl/E6P8s8HZy8HbWMu4VfdXnySBvMKF
D2FOXPJ+PBY+GqCkqnaoKwMuDUoRf5O1f/8PzC22/fLdpPLOk1EB8ihBPfIO+O4hhtFPsw+/4JXW
9GBqRBNej2cn9asrL9uotwmuy74CFjxM27OY5XsdlCYH3mVlaqPlsI6xR8QEpG/s7Dz4zDJ8idxr
PT23IGX5WEGkAUXEW8sUjX++lmbglC0fqOzGIccAi94K2Mnxd+qrD4rJnFFEgJp3ga8ntC4DKNP0
8V0od2SXEFuMfHaSoloZgiT3X7P1mwyUL6ANuOO2+MpI/GR0igtEfGFxxM9825FLQgOAwggjOtA9
kfC51utnNKuTWT7IHVfLCGWmtS65+WOkUEo99aA99OTzdus1OLMlDJB8iUBDC4+o9dgPjDRsjmCL
ihqAbKuQPboDqweLzn49+OMquSXXEORbJVHCCoHruXWQZlLH2PxrQf+K38UYvjrk+OEtp7NedYPZ
DTvV5n2BrA5yJg29MHF3pAjU4DMU1e7BShhyV77uMXAyi4RQU/Bq0hE/DpQvcb2jQ3U2PCS7vJJ/
h4Q4yyyvQVfIDwkpoVqiyb3zD7ox7FUZgHtFUIvnarqVxkXu4as9GUp5dOO7BZbJ05BR2ZxcoFZ7
y4h5bGXuihYQsF21Y9Rcj/r/DuzJkbTav/AaPuWAbqn24GU2CUXDKb8u6h9vIa8PFsnmR+YR2IQw
28tZytp/N2y7zrtMa5vH6WpiQusQCCNPDINxpi6Iqh6/Vyy3eRu2swsE6809/d67hW5JNTXAiNvF
Qm6XT0wYyD/lrGTtNhn5x2hLCCA8TIDUDZSKaqWcIOktLPSotyGJSPLqyBg/KNCGDrJ7uRzsgCLl
oOj4U0n0dTHLftHysR8ldr/y/QiWV56e19AEBdTsJfITpQo98iA6uMPctgPhCniP29sMZYvZat7K
eVtBn5L3Lk1J9oszXskb6GVez+hS3GALtmF/f53uHW85Iz9MIJi9tQkSNgzvp2UMx+mojMv8O/TL
2yePPHyVvuDaCTCMNnv9BVrMuuGyuEmQWkX5/UK3qoUQ6MCTH0jJqod3PVsLYKuhyPboq+j0w4Ak
MSCN/pzY7cgNUU5Ss9N/4mXjSLdkIluZRakHiH1nvt7Dgpz/HoUqY2g3isopq9adPIGNGpKKY9mM
7CyVk7C1w9OP8uujFQqPHGQGOcAjE0jMPuOQhlnRsiCPfhiu9LVz0vAOeWsQdNUlChJ7ZO09DLdl
44nubF6Zb0IHSEn/IiW16JBBhTFhGMpBAk9tuWG3/K2/oXKIENWHDZKyyftae8fjRiqsnu27yZ1K
3dkFmzI9ju/7vxclrwrj3hPZ7Wa0wJujP2kRw6q7Z13hguUT3CDQypn3pA/6ErSfg/hOYC6KhU2c
9Cs+xWGIKo1iiEcRB8ZEF/xs0UV3Jr5uhQD5fSQ/IJycYDvEJ1zYIJSZdtsJqJDxZi53Thkr3fud
85FGs5lCyDfCJzBNjuLhfhHVGDlpypfN3la+z42yhWfax+O/fPvmgIWkLUiAGz08OByXZGytTEb+
NvnJglxTVKVdWQJqt0CWw+vDqhehbzJrcpGWQOaSo/G5YU6EWPsZ5wYE3C8DHqODupZEO6mZ+uhO
JGADND5O/aOvBbdt6iaJBgDtirNsnrHkAM0K0H7lmhNio2/Vq9/6bx1mfrKL32kH6pIC+gJhdOgn
eodiKX6iixwQI7HtxIKfSWDrSEb58qtsAsQI/qU9ZuodPD6QBjswG+douHfMtAErrhjZvlsGrkyY
uu+DuUzU1e7FeETaIalBeAUqCwcOp59mOfhAzpd9UFXDaf/qQHfY55l3oKYlFNLBN3mB53E4eWfS
G2fDsyAyOExzaGxj1jM27rZf/ReIp8MHqCAQ7BYxrFEOSVPWHzjAj2ElVHzJKoySIpcBmzqotgaJ
IQj8UQFDE2P8LqYU9HNiTAHP9ull4umjkpWlyUSGZB9w9tgN1+yfwb2qweLUn10Mh2ujtGbUvUW+
JZ85NpNVGjxziPzgYwpznAxmwfRQ1QTGqAJ60F0v35AURcHii5f0HjNSi6jvS2/ivahEOB0iG0uS
zE1YOfTykBZU2no/FUnWj6rbpXVUjkSPbifS6uCnouGWnZsCxoYrysLYdORQw2ZU4/CDWb5m2t5M
gOgaIjtey//DVyXot94xBuoswbNycMHwU7rFvVnSlhKoNQtLbz5v3BFUbPC0ghsPIlysmhXAQBli
cQwrH4FuuPwNuXGhCmnrdy70ID/9JtxepKZfeaWvlYcl3VC0xln0iSq0ZtZvNpT95n6xTypSaDzf
ZxzWnts99qCeJwwgGB36JNE663VtjkyceFBncP1CH/VtsXKq5DKKtZsm+LG90kTI3FMQMl4jna7J
OCsG7HjYRS0ElMnuFQkP4JSkpYf8brdCxz7wPYAMzP/Kustgrt1/wmuD9841d/jteyoF4jdQp+9j
Bc48oZo028IltFPSeHAc+PMjYL7yuaY9Z7FcdjTWfYBlJJj0R8IPF5yIQqV0yShJpWoliaw+taJ3
INsuxIpZpJQMuugb/ZqnNQpLZd+yvVfm9RZH5ootqDgmnAWfxqISGdx4x21TjUYRXQae77jPWjXc
doELEVLKQ2Ic89w5deliHrthooZRbQajeD+pj0KxkXFDXADR29VsUlWzDNIwdyi9z8l7EMk4+6Bd
pfvQOsXO4YK6KC3SkbWjWwOLVIvnZTjOKNSB8ddhfCVZ+bR2fWQiQiSJYyATqgj/mQXMIzOS5fEk
8iUB6HUyygdzl70nhvJzGY+GTPLq17jDX2ipBX4SrB0Qef8urUzFomm9XL4nTFKM6iM7OPg3Ymtb
eIpEQTKsDjsT36QZCfZ/5pyuK5dstWabm6ZIygMA5Vp1JG8WU1JJ+UqO2Xc3gawC3OpuzcROI6UF
fRMUrlOK/bk9LntY58+7tLd6OMBGFSJUNSO2W8awoWsqB8qO3XGHXrR02keubguU3z0itBUXlDbO
u/JIPwFpw/jBOsZyeAwNCP1JGj+6Q6p1tXzXZV6QQELwYtx3JZTAgapGYC8zjwygEbH1azbd9tD+
ExqHh1qRgwGI89yZ5eSe9my1P5THJeFOPbCFhs9upXkCfNjjUlBZNLar6vYrw64Va+fyYY2tCNoJ
4ijB0l5aQE9Ol1fNv9vZE+68Q4lizNUfJ3G25qu75RmvhSWUqOrxKHb3CXEVIBEmPH47qnYZWs6g
VDVKzlSlWgGsR3JbIcFcynMCxAbnYRZGAxv5we2wbsOcRQoe8Qh9ztMOkLcbY8gf6MIlWI1mDeVk
S7vhvr8edFygC7XZkwFg1atwOGQRBGfnCTm///LmmekNvMM9qQKIGswsVy+nADNFPKwZMjKvkMrA
DpohWQ2xA3/7whDPdad3PrfH04IeEjhUsbCPoDzPqhdT8fqxIHe32NHzvzi3us8F+haMDbzOU6km
NQBh6kCDUUmdKEydXvlkM9KKhMJNe2u7S+J8KW2jgj5LyYEKWq8h6tSwqt3MP3kpQN5U0TwAYFLp
OkDylO5HxZHK468RA83Et4qy/Sq0K6xz2kguFyf3U5aNFLigOrQdz4CEdSQ5yJNa+qUomtT3B7TR
K8s4f+NRV+BSS6j+CCCFgfZ4kTOc+9Dj4mMnZf1lOgaULhqbGbbKv8vDiJmZJ+MUKCXN1KYoGNSd
eae/MFVrk9N3I2OFIV7EHdA6MRkaZ2X6+V/h+LOJNfPZweRrAoFoFP3JTZLhW2/5X3n+afZHBR33
UCWotSSz7BynfHEXswCkA3sBfAOV2VXXn1BktS0dJD2Sh0fIMwN6y9v/QPax4Txf8ayzda2LFOw9
3jc0oh5gQmKW7okiKSvloK9eJIwMSM80BgmSN5g6FNUtFjoKp6bt6YsB7YmyjK5S5vVbebUtFS6b
M+/8whn6aPSI6gwbB+bkMAtngFZUQxydGEuMQ8KdY21KN7VWcrdYSpzAdJu+ix5jSbhMIUGN3MOQ
souBAC/Qa5QicbaHNA4x3OWhAR7eIZFijd/ItIS7In/rOkgYwyQsojK2W+lshZo/u6TN/i61YT53
7GKwm6N3IbsizCCDk7Z2dmMcIIoh6J/fTXF3jk4JmywHl5hzqM6MdcrYxhPPSoFmL9sX3axpvpoi
pTWdoxx/IvY3K3TMvnCtU4cKmF8B8JauVGxI1pJys2iN23SbvQnoLHh+mB51wJgX84IEcP/g3/Wh
EmNKUHpw//OX6nV6Fw5iDO6HNFbvY0nWGRGkiRlOsNJBo8jHDJ5n160+njHeQrSmpLM1S4UQGmK3
ZVDvUs/nsC3Q9y2VxVUEkEfviGE8efV8GwwJgUlRZayep6ARdb6KfqMnMRey9gK1vvw4QihfwvM6
Uz/ZINci/lJobLVsrZ6QIiwemOR2JA/ceiIg3fw0eg0tkfn0qkGsxacbSg1KU9J3w6nMpPdxkzeH
iVW8ThGdSeRbY1cOVcZcyI7nSzc9t99nwk6K1uzQLjVVqwn+0gCR8RGUGCwQCaHq7wOge4NF5rFk
Rxkd7hW71ukHCg7OazsKp4zX7xnuF0gVL0f6UZG3rA38mK12dWVzWvV5162LIQxKjmVdt2cTEd6F
x637/ZjGHHNvmnNyPTxbODrerNMY8OnM3DNGgqo8A/R4Z8xt6DZZJeqTDsd2aBr5bu67EdLvifKM
r/jUlscbyoylKpqx7TsN9QetoSLgGKGpXdwhPNdO1Pq/5hNwAHTj018awKdgHH46PLx7PTeC1ab7
WcVGJSqIxoqbVASZdXYzDe8qDOPMDCPZd2WvEppXTjSB0SyD/YitjQuv4AU/J6anhAdrHzVAzebE
RlmnKm6Js8ZQ8JAy5OBVqTvK1NoN7Ff6BxmB0rrUt8AtvlosYUAjMyJxEn7HofbnxFDvjZ4utX2D
cyG607zXff4ZCbFn8SypBwUGYngtumIlEpYvG78Ssr4bzKXmDbw7qcSAhdL9SoDWVvt9ozMR/4rn
whe3Vg6I7Vhwx+0w7wmTeYxTbXxhxevucJaGM7xeVpSG/slbxe2aSiG0Nx3dS9ooxYrp7xO8kZvt
7Wqslise8BKyrYkszLfPF1jWk2LQEyG9gJUwcJdZeY5bkpPEGLEDUgcbAIcbng6Zb6+viWpZKUUF
JzC9pkjlpaU3bi/3D0BbH4+sMSeGX8/YLMtbDEATL2YTxWjxBLKme1+dxtgY+VnGP2J2GIrBG52o
3eDkGRoSSvf4noJukD6yNarqhQNkXI59vahC9++kprySEhq2j2xRi0SvtVPk7ZqPSjUg9r1DTxV5
iXuPjjH6yLrc7djvzME0YOhW5ar4mkfUE0BRJQSTynnPItFvozp8tvnOLyH+PDoJa8tO2LdhifoU
jwM1TTa0lIUkysTCF4xt/GfH6ZXSxCZZDPDT7tfQbxAsFpf04N4UhCuOdI/Bot2bTaW079oubONj
vlJ9Hd3X18wWkwxn0pb93s/sDVHOw4a7ALi/uSDAoGkIVBxU1mN/Vsx7m+ClvWhgdODEDY2EUm1b
U/lEnSj1ykNexbaLfcb8YBwY/X86Aj9SKfWLMvMc9cQqxX5Frnybci0n0zchTabL7kH9YYjZr+ta
Pe9gCblYFrdrQFQZd26O0dZHtB7gMUkg+H//64fEWBOtssTHUPbWQroAwOMuA3i6CYi0+2orBdp2
jak1VNaekHM23LoVUB1o8nDr7MSnHEVx/ytO4j2cKOnDOSB/Xp6Y/TfdoR4pHQcNIMZw4y58i7Ua
SAyOFp0yGeSRYXY9pp2tNbSpKhPPe3w6Iv2ANVguMi9Ud90ZP5t8x1lGsq2KSt4If7a4qErE4tQL
mwag2+NpPqhPEmM7YGTN7mYFnpgNmpRoaV+ew0mZ/f2Wz0UI713+CFzBnCDEx0SdyA8aCiUUjkmo
g8OpP94+Fn7J1YH5w7SsPCGZ3tpcZgUiiYYB6WohLDnXKXjlRhvIHeKr4WtkaImjVNnxUomBsaoS
emF9ZHSOeSRZm2bTLY0KlGt0Dmfi4O/+aSAENcB03rbmlyqFVmQjldikUPpv3nKp6DTjyVDhIS0B
MdfKZHgASKHXBLvXOqExYhDZbkcQvOGCUat8s0AmyDW+5iSKIjn3Ii8Bb7bVIGhg3Xp/Rpqqd/+7
OtYsZs1J9onNGa/bmUOthEPhIYROo3LvmKu6FpzU9OCMftbbFLp9AkBIQnsGqERSR9b19KN4EK/y
0zCkevN5fdkphzpVQ80gojct1t0gvf8ScOTMY0CQ4DF9Y0ubkSUy6nvLNp64rqXGp8hyDOtwmvNX
Qz1krePLARETJ6yddkNKZtCn39LEjTypy3dsQKwKLVIes0SRb67Tuyt0YfVAUHYdX9FPRD1KM5RR
Punj//KhYOAHOhdc8m7nEDU7XOglpLc1eUBtEAje8DQnuy5kHwP78ydkdgEM6Hui81lhWx+tJ4n2
4QGRGXDgCWTQW90iZFsTkeYi4xcVyxYqhQL8YXilvHLbUUJSiPjawqOjGZpu4wC69IAFw/XNWuZo
XNf8cXf0f80wGIHYx/OAD/eXNVodRAc1tzJFvYmmgXXb1OKA59+lrY4HN+6dtPjdnInHW64onTRo
CIHtY/lRU47cgmcYF+Z+4OULvoWFMNsxYOSZ1duFmqh+BnutgkbO5hDEqdyJ3Q8LD3KFNnhUDFWO
JyDPyKL8ITyV5w93JzCx+3cvDp0Aa8lecFm11OK4b2X6oarYfZ7dMRBk3Blvdop4uDDpbjdgSwxs
5/mbDvpCUrnioLkl6fwms5APf7RaeOyHB1gVW+Ape8xW+ZdC5C0gD+jwQVlY5Ypvg2SirAYlydqI
jh3fUebOGEPkVIN8pV9GixB/PyufuM5cJ1Dr4nixYhuGvmxh0nBUSftWttDWTZc7WFo85Z8SX++E
TGmJ/lxMT+rcFSDQKSDbiSlcGyMsUzCwbKk038G0pgpJjbrAdcB7+uaqghGLXowwRzq2UBc9PUE4
fzFw3ED4wgY2lO8p+Hbwlwb3D6npPN2N4EjuwQonFK3+6l3RVT5lOrM4IE/+9fdE5jCCgsoDvh/k
Atf+AnJW9EdkQTqWzH2z231liiPeepJ02USlZk4Rc1/SxEPo9llBzbecKp62Wcr8VFIBbyIxQj4h
LJNa2uEC9J+TRHZNEZXrLhsXSo6IJUc7hZUDPX2uZnAKwOf0e//Djvgt/wZV4DPRqTzEsi9/0QIT
2q+fxc5JSxJyFR03eePv2QQjm0XcaCzWWA4hBKGqkTlw+OSvvPX5EizNqCD3YJbMsv6iAMVDWjsk
VjHc6uLMSQMa4v8qZzgvKxuMQXZ8VaEzq0hwPV2BOl2dGkjBb2lWWu6pYaapDB2eDhw7IH/m1xjz
MC264Q5kMOpOmQh1AHlaasyqBqjACMyamVjO/Dg0CIuV6KhYSOejYx0bygHftRiA1+fPWHCSSprN
IypuFWDavb2HwiOPPGSgnP9DuLcz+qiSGlOBrzeMDaV/9TbFRSITjQ9Q4AFhHcPlm1jNqyCuoWn4
Cu4zgkvYdoYheX+Pv7Recxq4+yU/lJjSfbnTnBdPqh5NPscfn96LJUAL5kKW1fUWYmcpPYTC8Sdf
mpyfXENNDJWGoFcNWrStSi752XjwTEZw/kXo4Ty0vgXtAyzQuoJ61b7Se4wJQ1zEH1MBQLfQNd27
Vn8MKsS7HRebd8ArXFBd+HP3Mtmifyb01d8vGI0u3PW2I+AZGqgzCB7efIO2iS1siNIfO5PfKozT
0pLu9fJsRej7K2QFA3FF/4QmrjBsJEqLB3X/n04RRSSu2viQXwKGXwW/CWykt7xsL62hNXIxJ9B5
M3ECWgm9OrQ9SnMu1qujxCUlaGwttfoVP0oHmIikwpHq3upLmZxlXEvd6vao+LR/r12xWYtpFX7X
os8/aBa3M+L+Qh2ucTI3pNjWIhZSciNMoOHwWYLEWo7rMtdSnL0aFzBkYvRJXqhL4U9KHIzYYk++
mTyvVBQds7cypzIwx+1SGduX1OB9f9e5JcImBqDCf8gvMaCSEHKMIN5bOPL9HVsj4GsqCI6F5Z74
jw9bA+CtskeHFwgyIOHNm/al1WBXAZzRaahZ424T7lI/8xp2ol/izEh8350HhwfhmibiKGV0cneh
m+mLOEsUTuS54Hb+GUoWtJogeWmkiO6AFsWMuJLobVKSyOfRYE+eIeEgIQaedg0QIfWpCMq4dPcX
qIYsSY38uzZrAXVphmJ0jr0kpo3/ZHHtnqmIxIhUVaTnWZiJfHdfEJqrnE4wFbuvlpAQYXf+BQ63
SeK1m4mp9R9AfHlIk2sp96/jy+nK4JZ7veZD4xPnn4GHGxia5mDZWUSSiIb3HWbgB7OFJdzC774X
/kCOEdmBaJdb6E8L/aKeKL8eCgCOXgl+juGPTSKIz5xO1VQ0jnwit4qCCTRH3GtvZZkyyzUUPnoA
Whx9JCdK0+QqgWoqAHdnpdflBv/g7Vabsa2K+T0cmbekkLgzahgLgV7OykmtkitysJL6DFbeczQY
N0vOchizmxX1QFvOjNxf04lSumA/roTLTqWWBV4ikJsjqeIstgYkgiztavcNzDkSwodo39fVePqH
59U2a1LNi5OOJXrTcYbel+5Sfc2z5peav76fmz9c3Aaq/glckrdhnqMVYA2fOqqg3iOdsPnd9l8K
QN5Wmjn5x47GF6psMFAPeFc+anF6bZ8gq/4iYJE9wtQiVMjuFmwMf65tceVzL9uSSq+QLQS8wAG1
X52OakxM0nXRAHfVxABxsrSDDre/ewEmag64ZaipDbjrhCgXNG3i8GED1aF/mEAS6t6AakjUFFma
zuUTr1qaChc9P26oQxTHFtXbQD7eRcMZwHdEN/mCSGwOwwwk8Py86dlU59L9uwcS4Q5Cf4MGRur8
2uoC7tmhAs/aI+tWIrk6YUCOVShvbG0jfyKMdOzpuB4ZRFBQRX62VBBLuUUG5+Bg/M5aaKTp8tlu
WEq/LCg+E2wemqJjELKXuv8uo+u1AO0InANrrwFI45Z87pEyXiJhrF2Yuk82iyvn/HYDj6UxVZ9Z
eLAAMtBVORqGuiMxwEEiIBCKufWPDmZbjC9Xi9kHQfoDh7XGXRdvfuHudkAkpcNNEHS4zOQTnojI
Xv/+ySMViBJuJWBSPISkf9CsFU4LxzYyaqa35UOOyUBjnHb79wiTV+bRFAb/u/SM5aTAWAnscNra
4lDK46OoOLe8Zc996+pJz4LeW76sz99WL+JI6SyvEWxQh22csrLEDKzl6m2c47cXvXzCWoS98Le8
++p/2FuqcX5HtwVxyXaQwoxuYjovWLiZAwXKbVUYz+wk1wt4PlkWeyLZ9t5sT2LYbL3tX7nJ1olo
wgMHoNgmUevB9FTT0fn4YU4fpqLXvimjdiTQ17B09zSjGakaOmOrEaqh/qCOGwDUZPL6yQ/tBsbq
0o1CSxKHhpVQ00ya2E2pV0dOnB8IBayCTGa6fs5lytrjn/52ELJLxgM81HrbJEuxagLKl6H1nhd4
ORRNL3yBrkLEya7vnvC3DfqcuvkrmMpnT734WYVk9TLxVX2zsX5/ebOVrLjrFu29UFxKzuJ6o7k+
UJlEofXniusVW2ek6ySuHDAeqr/482JnahJAeCBS7WBAlWiNgib9jpnnWLTA9/nTCFMbjQFwAMVr
Q3uTi2c833pN4Hpx1XSroY+T1wJ29uwku/XLiN+8c3uf5viK3jFE5RpxZx/Bhb8+Y+BjJm/Mcfu2
H1JFkFynJQlypHcIylyoz5j39c7O+WIRcxPqHbzuUrRncEo43Dy9OVq7LuNOroYTBX7jh9ztgjY3
EP+S5tg4f9NpjeJtfvGixspDyFnIVQBspzMIvHTiEQTvBo0OjQraqb356tBV0rlriI3KULcxogTZ
bMQXhRo4ULLXyCHO4cKE8JrEb4BS/W6RECgUtlSIq+NnIQCDl/+aFMpKTGrc0GeYV2bVO6VAGQGf
pcEIxSD5SkM6MVqasjndNu1YBa7GIvFsU4+M+vCvkymYj/cFg8jlNggcJycYDBCTueanDPJ1LvGJ
yDXtv16Cg3VAjVC0N7MXBSho6s5H0DoOX30kODErPbV9QXxBYtPRKExDbGGdk4X/13ScJX/2glMM
MOyZwfXZ3TjtTcBkYtlsXq1vPlq1dNCCZWJ8+lJmhSfWXpbx4kQ92I+257ly3XjAiPUsLgoGOgBx
UKJlwCp49BwQuG0l+NIAwki5C79Cp1H9gbeVaWZ5b9PhmILxSJCZWuCkE0n8kcZ819UUj/BS0SCz
3bivbK4hXxfwpFQKU4UsNxaI5/uo/TuR+ud4AZytIacMy38VyVOkcDPXXqm+W3srx0IIHxhUFS9+
JBJQIz+CZ/tohEvn0GuMKNJO0JI5xz1THHvc8UTEM0oFGOOK9xbGW9CiLHyhkrOOMoh/oLbBvBI7
Ywi6h8mLJR4GiTx1A83PowxAE5VvmsNmMBaNe0aQqwVFSac+MEhNN1MQM1894RBkXf1YbSB1a1yG
bTIF4tzcH5uVt0KdO4c0i84UptGozQXOi0vjMtA1aMw2LMzs5ZqRL/tAr0V9k31dJ+H5RCNx1MpE
arBwSN1g70IwhYo9A5NLBS0+V8l+H9NjxMEJ6FrQUuRp3XXwlb/s0xvsEBAJqDZsbpWQETMRR83f
7m7d1F3LyuzSEyLYikihNLMM7v7IPxH5db5hWpqBwIDfWuS+a4JXkHg6uf60JPoYEw5Jjqxh7gMl
jxMMUNwVe5L7ZzMGDRUrIJ3dN/Qfof79CumsYsunvJXQPQEL44OzMb7gYXWFnfABfU2DOoHZMx/x
7UkoOGwKhROZQ9TSd0HrvnS4pIuBbZtsVuda6Sz/BiUZLWg8xAN4M/myx+fGw6OnOiZ04fvkV3fO
/2VE+gPxIZIOZotZnlkTQlcLvKossepvQZOaPrbqYLpBqtPQrOEXzy5nFF01LqZrBxzgpYGqioHb
phsppGyoNXBWHMJDfoY0drFb38ohD3QSj/O8exzT19bKgvnRYhNS2BXjFeskCAOUacgFfbJxgNeV
cEevxLF3bVj8eT3DhMSTgX95khY/Xgd3lOeB8/XZjKzGDCGpsXNjHgkXU7PtIZ5gn/qTKGJJMpiP
MSYSbPeBuyj6A+0b7sjYUtZE5s7YYwtbSaLE2uYtX1V0ewNTXv4N6xouFRJoI+x3S00XJP1npfIS
CV//IR/OQUe5L8HkjUIpEZ1xA6j9wtwMCNhNP2wAibLNEM08RL/zYM1XITZu/YG5BNSWCv1xYsTK
hmX1vkauadP0KQXu4rVZ7r43nRPFmdB34TMAvtKtFewDiQnaVlbpx8ITCPhP1zee+9RK/nDWPoF+
LwJZNJGEpU8EJoByPYQk6OSgu3jx8LSjYvaOjRinTNos8C7alUhCAVnI8dArb63jbe45KXKkcF26
U2dUpmE+oX/NvlG//zGVHltTBtZUYmtra0lJcPqb+s8SdQogcQtXzTjhO07/+HwqNLEm5vuCFh1+
0eAxht/A4rJhUO3rNjbH3C/ljpyfpSZclquuJvJcBy39gry29LXP6P16q5X4aMDIFmkCWL2bCEPu
6FAQi412bd0ZWgCkh6UIlMrCNo/bA80NU+RkIZ1BU7w9TmbtFBO/CIzhE5Bhe0BOoD/OZH9RBI99
F4ISB+qpeB6U4+HuWRnWFRThJcY/TMCi4kGM6LSwkUvkw5ogzWwSfkyz05oEk3qoLty3DK2vq9pH
3mtH4rJgBchQx//H4gEYGBZdwkulEyaycW6pUv+9sfCCUpjiBT3t6sfMo5hmzy2VxnNJFbNapA+V
FGV6jpu6hv9Xmbe94QKoUY6ikaTRE7X+RqijI/zxfFZBEwA+jfaaRjzIQ7qoblnOU/zZkSjzK8vJ
tJxWG/qIhhL4S+Qnbn/pVtdQsY9FpyMkLme212b7zXJnF2l2VPC+DxF0tYK/Kbm/iK6RhO5lKw/e
+tvLmn4FMUJCxVe/KxA682j/RzZxxxWaUncit6C76nvG7iXHRhJUS4jnykyHZR7buaTrwmP6Mo8J
skuUeI/Ilxg4F4cHdIwtl74guVRBS/4ZyliqpqkyMP5MCZoXfh/RVN8zM+6ws83RHdPDxqq5nq5C
2ddppJHG2B4yy/vhbtuAPyX8VcM+UDSwzU7zA2auYE2w8RCWKaxfLELbWyGR48azt5AgWdc5YOvq
2dysPB0MZftBaodPbylFwgKe8xe8r4CIvjKg7l7mtKmL4dzNpFnkSXbPJWFOa8Xe+qgDbALxrdBK
stqFF2EgVVpcyLiF6deJtDqprN1zjlfGp276nUzH49zslx1HuTRDZtBg90XjeNrJxRxXa9u3kwEV
8QAlvWC9lC7qWfcL0ZZFJpt9UViUBoYBaLRMeAc4aeqcwF6fyEpkFQbhWqLo0Jxk9VQkoncnaaqV
HZt5bVX3pD7Bno+vgrh9ul32sdkyl4ZnbewMLcHd2x9j4n3BgkQDBzMVVU8GaEC7WHHXAP2gjK2r
xwib4dNPoNvK9V3Yl3K8AYnHTAuvQwfMYe77L+0MZ6MtqVdf3lgOFR4f9ek/1iyLexizpLXk4ovQ
wGEJULLK6nITyQYT3dmqE5RR7r3bnHFlMA2A4CysoDpcQvNNhrs3MtPvhyvQKjfILtpx5BK5k7Ht
SYYx6Xdw9Ob6jZKqnShNKmQaibT7RfMmaxAk2XpeFciPFTqqp0FQ8Icnzw9H5hh+M1Fasy+k1zEc
GfsYo7wgsZ5zLv+Y+WhGK5gYuhYNturwrDp4I+pF9OSAec+hzfJx/+utoTlJJctMfach9v3zbjlf
60cpllyGtnd15HOfHdlXKjML+3Ws1S2TvLNlvC97CVaebFQYFv3rV0h9AUyXWdS6S7c4TU69n4jJ
8KL2TB2tNAtqnPFaU2FLxOgwApqrR0age+kHur9lE5KZm2ztpg2Xxa8Ee9fwwn3mmE7pYbhZRKEN
Gukcr6Pyvoj+4ZqMgGC4o0khcNFQZTStfP9jMet4ff+YqznAf7rF7rjqvnlCFsTobD4VZqbxurUe
z7SxTdbAghrUSY0kTmFFU5Lno9Hlrbl3kDrN/TzwrDSKv/IudS34MuQAs9U9hOPsmS6KgPtqOSct
/rg4l1Bl0dAUJJN4ADSJhQ0siclYLnZcFi0+SPplfK+skilyEpYLzhZdK/AKBI30Cv63R7Ou2ZN2
eFnkL98MXVUeEyuAOtgUJMrpjAu4lIpPopNK3Cwps1CxwkuC0xAPDY9+x1IHeatnQPtRBdkgmW7t
9jTuIPvnOm76w39BGmiBxMB+tO/xeXm+UEBLRkjNpWR+BH9w8sC5ekdZcwy1c4K8hUk6iO37lu4C
OhZzn4iAKFzGIuY+k5tgLU5lbl7yHc2GVKpOF1VT8QYwgmGJRlfob43XCP15gGRA4e6b4VR5P1Fc
d6NvTqBTbRf3SmKa5/wdz3p5jsLHr33fcvcEZLte6hsbWo6LzD44hWO+VYJdQ9vew/DsZyuwnusE
V/to1/8k4wdZCg7UpEzq/4WOnT2ldcWU0xRZFLorRfLWgteYmoPmKGVJ1ICSqWm70ZbouEzv7eZq
CWQcw7WeXgIsqsKpSPvZqqTLcJUUbX+McJ8Jw5oNkAcG3/Y162zNHTJtzW/Vr1rL92UzcS/Kxt1z
RLuFvMWLCBy5Hd3L1ORdTAIZIBkjzVbx0fd/hObqOOeFI1sKuEORrWpD9CQoslnZsBlL3L05M5pG
R+yulDAMjAE9Lxp3vEsdUfenTb78j+Cjzy7OTKPy37AKPTL/5RL0XwfqmAarC6xwhDmbsRurTiUK
L87SgY/D0eFNzsTRvvt9M8X7Soivne7esoC94sA5HMWw+bx91EbXjoftn9MISJyWrWVDE66fpWEw
c9WreIxDn+zg1sS9He7RLsc3RxGNFjVcxiyWsqjYPolzCIJEo3QmVNFAqKuUAVhOYEv5HBPUXVRS
m52yI8EHFlmOCpMc1DYPDcUE6DbmV2Ccmvq+24W3L0VdlyKz7jadk5EHq/tJBH5Mre0wFHk3uuN6
nSyQMYaENoxPoB4C9hjJHxUdpJxu3ejNX0u2AAnL6rvNKB+PbEzb22F+vGMHqwPrIWViaVQw8ARq
g/v9D2+H7+5I8+gWCv6edzQ/79CX4Zi6cL89EB+ZU8k2G+b7FeDLGpOdoYNgzNmSlt8MV4PHA0Qe
LH7EXtq4l8b6v2D3DzfY2rBQiDyzsHeAcMtmr2uQrG+AdjqIMpNrR6iQ7eGgbfQMlNJDAEcHY/V7
v2rQKMCZNrO+a33QkAXW3YYngO1VJwM4XipxHWL3U1DG76gUzBT5qWj6wrEsQNfNyYhG7kGBQ4mq
GVR22AWjXtTtKT8+yssktP+esrvQV9I8ga9P9XoPMZYyq/U/BekqVt/M1FyEAmugxY3XdbYDMcUb
WShl3BAW/7Rz4sQ1tsrN8eEf35SiI245xb98z6zR4+4riMYrbIBVQUR0BTjnAygUbWOFORchjHAY
ABeDr84Afki40X7G1gAaj3kbGqddvPrGuN8xLkQiTId14VKHdQSXNCpF/0fSJP+eP84O35STJZM5
/qq6pxMMwLbWbHjln7YTmLPEMdi9i5P0EMR6akj3juzvQ8hpZij3lQBFZWNG5AZC7pYfA1TRCTI1
0lPVM3fbN1RTi6OrOicHftq8xqtz4VhkuIbNx2FzbAlziBAZv80HfaKC6cbHXNEM5teG69SURp3s
CSquOe/5uRPWUIJ/ENTKcYpQxCRBUEKojHWLQvaUxoNCOxeDreHB3BX6dSiHBpQ5on5Lsv821OB8
xYkedcHWiGwONPoFS4uFKxxfYFV58vSmz6hRdfhPGIlhm33RFTUHDvguADj6ozOTeE5zxKhclv7h
JxJHDyJ4yIOYa0EzvA5Ohle1b9JDOAUyj6MPHzqrTAH5PGJz9AF+XgYUcRevt0lUo3qMm/FStUv7
z2HRtYrTfijAvhPNM3UTmqJu/TLSW5F3y55y3z6W7sB1qh9PhxCIhoYkHEWHIxIY2hJTqZXf955H
EvO5bqH6+JezEg/RoTxbQuL98prq25zrwLIcSVRYn/pk2223Eqd/C7mZx7UG/jYTygR4op3vbVp6
jvXneXa6mFg8Uc2o7/HUFwCk1aJt6IEr0v+h8kqXrXCQ16K5bBRgEe9ihiDegE2qbpm+djrfZ0uI
2ul0M+x3G4N9cv/q9F399Q8Pb9jG9Wk6Jq25p+cs6bH9k6aX5cWBECMORBwtrzx4HuO06HsaiGTs
DaLFgkrpyX1Khy0Gl47DdsY2EM3fPUYoBLnCfRuKMlaFhk58KDgHeZCmH4LerSvlCsHa5d5f1bxi
os1SGClDEw23HcmXSXMoUPyKuDzS00JoscQ4FzUsLIdZiXSNhFd+FaZpUn0A5njzDSJgxy6bv7Dp
OcW1I66YjZzNGcNzxzVZjxx1PT3sjayL6Icwf87LlPBnm2LXXZy5foR2JuatVmAqKXc4IArA8hzL
Q9M+Qq13t41byjZofiOXIvdb0mpBWETa8m8n7cNTuJtLp/kPgj7Veziwr/STSVso2TaVLPNzuam2
E2bl+PLF3bYveLVgmW0Mu99R3qlFmnBuDEyjMoGfLSlz2QAL3szXXlYqF2M1Ds6yHBKXQQ5CS9Yp
p33vTHYFztMWZ0yrcucwnnlqfQuw7j6F8X5vv4/OdZU6Uw3j1kBVNcyhJlSpYjkxA+JP/o4ogc+u
3yJuNpXOq28qbK7E0W4Rs8tp5+oAFqyM/1tQ0dFq4nL6cpCYnEI1kBnBFemTKzFOFT6T7xPOhe0u
n8rd8J3rIn9x89ZK0icUnhIEtLCN9f4TBEtmG+kOfd8sVZ3g2Dt6SYd0/rSNx3jUIVqJnUhgmuMU
SfVSr1QtdFCUpVh0yKCBsMIW3Vsm/KsGHWkJa5558sOrVvfaK41nqiKcQcpbx3PgNKY5yxtoZVOD
uM4XXtSGK8sXcKWQbZRCrVAZ2uacw80mfKKWdMzNeE9MjrbHNi+2ACjyDpZTX2mFP/bpeHHo8kfQ
mtu3dDrI5aFO6XLSQ3SJH3cQnHh/+gPzAyeNU/vFQEgs5dlMHJDHPssslkJjqby8f23Qxdydy1F3
a1RhzdXINXpiVjVwlL2LpAeuJYKouQPmma9AuN0bhgCjUyrp4BYWJw6TusB47/QUxSo0YDlSBK76
9O0n2wU6oN11OZz1NPErPSdwPdAWyElTcQp9s+oFraJS2VzCd+P31n71V0yAraKQnrKPWQF0uaLY
Nnn06nfHANmtl4dNesnn3T7Crm4eV/j7g1YHyIGVv/iNQYgBlarNVn5jlQq3dLnx7tOh8zGlIE2y
TUxqSCOjNdSJK63L1Kls80qxBlIShLUPYE8uBv2vIW3mLvRD9cXe36+JQ0FY/paebiIwFXHBgChC
F3EsKaySmcQJ1kZKJL4GjVu1bZmYRIVu/JWHBg/hQSfb8bSx9QmutLWNl75PxS/ZWx4kE1SChIBH
8mu+DVxyjUbMVRh5uUSRFlA7yldDMZeh+kTiBe4dGgDYLVJ42De9+tsxQJBSjhlqWm9uGb+tkn0G
JFoxmZAOxZjDB4zGFTPrpvnxuRTozVA4gZK74gEt7ktyHqaxjCH4iJC2d07J+jrD6dH651k8Xl46
anOzjaaKFHCl+A0EBMXei7JQjDUNDKHR4xiyrCcahia6sTLaGv8GfIvkisIu9SatryyUwcazYeE0
kHKlx1jv/Ykm1tP8Ys+VngYkKWfJ4OHfZnPo5tyAkRaRT9RnbA9rCEiWPis6O+NYQzo/lcTJrhF7
yBjqtNNCqh4og+wbE+G9Gdjkno5w/gZQa0ZAi60I5P9td+rwTEnXAu/UQwvXhv+n0XoJnVTwRqtC
+h5JHPKvD28ugxm7kentfpAsTTzrreAneOk3tpWx3jtloo3cN1NQp/mrw/YHPeqFO5aLhUy8RPsD
xHVkVUVILjBly6IrNkx/LasA8I91ehwRIsLehfAIv5+hiwFcziPia5ePtsghJLMZljvqe0L5t8VR
Zi17hG8dJNzxvdinNSzX9vekskxGxvRdb25MWQHeUcxGJAGoFprL65iHnXpYMDxrm/uU21bc9ndo
MtvpW3iMNOuSslNTsrmAdYfi+x/iKU7xKZ5s1WiDJEXKG+EWS2l83V6RS775MmCqZSc8WiGpMww6
SlDlsNnIKsc6LKR7CVoxmO3svRfRrTj6OBF0K4GT+GmGpziKzX39XEZouH7O+zw/Rh3gbNDa7KY2
TyBIPeOH2xP9U2sjqPLsxQk0RTXz03wiUusz02qcJG0Y3gTLT/OdfTtynH0XZDTjP0/6/xenDL+F
/Xzbmgy3KvGh6u41AACFV5OO8YNkVQQ7vZOCcT0rjQzyn/nb8FixQbkA05B2zFY+pb0UzTPCL3EX
jgdqU8mv1TpqXs8zJ12DtGS4NVIOPggaTbnONbhCd08zwbbaDxqNIuU5jk8U2XXDOIYwDQdTPBv3
U2MJff/r+8mv9WNHbWTjTiPFC1jiva2QkWvcNHm7tme8SFizurNrijLEodd3aRXOIpUpsxExp/8E
bb9f7bAVojFdyNV0g1IMmdu+qrMsRpE95pWQhyI1cp9Vlrs83MvQLZSrdQvqYKtgW7oQUudpgiAD
HUADBG4uATKehYj/nXm6U4SSgZZJb7YMn1C4Q5iCkhwPWcZQ3B87uIyNW5+DZqVvpafYIiOU1Tin
URAvZba9IUi15Kangcb0LB8LLzFVvYIIhfhPDObp06yFpCCWTUzCWqO52XfGzdxkxFsWfMrVvexx
I2+BYJBxzV5ra331T0h/vx3mex7VVb+VCMNMGlni89slHtToUU5pKqkY36pJTUjKguNAicyuu8a+
VKn/1iv8gg8uLXtsavL6/EsJfNio6MoD2aNQTZgIJ7eNLkr87slO4R/hmUL/nI5kBqcNW2kscTCz
LVrf4QQvSWl/rfbGSe+bEzmPiJbtswdiW4y5d3XucWbGnnA2rf5CXccXacDEL7fQ5jsElNhCeTEu
f3QsAn2CPTyr9zjOJzAPDcpnH/BY33t6jfH/tqBmYT0GDP9rrbkv2zXip5TXcR8Zc9MtcHn5YnKl
C2rmWWAJJ+0Y6k0ghIw+glXf4bedDikhCYgQ+Y4qhlAnsSIpZqpIj+vGvaQIhPvWkP9XNCOpoUgN
zTlblkF79gPyDzdy+fxm2F7XP1sJUeLuidIEE7aO0BEbfpzfyQDD3T8dSqwH/NAnXCL/9ZlGpmZc
h3A2NnA2DaSml+9SkBKBXP/w5WfTU5mrQZD11ejLkWR5yz2RNmZ5sZkM5CG7KuRK9k7eEb5etXYD
D3nn8TTynHV1Itd93Awea5zqBh4GnIKtF8q59lM3ojimQSIuqNvibIksMmhTvj/qUmnOQw8d949M
WpfFpVttqQQWhI/IJbaCHiOluaZugShcMz/SLuoHAAHxtyITNAiYNSftG2FxyVQi0gl2XHxK3G40
EuF/mRXotequojeXM4sp7jwhvz2c41Va1prXbLyi2/a+4oPUtqzIs7dFE51ExsptyLrIKf42LI6E
ghLDKwTpqyLPdr+gCmRwK0PnHTO8FJOzh0oOl9fp8cv7dcbwtnTgcOur3a9A7YwrP1jklCJBGUkW
9xi+hm11NXX5SpxF2zpOgCmrytmJHkWi7VHUTo1sOH5XimaUVEPykKth7dmmclQYHtaZi5XG1hB6
QzdCoKaDMzmbF7uN4lPTUxwigWpGbMk0Vot4FSun06EOVSFtedZT49u3GxfJPFHeqM2XgYDcW9FC
WkRkr2SeVsiVzppn1KCBgxQWcnacu7MYhdtdwpXFxj8HWE3jn6aA1mOCPreuO/q4ELXJqfMb6kY1
Gy94WM0XgDY/EZyczgZRa24BBhZGwxo73cN6zLcl1uDCMaX0fzbDs7qBlOQdkzpUPKQQd5Ir52qd
6FbiwVrtMYklMhzcTHarHpp3k00SwR7xolL4IERVbQUBll1GCclnX1H7sKSK+CnwcZiyp0ODiovS
4mVXKM1J8jvSF+32pdq0zYrJVNWbUcFo3IIBneMEnGXs6Xc0gG6UzxfbKeSdRgxi3BnDO46uGZWt
F2eDbmf1i/817gDQfBNQ4OhlDqYcRrKZajDAOgW1kx2NMfetmjUD5NhnaHkwuZ5goytYR5KryjbE
tQyO9jvRNewuggYnnpXIT3AXOqQ/xh0ZjNGwkK4LkztMltlqbpxGH3tpV84Af+yy9M360yGVPnRw
cbEsI7hcPA266ZIBOigWGBE9yrnMvmp73ZazetpQetzPAx8IJQCaPed2+Qr0nXueulyueVQJtdSf
ye4m3cfo0/J5k2Voal1JwziEiFf7TdH5N2963aFToRlJgCzGM54YThUy3Bt7Lmj3ehKQvs+gTsRM
Kzd1NqyjmiOZBmdab2iT8XEQa8cc4hvGDYeFMFgKbcTDhzn87T15EfG5caiORw8f//xnkQMnaMxB
2SIV8ZCLxr1wunxf5VKCWRtCBRdc4AJCyLhSv3HrKyR702xDbujmhHtDadx2P17823eXkYlYFN39
b2gIwr0aq105cm/c7oUARsM2qGEhCMJuDO8hofC0C5b5cgY5BSU3cPKVOE1/5YOtIW2Ru2aNhCee
2N2EgnDWK9CtEmbrBfGSTR9K2+sydgw/BEFPqlixeVll358lDvak8JUcjrxvXL1qJbaiZGpl/9Hp
XwpVWGqkldovrXnhsl51DenWADzXt8VmaIRAQFUyJODKlBghttYGtyd+VgScQKlUOMC/aW88n4u9
lSGzgGH2g+Y9+gancjZ4/2cRAKv5KQAgBRnDoBfZuA6J3pj3mOfoudx+j2fUIVsC6oQXtV7wUOpf
QS6L0jiqsKFys27e/z/m3cfZbcWeSr6r2kusvUnplHOhXp2+QjyVUtzYoHo0MZiz3ysj+W+pa479
BxVH+KU7efR9yNKpP2LFBXPHYQO1odxKDJbo66hDr3XBoUe1SVQYDWty35eIlbM3pRIXZ0kthobV
e3frHoeikby7JfjW0ymUjBp+LFajNpysKORfLZ2qk/x0TvK5iDYEOCqFoO3Y01MV9P8BefhDBQZD
onJ8pOW4mi60vKNDwQVE8/HyXTS3krhhcD3IkbCr/0sdiXdSr2B6RNA7Dq+F8cdSEoRUh286WeKA
gkEBopUrnWWfvFUC8Fn5sMRlVXtFPzVQcHI2cVqsTrax4nLBEuKKrYUsP13NO/vCxN0fGDpakbTY
maxh67VziuDrE5oCoeAr+GnwuBIggDIgurWItWwz+LFhq8S4Ic4VtJUPWv6R6oQ3/s3/K7mFTK22
J1plmO8h+xKldyIwMuySMAoUdUKNShXNoc9+arJDAOYuHBIHDLSU6doeBlCSmLWVsmW8UAMmhL3h
UER6hOTXJHqsvj7qdrlszHnKhIgQ5Ltd25zOJn7QaAl8Gijs090P+SHpRf/sedAARwJ9VKYsYUNG
P4PWPkZtgyAB50G9wiDv3es7SiLQ7mpO1/jRaK9gclKUgvTkMejRjI/mA0+bM+MYBFii/sEJUjUq
FXJc/O9l/k9ag9lBEGQon72eNSUbK+Kl1bPQbJtaJNKYyy83/yxOyEIYF8Sfgc6I0B4wOzTVT+bo
j0pQ00jIiyGkiZ+b7R3GE8ELHpT+GF7kj/36FAGnBwGdPN9lzBUko61c8dXBpaf1rAwehWgER3EB
PZ4Y6U88HH9zaHVcBkskO1WxwvA/JmvJWr1CxAgbmbca/PJNqtSuC0epxpYF2M0Zn784VE7YYM54
IicvxvvFj3GzsLFYisfw/KkdJPdk2X8BiaNFm6fFdX6rJuga1ykTRzaREhESUmzOY6mx5iuDFKe8
sfgQT2aAyNVStZss80y3C03G91XmdVadKGRRHbp9cdI+ylQfrhp44zbNY9hM5Y1BksIjrpElQCwR
NKz0BzMqBnXN4W8REB+v5ce6CkDLqkgUe+mcu3S7p9+Sw2KXTfcV85Xv1h2VmbJP60dmIVgKhhnp
Ua/6sXsbuqhVdVSpbrEw7kddmFOLW78dlI+3ANXW4cDoTn+eAveEhB9VFS25UCyf+I3ohe8xMLym
C8RSmz4B5eue8QczCOkb8vkxpnMu8FbU8RCEfPI5CAv3zFLRYOCWptF5/XAU/4x6DmzWMw1zkTha
ds4zDMSMd6KSQqLbTcMfILQeaFw/pHBu9+NUBnaoplVVWK42aA+6txAfoDJoTSa2+BpUqaLw2v7s
R8JLtG82PGF97uWjtxMgaHDU1qyrlA7MA02PIHpNhGAU8taEaVKGRVbcnuRLqnpC31CdCmLpwl3p
G3fjO/kmgdM26eY+zQW9euWqEEkJw55kjBLH8m8P5nAighz3ZhKayz3FFwNOzYZDeSNOUu3FFsp0
YFQq6JFnng0wXHhKEMERvVHAWbgYFNLkVhZTb2cqBsd7ersjOWc7Uag+xuFvkWu3Wuu7hCZ3QXEO
S/KOs1/tWKnNBiyjHxAXFvZa4TUTohNRGVSUydGEVhi5lPl/KYQ/jwlWm+Q+k1zkXqmg4XUUiG86
mWiEm0ZOoq5O6jR5LAuafviOa2vZfmRGgvZN+J8gKQS8Fz936OzMpd3qiFON+3Cdxkp3Not0Z6ar
aDfdG0/a8gUlZN7FRb9DSKTbpT8gC4PYv6+yrgx/vZ8Nl1WKkTIkO5FPj4Gaonrr698G1gbSSYhl
WFbTPTnI8r4hbztwhgclLSXXvA8Cz9nlriQ82qA1sU2KUUqgPRNQ6wXxs1q+wmL36WcRwxE9BRlp
emI0CwM/nXWOOhVnDX6xivL0Sf/SZpEmXSgDBHZ1VgQ+QBKksDhKH54/QvlHzjVg/qUZ4Gp7+1vm
7+ryYTuGUsWh07bpIxdVHynylLJYXIiCF+pCC0Eg181jA/+2WvNa9Zsbxw3qKJKx2eKheg4wgOTF
2TPbE7p3b3rdHrDDms5D22tC9i+xIALCGLNh26YXlpA6OUHfqvJYQdYznn8GruOlt/3rIQw9+WJw
9L5QKgdFGoodKGhjo+4VLpJTtbhJeWQ1NCRz2wKYp7z/aKNQ3YtFeQm16RVCThe1vpeVr2ZeHLAv
QAxplcaSvIMwmbIXDWnsvb9Gi3J2cBjOGG90ttAZTFaI+xAQFA6O1LDl4PhBGpoeRWa0FDWc9Zvz
CN680N+X5dd3sgCIWZrzYQzUn4+dG89+3PIF3WnO0zsmfcGsfBaCTVLNO5r/iUb9Y2bLg4UFSbq7
D8WumaIrNeyMhedGQWt7uN0+ovy2pqfj3r9tfnvPBzZEmhiuaO5EQQbeFXWo1g/ctlwrheDeSfnt
f9uPkgapGug8jb4KAskcrd5ZRudjoYhAU3RBeucl7T66x+xStmfXImxDjkTrVNkRl4jcEJFIE9vI
kPdrUVgEm2mm4C+YGfBudXC0VdnN2n9HF2s02x3ptDcZTMiRKpzhqI2YRIU3DMLS/qEkJ4I3DST3
FYNtSSK/rK7V7lWxMa0eYr3MU/c8dHAdttnRD00nzEAzlMALv527wp5X5rCj/Kqqkf7amaF4xUqA
zkVoHy2jxcnDrn9/mVUsVfOZqJafC+ZG024Yu7DstJlTL2xiYeP0dVxHIYmyH2ECcPhkrD8/6awJ
/3okke+B6A4gsVEPjTr272L64OhE0KBtCia3OkgMkyRQH4HHaQpwFclWyQo473LkcxbHWhDZeRYe
TbHsVl7NCnQfwgd7Jc6Ua/zZHpzeNOoHgLL325PDT16ibDkS63mFM7N26RhMk0ICEljY6s/hv8cR
tNCQZVplNPTUmuxqX0JBtutX6jenvcP69tW2aVxTXoRXTAAv6W5mq7UVQWohQDvRN+FV6ZfK9L0X
1i8+9zDgudqHq4Ht1/iK9ucAemgOE6rVJL1Azmfm8ztn4Jqih48sIDnKHAryGSX96HLJzLLkemBz
VgawNNphL0/pg7dENFu4boGX1+W1abgcronOJlGkRa6SaGpkhZt3CCqinVVTyYadEpNlBVdL4HUN
92M0CuXZ5EvzGh3lkkVUHzGs5joHv8YU78H5oEc6XrXAPhdImXn3bscDDp3IROijiEuyOeUUo1hg
xnPvMwqCvoWWf64sZLofIrQ0UNMjryNmfim5AD2h2oC3GdV+6MmJeYfSTZ+u2AymFxlJv5RVNzwQ
uu2vUf+VkyRN+fJuCKKHyv9Px2Rz7Eg8odU3U3o8xQdQkscBTTsWhZ1Fd/vkf0ycH2Qhwzk0K5Y0
XkrWNJJAmo/bG4XG7ZSnbxiWqj1UIHKueaSE+uLAXL0uuHpu5UEopF6uUrjsuyiRr+qudv1dv0jE
eQBJE3yWSA0hqE2EzZOLWgWeAcxS3EegLlQRjeBE/x6Qh1y8bKiYIKQ88AG8/BSOLCyFQKavvsSz
SW2PtjlwnQllC1eBa4vCw1j2PvKFsixTQqsrcVPY1ZikljqA2FiXgbML4UhwQ7jOr9gds0bk6R13
Z6omlK4UbyGUx+WifICjIFIMoSQQ9XGjxFr7RxNLf8OzaG4c/ubDnjrCN/D+8RPg7ZmCRVXYcWlk
4JTaK5si1UqeoEjD9luJ/W4kgrSlqe0+qgbcHFevMM3Cq2SRPXh8ppr6dbbSLn6sw+Z2vAvMynL6
iE0WSrhN9vK/M1RDf5EeWDAvZ/LDSUcH2RmuNTBJTrHBnBwkgzlvptEJNneJjnpLNCzeWxlGhyCy
0R/Wc3QFzfXG9xx2HT7Mp+GJKZc4s26xWimLeT09LdU6uyRmPlSNLjvmXpctQa5A2jDUhx/4f5ic
DjvQD2O2FMTgWaBrKvF7grLtUGMA5qN5xCKuRjRzOEPFNew58zdW/V3JYG1tbQUzvkqe/mwH0zqc
+zBL60Rjp98fziMwVuVfs9eC13RjBmW0Nm+yQAcL8ToI1pxzhAUhFWFjeGm3TC/k5zWF9i3jLaMx
6dZ91TVoNMAvEdtXhklr38X9gLYNEWBXOL6rFHGeoiTTIPlNh4y+dkO5lUujVmRN/qRztJO3R/BS
YUI493zFQrYLZGS+91n31+7N1Kf+o7P0XhrQWEqPG83DHTQPOuBQ0SgRM9lWKzJQvB0rOBaZioao
xRwZt9C3OuuqqeVnxR8PxHHo1TruAR/uA4/q4mc6vJzOzlsxgW4ZDxY124m9MrlnWtiRbvXGY5Xk
p1n0OlP5Pm014/EZuclpJxzMPM4/fHmei+HZnCyY1ummQsLlg0kwOIwFpPbtgcg2oLQEB2JvtSEG
n8OeqszEjN7tfS0N+Vat+9P+Ip/M67OP5VXI6XPvOXnB1l5CR7PcXaW0oBTO+NPRSybnvE7QKpIc
cmQigLH4uIGEFG1ousVY5ilKTlimr8A2y5rd5wZ/5uMAc+M7cFpt6z8AmJKoRGfHEIKFc8Har2SQ
5RkkllyVZ6kyLD7iqLD8+4aXsgqP4PPzqohvPGHsnLz4uD3NodFBJ464G2naq4S1Z1NBDJBSxenr
RhQ8UvGoi2qIEP/EttOGNwl6FJVahazAFVGjxLrZwPSvlaZDBNCLV/HeQPTrtiZjyt02q3KZMO1B
BajNsgvs1QXhTsiKALfQLF2q8YeNUbN/u0kds5qOT365lApl3p0hgzypWvjSeZ8HAwEilvb4EBp3
hH3+BjLUQUbjEXwiJtbRZHe2Ep9Y2brnqbX9MeQ7oooRZy6Z66KNR6dPzXaEP19wRR11IPeXdPNc
ESzKN8o+HCjFiUBIejtsiFRgbN1BbyHe3DAz4tgAwFjCkADZ5NsNqVVDp0aoaHDmxM0ZwTfrp8gY
HID101Im4r48BU73n35s33Wo+yJpfRam1CR1u1x/VvBDmGkyTiUbCiT9+msKCOezLRUFWIzyvNe+
lZAxkJ1MwfNxMoh1tKGqM5No+yN/hgp8/LHPvxrtbSXg6b4X8nf4b7sbUhIh5yhxqoGxg6NNVsur
6xS15ntpywTTDzkx3sgW/muEednEJOxulXcNgqA+eD/GTGJMMZdfmg73yI/i9+39vwQSX6ShgmEW
tmgfz8K4zCd1LJkRgK6M2rH7Sl9IYGnN8YPu5SBAarQrborAGPK5Gf/YB2/xeJ3hIQ6IsnnhohsK
aralxBx1K2d2bvF0IL5yAl7j+OJVNXT0DgXGTOYSuzhNsUfkiKps/v+ve75vqfqp/dr9TRas6aji
Z1mT4afRGpU7VxBGXtRHoqz/lLuNoXF9B3EsWu3unlva2UtsbF9fOIhdncH4yiZVUrOhR+aOmDpQ
6CYpgsJ0fTa+2vpv58F4RSd46Cj09YAWTUYwtWrbUS++JB4pb16BNYMD/nS4/i11kRYQtdJtFHVb
lOZ18G/QT3fordRlTmbod8Iu4woBr3V3M1J0uaICFa62WPPlDlLLSTwHt3hTblbN2UoQdyVY1QFv
HE7sjL8uXRcpqhgBOwzmCctwHg4SXQ6hPEyIdA3TCTsSlhN0KZYj/3LbV+AI0yEsN4008nvQAWUT
qPraFd0j32DT0JFaaejVqjpSEyw0qiVNKaUaE4XpHYM39bLQXXO5dIyt9fG/UEhw2q3hZRCTnM52
HdxUYk8E9J7nLCkSQLKSL7/OVxnjbv8YC42m/VISf32PyCqraIm7ZaZpcv6GtEal7FkWlZowCwe+
iPJqmuiyq5s/P0UczkTCP7qjGYSbnGEO4IR06YNpwkT+bJvqEZIMA5NNvLBgCuOGnTv11cSjnDXL
oHOmyn6Lw7n4RFaEMLTQQl4XtJ/nXpEPOMMrLYDQXg80wI362OlBULuMBbA1kPwQyo3sldpORVdB
c+sh8DoYGJ/IL3gsASCkgqobCnELPXF2mIVEPhiUWtw9LbpbRDYYccUjHcDg7kr4ER3edaROkR6S
LyIMt8Xwa4/PF13ebRpz17wNi4xsN87maXXrNx1J7e9t2mSL0p51dsQ7pnZFI5WG+nqp/pfYYxRO
vnZrJvrNUmmsk5d+xEw0p6SYf5ydXPILmwF6xWd5rIDSzIqmHuhJ+in/fNpYCblsxZmz0DrNwxUp
/BcBkhS03k1q+3YuWJBNTURjD6Vu2W+hSfXCrJi93tVZtYX0bj52IPG5LvByUlkymEEn5WOXIYKH
UaK66fPeYXVY+xjJdFdSBuNXeQhev5JEH0Sybvm+jVMG2qLqjzGWin7AoXlwZCL6CppVIbrf/qq3
mhOyU4czvvhtHq7PzUyAqkvgT1vXyOT4yE7gBxiFKuStoXFB7wifF1fDc9M0eoCxgvRGzvVl5GBN
jp0apsDc29wkAFQyLLhDfFsfyl2BuQHWGhUum1SEq0tSE2wHh3sydd6qwosXn/SMFU/3ugMpcGer
Z3J9P3ZLzLN6Cg6o/ELegEbvTAhgyfVPcbUy/0WXa28HkypQs0y72mjxgUW+AkHq5WMAwsy/uGzp
69orO2XtVD58Bpg8b9GMj0xBgMbNImTtC7XMw9PDpdF+U6dcYmjcHZNfJEzecsbdlXS3YWpYBGav
B8RjzorEPowEDZebu35B3qXKYw6pyL2ONc0mH7wZ9vM2OqqkoLPLkpbmGXU59hBjQlCYt9HTLS2D
3StQsqpvdJ2qNJJNUA51WDiZ4AKFJAZs3vo9qiYomlQH7RjoQuYzgbqYmLuQxWZCXO2c0jNFd++c
XV5FjnETeI4CR+qU0KiSWhTe1aoUn11VeUqkaBWBc90GQRpfbLHiOid7os8uULpUmfEHqcNcLfpA
mOWZvdFZZB185sRuOsAJ1FXovf5vsISd0f8hXAnWMYyYVU+jM9TDRpyz0VEY7YzCGgqv+5SudjVa
RQARBetoEDkW/aQoWwKb6lAWaFHeKRF0XmdC2GywTsO86CFEKbMQ2nm8c3KlFxicCL3t4V7Ycyyo
g3SaEWSYcE6IeVW5FFGhlVwrjUhA8SIBACpje8jIKZf1oTmuuf9uWTiVcdMXKFZSwcTTS9Xfm8Kp
8j96DsLnHMaxzpILp2rkQGV66RY7bw6D6k4S8kriPImZftfrKabBFEjl8Cwn5XAqwxvyPUsbb7sB
5No65psyA6dqx3Mwrycdzux1hOjjj5B1jHwPRa7Gt8lrAPlPFvpPIKv+NMxTZ6tnctwQkIPHAsXb
ihbS0PzxgAlq6MQ7m1d5zADu7tQ1npsRghFYvApzJ29P8f5jewPIva4B8/xBo+Yz0IAntHMQmwqK
4ewMeolqpXUxc7ne1X9srhI2/npeK/Accf2yH4sbBD/zVglWqK6dodCOTQlKLC42PM+dju54CKK6
SQMTDlORGqP9et6vALe6o8Nzf9ruJIAqpjJI84ay1Xjcv9+J5D+stMI2MkEpFwCZWb7Fn26WzGDC
Cw0Wxf5krCcEKAimqGock61W9gFafwl+gxJa6zTT7nZEMbYRr0clZxjgiHHEN4to0HmbUFQxP/EL
hV4c0j38J5Bu6tLzaDOdUdbTFwzcmuUpQFMGDOnSck9Fsh34D2qAXrz43+DA7eiUW5FMPZZUaaij
ThLliOjWkP6cDOYenfA6radDp8dJeHhyneUK6cS21n5YbPJGslWomaHC84LcUJVmppd19ZoA9jN8
MaI6guZmSZ7VoZyvPJFifI89DojtNdMoI5t+tL3RlQBqQ9Co0CAEpRlAreWEoKKki/P3OSMztFWa
rk/X4dOixytN0ubIEeNtOPH3sBHlaumc18PkhE3N1FkbklGO5CzS2F/VVK+BGWuMqqBNxaKgKzpF
qY1IVMbAPMLysDvFnM3MZKvVmQao+I9bb1N/X8RvF1khO94rWtVIN4ZpgmaPI0Q+IcDwZulK2Puc
NEsxa2yulYd0HN5mvH8xcb01c05T9mwP67lwmL5/uP3BQP3ho/daCab3o0/hax3CBlUMPOIy9/Ck
2LwK4CJAPkwNxsWtK76RRCTKmSgy0PSUeRFGOVWV9tWDkgXIOaFN7Ks2/bwPVPgq9pyyBhNL3vdI
DZ95ycSciXucPx/et2na0b+bXUB9AmyoB4YRz2LtZlJzyFVT5yaikD4Uy0n/wR8PWJ3+ZLmWUaZ4
MuwrCQ4Q0OGO/BkFvIjYuNrkP5Z8V9l3Zc36A3ClLUmZXty2NBIw36PtdCOekrFsE9er3cbaUwFs
ysZ/CvHap+7pyjhRsEAoxZpeCYUq8xBIUzPlvGyYN/VJ//H5T+a+WcA87RJa0URgusWAipyQ+j62
fH42vwzpsr2UkZ+8qVPFcKmeyAdycNUTl52RLkZuLPFr/53KdrLUhWHHQ0FOqUf1TW3j8ALNEZzY
lmVXJ3unUu2bptLoWU2OswIhYTi/Ba1o2Q/vBBGTz3eMtXo/2H/OqjQrUprDgsOH1uxdwtGOQf52
yq3E3E25CGlpXeHBs52qpr3sd6UwjEEtMc5pcaf+siZxB4/Zla8DbnjQy7kYnVwYR+WCHo+VkySY
ofkWIMZDt7JWWDBbVKVhk1ozFDPrAB4EPRRIbViIo1rb1CJC4vBuDuYlmN6TA3AeR3CXc9T2Ua2U
1+PAlWIXM12a05ZCFb9hugcyU7VcAFwNv0v/fr4vIXdIE+RsNYo3f6v8ZYkLQx7NqSlLTfha4FnE
M0Fzk26foSQISZAerMunfeZGYZWxBNUPff99ILRg8KlrG+nomYbAzFF4RFETrQUAyHugyWAZWB1s
Tp5ttAL6oUB0BM8WZKNNQ3cW0qHaeqzwJodZ1B3L7XA2yqdpcbpdMg5tnygaQCRw50pBqOOsc7o5
TVo0WP7A6DAG/rOPVT2OaRbmdTQ8HrkXgJzyaAvawPvGDiod5ryuKtIsmIUtYVE8dg6VAvb9r5ST
4I9CiBIZxK9LHwaUrezSkIYxDyqzhBQwblj8E/j/axlrgcFtZLGTNm2rIBMeRs2veSiBliZiLs41
r+ZgulGbHgEPEfuJ/e1Tdmmc3Al2YqtlcfEY4TSOVX7czBB5wq+IGLbn/VSL3bTlvMvk0gEH/6vl
0yOse4PmTcqrEA9C0vdSyQ7WFHGQO/L4i6wt5Hw3mXq7BZ41cYZgWwktHEHBNFnZnQa8YJIrjC0s
NTaIgJas2GmPT6CYgSDOVtNROzHRzv8jxKDrMbcgfJLomfxYqVdx4lvA7eEap9jjuKd/Lc3cTuBx
UnpTU8nIncpAonKhmsbBb3VkFVf0+mz5NbhEPP3gGZhAtcApqF3Yga5VCCMfwMSNNcaUjCodnNFH
lahqoRieikbzXJXQmGlYow/vjymBRF4JzNFxaNY+NwNKZ4GWI1I/En2bCmMQbcFrM52iiq2ZDNKv
PCQowbiTDLo61wcLq8m7I+DDo/4HsdjPNBxSyWfnbDGSCx9mozktnjlY9PMjb2uC9FoKa9sGvIWn
ZelapVfTqR08BmS2p0oWtCrH1CMrPrrHU8BeRKsxAU8q1QI29WN+diMFcEeoPtu0V17EqxgCosZh
6YeO2Ylvbn25Qzy9aIQlYSux9I32svEBoqFB+BBafe3rdcCKUbBzLfk20ZJFqDF9TEFT6DvDymKG
qT3Lcnjb74nnAngYEOGZLFCD16ohqDk9s8EYxMHGWNaQrOG/uKvg3uqrtdqjGemrelvM0cIIDVtj
NHYa5N4YEUzeF6Fd6/SnND/xnvSUjeKaq32h0aEHfmXzPp6rjFv45P8tZwEvFgzPp/UdPIidiNe+
2F0LvCoIeq5Y0IlgCbqe1HbgFVaqcq5zBtIjGX4eHMgO4gXbFsAHh4V5eCT4L/vFXdbLYGpyX+9m
zW9k1CIhKsnFHthHJiEZXYgq3kiY8VdbO67ol5NrAPXpoFF1WOA7Hd0uCOAQM7vlpc8u9nvr26+Y
xlkZiZJL8A3KBT0S2K9hk8QMGIhjI8R8bEGUWIQO16KzKvGvDo6Mbzor3bx9SsK6ScGhvAKKgcBM
fTOdbVcxQkrOvFiq8lwM4iUuQr2XgHn0mfCk6ktlAGjX4aTtq64i2UP+Sco/A2JyWFsEYkfi6oz3
vjjHBw4e5Hmmmu7O7o8F5a9U28sgslkKN0jiInBOOkvlZtBTYDRWz5mCWArr+Y1QytH6KchazvpS
TpBPHJMkAJIn2q2dKdLim6E52kI1flYEH84Jzsz6GA+pk8GMCrpEZn2jL+Ca/TPfMCZf/MTf2/wa
XwlPwOhldKYpRcZkOybGIYYdy3p9bUmkbW55AlgGPF3FurBKpl+bkZoFB9qBTs7ks4ETbjp/Z6Do
W78ce2tvojSSHg9KRwUejblk24CWdONr7WlZ4mOS5YuWxoHy9ogiU4C0Q8q+ILWNN+mwXIbruE15
jZwrxGfcAl3Jn+9bREPU5Ck3QWYEEcaycvv6oPKt/PB2SzezbjwGsnIGOd9rbiU0NujeH3PyVHHc
qbicKfzmjGQ4MnTUET37C63ctalA14aW/otLKOcT0mI98w4SRsqpqu9wpdekYzQ5R9fyXRR0rR62
3UwZZ5gpEgUkIqfVRQJtUJvIEQtO6bDfeyJjSeGUo6A7+nnUMf3oJVBwub0sgrdCh87JHOZzy7IL
Eaf015NYGnoewV/uQvLqpi9DKL3OwEUzkRsMOqdVp37pX9fzZQ0NY62BULECZTgi7lxQAFdnlQJ7
NM5t5N7gMFm9E/W09SRFosE4DWWZi+cHwEo9LTy8GblvDYDc5gKlT40d6tPzGFMCkehTO2AjEKPT
SV/KagEaEXX2dCSh5acthxsB9L9E7QA754P03p1fQMzlFAV8peZkWwr7Se3LawOXAWZ5ghA67vzc
2x0utDgmz9eM6rEHN9VqZXDGAmEj4Yndv7DlNxbJjcfwlk+tNfk0Cs0Ib4WN4Y5mEmSCyJCK8GVT
VCmPQ9huZXlKSDUcLXIoPuwdRyd3sgMY/s8vhFhcxaTMJnqF0ikXSwLD1oK8I3Y5TQareRVQshRR
+WOPblD391AyGKFz5yYoyC/XdT7cJlKJjxIZvJ4kTC+0mA9NeFhKV336U/5m+L9/J7W76vgpRcKU
t0MVGsR2Ky9b4EYUTmoKdK7ooava3jujo2H/ruGKY5drNHWc2FKneiy6CaPGNQnH1AkH/tujqMrd
g1UpQgAaEuPvjKgvKH1cLG9tciYpdN11XbNk8Bt6896HxT7sOw5PckJ7LJo9HrSIBHK26E+ufnkm
snU6wD0zd0hUhoxV1/9VHD6kLo8hZT/68cSf+ukMhsWZHnorbjZ/NSlgVApuTaPapjYO1vTxtU/A
wyBLlQeZM2zSg4Gw3zWx8qcPw+FRkgdvDyb7w7y8SIQ8MCM7Qoht284MRwO8iv+mqOVILST23gq3
RbClaSkUd97G7rDgr+W8qI+rCaVRGgLYHcxvtrrfNBIrO5/vTMwi4OoVCt6jR0iL21y2HVufNBg6
CvbDLBSIGhJ6uuHEkHwL1wLTiNaVVBCqXQ0Jz9sYDimeWHhWH6z0e13ESq4c3Wk0xRrrwFhiHmws
Gn2m1rXOqNXvxg46UexmKOGFCZxzrM7jOAUv5QhkzSOrDzHn7/aAxFk2+D7QydUPeVgHAQVz/RT9
wrf/72yGS6Q9GPMR1fIokm9fCSrphsp16vK98moZp+v7AFMo2mag+g6aWqKC9mOUIAL8TlMn36U1
EdfjeH/6yNA9Ljwi1P0ayESfg5V60TCPtceuantv8gGiF+jRtx9UjjhHDWwZa+QlHAeCJz6EVzRh
CWv4bVwmOG1w7AWFvMLFYdQHCSf/Hvv75GnuZUYHEgpXsO0puszmGFJyHHA2sQhAQR3ia/eZ1M7e
KGkYGTbxCbdusgSKIO++NJwbrjQ65L+jQBAjm4KAiUqc76CDjlvwbaDQDrPATXOWMPKFH/2oNPub
TBsILme3ZP4iAqVKZohX7MMAPnb+QP34PYzsfLMeOcoIDB8OCXPhjhib4TDtRLvXEEcm9jTjoKmU
dnK+O71NisMviFw3pvgXVlsV2oogas9Si7SafWIsSetLauSy6SqKIPuhVM++lVl2sv0JieSjFCUU
koIHuEzwU8AH4JXsvKgNbLwO3hTbol80i0RzsjDF21g1BcOPkxp0jVl2qKgbqTWKMBPRCxCbPQA+
2jkfRLqyHC0f6DiDcwOGj27bISUlRb3hUJ5QdnoQX09Lwp9KTE+xQ78icxPX55Hy62I7g/K5HtTf
KLDFfLCVQFZ36WENOeMO0Ep4sDHKprftqbnMdkav0P4DakVDlrZJ8YQxuG7GkZcK6LEZM8avEs8u
48v1y/A5t/sgGABcjq1a/ST638jjlvlxRCXx3LLqpWt3k3RFzuc6Y2poGKbNOXJi368lynis6r2G
FcTxMq1ggvGPsHI0eVeMjlxMPg9qZN/sXNHv24JiFyR3p7NoDEyrHqPdOkm3qK03gaHL0issAEDL
uELKUI/MmrLcGtlp9lqUIcACIhfw3az8C2jsoeYnTYSQzHT6V12dmLhYqQbhcwcI3VNoGydxX0YA
ZNY476Lup7B9IhzAvB5mfQLUKFkEb+s0EjRZ3ACVULSRVHPdMOw6kPQ2ptDCg5P8At2NKLG/2s8q
iAV6OEG37+6ni8O4/TIK5OcLo+p4QzzTWdiK5aFHt3aWvgx9kzEtNdsriBylOl14JmhNwXrR74/a
mRFGaLVC5EF5cAn/dAAyK/4ermniqcrXg5PoACZWo5B4K5uk8Z96LP7+HdpQQTY4ZtvyFLAh/Dpk
klNvQzvm2E3VB2fWWluhJE6pVjfpwBkZXu6bAgckB3E9OjsnSZ63b+5ZvRlSwNVNYhNjgQFjNo+A
g/WdBbfSncWtvH+GXYrTUaskm+12WeruqW4CLMCRPAQnvev0FmZJ9dQ9IomTeReoChoZknyC94Cx
W9/GG/a3JWNGjAdFF7NZMJovCSBqMV5cnF2cIrVBhPxMVPhawX8NKKAq/lVsQlILEvlgig9GmXyi
83pC+m2z9s2QXXtqDdUVDu/A0F/rCEmSst8/lNoaR9UQdBWlB5gam5mu+lJi9Zur0h+1MX18iB3T
mrY9Uh8RuZ2Q6bfmF01FNsHSMdVqmdXRCH8lMz2If0Z4do1Z1iI/waOgxK6g2HLT0Q1xM8pEKj1Y
vNcJSV04h3Tu4TF5ee/oxYx2PqinWJUCWzOw9NjmtL000+0UzEaQKyMlYV2/6rMSQe4xVUkPnQsS
kJeOpnB7BXXErXKDgtsJdTK7/34wb7HKbm5VBFJ069P2gqispeZu/J7NSf2BaDjJD6p74dVQdLaI
jesjvSfiaRuwuTRVDJFwTrqR8hpeycb6oYzeVs6oFaOEY/vFgbQUFQWsNCKIOvQFz4BsMgyKeg1u
zMPHA+Nex1YTkyKBvBY+caAhybdVEWYJuTXP9KzMBMuwn6LQhHFJ39GymGPPJia3wbArhWV93v5M
cEA/NRqMV7HNCfFlMxNOcjzl3cdY0Ofu66a2+/3eyAPyBJFd7SKn83B3lGnZdIDyFIT6XcOj3xoN
bF/hs/ms/+eZODJmsy/Kto/W7FKhaiPixDzfGy/pieoRVuTGvpRlIt/NDPtK4DJCJlbo7aiVDJin
pxL8b70isBwrVgMjJxqHBQ6HO11hY2DT+JxX6SjpCvaLDbfT1bp0tApBcYesZbH+EgxnlkMlc19I
ApIqNmknGVNp072WoQtkH62iDxZv2BwGYcS6d8VHbztaA8iGIWJf8jnePZ3jejUKJK1arCy+JX1g
lTO1unYyQ7DqDq8aXXila4ikzi3+juhVZ8EiC0aSMhxxHe+dm+R0pp7Rqo/8t4KXXaTbvQhgTAMr
1LnJYo+LH3iHutnGOvseldWzDIUpEDuPxDY3s1xW0ICRbDRIX52Exga24vk/rV7pYm3OmkKN6hPk
sdVF85xmZBIJiMr8gnU5SjQQcioGpwjA+jVTZ+3X3QBcJKoCtVWd9tU6vCUlq3GNo92+akBW8d56
T8OTYLmn+pJyUSEfeOtnw7N9q52Lxic87U6BvPNa2bb/Ct+8OQsnalrVG6h0ynYlviWPFhAO+X9G
Etm1WahlXFZv0CcJ5nAj9d8Jx6jhH9CgB2ZkuOdLpkUmNIfh+cCkGkHrASETDFiUWjubKHAlEV7V
ioMvOKjUVIpLe0MHiCZM2GSHAzng3HIhFpgH0bsj5rnC4B1vD+GlHcinhzdx03JrKH88gawl33dq
u2yIpMJuZN3RoNCF9VUGvrPcHSeg7+SKGKHBTlIkQUbPj9CxpN3OVcKNKD02jctjpLVI76s0AH5h
ePQKS2L67ARnfOQA3E5Obs5lXZ1XUP7100DkA3u1ZQf2Y+PiArDEVcVAALXJaSsnVa7kxhFrng44
PiCvZfsqtWE51c6IO7/CxGTQeUv8XoNPL/DUFQzXmWMWbK/mCHnxZig3MC108wzh+KcZBozdbVf9
PydP0Clpb918LhS3zt8k8XTcetLPt7VI4fmlhksxoWUE8jR1ZvlR5cL47KdNExtOFkhHmYQE/X2t
w60xD+ZCvHivUdWpsD71lkBpZ/SeJSWHiyaLN87t24hzY/mTkYyFyWOn+FXquF1YihTJGzz6k243
I67AqFCmZk/WtFTgJvYgWFr3VEnLtJkVEVKAmt81YhpWdMWiH3DbtDlGAJX8yrcjGK0hjqnGwJ5n
sm8H1aRwkZZyJFsFhulBpStdmYEKhk9s8FDNXD/oEdlvSCKdnSxsPge9nui2phc0SLtBQ0V4jnHL
WwM/uAiMkD2ejSbYGIO20y4zVkCQv1C1LS2a+q946HToMmGfAehNL+bk2lgDI/xreCNViLpTi/ik
gYnJVBo3tIII5FReKsbIIej9y80cefsLot93Qqx+6MnHcvFDSa32syqLT3L1U44cl3hyhIvuF9p5
yZfYD8EgNUDOzevbaWl/VKMPNBfoJW/Cp6q09LktFWMV0ZbROsmJlrvLc65Yw38s+EbxApwK2LgB
Db1BO9gocdOz1ymP4iERQgyr6G5feEDOWh9nVxKV0mZvebaSeUb+X20oGn8aPd0UiVyTERlAoV4T
lGgTQ8xNIZIdGFhaFhGY6JMZebCoI6/V5YgCVspnV3vlwLgnn30F3Pbr8G8l3/e6Ne1qeS7H09Ei
uAfHaLMQFA8eO+8MyK5hmK0gOHC5N1yvf4dPlNZTKkm9qFIt5VfcR1iEQEbuuSP9dwlX2ih8FYIQ
p6BsjaNYptuiY2uhj2cDp0e4mfnDdz0r65pWkB+uW2RnywdcQBwrCBOWf2cK8e5P+Zep2GiaBUv/
uC771gEeCSo1ljxNwP5QDYItCeQeUJ7tYi6DsEQYckdkISF/mXndwukW5ekDpW/ewpxKQeg29mmB
se6kehFZQMa1npNq81do1UMhli7C8obY4m2OW/cDwe3cknbPRSmlkB5qiSKgnKQoaXuudLSomZXS
V6pRfUGLQ7DV4YVCDUSdiVv/TyZ+kFQjwLfBaAReVO3F5JGzJPDFXR4Afp19i8uvz3V1WCzwgPX6
Hf1weuasfEm7Gd3i25LBX/zT3eTB3qOWbYqmRlAyXswJKS51zXlyA5lrT+0M/9IsCzP5ynSGmzu1
vCgSnIPZ0tpEMB4utCL+0VWrGaexKne8dnOvtXCgW8pbQThL1+TIHLx0oXR8681bxmweJiArQX/Q
aZ1GdHwYapoqIVt2P+FIL7vByrB+zzjQQmtI0/Ky62uhZl7pIbFZX6a1D0LKawBRdOmx8g+qTTEc
BjxDDHlj4ILGgl45AN4BRJ5mu/c5nKv9njoBovz/vaTY869r1L+7h8ltQkHjCnpUxmQZhnmrHKMu
9/YARKdyiaubNXmRCpkNoIv4R2ZISoPXsF2Bnss3aeGq3DlWY66LpOL3d+EwdJb+uTkfI8m14LJL
FVsOw/+NE8LSwUemZL0adwMOdOVes78QbRtFM92a99yAmwSmZdAqnTQiVcg+rnA3UV2nUoPyb+WG
5y29Hl7NlS20J9S2X9Is+d3CsIA9cUQ0hcCTvRshCTykn1qDhd3yrSXiauKj8cKstiOnAQwGek3s
8ptM9almX+lo4iiC2prtNQuChggIY5eFdgj1bYTNtIteXDeUkjlu7bhdo9PfGTDDpGCGXUFrComS
vKMsc9jScaUQXs20fEkqREEArfMoCnnOIs6dzSL7prGHS10VT8UUDyN7yTQRIYhBFno3PieTnY8f
sY2heacoRf1X+jdRhjArbA+tAvmxZZP4P+e13YBZ0WCQRoVDkbE7gzui61C5LsjPBSffc5E+BSOX
Bo+sMoguk9mMNk+APcKbDMZkH/ADtSuPH/mgGa3BuD/E+cD3lC1O8zCF41zUBK7xpRl9M43U82c8
FmjdhfATeyvxG1BFo0nAjrUXnt+91L+NJ9HaN6VlKJQSGgD0JPAM/9WoMwYwHLuIxXh7pmr1OlXl
4FsWEU0jxcJRgZ49Mwo8XdBplWHXpEGJYhB5fDDjZoDAlcK6LgvujtHGzS80WkfLP/6VYmyNwsHl
hs6nSqX6RdlyLvCeINpn40V4mD1CHJ4uO/VWhGrCtCfa3NSdD46yfHE+2tAfHBlP6PA5+o5aLPhx
QRJQuPhe/HG5xFVu5/5C6PP8D68UOFZGZlFmlWvqHLuU1a+d/jVSS9DLedaLdMxhca5936ADHTNZ
vw87DuycpjDiFa01v4jf7ZmzJCirkJNWIxWcBwjqIFh0pAGMM9mGuZWa8WQI67m9X+zxLW59XO6U
cJMz36G1+Q1jWJw0HfgqioiRRDgZkNCoQProB79u3OEdQeR/2RYpdlosKkIWyXNKaGN3gWJz68zH
vE1TSN604PlqR5v5UIGEX/QUvCzyqOON4pzuAwinOpPDc2J+E1lbSdCgVQBSW87blmHGbntzRtbb
r62yCwheh9NDYAwWhukT3MwLvDFBkHUH9CPSIVaEB1hUXYFsYPo+BnR4s8U0CMXCz19u5Dj12EZt
Fa3iG9YDt4RTh0M/lTAVU7Bgv8Kyb3dsEHByuUkoQKAcjK+FBa+NUSdO/+qMXAX9EVcaPvRLNM2z
m31sudVM6QtAQcp9QTc8Jv8asp+BsQw46PYyzchfXkPUtI8NiHZOazcitRuPodErpjPycZ2H9uJK
KwUVDiV/3FxxhBTvf21kBOUz3bYh7yNU4KrALa1+HcreM3LeKEgTPUQiwzmtyQPlpDTMqhbwTFeG
4e8muVCI7vE1cA6psUiDAvI7YPo8VJBZfzl1oRIBXjp3awZDltwdD89gbdFE/2JJZl1QUbsBWmc8
VlQMXd5DMnLpFFaBUNUE3/G8v0GU1MAQIMuWXy2nHLddGLTv70Pv7jZKnYV9YEQ4m7Jy4VojIXu8
rUAEmkbStKZo7aKhQn2ATVny+vzzOTMJE52+ETU1Xpm0j0MZInRBFjH+PKl2EaABp32Px51Xhs21
5aVbgAwssKQgCxNT+HaI1g248F5ajKEaJcHIXbMKZLnhgMD07k5yEFDJ+y4qMin6r0UarcY/b6y7
8WWOgoayaO/cxR+4qQr94dPMUt3L0rGfZqXI8VC6usGQaF0+4wF/Yn/sYuKzuq/5K4ADfn4bhKVg
k2cgudXC60oR+kXsEPjIbmuuEBU29bVqdTsig+FdrIvZlGD3Tup/L3S0jmFXZI/7Lp5r8/qmbhX8
MaEcp+KIaYdQRedvlhAVrvQ9TUcq8z+I6KkugDEW8Dvxa7F9n8Vxs7dRKirQEVlqCCgXRpxXa73y
LrMW1ItfYaO23IK471tnbJMXLM+7K66dUtyCDIJwWhqHqr4t472Xyhcvlxqd5YlcEGTdVdaLqU7n
V+I0hQRejeI+E4oeTmVVk2XX+85EU7yT0vW7x6/kbajRV6iNmzZSy30T/7h1rXiafb3lp2b5LRc4
YBN9aZ1GW6X7c3Byke8NiKl3mF4/ow313qa9c89BbbhuZEx39BenQOpEAnbPFvkiQ16tQHWbjksw
txkiZ7+cKM/wSryqjOTbPKywniFe0DkkdzxsywiOtvYjYVXvPfAkjMlKl6ybu+k2E3GKD1Oxixlc
WJ1NN89xK35dermWZZeNghSQZbqr71w9N4Ap3tc7YFm6BrCBGXiXaXpk9lbsl7aY4MhfxkPpGqr5
jLr1ZFml6D3wUDkvy7I9D3MoQd/DyRDjJ5TlUZ0SHAPBCqk3jsPCecemzIsS4NMTcuI2zzzQHcDG
OLSkUYhNdCB8KEyv/aK6AfX3Zij+pQ6NNYZI625uSnIJXqBQXK7X/U+dHkACl/VWL3InoRqBcmjm
xbqzXSWgYXKJsxwn6FI5+OlUmb8LSgJBnyQUkxVcOHnVFUGZ4KdrsH7BpqIjpVnvO1DvGHC4iDqu
OAsAMkv3cOLeGW8R0AFwwq83cRjZ1wF1qed4K9X9MpSVVztviSjtMIsd9usg8B/L5nI6HeLblvOM
xSUzHIhSRnM+4IhE0DT9cn+CbghD8QVXkYozxlfIJVAE2wQmnaD7FiIg0LzCqMil5Q5I/viD/1i5
h/daZqmmPDq2Pg0BNtOLjmXX7zoUM/Ge1LddE/Q8IDhcswa5dUUW3B5SuQzludU4v++MSFJlPnhj
TnrroQq2j/AojHoT68IogjGt7ebyhD0HxvI5r6+k/dOs24PmvMWdjb0V1mJZ9wIe5gk1gcJK1cxD
jgvHmh5SGF3fv+1lw3IaxF2cza/pXW0pQJKuWuf4OkKUh41EFzcENHrKizeXU2xp95ZndYFqD4bt
8MJojKibaADyE9HaFnoli2WuDfOFRQ/PWGbWJq22f+dfo4Zw2Kovuq+OXNjioZhdOfqUY/xktu0l
36GWIQ3UJiEcTlEg6ztrxtBH2L7VIYtYlIMb482acc3SY+QZHpior21XzKc7WyRFAVsA3mrYkilY
cmw6xnHsRs4paXwQsXdIy3Cx1uIFOhcpmlZYn3FgiEiXvgHNExN4KyTeaskj9O36QJ5OoS0tOypU
OhcnrJjBjItGQDGrYNBdxCqQ349uCMV3vBmTj8kA9Dps+cpkTGIL4OCuHRWQ4Nqhf8KoTK5/MI89
6w9/pON/aXHBTrzrZf8/l5RWenM/VoDC5Vk4mARClcD10DL7+Inw5u4SOWwt8QyvExRg4Vqt/xGy
/nhBcrQR8PVDznNL6Ht7v56kW4jkuoJS7OFvWe4XeUNfu2KixcjNKFMn2AwAU1X9tr+CEdexOMdY
2VQCOTYYOpC2QPD+tkYuj2vJD5WjcIGZzSPJhqOZq/3qKvqtFvLzuo2LWM1dBt4CjjnLHBSm2ovY
rcG0ubBcsMNf95BT2UE02Nf0iMfJGYiJKTd+pqOyTNC9VfGZw7mp6CnN2sBaULv8woAuonLBL0An
272xfOYTm0i5DzlIMuFNMPru5OA7lj9e5HrOLq247rW9TOjPta2GdkV5Q5h/1oMBwSL8sv6s+Z19
AH4gErsL7cZ7AtecWmKU018fKRCqBGy9+gQQMOulBnVuleZKNLo0V5LLqusYMmydSbjERyPs7Bzg
0vdKRmobZqrnWY77cB9dqrElEfBw6t5fdFUGHx55AK+0+1KPtJ8cr8AatQ18jjMi/RMwXOYlCs4B
YUe8Gu4EhnVfzWGe4/B1pKVJiNrPnR6nrdNBYZRSZL5+uAxxw1yK7S64fsqeKJ+Q8y8j+BCdl09R
Gp7thNLbSu/kBck02sFv7WCpN61z4Fz8ZBCOiMSRdpl7HgFOJfR5hKoSgi4ILafPHqNec4ioYn05
/+R/R2tNCukmiZ6NsYar3PUY4k7ct6FJdwnoAgHEFSsETuRPkiI6nlbt5mefhR2mYRn3a3u865H1
Aw96LEuz6rjg0J4keit3OR0jtLFgZwcdV+yCL/9IZ0JVg4XqTckxOKmW14oEHfBTwUV2vj2M+Jp/
CjNBJdeFfAisfIwzpCHs69UdyLug412/y3Pw9a7SRLbWBSf9Fu8C2VGGMDSSa6iCHFuHfMmgLa3A
JEJTdh5aKrHjVnOZZYr6Qv042PWChUHkuYJJrd25xeOYfVSwUvXgRHzOKRLASP+bodvjJ6Re7xaK
HZ02YTE8TU1QM2O1AZ6rhCBrhrB2spLXVSw+EalWySlwRTGzpUkyud1CRHzspg2sH8135xonaXnC
qnkJTulcL2lGcDybj23daPYwbfGud6oAk3aHKxprbQRzVSpGc292q0nRA1KKibjiMFvHfeOhOMaL
pIBvx9kttxUhKEdbGsbPTajpEzG7NipKyT/DsiQul7Tvm+Xy2Wth3KhVHT6nhvE290a/rqbGbnZS
UOVnWyY+WcFHfXfR0k1luzXNXuB308Y4e/CExbdpmPzxSBX0U6S7wP2RQhwoqVXsYFgsP6t57wfP
WqOPPZloT0t1IMrqGvrP94YKIp1Bb64dAnXmCLkVxWaMP9/Vt/tdJXQ/nM0Dl0shnjbFuqVZ1Jgv
GziUUCo0tkmGzWyc6E9Fq7MsU4sqrWKrHW1GfGRFAn/nUJ0RHAlktKXpCeK27DfReax2Zobaax0R
sJ9sg9XFlPrkjbf4IT139MN3w/WjfJOTDNJGWBMEBcnxuAqcBFwWG+oVcmuOn32Y/R1l/KQ3rCTT
ECR5Ew/VeeNXBnjITYIbL2wI0LuUPyCK4kiC95Cn2AyYZi5Iicf47EDv3AJDcxUQumm4MaTed0Mr
USzMcmXYZr3OtIyEwOfV34Z+3lAvBOGOgFsHmwiktZ8jO8c3OEnDj9rscyPU/jAu5IG1DCxCROf5
GRc+f/8CvfVtxWq3UdA9ENS03PcjCAUM2Q6w8tOuFOjGRUcng5FaungyM7DPDnKX4MY5EJooS+VK
bdCwTx3ZiP3TWJzv4DjR4Qutaoi4A0m7w1B7u0qxXGVQ2TS3hVwrnbLp8CEgJpFWZQgIk7f/ZJ6p
T4AfyYTRIklv9JIrP3J9cjvB4/QlAqxo+bd9Sa1MZVLVF/NOxW4eeod54NbYMQ50AxJO4T482z9w
fc0JpFuTjV1ZLq3oGxtZA+c4tiM9M9lZMfDb18x2Nsn9wLQwhiqBmP1sjCpEvG1z6KTlUZ6EXB3g
DwXI8JTFZnlTshfzYRJvj4CZO4KnIhnSZsS4fh9Bax1r0lzffQtD9VYgneu+rQfad2evQMzwqxQS
dsOYcewDda64YefP/R4i1J9wcxm7EqaoBjzrOw4V1EIIRhmNrIld0e7o+hSecRgiLjcmHBzs8GCA
NiU9iB867VkSDuELl1tbK1ZX0a2afuYLGRXOGP6OlQ0NvoWtdIjZDbzkZs66puOYaXM1lqF0Qa9u
gOyjZMZI7l2/Ke0DyOUsB0mrykd62NpIRihrWQCdY2YdUyvzTet4WPBcdLSRRV3cqRy7bf5S7cci
Zz0wCD+51M9qIKS03c3/+23Rx7Qw3OhO+3El118797q3mPiBj9AUcm0hqaODYZjse4hCqyRPwDt7
YBqE+0w59vCK6YiQUp4jpffptLtMl+57quqrGmLrSbU/IBNL/vGbMS7v/+6WwkPC1cvJ+SGPphDK
bCnIGsJPoN6bQolOLfpIh9FOuKs133On5xuoe69diVZXF5o5H/H+YztNVn2gVbRrYLtx6nK7F9Qw
lIjFR1yg3s3Cizc5jYD1yq+U2WXLBmlU0UQFruwpyhfF0S/KyTMaycv4scKiIeswG9+XUZ/10g/7
e5qmkd0hqd1KYI5f2sI9odueVYHiG1Qy/q/KdVBimaiMb56RtdmlXpukc1ynh3M6S/NnNC03MsKg
UyP3q6Jv28s4P9TGNvAiJkvExAUXBty7y0IRCZ//wno4a1TAxtmHkcQuetNmTkCjk94AXkZq5Nj4
KvhekZG+fsBHgjR0X+pFdO3ZCg5dHdi0aynWb17RZLLA8uiJuQ8duhYFDs5HLSvtZJEnTaN+hLyG
mCz+BXF+v0nR8BqqlLPbfRgWrVkgTHo5QMcLdwE9AKplCeHQxp4v+NfakJkzGPDJyx8j4Jq3cbcx
Q84v8um+WVRfbcAP6A0lTr0o4RRFMDjuGRtYPgNbNyeCT9DL1ydHjokwCnloSAj9Ar2ixj9v4Nnm
DQJCjISpcZ1fjjLCFM8tqGk0EjigK9kNyGvgvTcW7H2wF06RWlbi4P8Zy5N1JMqZww/peGpKUUxu
CzEI/lhk4D+7PqXg6/NvSkKR5KEY7U98hORnzwv/yzN9LiE9unv1oRxroK1SrTaKozGbcrPwA8Og
gYVI9B/FwsVIZ+9KWVPdWQ5uNwTbYoey4o5Gn+aAs0jKfQHPb0/n6K/ynTiKqcbRrzozTfqRVs6i
y/U8+Ro/BwUVlFRdmkDCjAPUEv+s5Jc5/WTgKZSEwhTI6464ez8SLcFc125UXJnXmo68GYEb+hrm
IdesmUKdyt5b8SuxMvOCccy1/oYuH/B/3U3InjFn+iXM3Vw409CepbdgLVv4tfn9gP2NcvjC9ktG
Xzq8b7c9jcoX+PZZSux+tUWz06XXFYq2GDR7xiVMCWRfzoxpo6rpmlauizcog7maDAK+ItPNpLTW
neyWCti33CZ1TNGvfiTwwjEoQPrpjzOXRIpBK/k2bVyMNo+qMiH21pllYHmTfstANlAb7unEAMZa
tJvJYh6w0oK2x77IdKblrQXJXXRdpv4YdaTU2EQJWNQjLZrkQaVBPAX7apckcp0ZWEUzISAqjqKn
TaTmF1eI2OepWl8GTv94vJdG6TkZzF7b4j1RX7hYk7o3IzwGMPoh7NYBE0dQF71k/P0god+WWbAs
rWCpyQbBEMQ0t9nv3gQq+ROwX1zpuBfwSM7gYAJse8eK6WPRliaAr2W/3vC3gnsumd0/C4XPNO7d
RoWZCMgOTlOyjapM8oAHkAZiMwFqwW0FqLVfwOI9X2eeVIkUXkINSejm7/3Vcc/+oTunQ9IbYOEo
PxEAW3Iilsb4ux+TR8xIrjI1222FZf/dIb2UooS4DEDrYTvLGPEpNe4UxCtPTwHQ82jqMoXTcCpl
6+6WG/jiNkk95rQLMU+G0Sv0elKYriJKNY6WxsuPuqdUc5pwm2UvJVTur3ncm4c9HryKh/tk+1Zm
FTcPNP5E5FuafQAHsEhp+s5l2BGMlIQV4YZck6zkMjK78H1qHLalgX4qRDrYENtdz0yKc4j31Z4S
xQpZhCbVDomgAQ8MlJyMG/DPb5PltTYe4KUowjDzB6Zisk6mjsZHTR15UQ+vd1a6SGhWLbRHM+tQ
RgqkcpkNXEj1cCVDn9SWNDGVrhSRc6LTq4QfCdXCXpoBTC6b9Zzii9gqhJ4EAmaZ3yzuRD4m9O4M
JFAwzuKtJtG2AOWwd5jOJpydprabfMxma3wz4bp/JVb5v3gIYX9f2/nqboM7WmaSOujoWcGWvXTz
uqbW7KE2NWfmmwEl7zNbPP54CoqcMASpyrux1BzicCQDmoIqb36my6LcYZSvhUE+wv14BYRRDGMW
bqe3Q1zKE2vxoui5LPOPimShfa/i50oAMVcfiJTfYGsk2t/NwVK5KyzHT/ubo3FSyM1cu5gxunzS
y6O97o2ifWB1y+oRqxQ0qKlIb073oV2qPC3Stu94XH2yOxAEwAr1MHJF8RLZfzuvCl9ZkHXzYypc
/DlLp2I+rr95LN85ZNVmuVfO9RWboLKULfpHaCIqAlwyk/MeoNw7VS37Lr6/4rxbpHqcWrJHiDPE
lVnIYnGw0vkOOCrROMuvQr5vrZezP9jPnCRuOSPIWxa2HJqwVbF9sTf9OCqmAb0M5zaHGmSaLmYN
pwxTrU5Ks7zFjXdXGHv+riegItpXRBfe0PgkaN8hJKNVBJDkm9M3qNr2OJr33aW8ufl6X53uhcP0
2Ou2fDv7UPyIwrrhNtMSwtkOQJhpWMzCA7GlwHLe99nQGP2zDaJwPekh3nbdOJd7nZlYfuNbtExV
2xGZEfr9uNKVsSWfvmkS7Gz2DeddjhnztIxUXL/dh0BnNNk+85qCVYRw0hQqe+vQ5SSOe6iMExBF
0OYuJIMmcqISJZzcHZwaNEwi5Tqpw2WNBpEy0QBzryWr1kAkHDL0cg6pBH9Zl8XuUK+aS3bk634L
rCL/Ea00uz2fBFQaG+N1SWsASl5bX1iYcOVjTGsCe1jz4JpvGGl594LQqYmcjtiWzFQMWxsnM87l
2uXgKiU8WRqcOqO4+XEYjL415fPluZMWqGzEw5zGXtfzaR1Y7c9yunkQbsar5q5zREw1n6eV7jVD
qfFvYwUMty29jbrTezE0QsADE8B++8IcG0PQ9eBvPfH+E9C2QSLZZMRInnfX5FtFfojK3HpYQlHr
VXyd6+t7W+Cx3XqcFKrQnbsUQkUbCqyrlyrREPtox3S925DPT4C5MXPbHZjlgl55QP2hykrnXzPl
uXPlhfcC9G7kH+VPFz3ZqdQQMEwlM23Q193P3kmIMsvBcp31DZB/J+DnTxyKvNvhLxQ679XxUjG6
gdXu/Otr03dl9VvI2xfqPzL6DrrWr3BZD8eCjMjWAVY7VkjphYxt2OuT26zaB4u+NZQnYvZ8asdg
9Vacn4wSDcHZRzrHj3BpyzwvV3QEMBRdJg7Eb6PsgANXQEv263HcZ99wescL2n0pcQR26A6zlgke
/Nv2h3RBilUQObJSdYufaYS65CF4nqTogLtslKb2UNT0zCuZ0/UNyd7FxYtEowO792lLpqfswr6+
nNFDQ0Nf6EBaoMqxabGCtbxdiEnZSLqclw2q+A9YO7VyUGi7XgYlBDadVrvl5bNyxnvElxlbU0t0
9Usc+E3fOgJjwrrLzCAuRBstfDoxrmIAQ9IsDTijQx06zjAqr1FFKwPrjgLYyEgZbpo/+kaKwTX2
zPmLHrC25ZW+rcnmGczJrbgEsWKkTiLgh80vu2EyuJuM/4uHZgj4kdnaPqIXzwH2rtQw1sNyKJmM
Gp/NqG2p0z/8lxmJKT3SHrEULKV/taFDbTmSvQXsvIPc7rhjdWJNZdQNU0T7M/94Wz7FE3uaNbL/
4Moz+pdH3j/QOtapHkUbWV9Y0uVJWOm8LISRCeiG2OVI0MpSCsn7pJ2L5Co7+wiS3WC5Vz8kFHxN
aO4Gk7j9asmBqK8J0vaaqFJWfrv3qDphN6S5AeENYvJFiv8H7l93XM1fLGI0wBHZk0LyZdAMs6UN
nQEIPfGza36cl73GTHxBzQPgsO/DJa8IoJLCSVbmn5sqHQ04Plzq6zziPoAau1Y4/yRL32A+KRJy
mAxYlJMtcEUk0sbuvDytUZxNu9Am4J+EhjhgqnxhDZTmz1Um31VfwrNUB72Q+0rmyTTFPyDgPNPF
Qqzsh1cvJ5+QwKE5xofqyghaerWhiUMhScsTefap2ZH2r40lIUaDZA0xzdi6bW5El3l9qnl3uJva
FEGrqdDFRRgkNEAkaajcdlMnaH6YH7rw3NtBvRwKUxq3Ft8Np3GuOLBLvafYyKcdihhkkww2qBuC
yZZnx3KHqsLtW9jxn6JVsvMAomq0TxavpdQd+TfU+7Hj45s1LQUL2Ts7pq8laa92Y3Ea+kg+bDTi
HNh57e/uA3OS7X5PXl/fVFwlDsThYENHTFS1eRJtMSWapgApo6V1nIKy5RI/cYaHsPN4cQIW1VAk
CJCwo1BBgh5iaTwQDllUsGZR1dBFGWkJg1qidI3Z4hI7PE6f3htgS2ARaLw8gRyc3/QqAYo7j6XH
a1ESa4rom8XVFGUrNwUNTBB4qY1tE2R9eBysGoptRdH4ndz6YPeZcLtfvi3z3/KnDUbJx9TByqu7
gJRSqxwY83y2Va0RGZABu7vKxCymTrs5kgo0ukhuqk9Ru0g0/Fq9+fHOe7Hp3RP5aykkS9Fs4LwJ
z3DDz51Bb9Qu5irpuXLyxLrQl2YYavgtGNA42rdtxtEjROPwvtfXI3VuN67ntk/NBChlPcJAYU0V
YUqMU0Kir1pk5tKnd9AdR2xK+Of+AhM07b9mXm+fUUsOs9YfSKICrNKKjNj2l/LNmm+nZKZ/YRCp
VhNekuQGXnXwOscEijIq91cYuzvIJrHCTCCumKOmUUu38yyx5jsKQvI/vhkXylNSjATjbQ8rCmj1
kDhbg+3pvZI+1/qGMUDg8S7y929/ujQNahpST9DyF/2O9A/ZuP8QErTrArR0hY3Qw/TZykezPhcU
zauMeBYQNnRSeBr3KbacD9lDRVAnVT8oFhCqo7PXKtZB9qCFazQIeIU2k0lzsdv1qFG04J2kvnvJ
uGp4SMOGH4qRjaPkFAb2Bdv+RZXd6fjDMNMGlKVn2i0PlQnPf3zWIX7uJlvHdHTezuJQh3wf/m7i
Dftn8I2Qde52wPriO4P6obmrjiXbI1rJbpvNLJxpa3JR6wpAk2rVjiofUDbxisDlq/vjSOl+lQP8
EfXC+j0396TLpM5dp10ujJHaRsDXQ5nAX8OVMwFC+sd4Lhd9+wCFlcbPi+ttrnHadP5CqAqrqDfI
hXJ1+wbkM8hieqxTcsDwiL45R0B0jmQ2fRo+yp98ORfd1eb5enT5JRRfbKdxDysvZ5d4SShQ/c8X
5z/T3NneJt12AX09pDsjIGF2VPK/nOHj/TPUYYbfGbr+44FwP+z42HBw7YvoWVJS4Tdc/fD6V24w
Wsgxp1U80v0ESTK4zKNQ9zRkiOc8sJm+b5ILOWeCclBpMlnbQMKvH3/CvFzdjgFib4VVwwB+FXhM
wrZJJCNRz4n0UCBWUbT49iGbNnAWI0cqcD/KoRaCEMnbSpIoywNJYB+Oqal4g9rJh9sUn/XNsXYg
7dzj7kWllo7BGGS5xNBnVckoQhS0YPvbI2tea1PjxUMBDtg8Ift3fha429uWLFlBOooawr0fyBk2
qtLoKnhLBJMfRCda3D/Wm0R3uV/0DbS/U5COxYZIrIK8Wa6BML46WBcTK2cG4XKhdYTRX7jDKhpR
oo0em6H/LgoIwGxc/COBUz3J0fd2TUYmdaOgrQ7dtkHkZqhbScKvNBAAJNX8HnOhVJP4fAnyQMPA
2rBw9joU7bvxqG8Z1sbGRYWFRvjhQebfMb3l2M+BJLVAwgzMSmGXvXKwWnLhKdR73s8gX7R0yRZj
gQQLD/AiqIlOqyH2QbQuTujL10jiWYt5A7VKgtqUKpMTYu3gJ/6t6IttpLzBYLrAmuy+F+miRiaU
SVc7uzaoephSUx7lv0hlG9pygfkDSk6geflIbUlIr6s0Q7LXAVfvm4zk55KrfNU7gnlV1g8E47Xy
KoNG24qO9LaMGCzznULQ0xAMfebVS8YfewIETpEGLHmNTVvWKn1LpjJZK90uoYCkpiyuwSGKqc7X
mkg51i+36G6Dybag6mFJt1prIwYlzmP1gXp20f01SaSwIdj29RSpHvn4bSfTqqZeGqlq9/gmGw+U
dzhdOQ2yo/E4KJPQPivzkUoeZxN/3d0T64oEStjRPVYq4mRpv7WwRgdkHyohOnaCkNhoRlRYI0Qv
KV6cJFno/qU85YsidNHXWZxVrduAhNQWT5SVlr1U6BmRzhOKh5ItOPSR5HwOVt0UBVusRxi5L38r
6V4XxCrkd9QqJ/bpAVHxeF2nARUiQYmX2xCFMyrm1GTzEnnG/8lP8/OfCZ1haiIhGYYhNo6S0S6q
bfxU3bOj/bP8ehe11CFo+kc4YjcC3KLfYPxC8BauvC/v+23z4QeWI3Xg7qru16PTi2WzM5IP/5nM
pBYGqgt/1PHbxd/OEPv25s9ynf594e0KDM8cVrqmWlPxIgoMNvs1TzgwK+AqBLfkn5pSeUbqHAgd
zjbzT6Nw9NWNZJu5pm4BfQrzbGuhqLhCyaiR9P35gr/2b1WUQtjj/pxDmODt12M3alhf2bpCV63U
TNSRTkZSycK3GjlUvU38i3bssuqpwPgupxgE19DTADzknHUyOPxJXKSDcCPrZ1SkBXHqYI686G56
BzF5EwwgVZvSljf5c6DD7nk/Kjuay3+c7V8BhuUouHqW4PdyK7HHDmqOByrYlNNFuxg5Db25oUtw
WW/0vfkc+zrP7rx8e+Kn9O9lQApxafgFkMcId7A9FHhmpvK6ZC9ik00WWD1MhjWdtrKpAILyZIuT
PXzvcGED3Icp+YjeP2xhwAs4H04vIZ/ymLtM4rTfOV8PcRVDDwi3ZUyquoPFCNTyfuvt+FUljG8W
aSynHj7vEPZmHVQxGZKbo+JZR6+JcazUvJEMMm475jWfQR5THJTxBMAW0o0VcSi4ot+AJ+rMVso9
TRgf6GaEJkHvHC66zlzLefbnqMGAs7tvU+eGmiV96+gym0Y6UYHAa+dxroypTmvUod5EkkQr6U8i
WbbmH3N8eb/CGVKLvxWfNAw3355018JwtY+Ol04DrsS+ArScY+sTLOG0t1XlFHMAxLSE8GaJswTQ
0t6wLl09zFpNo+ClAP94BZtwP9QDG7S/XRUNAVlTNVnnJOwAKSxUbUXxXxeXfptrC+ljfPYndnzf
iW5SFxMlrlLreEdrlyhmDVoFj0xI8WMKH5T12DqP3iZPJ+bUtSyY9NbVKrHf8l7P1qoQsgIVCw4w
SDA+B4tQc18vqCVbp+fbCKaqXHmu1XXvi9OF0VylEsz7ApIYIZyZ3pVblFP2OeYquMfBn6h3/rSu
PfvnjkD1BVjw/CY8TFWBlZWHPDSZhMy2Egi5ANprl71abevC549DRMfWcLLf0MIrCuxdeB1da01W
EmpI71Svy5+lVlE3/stcIwstaNAE3r6L+ucbFf1ujz6HISYI26wL0Hul7PTh2HOd+gFjF849KlaL
82aB/e+Gh0+LuuXzx4jmTv+n3NoVHo75M2r96g++XpIgjdtQ7xFbPAxvuHWQlcDZ1rmN596bwOl6
Ti8fkKP8mwGg+vipZ9YawSlyakO17HUmEHrBfn9eMUOvE/lNW//oI7eodTsEdeji+6BLEg3kDUXk
FLn5VBGVTfOgmSlEi07Uuwf6nYDLu7z1TGcegxnnNcd+8FFpYsoSkFGMAZMa6cRvxO4YFesCikz1
0mXHAFIPlPaDfUulTiS4N/u16LY2/fs8yQFsa9k3we3yF4DOu0b3AM7oR5DKE4Xw1+igx7KhwCSE
1lEBL1TXIchgU2QSabPB5dXE+ojbZ5dSNwA2bhF+EKE7XaXbkq/EQHOsxi5buj82u18GuiyCgyx9
fiFWg+MWcE288qJJOuJGaOQ/oM7OPqfacYQ5JHzmkBA8yQXq7hBYpsXDcztwprtZH/QzFYCbijbu
wOuY2MojwsTTEhxSR220puMRgtyrWGFXcR+reOEKYDRxUfXTqDo30m7dQUhigjnzsCXuTpR1tNxj
SoP/dRx6U9IIng5sOXPnAJiIBjEk5IYWhu6HRJSTlcv1lcVuRmioTkOXnQW8S8KGZ9bQ8b9ZpjoU
W+VtKL0kvrnnzm3xGdJa+lH2QqoHti7a3Wl1V7/SrLARAEj7nFOUbszT0EM1lL+jUBvoGZn2VM1r
S2fW/I1A8j5tzUkZWFxowx2Hd9TwqXEBjEJc0RWPfEEpW3yYuljnCHbVS9g6XyX1urRp21U9X9lA
tcTLZB3dSE53Ilbl1twC/uXke7EkaZzykOWy8fLJQzg8TT3hHg==
`pragma protect end_protected

// 
