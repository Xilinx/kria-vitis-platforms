/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
bc4WnAkqx6dlMsl5fn3cAprcqqxHUHgVY/ImIQQum+cRAB7ouhGGGf7iFZf77q22uZ5IUqV83Quw
Hyk2hoLyHV1tsHXgJxRTk+FG0z8kNO9UiseME5aOM/+f1fcoxpdwoF5Nb9O6O9ouJZW/9wU+cOBn
deDxs8Fe2cl/gc7w+7aUoFn4WojygKnIaeby9NCvgShnH90A/5GxWomjUdPAdBRy04fmF471qpG3
rcDSX8G6arFIKQEh5UwVCLxQIuBK6e0cztUh2ocE1tgu0ybaWCTYOjp5wNkYHxW0TxCBiXthO/Y0
21pIqRWTmcspQgDYTjUBBMfo4xnplJBqhrkXZQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="ASJKkguRF7cNZtn0GfYOwaRh6RbIlcvsA1oAuucVfb8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1110416)
`pragma protect data_block
Xy3DKr6jQ6T4G9Vc1bujRklnf6lsD68FVErHx14F1ZHaBo5PcDbwpU5nGyPad8W6s86m/zkvlaYp
vGU6MSeS07nm1x2uA9sOs4EiVuOKcDohq3JnCZy/QkpbUlGpDibwtULF/94Ipi7IrWyZ5PcKl2T0
Bk0fWHAy0/QvBGmWO2++NLiHLk9GbMSj84IWKLgwDHjpo+L3tFWIiQYyIHnyORJS/Ox1OjLBWkz1
8Sg3bJ9OBhrHyuxxR6b92P8Tzxt7bWuiEH9oj2clCLMrRRgYSX6lr2+JZxRp3EdeRZ7UY4umKL5w
7+Vg57M9oL/Bbd8rjaWaFpQFSxKX6bF208VK1vJuZyRe0U+/a0+r5rWRsRCJX1DB0nthuFisvv5v
f5n8n+WKiCo26jQ26nvy/kqtMU1bm0NNkq14th8oH8KUUHKoGQp6sM9f/a/26U2CERc4GBk9THar
jm32z/z4LRYGcjtmyOVKiUtm9hmCGtd4Nk3efbP11m//gIAwBUVAw/JaUlzqxzTBOxaocRgPQ2Zw
sEe1mzz7lqxUn/OK96HmTkyV/++cgJY5j3MOYG5lUj3xdM7uXPv+/LJzRHh1G6MnkUF8LCGlCaNV
dLflB1E4bHOxGKEXIed9v0ISrRatos6Pxas5MBZ33L50xZLLS6icFVzz5ZvLT6oMEFoe+s0SCkZz
Pk2kF51sZFmDpny75CaXlRBi28LbHt5FetIMwDxEQjO7NGyYYYB0DRpfHQUdzMZ4xOfkD5wwHjcs
fhzNTa/zdmCmj7owG0K5gPGx1TU4mTiVi5IOgAJNiLm9zhUzb9A3HXTIT3x3705/Tl4VZRoherqX
4Vc8L2qr7arcBTtQHvjDmH+oN3cb0DaA7LidE90N8DxWYlv6bSzRlClTEOD5xD0GQIM0JOu6AtmX
3l2oP2yHsph67JGMxWu20s+CBxdUCQS5Wj/lfDvdIzY+0VR7wvybgjpDm4dPZthgXkFiIt/swenN
Wj66+xPvfWjlEET4oGopr7wtKIWYHaBeZqGv9zWJZU7IPcEB3vLXmJBQDwlRGka/IYOIXVd5Aj1k
13WgPiG3vy37jP2M6a11wxPeiU8X/JpHNR4sE6oqQN3lUTLKGhcgc2hFTbtiAnyDWHnpd5EyFD/o
MITLefeb1/9yjtHlvyyQVi+Jlhn6CWBK5gXvyQO2l+hKFENtx47Hd2YRrTUHOKA+kOBXajOHgV1C
Q6+LtJ/DblxHs6spdTN6+fbnc3YhXztNU018kI/Z7rFvO2CJC+1VCKsrGsSEpNavqjmMjIr1eAZk
EsTi+NOjufuQhk1O+suQztzFZ8/DLw4JvdSd2HsjGmwvxxGNDGoZIzJv+50MGc0bRIZdEdqv18Ao
wPJdhF63X0pnrm//9HoriDeravJ3nkYLQDJHFWIdwjuFUvg3blRqMXrgMddFjoe94VJxAWU9SMY3
sHk+KqVPc6xsZk/fnllBjEOWWgqXEsDtj/rQuATIB4Gu+//0HPjm8XSedqHOH1Yo6v8cO95Id5Q+
eQXRU3G51FwovF0WLNqBfDFJcKrv+kVVr04AVDN1kCyQJJUsj1I6v0ZiG6PYXga8qMzzGBDABgIy
cANoAaYhPrnLyqW8FKEYlxv0wuoL8/RwN3zauG3rgraa4FDVgiygKdZxUrinZmwSUwViDn6oniy1
M2v4MDwy9NiCuwD/x3QZaSHDhDFFLJipECXIdwsCr0B4zZ5nQadSm9tBtkjjzMlC3PLzinJPNp/5
XV+/YBp0VEKJEJmOYKzj4k3un/QkfO1RyglEFh8SxXUNvyU1i9n+58+0FGJz/uDy0t73LDzEWBuV
4SIZ6ZUaJYo+EWgfVsQDhalzN+zr5TuHfcjMULert2LuqFIH88ad2DNUz2KNN1AM3sP1eIN2Lbum
9/dGm8ZIUZmNHCeQVJhJKXLBlcUPlik63WsU12VObpmESh/4s2jndBxY+87hklkyg/Fv4qNAWBua
2ZuU3+/I/j3KrjgxV/YJlTGLbvwApBIpw6m4s7y+ronSiJL1E3NfRvXtR685q2wE78mZd39UOTMF
LW7tLPzcb9/qz0jaP1al/MpFRCCJTwegxsuM19mPws9nEWQ4tziP77tUIsWC13mMbo2HxZbkCV9W
hIwEdbwz+7WreUPvm4zV6K2inAV2DtPMlubKTDzjTuPLv3YxYFMQGtPDeulDH9QQ3K9xX7R5lKnv
b9Jqtb1jRjM2q5VMWK59M3hQnWymOEMWjq8Nr0m9FDnYIEQX3X3gWW3pH+w0q0bcSxaAU1cS5nua
RvQDJMfR6fqXUQXjrCeJcvc9nA1XcDSTJ2F3NStle3KnS3Iw8sl3P9EfJgiLNWcmSgh2Zoa8cwoY
GOXXWKTIPvA/7RFlRnpuWL29WuSwt5mYWc/FCirNOqa9Uqbc2VChtvo62IdxnaVA9oPcB3lFxUIJ
LAGV+HVT6HXt6Sedd8jzKfsKQ8RpRbbRj6YbfbY8Q2SOsnBCmdK0TJcXUsqY6Q7o9QE60OFL+sTa
v3AY9ZGK2/pDhRxcVAutIfkPP3HruwWNdJplVqa2gCbXo6K9Wk4UdtWRW8wrlTmQmQl9Y0UYH45u
l6G/ohBiFY0j/7Kqcs9AydAbfnh9/HLiBnJZg4cUF7eK2dhHEHJQuD9VpD2gchX+SfM7pRqgqndG
g+e8jSYC0/RxeDN9nh8pDOuXSw38w5Vd+3ODTa5jsiXaXDXfSFjPq7clio1y1X7JIcu0fdMIZ/j0
nzOOELXwj1pGMAW0Mx2R0V630phA3pmeyMzIukRhSI0yo6DXpT0PXehjw/JXf+6o0rEnq02dekns
FLDRXN+zMOUJcIU+x5uFfEZkowYgJTSNXRnPBoHy8h3G2I0TRmVbLR9RKtjAjoDAvL0GMt3jango
jcHC8A76ID9oMaofXXk/NR8Qyfdw3X7qwGq6PK3QkCAMqotce4NKbuNpgVkx+nnDhAsAzjv20yeq
GHaaC8wRagofmi4l65nurYaHcbvOYSQyT/5iiAEWc/IURTgHhsKtE74x4etTh8JqLJDo8h4d4WFT
/a83cVfWod0gD8CqSI9WSGtUQsLZ7qqCQAYCdfokM1hkJ5/3j+wF7iM5mZmY9mT1opfpdNcHMoE4
i8VWNcEW1Cf2IsYooU3AqayWQFAqg/cm1IJT7cqzm9FGgiAbeHf2M3fF0JfeGKARmkcvo7kJe4HU
hooYIzU25g4APnqKCEUZ9L5iFc4TI0yxWOTTOYdyEfGTW3hdrkVqqdmuvAkCtE78lc+I1QU2x1Mn
OsyUI1OomAweBoFe47Dbvbv14wKTSvfS/PSV3oiCbXSqr7ozvZNIcwujok4L7cGekr9fgV1Qt0AM
oWUZuWrQKBQyeVNVS8nT8GczxqFeab7frgMBzR+bnL8TLiNZxoVtbkR0hY39FRyaPbgsQlwoPTVS
IhxHF/fqL+hI/xvcFfrNvKWKr4QDtWoqVtTCDKYl1IHuAMb9CcI+DhlocVSW+ohK6ueOWxe5/3ui
IJVgt8lfalAwcjsCdel0NWXPg0pFCyuAusdLZgllKyeahavKizzZKLR5qdnuwSqB4VGArfk0aIt1
aSwKW6k5V11oP3Qc40f8x5gDfAQhgMp9pShE1XJuWuW5/zs6Cpx+lBWhDwZrGzyHNzfSE2WI78vF
vzWi0PEugiIIv2PCcsWBinh92q744Hic1EOHhfvpUd+LrBPyKStPLX6VXJuhK4s0WjXHw8hKTmhz
VBxZ0N0Uhd5XRNppxd/oKFOyrFfWE+wSCVIFzJhiU3H+vvCtivMktqdoc1adoOT9Bi7l5viO/v/9
kWbWLN5D8u+88I+1wQRVo6A2KxXXR1iFqXoasaEimUHDFE1JinXGFfUjZHTVr6pBMJIHq4EpF3wX
aDUF/uhNNMFEsPATThpFlzYcdN0VJ9Gkoknkn5cFbCvz2/E39mhop57I40kIwCbbxd9APAqKS4Sk
l2CoUelKxP3KvOdOgntqOeLmnY2AJnU9RU0opk3yiAx4kd95n20KDLQcZdE5spu92xRAuWxs4wye
OQiHPvhCuxmVcL1GpTRweLeMaKUsgUQDPjG689d5re+AY9hgcgkeHnyvk+HoW0AmHVWup6z/FeS0
MPSO1CBpHv9amGv3vCfX/xOzAZ2InEubSTDT/QNDrUuZqUsyQtGEbovn7RmY0xCsrc9wfePsq44L
TJ+H/vObj3FULMSt/RadozkxCW/uyJ0P3AXTsF3ECD+u5SiiQhRIHu5jspiAqWqG/4IdClOntmrH
Hg/vDWFP3f9clCU+O2sxKo2tN3PVdY8hoeChXISzwRBnLs2aldbj1amtc+yFl4xKdfj+3AvUX+ab
7BqKWErAnZfy2FsRfcrh5lTKOZBTYUE5GtnvQohW3hoOKZM3srZY/HMgios1P4bYwO4bICQ2OnMb
JKWeP3cgoOol8KbZhRJ/gKq3M3KUMIa2KMM6sgcSQvTVgB8ncy1zSlmy68M0iytCWLX9TAaeGbTn
44m75aDf/8aS4ewYL61/FdyCLE3Uu0ap84JK25LHfoJeEoU6BZ7DGGmPBUXy4ri7uCERNZN2eZKy
x7123k9E8rQCNM5OwgjB2Am54MNdZhai18KnEbmsnmFT1o9/O8sjrJpgMPSp5RYj9fHYVkjcnyI+
iaJnuw9B7D2RbsXgjzBinufinEdykomTPpLUTS0yzcmVIwkf2ElujLq+XGuM2VF14lRkXVM6af6q
J3M9MWcb980JO7/ZEky6BKWYTDCJyVQTN9yQN+yaoFSUn96YopyB/fg+RrelZumHFW5Ukttn7hdg
fVqc9GxHLy4Rzy19s8i4t9+3hq2kT6w/eaCy8Yh6MW5WFigcnFC1DJURTq1fFNqnsAtM/EQsECXS
Mmw9XmwlUfXNeN5rQBLZfRk61dtWKY2u8h13iN62My+4xLtnoSlQN5QoS4UEa+Q3Nh17OZfjSIcn
s3D3msLl7ZBHfmyLG/0j0G/HmsSItS0qD35zC5wXfqSHpdybTT1exW0yeqxZq9tDV6g/XU1QmORK
UtkFEMrN2dpb0FlSiBUvnOlaPQWl/8rFQFpzM4sbFcXQW4NsjG9FTUrYf9EMhNJTbf/OF6tN6PwW
9Mt7yN9vzyyqp6FJ1GrtZhzaZIK8kEUx7PlTJ1j3VE2MbVatLroAGzUU7qwxB4gP6k9Za+NH3soj
AryzndZlgXXuLbaz64kTc6Fx84hAAE1m+a7BkfxRNcBO+32+foN/2ERuOteeFqUs1H8vTfmXmlek
H5+USCI2EflxjxIDfMKgVQaI6l6YOtuQG/JBJyorKaM2/qWvKC+L4pICNysVkvTx4wFc8TCi2jYw
uU3PawNl/FjbJYvYKbGOnQGm1CJlF9Aq1v7o8gLZo51ZmdTMu1ccecXohNiyD4vwNlMPEuxo4/Wg
hwCrxUuS7azZmftY9zdGl1oBeD45oS/FjH1Ygo6au54xZze+Ijic7QT7sFlIctq25lxUgupHMVjC
SqhxOFrnsYwPE+VAGw8kNF8+cl25goURkoHojGQ/Z+JE2+9laLihqt343DergLBBYFHwaRUQcANb
OmTwZzn8B5d/ISYbU/wVVOao7iv3xqSSAbiqxqkRxowdcBpus0p0BYrtspxGFYoLceOlzJihUxLb
RZNRcwuhBKZ7PMT8rrs/hl3l+HTdsUzMRNK0KEIvbgVHelF+2dj0S4h3rBrLmiMUVfY50vOPBBnz
2oannISaIKjy5/5Qpv2/7lvUiRAW989z5SA62GGrcxqEzow2CXOiyqrekKbcYN10/XN/2m3xaJup
ws0gHIWmA6cxeIzgtFsbBUQ3RunWamazFWkABm4LYFcYy+aZJw9aeCqvtzj1YVn/Pl9xAtUexQPm
CG0Q+hU0wkVrLD2CX4aQXFeR+Ch8wX9VBM7+kMOHrwjT8vMa+saeCMeAMBYgWFDrzWALb3vMxxuB
Q2jet6RbxwYFA4xTm2YPtPoQRGibNxWiGBImvZEQQamSyHO5bVzgkgUEop6vtthMuymBqSIkzdC6
4TtDKpP9qBUM3Vtd4j8eOf6ihC1E2cU/IqPfEGR792tFR3ALHOrtaqGPoaJwovdH+G4IFxlr9aqa
lyIv3QguIr7iLDdvRP/bqR5s7RaTbToxY2FZisBVHidQBiEPULMq7ULCI0MJaIMpZUDpkPx1WSNd
ppwpANBLTnrSpJVJp5/p86RPTCB6e3v1WEP2b8r5+YylKipQN87YDsEtYqLsRl2mEStlcS48Zf//
8yRahFBBMOSSsF+HpLH2+bsVjpqhzsfQOyaRBDpPt0pqmdAPgR4ipK0JG+2pNZd3S/az/KCzEr5i
biQzFK+AH4i9q2VapHuvWxGeGE+1HOR0iAkGRiezob44tc/sbAtamuyNgjNaC/qi/KcKyEsBmENU
nqXozztnALqXicv43ePvinRA3VB/e0J7OEEKQjkDQcWIswIllnWirjFaxm/+XMwkw75c1lANYvRk
Q/WFLndpVWiWrwt/rNOuBEhaC/tGKS+XlUVk3W7oeGqSe3NK7SeY6lgfKh6WuvJ8dq1V7XMDlxiN
jvRYbCvwjlKR0XsJMIa7cKHluD/+Bnjdr/w6/5pxjJ9b3JFdMd8czXrKT0R58/Bqm8HmmV8kTIqV
cUsqLXKzEcmz/YNAdjHiEpecbBy+W+9l1elQviH4UEk+grcsBbMdPWmawIBvHSUB8xUPignSqm1p
AL7l4onRRhth90EIDN0+BlK4MEQPx7zaJP6nG82U9avxZhyJ4/TOhkuEtIlplrfeoFIVd5KB+Hqa
Ji2AVftZposWkJEbtoO148FMeNTtVFiTJRvpoEoSxP/7ezpxFT64tR9B6DGCHcpgVuTtTVVodCL2
v5U5dhaF2qQRQgvFUPV/G9jXLMYSOpZCcAUjLwaDFR0p0FCiS6+mBl3n7KNx8sPQPYh67511OgAb
DFk1R5ftLxyf0SMxjo+cHoR8/dQA5j3N60MraGAOPqKKMJp6sVgR7r8YdPW4P1cztSp6HhK97Jb6
z15cGhG3mNtO5yeYOh3fsUuyurgmETNj4Vf3fNCmTZRWweRI98PfRZY/rY/ht9ob0BDICkxrjNHf
wKDJPU72h+ySgbf8r7dAG2MS/E5vyQq9Q2X3e5wUOhyEq5d6kaFfZnbpP5D2jzayJUpW8D6/8MRV
YLbzAkWkrXXQ1lsGHGPycSY4/Wl56d/wDslmhvUdTfyNn79NxM6NHv9QbY02cpzWWu7XHGYhq+hw
ttwjiJeUjmlu7277TTtCEHapBSF7/uuoRnhQzGijR9jc0lHRYTgCOPJGcb9vwXCNpii3YvG+LVYw
W9sz0Buv7cItoYEkKL6ixRsG1APV3E1F0rDd7anz/2hsV6Att5RlNY3QuBtoYnNYD083S5+xbcGy
+xqD3S9gRsVuZaHllBLRPG7czp926FoHo7xPHkBEojntmLewY5EaNQsqWfecrxfSa/l0+RTnQceZ
Tppo0KEe3pJdYaW9TCmsJ/1Jw+gONPE7P2Kn43ejR2Nh5ySmgaeWHsUrtZt7jq1HIWujN6ILHr9X
5GvACXgdoIB+D5BCRKJWikxPZianHhKk6cCqxGG9NFvSdlk/LFW6+zs+of0tGHVA+4PadsueP/Om
455XdiprSh6VjkOonNT8giBsWT9CaqR3Jj3aQPuk0kZkv/OHyeQhrk1CHLoDb4h9KUHb7G3nLPLN
5zs0LfHPtzeVdXol3wqscqB+A8SVMHMLjYyuzLF11YwwKuC27YdSfLEW6UtH5IuGEa1CddNlR/2C
Yr2rsUedUbDMYz7KvhdzPekkKsryQtkq8vU+sL9PuhOxNjQNDBVo9fIWTUpf4ZRUe14UrcftcJZz
C/LtcGOOojSidjM/GuvUzR9qk9ImFrNwuugaHmNjMr8DfrF06SoK4BxULVFcYVN12jQMxutT0jEb
YsNTsbHZyaLVVCKbV4044PXL3odXxjEJ7sTkUguNEZvu4YZKWvHZGNgUkxlAqCjd3L+TTHlEiFlv
83LisRe4UdjX+w+aWMM1OV21yjtdxV1t8/Ukr03Nfra9lgmH+xO1kXu66tCFANfS9lPyBtOhUeN3
bCVDWHJyX2DiKkGOjzlAI1nwh2ncPxn9sUWFu7MYPBqobnyJ2KqY/YeNxoRLFXl9G8DzQneRNGs9
0al1WLKx8Yfsow+ROl79FLD8cmj5zT9zvn9zj12B5kHailsIr2BPamPlwHLvAJh+dLhhXGm7k3na
SfhwlWW9XeLIXLOilrmJcWmKRGZk3n0HTT+hQ0MPXA3RkZIPLZSQwkF+jWWQxBBzC8y6BCQh/6Cw
bDFOxl9a2XiVZuPFF6aewpMMFE40GuzCuSoFZgn1lalgqMacN2I01aRB1s14sKCr0oB4peit6Pba
57PyAZereiWYOrxRXCed/i2A55Ix+JpudBtRewi/vLf9iAa7EiT4CR7KYdXCVznJNlZjZD4ka9Bv
nA7VqAOZLHLVxDlI8JHKur09aSiX4cMhV0GNLJOVMTnYRe98SZuVIuh+1lXEmeSRe8E88GA/D8R7
DKX1q3IEUfBW0Z0LHtMtI95LlWDEIVYk7v5MMdaXpBdus+60XHv530U/nlnG6QaVizuYU+l0HCuk
bNCYN7IR/tDaKcXYB8dpuv0+8nv15kiZaqTnXCQKosCZmDMiLs8mDvvJmxu8ZEWnJJMMy/YfBFOc
xTJbf4T+kl5qRgGRoY6SEgfSPtKktbmLAtqyjcMqp6148Qok+kz1B9YS/WDBOHh03BR0kiMi6o1w
XBDuRLIHHimzj0tZGYYLbZPuvsd22BJu/HfwwV1F5qCo/IS6Ndo0GQgDU9OCDfNSe16JWrNCnLnb
QhlNYRkQ+qHI1f3OmKxtrCyefD8dqa8pwORQCF+RWeHy1SpgI6s5KawmLvJyahIFWo5URbzodI7u
/0Nq84aAJbNek+AxL40uGC5UYdDnYX9v4s546VnhdhDoM1zkh+g8nsneo7hkUUvIxKaSjjCUAq8q
L3zBRO+LHz3eRvCrcKMrETFKBxUcEIUBtfWVTh4o5gMsHWxg/CQqVWWf1KeTWGcjGO7RHfqUl07u
R2N8LMFvJ//MBikZtYmhBDYbntM6gTJd/LRCoXBx2eeboQIF1Ih6da2p26N528fQy8z/xkOiPPPf
zMycd41sQq6pp6/ZhZnSBW8Xu4FE0zxWTOU9TRzVGhHlQvZzP7OiUnTraliJgpGFe6b57VgSg/0v
D/g1JWmLyIxSzRAZLF8dPBtHekEoBGjQNk9PcgG01VMiw7KqH31VN1GbG6kEKL5cX/ansLW4BCYv
wpDhtePQekO0VrN4fDMmQ1H17LyEO52YU0tDy5cHkeRMII+QwUGnm8g0ij0dmek8iEXfXVHazMiW
qqFhm0ya7/9LCNP/NFZ/5EcOp8ZgqJJaLDqDkQ2YHgyQ6O5TSTRKHNMnLmObRnwCNSdL437VdJxJ
92pcIgovkpvCo7d+l5lzxS7WYzXxl9u+n+wqi3R2u8O3RWrohQ5tySHZ7kFkngYOMrZZ/5ony23m
OvwQ5IoaYHQnmZBXdLSZzTNVXVeGfXBcgnS5iPuSEUJiu6D2AFFBpHCIC4ezgh2uxfHRxtBL5gYu
1kPhXTLGxq89BFk2HjmWzKY9CxikR0Jo3rh1ZrrbYvJ3bda4KmmdEJBewyDj0GTldEZCsndxfkvM
rZexKExXIOnQWv9D3R252+qABuvb2rYCjPEJVV5UQ/U9WMBHaywWlrQtHptmh+McXsL63SRVUCpu
8YCrxCOoKvhECwoaRRw2ei2ayhGP+Om/RfGwWQw3iNH40v5WMKXgb5hC0GHBKKtZyHwqrh7/78qB
NUsydVBxtgg8kZ4fJH0rS82yDZi5RvLgXWqeEZlyQEmkElH+A1O8mY2GFJtOcuY1BGvCW9Q0ZA4l
RvAyHga1EKP/qQ6hXr2OqDGKKcyNZ8h5a4McAcLB8Dezb7QVi6KHliuil4ifXU5VJKg4kK7DAtHJ
OJHR9VprsXYQE4SOYoGHZ/jefQ5mn2jJItzFTFfX/Aj2Y/zOY2tqdc1umYmTyzZ2zma5WfLptWVu
U0VTB2T9GZL789TXxFe60FSobWXn9Vk53C+AiV5HC46EmEsbyAcIgUsOc1g/fJeY75JBz9KG0lxW
TjpkXN0iNSwTap/SEs2os5U1ZABgROKBOMv3ogXL+fggbTQdGu12c6Jhi59MByUgncigvQNY7SbC
hXZn/A2FTFBTbEeSryAjEBsOOb1E+k1rpB6Io3uxU8V+bdBvfMiiOw0loj2PEPGQy5HzXn0EXFcv
Ua7gH1bFBiIuq8pqXntN8rZRh/g2TRDe0ldny5sjE+19klNCc6wSM2pRL6mEbvlvITLZWTQlVlZ+
Imw6pn+xvcUQfAHyKa63X+fltl98jP/4IsL6ZK0Br5WXF9ABlVoEP4UKTgFNUQs2e5j+Thfk1hyM
jY3WV8TZ4wrymuD3hs5jFUav0ENBFc9jUEOADFdJ+HMEj4LJDPeghWmsl8o3qEIkpmnOrWM4gKcI
PoF5V0Oj9WYCDnTR8naRRIs6XMKWRq6l5N+Q3CJvA5i/VCeFRvMZI36Vs2XaVanIvQEcmHagkMm6
LrpRPhgivr1Tz0QGlvfk9TUr6Yiqk/dB/to04mkznjS3pWeho/6W+2ZM04zTf3TXTKSzcc2v7yAq
TY4+9U10JqW3wsM5FI2RchOWrN3pN8amVgfDmlU6oPaBazXgZFnztYZ0SFYSj8bF8uA4hKV4coXD
0ZYdnGtdanzFQOo35UFzLDmZ+o+Ia0XUXZ/4/Tl5Ghe5dunSteBxy0fWWtitSnkOFfTHi8fjw3kc
U3ajxvoPWj30Z2dP/UMYMnTBFLmDU7K+OiRoW2bAo52G05hBd6VzJCD00H84qveY3tI/g41lSgI8
4WdN/9SnKswLDwT2QXoDnKuhMcDMzegnnPelGI5XLPZH/5xbpw5EYlzFHIBSyu3NrNtVFo8NtX4O
VYyWXzI/rhkA0e88u+0rOZZTnvVvqW3PW9KIlSkU9gB7kLksPDSJvjcnLiTe144z8qdrvqt/n5gY
z6+fX0+V+M5uBpN72H6vIwEp150FuinFfIIqfAE0QU5P305itgsI4+XayKFRV69WTGdtWaiZIyeL
hFk0z52E1WeSJA4xa3aoA7kmNCkJ+88t+OxIvEfCn2T/Fp5vt2Om7IfbntaNBEU1tPoP4CbcffK1
fYU/PbR5uTQ/eJ8ggFrpXFP/ozr3aH0DlcPKJgZql+NIBQr+OHPSDwGoqQozvgbuBcY3HA6H90Ac
vEJ31C5o2yHJ7ibRVpNIE/ionVur884SwrmVHrHuVKG3LpDBpdmB37rJeUEcdVMoaUaHHQfB2CR0
V9bDX3FqAPTnRcqr7a3LHv+mhMFn4M/XAPGm8OwSR6fCMtTYLEk965BR/oXCG1tKp8YAs/W6s0eI
RL48gG7n2JP2dFjQUtZsuh6h86lMGw6dc0F3xNonNgXUK4NvoH0B8dR7/Li5g9ku8eoWpR/YlBQK
I7FikpTGGNHnGgJx6jGx2HvOFM9K7iUwB4pVF6jJpgftAK2RKYD5WLIm+jOUgLXxzSYeObwKS6LH
3hM25iiD/YGdXP6EY7vZvLmwwhGT9pGchcPF0lm2AIEXRUhwFNAG94xyh4D9Jto/cjMLl3ifYvyz
afiWefwsD99gCxYaumWj5CVT4Ab3N/+NvIQkmF8GqzUy2nv2kY2Kp7T4QmVX4CM3sIKACQ30CR5z
mO2eWdyPvqZEnchYuMNHF/3KDEyQt1KZjw/xp8UwAqUDrhUoTaZmwUdV17vbJ5mgIQNA1K2gB/HY
WAPTI44toHVOyJLxKMzVXm6qNfJ5TnJvljE4L+u2qU1D+3QhoQTlAeXad2lNw8NBgi6e2Ws+Z0P1
5bI3W062Ca8YhZu+h5PSUW0Jtz2yExY4rbfUhEsZ1L3BSDneNSMEiPwZhWuxsDp0EnyZmxNyjgFI
MEqUS1HsbVKBMZ3y2/MW3mN30sG/hoMKq0GId7rF0SFCxPfX65MN+kzQgGh+7IAGrqIC6+f6izGF
Yh6xQTPvqvlzw2cseyGUeX7j6C0xnEpCB18iKUf+MfC/JWU01M2Issls4dBBjZ4iyAC6vasbeXY+
CAdobddX0+bP6WrfBlIwSY1vTF28P9YO+E5+sNCSMwHcilPILSroA1i5FJ+Hm2oF653Ctv9FM38e
PertBoFPSXWnVzRiZFU9SEFdl06KY+M3pYzdMJOdB874ytQC27dd0ltmXRHSFifYshoxx3Zgpdz8
CzDDdNP0eR1n5gbWXjm1HUB+Jqn4UbMtBMhMymhfzWGJASuIOEsPQ5aRX6ebteCD8jlbSh78ioe9
gVtpQfV9h/2kgBTUc45Kon/G6wYZOtOjIrsj6VgxrYCOeTCu2WgQRtHdzuH4cBWO8ELpFC/rij7l
zwNGjeNAGMmjzR/wbg2fYpnql8v9NwFf/6JkxcomJ0iaHYx7dsvDAvxxvuGQaafKdAinLYW0/ROO
LpcyKNSEKKwJ6PaLpfMVJ0ccaghNQMKbWQgqbz4zok2nFpW/CWli5ig6d9G5QscTjNgHVbwhC1wp
UqR4DRjdBVPGuTSBYhFgcdxY69j73B5tR9opZxOAnfEzBvUQMHjt9QvQKHA7lpUXK6swsN4ovUV6
LtH6uBBRhKINa0ORcTkUnzqJ+l0Upb2T251dUCbv80PTfTWsUvizrpsM284/LPSzZKw/8uTkALQo
ZLkWbgy1DPVMMZ/EHkO1YFJZAbMEOxmX64AIzKlC6SpfVISoE9BpSuMYaZz5MmMtLdorx/PpVF1N
kGZF7slQuTFMja/7QODuvYy7GdIMezHOJJ4wgofOuKp1K/ugjEmrkwjrdji+qg/mi/nD8gxGh3ig
D9nI3yRsmYgWQQGZ4+AoagDVtqcJBFs2h7xYlbuaUfyMa6GgJsL7jMXzrCagM3VPj6Cl9E1BIyzz
YwWKwvLqkNAtTaqONy4ww4yyqQ4UR33+e7OmNPrCuxD2cHJLgT9vJ8P6Udx4+WmvJAf3yKNWtE7n
Xi+mmpbwEI388ezuFyegFKuNYX8EGxr1OmZuTwdyzWffPiMFM6R+WZTfEyZ3RvGXa1nYG5XnTFBF
u8ABzQ+cBiRRKO0DGJ+Wxv/nGbyS7tGS2oUaChfKfhQ/Jv9ROOQdUBbvqG+b3Fk5NpkuxV0m20Fu
4kYx/JQYTPQgZPHU3DiYmeBcoVAICbWYGLLsmip0AtnKXWqrQxhT7lQvU7h4TeugvgdU9XE1IkRT
Q3P32tZpPuQ0mBfLE2xEKKqO+0TBhpb+vYDPW/cJyy78vSc9SZE7Gym+4dX1jZxHZ1vYmB2DyJmY
vdOw/Hd9NaYpCMIsdC2wViT+I6as+NIQQtUbvBCROvEd6al+oKu0erfIzAnEH0aJyz0Z/w33IQZn
sX8uKhY7yDKn12Nr/LnVnZ5xcOeJgy6sWfRLHPte5BxICWCWOU9Pil9xKnWL9+JBEP1ejAzUzhPn
3oGFTCvVEKYVs7fSz1n6uYLrMANRtOYMB3EaHdyGmlnQSKONaGNy9MWrKj9yp9FMRY61PtkrjBGk
E1QMhXQ17Ja3LpbowmcOxXaXNd0JlXfxxcKFIlbbnE5LsE8ps1F5xgSbkcL+vZnWWBVDImPUZmNQ
xKh3cOZcBQ2GW9yKGoczmKWluwpVFxTHVBeZAm9pVJb5UYX1iwOYAPH5bqbWc+CbltNvlTHTesjT
Fb1c7e/7jjVUvj7XdruIGFOwa+BAgpHqJjEw1MouGrVSWekIEQdckXrCwktGirzTKC9bfJAl+LBR
aUCDKUqDQ8lqocbbhsCAMvgvsRPRLH0k/yRZWVBZx8NFuXzkgoSl2bdISo+uSw+elQevnMIg5LoK
337IxaN2v01W7iMwSYSUmtHLMTsM0GtZ7XZ9eNPC9GOz6zj7sun2y64gvoEe3t9pdLiptGduCzJ+
Z/dBvfWD8DZ1+Va9b9x8RuXzlrEnKDfhHFhzOjFj29Acqn75WNOr23P3U4yxatrfejJkJ6H1Zamz
AxSnPpJWW/7kKJKTnSU5Pa5ajVieYMb8drP8wvrJ70ul5QjrHytJDfMA73+wq/rXOcAwE+SgzKX/
doo3yqsfU765iUlhc6thi6c9nXOdWpu8JINE6UjEItfYe3FDzIDDccoPAa0tzTqlCyi4R0m/YOeU
mXNXEf0xE6US26TlvgkOGNIK6SqV/FBLWYQ+q+tE4jcmhUUuoN0TrDJlqNGWfG6IHja1Vml2vx+c
41DA9F/FWF9PJhoXtUk0BLWx1uQLCJBfR5v/GqniCWgSzQghJK9MI+HdFrf03q6pgCPXbhITSu7d
Z4TV0WDFtEoJjlJXolrVDvRo5W3B8zxLqkAFiO9N/dtKI4IS6E6kQDC5mIUCWo/0z4xYK0zOxZEQ
IAWfyHB8r+ZqaS6ff8HGkXgdnm13JIgK4zus5nSCFBmg2gfGM3v+P5HqyJgOu1baHmjYGdIqvh/9
hcj9jfOkz9tUuSioolyMxuBf9chLj2T6Lond5nfiafdruXgpbtMSxc/Y1hx96rSgLM+Jgp+U2JLF
6vpj8avc5SMKO4eMCh00dehcxPjbK5IetFK85kmRAno4M05a0R6PH0LoySeOA3ktPcbno99o6tLu
CYyH6aBcSbBtGJyUfPZSlYi1GOcaRWiTdTk4CWnh2uVNZfJRpkqXaQ20JCRIrmrzfCMpIqatUfGU
UrAxxJZ57HUCHfZSXBHhfGtzl4u9sdEs1UTJhN2MRj82dp0vP+OJ5Lg9H1ycg4yD3BuYTuYtdmBj
oOXMtuVw8wQeI9kxWo4LO6TW5N4a/ZNl3HHU4n5i5N2ryv7uphGy88KqoavgYGw4XewKOh0FypU6
tyJ3FDNMpakAkX4rGKNPtI0fkkLPJzSCrF9rr0gV4OGlyNucewOOd9/mJM/OMejYAdDWQyjb1tXi
MeKCjR/OPPdUuDu/XYxLrYA1NFW84rjqI9RAc6SL39sfnj2fgG1pGlCvqju6L2PVOtRPYgVgKlom
Cg1oAPwpu0dsAA0h7BnF4RKe2qLcROlWNDFdT8u+Zbdze9N6I9uduWCwxgYMF+Q3XO9S3KsPv0z4
U9iZXRd0XYTgI1Ro2Hmn5v2JcoWT9VwHGf/7kx6ZuQL5ZgtcQMUD9tC4BPH6hd9QofStqfHYYnmh
Szq5MGJZidRfRaZtFRpCeITNGQgTYhWxuowAGtv9RDqwSHFqJTVH59/znuzGuVVzlTnVXxstoKvM
6zTRUdI7oYj53D8gyWoxQbcgtW0a/kQ+k7JY2OQOM1HeupFAT6N2JB7m/KBjewr5QUABd4H1K4z+
i6ZElZHFXWb7DSNCprcZt7vnlEmqZZznmalh2/2wBTfn7UsGKxPYz865nuKnIgmlLCufFHejPQIi
SuZtgfmG/dOVRXrdNkXREhIswtXQS5WpQBxBOXVEc8lUjw4TZTy9z5G994OfEdjR6c/+W1gfrqAj
r2E3X2UnNt/1nVAdl75DIVjRw8HgtKquqF5TqYqBPwcuzIea4ALOwukPimpGCKEAtlmaJmE+lQlR
ov/COZi4QAO6MjgeKZezh66HB3FTgXUtJ+kESZwWUFsjnU4lEMJbz++bNNPy0ned5L0I+2OKsPbP
LL2bM4CWKfY/f7RVeU1ufA6SMSiCOG0SfoKbVOAsGEZV0f28tOmQh0jrhXV6vRrKmjyNoZnU5TS4
TK+MBtSykGacfIv02RfpTQLGJosGNy5TYDuPfQ5Fqn1rLKPumXA7ctKRuQjgqnLWukKs0BRLOhBg
ThmCidBwOiCuI2or8H+uP3CoRN87T+QOzy52mVytXoRG9cHJQ1X6V+tVlSu70C0m7hx0HU3JUZ1O
L0SRUHb1esNrvsES+Isn5wsAagqgVmVz8ZZ2ckISJsFn+4gzijb1ZyvaFtUtBtD8X0kW7xujFPej
YVUFpUmnUM5YtfjNVdxhlQN38g4q5hm3aW7RSR2Ug1lrwYdrHxo24X7NxozEYjrG1bgv4NrqJUQN
DAFqj8AChT2cvhEoHuwR4wBi45PSRGQzuwTDKbDjL1W1eQzegWuf+2wvAMkqiq9G78pzVGPTOMV0
kplCe2ONRFu2Jfs+CeHGPbdKiJiJwGMEJsZULnBEO8OSEOAS9AonrPEvXf0A6ZUrDh2CqtZXbqY1
JKoJDxRr1OVzwrT5aWwckspMiNiXNSovn4/SzhZOoLifjUr8GNIB8A6wAMfA/qY5dPvgnT2qMNmK
8X8wnIIC9uNm4LWl7oSfM0xBXlyE2tweJsL6jnwY7t8SUEHlPAIScbOhw55QTL4pzveJigtDwny1
EBUf+P2S0Y2up0JXLf9JBXIv3ZD3kw+RqXcfMgnNzrv58XQv1T9BZK98mjy31jnbjvN2Xm2rDIlz
mkzaaoUcsuD4/NabhLfj/A2ODw5XSPHrLmppANNDTtG0Qc/BrdvixFX/8yyKyxrYmaPexPrViEb9
8dXDqo96RIlzsrQKpGVgGgd7zThxBV0DbGRwP3CKUPSSiSHMv3q9lGDNco+bCrXridDyeXWhJjHw
5A+ZF2d0cZEJRsjvcK+j9WqBTMB3FZ12W9cw67CIVrkz0M3mAZNNePIHXfJxdMif7u7lQgwyetqg
1ywQ0ILULrP0Z/4zpq/fFMSDoTkj4XJCPAM8H5UCaipvbwDdiMh29R1E38fEmGdXea/wXJkfkCwO
eL+WVXtbXgwU1yGvjRjbgJ6b/GAc078gC0oFdW5Uy5TDZQs1693mYSVWJqrIQchYnohaNp4ZDSbZ
mnH0nI+hO/FCtUyNdD6dAHUjPLzIFJjJ7HCX81MLJypnwhY2sPSmUs27rSy3rsVb8pQRruPHFBkv
argtPSC8LI30Ub1nYsvbRRR9aAoqeXF9Yqn4pgDeLSK9v41mkPAGjqdOKCzbt7a+yHM16H9pjmUn
M1wWIY85H8nbUYkifv2t4z7ytzeaAVzYuUoN1wyh31/er9VPWBKw1HP2nHPwj4pK4C59d9CiUCzr
o+jTVipAmLKT/jtO0SkopfsO1WUlsnhyh16XkXrMgeHk0x0IytToak8rYveDyuxae1+nfAAvqm6y
Frspf8IEBNyLygCgIOCCkwL1gvEXcQhaPOyX5Nk7+y3EeqqMQ3flsYc8qD2qCgYqLPh+yoO2G32O
GzUkUMq4fRLEPo73y0pAjG1clnx646UVry5ND/AY8Hq3KaDDx4faeQT0eeaHTtmWjFTPOydA6V8C
Wcy++8i6DOYtuFfIh2MLthAPvaq8hp+sz7BYlOvMrh1BDoFESCcvFiySae+TXVqp5hgI3bHhlKDB
/w14S3yP4Y1R0M030XPeCawjswOPQD0k63fDD8T3FTxsC9SDkzRlkiVH+n6f4I5Uo7NGx2GH19zP
aUYCO9jj9fJJmkx7lTTLEWykc6s2cZdpihMwQa/o3qatzarDai3S6km7hgN++CMun0vwrVVKXokE
cKMurhPq8niUuytWCtg/U1Hmc+ZHBDhuhvtfJd3FophLV3/bKBNwesoNo/qLHggKKNuPEkWUy7KB
a4lEQNLlX6lkru6ZyDzx3VUGzIjpb8qwH7iwGtzhTSHsN1YVscAIq//+DJsAJdYxpEIrHQwiV7t3
PIKuiI3BKP0d+iIaUwAkowa2wz97sCKKO0+DdI2xEbynyt97M3/g3HRD7eAZ6E2Zy79OBsvm5XaM
KB+EV9kta4S1w8hSvgE0TKEuvh/WAOCgPUKpPzuuQ6X0Y4T1Jqi46f9LT+BrewRSHki/ueUgRpuc
QSZmqeujGzLj3zcThiOh3cN2bLPpiIIsIK+uucpKBDWfDfjHGhI0OGhtFhTsf8JM3yG4ozZvN2ad
t6Gbu1ht53pF6pVYYxJMh+4IhkMJWSJ4uHXMkTvSELbOxxFbSR4FtNx6ELP1KCvv2BCg6cOjM8e7
mA+mJKPOYHxpE08PqwLWyUJpPfzlIqZFMnjwoa4959peBn9VgpE3mleTGTdySaCWXcMa7SfY7gq1
0ZlE/dXo3YD2YBw+cjkVh2FTWhkaiBGltkchbDvuIdu8XvHXhkmb29gCQ+cls0IVOoB0iyFdIIvJ
9GTa9RZfMuOsAKhm/H1iiFy2KFea/yb3THgO07+zIgIQbaerzVySDAen21IFujfXtIzWPwO8Ie5n
EO9T8Z9T+4O6x3WQUBXqJBx2cnnw5JUZrKiGGFQJsdjY98sOsIa4D7K8vhHWDfh9uOLI3iN6jo3o
uKmVjM1Rv3mMrBXPxSbYrCnpGC0hjaaGLZDHzMxLv1pHaRILubL8p4rKTzd99vlvZvCKn/JUIyCN
CfzK3uJKquq36D92QGItux8Wef+9jMUrVEsCPwJMYsH4xVd4LoDg5u2vCXB9eqcoJsuB2nZtIZ/i
4+NjTMJHztgljiMF8OMXkovFJh5q2LjVCkrGO+NfNsj9IMvJ5uF+lVhOPXg4oykRFdSLe7dF55D0
aD56pJX5JKWfAalckUiDgQhFugb5fqvbU+SZwhyLHHNNvqCgswWcZC7rg6ox9Fg0rQGw0mDOwIQk
rxHZH1KdbMJkEzo9XdxCbEZbW11cI9lrX++wp+1rMKRAsX799dSS3r6p5Vcip8798scR/UZYSBMI
HFQ0ggvJW8/89or6B5+casDFqxn+mlAbqMS57h6EgPT+5tZ7yUvSRzL5R40zhqcWivTGom4yakLn
pt6KUJhRsjS9uiZt6KZp1lmAvZ87Z8L1tUqBhUGHz7TxlzpGynTJtvbKH2entCdXq4lmStC2lm3M
nE5ZNu/1wbRVvhWzMEDb3tqq44dmFuuSeVduUHr4zx6eRvr0a+NNTv/xbYECdoL70WjPzCM8t+jG
Zg3JKVxySSs1b572UdKvhOmzGuNgbDhvEUq5DfaPYhLsWDFR/j85wFcBMFxMJOBF7MS4sHokiZOX
He3/JONx0Gk3Ef0uEC7Is8GBUm3VdeHA8y8ylHEIroirMqbeZbZZmYJ/jg7rzt0fBv60YsT/yW+W
64zKo+g6UiF5ibtJfiVfrHi7M835mrTetgiZrn0HBXMBOboJ8+ESORG0M72H5yk9tTRuHuymB+4U
gFOBsDDDGa+wbIGMSWb887daXCAVQAkiKWsSvWqOeLIjoAswMqAHc/ooSpaYrGQ5jiUAtM+j6SpU
dZW37rqNwlE8XXl5wa7DQIFqK6rakYgB03oqgG24tbW7oEgTq6crDqp/ixOunqOV5ZyK361FbBBr
l+IwZTC0s/cE3x/8KWM4WJdVJxWQvVoclv1SkAE8hVROmqRBIhcLZUCnu/VXxqdHSIoMLFji4W9X
Q7l6AaJBUvCRN2UdztMDbed7Ko3l4s1rnMIvpktVR9cNlBmGNYNAAWCyZjM26TqDy5KaUqqDUHFu
ig/HvRs9pdWG59cMjkzJPIr2Oy9fNTI/k3G+9J0ZV17ExWKykvCKQFVmG7hWVZ6Eu/XA5nE+Vedl
S6z8WqsbabSd4KNFd7X9JiMc8DKzLdQlfOp8RYcTKRTZxwcsnBfXnJheA40OFd4EwQGbe7KQrIdg
8ECPhxY20HIE5YrWDrFUukUwvT7hpVky0a2cTK1vbbttJJRtcdmMHaRgAZBinJ11PbX9HxiuXHlA
9fJGbbrmSZu+ojRk53tYFK7kwXag3+56IHa7mGo2KZEjOfdv4Yd8uL+J3EE4Ky3KW0roSgiu5Guv
Ls/OYqqeFxhiSlENbB5IJ+HGS7qXtmnnepPa1IxObUHsacYaAPY9jdeA3sXf6jCgy1pjcjHyu39S
oL803FEmo3o8yl3oqNrdGRhTQP+5hRNbKloYZ7+LESmW0290Y/c/Y3XU5yAsiVcLYi8EvGcm2oc/
ybliqkoq/RyWTcZXr7V1G52HQ54X25r3rcF9uMKLVkw0dG+wj502P89oeTxsjGeqUKRZOcOG7uRp
5T6QIEi0DthnZY14ZI7w3O3cclnsQRidP9g1BeVbptTAK62wArw16RF5zA4isR2sHVRkbA1/bKdD
lgrWD0xsBuSQy+h5e+EKye8EcMvB7oQMEV00NcVlZGfcWldlAg8eM2cUV69kAdxzeap41YiBoJx8
TNhGG8DzsiQVrRoIIpBzODko6hers+lh8bjjTNDu5IK4gXAQtVzIMq2Je6GZmmqI+0HBNUCU2j+t
ubQ5GY9VSfV4OvL6qcCl1e7IB9Pzj6uw7rgsQhykDLZpH18PTqtSg59Pr30+pqeaxXxqH1Q3vwGK
+03xTkuBUdZo0dGzQVtNWb/vTvhd69IKY3srQ0Zx0F7arRGCu5qqQk3SuaztzXiBqQOXDAlTI2Qb
DmCEqIHqXFxh56YBkjUZWNEgBQHFp1D21aeHeF2lB/SKsPXow2d9c4WojNY4DYiX9b8fGfmO61zK
4XdsJfRLYkZu13eCopzuL+kd74UwSYZDYwWxWPjRkwO6SJcyE71fUlY8TYWjNQxjVwZJ04GiwYaH
FFO+ZXrudwPzAdh1RK532guJ0BEaePwoQ1gK+aZXfgrNinZmLvuNDVXuV2pwYhHrHdeZknxERLiR
NQCQUfV56F6Gu2pBoFnbkQmymsBIif9eAZ6s+OJolXL78DNPXBZhy5Q+CElTNvrVXEfzp/KVy3nZ
2Zf+M1Max3wODcAFHYKmJ4RLgDwNtvwB3s/9d3HzwVLm9Etz6ryTSAko+yOquwDGLQL5y0J3XsTj
oGswkmApYpKqAvJlfQHTj0QiZM3i95+Y5T4zVF0WM2/a+X3bqMLf9vRDzBhIS50eXVAOTcn5NVKe
urj/1sx//WQy4BMEvdzrkXmQ7EenBsDJuBp4iWeRiG8azoL4z9Zd4owYOQHrw+B5nQLJYIAP8pSt
CN8INps2oMD+58DBFmVDwOyXgSAZS9GUOOOCwAyIbFsb9422CDh1eEYEuXYqVjL0XSKS9imu14XW
84rCnszJAqpixhzzBjw+LnCmhGVADKEL03bS3U57v8ay+tgB71jC5dbnVob1XATOhAaLEylfmgLb
hyJM7HqHBB1gfNC4uL6jovnJAVDYpW3HrtdN+Q+bP8BK6sAPHl7f8L2lc1Awr2UFkcSNecNTw1IY
HljNNzupRJq0iikL8CwNssNkB//zQAIN2qJcJMTHubHV08vEbv3PfwIcG1hndVREQwVtHZyvq+tA
beWGcmn31/zjkc/pWbz0O6Sc21oTyqyKyVn/PHK3euSHLF8nMZD+PryDZ+QOOj1o06u0X4cl8qo7
eQHMm0QKK1B8+gXRZSDwsQxcQgr4Yr9A/w2o1azhVCvbn2zuLDNfGpC3rpkXI8Caiu086gahQZHW
9pOurnEfQzbssBDFim2QFkXwWdK6XaTjpHv7bGIrKlBQggPoqnyjUVkXGCJh7adbf5qK6rR8i4Y1
oOp6LSjY9T41hPK2m4FqNC+wx3/Cx8ZEVXwokDntGsIzVuIAvVp0Q1KE+Chvt/LyZSaRfrvrplYl
9715P68trKOSkskEEztmhzLTkj0oV9+erna9V/8HLMaVNaLz8CVLjSv/Fu6vCSe3vJP7dpL7vSEi
DjRfElW7r7hIti09ZV1ktoQn2y1ixf//UQQuBHdzmLDw0j1t/2QiSNOynEOdW1M52/cfojzBpNol
wQ4N03tjj0lK0YyhOXBq3LnQnD7WfuYKTj/NBOkdTBrpzlM5b9kDnB3UJVvxetpbQmV0huLp54jY
jSD+/VbHqDbGhOYsaoktqP2kOEiYrDLdvzKVngqmanlotMGWOIEiKoEDmGNLfpICcZQfRgBJRngI
t6aL1+iIu/aFvpPCFZ47b8F9wih5rUVSJaT7fvQkSvWlJpUT1r9pFY3+wxMe5wZcwahLFf+ukZow
IvrRXUEuOLl//K9hmC/oOqQwDmf0tV5WHJB4sgAJj/SGzaPGyYOKYkNmuCE65IeIDc7HNWPkBGQE
N0lzK5APz6TD1U6QmzhDj87E3yAbJtyCXeUFRGVF/whBqrFqBeCrRJwSJS1j7KWniz9R4HCcyDNL
MGtW5oyNwKrfYkQHJJurhBQHhUGsvdLRPdDK179wYoSbph3otTkJQHc9AX3WaWixGLUYPlVoC/fM
YrxjXHcMHykP3AqvFxoOoEYfdS5bSZrfc/MAHjEAWgGERKEp1jWLMZLADfxoO4pankHDio4N5c9p
VQtUMR0ZGbvP/NA9kVllch1MM7V1pTaYNiuzC9qza4WiwUakGsS5giACZscqRrO0Buv+hg/2OwSD
+SWoNi3yhgJ6CJmXRXT+ZB1xeYP+H5Xom3MMovL/MEaReFl/O25Mr/UIV6aJnBDzzTGWYWQpVpRr
V8YksYmF8vzyXdh/rei2EaD+Fdgs/MvjOrOhVq21S+2Zxz+z6kMXBlxqL6NuyB6viMUjC2BkbtZI
lRzbqe6jm3FZK7AreW4Yop0Phd8sq91jlL8sOX+l71/v6/v6ZDMMuvsIZYHz4AzoW5f4wp8d+qMV
Uun/YA5oscmodS3g+nVlRAjzglbdUnE1iNQmS6qZk1f0rou+5aBjVnBjfkaPHjy28trBGxQW/yez
7wiNDBuP4hKnb2LPWvUF9YozbAcjNJd1+QXn4+wN9HWZluvmm5ImAXfXzcpfniKWNxLbHL+EDKjP
yM8KCz7o3Q/JNcgrU4f4LxPs3ckwjyKOBg0MZ7YUbvcq5j6Dr5rGYgyrNE9s5CgdZQOfpR0W+qmZ
RRA4umQv0cqCs/+Rt46lsf+ee6thnmxM3vxmfwHW1ALvsqOGt4rCZXxunikCMcrWEH9cbj8qWQ3H
oGPE2zkdBFnqRjzslYEDSyhf7jspl/3QivK/MP3Jjy3d5mZGo+jbXv70hsdibkThjQuXOuMTZNW2
mTWWRklv8oBGLMp/U0PpPVbDhTWJYhuE8PSJqYc/XNQ2sfbbhmlouQcNrmjKDFoXlzVSLaCEooVt
cIe5l8Wp5bxsksAMz85zkQ87gE4JmfYNRlBv0JJXrYKeUi0hh1itkexIfb07BO4yslCY8Uqt/cCo
ZCxfetLGhQsIOscbgm7YrB0yQfphnVwRnACcLubthz602Gk75Lj6n+XiKCUjOoBm2yHeP78EM8yE
rYGWowuZ6C7JZPHopajozwoH2D1eXPOsP4S+O1xVCSgALpp00cLJdq0JXxDyL0KUZzvk1xXXZWrW
exkTbhrEFTLGib+cTzwvo0rXFLpIw7xyr7LRlFFBo/qBGMIdeIZj8aviqTqADiof3kPYyAJoShMK
TY8/hevhF3KDYMihdnACpzHjTyNX7ORbUqWK2e4A/JrgCG3Gikt1wHhOCDrcOA+GsrW2qR2OZNfI
bGPh6gITg7qkrT20u0LSZezSbiz18pZucaBso6gBwTtDQIIH5d/SnyrLNyiGgPqepmyybJ50yFPK
x0Re0Tcq+ZYLKW4zAK4PppPWjDzOLfVaHrA7sDAM1VaJb94KPYXcblUSdv7ht38iQPasAHQkZehI
S0OBAB68bvzyJ2KVWrJOEHio03Vi6fsiT8iwxEhWS5LQwDMqB5czSlS+Tv1N/uoNiFB1ZYRLWnvS
g7ukSu7rpGmqvaFrTQPUH2ConnWa51pL9e1QkRSV96gu7aRKN8OTz2gm0UJurZidKecYA86qHeFu
7HnncBXCvzrKkMm7TVH3uqConr6WpSrdAsrefbYmMOA7V13Psx9eF6du09DjiM1yhxQRpDglIwKj
XLoevfdSiRYDW/+0DN8ZzYbQDStJ5gvTtMz/fb0UOkCRx8Pv34G4yEqFNH5AkQY/hdoKPshUyYUQ
xuu+LY88nI25sldsPP6w7S4GKnDPXKTJTBKfe2DbLcmGCZ5udOhGfN+coWM9p12F5BfRL7/MvX7q
5Rndhe74/tYGy5gNkqir76T7UtN33RjXpLF4QqVMXv2YLxQyOuLhB3IS5y6IXHCUVpcov/0zYljd
qAe+jrPnsImTfcI2tcP1kPzxoV9d7Cc+Lu6U8UXd9hmCCBHh0n65+RJCnX59HTpVTF/ORfAe9/gH
KtnXL+x+VA9vxzxfexalQV9IqcZEBfEFkvXRhwBeX1nTO6htUsd20Y/6m6h+JQKFa+g5wa41H6Bp
jXJw7MagskxIQQfvhHhqXDlTwzuUUd7OblGzscMejudZUtazEYz06oLlHU9FN2DN2RCG/xVF67z/
x6TFNrta7dLaPIAxjmIECddtDlI8/ay23AnONww96UxKJpRq4Ur81h9TaHLhk9kjyTajD8dRyLKs
0aFvcMd3O8/1QbyntMxXj6QKx5jupDoh3qwR745PJd0Iplp0kjRHVANEnf/2j8jzy+U1jeDjC6ok
aOXXdRsRHhxB1rd/dh5zi1jCs90smnsl5azWIwej8DjW2s1crHXeV5/2VXx5RLK4s72rDvLDNhhh
JEggEao2nOI981ovCBYKSnHgEyIuCbC00+QbjR70cML+C0VD8c0/CiBUhqcfXnFp5wZucxB2WaOW
n8QkK1c9sf8p+F63PpklG5sqn0y0PxyuRllQf7ZqTzBruW2Qwb6O6ubwvYOkxYcQmQ2dsUBXuua6
vzFPuhYxR3+mjc1uOP/NeVnSU7ehoxCwVbsnP1gcorcadQqRqpAaGXPZYtSq9k5G9felGxuzYADN
iLqESlwnt8YsCiMcBfBULHG7RLWh7g/zZMVTuIbMF9DkFwiLlg/NMS2ciJe61fce56JnVN06Lf+5
OPO4HRWPNvxp2cugkVtJzgzHCrCjY0p0uf/aeNiqrfsce0RQVTDopB8+fY0bsbDCC5+xb2L7rEZO
WS/mheBhj1/lwIxUTBQXviKP5/S09Z3vJKFNB0QxVAfZ4wolGxznqcT1vocBKu0HnbNQT5ukB3Ds
Vy/2TDl2/fVQZ6Q0HvVIEaHPPwvQBW/Dn73RM/OD2Kq7OEGn0D6nH9lx27pzwP0xtkCtTrKquSXA
LOlTp6F3FmiKmYZs28189UZuMy7lHytawRrckvnyb6p+QDgQFrNTli1Xh4H8nlB8edLhMQcQ2dxc
RBpKQfxcIKHs+pPLOzFiKVFyauI+TwKLnRUS3F0jG1CYWadmfVEgojOzjvKmesnjs7P35AgyIVoC
Ws3hjt/MOdYUh4LR2Axk6+2jARvMrNCKMvzhaAsdgP/hZE8TMW9v6pb56TkV+oukh4T86OVR0UOX
pmzG+vt1jU+hOAH/noYNixSjAbQwv/r1jY/ihE+HkFIe75uF1UsNwoes3WTzkOO3qd4K9679sa9I
p2seXdsxkgPhShiT6sCThXMwqaQeC8u0cUV5Nis8G5aZx9L5qnUtBmzJemMx7/WBOmIG/Tyx1Qqe
nO7LoGQXA70romA1lD5gCbGWvwNB4nxi3jSvmlx5rp1kYdCJCHkIxzqF2e1z8FYxl2rcEsyuLy4E
6PiFEe/fK2lQ18tQ+azIVi7VjA3ACpp5naToNXmzkAHWgFZ/fwFaYCeBVR+fLXGXU46lpv6ASGpy
bVS6KvykC1J55mwEgETvbZnTJ3MH+Lyu3HQttc2sVgCsxAnKdyCNWiTuF1srCgVQwhQAMwAAjKg9
ThaMbT2jWieYf7JN6/JeZDal9s6AixWVPkPzadQ6TRJFSiESpPf8eKYZb0nYt7Nxl7/wcui7/FNF
depeSYXkmrRiCqi42vwpxKKSSXQc4GnVKkJ6wS44lio6sC1Ros9+TspPbIYCNn7MKzbfnDIvfc1p
M0xRrt6CV1GRffLztOKCBNKqYrycLNqq+FlToxNdnuzKMUrs4j78CXJTdj4CXPy6yCSjL10C9aFr
nKcqGcuJ5lZFpZNXsFdBmUmUyZxOctgxaISk1BuBoH171Y6q3URa/hFkZ/JMmWuCPpgVTrX0lzkd
9c/iMd0E68+BDO3GgWEJPYxism1mVO/DnsFBw4o/LaSWI1D4oFOnBeZg0EPyE8hw7Vqx5iIFVWsC
EWa6SQ+LWLINdorf3I89aDH1rYp0NXIQSUqO1lX+s8EwkB8I3coE9Qw7FwPJwenPXXr94MrQpo1T
kFB/4uI9vgc/6A7zgk2aeF118kPF2k81Om1hzUsMyA3h6DDmuCHPLw/9PxzWdGxpm4UiThnOgTb5
IUYKLR+5zW9YNZfnNScU8sfb7IuLtjkvHKUu+IwbWVYnMIf38GhgVbLrPx6/4kdKzyRgYRhD0fsN
fYEvp/Bzga3tL06uwJsrpJMwFItbP0RtVg9cvnPRfxxE5ZXrFMqC6V9OTNXlcyX5G07wObvWmkg7
t+8naHpOdZa7mCTCgIhdI0hG2bElz7KdYz+59du6EhxMHWu42cpYB3lxM6Jt6MhZUM81wMZiaQfG
pGl0Qk59mDOxPtmRI9RudhHi+q0M0oJrLssy9z1uYCEgFTlnsoqJt2k/sDsMdogMjRFaXTDVSmB3
PFVObEUdRzuYL5za1O6x55zZqNnz3uGenF0y/TkoY/wosQo+B6qbnSupf0xCj+F+JJo9uV3S43so
e/O/YgipKyxbOSOqizA3D81NMS/EQAyy9Hj1seXz88I9PEYbozJyNAP+5wQXzjBm6mskogstVRQ/
36JqKTfO7Lb4X9xVcYkhRZMoO+y7lN/znhzoiPnRg14Yh+iKRFsnGAI/gj3VmBP7n81xKl/QMK69
zpT9yKV+oCP9/vWyzd9fB4UmhzJoqNIsXXQ1gwzLTs6q0YTNmVY4x1x7qURUJ/VQ1jJTPaqeL5ec
LZ54w7Wa+tRa20CPn8kOIfPfEcz1hWZD9YM6oKJr285ivFNsiknhFRa3YJKUZAmOZg4EayZpoVA9
+SLWY+zb/GNgeX2GquRx8yyonJvF0JihqMTfxfVvAQ4UJ32suZnZf9FrOmZU9TGAmSVJLFKhB5Tj
y3t/pMpH8v//9y+xc1pgR1EvS7Tmaxku0HK6wdBJzKabDNIKh17/eb6h15qnYTi1yMUHqhRuQ5gd
NZ0bW266Eu9St5lltTQIYhKUJuhMjd+iHfrJ3YMrNnSiuTqYqop/0v5o2gzcPKXzDTaf3O3m6MoE
0IxF+qsz9bXDuzD+1XrupFez7v8VarEo7WU3YrgMikG7FyOYQIAIVYO68+smsFpgDqPgTT4Q9XQn
ziEJnhUqbO71ZUufxgFZ3wyRqMM9XOgDC2OPyOH54aXlI2RAQQKdVa91nKgqvu6cSF5XR//Wf7j/
6NCtIqBvPzxxs9fEjhyDjeWpP+HEdEPqSWaOa8hSjhVg5XNEPNhS997N9ujIkL0MCiKisHYW80is
eYuCrlmCMmWZbZuVP0NZfr90ksdZE8unEz+cg6GZl7DZ7zxeTEehqWTKHancv8WlB+HvkAniXTwO
bfPIscrlIqijNaE6fmIO3inamEG6UOniCqjs2ISngkFsEQt6uBt4uungImDw5zd6WfzJNEqPKT9U
NKz0MnC23/34TmSCxa6B8fS12C4cbN/JQM6Sb8DioeVVx0CmUG+FJchhDADWxH2psSNiopWhgXMf
2WO5Aan/PRKPgrH6FOj3MbCeEF3UfraMl2LN7nX7tdDCppo+6G8Vaa0pl/NnPRT4iB/SETYn/GjL
baTo7gvtItteQpYIKuaXdf9mwoj78kBweA73NzTcozpSlOutcXc3i9R7FrUUy/vxXnmlAJpEydyk
s9GhqioJT9U5uiMOXBYuwo6AbvErwD/V5dowZ1TCGwM8mdHOJX1W+CQgVpwEBnbqeyP5GudO/Xtx
AYmHqRh1+I1wwmyffWLQd/SBxzT4ET1My19XO3CmJylx6tSmW3biL38a5wgQHOT6uM8Raj5g8vJf
MdAupRS9htu7pUd9KAb5BdD5DqhOy+e7tQmaf39AgyFgNoGoym4B+ugvll3orjx06VAYZIb1CatS
qT55Fv9VbF7axBJc5Zzts3ZLD+/vpj891n6EgxjcM2b+R+xMCOET72myzE9t8jyNW4h7Tn6e8oxz
PrAQxqZ5QrJB5ZCzS2gofD39VUv8z/AbayxIvVyx+QiW4y39Gt0k3eQyYk7/HBdaOg/6a18t1gjZ
2DqygZs2JiJ4+fgknXJlGg5oX1EJgbF/EXw9CU8UhemYOhjmnbspqM4EwsWqYlrSueMXyfW+Mmch
JTh8URMsAzrfec6gR523lQZE6wDjkDnO23LOUqk70Nfpa94depBnr3tDWHrHOaCEF43Zhv6VrbDY
7xKKfxpSySaUC26gLh7oqAAt+k/zWYlNC9YWOJ1zZ9lXlr4NIl1FtdLZCK9Qr0iHqwF/eeD6GWmf
sKL72HFU2vJfq4VXN5GeWkkl5aet+uglzvvwNN1RpAe0o2+KRgSohJrm5emkmdZij8iMvRs5G0xy
4srjHsynNSsLLlKJrLgOaNaLUFzIrJWiM46CwM8pSTYZvlgGuMb6O38D0Ep3gdUskAfOHp531LyR
WOduMxqn1GgyIo1mzLtELJjtKSx8sJ3qVAJ7pBAS6fxXkQx5I7bNcDAE18vT/YYyR2VIztdDWdQv
CixCUy5BZ+nSEd8b+kG1A/5aElnyZJIQGp2pPBj/XPPfWi1P5shv2e4d0jFRTcV8smkEzrRaLJiI
BpQQ4qmKv0pfY+evSufLxxjfQBFlBfxTiTFsZh36QiH2F2S6qpmTbVC3T3guGhi6OU3bULS8EmE4
NUSC3NCKX7GCk9ArrZr2S0rjIAFidatoYdELvJORwczTg9W2BkcHld3l7WU2UefgP6cnzzI7S5jJ
xcw0MtdKE3llF+V6TZA7pIPcNlfpv9izwjyXj+sobt1LLS2R9HjVDdsAyqLGn7SkZ1eOhLH3aZwG
F/g+RsznI2XWd0xgnPlKhYbqZr4GdN6N3mnlMYuQ/aaRJV1vwO6BxXo9oO1faZFkoElxye2kszA9
pXh9l2LZV+8fR+alAPxTj4hM4NcAkXxRLcaWlEVquxZNTDMgnXNZhrgwxFafUDdDTeJQe0O56DrY
Kra751z2+QduQLbwHAV42WEm9eUsQGDWeVZ8YLK5KqCaxS7J18WgRqNVpB271+ogXYoqNLIfLUcD
JRHEAdxEfXCufkdxnAEbguk6SWay1gQMma9WOjyvfd/CRFwEzesNhuI0v0k/KJJeMmciMHhBUTF2
9nGEldrLvaLcE62zae75scQ9eHuwwJpU711q2T5KGxVcB0f5TlvnxP8+F9KJgmip8xHSjrzsQ6B0
bbxtNIDWFvied+Diyo7pUUQO14hBjr/hZhx4dc2TU/Juwb3WyQYt9XOTnnoWmZ+pL7vK85po8+VW
gmAfbhIf46wLoaEJdOyXnM25fNEgXOPQcceSYynuHilehL7/yKXS+RiHETP2vhQ7CX57XS0hK/iG
7yrxM3ZQfzZXMcr0vrZnRgvinVXGdPJodlVymqNkiySJqL+ZKpu7QuJTwAaOgi2+41U/LPy6XPSO
c3uxRaxH0dRvgy7oGPQTFeiMTpr8N95iAx5h4/tTOix5vXW9+xR+qzLCrmnsKBkmmNpnZ2hbOuaK
fiBmx9Xlmv0inreQUuHrwyxr0mzUN+W4cqc5I8rXfyiUsjC9n6qUXJXDJ29gzDgkeiQApXDzAJEm
9/Qzds6wz+WLgA57kgJ4Abdb5/FUlD6cwh4ho/Lo0FWG5GySPVoheVc7wCKwubuayKNms/9aE1uK
KXnREfLNu/vfhR79RFkdrfRU9jJCRWYV4K/YP3FnCl/pPsSoB6qhUskS/9roIgTYRpxF5or4+wEM
VyaRdNVVC4s6qKpz3TxytFB9Q9cXWn2y0OkFioUHFkhiwUD3XiO+knWQb0F3r+9X0mLZIZ+ddf4+
3D8eIG648mzT1Vf+xZTuT956ZoLnIDHaMN7bLYx5dWO6Hr+XCHcG+XBp69Q3ep8KDrZhhyibWn2D
cnIqCjErMBkwjREZwFqQiTVg0K5odst9VwkxMFrs0InRQ3ad01zY8SZ2cqxlCR5Ddb39zDwHBFLO
7S0VzTq99S+tlDAc3qbktbPwkig2dCQm77ucEZgF4FdIERIJv9ag4auEDwFnocZr0fJnWGNe58+w
g45hAchDFmdvimEvcL3WuQx4nMJVcZejz58qXKzvH4IupYWy7eXqtMLqgOK7VYa7lfOW8+sU+554
RZdcLmuiWvxljKwXnPK+x3X27CK4d1UHe6iwk3hin6iTgzfi/NUbVCf8NXmEnBNLlBGqFCLQ+nEw
QKOXS0SgOlbkKCWVsGuJLtEB/t37I9kIGXavjGrV6XVjVKB/Wq0coNiv4waXHnOGxiFo4CxUzMah
2zcZCMHSyIfFRSTzlirCVCQL8CyN/T6bjBhQhpvboVv3OcuaUAjjvnopuaOwADUD64a8rFLSfZrC
A5smNa+YK8JY3KQRD4hHgV63wOiiUZeV0AwGKHMtOJ3vQX0wEMeBBSF2LCxp+Ofs1gN1JY6kkPun
v5GNUsdA/s3xYS8VqBPFIBfHiev717PJ5o3NqFw3pl6J/uKT8PIxDBUkvfFGiQgSAvMSOwZFnIzM
Rk8FYolDVayKBZn2UoEZZpUGDtRSQMr/ruzeyWOUdSWGxULMRy5V9qOmPz4sdkrvrYLTluDf1y8I
pMFONejcFC6gd23D3WvGfl+W+lwdZcZ2JvIfWpvPZWsxt3dkNK8DoFLWwGQsCDEtjzrQDLxvgr4z
4C0gA3jDTgKTNQxcNeJ97uEuCbsl9GHXpn5dgzeFx6x238QtNfTxnEUHtOINOjRnIQpcwFMSkrtb
MSrtODB+g+Eg0cUVL/pxrgHQnuvcrUmweF4MbhOnbdfTP1p7JOyhMK+hmAHBqVWILGyDu9dbHPxT
l5mg7Rrbg8RU/gZK6f3hpZPGEgh1yuM+tKnXIAbQFciqZM43Eoj9Hr8wPj1EoQ+kjm3hRqc1sZBm
OIIKNO8RMncOJy9InhO0NbvdRv+03OODeRBxgTLNUhaJQRL4gTsmWYJe082mFwsyqka/d8uxwLL9
5eGZfQgqeGqqWmJ+xTSt2hNU3dojDpIf7uVzxnMXbOda1/HfQxTTSQbhRQzYlv057jeHvaqnwl2Q
uIOcNrTfT6574ibNDG4H7AJf5af5qmJ7EMBkFfwvB1MR/JZiIlJ8/zlxT46hAgGYk69+eM3CHuzA
ZooibYqR5wnHCgSRukafTDv9i5MY/eIbohljl7dSClHNDEqVh8JXslHLzOGr14/gNbSMD7i+TMaD
e/+1weGEWFM81R+nKdCOQJlFqfVoYpb+2ECKLF8jgz5Pu+V5ftvegGQVYt3f34Fwt2yXAGJ/7+/V
eqzy4n3n31jFTcrKlRqLRkcbk+LZEMwQPceG2GeFJkt23pfDhsm+8qDmzjsEoONG3wNnM01/pRPt
8P4Qj2IB2x64ijE8QKOHNV7agAuzJGLwmTYPUFk/2+DKlabLiWSRv9gufwbfjITHkshG9YzmZUTS
dnQZ3qr+WNECKqXso7vKzg83DMMWzUdkDdggBUVZEwd1TVSZwtlOwce2m2XiSTFMZ4V296y49x6Q
1QjJxI70QGIkE3mDsI+bbQtBvcM6cFOk830GJL8jrhqJrSoXoSAVuNcqAhpOI0AKv/ZpacPlNWEl
ePhlwgUhGskuQ792kZyVbkM/JMvBvOVNKfKhqy2CgHNFEib+0R7d0+nyqC28ynJWjGKUmzPE5zM3
NSwbM2ULbDID3GGAEJrrac2ul0rZX1LpEH0Kpx/8jqrOwrinPwC1pCf+Z6K3VFk7gChFN+/HcenI
8WN6gN+ohTvqBsJrpZpd2NjxMWmIHgNj88qKNxHl1OJ7EKh3WkQ+7B79J6B7R8ZjKrMQhpcSu2C1
d0K+izUmPScHclnQSZtqFSsUT+F5Rtv90Av74XkhJpA2xYZ2Y1DLSEmjAlXU2h79+auUEz4iBDXa
t2B/HZ/ukdzJp0qkQwE3Y6hxndwy5LfnP/Bx86ReVewwpNkCOPfbIVNZLqMUVEG7M8XE1XmpnkYz
X8h6UO0i/E8h50CQYk+2J40XmAfyGrlvfZGZAuJXIRXKzXmL7+f8miWDKUuht0rxjIs38C1dMYX3
WWFqpUFYSzP7YFWUiqBZ1cKUacd+es5KKvehaGL9SH35W/pw4jxV6rqcvxViS/5sFxYpUgHVagqI
eYJk3NwcAV8BsJ3+yVBZ2PlvckgdRK4CqcXSDIV8dqjkMuEP8DY0UgHUanQeAkG7jMLML50tNeVl
aFyn+1RjAQyFtYY5UYb1HPVfQ/TrQRV209WeA2NMIFb3uGW0YHhZ0NYt1a/0I83xqLEzUGjh5wAN
WJdF2TtALPcTtP67EHNckpfA1SkY+q3HUQNuQYVcl6t1qujSmjSQv86SlXqTEEsdFB9iM8w/B3KI
zNpqnXn7bKt74/Mf/0N74Z7sfsmtSEouhTQyPQIElL133PHzPnCVcc05sYOpd8Cqqu/8S/ncpLVQ
AfEOKQdK1juwGls5V73XU5LbkSOPuvFO1WSZjktspZjZDiES06tHCCMWidZNePwLnORTQHLt6xvs
w7nUFVItu+MGFnsdNpQQjlMM7RadwMpBUWMDgGw8SblS8XL2l4nvnZZ0+486bjHMsv48FlMQymDx
9Ca1CLLjpNr3Vkj+/cNHb+xJz0TWl9ypQrcWfEXGR1kYXAQYroggr00GErkLSz23oo3uIaU9I73D
zWigvPOXWmxEkBCKKI0QhpXhdHSV0V1NnzEsvujvVcgty4oIztfj4H/VY05Jn4cSGdQz5kvi/Ud3
m2syhMRE3FwX2e9wjjKMBbBPSZmA6QCaAjSyiy9xtaU1dWCo6yzZ4fGIpg28coaV2EZv1R4MklTS
Y9cEeGCz6FPsPoFokzc9G7cgBgKM2qZZD8kLmqpWgfMpwN6rEGHaxPBYiXjLU97pu3hRsQthihqB
6DcwTsP/SQLy49/Ay/CUW/J96OG7hg7bB+nAOmI42gN1hvpjetzI9p/O9reD+qaV2xFLqs/+bbZe
H6TuYjzE0e7d6gJrQhKiZauDDeJvW2eIYXPnFnqjJeR1eVmaGlE8llxU4To0nobXN1z/qSQlHZPR
JgHK5GtKdLLUF5dsBVlk2hH573VZ7FKXqVrxTCfvtSt6J3WPNlLFMUgyvUPst2CMZsjL0LHc54ti
ZBHM+NHnXOEWENpuf71doCPZ0Zzt7tWnoITGFjI+yV9VVyVdj/0s8yRvdTJmvPWfCwZsRK3/8NxD
o4XoEd4RqpCH0WCTmYlSJM1iYB8ox0NiNcuGAwMw06ZxK9KRuO18WVAevvVAABcN44hpLwuTeVW0
QBczVxm+kCnVW3OUwfOZ3NjbaU2ofBPCENib/qk2onNphTAkADgaTRSLoev4wFcPxfvczvVCRpW0
iU6CNpUDzYBYm8pNey2korvgR1TB3hONMXlGYYm2SAAlmkv4qhY2nn3vUGS8Vv2iUj+Q9DSHhm6G
c1nsyIG39tGmSddaEToRjCUjIAkjtIuq+uUmQlhJaunyr0z07wmUGIMna/aEzr3Qzfs4+d/Y9yvE
c5tkYC0FHQhl9QX/3gdCNie79xYKHyXumaNPIpQ4e5C8pnRFnruXayYTw4RtNH2EXSdqdu2XhXkp
Z5DPtqSe108jXaKdtrQBHJ6vhHDJUxGIzBTBpPYyyoCAnHuSuy4MzHl1KU25lbMxsQlsHqVzzOQx
BIei2ksOenJTzXSKekdSV9XrhMHGGAUDDWbmfY025A/Uw8wtJu2t86l5/9r0ZPY/LIL9XXiZgDF0
lW0vS1ogaGqI/nC9nX3nv6GnkiH68M66JhXAcVlP7TauoCuQ40O2vahAf/UhAKS8J0ODxgIFGzR3
DKGJK+XtpWboG3mshkcz81Ogk2/yURk6C30JPbqR6iwV1EPX+UiTKSns92iI/Hc8r5NGsTnCDseq
oKO/IkFBFGZXdmjzUN2iMCCaKytzwE7M+AFU8gK2Iero8xzDUe2p+iVqvDV5ZyNFlj9DMHHlDgBc
xrJWkidNMtAhm3NPxohS76l/oC8W59dSHv9GxodIf6XUKhJi/96y9PRrUYLe0Yk1BWcZ8HQ8gscx
1VTqV8gYDensa5siTrUy1XV0T/4w5eg3sz8o+gODZ6dcufhmmF4ddjRMff/xL5Uz6MuYVb0jdD8D
4fzaBnEulAlWFBKHc2TIeUFq6Sy/hdKscdp2ud6GlAvVBGNUHY4E/cwXte4GtVgI343H5kZ7vro6
H72veRDy1+0w+xZ2XcDAm4IzEoY2wyl1G1axDtQwBRRAlkrvZRHgnJQZWWb87qdJ/i0wGhuvxNuz
uD62+TEHP6Pb3sryHsHfhCaIt05bOzJh80HTojM9z5PrOQA20ix8zEDEjalIXti1cTrOYh7zevx8
FI0hFOJcWKR2yOFfAw6GAt3VChD5n8d1UhebQBZ+ViklHhfIlgCGekCxB5bZghx8TrUUJcY3ooTV
f4C+f4yuZtf/NinPMv/svJ+KPtFRfRgF39Jcj2dTFD5XtWRxDUmnN0E/Xi3feFmloicKlq3IudZe
G2JUj6FX12rM27I+044K2cMzisL3Ak+J2GfBtUHl5VwGV0HxA5x80FAN+mk71FAm9LmWIiTnPc8h
Nh5VO0DkQX/kI8wOzeVS9vpUrW7Q81kOH/ukskRFK7sWmj4e+s8fqsGhzwZWwR6Djh3cGF/s82bI
yvqKO/Z/5TrDtD3PjfKFmlI7eYQvwOXa413CEVK9ejTAfKuGpnQ70ir/g3Ve5wR3gG8rmwHXDvPk
1B82gjOeQwYbD3BQSdBJDhCRSNpsJrRkgdcCSYyydk8wTpqO9n7SElSOfpnPVnEW86N1lvHMFb1N
p0/BWZKx6/9VPQoGyPzA35cImB7rvqaXcQl65EHmOzptA4+/7XexVYcMpnE0zgbnj/so5XqI2TUc
WCktBB2oL71tlNlUvucc7z3J1tbafZgGGCydP9H/BYVqUGYEmP75hVpASYnDbkqYXffcjg5hWlrv
pbasa9AebC2p4WZYq9PCMHdWaNXyRwgHIgoCq5U0C8m35P7MyiYyFjr84IZIWiQxwBzN/t18uLN5
uqK1gZ0bQ2Vpvns8gIGEma0JEt92ovmawIUqjOUgLNknylQYdxBPGUlnnEHQruhyfAIkY2KrhK+N
gqDmSj1X27PR4CMW432sYSDTit0HA3rDQDzs/gyzDvHgUx/7mv2/KFAv49UwsezYdt5RSmJZ47BK
Vlt6WVYLlMr7aSAAqBECusQft9jpVYtv6gqnxFM33nBtD0VTQ6GMFOR+yMhj4OwzyFWoRWlGzgXJ
vZ7AWXyw+hEzYycpSjxFGpLn/WpqMnvuvTirszplSY/2XJMBpY59NDs4XWlgZF1gi/T6WxEBt8eR
woFsZ9veUzWu6E3DIFKnYOcTnPJQQ+gSln9Guum8/YeoJZ5CXkw71F3TrP8WQRnmyxiLn+Ot5G2G
oDstsP+f6zOHd3umfO3ybxRz9vHQVDXJlhpCTSivbTGWuGgfGKI84jzsDTJgimzkxy/R6Zr5bwcT
Sd8cqu9CA0/vVxg0UEQqNjHDWa1xTwOwVhhrh5PyaLfhCvScR//d+vVtftvex+5RQnAApN09ktsr
HeaZ/zcGbGjViBDmhWEhPtkiH1S7vincRjYj9vOD+ER6lE/KHAnFDCblf9pR4vhZ33RAu0I99ZvO
IckQ0F3Ciyod9ZusAWA78J2SA8afJFfpWxkRHiqhmAoA3qFmUb120QAPXNbrWboDqvyDdqCuH7UX
QDbyOdV03giSRuWzH3KN9h6+VgT3htQGIy3W8QttPkqyFYwHcrFrg7vgohVOHupr3NY6o13Fzy4U
6lwnW02uKKPtStS9ldt0XkS7wZ5Ia/pC1koUNKzYXbsOnMv7gzzUtvXnzXn4jvYwawy1SCK7IJKu
i1PT88iP6vEXsehHf0j/SPCkmJWoVbngZGxii61XxP8A9ccDaFueOdmfPEUAUY/5WzBRR8xJlSiE
cvY5WAFFuPsD+kx1UpfPJESCrGJDH00aZYx43RGENP8hS+B7mir1dySiu1SBiaiCB848h9uvD2xp
GYX+P79agmWXEpnuQi58bbAVScKqhBN5FKWuP/Q6ofFuD4E1DVMg23izvB5knf4qGmXw+iUtH3V7
83yUwY+TeGSocYMW1qqO3cx5SGCftEUf6wcc7Mhyh2wJXcg4VYSDHMP9ppPQ6YjXdVBND+vQWGNF
pTBq7bygDhO/tbtFeN7ZSOnK0Q55xqatomOtq0ozqP8Z2B0pYA6KApPkCgGrw7uhYi4G9k2eCMh+
oXjgJO8JPpuF/zFh0RIVOroQCCyhtS2eobdqSfmuV88j92CmZ7dOvset3fIK/oPUrXa+p8vm7hgk
TuGjXFoCfHWJYvEE9cCF450s5oW7uema4kVRvohpOiYwtcEtAj/urN11wDwJTdF7/SRCssg5I4yh
SMgnoqFv0PiWaISlmD5TAPuj5DJHH0c7nL62kdiA9RWjPylG0AMxXUZwnXVWrphsi+fMTPp/cbQK
zCMUZvyrOVBd8kiH3PXLwDL0VoC7eEZI6EMJDMHUVD3zDzKH/4s5xxHMb0z0a0FbvFz3oq06CES0
1bfEiUOKy8LQxrQSEoKsKjgzzfqQI2P/EbvO81V5VhJnZeEyHtR+ymY5o6LK1YyHXkylhCfUR3+V
kzsxJUY6xzMfjfkhx61yi4fOMmZPpdw2Bpb5ismJs4QeeRMvkzog3Bc5Gd7ElsxSSstWoDfDMhRy
jYABFUY/oQsxWEZmzW42DTBA2KjnwD5CJs5WjksV4fPj6O/GIQNAS7Z0yrQi7zJais2J+0hX0bRy
iwy5GPOLoVPBF8Vm5sW4J/JADzavlUwro/wailh3H9a6eOLWWP5WuEhCyoJKG9bHGtZTA9k6MS/G
tkZqAGWm0DkhbCoKhEwOo7pOM0NZmMQkW3Po+l+rDDAYUl3hQc/UwjzMQmw3BEg9AXBKNSdy0fOa
ZZMzzk7jZdKWS+a1rykmC/CMUb6/uB2QSRg0BhY6B1PFXLFnUnv8CQbI8Jjq3jJL5oTWUDfnF98T
HL4KskO1veAY2JRfIzjQPUGEyxaNUGPWoffQBg7JnAzfUHipnbqra7oKm9chyiVM6V8dP76myj/F
4Fri7+/JsOEnfkVyrNF6hNzQK1aIfEta6gjvmAC4eXX1nPXDHunOU/oRyr6a5VxuuyCHYi8jO8hC
mLpc8YRi1I4fJbegRjgfz7bTT2wTQ0wwKjgSbe5T9aBzAYQWMtz8ddDQvAg8Otv2SiRDJzq3TBX3
00ZzhXfyUTjpDouAD5qiHGgeqmXH6hcIupvHpIM42D/JAnbz13PrugcmK9QAeO1HBDp0VEDhN8mG
oyOSk8ctJ/cAonS9QU13mI/CBtZM09fpOg53lGoafDeYL8J/usRMBiXfphpmPDGm8XTZfNOi4obZ
kq0UD9mOiiobeBZoyEMXXKu/ljxCNPQhRGo5C+niYjiLVx5/Bx/HQplGGoeryV2Oi+4ETyl0XWP6
qZPVAxE27dJACxWhZ2tqVyvIijgV0174747nBgtnlRPc62HU+BwAebwwVhztKZZfWM4W6ieoBD05
MViBJzZRHV8qT9j5lCzjweslwiWH56xPKlDvBnX4mhD2WoV72R50RSc3kK+LY9/yjCfHEHxL3WTU
S6IR9Vd2JBo9Seb5EvIt7J5pFVv2D9tfCaw34l8bbTFsB1J7s5AZBCteOhKTmj3X8cL6W0SHY08Y
8R1OS1pYd7ucM/ZiugWchBejBkmE/ZHS8JdXbwN9oQbCyZDO+QDwpCaYFykv2LBBR7YacOBFNHbn
s9SMiank9yc7MrxbD7+lXiDCiQ3s54UZ4D/iNgmdMTwDWBvZvlO4/uKyW2pMq8Yjc8pWTD6e8T+G
ya57sN31vqP3MBMa4MWs5sN7tiyAmOaRpr/P81hfq+muQM36wPjf2Dk+OHVWcgx/whQfKJAItMs3
VMVzweql38Q3Jy6EKX0yKPbZ9SQeUx9GHFw05cFWLKdb3qkqxNKrQPshJCPF/68guk4sA2JUnyjw
YOIZvx7yoGZkWhSwmgmGc71JnoT/fmJnNS9YaxYdQ9o6ttNs/fpVQogLrvyRxCq783QG8UayHHil
Fasx9ykw+5mh+9ta4XNvLvnQSH4AYjEFprC6H2vQI+egWQiAnulhh7RNJKnbnNrp4oeiEVIbRBEU
SMscdY/cdxuVI4vvLaYCTMODz7+6hWAItGAlPOj17Va0v6Xpt56fqxCfpQhko+Aqa+lpCdsckyTP
OMaKvD9DxOw4osHnl7lM05Ljux3df3sDWbHICTkHit58VbLqG5flUH9fa2HOGJtZNSEu9g2Lzf0Q
97W2ZeWKXJ9p1ahbhn5ifaQ2jvVQ6Z6PY8NFdrkjLMAsJFH7n80nHKQuPgZFGMm9mFEhlHVKxZBN
ydn4WufaEBtwd1qzEDu1W5gWL5uM4jxXketn31lHOaSq2Yggr/E1avNo49WkxHq6+HH9E0n6dtGk
9sKjw4HVcZqOpaouhWtniGts6BPVvv0rLr2dcwJIPJh7/5q5n/xqvC/01YJEbVkdJ3iOTukia60S
o+jtqVsMdool3plTH5EAyeN4jWcHH6ap5VL8dP0WblqPHcyEGRZWLYGfQqpnd2vUQdDkbDQqmJUt
+KQRxQ0A+zPEutDHad9yFEc+DkqWEKLk7XR4qos3/1/Ez2zYlZkz8sKI9O9ScfySpoPJYncMN0za
dzp/x3DAnYB+8Y/sJ680IqWIZ+9Lr1tz/RHWqS75EReTErhkS5EEu4T97uSrv5BguS06K4+ciWGL
AHQiHIhxveWgUaRdY3oDqle5rYEnd0fBcBwhriA0bbcw0KxxnwywozF4uRBGnIF8dREyzXr96WDP
Qh9Cl1LnenhJviN9KaLp71Winlr3Afm4aCDUzgSbU0WRVArT0ONjzmTE9Mj5KRtiAs5gv43mIgzk
7E5jmVdtyG7mrWz+oxyMvYJphndSkOYJw3r0xwslGfuYLiA02Dnp5bMIinBgT9DsV4llwF0UkZFq
HGVliHG+qKf7yACxxXIl4k+LtBMUYdIlREQcOWH1g7nGiqu0De81z0oT80zhKPlEDur/7vSSn1VD
nKFCtYkoRNlUFTNdi/fQ9TZQypbvaZMgJ4bfVEZPpWLB9EvhcR7CmC4J5EjG54bbkQ8fphqeuqxY
LMJ/+L83mwqMMnjF/LYI0iOlVvrL7aeGDH1zfv+Mt7B3VAyHyDMYm7IbhWL0SBzWJpRNO2Gy2+Am
zzz2lLxyMd2hNfFpiQjPnxEiUPuMM48RkUdEIrYzRYzAaehGHDi0EgQ0cGDdZ/NA6Erz/Q8nzjw+
W6QfwRRlxxvdP8BJ8WUWlCqgak7LsB8FyeSJ9yPHiUsGAbKCSO+nAjrNfCoqTlJbPAsY4hLeOekc
o3ebdDkGTFe9mI1FbeEmKr06x5AbAW805Yzn6t/Qy8zcBVlKjOPMNSPUCkI/Q3wh2ALf4JGq0BHc
MoAOZ48NpEiKHbKNNXjk4Mvqk6cj6Y4urRpzbbdxVn0jjhA3Fm36GBUZgruFTGc9pXg4jB6h6Blc
V1RmCze1dCg+uHoFBLcmuWFbhhS9MRQACHw0JDQqRD697utr6icKrGVf/lX/ujNpbcqyiycADRcE
BS6TwIFNvDiPhrwVtyxLWecg3aww/5xgynyKA/52TTpT00CoiXQ7wgf/GXZb5doooL3ou7+9pIgE
+k4yrwP6okWyhaeNb6/AVC3fylW8LVkbSrM8Ia1y9FJxgp3DuNYbbzKQCceMeBjLGh1g0Z0WLWYW
ofayd4Yon5Jqq1qZ9yeJdO6aEKUVB7ub9Yi9UlSatH+2fd7rg+IkzAtF1Ak59VZjk+mP0+1PKy5+
n7syqQ4uas9ymDOQrym668uwFSp4hqWNgixLkYKwXTxa7Jm0CTGmzxYkPQXOcNpbxXpYNOR+LYSx
FXDcI0szR52jdzowl9+5OdSzRVD1eUSkNsc/jN8DoLUqq62HHr6tcMaA0GP3cpHkeuD8J0z676pt
iuDZfRkOOC/XexRfHihfFCk6Nv6j6LNZIzxGfL96sIHwiYAvw+3X+5FHyMuX4WS/fGMlBvgtduHY
9Rr5q4lHzyn1lV4mu3jJHUTjJuFb0h6dqphINI8IJZpZugW5dBblTW2TGHJQnrf0e535gf0yOcPA
ilcj8sRoRItbH9V958RcXbSmSWsviXWTaRrDr3MaVI6XZJb0ogEMmApudxGUpjVgiHO9k2M+CJiZ
cASSHo5wO9SPKSnw3lvOxiqMAaB/mnhOl9t6YFzYMlSuBM4w2KVLa1ejRfsFZSpNvO8C1jvX6OyE
Q1lbgkMMHPhRs/3HGTuBqIklRSlhuqvy/C26P37+efRz3vNtB+/ETIe/nuN1d55ZC9SHtRJ6NSR4
tNcex/+5diN1MdCNpGcJwj1QXThVzdPpS/PgXLNX75rkBlhsGBF6g5tc/dzmmKAvFpE/0uZgSHew
zQKwXHcvBht3KQWpfLhFHsTk2A+WvJ4rvUIUtQZ9vpZ8mUebUqMGNPtijzDlXL1UHtkBy2B9sm6M
dEF2H6FKD32lxKYNOes/RUgrA/ifN08TuuSMwaJher5vv45LrbVlDNB2qebspB85RsXCzUAHSV+E
CbXqPH19fqd4t8nKGVtzM00ADdfGHFSk8eUNRt3+5BVoHGwQIvtjsfod67TJ59R5zJxaIKIzTGA6
yRFAnUzX5pKff8JjTWOot+h23Gf4OVpLAJmP+1BpKM6cNMKX+wQs9D0MuPQorM1w5AojrBzs/WeM
8A9LA2FniAuLs3Jb9LvqaAvFcdoBCYu3AxCJISzvl1tWrdnTK0ZHlJCif+JNPatxeidZ8q4kJr7c
R56XZFMQ6t6MgZ2F52DWBbos1ElZY6fVMvRu2GhVcKLRQNUwaBV6l0ED+S+xUraKPUkPc2uYR+Ji
kUkdtGebR6eCVUE0f+J2A4JUOtt00nAW5kz1esACNTd7q+/kCRxqJrI9DC9FhUUyi5B7maQ4nq6R
GlAmEzBVLhNR29/hVmgNMwXBWiBZBj7m+HYN83MvI6fUA5dCFLSTv4+XDHR+RWmYUSJIrSQW/yUp
G+qWsPk9MAF2rDjdM/jS2HAHUKFuYeEsK6T8h0IrglbrMvijrBn4LgiTVhBd52XIIwhaPSMk2eo3
8gTSMle1nZmJsAVqflgdUWcl8/5I0tQAhnXc4bsRiePRfYu5vUQ/ACEeWV3euwp78BT9pot+p4ud
RTNKNw9Bf2Oehv8T88WRnda3hiQf+XQ7+K/AzMXcAgWEhh8ZEh2W0YDO83fsts9AbTZC7pI6qqWH
1/vfyKZvyIihUrd1uCX9kH+LJtN+b32Jb6N9cBH6AwGOMDq0PHVpS70m2t9ZxsZ/iI3IJe7DaV19
RgQCi0X8Q7Vg+54e9G6BK5Oz0jhPMeFtHucRcXfWih4s6ibPCcX7UnisyunYYfe8sxHO+zNwzAP3
lFT0WeixrLORudzm3G6fTjN8Tjai+lqh+IFruex6TZf53yZ1OzjXnKzPH+5tOUPzGJmDX6Zh6ZGv
SBHN1IEpwxaX91RAre0Gg9KY6olYljEylxBX1XfxiCEUFstv5GzlaH9Yclp7KzWKz05FEsg8ywZm
iJ/m6RoP1KPMgMIAApyEPdSknnVDDypIYnyfGwkc8AF0Cyt1p+iMMlAuH09ACTI6alCLHITzva68
I9NNyj17wl5xpSyYEcw+0OumMt+Bi0Sr0IABaDilBxeb725Qo9oQJbpEn9rQlBevJTk9NDON6faA
M3OIxqqQWz17Dwy6EfeiJjehEx0u3kaSSfEhBdLOb/J+53lPaFpu9X0Qz0ngXO5vuskLg0HZpQBW
dYDFfX+0IFNZqsFSsvtbg/kMGKm38x2AMw1mJ6dVCo9D+8pVaXaW49twRK6PEaRzgVcjJB6Hq5VI
OCQYryeIuMRl0ZpuGBO6x9G8DSi5TY2K1aPG+pSo4OjD3eEU9pldGTXkWYZvDV2fjI3NdzWpjp52
G4YC0mzLoQSQJfEDX2ekUPKpycyXlh0Ides0kZzoJoPGs6tezkchEOQL55kJBDlQRIwMVX5a47O6
Qkrrp7IfWgl6vUEqvr/chc2xy/MQCX9y/J4yz9DURvuqNCE+OEnWD5KGYJBKE6fwpBks7/KCxWyu
nWRIEbuvbREBeZuoQKaPWwVA8xKCjB6Hf+ZdrO5SeiSnBKlfpU+Px9c/5Kj0rq5AQ292jwmlAG0E
9m9tfjqcgymNOeQu/5WVdsCHsZvf5pqs81VdUegDi3uE/ngYncMyX++4+T/Hpm0yc87lS/CzQm1J
cRorCg1bdwrO7/bRqrReCx3pcCEJZBQvkv3IFcI8bA4ZC7C3tZMi7BYmbl+jASwOmO6CxDpArdSg
jXtHFtXoQ7gIVbzqNCLT1qiwZ07cAdCKioolSS0JuL6iakkRFWskduZG6lVd2MKrf9lUNuJXMjJS
STRqMze+oxPKaDVORElcdWtfqTLNvA2dm4th59EiWDlq3lMQz991Sul+2HpFxVrd/8co+ZnCddKV
tEsh2xEZI/uiLAwQqqIu+JCMznjQWwCRmyqNIwe2W6foIvnHm7LyhRsYafMjbnDUf8XYCqnjZcOm
E8LKdqi+NmekMQRtyc8o3bdN0CWfi5IaUkuJRpmIMawCWh1iZ43aB5VQ92Uh91ZVC0ErEUZVgZv5
SK+W+UGJo+1sy5MfeBA7CI1JUwbtcNxl7u9fiRZwF55nYsGn6dUqXxNAwIoQySMrUah6jtou7DCK
Btz/9LckYTz3qUU5yO8Cl4TBgDkJQGshR4zbCPPKDrBRzAUo8FizS1dEnjcVmtdn4TGfQXoimLWi
/YZKmckbFEOjEHU0AIi8QjYH8PSseOC+UZQ6B1Pn332MEo/aqYqElUjA7Ve+mBMRVedPw7jvxrI6
KWjQuHBHM+iP5oeNA196sLVj12MXPsyq/bZaJqWIq7UEbmyJ9g0+ciVdmUkTKbtZzibAwP8gylo+
3iFHsr7FJk06pxz3Ir4v3j7zrZfDsmAZgxt1eX08ss9kH+zxoy+EOZKMK3ajGbVrPRZ/J4awm4UZ
07Y2Vqd/GeqlTLsjNnXg2g+/YniZJkQzp3g4NGvoVfQpsU/lyxW93fo7BZGxr6qZYsByLZDp2VSu
PcnE93AlrzSizYu7xg73eAPDEtHGPFQ6k06Ds4c33/cuQnKjSkzzZ7ceLTIXXz4SitVt8p7Mm9CW
P/JQlP8uunGHQvk+cDl394ITX0Gx2bd3jildVpvzYiH7i9POR+Sf97WftsQeuuwwlQEvKBeabfHj
Ii+eqUbhCoNQdzsxSjXj5QmEGNQtVb/dW/elbGuAHDAMgzdf9BYNsTCyTbIKzRyX+psanQoknuw+
IyCiOYaotnPrC9kJCeaXiC23QOtslVnEh5pB+C0UT+kIYyU3vRgudOUZcmZuL+ZFDUL7vNZgmoNb
aYMJGXdDWY8sl0JV6MelfInuRS72/H/Snelm4dZw09qCJPr6EC8YRy2t+JkuuXBXRnahV6HId3Xw
CDr7eZhCg3OhAt9O5SSaUfh211WnjDDsqtSnMMRcb77hpvsf8YzX/oVYAmoCjmAQsNhYZpDorhAi
sHKeQ/WmgPPBogg64AaUGHLfKm8Py8+Gpbc7E/H8tfS1E2smZiQ68umOvsjCm3UphkdzVT69kJkA
xiNBpR85ZNB+dWG6T/4pRutBD/6jtcKSv9Uw3a5Ggh6IW22x+ni5hbSgC6tNtK3/mEnWbemZntHF
MbHkADrNtbGDLVt3hHKqk/mCplFmwUgpL3XZaYiGdtxKOXBKRhrCM6QNEzLc3r/Tznkq0y5eHrPy
KAv8f0KXflKvhC3jYTejtGZdJbT6otRw2AHq0gElg7MRwPfoeKu2mFTQmkqI5KS2OgVgJVg04hWc
2oth199VlVt/C46D3iifYkPKafTJdecVwmQr8LYrhCNM89eU3BJnwAZB4C3JU1Byw5M+nb6xIa8q
jJb6sWA4cq4b2XKCFPdVi/ClTOZxBA109t3jf1mK9vM75DkX2461p304Z5FSMEPe/BxkJo7twH3c
3/WqfPXDfUibdfQIqikOqNkAxVU1YUPAvOFxp/pceBctLLpyXxpEBwiSJ/CfmdUSq3qEHbP6pRJc
NCUJFhEVOyac0d3Dl4U6myF0hxn/6a/gn4m7gH1cB8xN8xXH9/w7gsSmA8hJZ0pQ+tZ/9uG9COXq
ZNOZX9UlZu4LwD8j6KC5oI8LDFRhzqowZ1ylW1kjMgKgygZcIQKtftEcvqY7ShnpDYute7VTZ7no
aDtY5O5qgDv6vx5E0r6PNhQ0Vcy14MJdXHu7VwzT0AoAcn3EG1eqm7kRdacnnxlLEAHZ51xrj3OA
aBEnSmz352kh+0jKqVxzvG17zM6VsSAXOlNZwST6dZj5l/LUJ79eqdstYavw+DvXSyDxhGtbCSov
e887TURcVob8tFLADrorx5A5k59mPtWoayrS6pZcBcivB7YcCpaMg4dzNgfD1V+cvF4MshvU8JX2
J1rMrtbsPEI3p3vfQNxkfKt7NBocwM54ouzDg1e/O/5TH7Ep9P4Y6NSub/0Y+TCmpyjrEXt5ZfVQ
maTjBAPPsOlbT1c7i4ROL2HCrcVqtMBs+/S/F902XtnsPn24wyw/jKeu9E52FhpvVJXXQbhfM1SQ
HZKiwXFp9UPI8GQM/35p9qjWJ+zaJSp3fit7AN9lun1v9qSmv+y8jfUIQ4jeWAmQ9Z1O0Bv/HONh
RsSDgzZj8pJJ99rsM3RXqgxReK2T117WEJ4P/cUDLQYcwBLGdWmJUPw6ulN9zEW8iaIrKetI/KNl
rSwT732H5pj2+UAhu2U6M7DTCOgmSv3LrqVn9nph9El1ku50GvZBEPoTd8B+itnFbtat3JczJXz8
/YiTiMbwwYuQPxhmKGBdj/nd7LS1RSsYpLzEb8vfFFBqwO1c5XLT8oPIkYN14SJ45Gt3a1dq+7ur
+3ohtCYp6WSQ+/rp9AYroChGt9bP9m3hUZGR5waiPp6T0ur7KpNwVDyjfH7VYxhHaN6lbVXzBt2i
tlHSqtrL+HyYTVXOKqZSEDMmu3y3SSwHdE/T6BL25dmFLC2LnWZPQGj05jYwokHikC5SzfIYSs51
EmyYKy89VNPyP+ttopfgDm00lhpU+q3bCogTII3dF0Y6U6qZyV3eaY6Na4JWDPLTUClIPTEXnIo8
Oa0usjsdrCeIsXD03ojaSCDF3sz7iuX6sfQJrWe5AT+trYhRtp+YprJ0onbogC1ki6w5/gGoWQDY
By92W92s+Bf9elPr+Fu8ggND5tHsFX6TVCdkZAlmn8+12qJ+pZflWl5jpQNgBRYeSRHLKpYtNb+3
qCt7jSvhxC7b5wBuO1DTf3Zz9/KG87qAOYRiEJGmuPWypJOag1czIroBcV86od4GKRqdJbNZRS/o
WtZ5LV3PN+GR0kgTlR204RPX40x7agkoFLWO4VKn3EleLv088gu0RnPSD32ZMJOiHOHuyBpK7DtI
M15AMczP7egEU29MsFwmMa2pZfSu2luL/7T4+Cs+46KJjbKCk2KiCUUZhxEewXfjZmH7PAOw832x
+sKejnNgeG2oHjV5bEBNYCKLbcgGCJJrDl+QiYB667BaAQymW3L2Biv+QlfTPTfBQcebgMbJ6O2X
aJ7DAjT1HH4G1lX6vXF16+NkVDlb8edV0+CN8NumImdIk3pK6Cm6fTTj5F3JXbSi837DBk155fve
QjpG78jZZ8a+GmoON8N2I4bNX/4T1db9TCJGXrliQtI6BrSe5fC3HjCjCw7o5KNhtOkDFgZc1uw7
8+pNfwlcd5lclBtF2EpcTt3OVG5n7DuDNxEqW9kktQA9A5Up4lYLSmr5n0f34thJpRRXg4t0qP5p
iFMjuDYnIAEnZkZ9cLoCPWotqKpEapY5QB/i4rKDB4OJA+DhBar5hTxDCX/3B1+nZxE8PHa9ns/g
S1vsOxUYcnYkUf3J0nm9y6iBfxHR3Q04L4nPVeYLn7MJvkhDILy4lmOaQSbPBZobV8FJjwfInnvQ
CX+85n3aBqZi+ihy9Xn7MgjKQfNCvj0eqW5UuvCX4jKcapcxpWBgTLFe7DGsH68F2gAaleMm9FMV
ab56FBMMi2Iq6L1/Hgoiu0ieMEKC0PgT1CkqNFKxD/2bKkpUXFp/lrQNBxjNXus8pXyEfdxzbnl5
DZ8vwICDdQadlB4zu1DMwJkquOGCFX8/e8rkgciCc/fE02qzc7PrGV+dRT8YlDp2f4hVRNqzFmwb
2wf9WHyQdgP2qIfAp5LRSIX+4FK13y4gSNoq3WNNZZOFid2ikxJ6uPCMMCNb+qV0ELk+o9YwMn1x
w+aexhw7lfYWRWPaTdhjdKZ4lH5056iK4xo6qxGAKyEl9zdgDbEsyjnG41/gvzSgWO+SXuQIcno7
p0GmE5yO5EmO/4a2NHn8R7a/mp2XEu7yxLN/Y4ISXJgzx8dNOihBbflEwaPDXlcNpT32jv2djRfd
H1Rjyv2kGCxEztRnB373NvGe1l0HzMdPJEhkx+JO5vB3rKakI56fXm9eNy1t1fBE0ukUiZBCgpsq
OuPQ/4yPzTtxXIXAQ71tchzYF4mw8CFeOF50AtA+tWfNF9XqX319Iy9FibVnrQNgpNB3aeaM/Cug
Vzz20lrsEm9MmI9v71TY0Bba3vNVCP+fHYwjC6Nivp0B1cp7IZSsVSPBEFeSFi5Z8W+nKnLG1LdF
PpMWUN/uxgPde96c9LsnuFRkveHGhKATIk7UsZ1kfe4NQqXINnCm3YHrL31DCnqSa8Hc/cB79Zf6
PuyHFjmLijFBpFbsCvwi8/Hx4uqY3BHiv9dyfhQ0knQSef9Qwb0uIp8FbH6ITcW+LgeJ9uAFXhn1
QmkBzEEQJEphES54zZrCKeG8sYQ31g92nlHHXRlPVf5Lmzge6T8I39RJTKAcWsoGEHESRwPgoukp
AvMmft1qhSg1G3fg9x+GcWrBihIY/QcqlpN9X7BVw1pL6xo2mVglHkD7oqiITUVe5KRkFbHEDSxu
wn875MjQmYJowpyZ8YKtD1Tyxc3ToLO7DIg8uTfm5dmvsd9egMxE5fwkvJWxYeWcKWwcone9kh/c
Guv44TQCJIWmUbI02OOd/jEZ6tp/8nRmQSimBxbUEnG8eV/SCVCRxI9cwDOHHZO7hoMaf5sxW42t
bvJj3OzQ9s2qvo+M3Cc/8fsFMFxdfuTnXvmA4vVKjbyI5ksRf8H+7cx6+RN8IF8mVO8XULI0B+Fk
Wrob9PD5NlAmfMOiYu4Zlx0tGO+Gf/JSr/bH64twJKkJh4E2cFyluqMfAnIrsMrC39wh9S4h4ZpS
hlcL0biOpvN5EFqIYSZ+OsXonro5wd7q1p+JxIzcPvN+id0jNUScuV4cavC+XvniU81DRAcsWXT7
FEMPtwHvvrYtMJTqyAWY9G7KoomoUuthA3q4CUaYFXSXljVakIOiyT2woaehbkqmfrTI5HQwyUXD
OTs7Y6tNE9SlpNvZrWV542szBO3X+kqQEH+HSTEi069/2BdTdZpcP6weEb6TH13/EsQPD+6PQS0h
d089S/Bx6llmvsuHu6IzgIcY+zOVTp+nDxBhK94TOfdJrgIlmTM5et1dWe+AqiMfu+JvLCphevgU
iqCiUPL7/M0bw8t7Lbf03Y8ghFtuNQi1E5/+pFQfM7uipasnf6gJF7CbYZX6eYMTVljtTo94jyOd
Z+N2UN3nRvDp4UqAeq59HGdRxx6iutJMy71iNdEsS0zdTLOYBZBoc0/4zba5mOPDQ834CLjAYVZX
g2fG8JkuOkeo+Nf/x1npgNSFZeXemdofBRymnwsBnwMDGlD6Tv3G41y3RPYYO8S/XQBi1fPln8WM
t28HN8u3qP6Gjk/droK1b00JTvHrtUas+5DQHuCsDrTsKn4blFkksL6Q4ATLmxGieO8cYnRWGRjW
XrTEmLSaoyz6IHOettCN1dthDlmvlj+8vH4gfJ2jvpWwXM6kFgaGi45VZGtM34Zy46R97lm/Gr0B
p3GaAAputNfjJYPhiYMreMPAfenoHajz1HIxTz06VeIkLlnigKJv4S88WcJvqCj8KNcxI7kyUB2V
kKb+RWKR4g+BXO7cNPuhEhHI3qX2BM+gA9/WPmbiXe356jem059X7xIpdxmT1AwiqjIgpqARrL84
l4mpGaKfwe1U9agQZxPQWqsl1hscBDd0fQGj+sZHEQfoomddB9Ff86n52MQS8Bd6bz65lD02Ts4p
GknF84MQu6vIMdIkGzNOEfqgCdHchJOffo3RG2YdXcR7FhDHF+USG4jUys/HO1lkmnqTcjOfwD/5
uWIkx2T1h5XjZEMTm7iaD7SJ0vVcJjfKBqmJrFWM3+c3MVpmdaSLTYuZ1mclRPt3Kkih0VLRfR77
+ko419B5xKp3taGaN4uSw+j5OKv+ygTSra6Ruzd0pbgwkBdrpk0D8cXqPM+eQUVE19wj5uIk1F/+
pOaSuuznqQw4lqxlXwtHfqBJXCamPu8X16WdlD/OdvICgMmeCd4tprQ33/MdfmzqLIKZLi5WywFH
4LtzSk0juX0x5B1cqIqVBxhXHxNv3+Ox9+Ny+Izn9zAOYRZMxb7NdObtL/JAcXHkFifEhf+zEFBu
bRCc37iIcjnchf5Gt2s88zVm22I6u0tAHU+36wQvMA4izyr3CnN7uzvyft9+WCv08cuznDPuDm6Z
FYbgaTx8Fe/ODZ29Y9PUn0MUnAeD225Jf1MEzht18RRdxGD35iNFJ+dlbR6NUmqzH+V59WRyM2yt
7A8Th7RThsdvHQSSYe48hyuFSKfJMQKWhktSRMvBcuuvVajOEzmJvs6MTwWunU31w78r98iFKtim
owd+6QjQ5FU+QD5yeIO302ccHwAPrtOnKY4IX9tD77fsXikrpfbhYz2m7nAuMwWj9OWZwmWRpzuf
804DXD2+oueNSiI2QfcTCKQqZXQil/vKszHEVQpqO9sBNNnqsgORzEVS9Y4ShcAHzH68eYsDZaPS
rkvmM0rPgv2M9nqyT7FG6mcWPHZ0olOTYff2bwjPY7ndjOT33ZYoGV1PiL/Xaysjqq+TLEX53ZdJ
ijx63n80C1M9QLqeA4oRNHbDUX+8tVEeTgK1aSBdDDTnHg6vjpZqMsl0oeWV/NzU8cQOdkv+t81X
+iHvIc8oCQAx2CiZluAgPok0BbXaeCam1wn75I9hD6KtG3tw25hNCXnneykxF/uVsWi1H7tWfTXs
f2JiZ8hg4qdJuOr2u7Nu7P9juus8O1DxUOTPCYsMoGEfF4i9Tb5NpxdD1Z+XTM5qy58A4fNhVNRk
Rj/CMGEqQF7KKDlyMjYAItttnRf4a8mzEidnaBWl8eSkLvbZ3M+U6jfm9vtCfGjLNCNERpfSR1tY
Ylvn34XhnVlRePTEDsXGArAVk4yl/+tkmPPFYH905xqnlivMu4LgM+1800s1d1ehNmTpx9oCITlG
3oskNVD7AG/PqCDScLIYhOSXqCu0NMsjSO7bzE1262kVQQjE8LMbYrb84NxoAk0aEUN4Vy0x1Mw4
EOsyFq8zOBHpXuqyG+Dpd6eEBlb/fguhXMrNOeDhO2gCNWTF5/AcYcccVCEmXWi9yeuzgY/faVIy
mzujYELmWDRmFyGxNoP/D64RllMHGOGD9XqFKTq3T2+SmjMY1og5PGJ6uwal1qjCZ+HKfzY0gn4/
5sogfrCWvuqp0SpKo/RCk65XTgB6GpdomcyYOGVI4Jlt0PaIkIg25P/xnRVNI8sqbuRPL5IKmBbq
nOf41OX4shVo2YfIMfQuiB/Y7lX2qfYlsOevjR6L6Ot2I5SXAzi2BF3x8gb1g9cjhyl7w8WH1T6e
zFs8i7KFtkpF7wO4zJt9s5+5Pc8p8CV6+hL3YnARIUDVt2xvc7KGuagqoT+iyk0YXsmvFcFwbPxS
BTV2DvxBOGRHisUXWQ7bhT0LVrE1Hs3BaRTcdZ1hjRlF+4VlupCNIuJLterEEHir8NJsPFjpqO3u
UXiKcVzz6cVgju6Ce3YjdeCbKDu/iqKTB7kKeYTTGC9TXNsR2EhNnDJA/eHiuYfjdjls4JQTbkII
Hzq7IkUngSdQoZhOqNsw5HB+cIW0jlEI1V/i352cx9aA54G1YfIm4EDMAVMJpeusbCIU2OmyBXfU
ZlCcCJUhq+KmBvQuzLKv2nhjbKVKAq4IAb9UfOYqYMl/IUPrvBAUP/fpIiJVkdvxnesfzEga7hnr
tx2JOgPw0WpRQkqr/+YwNKDgOtTqp4oGxR+4vHE4pRtMikx1TH+XnHWXH8Q4M6G2fS3rZ2D5Rjek
Wx+YbSQoXmyS86wW8Q5AkYd1SFUDc+XJCsmK4FR+Ja2Lx/ndH5+d8m9GyFd4EWnEqW6V13w+LEaj
yOQc38CPwFCGDI0zeB27hCrkSpi1u6yxctlDvhf0dxd7gzr6tUnvquIs0zBDD1OLSYW2o0zuv2Yj
AShM7vercodX7D0fapQYgW+jxmLWMBcSXJb1hs9zUu3me26vRH8Jp6+pJi7PsvupijRhsbecLyCs
PFK51gwzm1lxHi5R94R9827XxvSYznjnFHireo9Pw/GmSUxLaGKnC0Nm9+YaH3fAVsiOmije2txB
220PZd6bkABIqXb4WtyNBv9x045XCQf0QtotVBPg6Dy55FsLRQ+ERrocBTEdc5tHUxwHvmHNdNC7
gObJwVpxBNq2SsUT4EawXiSeMKWDKmCLzrlb1u6agjxJMr5op7jqUOw1fjXcbzals2MUbzsb634Q
mXnTYdVAV5Zrw/YU8ZbDr+VXuj4AFCzPHw2Hd9d84JNpMklGRhrBmKCvO4H+S//hDiO3K0bBWV9V
J1npK5yBm3Usz/2XoLEOhk/IeoxL4jWPKdG0WRzSgQm9Y+5hIWZofBPP9HWE2Pw58//LmT4dgiNr
/3GUD58vCF/ucT2ezInEXnkYYYNT3wV0pD50S2D/OX60RFoxVDmsJV/s1P+I687+Rq3LW1DK7Eo8
2KE2GTYFZEx6uRPtyN7eGuZsSNno8Z1/42MXnzFUr0nF2vgRu75QAncdaNJloRRt9GgcxOmPlCz3
ciM+f+8mg+s1lCU89Dbk/SqWjsMCltStmXFMqIQ4U2nabh9KeTTODcB8RBl5WjaA6kUmSskEnkOH
Vb9idIA9X4+FbebIraXg1jRzDwY8ZMztEDLDNsO0ayixBIJJa9teD+IgKBYJ93WhFs9Cz+dli+Jy
IpQjbnxxiwyFeTVko++Pb/5/DTXgy1U32LF5GPqpDaO8ja9OC931Moj9eBpdV/22/RR3mFyQgulN
kVkgidHj7Q1qRazfGEO99lhe8pF0tHxm26LAPdoEl9IYDUyBHGAywQu23LYBIhyMORtkKp3lGWNs
HJN27JQHywFE+rOqDH7ai9gXreEKXpkYcv2mIk83FOKnq2dEvFtLUjr9DmgItoKNwDSiizLMIpTU
1pnM2C9hLFwUcHI0lfL4JFwO49hYLuXLydAclkcLUVlZBEWvP1X3TTMRbE1g0dQ3i46NJCVNjCc4
H4DyygMEx/gSVMxeZj/xAD2VoOvoMHGRt91XNhuyO80cFlrKHT0Z1v4Ne1NwXtMrJKIRsnGfGTVg
2jarH4KEd7Z+OsSsZsgKf9UwlQyRtQmi2LU7kWVlRBiGCp41/RjIz8bnCR2y1vWe4ralMLIW+jsh
UEwQ87ejpFXe963fpvDYdlvACvW0lWi2YpSO2Fs6WnSzGo276QK5UJM91dhAG+Lrgc1QVzeFD8SE
hCG/LoVMXfkhHIR0vwg9MNlgnmnPOm70aKvKKeYCDWjFjOJ8UXkeyPWJt2qV/YUx1KJvbGgmj4yF
wK4MkKlElo2gTQdnUyWuz4uQ0GhXl9u0S/LnwpNEz/yyuUUUgfitLxecTUG2MBu6GYelhv1WkdUD
74nGwcW3eUK7bOEY3w8wC1QRCG3zNB+PKEHMkDDp9QIzpnTNSp/v8dAvZz+1K3qU1ReBVfVnWCK5
9/jaCyFRfjarHCdLQRrswBS/O5nAOtzQNDH8a5DfMBfVv1KWZCBdiPtDejznn6GcSjbx2sVQ5cVT
cNhLprrgdt4uqqbebotqMFvfChnigWViIMmBa65koOHRlqM26obC5X4BXs9YiHPNA0gfEVqdBMwG
JDAjkwqiad3ByfFMCaMSp3aoCEJe6L+0sNOYPqFPKimLHizWTUm+3D65u7nbyni6FLuALTmmTV3H
dvOimridO7jTuNpicBQ1oqUOS3aXv+rvbcIxoCjbJ+ZG4NFAOwQ+9KD0ESj1XwY7ycG93d1PJxXN
fusJKZ4RE5HvonWXFLq8QiNWVFWiM1Br5p2attHmI3uz3bUikmGMFDR6jvgxBL5vq1QV0f5gvTKC
7P4g+52jBPnC/mi7gbWtNHGe49i5Dor/e1XN3Sa1PHs8A/UreElbF3FmiCyYybVKLQwgsdH3U8mG
irEtHATvlidpJH37hW04n/Kn8KtCrumiX9HZSw1q/IQm4gOMMsqlHMaQilsvtS29mpOtcCPSnbzj
Jm2PXXAzPoK0vpip8b5JYjqu9HcuiSzum8v0P4dA/vxuaxv0fhA+VItuHuUEAbwiRGafCPH6vpJa
tTBtZKNbSgZFnV4znvooDdes4jIFdOBTXLyRgWhoslndfb9VtDLmzR4qP8fsg4kvYI0wokHsZNB2
lFmYqft2hsdBRAkQgbo4mHemo7ndha+pGDypDUws4SCdtUQoY5eaSceLsp+b74Oze2dGUbu6WfxR
w0zC6akPzvPKQCYMm+VwcGA7T7bxUv6XZQqgA80QBPxYe4yi9ZGvp3y32TAhgeIfHgvPF80pIZGX
ksAehGeZbiZNeb08/gdb2WZX4uZWoQkwHYxVZV0ywcmynS0cMoV2hyNEQpKkN+ZI9JJC0xmGkhN2
yancsUnXnVUkiRAyr8O7LuJQuIU4Hov4ZY2rgfXj7DJOxlatKtmznzPOFRqgf9LEu8XIf8QOxIv7
teYrs9u2ruwi1m4eGwYJPEWcDeiAOsNElOfv0+/xGPjgi1exkQak/5EXS1GHT/AevI77AITSn0eB
+YKVSrQ6uanmp6KWSfAhFarHwfCTWmo5Red9R+hZHt3aO4Qm3QH/Y+vp2Zd6fw89sS8/IXEXvA8S
phUiW56ihAT1Ho6A3mV/QYyCVP/FeQfEKHVQdOM4pNauJzIZOZdWlQrR4P8Bt0wmBbd+H/SvWzeu
D/lDmhhQ520k2p7ioNv9pu9QoFtzjdLMZt1jrTiC+yP8yn4AOStAbh6X5Z4yMRSV7AfCa6B7biQo
EzuxgpZKDqd3mYElZttBDXBrNf56pSw2aomyyweRUFELiP8TMFJB4nAYzytShmh7z1QX3VGRcpAr
FF2FYbh8If0aH5lp59PWydsZVrqSpRLif5wl9gNEl5YEci1+2SHiCceDcvrdBdO1gl7COKCFq+x6
WKjF0xGNR4HRNnbeCoNuLTaa03F3+GSwKbvuB9TOT9VBNaRSO20APhDBMH9b8wdgryebNHkC5b4m
WPfZ6RiHRlDSDbOIpj3/BXHpIRTq/Qille9sGjoIBNng/qrY1HlzwXfi85i4LJ6UdIgH7PxYz8B+
iQOhfvx3SiCPR+T6fmy4ky/2zjLEST+Y7KRpkTqiEf8FiqJnE1yjtYLZH+xKfCOCcraH9kiZEM0U
G0GSDIihoM/4AFdaghkyrkWLQWvYrqwobQ9losNpVKXzcLJTNMIURzkO3iElcjM4iZpQTYsz+DM2
iTHxnJ0xdWGpOi0CDyN9OzT9h+svklDyu6NN454SLMDdUi/d++5aNHwB4T1MPkMK5MjGyLZFr2rO
dSXukq0PKdWDreNuVu4vLyoZaT7qeXPYqgkZ8N6tAO0WhyFBzZbGUHzvQTEr0fmOUfWoDVTny7OA
e4KltFu1mW4A24hPfsuua19NxOZMfWWw2sBUBzloisq6RJ8Msb21JUKIpcDQafXKh+KXBnE7pd4i
5NjRUcgpVReWnxKOA7Yv0XA5DWlr03Iu7xhiutN86MA8TbvZvUmd7T9cINCd96OuIJT/FmBX4Cm6
5upGpmjSEJpGKdJZVK9DJoOi258QjRS+9cC20/Ougph7tHWXb1kUBjqBR9xjGdiGXbNY3mbLwGvG
Tyzn0cXMb1BhvH82Gj4j2ep2Q94qtVPN6dIOlFWzPlhfME1ySF52hsSmmJy9XHBEStwLWUo9jnxh
pBfr0HJ2jhMPRPECIvweX6EKfxcHo4dikJ4X/epdrVlHw2JADAykMOhXat5/pqe2u3BAXqsQlvdT
KxoMbX3qxdUH/1m0SgeeFRVCtLJiahOprAV+LReYT462goGz3BNKPcW7cYxnDWfgoQwtylNiIXT5
A0HqGU0NYw9WwjTjNMjaowZwmpijPc8tnKwYAH7MeL/fr2RGt9lCc9P7wl/JyqgLiS8arnZ9HRXJ
TD42L6ps43HJ4Lwbonk65XjwAMp6kjqSlm+SxpwZEyF06GXWkMqHBRNmTlQxWYTIbvHm4wcNJYQy
PpkzktXE6C9Ph1b3+rgOBHO6UNiEHh+Jvd87padOnOVXXHV9J60CAHwvaF+8xdewKgMCfys7loZ+
VE1xCstt1XDTJ0lSemk7dorLFA2EnV9H2mIDhc+smJi3uGcDLJ6oyiyX1agL8rmJ/tNWi+xe8Mbx
uU3G08oKjzsbmxlOhkwy4PpOaIyGpOMwgtBsNIJmjf32zpKCfAilDrSUQ1HletDWE3OddsludwyB
9FMAuzTe0Xz3aBl5XRwnrd6O4DNW8T8Lu0w0QabDBU/YiWjGAx4AHf4WKVZe/y2rQTPFvDH5z8Qw
tgpBHedy87eDkd1HquKsoujb+bG71iZKyGdfLESLxv+fXErsp0rJvwpIftltyv9TR7KKDMMA4ezt
WG9cXdaf2kDqAHhRU5P3tGFIswhL8+dTrGqNc6PlCjxlOlkbz6ZnBW0EmmrHmfUBHLKQ1XDcS53o
HJqjqO5XusgXxF2S46mtwxvKBhYhfcBqLxgBB1SmNqFVX7wPKOBFe8ovtLqmjLmGGlps8KWsj1q+
DLtfgdESIlKQ7gjCmfNXN0HWL2Kd9gdB8kbkNBWEiJvb0lj/5rCN3oGAqP5Y6SHC+hgllF/gA7jn
SeKCJlo+Gr7UIfFcPtWMkRuy3Eu1rOUmvKg4EoCSPVA+Lg8A6sVjB0+kQ8duYN3g0vH7a7Ll35qR
fLrles7kN+oCkn4Qn0kLUPKLn2pMM08i2PQWZ+UCmiqinwJwTtV1jXFao41H1qVRAWHqgkO2GfEx
kqoqVIOp0VrN4w9IQUx4UaqYAc1Agt2WZ/X2CmQeJqJ1Lww81cALiQzv7bbMfLlnAvoA4a9xUbBG
iFPvMQBj40+Z8gJCK3IRjXAaTKS+HCEGI4FEok9C7s7UJM6rHX1Z7OpoI1w5EwRKPnLT7bLES7zH
B+UZAVFYfz78N0hYTNaC8xWJP0/EvRQpRYDu0rQ/7yR2+5hsqC1jB+zd7/53j+MeatEtwV/hj3e4
uXLzHJQxD9E+3QqeeQJOXgGdo1hX5w7K/xcx2HyC2GLCdnp43nZtGfRybhZDfzlSE+jQehZrfaJw
ER4j79ZTgamnqAymHOir7PzN6k9rkArmsPKlEgovPyYeRVo2rSiJlJDvx1kz67eDzCRIxvNlzZqL
RRWQY3MIGxAuDILJppAkJBOgupjhPKHGhWgDeDmrMPZ1n51HvJrahm+Tv10E6IHQRw2HTrauziQ3
WaDCbRsHd5X3zTmTxaFslr0S5he6K1R1oQPSLG4XxuzZU0Uvre3COy8L84HWn7obmUAjUjFrlUaO
CcoaAFfwTdyeljK3tjvtCsQkrxsXkXsvN9l/yJYA5F1JCLy2HDJYEMAmgY+WOOLi0z8LPNcJdsiU
D9VJZLK9NSITjxnL94Xrn2GTfVTyTN79FDzcKtW+S6cU5d74BbkhU6b53Am4I+qxE+xzJb6OGyWb
gRdNHE5Z01R4WjC/ilc+iFXR7dgy3ZuEm/4AmelruC7VjOJXtFvHR3Z49Gv1lx1GjBlkJOw3jDsc
Lfku8hByjmxmkDj/4oHUTdR3J1R6B2u0Th4QZbEZpRlTAlUBNmbmAMiAA80kmSWrbGer6mT/FRlc
oab/onMtFcB+gITPwYvi4Elu2NtF/t3E7Gu2bT7CvzPOeZro3Dk2wbHXikHiJKCdZy2df11XLyJo
OPRzHNnZM3oc0+v/F1OxXCHbZaV5WGqK9ctV6WqHRWEMaMzECu16k37zS3bZCuezS5H2DAikJq7J
ptnbB+gB4N4V3CUNbXX42qRMfOyX+dW/QXw/R+sTpp/53bQByraxb0fQUEoG6uyikN2ZWaKM33eh
uf4qSgroPvX1RkMHnPDiwZ1gu8Lkw/knYgiNcHN+5b7nGtiI44zuscvWKj7WnihlFLGXbZcdT62L
BhN4FHLolaZNHac9xi0lWgNsZCaEYh66/fbtpxc6fslIjmRN+Ygjs10APDrsbfzerrO0oET8O2/W
4OXvQTfQGpvBS55p6/FtYKaQVnjbs/NgVeIBHX12WfZyfYHWx3VM3bsD/w1/v5J11jQCrJTa3N9X
oOW/GwwL9YjdeVb55uvUFbdU2PpGQBEg/SuyclrY7/kesI4bUp5PFPC5bqAtbrs8zetNukXEQ9BB
YCPzRHGZSUBWU81yiJUdWEd66yn8FWai56y7M3z92zIDQOXccNYimJHgqwB0mkcdzXLK0IioRDZ7
PcJCncU+EeVwltd/6mdOYNHH0FaNezwl2H+8y2fR11C+mDYf7V84DySjMZeee0wdIt6MBV9Ee6iD
5L5g/JipG2skd9l3uYNy1lqgJL9vWWfNTsocy6JKMXP0IWsklBxCynZOq9Y5ztsCxPpGlcEcjVe0
9W6j5K9hinQzYG99GzbMBaWylI/pDiIuq4lPLmn8udmxRHz9FjlJ9c898fL5vmHchVzUejsnvpi+
gP1Ge0xNNMPkHtdzSwlex81tpSPYVbzM2hk/cbinab1sjOiOCFdghehybpJI+OY+Rch4uc4ci+u/
frWGbrKC7W5Y7dW8jp4aUCL8RJo47+ZzMYp2E6WnYi8SUB08rjL/em2LZeoz4p4KkXVBUwnQvZuq
+WHLQz9yg1q4C0Q64aw3INX2BYDkvcRE7GlXndXfvZBOTsOnSbezrWfUpfr5BZhRqvb5k0I/XOl6
LfifGwb7ZlAndkj2zvufncPHjG2nX3XiwHJ8aaFK0lK06VyyzDYGhUgpFFeOibW0maOJBUq7QXmP
9P7hi4FlZBULIwd11Md+1ibEM379B+RF9dBDDG90+jeGH5U39HT8vXZw/fX39VIAjBTks87Zkye9
axtlxmKqkU2sDXI51iybX0zkfPxLeYQuWpCzWXvB1SWO1ChVA5sBvg+1GYF98bTjkYPKvg1Qa+vS
BKwjPjysXWcmqP43XqJkNr7PbGVvW4HojCOkKoUZEA8YNeEzmeDEX2eUiVNxzKKNp2RyzMjuTtVZ
yqV+vFn8MlYw/ZSG84/drhlKhXHkQwJMBbINgvJbFZALLMSUfl78jRqJo/B+SkXI9DyKKH44kGHx
Jd9BKt0CAx6qAEiCGbLo7BfFpqDYOdNuq/SIQeMtFlQ1DIsucOB2tNDwCzSekC8g/5ak/KJztIe2
nrQ1pPo4UOBm4/z29o3r66s4IdCxpdc/UwRqwN1sZCIaah+EokQgHjzeT43ZPEyMlZEYLvVPkehb
rc7QRz90FchlsYYAOinPnrFT1Gr6OLy2v7ZibUrcRsu9i2ZBK8lFTzVK2LUHB28x1AdfxSsBwgR7
hIQPBPC3wa90k/ohQr7BTJJce3n3yRggHh/ARykG1QYIL32PJbeqDfwpC38J10HhyadKxd+JTrKU
PA8mSdzbRnmHPoKUAreYE0mBOG5O1ak+3yMWjM55pRQalEC9WVYouN4oyrMZ+B4YSWATJreGkfDE
ZAj7S7Vh3JYquhckOxJo/orb4bASbrHaWO9F4GJjkS6KtY04YhQ4rH9jMyHOGFDaQ0Y41lmyKstc
MmXjR6/fQ/kO9IIRWxDFUL35fzHHSvtq1Xlo52JLb69HNd4PXuO3Ymx6/ly0jjgSEknCjdeR6aXd
iRCGEmjMTaAZ8Sp5l1kLckFXIYgp1rshFVtenhOOVLZMIlnCytN8yNdqzJElSOhTH5cZ4VLhSvZE
Mex5ot4NAAuskgbD8oOLCMR+LjKEprPqTe1c0TMiIX21+fRxImvgX5keDdJr65KxH9Ds19rktEqI
E2Nog43pidELQicIK8aiOKquX8FU1D5VX82732+1uII/zrKZJhvD+QBeGqMFAWSja/MRy5SwUFTn
XOEkluPHKGZLfBootUqnxE64NgVCbENlMVVluxR9Ixoy6eQzvyzq6ocKHRM5AXNRpvqlwozkWPMu
gJ8J3EjCcAwMs/C/yz9SeumnCC2rAc/B9FaY0OkmRp0qRR/NoX1J9JYHP4rxE9OQEDOmgMuJmNUX
T2HVLt+btwpYUZzQlnWze1/5BvCoL/xg/pz9Ea9EmyNyhBBnaVy2Byh2Pd7znjTrHuUlrwSajSfA
J8Nb0urDUarAnvyn/pMkoyq1CCPIDedL3C0DPSMsf+QwlRtPrGgluAAQKNgyNgF7EoLRct7nhpsH
Alb9dC+Eyz1QLiSDcxLfktxrXb3JFQCBaiQJ5J4LSWwMe0rN0kG68XhNGWhu+uIyvio2VaasRZpb
mBCgNG1ff15QMMPXKZdw7CsjAwxg0SUVePCYLMseVMbxVTtj8xD2on7Xxg3iiF5y6suQOdi45J4F
c8MVuwcs5AjXfZC+uCy/WKgwb6zqxYYa/mCv13DY4OfzShumlruKubLyn14w0963KD10p9J8JQAP
b3wTJBw70vKF4br4vcPil7sBOQPo709z1lcvviF7twEe3VBniHJGPfJ0T+iqWLj3ubyr8rO5kRUp
riUPxK1QAyq/Vfhay2V0fRFQwCKGQsBmsgkMgYDQdTiegoRKZOk4zy+3MhATvA9oCDYtnatA53Ji
zvXNQR4c8TUgpC6H6f/WWwkCI8v81mgaYAuFEe+N+G+MEeku+GGMbC+hkZ8WTd2340Ly4tStCyi+
hpD//MIyS4TZCwUSa1x42RivAHDO9IjEKOJ0Vvn24WtIPKSSW6orvvwqxoxeb0so5aoJJehVG2vL
lvG8mYcCV+jbxljQ+NdItur4hYsrFH8p6A+63vXhhXveqoKARSNIDlz6NlHrWg6hkywTT/6vOizG
1hhNeJBcnLVURLnI9duNYeY7nX7RzdoqrVw7T7MTpslvNsth2hdrOG9PAUSDZIc+lznGLMZHoxNy
6B/OUgWrnHx/EgpZjTBY1+EGs6J/IOQMlg1Dhx0djYryCL6/R5WyPSDDy+ILsaULglhHEBJ13hih
UTX0JknHMchIUivfsoeJoMSgVYOctj0TOKjlN/OTKZLya1DpZ2KLBXqNZiaAnQFnehRTKpVIc9/q
IyQLyvaXz3Uv2n7fNwBmUDjL4AYG6ioyeYptF3JjProi3o24G185S1GGWUHOAYerJxBsYW5ZcFyb
5unDMBZ62U31HW8FEVX2VbZmil2cRcesublfPg/QvUbbBL9KZZA2DEDhTOOwP+PzbqehuSo2/cgK
sNBUrfxmWZ9XSyE5l3QJyN6+9cSYvhTi+NH8ABYQkQFeIr8v7fEQ32w8yuirYWrx1lWBl3p7FiKH
sXnLK/q0f+vwO9NaBCZXOg+MFjZu7PlUGeJiA4VoVLB0PZ8nv/CxPgQHQruERoNjLlwyTHaJ+3Tv
AD/fTsDyzuWxJgUst7tgw+AgC0o65oXQpsY42OZFpNq2omhBRUy64hJ6PL9gULRLSpG/Ivsw1J8S
/KE0fEE0NuYLD5TDoOTZv2p9rpl5WMtDBCdjzICiG8aOlbEjSVnlrHTYZtz//Xg/UQ8h1SW+7ybX
9JHHXRgy0yWDt1rVPT0EhTFjC+sUDuFJM9FFF4CaDvNtdcVLN3fuIIRBHNPRvrR40+QWtMXGsSR/
FgERY7mzeHz9Qv6LGyB3V02jgNaiGFb+xuPobwnb146WtX3BXL2lASZpivSndQCubu0mE7/G4oG5
8ligxTFcmuj8VgG+uls4Lvle+X2gQsK5BJTvlrdy8BfseVwXgCsnGRWM33xVCiU5eX0p2+sf7t9g
3RCb+W/iLubSj+vgwQv6qp/0/+KgUxJp1O+qp8GDoeENHuWJYvfCHtASGozFhfgwDHHSF418Vumn
V40lpnkgfuusYqC65UaXTIUShY/bGrYbFi3APr7BWF6pb8F//UljYDtJH8GOkeaYmffz47OqRt8t
QdkB77TWfANTvEhCk0tIcn2U9qZi0eHFJHkfIqF3FcyWIO/B+KAqiSgH3vpYesdaAAm39KiHbIFR
6lZyk6R+0on//Ht31P6NAZRgsD/46eIqZT2AAOKBr4ucMy8tVCRMAnfuFuc4RoAeWnpsdpKHSumI
TYRiSB47rXi6bcMdOc5a7AR41QiH0pOQn94gJtpev2+jhGKMLb1vChwCtPGStJsytHRQkocrbH6g
YEaIhXed1cqi2T6yCtclGbe+4l7XzkM7HlEehNHyWGBQx8/amxTz+IL13ed0e7gocBmVZUx36v8A
wDo+C3DT+S2iyjqhSRpKNfoOWYuOwRPBSwasxJLI3wyPGncCSwTi2YPwGwQLceY3xI4NkIk2E54a
YtO/3Vm2LeIZgUUvQRLYLKnCTmPHmYt8/sg4TMD4/SV+M0fSTBBlcFNfBwvpT0FVDQUnLjSJOw2C
8JYcfsPPpKy/SqOEjOobetenhVeMW7BZchD/qoHjajidq/1Hn2p3h+l2zfNeBfbyEF1HNqXGUUoO
ipM4T/MgL4TsZK0NRI7bd/skrQA6WJ28QZnRCqs329mcZfG0YQwfQLcDlW+L5sYh+1Hud1i1XUSv
+MX1UzCEBo6PodnpkNi4y0EQlOS92ojEw3mWyX2fRmXXFDWKqF+hBdJX2tTYIOlxWpg/zYY25Ft0
zuAnTN+wVkzkTpJLIeZI4+phCKAx+7w0JduhF5nmo46z+k0sdmRz7ZTtpXtS7qgzkPr2kGFn05Qt
UZeP/QypU021l8wCImk29fRQJvPsoo5+SAz+lGIX6jMH8/xD5cEum2VKKouMxW4MXJAqnOu7iJdk
CF6F9LKMsG8tirDcrN0+AIfeWWcsrFLxR6eh/oubavpBk1jh/HMJR6wojrURaab8Tv416Md8GI8O
Iol6k+c0F2FfR1TRVWbRb5PAxljmXQHGw9iyV2iUd+JYlNkKAJk5j9g5Q/BNJB9mVANkxstWqGqu
4OWiiHBrk8wRWllgezF94eWREf1GQPm+hkVFnx9uJj91XXzcfM0bCrINr4D0BXKxqleOkMe9cVCz
EP22yT1lofF0zrgQcMdYjiSH6iI+l7S4quS30JK6rQ0Ny5XklHq/CyzUrX5CaYYs4EpIO0FVeXfz
KRDNly1t0oCmnzPa/I852OZVrJiDifgtAwu1+gUQsx92v+UtUSC8xrKVQcr+yLZdd6Up72z6Vum2
ZC3Edt8zXI4PyPvVRYrL4J4uYyVaknu34yaWARS/NoMyLnDKZILG/tCoXCqaqej1konuWqgGwKcc
J2j7Sng1ykhVuDUdb9lTOU85u7z3ezpo60+wdEII5a6g/S5f+mPxLjFDXpE0ZRSGYz/qjspXvg2X
kKjO10D944tMLnCnhTbuoYYNUWD/my6c4MijwF2isqe8l4AZrKvTw5FJNImKOhG9kNF4URS9/kI1
tt8cQn2NMfDWWl/4Xsd+B7PWCCSQ78B39L/LBK/ycTlhU4G1336Eno7SfULrL0GWXBKxFT5CCtTj
gS+qai1+qLHIQdrDmjj7JRGPqmo/9WIXaSz9cb4f20CyjMY7k5cEO0R/KXq5Vo9xH3rcasoqYRNL
sLBxk/P5HY6yjQclOCXdRj8IUY+79EHE1U+0+w9IYU6OYWe/rnvrVRsT2NtBZFwsBORpvXmRhZJR
8Gsbea105paY65ze5YbgwV/IEmIVG/0CrV4KWetiS9X4YPDxIBYsuXsq2fwlRbhY0ycYzvPrp26x
7qD0WIecdY9f4q1miqOCRGg7UKjd09u/VYT5NhsvQIZeQ0Z4VCChv1uy93uBp4RHqzABZaC6rEJV
dDC9HqWyDGgr0FfBF39ttLMlqYEULICXnWKz5hbhScay76UXYYI2u1XvUFUCVMhjw51fag9gJ4r7
UHQkwTk/Ys/bxzMzm57TX7BY+ydUoZIzV1nTrHpsn6ezptjRHcwSrmmddxktgCvdq+J6Na87mpzj
O3GwP9cSou9gAwvk7rCvqlG07mrY/NXg97PFninjk5OdlNlFu2PkciGwSh/mYtqlyu6Beqf4vCwb
ljMy4ZqDlodBbKEagYYGP9Y41YBtE6hybLtZguGAnI7rfI0ZuUrR0eVh57rv1uCxh6IOdQSlFkJZ
0FoFHDJj3J01663sAhEfNAMIRODUyvxY7P2ksMi7oBlpfm0rOqTbCUjkX7Qpa0r2flJUDpfEbpkU
Ilu9aXLsHmS4z5zathK/noTWe+iuzvC7qwVQ1VqJnfDK/jPdQexiw5dQi6GR3VRAUcAOFmKI/8tQ
PTsHCu21AkXP7mU6HdEEeJInPD5/sbBHSkup3hlRzlXPqOJUb+ogK7DvcI1RU41whZuaBU/t2cik
Dhtcot97pN8ccD+IAuaG+Rf+yDB6ickWk8YKXf/2wX7SdEI6ozuQhPGrBe/h6mrqEsKn2MwXPLHH
QKlCJmYwN/k2y+XV/miuTAOqs/hKtR4AiiIpap7cwA/ZDzrrfo2opIlhkNFJi2OTf4pLSyfjCqle
6+nn/Ws/oGMhQ6CSU2hsR74BKBjLOQ6yAMN3acLNtxMWLraBR4yL4qU/55P/XbXTrrOhus3okXNF
ltmFDmWDRsrs6bO0mW/L019kIisUG8n8qcvslAwhvXCctHx5YvI5xtThOVmj6AIElAxbN3xR9mjF
b4eSJlEkjxwbizpeRCTW/Zy2b2xhG40VYgdudd22ApuvrR1z8bLWlQhc6JsDqyPmxIo/J5NPDrsI
devwh+PLCjdCZI8yacyJadPElAavKj2KCS9gVPB1wXb1nGcboGeYQtVwQmavx1TOtAoD8z/2r5aI
y1z6oFIkrxTyK4PZh3hR6l8kvWBTOrJlJPUQWEgnr9cJYAzh4DXbLMyjyiSpf0pIntGKIxbvp/5v
cxnHCJ5iPHppwyhdshEGCerjXxD7I9roRQj+x4VSgT3+7R+iAjSnnDo3tAci9iKOOtSR0w/mUNB5
mzsUuWvZ3AA60NIqGpLhBeVGhLtQVeR+jg6LLnv8g+C5u+ppnT4US1RdzydRjXxeOvI/b5S2B+6W
eoWCj21bIaMQe4slUH/jo/x8XZUom/45RJRdgoFGbk9jegG5UJAV5kiSwCY2UTen2F512H+tEMbN
95Q7Mlrw+jgec1MhcV8CQpJeHs8pP550Xz2ellMvKgdH+Az7D9ILnF0O1bZ8Nsey1i9aU7Ocj5XP
YxY7iKGe/UoydHBqFUHy89wkreND7kCJ0eP322/pef70gAGaoM7P7ZSicne/g83YxortKKNX0EJ/
VQsD2rzS1UNd0ZDVS/AWaL73xdKAyYV+gaFRn9vJfnP9u0n90Nn4wf/xDNkISPiqWIztjgcu3Ljs
9VZmriXERl6H5sB3bRtDqWhc9lHU41bDtM5X8RAA69p+KMDcKgpeWNXtWZev8s4Lxsok2fnD6WKU
cTP4nyyNxnA5sSHdrvAy+JaS+RL83d7QQzv95XtGrSz7SjmMbH0DdwxIqyItJ131qM7Iv/RsHTWl
ZiHG8NRnQ3miVF6nH1SNf/IjghbitiXgRwKyrEMetkmyiOmWGH7udW3fDbDX+fZTZF7QlvbuJpBk
aKVXq5K7Q1vtsJqA0jP+gXH+kJ1HCve6pY8BIpv5cO8MAGfA+aWzM4kB+k6j8sdO2+VNyQn5M3G5
juh8G9xGDnS6f9peRMtoZkejZ2S55rneZ4f3CTA/6m2YZPHG866YK9h2tmiPALllpd7BFEgq+jWK
TLLSVsWsUa+V8y6dbEcfG3n2fffSPdG3zjXD2rhe9E94/u9ncaZuhQeJf2HtCu9XFZPWlDm74lvi
lQotEaBCbaOj8b/hYma8BNg8F3w/y7K0hyo8F5cVwde2KCyZ++rVIoT24buLTHAwTvd5mRQwMRvA
2NF8dU7dmN6++buQo0iGGgep7dXnj4rrki659lzKtIzV4bOrQfRfRl3MBRql+vsEJeunLXBmc5Om
vY282L799vp+Zt47eqNl1asYJ7u8WtwdgnyRG5xZopT7+B3jFCR8gZETQMxmEP/urqvxAhTcA9Yl
21aJmswJdazKGpA7GtflyQEbw0U3/GLz7Ds52h8JfgtrpWiIuaeAFuOFGFAs/lbByk3LfCY6GXoH
T8sOP4bgs25u51F83hmEEuPBwgzvi98zFlZ61xOHTBsXE0XvviHCQlDMAB/zrx32NGZp/4n9W6el
3ohvRJCruFgFN5glGsu9eFMhIgfIXuMksprlBMDItq3ZMuei4Q7zDclcx7lVDTzfCDFyZWeRlvoU
TiKHlkWgfF9B1E4aPeP3VVEvC4SJ5z4H8rNi5t3wdBNIzIzBN2pdUS3HGvLBNZ12C4WQ/QqIhT7+
6Vpw7lnsPM7zksIFksV6HJvFv/m+8wOYkaxnHIvNiKneyV2ybVvAHkHX7ROUhkJJHmm3hg3DiMNC
rprsfNxs1VCQRYBLPQyEG0FdwoMM2fS0K3vbq4rf5YIRTC9G2O067vvyz1G47q8vMnOrpU5hRlTI
7RXHesxahSH8umvF8Rk9tr4fo+rITNLP3hgm7r4U5rnmODSgCl0ORdOrfZvsKL2AFLy90xl99mRn
rLzdWJylenmB9rq3HFRNKh3/1/b4P9ZxsdcCURB9+AjgXAMSn0SJ7UfkllPB6TAj1+/ZdeDcNhtK
+jApCRpWHiT/wYnvtK2qwNdtIRR+OBf4dK9opAKsXBhotlVPacCwx5CVGpwnhlr6yOYxDxUTOSuF
lThyjPsaMExSjf8nACTgrtwhFB+cHp4PUz3Mk8OS9iZCszJb3J9OS9dW0WOU+ULFKMGdKgLf1RoF
/PHTLmXcbiIu99V1OKFIUmJjzFotKbh3zFpWgQbn6JriezBavVS/x1P8DVFkY6mjgcgYHB5fAAva
ES+9CWM6yk6zlGOph22KIKLr5/1MeFQooJme/xtpUHhsBZG5pAWi0aJJRDN7mkEinRYgCT3TBB9B
r28XyUOrT7xLtVwaaGqdEbQfbCqsIdFFXLtiALV5CL9pzwY1YYBcoAvLNtYy0HxGbdv0rLIvo7RM
owfDkI0wTV5AZxRLHwO2T8+GbawSlxZwensiQyugLfJgiAVdcdO6W/LebisLhVDwCrWsI+xxYQPi
cIz/0VEZBSgGQ5pEusMo6Z+SVGTv9cJmf/gbpQUZQNj8V4J4CSye5hU5c7Lw/TUzrSsfUffhQ7F3
8ITIuH+Rw60lIIriJvJTfojONpLN2ZzMlQ6XG6BvI6mdKtP/zN649YTx/zjNomjxlgb3wsKnClmt
4QFR1HVVvQM1d/k5BrL6gHTzfo9wE78ibncAgX/pcSeEQECUqEj3KkgTiJPJaahFcVE+b+CXvjyv
vJly3WHmqR3E8m/qoV7WsV0iRAqALYBGDd10ZpXo9MP1P2o6aIzKk8Ko0cjHMIA6hmbrMn4OwOTg
+t4zcrkhHbnA+5fV2Z24bNDqzG4aH2kAMQVbCaMy5oRCIk0ePX4Z6VTCj6ZrjKtfUSYL4AqAdB+V
smX83OFW0Ika1K4zmiROMKg/70cRH3yEBhLS1UDNJCkWs3o5wF13YDU2ooXFNLZ/iY0eChCOegeR
5xkOg1kksOa9Ou5XctIKKl9YX775TPnfc2H4+K+21PpEyPT1aP7QGacptTv1ZsQHSDM2l8scXkol
UOqIbaysmvbjfLANZyV2CSp5275KbB04W9dffHiqr9TXv4/mM+PEFViyTTPY/sWsyCYzGmN/yTOZ
d666ktJtM/vfLq5AN5mmF19kEVILUGshcItyqYyHBHSXyCxJRC6z6VZOovuDGC00IQJL5Uj2v+DK
2E3xAoGqhQ1ei8YGSmrAnUDaZ1A4gTAoqfZztmE8RqQYol1xs4+vloHurAlNyW1pmkVN36NXVV8H
Jp2C3ffuWY51MFUcMEW0XsNhWKUtZ1sPGr/eHGyJbUgcoA3n7zMv1jLrib2uIvOWnT8c66xBvhcx
QQ6zF0VntKXwwk9ZgEOYVifmqJVa3Psr4oyaNH6CMB+wCy2jK1qQPhsbpFrW1kPI7pn0k+1Ti9PU
LQY8gqv7GdyW/wbvv5B+axQ12umwzIhg/PblnPCEt1+Azp9/yWKXZ9/eDEzeqRPC739ekd3UytP6
K5Cpz/BGnI7jQa/Vft14QDGXW9SnR7fk8qC1W6fDU/02aL6k+lNgWsbBnTIrVdc8et2nC0xuRatZ
CafbDHhhmNdHApxd8aFifzow2Wd0mxLjMOVLAR0M7YPKSc8iy7yV5UsvYaw9oEsqYRb8oQoMSjmd
a4EeahUYOvIpwduZVhdN2fvp7vYV0uQOSHAUicNQlQXivPcJrAU3xPsmTbbCXSmzi9mS/m/s5e9b
ZrHUO0V4WiYp/PMiZZJ0PuxuO/fmQwgyFT+bN2sVQP+/kQteQC7G/w+fNpfmzg+Kp1/smYCTlsrX
HSwinUYgdebuiowztZY3f1DToQO1+NQJoB2UKgBwMXKm18Peilkxnzegw1CfK7s+PVGqiKATfGTF
eq0lEQFAzHbH6TWjyXCadUEkPGthxuVxVPMAb94DggMxJRecmJwiil1pynrJCRpEy8GNZaYEWFTk
+t8wX9PcW1rxVr/UW8ow3HcVWHM7+xzRsK4RXSrv9RsEsY8muAVcD9Tx15wHvsOs8SS4i0U8uk3n
YBA6kR6CtIzvnS5xCsxhSsRUceSzW6QP3ptXRKVi5bwmITOVWt0QhAsyLvlVYFOtFkG8ohcpUPux
4+j8NxQ7i62j7RMsh2Lg3fZoFq9ZbrMOSXe62UanDZjxUsfroK0BluyKatK80G+EtNTfXoi3H4vi
adQIijujyEOaYSmFy2K+zz4F/QmZ7mi2coQndJwlrh6RQBU1t9kMxz4jHIHoN2MfrLPjWgWiIllu
ZohLOTYYJ2FZ4giwazpTIpK1u4PpKFA0j8hGEohdDqO7ANuW1VsJoXKctOB4bunfGItPLvo3oYD+
ARyV9TsTn5hnjzG1YYp21ZzkOzySFhW0e82JO71u14WoDbdgQsxWTH9G7G4UPWtkMaxJsZJM9ZAt
urwhNjNrZXALSnqOxIXmN4VlLkiG0uz/Mxu1/26VsSQNiDtaF0lVg5C1ozhhS70RKw9T/GiB4FQU
BimlkN0KPNyMOP4TVbJLy5mkclSDMF02Lo9mUscYXz3/ZlFlHQ+q+6aClYLMfeXs/LhU4jmRlMJS
uNf0hBs0z1sKO6Zbdw1+UCSc4ko4T0HxT8L1tOa7vK154HPylFGcL5vwcjXV+/Pqc1Z7fzOa6SYU
IEi5keSHCvoLOutEVBvIUwXohFipV/qXlr03P1S8MZdFAzJT9MQlRWV/tK4EwE2NfBpZSDkORDQF
045u3r4lHXSSql0e464FTZvAwC+r27Aqd/SJT23qKX/3Q4+FeJVwjf+cZwRxDWOizBqN2htCfMvz
IKATsWUAGR2yjn+RXu/Y40cv1sURHGSRPES6SBTcMcR3C6JdZL2iLSEUVRvkvVLq3ILc+0yqTd5t
7goU/S+xIK5/dKCygY5p2w5tim49p0nLrs2cu1XMA+CQvHlLO36tG+/XXyJrx4u05zxz08sNWFO7
pGmCGt3Dp26kWivIjqKIYDLOs4Clq62/HtX8UGzNyct8MulAyiZxBhNr7yuFe/6oyF6IIeQQlHH1
slFyzkUEaQXQqPo/swjbTjG7F/0lZpfFz4VDreoOtd7VQnktWakuTZqizCM20LV88WyI4+1ncCUt
cKB4FLDGVqxWrvwqiCWnl+HYf/KzljjytjwdObXRO6MMPROEF+FnduCZI982hOOnglmJtLgg4nyU
E9Cfuj444ETOL1K4eGLB9ayAN8lcpfaKtJtYLgJXKDrmXX+5hr6/p1ALM8bK+Ug3kTonEOYanHIn
5eJrQbaCr8EFl0wMqRSH/jMA1Cqfqqv/QRERp4NStJAjY/VCqlQIWvuzMQGEJ6qbNs251nAHOHwS
Ca26/IHoNgpa6cj7w6T7it8gd2JLy5U0oxWqPPNkpiNabrJyiFOFy6XMaOiCJ55pECh4LVbkTszf
9hOtEVy/mFRKxQ/zKZG6ATCY7CCmtE/3REEdqc2qQlnJIFZBIiKiXAngnw0gjbRnAWv8AuHZTVGm
nsMFmUvOubpO/6yr9zHqhH6aZroHv+wWt93UIZuYhUrFP4BDipB+rU+tfrVAjdaLEcIv1ee7Zvuu
ywj+8ef5JFdyiDHkZACUeOQ/FdqwjT6ZiC0d9PoMKqGuFgTys0C/7AShq0nzZp2haBvHmmGwmJ9T
ZuGTkzQ0s3b7NPoeZeLAxz2LK2mmtcl7QlcelBi0jU7zjIOdNnSlAEp6yRw+4mRyts1ZAwCjNWeP
cQ8FtXBb1FfoeHzwgbJo13v3evbSAhgw6trrg0ATH2tEWITzyMuVyvbrVL56/yTbeJXME7icXzDI
jo4mHp8nRPI+xakrt+Dy+3KeOmXJMxku1AYgd0OVdxqFRpL/ZvqwbRdq8+XIxRDmf+Qb4YMRGoq6
zevEhDLGnL6XzMj0qG6afhKPcC17MVStbZMCy4gHqiHUwGXD9mghr7IUmpqY9vAs6skuf5fJKQA7
ip3tsG6pR1j68AGj0sIWp1WCY2Xh+DV5/vIVt1CArJuV+rByvxIQlJlnD0VvmPMPlc2v4L7EjYu5
Jx3cEfUayfHsL1sNcX0sHMFwaxLM8ZvLBfUlofP1iozCrIwjHo/XZXagbuQ3Inl/0gyWqhq6fO0i
DjLKOs6vM/rw7xo9uqCc7uTYeli4ue4F2bHPWZSE8S71veliRt2Bwl3MiOEEiDZ03LBpzLnVHcr+
duRon3N/+ur2H3Ot05oQymUEYav7LR+YQIQ7dnUFn1Q5X4OWB6vsmjHitEvU0aDlgwtR9GTNTQ3T
lmPMx3XjK/LhUyrJWjDkUqcC1ObFbiaQDZtj6SbsTfv0875NbuSc/ebSxaA1d6q4DO/1YVIqVtvu
nffSEUnf4XRhcOtDgTe+HB028/sq8iFUthRGzsZAm9aHRCG3LHRodZCFHXhPNs6mwEm3VWxY2bwZ
LERqM/yze3OHBIcVFxEfNgz+ekJzC+AG6sa3U0JqQ1vBjr9jR3KwHARrY5Hv/OlpmxWE+y970s9H
KWBiU2VacFC+0lJp9n35ikEYYKc4ihGzRyww7JgZpXqxx+wB2lA4q6kKEq0cz+AbKu46HhV8BQfN
N1z5mkb4hFxvWEzz7FiKKuwIvv+j8bosGI5VUqMyTb3VaH96yamqGKwCYAC4nofdWazqVgGf6ICV
9wfudnx4HueS0ra9qkIUE9FuqHfpnva4tVK6d6PUxcR/S7K9Z4R+WZU0phxTvdbSILN3d5SikppF
qC9RyYK7hOlF4oA1VM2xRCHYDZHP3urES4VUSFUGWQuyehxg0I8HdVhpu1aeBlEZj+IVd/Z9CkXb
YZijgefuL6pTRdD9msPtvZg7H6whv8AbOJPcu5B4V4/G363og6sDh3NHCneJEWM+UWdBOpYCwnYU
apeMsWggS2qJC2FRCmx1laM2YmXeSh56T+wtxLHgR4ej1UtFYG2tebXuFkHGe88AR4MKhK66KBIx
VFk3len2IcwiOrkjIt546BBIZg6nCPICBNkL8FIXfsthpnFZXx5YMDNfUkfNxnY6KH+Xz+Mlfq3T
5RVpYXX0+jr6yRPx+No+d3668UfS/ZobuvMow59K48TnCaz8Ge9AteeDBQ8LjvcuJwK/wbmb5f6U
9Ybx6wSIbqMMkH5HdAA+2PZDffwPHyMOHmpzaFMdpuQNTJzZA49y0+pkxepEPWw0l+UqMZq2pJDe
I9sigqcG/hHR/Ep1j6IZuw4KoyWY4cp9jZRCs0JKs6m8wsZANDI3a466bKvr0tiISAVbFU2dCDSu
UKvRmU6dVsv2wFes1ts666cFk3ypeV4+Oq18WgvjJzROsEFsHxOkU0B1s3x8h3L2mn3zhQcVrZg2
UIMwsXq5MsASLNeU43gr8y+PQ7RQtDhSNj/31FH/lvZM/3FOWQBknlVxvmk9dYYCwMVubiKZUiLs
q7f6sNOYPOq+MuWNwGQYuEBpu6KhgDB25awNSoq7vvavs/7ndmZ/wkAluJSbbL/gRx2RSrC2bM8u
h2L1MwF8yfQcvcxDbNOnmBhZ22A074pUDb8ufJvx/6sX3AJRRZP11TIUDucjP2NbxdwrKrLk0cj9
eN9Qv/PuiBdfvn7JPQfFsz7xaaLVtcfmJaUMSN5T6tVwOQIwEbMulBNbYQTUsrx1jaC7A5dCMvkX
rIDYsrtsET/qMbZFKF1hNIEDdd1ZiGYSsgWFgKg2B47SV6/CB95DEC9Ox6cnbt/5arJOwz0ODOt5
fNn0tXTNQG1E7MemTdp/i1jZjsq8WcOUe1TGDbKtsgEpMAFf4ltVY1Rb0d0Rat8kuh0VFQGdaVJn
hqjq+FQ/LJUB/5GCA2sgeZTVWXB7QOLwiV4YD2QQ04wtl0n0k5oUD5HnRpgJt7xFxSJFyNVswA/T
H8UH7+5JrrG4BR5V3Z+Zx/HD5Tkxw/fRXhySQ4OxPLvLJ4WpSz/rIOUrG24xzEIR89GzNM3zTb8e
RYmxiB0gYcwSNbsvgF39UE+C1Qnlq6OvidyuX7JGpWLaARMYbaFJe2UARyIShXwOY7PUjN/bc1B5
/vqOrBwInGiDggNR/8b2Dhno/K09d8R4Ba9R1RCWa3WnVVblf3NSsO4a0Ty7W4BJ6FlOMT+ietkz
1V8+TcPht4cblXvpKlQItk/sYko3Cx/RmixhdUR4fTkrPrTqU9VUpPrGtn76Sc/q/oVAwcDZR6J/
OOLoMNxwXAB5B02PgYCnQKffaPiRBWc4DRzBPVwGmBXku1kCZ4oaH21z/roupYpbg98+KJiDmJH6
t3q5cHhULGqouXZ5/xFv1ewip5+jg5ikz9O5r8cCwukT1Z9a3fPITY3wDxCfyqAccm7W9Te+Opty
CH5xGhjJyNrbpIRpyz9MVl/aXv8N5hw+w26r20lzKvoif01qspIqUsDWPFcBFCY/005EKtQLmx6g
vC66+++MGUKMHLd9kY0zDjmekOtWa6wjGLnljU3YjU6FtCUoFirh14fn28h86P39jWxvRK7xE0J6
mEVjHc64yBpuUtrXiZa8Xj8q3TpG5JU5X4DttEcsQ8lhHRVwxaw1p9XSuP9Mefokm1hbyaUP/Pbm
aAgITd2eXbVYzcNwLKQDuMcaLB8njxWB4MklGs8pW9eR0V07PirDEq1JInTEUIz8mmHCWZ0sCOS1
LGCarQuBP14JEHPsm5lX3MMkvy0q899Uoll0CZyyOFEd3QaEks/LMmRAUOH1QUKRE2A7L3TE+OF1
IN4S2UrA2aq61cPRhpMYiB5fYwGCJkxXig45cGgrxOs9Ht9WxVAsT8twVUqZN3ZQ9VdT/xp8pnkV
WPzfZTWXShZ8keUyEqelRXLZJ0Wp0sc4JIEhVIsqLJ7fEo/RN4/S3516eg4Phbbxll2JJErRYNs2
87zHu8mWqaOA3DuXmGCD+95HnfFRrxIOLAEEy7wDrQcrxbnVatGtA1nJlazVspPvwxT9LsJFE+Lf
R9uOxtyxYa0G2XZiVZBJRQD9g2VRW21ieq/qbWeHTYANzSJ6wGMKcjFoN/ohQIFixoG53GtI2vhL
LjxCWWfY9xcY3ceo2zgCpom7EBZl7vlHKUBQhUaUdeIawjOKiqk9s79P97iT3ysr1+eC1/E95zhS
z5cwh9Roay2JXNzUHWGfTlg6A2xbY4KB4awTq2qaCE6XKXy4lfsOlVOvLvFMZ8cQDU77qNINxrJy
NHhvUoOY0M9gK2WtGJPvBdnH6kJC4V39d2NeE7qo3UlIa1NcBSiqfMFY0los+LRs59yWdF9gWrQc
bPpjurqyfBSx3cKhPXOfMHf93hKoPLlIgSmSouCT+e5XyQ5ByzORBHDbNy6FTqsKEMbEzZ8ouUCe
vryqlERI6huJ5KRsZA8qIXAJrDZTGme7yEueawEXKtDmRVcb/I4feId9L8vpcvKJMeWJ8xQ4hT7c
mtPgXbZxKf57SxE5cEy42N+IdeRd9QHLbLwVQbVsB/JlygLE4t/gVthk++7wyU5uoBVk7T12UtA4
INPqyZra5PEaF9n31+iP6F7bvMpk3JwMq/T4GC7gBsZ8T6usTJERg+Uwpvc/HfWPNZvOh0h6gj5x
wyA0iYX5nihYUnLv1kloABlug3DH72B74+0+/TUzsHMY1v12gc0ShH1em8/yAxk64zx7IfmzP2sN
ObSD9MMz5tpm+CHF7j++M5D42TRXwGOZ75NAS2EonbG2uhFoMVLD+7WwxFE84BiJEGND3pesZgs6
02JvgF+PBmUlTNdw1Y0kfITq3imzG/5MowOx8O7I3c7zk5IUWbHZGlUKmAXqMIlrS65VyJXqKyw9
AcGZ5t8WH62GHuPY+AO4TjrsXpe5RTWYMycxKEQoU7SrDYsAj1v9FeOs2SRKBND06oZh/nuCvhGM
uu2V0gFfzJlF6J38yz3n/uaiBJ3i9renfSQZln3uDZ7pV1FPvSpG9yTzaRU1/BirE3soodTCbJ+F
eVkMuvP7jsvxPJxe9dFPBAOFF1IrwZMghfTwQfwe+85Tvh8Kmi8MyE1Mb4aLhYAzj/xZUyfhu1nL
Ha0bfcWLAadmzUekk4DC6cR3racZrfwij0o9daLDbA9fR2fN8ae55x5/F0nmCr32Ls1hW0e2H96Y
oYs/YHZdg861qp2hxMvjKBCIpRQLlpcKKrmvj7brOrUAgDr6EY0C3dqW73BxspWc9FZAqO5dlumu
j76UwIABxiAADEm4+Hp8204UogPWFbvUglcI8sMKSZc+FUyrnIxKE8HpnddZ/thYL/hYjJgktCRL
1VZlaEkBE1J1/f4tUKZz7tKcuFOXlXZ0TEYuu67q12YF9rbyCl7xtt4ymSBhgEQyljjhodWkEW6G
GSa01/YGNArqJSVTXU1sf1BbW0FtYffsNBzzFyhpnVBJAQ39DigR/zfID11LvEudhoplRCrqs/iw
tp9r+PV17l87ifLqixDtN8uNz1EiC+GLhJIoJYeFh0/6NkMdYJ7zpgdO3C9r0BERTNtKxe4WUmmX
YBVqt1/c4f5oqo+Iqc1enk0fuTBFfBjcuqtogf8d8ShfHai6/SCprisGJwjKJzgQBMl7Zq9iFABH
Hs9/IibZY7dF71AsxaqtwluTQWGvIaOYlTnaf8PnSoGr6AEHu2qU3+epEFJzEXMBo4U91BptyKKa
klZ/N65Zz/aUYaPWc+O2eL3QhvyjX1QitpcEit8QmOfDp0dtzSTNS0e/ptlfZLzF0zvX2ECcvcK5
VTJihSicv2YryXCAhBhrX6dYEqaY5OH9pChnl57Xu2ofKt4HJHh8/INc5xJAa6TDobXhXw24A6pA
KtGEql8jRGbXi9EHY2BMRcE7+wnipQi6ACtoHM1x4RuVmC9nNRIoWB0Ulan59X3eQju6HH5kQR10
892rcSegn79btZ+oQxdwvMwrXHUbWqN7+PiHO5NRaAbWgpGAXu18CiPFkB9SFqBQEhMQ66CJxHdd
NXnZ6VE3oU20LqoQ9SWEVBAzJsQ707zGayrvdm22M60shObvIe6S0E8kGBltj+fTwmhPOdYIkpuF
FU3/1c9ODTBGYge6KCdYFrK2le1dqyefaZqvQdXxPUOgwV1jz0ki8fdM22jO5qyMpAUwS7gDKiN7
Rds/SHLgrdDSnkD0cB7cp14EOOo2lH0r4MnTfkB3+Mnel/E6STtN8/CNmjuBh+V7oRQQJ5tXaeGv
i00TaL6moNkNJWNoC22IctEoWvsAfarqMgh89Ode2IPTIEEKctjzRQG0knm9W8eCv0iaZkKJrH+D
ZzgvqqgJwMCw+kcXze3yIKHXr06q5C9KjTaXmBEGieiw1osnX9SY03K/ZhMZYMqqHFOHKQ0kJ9qX
BIac+9OXLaWMEuwagEYK6fq489SQC8rFfMRzAMUlQ5JZFhnbkKI7Xp2hQaK0mai+VXoK8JoXa5CJ
x0k9LsCv4bA3wbH8a6EXyO0fmhQEu8afFTnfobKc3U8kSU9UrNJhkKEw/wCdBPns+2J+1Jk8MP0g
XsNacCX95QaDbfj9YS6L3bpo+V7p11ZY8urmDYp/fW0ipHCsxotJ9AQ+k6db2WLJJNp+DxBmK4kY
VZZRYMUyM+sXkaJyXhEHrTypaRinqd87Dyd8xezHwaDPbBpwab6peRTaA8hXnwz+0fZAobck5DBc
rIRF6tbVMmmhZ6KaRCfRB69/JHbEqNp4JW/K4jXkgghJ1DL+QooroqGTi2JG6wdiSbXJLfqgmNAp
wsYjkSuJLrsJP2YZ6N21Y2xOkxGVvhmJpuAWRht+FRWwvtULH4YxFIrzT8t61iVzukJmlx4HuvYK
QYI43b5CdeGp4c5X90AeQtXx20FVe005Nmow+xNxNSvAUtZxXrtJV3qS1nvZiY+Xs583z6hFiv0u
Il2PNRhHvz57oYzgHC2XW/+WDIprdTfu+epyXi1E8oORPXJHEuxyBPe4pERxpxT7pzARNCZRnpa9
db45GHSF2AcsvjOipHDv4t5P5i+Fevk0SbV1JZ/VXVBBJrziU+251/pqz9JDKIt9m8/x2glDLXVx
m5peHkqEtAYsJ/qxeH6UBolCKIySlkZylNel6wsQEX/E9j6UYYH0bN08QhQjM1QdHJ2fATF5ajFj
ej/QgwizeCufSKevCieKf6QfgZyHtQAn5cesyBuLmmxuENHF9UhchpvKpJBbm60MvB3InQ2rps5m
qtGequUc/zGT+LrAG5/FhgABdg5yUTwXjAhwDcYtTr2jZLcyKyTFKINRWvP09jVmw+Erb/8hCKQ6
P2wQaCsyUl+D1H5egOH0c3mrbEZ/1UWPKbTz+AFbzGllE9D4NK2uBweCmkE1f42iScSZriLlBKdd
T9N6UXuNA7BpSxWPUluKk2rBf5SG/DqtzIGE/CMnjHWqcMqfJ129JpJBm5eRaMaAM0dZ966GtnxX
SpPQGAga7bEoYVDH3Gi5lETbSeChQNaNeiVyIpEkf1ur5Kt0xEUdsGi5ccLyIqZvuHDFut5NLF0g
j6rNq/UgC+PwPc74zh8V7OM9b8hglW7C7A68/YCPBeJ215XtHNoveGIjPWLoCV+1PC4IBXW4YMZx
O0apLzPPSS609YkSHCeoANXwkU9DDsPfOzNC13/oKVbh40viBjUR+X/k7Thobvbs92b4IcoRYyGL
CbCCzoGbnSFkBMikKUxRDGw0AUgX/aWFbTU03blaTHJ50m+2DsDb308LirygXjo221pf8sW6wEc9
yFtqcXZ4TttJCHhFb2kbBhf3RoXYRYLDokVqWOlIPUG259oeHzp1n/bDeAgKOyQYuqmYsM2mnXx8
JaX3rRNQQ4Np0uCCA7NpHPlihOQweKKIi3qbecPExCQcdjXBe2IbaTaufUVYngMvI0P3i+FBtFQ4
DTkmdB7QPtX4RJBJLumO5LVC9wwxxclLuyLtVCuS5I88b8I9LQHmacr5PptUeFaJT9qbdHqcRlcU
zJVnsYjT4O8mec0OWypRAB18uplsD5dJ+jJPdxyxteVhdwVTGx6zpTCX2+ZLZ3KW6p07dHyo1wr7
k4QUTsHYt+gifrDR1fiYRRZQenCvnk2ZqlcjGbjtax6qNO7gaqRgKI5WT9+S8KRLCzELHAnK08Zm
5KsSn/4tCf6DG/LgocAtx4mtMAnbJTIG2MKqco3+Tj5OcKGuOjLhb78iNRZlXAalJwzGQG+Uqgzh
VLGt40NZYjAZDwc9kKAw51PrHpyfTYCTqs9iRpfRdfcO+DuC6xUNppw7RaT7zV/g/PVOVEmmZM4P
ri6MOKv6i8SPSdILiNg9twgizAbHaPkjlXzRbDI7iHGKL2/+Z+3Ha60TjKSNBEV1rmkquSOunCq2
5hmJfH/zMwr8fb1XX6ajUgdjm6uAhyjNVeJ7YMznQvTz/fd9ZYz1/mGLubM3nA2kBBnlCofU/T68
JLopbDz77pK3oV+wu9CoC1xe8UQQ8l1ZlEsfjOhn/TGIofhvFCLs9es3ZZJ7T0CQbPWSiUWnNSmN
cnzpJA+KfCTjPqE/2AQTO3bOCH1Gs5N3+QiIJWmQdG1aeUXUwmawHBhRlp/SDeqX9QIOtheW/oPo
e4YJpAS8YOihGpIwCJqvIjkMh50wdeRAZmZO6BLZRCzfe5hku/GzP/YjfhvtYFv/bkvIxOII+9Tx
eF1AYsp2Kgx4uSstIjA/9w4WbbUXFhEHog2z+KZIt8S/0ddUihAdF6a1blWM4zpF18jwdQ8CURv7
NLJar1Ub7Rbho31drH3kYxEQ855qRXWq2OolJeRBWYrpYBEXh66ZYreCC7CgGDeN0587/NVn8lqE
WhDlm/+Pe8OkDDX9EanTkTvi9y3owrpNHJ5UNQacAEQT79qDsi4NEF8uVC1Vw0gNjPSRWE6BWP9f
uX16lYvw2kggOYaTj+6cOZsLpEpQT7S45/BqZiFozUP8Xe/RRESgk9LgMlW/0c9ilGfA2/VUi/ip
OBF6yhb0tHkWSIelKu+2ADexAqv5LUEftYkCKgT1lEo23hwiaUMqQM78tm0wUIq4XpDWcYEDkyLT
8G4XZgDMeQ9EUlr8ylq/n2wcZLJhHtkmPt4yVacpy15EU/fWH8tRg5e8MGUO5ZFZXECdnFjyJsFc
6J20Dse8wgJRUZqpQKX+AAQy3YUVyvzxlByGA3uqCgijyxPLtSjDSYv9cs9DF0gJRgh5kDxuAAEc
0180yhgzQKqAEDJ4tDYUEAs8DBQF6rFa7+7k8iJV2xbcxwYZUuTKJUgSDI59IETZiYV+Rq69eEmK
d2PcBJMiyv2ip5BGGqu3y1BqlrWJmcfBfySdbo3aPANAd6mgvAUlekftfPOon203ifuw9WmRBQU4
nwtwbIkwrj2Yve1hUiA+uJSlQ195ev7Sb5Qhci1+dffNW8ZWdCeqXFn+QYODiKvuH6adHtQfcASe
MbR5ZyXg2CAaKCwILzHtBzeUKZNLQ1/3sKUIsiWunIEOI5JwsSt7SiWS4VfENmQWZkigvqJVofuS
sB9dfUGwYmrh1Fh5xiDNQZ+x3fA2nSxxQhFebR99Cz0zqRZgdhlNqcJ/bqT6Rr0lq3pkIPS9LR0i
Dc09Juxahl/U/LHeeZZ9Q+aosrqUmEznry3q234cKLOKTNBbRo5zb8mHwm4HBxF0Q+wBg2IEFjTn
6F7LNlgw3gbihEjs6fK9vORm8WV2233+s6KOiJDo93e1KpJaSe1HMBw8D3zjJRqoBU3PxH798rDC
nRRUAhyWg3I/E6d950IungDedAD8voyp7qkRwJJ/9MED6yAZrKa3qCMg2+U+RHQyP+kmAdWPkMFO
nb0loXSeGtwcdR9zJg9yVjciRVQQr0xXK+N6qZT3LEGrzmrU1n9CcYS4Bq0UxHhpiSVll6hsSK43
B666brjAJ6ukavEAPct65Bn2xKpaSoc9+Wd6yB5sEIwK+rwMzaxaaruK0h52/mnlvINuap6pfdkJ
KfvDLo267PtOz4u/1jkS2kGeo60V1+pPM9FWzW5Zfhlh+rngabKhzzFssHNe6pZYXylpZFG2bKvt
nrXyo95TDLfhMY9OKuQfAsTzQxEw3e3beam9tnZhltQw7Cl6rkeZlnGJcmsWObx+3KPKoO9hX343
oEvrF5C6WDSQ6t8nYQuT78Zm58njX0fgHx7SRSetNbkP1g+VOf7lxx/1X1jNEVXhUBPwl9vjn54V
w4Q0RiLV8rBhi3dCT3CcB1vnNbAArjZ+hwrKCuDWxL0VanWSLguKtzNRRWPJvkbbmoz8sRG9D2v9
EhqinfkLjdGRndmG7mIOCqF6o8dF7P1HJjuPQTNrfKBf1DI1B390OgVWYW+kd/V2HYDjTg5+H66b
oRjl69Frl5Ai22nFriSLxsSTUmKCrOQbEmPDp8z1jY5yPz8wceyXIy70rO4jwWk4zL7y8KiXokUL
aPSCVPbyYbryLrtqYKHOAcHqf7c+smdaUgrHHoRhKiI9r2gDtZUzDMtABKmD/dIpLwVXRlDtnthA
PeXteW3FEnLTqvTdZv/z/hdVjYJVlzl77FLUEjI96gxeYZGFO5H1HZcCKV9OE/nBHNa3M+Gbsx38
mckb8t0xPfT5lqzK3mUh5FXP2xFKGXLS5ASVS414wFG/uzjPEUBrUdKE4n//2kl+bBJwokqapXFB
YZ+LKEutQKPt7XHeaH2kWNtC0NE+wgDqUxIDmPW21uNu/f00bGXV3e6FXVIoi4g+Te63o8m36QGy
zbgEQNxwePqDaSo5tr9TRI02hBkZYNBexCA/m7eVDPqaYM5kWXkNceWORW3xDl6Pj9pGMfI/5uRk
fmS9DAM/bXuCpKTb54EY4utGetwJlmm4HjN4QY0ixAkp6k90TEgpU0XEtxhFZloq+T1d3JB8oIaE
0RuKmEUMT5OzqBIWlzazTLC269L2ha1V6csdaaYFPA4gD6wgvH0/9ulq37q6JWb+bdGr1ovwnMjW
4smR7h9AvQsg++XvmVpNmuQYgiR6Dnq9Pj911TuqJjUawkCYj4leItnnZ+/o83Wtph8pQqO9fctE
HBLA1GiyoBZi7dOPg/VZWMBdTpDRY6p6foeHlTLOaKUdA3oxGXR2rCZCjpikJny0PSGvVs0yIMpu
QKa7vH47UI8621MugYTwkFmRJY5QK77GME5STnO6UglvNS9cWKh2EH6vjR/0bhzkS/Do3rxC4KeT
pgQ1ukezXNdQ70T3HE0ohvfFEMw4Uo1MGNhcnM33YpJJdAs39JGiq03fbZcIdSu+T0X/hhAVZRBn
6N5cyRjo6GYkgkOSx3EjuDsLVOXGveURss8psBDz5z6I2Wl7k3ZVVXNDo/2U7ceZLcYdcaysvuDd
ZZnDIzNVZRrFhK/sAJp3xgRzVb9TSZmlTAeSsCScYGcwZ0fMjldU/pF3HwFLUebtyi5euWV8f5VJ
xK9c/EK+L51xcAl+j/Tz4UwqzD3xGyym5CgyupByTF7Gz+1rK7TeMKC5I5krK175H9vHSt6HRgjf
2oYXvr7UP/SQdAY+WFW0vbibRoauLHl6EOnhGBSEk1OZZjZlVb6CAFVveUiNcjuLdZEEj5CGzBO1
gYfxd7T6ezoz8AvDcSJLB9pfeS/ToScHUiNfhindoNoTa6kd+wj7iDI7oCcnjbCZ8m6jxYbuLYrf
KDy8XJCygj4Q6IMfXlZy5n/T1OA/eroWHENmNemaT89SEcQabYEU+/9bbl62/UYj+lT9wWxoKEXy
6NzA5YTELN5QBKwtxql2rAFU8wiPJZl2jDTLNExoem8Ary0BMEhQsQn55d61wZeB1l9wvdj+EGV+
SL9G4r9LKSTPj6qg3qeENZwT1SfeyqcuPlLHJUIaPzt3ZEcUjO5c/n4Wru1X6Kj/ZyJXqvuz6Po5
gy6w7hc2vfIldAYOCDPU8hSKrvwqK9W8APU5i3hnsWzvoLHCUWWnO1kEhHodQb0UPfoLMLf7qZnP
bDSl89dnDjJ1vZgmP/Hc1Cg113P8ZhFTwC/YJ5gxPVHxcC9OLr+zj0tbdJJj6lkjwyZnTBMxH12g
Gfpx9swUri3SCGXSUZDfZo6mh6h8FYKclsZ6yKGLJWdipEynbFH2da56YcL1Gt/yyeUsJu+H3DuB
FG7WN7Ll/5x8O/OBhmh7Ivgd69U4VTg0u0cD6qQyFtfoKzVzW5StnuJmfI4mHC0oOsoVV4odcyx0
HVemDIb0fMyzN6tutjylTlX03XDyb537P9pN0mXdWH250kiwe1Nk84DCaoud9/YXaDE2Bw/I/u6Q
oMr8cplbOGQmYtJYM2v226dZ0g9QOYJMTU67SH9wPGKerawAN+ldQaTmThRzjrcsriBKHRvD6NbY
VCEkifH7821kc792V7vmUajBuBser5bqngAEdvtXYLholPQ4R1j0dGyOMXgdeXXsElLbJZew0HIM
O4ikQVj+DxpsjpmBsLRclcfMylxjkZP+0grJG8Y0Q351uP/sK/HNhKOz98mhdbD9PIVDY71vO5C3
7p9Yd0xdqdXZKsbR2cPyw/I0k9CtvUSLNFuy3EaOfKonQTAX6/9G+YwUIsc22EV8Adu0X16FTAcI
u5TKMVd0WTbJ+qNwbm6B1foPuNpnh3ivAnxgwyNkxyECzKZiJuXOcI7FGKtgGHjPT9iJgFY40bmR
gc9ne34BF9GlWpXxGeu9LQvb3GQ4rSLSliqJril4xfbdqWXtGV2axcBM1Mk8QXBhAfkRY1kg30Zj
kbkEq1r8OTmOysy+eA8D8zVPGirK3WIvMN21a+uRWsVUdZWOAfBj8N5xHQyrMyzBv6Y+XAHJqt/h
vudNxglZY/1zDUZWWbNnU0LcPxFLHw2I/oWGwKgGMymkqdfs6wPb7Ojra/hsPUoXtpkjfBdnktnY
ryZVLvqPeZO9CgnFqB1kPS5ry7TTOHqJbjUzVPszjXT6MQR399eSWIbcnev0CAOnvvKLJ7xwxGv1
ERF5Ejo/0J1fdRDlWBLeOYi2hwQp1MrhouDfV6k8oPHEVBy4rx9+WsKIW1azPlrXEMmXf5VQb3sr
FZcnIRzDlSmwqJsP/iArgrAbyeQt14SUf6eZswM7rQlKcgELOsoW5Vs6ZCeA152kH/JjUaTW7C17
V32yelI06gW+D/HVyH+rwl35Y7D3rEmuSnXbWiIGSH8Ig8b9A9Tcvf1gjxPXvG9W9WuTe0y+8cuQ
1lAXD/rKwXuPcFWT8/D4+q0DgtXEjXhqeXHU1hKY7+5vD9poqsHAHJxUP0A5KngRju610C5EVi2B
R59Hi3bSbtNOLCLIw2Fd+8p3dGvMrXZQXsRUlHEPrlAHdqUJUASbUBvmpjSPVMzzsy16n4l684Wn
Hv4t9T/ElRucumRcAFEAa4yKP6sPCYmrfOs4hmh32CttASZyP/KJqyrHNqBPyuBy2BFF5kmpvzLi
EThvejatmZvykyqf8iCsA3e08N7yZH6+a4k9TMfqSexjsclEUOGdqfcTp+ivV/5uKK9XyrNl1JHc
2y2/oE6YtyxkN7SRyF4iZV2mpRTA5bjKxg9vV405rijFWwWGmt9JINDErk7bIYYzp/yYsv4R7QHj
Kpwlb9VfRmfUMtuuaFvMcnjFp8pudt64ISkbQ0G0cm2ZxrbZrMzkPVxoYbE1rZSnon/cJ2AoCZk8
bI3ZElEvIQmRXTlh9po8J82T0TShPRtDW4emnwrV7i5ud0BE/qb+PM/7Go1QUMcl0rHM9jZwUSr0
TQVBrGHiGJTITnyIblhTGpqAkObsQtItyY8StKnDhB1volTOIjYP0VYIXL9KiEIz/Ytm8F25/w7d
JwLU/mHS10KBGgj8Ap2tmGnoKrwjyFyh9QfKQBT8Ub91hBCnn3G0TF6YtKktChljwJJY2lpB1fKc
3ABDu+AtDPc1eYRZvs7sRuhNyGC/QsDn8vBb+qPGbJttfae51NBa5A5mULP78eZflMqT8mAlX8MZ
7nBM5YCygSF4f9L8DA3eQARmWavpRpqbCWgYezMsQzJDPhtCCxG0601UTMa+quuQifTlaagEwgE8
W6AFE5SVxKWMZo4mKlEH5WLf6u+zj/S4Zy/hnorMY4Je354zATQUfHayoTbHOjeWsqH3xSLC0CF8
LskktlJ540r/czLtlpZVin3S/BqT/XHC+Zz9SqQ19mlOvbrzIQiqZZeXj14VFGfQMBiWMkDUYD9L
QgzgGslGBHNSenY2kzGr3rPnDr2vRHKk0kJo/bAV1RZ5CN12deoMm09fIruUkyxZXyavJCMqPspj
oskhDZFOQkrkByHEXy7+ChoTQTaBScWU5gtcWdP5xggGHmUSvA01y3K2+78KLFibI2PJDO6xAaTQ
oHGK5jfEiO/wFB22oDrVAdfrd1bsIYZevUSB3p+yXm7Mzy57ZoSnkf6BXibYNbhHJl792wyrdVsH
YWPj97DCgM9qWobJTxEohGxIS7GBou23DbpQvHYxzfoI+xi/ledIiKjLymZ9j6HdvqGkeQToHOZA
7gUM0wwJP9x+mxMbKvofhNoyx8MRzO7E+PrGloHbI7f/13mPVQZslkuyeUcj+CixchAWQbjW6cy9
hkQmG2pb/jiXU/KXSkOHOQRSX8MIjQ9YVavWKKBdB7vxX6RIoeSoUweMVOm1bRjWcZMO/By+WBDs
5VLBalEHsOmRLPUr8+yFRR+VQZDzKi9S/I88zZO6DhUU5oBxbw8seS8CILCQt7Gj60nIXDg4zhnB
7dGSYUEsv40Y1FU48Mw4cBrkYN8//yc9SmeiuXPyE9vdZFgUh7wWpzTr2WTKj7uo5KsnLPyRBh++
U725HKjbG1uUNzqgHyaJayA7VwewoStstpXNE/DPf9Miiw2oZe7MBMdamOyMB7qjwq0ahnddW3Rt
sgG+2WzpOB7tTuL48yE+6mQ3SGklzID5Od7dDSH/D1jrdGhOolBJrDIHWnrpL2DYxpUH+7Q2+lW0
ATsOGXLnk98oA+G87SrhVU5rZQ/MGz7qiZcCRKT60DC21xUDJjJy1ylpV/FxtIifwWeN7SgM/ZXq
3HYKfrjF2KneRjqe8P35D/MHkkUe+n3n/uEwNtWiCd/tY2DxwZqrLTKd7mJdY50qujgkkhotx+Bb
FNJkx8npBXEb9Dy93CSFRQQofwaMlgbifSHcLwsuIQ0zC/CE0xx8mfl9dZZJqN7Nb7HRepD2+Wld
BVWDQ17r19T32SL6N9OaecNeKoWifZsPgw9+ePRypMnrTJkH+ZI19rtgDBO6b57BbmUj1WT04WYh
SupS8NpOPd0YZnIPr5vsUsV04xuh7cA4MgFRsFHzukRFoOYljD5LTfzh7bgrE1ICUvXKr/aZByxE
pExC9jXZF6VIWc8RjJjDLgEXwMjVwVidiRFmk4Hkmp0zGr3r4enga2wXIf3C0Xl/FoCCEHMHwhat
+mqj8uX0cABMjOJNKfkx6U321HNqy9q/NntZVQiRswJpmG+L6aECJjNgw6cPAS1tafJeQktLVqSs
OVJTog2ZX6/IGmYMLRbZcoRkhOaJuXqK0nBgMka9dtJ7/EU6Wodr5IiLlV+jQnHRL1ubHMmlj854
woKT153SupZKpnGJmawmi8wXvXuvPa2aJ7oaAzYTUz2hyNNVhWT3a+MT0CO+f7JELX8066WQ8leK
7q1KnW7rzMCSmMoYGT0No5hxxHi3jhkeiZ2XsgTFMe32XoB01579OF8X2yyEHLfbJp+iwLhz8ukH
sAw5KoPD/BV9cEbx8nmlErc5qZWFGC7IefMdtJdjGItdGTEJhk6Mf5WiUMEAnisNYYPI1E4QA0ql
+EwVmjlP+K98yVVFhtdnLLyXfCHdbHnwf6q8OHQu2SY4QlhVI2qASxShsyz1HN3pC2ZbroItB+UI
KXGbxj5b8tFLQUGh26Nes7cwuSAvz7yQTtiHj6JkFjjC1L9drK8AshtWFnegX+EF41BnMTvvCH4C
3oODMvokP7KKsOyefVapE76/1Q72acqpgixMW7G3FCeft3E0li8at2lNjnpPlfjG4OW+j/9AcDri
i9rxbSqBsMD7/4F039BZDFGnL6LhBFWxBlMTlvZYzQ2PuwiYc/JkdJ5WjEgY+yzG0aR/OBdPpP5v
IKvqJ40Lh9+t6KRK2zq2v3w2BG3oDiIdFp+spd4GlUm5N5zfzQSvpgF3qTr5hEIjNBLOSJJ/t0jr
7PzCtW6RIAheLmLxa20uGECY29F3eW/dIhdWrRT4KnVF0l+qYMKuKkeaFBQzA3I2rJSUh06B5S/q
WCQYzKU9MmCpxKOnjE7mvVpv7txxBw/6s7GKmme2AZRl4J7SQFPtyeniFq1EoYz9gE2knpKGz7Gn
ED1zngVDdFsNt6dIEkVivUK/0yKZ0OX9r5jH+/TDnSCz+B3cT4Bt0TphDjJglDn3oRhZWKYhf1Xw
ILQE44CJbYA9esWdidx/17Lkjx8DgLAw6i0wkO59Dz47nezVIrwEc/uHLisicy18CdmaH5C4diWf
4sZ/E3xrRYj6YVM8lD8j4op1J/vbsHjnjFr6N8TFwEUzSP1EGqQoHoNAW2/YWTqCU6LjrM/gWDgX
5xw/MmfWwW7lzTL2wkrWIaDCOJnN2TAPvptXEohaXluVCGmP7uvLbfLcLaR0x0fHqh9emfcSsACW
6F9ygu3s4NedANpYv6JxJ6AskJk7wBRTpYMOELnXvs5ob8yaco18POXSuU0/gK4PnN1kvo+1l4X5
jtwKH4MK1ftyQe2GC238WFvpEXjbqg7plRoKe8CWVhRTEohQbhTQj6h+oxO6qoj0680M/y54blaX
L7NG+b7TwhRlZVL9oKcVrgp/PkDIFS9yiWJysD5XU7XB3F1iYWdQMlYN7UPZTaw/Gf3Ojl3Rr8eO
t/yKrMcYytpcwbKcnI4JwmKC6+y54vxkUoilRbIth7XKa/InREuEPkemna4YDUsedNs6gHW6552R
YcPDM44Q2gDYsTWZnrjG8yjFanDWxX2cwAQhTyY0uyFwRG4NgwakNW6O939ULjAUlRm35aojSBKV
ywLiNSsebJQniW5bEi65u3R0r6aevYsEZuR/gDh3XVpMNzAGMUqXu3BgKswQbYf4cxAaz4VIC6A/
ro2rOXft5IAF5CGP2bxwEa8soccQm3DCdxMQNEIwhpt8H9Cdgur28hGxMMnNV0pxCGO+rtVOImED
LS/pweMDpcmvyNFUxju3t47jce7SM8dxNPd9iJjHJZalUUYeR402w7HFOo3b3tDEgVo4u9xY9NT6
CkvbMw5WZGeNsyNBIVv1y7TJvlP8vterngPEIjCy2v+9u0+ep7UX1FXDRuDJu7kw6k6Zlpb31Sb9
IBn/+jFSr7nFPQ7yW924mDRd0OZJGA/yjLD2DwxcYk2OOgjKiYYoh3yJcWLc8bWIbKOWnzRJIJPY
DAE1XXEV+zeY2a89fTZ0jBoktst3CMPDfPUVv4IYMBIRki41bEGiN3Lt+U7rE6EeEbIiS0nxyFwI
k32wynQL2wPs+Cg3geRWDexN/tVib4qC2cMlbBwyVHPNpL0BR+cSH2n16r9fKtDJgsNBgNysfoAe
OYOcyizcOZkJtzb/jcekblKyQZN4kLt6nQH2P7Cy1E+dP1Nkw8Vo7iUmROueZPOCLjRhHFstuO07
/iFyn10DcxwtI5ZYp0nHnxYu1H70cs9Ehm0zbf5Nu+WHVQaqDplrLw/cSV8lgEz5dGJn3TOD9TjC
yATBw0BcEYiIbWntyNva75BZlX7A0446Vz4N8WPi/YTPgJuG8XhxFy8di06ZpD8vligJ1rD6ElQY
DzO5DeJlFw2yyNIjzQzZKMAnNfKmk0wDjbC8VkvDGWMVRF6oxsacAZh3ECar0zd+1BMXNajE84xA
Jxex6xijnSKWGMqEn4bv1m1zOfX6oxuIM3GcUCz6p7PZao0Xqgi1vJAgTRF9di0FQGIEY8afomBq
mX+otdoWAE1t+ElgkGuWmBQrXCMo4ssa6EWabstVxvG2Jb16XvxeXwPnY8YlL5FfTRpWRuYYE3L2
03q2iXIP65dS9kphH+fHVmlNnhWI3yRtqLc6wkHoNHAfpzwbre/Np7bbGIeOof8357/w3JnC+kqZ
qngifOX0M3Zh9H+YL38kAdadNn9elPnGvpalAu+2P39Fvn0M24W/x14J+TYXBCX+yv/4CqIL13vr
84v6R+/McwcdgeHjyM+DoiaoPHMsw4OkvVenfIEyPB9Jdox4FU9/KGvB4dezbvGGyuXvmoM6VJHr
f5c/YQfpAfyg6guIgToA+pa3knMgJs8h8OnVdPE4XpsvHD1wTsPoqWPbOEIBoj55Hkrwg+F9vDF9
JCbvJLzmSFwzk24cw4ZkjCKQo92QykQT0qnCeVpO9bwumE2UxPJdZF6Pl0+bAWDIaWLddu4Vpftl
S4ku1UWDgPs04msgCgvnKZgLVyl4OcFqTRk4BnDuiFE5fUM4WR5PuDYaOmxq/14L9klrOggkGgd3
929FeqVyMyvBiqgmKZzdkUPmcZygbziuvdJ1fAqsUVtJg7nBRHQjDwKVpPg6UbJVS9fxSHvJhvP1
xLZCrkzHaG6Lsy1BjM33TsbXJ77eoHbdhxndicORUEB6/4xnIM8THB4i30WihCwFFXZBrzc36KsT
2BEZtJUoxsq0XPfsvX2U9W2a5gg6d3oEN4pInTsv+3dMpS50zQnyVy2Cwwz9t+PTOKN06plWOujt
UfoxvRVUQKxymtZ+87xn2TGcU1VnLPBtRgQiezUXAszY4xEhrooitIXPFNy/ZzhsynGm6cD4fSAj
WPToWBHPRLSdq1+PjBXk/ngrAyz3DbFiqHvgPpzniN3IaFD6P/qX6Vp7rYdpjR8M/FPknEyyvTKy
IdMXl3A2twz+Zwl5YHwr2/ciUJYnRuJNNYbYLEcR5GpQFko+YHHFlnx/N7W5vhTX8/lao9dpei19
VMLNK///z2/hSNqgXEQ/keFjDJeGpuDt0G2r4VLjOTaA7EY3XOgYuY/hRGxmWASWc1WWtsCd3HNh
QeMzV6T5VUrcQSlhD12rstvqfwQlLo0NjfRSDqZ8P03qbXpfG5omOJ9IH1KgCx72BC+wi+W+6Y8u
QIAwV5u5Vz9Ok3w8PfOjXNDrfaWczp4xFpRxs3nR+GmQdbxQGeAcFBr73qJq+5frIF8tBauCuE4m
CmEWqNRgoX0pJ8lKVmmPhJJhceNmhurIZWm4NN+m/74knLSXz9Ibo/Cdl/+ZrGX8hw+MRux8LGh4
/64fvyYV0lXGdVMwXM3qIABdXCJu1k4XzjBMYaCbb+G4cYTFC98qFnMN0ldocC/Cv01JOBbTciM5
X6wtMSSJYrArGRO5UhvPHUdUy23CU5FVjWs2kPqCqAlIFsS4PP7Ca/QPcxa3Fdjw/M9Irz/NZG6W
Ku48j9NGoXYNNwszUr5NYsusrzkNunn2PDYBUtlFJE6Xj5RhI778oh+XtPOcKhSX/QeeKZaVH2UW
wcLmunJzdXV00zndmtW2TCLxdkhgINd9y8UghPul27Hw/4RPOv2teHb9L3r6V7d6ZBSi2HCNwgcI
v7MxWc0t7Bg6ncPX2ivUSVaXhjRbMVcSNneuGNt80zSDhMH2nttVdqVl1HniI4ERNXjBPTsDmNSB
qScGk+d2W0wMSL1Hs8IpblbTobKrzAWk+vRszaitnUAx1civxUrMxZGeKC7rtyxgabFb0jN1tEmt
ZA0ABnNkjkLqgf8riUQdVz5csMIAfiyu+xYkqOvTCyy40WR7QfwAGfow4wkyCUiJUTyxyRX0OlIi
X7gzpjsdMdOoou9vm/g5/NQpvumS8pzWh0qoCmkREaBam7jTzCoCj11frxVHnxhESz5vNhXMC0di
3xwptxiCnXHHf6k1JL6oxvl/Mg/Xw5seE8zFyrzRJ3D1dX2meQxqFfK4lhNFvomrS03rpBXtR81V
GMPH5p904RwV/0IvR+Yy8JgA6kVC9SLW2QKZkYDe2GP3SPWd4soinFNh4FFZVS3wydDz/OnnC/62
U+2Xz8F3dROnUhyc9us62mQKuhuWr/Vu5LEVEsKPR+euauj2Jd8GkZ2hFzu7zYcLgJHD0EvSvcSs
E7nQzspHbD1vpxlZ6yp+AuNeHcAnLEz8GZU3mofPQWLDM59aJh5Y6DkXEogMVh69+yTKYPZGZ2Li
s6juPUT7zEXrgDBUGfk3IO0jBoR+W3RC5HmvKcJ9PyGjxu38W5OLsNiXj1cWsBA8NTAZtRuZJ1Yw
j0KATadsHfhZal74n4pHvYTmYe16iWpo1ohzVsCWdWzHFE4EfvYblMzikgrnKZ/nr7pRD102mHpV
BxOB4g1YneL836uHQV2Bjs02GbTJ+NfW+nk7pPwP13rKSv3Hzlk0DuE1VmsQ8u46LFd1KwTtU4ns
RB3j6dNDfjEJeLVQL/mU1Yq+1iVwG1cQ30bXBdyU4SHNXc6gDmxffhYcQfol2OjqYoq6y1GOZuk9
ZapzgqSwNFSiTD+rGRvgVlClaPD57tulJXrd4aQiIY0TpIa8rk+56Skmh6VrOOzi4d03ZbdvGRtA
Jw1XT6eK2UQ4SaNXhLZD1zQ+TFU70Y/ZX/uscx65DrdjkY0AszDqPi6Uz1WOGBLkhI8g++4hms9e
mb9Wl8yQWqB5yP7X/7g1s+QLLTtH+T5sjlDK/o5T7G2jU129FzYLPmqkYGFChOi03iIe+CIPL0AS
7t6GJIk05781NyYP1Bqf6OiqxtJ4YCgMW1Ha9EFeJq2w+QQUASrz18O1rhrUHUAeGUq6QYeCcSv+
NtlNDq2iTK7lQscbpkVTpNZN7497tcVHFBqVUlzO7OC5RD3hEEUThHdlp31ooSTsbSBYfh/ow33K
53bGBPI89Q2hNQmSu76dmtZh4ne6yvPhNhYlT4pflLu9GgJahPrVmKM/2pr5JJq65Jx+bCABb1OW
tVoUWTP9iLazVysSkPoiIBCPNKr6rKXkjgjuuuuVjM5CPvhHyVIz6grHJRXzI0xBeLy4otDbhk/N
UPGgaqYUn2Kvz6RA13QupnV7j+QhQBzxNbdJrV3x0nWU4sNuserYv6q4gel4bdadF/0os99irjHz
XEWVBIwO2AvJOW2eRnFSS75hq6QWajXEoukoSH6v6T9vykvA/aHsYJcwgvwfE4UeHxzDYyP+kTXZ
hejcY7z/DAmoik9SqfGtRTn3HfT9GCnGF0MiHVjSyG3pYDpWm/PcKo/pQKcYgpJ9PbY1aWTSq9Y0
N2gyxet64GUxuDCXIPcc+hZU7U2ho7lw6Bmr5LPuj8Rz5acWtQrWEBt/e1YtElQGnaeqiRTYcgU5
BpJCL+Xirw1CrmEowfrn9WnVXDjehAg360u6sgT7aEBYlIb3JFQazvR9AWTW6dbA6CN5N17DE+WJ
Hc6XlQQ/qg2KjZKrYqYeMfP4G8/J8loMOxlZzxT834gQKCOrlnFmMHaJWPhKSHvShtY7Ph6gXeOD
3rkKBkzJ3SORm7yd99rsnGCRzIqBNgGV6+RuGmhRmjB32AJnQbzS7RV+zK5QrHCoy35U9myJKCNG
Bc1tl5pER1YS0y2Y6Lpfr2AyII7y9j08AFi8BzfRpmJeeIDY0MmefejsLgR0Yt+pN/9ly9vYkoKK
V6oDvOOeGopE5/dbjWffDTzUKXNZLrPUdP6g4WSanEz8J4eh7pHn4hUc47qdqJseeAGK6pxf6qih
8A42sDdgPD3QiOLU3Xqm8/xJqz0az1+xij/w7867a/tomph4QXuPqv2f37ewjrFoR4BT9Qy01MfW
c849djbG+pNrE7uyVeuQhV9Z/AplLqWUrKI4h6GGSVpBPYFsPQc7Z3GeBvUSeBwa5BhfTGefY0Y5
xDYYHGNBl/synnnqbHcPqPtO0eYOKhsOdTJ3pwjMgHSApl9eNIAdlU3ZuhfudyizAOeqMh9mMO4P
4DM6CJElaG5cTQXcY0WxcSGNJiX64klQR3/Oy5apTSoWz8RM7xjvCy/tz57MHjhtOVcjOL2NlwNG
gEsy1hcs8jo3eSOlWNICHQ/ww6408opeDdDDhIfqxa98PYrbPK1EZmMFL1PzbSwxhQXvAaqUSldT
OpAqw+oZq3/dmiS0AlbLKfomt9Ei1sxo4ChCtd9Qf/xFlLt7Mq2nNVraHAEVDY83Jfp5DhVYgj56
dfchrfYx2Zdzk0/4d47OW3EKfm7RcWOtnajWr2S4dXHCY2GZeBXWxqGgXlDjWmsod+0TTZPPieYo
dhenzPOCQx4MPreAPLT98KXRgecgVvUI3fbjLwvjXgMiaKxPxij5pSNG1afa7n6xEWWPuZ6VsG2p
Tef9Qb9K3PavipeSobM5SJ5rBRQuij3a28R8GtSxwY78F3feoweVZ3NEPvOtBK+czv4k4LeY1yvu
Jh7FsMLY9Yod1B8CGJSQEOmGO+YPkVrLeK0wBQWxQoSLoZ06xyb9TVxmReR/hNjmbiDiKZsrRIew
g+MjgpDiGgh4jVRN2kH4n52viDQD0UL55/ikYqFmaiLq8e9salD2M3gWhl4YQKHDAIGvK9zUYYhd
Wz283y7cuQJJVui3mhv7sXgVtFdn29gjhemioI6V1Ur/faTQcUVNeEAP8qGU9vBvHIx+V3/IdABy
vDAnXL1iFBRFKF50kdYB/n3q1/snDll3Il6swLNNvvPnKyt4tniHDE5I/3BDwOEDr/wVtp9qfWXw
H3RB2b7cDIvC3iGEs9V/kj02wv/9GGcNST8HsLdf2rzApPJ7M4CY8Y2y0VLL1jk8qTtOKaCnNrDd
kWNOHFSQLg9NoShJvb3hmOUOCVvHHQVh/+ZczFJsjX4luUV56I9Q02XuWo5wW5cNkYif3Yu5eHO+
L5qlb3Wu4fmF6XTsQ4mqxcjSHL/MwU26v2BlMv07A4MV6206KXunGewvjF9EvmlUsNsgaFS9g1er
pdh3KatyMoUKEc0YdIDoNi1NikVTZcrY09Fzb0wyK5rKbDPGqO8cMXHEHL1vHuvvx9cWbzGqWR5Q
YoaWw6uloxymfEi73L69f143V3CvTQWx5tCOo39X3PpqsH9+nYTXqRzWux1TWyQtHlU0XOUhnHl4
dRJfGHhbn+eEzj96yjZ2cz18ieC0DlUa7w/AorItSNCjFw6smTKC0qQpyYHgcpkM4M5btFIwuF+e
03e3FQ/VJ+GSCpVeCx4ytR5WVMbhh7UfhIQWqk+UzPrf1z5bvtp98SSjNSLusQclsVdnteaWJ7k0
V+H/qyNwG7b+iMjAftYTeCn1ZWYkcs9vAY3JAjrNpJAVriA+CSQB0mdLSn4ZDvOTdc+CIS3ozPjd
jqWL1T9LQaUUfOFFRz9k3PdBAS1UbzSnvPvbr0AeZJw9JwvXEtZWLAIIhxPxwV6OR+dcNnrZ6VnU
C1lPyIB30fzA3Wy07s4M8GANVgdRzJLdfEn9N+l0/LCFdAgFC0pjVBOGWhQxXa0dCXv0NTto+e1v
vODHwsKBy/Nv461Tr6iqbzrn/Bp0IlmpOVliYm6yJQqxew82aST6lW2LNHpc+3QEsSl770hTHQzy
eVUaXhgqT+vc1bdomkwejql3FbKdQ3v7JuFLE7ScfZdmdoctItKJNEdI7r0DOz57dilTsoAirzb4
Z5IZJ0nWlCHUtdcuHTjV+4qaxrXCN/3EWIx1oobcChqUcksjVZ+QBFWdHWZSIrHyniyi4TKUBdH/
yaJcgBo9ErLYwqvT8/HSq5ZW3GC2ssleoxhZU8w32lTZu5avINEmOlfvnIGhttMwJypUnSYyfnTe
03H+JNj8yqCPtNpr1ysvmALycyehA1ZKobaMjm9/Iewry7hrDSue+2xe3q1Sf1/nFdn0M4Mp+aEB
EhH8cdpnThq/PPrLR5xtmhdPadDPyq7KFfQI3XgKLDCAW+9cgHDOg/yRTSf6+Gzx2QgZ6EwsbdTW
5SojC3vZ91IXr10e0VQP3sdCWbDZ8mFXxW66jCvpNaWZ3Hca3sa+bw1cGkHRuM4KnC0IUvSLuaWT
a9ugeZoObUyDMbNgq8BbSMsP/DAueMFt+aDFi2j60StDBntabA8Trg7NCsp24wIxue2laM/QlfrO
LU7gbL437nCtNI6maI4VK/gt5GJ705J3chfC7DIdOADvsxRzln2M0U0fO2RiQ2dpGuYcyREysnNx
SrpOOJOgmfVldmvaYZHWlMY6pl3fx0/dY8n9mr+nVAXOSCQX0mEsGJGe9O+m5Ugy0LWC3q8FGLgW
5GgWQP0jNGk30OQoFqcoazPK7pbIgHeacnni3c9sdJK8gAFL7G98Mp/OnoLeh2zuD/4Pm9ZH3veu
KLD/vrokQxXcerAxzoG5+R/dQGyOfo2qOT8ek4owmSIqGoTDeJmclTa+fMKIy+VBZuqRcP5u0Jf+
5y7cVkV7r6NwSnGk8bFMPysdeL+41DQ0QZ5vNcYjBAAw4108U0teOwy+8EMZcsOpIkE8mZ8SRhJ+
8xazPuE6UTZSZI2x8hoSvRb71Q75LbdhQFaN/HYRFw7bmNsQfvZag1h3B/xlcM5wVjjTA8hFEk4w
kfMGw9QdoDD0k/7GiBpJvS3/tkaVwJvw1gf/qUVLcJW8DEguQSbEPW5L4n0q+J/qvw+2ZAmb1yMW
jHhIqLBjCMK/qGyP3o51VstWiUD1C/I4ePnIVrRYnpFzkE7uHW26QlTKZW1TNu5chpG69EA5j8Am
2FTLaCDiSRdYBFOgyHlMOpXomKQo5VbiWUF86Z3je0pyIciSOX9cVdJtD7M72yypvv5+DOfT4hLJ
QrnG8rBJRAAeFaXTUqOhJEF/Fc6vJZ6PdiQ1zLSuyqEExR6MKGOJKiL0oXzYZ5PPU6C1sOX5zrbN
1e8Ob29UBz8c9qUT5jdKDlJfc9BCeMfEaYuRZs45EvUut3Hde1QjKCN4Reu09BpEIj2c4vgZe5ph
4QjUPLIujOAz9iCexHJ+8NLa3CoISDcH8m7tFKTfni0/Ith0fxiiB9CmGRqovY+ZlHxKnc3ACDcn
/glBn12FxuG/fCcGQv/2M4DRI/TxG5lxgwJMpBS2ZR7l9CFL1AFiYqwyxfY5y9KAWa2pG0ZAnbpU
uRk8wBpf7rBjdL20l+FUMkINHNFzY8piYyNRV2njyIhmv/BQQaNl6JDVsTqIMhfph0+imjrWbTSm
EweoOfYTsrkOgUadxyOTs6pw+ZHh4azJieyAq5MxhGlyxBMq+MFqsued0iPVuQ/pz9LmGLUEwfB6
3PJxDMULq620OJukuMVk6nMenwfDI7lEpRpSX0ipzocecm8ZGqepMsKmWR4hJeflIUCtMLMpYvRo
R9vWisQQHmD3ZRbEiLN4F5DWbNA4mtuI1IVSttqrW2RzzbtWW+ZhXMIEs9B9tdjdm2yW13E3i9cO
0bJ3K20PGDlyDf9wVLUeCt4C19j/9cGBnfsFlFvEgnMu0FiEUj7iwrxs8Dy4Z903VFvh8Wf6GOeg
4bM+NpuF1L9HFely1LN4aRJ4fCcVqeJ8zgqVGmJxAEQKFjLWTN8O8kOx0KzYnEOjJy6fL/b35tWc
B11LeGUEWhkKxHtVI4O83tgb+rMzvOZJJG+MO/bweC64neIuAxy1AZc75WGaNRF2y2TR3ssU4Pmk
Uibk1Yyo81T9NFSqP1dBXRg4Qd5FIx8eBP7YPwOujlAfXTfFhXCgInUAgdUZ+Fyj+qkgmIN8pcNT
Gc8ksksJyQA4X3A3w9ktr1C9WNQwJrIbwmZezxtyhSZrn3hIwX5uIX6XKpeF/BfFfQFQ4z1zEu5M
C7VItVK2kqNFKHEOBL4K0zZ40onOv+Or6QrshGppqqTJefeenGqTffirWnJvelb78kNLvcpUB6SV
QytXVJCk8FIvtcFVupeGtnvkruGbqfEne79dbpipymOc9U+tKiOAorKmTkkVJboFbtVplWcHenPR
QTiMLmDkrQvjZEonU9rs3hyK2zRa3G0IfQVT3s9A3OpNnUnR1nmITCweZTgWfVN+a8ovaANBXmP1
ArbPIDADh1O5LRntcKWbluBqU3XN9SClVfByyUJ04BHWTcLTckzeT4UvKqubHfCS7ZBNh4aAJVWI
9O9ngOTYnk/G/4oyBw9rTylEy07kO/Q+3/oYnLde3vft79kjxPZXUer72FV0y4X/+MFRONvppEpO
Llwf3NA58da6P0tpi+NF8ZzVZDJCN265wewiBZtwVivZEVyGlZ8mHzaMiR5SFeqkeAqXZTxDUduy
oTDJbq8W9R0d3sQ2u3a37d0v6N6j9SxUKSOFba0hzcrwFOq8/rnRiiw+14Ajkau8Xg8yZJt0GKAN
XQ/t5Y6NeirIkH//oXjXkTp3pk9KyiIW1kDE2Vh3U+XMgSIE5OXI4vuGvY+atboE0GxydvRzlJ41
kHoIGYyFp0kQui4qwsr0XCrDgCzOLlDmnxJZvwB18G+3BFXVTfjac3N0rQF52JkAZhAME41Zlhuh
5qzpOnnQmB0kIQdO0wGLrcmXn3IMCnbhiiXbSQnzuf6AhksiWAwEU8vug6zsPTtz8/PV+Z27dgCZ
T2TSqKyQXvAWFldlR3UsAattAV0GPtz2Y4ZL3msOiV4fKTaOYjS3ghcS8G997BVMXFYluAXHSwSu
wCatxUrMU417tn12rud8rGNbcq1P6hTHV++y27ovilVqFryp1s4H3Z1BaJDAdvuzrP1jdllGlbuX
DSqjkNdPGVX0EC4Cc6/3oFwvr5S2dIYnoPaoynk0c1P4ZtLYNcTBMydVIeVt2UGVUiC2yFY1d1Ma
06e7melmazcoEDGLJw72zWXrpsLG/b0lNSj80IVaVUAVVR4Yoe0gnf2byl0V1M7wdVlLzPGiPrlG
zjZn87ftGBjJAF35rh60i74hb9XNb+smviuJSp4qqVgVI0sOMCsMb2Hf7L91QoyqjZy5wRgVsrPx
YTE+E4BQuOVnD32ibZgp1h5eH+YeDfo6dKV4UuGPF10s3ZhFIWHxGbbwHA74sRcUqXxjDSp9GjiY
8KjHledpOT9yu4p12t6LNxCfcFmmX4xwQdZhO5gzKi/87TyuC9R3pmPrpgCth3LQiRW4/cVmIqys
GLWRcVLEkxITPBX1YF3wzJBFOVOPSazdmahfob1iE4/TpNC5a94coIPDi+ipT6b42LzVoK+vupHh
uI8XCghLFL+fYd9/a1fyi/5hayqZyVxVZ6O58SST8eBINu/PbZ3444w1XaKdsj39Ie99T20Qhc5C
UqeyxhFRBl0uYJLsKFekS8GGsv+Oy1CyalrfnA4SLP3CubE+PMBd2smWkV1UwEH4CjOOkuwdfenR
1YcefX6nVqCtTNpezjSeWIj2hY3t0ykzrj0hcLq89cLOjbO9CxUBYhUSKeKvoOWsOy2I/5dg9s/A
GA0edkAT2t5/8uhnleV2IqrGKXudosAH6/ifoAHSfgMS85NNuSLb4mzJl96+kinUJ5QPZE6GEq/l
JIYdB1hP45jIJ/Hb6XwzljyyRX6vYzHy0+6maha+fvTsC+PsOA0DIVVp9qA1EwjvXR46H24BSaL5
1QDC4XRjyguAB1CkEIIblf3ZLutXpvaq7PriUsjGgA2o0BaJBkUmS2AN9LyttxHc20ncM76pRDas
d3a7lu0I/AKRDZ9+Vjzwq80+5zzpGgSCqwn8Iz+hXHxcE/XBZ/+cr3GjG1MPAYucTYYJiU/+13mc
ax7nqEoS1+L8IkQ3RPcmjOBQ7DWrWoz5zHueY6G/M5QR9P5wkg+K9doKZVV31VvP2FbOqea8g6KX
MaWPF8tCpTMFGuH3Qa22ztRQQMPvE9v8hY0oPQMgcchM/OCGwkepok758lKm9KXlgyhhhjIk0cwn
VzNv9AiKryG8wR/4CkDvO+FWXX6T/ZvQfypA8f+rftM2fLFAe6sjgXeFblSvnL7XORPM6lM8DqVU
qW8hep0nGykOtd5o7PLjl2vK3SdG6F9LUJQANq6gxHfJGB+YwDNhzCYiw6EvoygvviO2xTGBOV8+
flcSVC7IpnTF4ic4s24kYmhDVzJox8F/0KKhtYzSGWhp259F/nK3HF+QzqgTca6iMJtP7OVYSqmV
PYTecUo/uDOOijpRhTFA+hYB9xcKa7G4TKx3yuKieOMdufvzg8fDY5lDQg7BSTU7EnZ0TMxqMn53
LAhemSm6DbAHPJg9t031wlIeVs0D/k/H8VzmIIV98ainRA3vxaLj8X7y6NAcPXHkRjiYO02rAHCr
3ZS9FEdN+9/mJzNHSUhhOshFMM4aQRU0RO3cP9RrwtqU8MNG4xXuGw4/DZemLXKDcHMQWtjqUNRf
Zn9z2ggZl5f6FW99QL6btaQ5tdGvNLGAbna2Demq+MXNwhnOEl8xPR3YWXR5RgwkvIBqxHDKdTdW
ubnMLHoGzxm5quQd6+EYbUMT98pOatWBcGgpquL0jFWfoNJof9i0L0hkdYl/tcC118kGcf4spMsS
kl/DGNDCoFK9VsVWBQ88RtlRueojGQvhBJk3ixj4dChRqzuqPSIpvTiHnY5dh8R4SdzhG9ToLcoA
5yJI/C8arQpuaPWezOXeX+BXEAsPA5D1wcXD0ejzGoDTZe1/5A5SIbJtpFdU7DOdIDhOV8OZ36FB
QIsJyCj/SJL+oK0UsgLb7qGirH4X6XyuWsv5s/SrDY+LelaeflMghwTqJM9x2fSxcl1qYj67vE3D
FZuzfZKN2D97ToynuDhGDZFbzScFHf+Se9YiNXoylwcezQ5xynC2A4XMROGQXG6o/o0esyiPwoH0
skS1BbIdl+WwYLXoK50pwhRsuT/vnqJ46bb4IDmE96PwWDJGWcZ7NbAGMu2zHZE7iiTeHFuvpb+Z
rp39UuJPooTdUnNKuP6o2w985sDwyaOsmpSBDyqX0D8nuZri1bIKYG++xB9VE4aoCUTMRwUG8Qly
B/r8HF3b7A0Z1lidtcSol9I2O0jifoSLhdCbSVWXjkCUT7TDJPGrBUJPSXlfGKOcLiXvdRicOcc5
fXENVT3k+LSPa16vCfoEy40BPX3cdnzsAjwtbAGYVmznKQBu5Eit3/oKnBe26c5kHpw9RUDLnvw5
GJP8aZSPzIJX6qnewvQbMmxaio7Ktf9I4nEz29zzemUWJjJtQV7SljD3AypUI2mWuL/p/nqT/woJ
p0WCgXPzbSpW0WrXcRYA0EaHYAbjEgPUTdhAKuu5+hVRbuiKv9qvCzmmGsB5MKieLv4K8axSSx5U
mAPRRiNSOj2M3o7GK/LipoWLRnRvuSHT1EjqDcnG74TyfCqZ+CZEOml6yAxNydHMrb/Sy89ht8Ye
GfSdhdcZ37j3lpCspxK8yVfavHcPpPYs4yXzfb15uCCRcbroWiCbIDk13PnRQuyVWBndLF0XxfWl
UD6kgbVDeAk0d5XED7lpx2IvVPTKfte+bfY4rVs7vS2CeC+gfZl5dZ16kT2+4jHCc0E1J6X8ptml
JN7s4h7GzuD8fUOPts3o6eqcls94EXVHq5m+B4BTuUvoovssxjL+EwJRfRa3mw5/zb1/dPsrT/ld
nf0BwcMf6Va0vjqSGcAKxa39PQ37nj3Tmq7Q/Rbu01ET/rj2pleinZqHk7VTcd3dp/Ce96YC7tw8
6W2vETF7OmTxj0J0JNIhIwVNW8MWQFzkgkElxBe3w3tDYMNwdgjXbBAaH9FG+afmIXfhmrxqDvdv
mdwZKjoU2Rs4xCEVqYmkgJmPueov0zBEdKeFlQ3J/6MWISTEEvWXicPisX7EXWwfg1kAU5AFc7Tr
Vimxg17ctg4PEmidzWPmNJA1OOQDbtSvhhNy4Zi3qN9o4D8e4uZxFGnH56LOlGZc1pmvXBL09VNa
n2rgSWVcnBHTXeKBaL2eWPeFkUpilek3mDKT4lX4fkHUe8u2RfSlm0AqL0DdTRKiCEphMcwgIJUp
61p9mw+hAX9duUaC5k3wRcPvjsEF7840OVfUINKmvMb5wM1ST3J2GNr1YfkaUYRIWJwPIOrEdLxq
qcgtTj5iScU9UMcp0KvXRyJb1T2A6c20kwg8tuJTqIZLH7UsWc98f42Ks0Ftdm4ZfZzn/1FKhOKG
17MUatYz6LwDOBEqMi8kZqLBzv6m4S5TY5PpnmWvc6Z+hbI5M5MHH6y96ZAaBkKJ1sXHnO4xEUUx
I2yUvs4iCtSv+JmZxiUgXzpgmIsWyPXZlMH1uSFhT5VQZaht7NjIQ9rObth3umb9digvnAWJEseQ
cqXrZ3qGxVae1ZOFgeL1u75Bg8KoKVYKC7PoyQdUCNOMlZo/Hj9Lty8mEtgP1aaToHHdsegSVg4M
4cwvwYkRePxOExnoIvLFhfrlclFWlS+FdO/xFNEpVMqieRJcTj43MBiryyeGKd/tSeKdytuI1l44
gO0sAgLoqEpj6nrnYk9oWLJbxJGdu0sQLP14h2AdT3Iuw2J/jn9qmUXzILYQvPLSB6+KmSa40sIt
K1bwpM1OfSkc8mPHX4xQAtttocgIfaiP/zgH5mmWAR3mr/QJlyiQ7SQIHDpT8PEP9j1ez5960r7+
jAhFQ9f57FftofVh0eu6t02ebFG8RHb+zR7Q6RELbsnb1cU25CW5N7pA6qIFubWYxpV75FQHJ4cD
HsIvnjYabzqTcYGmUr1XlCfupakX/4xFD1rp2cFpgtXe6QSQhWIYncPhmmbo00VrYvFovJWBXB9G
M4bHrRPwuhvnH2ce/XwBAbN7LGoNe/Kn4bZvXLnuF/NCdNaJpy6mrjC0y/8jc9+42W91WV5EGoJd
PRosVn+s6R8RL5uYNNl1G88TeiZlvur/R87Xia2dh7m6p3BWCSFy71BLWJBeBW4OULE4HZjgXzP9
BdKGn16ibpHaRIIK9wciqEDn/Fayudvrw2erQ++ZRrr+3Loju2wGx0J3iCpDM/rXsAxpbKRJfbNh
D+EnzXLQ1UgCPAuftugNt3HKTRHKMCi+je5QN8/Q3ttoIbb3v6rOa/4ZsB2rJpzRxgkUz/FK3KXx
SQlQ5eXz7jJeezM2v4j3opiBJyQL20nLtZlgp5BqiCXvshUcX6af4e+6Zy6lFd5JDn/npddEeuO8
5fek+FLsKujmCfs1xqSlo8N1XmSGhfhs4YZsY1bmdrx3D+HEfZvEH4HA+1++GBIam1X9BO/d/l6C
7+SP+pPpOWYryLHA2tESAf4DVfqLRUE0uzbxAKtSOh/YPNV8XlFvX7JtS150kIyYPYiX5n63DlMe
uAn+o0sbUb0xVKUQNcz6WkmsKtYF1wly8UUdbwYWpJnQbiEI/2/NFdQU3hC6D3KwY8/lwHzxcZbt
1zGw/8f9iQVG4pWkAovuaLNLmp6yssV5zuQTb3KyPJPKczpD2K8735yZowBdGF5JMgAXu1xr5t3N
pOvNpkjkZkkDYr9G2P1oY2zDh8bxvvHknAmcSGBrM305RuQqcKGWX9ZRKYQlI3puyvtqOqrWYVMq
aIs9BRH8Dfn4Xy+uysh9l+w9yyJ7aEs92PWCgz+fmvno9/jpYqL2nUbyOXwjPhihDfo9hfHQKn1A
oFUy3yS2s6z51T+YhRKUMfdglVI+40Cnk3qY6BOJcJTBz0Sv2y2PoILSbjOALveRRIcSgSjKkcj9
JxAfxBr7577plCH26FwY+rXd3Tvo+fUlBmgIN67uAjHzMgPkcSfQwR88MxpFh9ufcPhyd0GpsuX/
qsNZbjvA8Dr9TRTEIHUBR7nDCJnarm7HStSNPd5PmjAuZe/VlR6j6+GJoEH8NDxnlZNYAN6al17c
/LoQ/qoRRHeKI5sDFtHeTt8oOjqw0bHpAXGeErph+a4DxSmuVX5TgCFenCWOsvbmPyOauMQq+NkF
3I5eQ1OiiQNlQTHvUNy2KxHOUzToKLQCtMYXGNRgCY0nYRvzfAAj3tFE+D/4oLVbJ208s8gcqxT9
v1vLUIVr1pdcoxFHDQqn3eB88CJnsGymLehKYjQR5SzyclQwbjHI+6W+tZlcqNQdbDMJS9hluwEq
LgWR9LTyYaA7Oe/xPlBZxSowGL3p1WcWx/qzR9we08u6zkxbRlcy/b4923o0Jccsklh5jqQYAlYc
w1YG83sk3q09K4rPsojE2A8KLhJCJEtCoa0H+yaLSwX/SuiKfj2xSfuOnGnZXbvIfZ4j1tRqUHFN
5ByCxHyMYG48rM7mj5KYs5LauEJouY+Tc4XU2rRRj3yXC6lPe35eIPKTdx6CAW7UNssanN1JHnLg
ShzHvtYsCl02H4xZGinhn36ToaE176YuJvPH1fvYBiRFC0vVzrpcqNMj81/lizZZo7sTfeO0CxBs
X5aDKeOjFPVDeNXjqUJj9OZAxHyb+WE8lKqKdcpXCwecDu6lIFtFr6O5oPLMDyOiHDpuoo2UofQK
97wD1sRfOOb8QBpD+xvSgSJvVdksx4VmAkfFWsZ4Mc8VCJfhA740gQILZFFKRrqzUJoTkxYuwzz+
2jxmj/bJhadjN1oxdd3XGM2MGpQtp4XzJGFG1Iq6JJUOBtAs3LHC9bTAxMl9Gqra+NYqWcLSMvvA
Y8Yb8ELbwYgsZyDz2v/v+YWZ3V8EfVGXADBGvsxqx5/aXo7b1kcxoC9KNR6Man1LWiIlzpv8igC0
5uCh3cCvqAN6kkiXLcSgWB674nBxkrT9PonooDrhbXhk14SdwlKY0WlR0P7QRBEOEQMmYNPONjgQ
xHoyN1uI9HumHc13Rtvi7y6a/RWcX3dWJInW/0+Zrafp7vLTDxmMu8Measkc4tH3jkF6Hhg/3l9O
j4muEvPd9IsqwcdAW0Eh2uupSc3wSuDLktmsP6tdiDqTWEuyb2ST+j2FT3IlCRwml7V+HR8DQAXi
8OTUVJWxUGYYBxGyrVadClLYGjzSYyPocVDISOzuffhw7QgzMdCof46o44KwORdXgdNF9owcwlUC
U+fNtSZvIsZNvrK7lvvZjMwo/Ul63XKcf9zZ2VAO1rakPK3eBBFR+gznI24Ay9RqTczEWGYq9kdY
EE4pJqr4hH/VtUOvjmlbCk60bOZa2Z4CHyxO3rcFLLpqpfBWvdrW1UG4N1LSA5+ZIu+PNx5U4++F
LHXGd6XyNGJRQ/opFieRrV0qnLqYXO0J8T2fwyycesmY1bPquJzi3GhsOH6BX/I2bWB79K6UBmDz
eDsk6NG+ezyhJ/v6z6IUPQn1Eav6AAitMwqlKnaRxC8I/iB7x51eAU1pI7p8qP9mz4qcwXXOfyvZ
gw0N9T7FViBPU3LXkvKjCmemcrkNPzAr+I0SRS1Y+BM225PqvLZKJEUJuU8PNnD3uheb+eiEQO5P
9CsKm7GafvELG1+Mzzr9G8BrVO21t/eSgsyhe/2fb7DtptLaKmd10GF534G32toifQXUIsoPA0jv
N7QAwE/TcOtdVYgh6l/Ipz53B3TJwtcUTm2UXQ4I0TEpP4ETJAeVMJWrB/jtcJNJXOInHhTYFHRQ
nru9svs1BTjUYzYgmUlYLqYRqd2+EwWWY7N9CsROT6cdgWeTowv5NtKsDRCmNEh6/AXldvbEtkLF
MTn89zBcAEXXxwFjMtHzy3R1QFIwoUek3bSwp526EK6t18rQAuA5L6nSps9dnJApBqtwDnFTJUBc
l00zwYKxE2+L0RwRtQs784AHDFU825H7TJ+nVZnnQlh9egXjj0qtNK9Qmpmv/rsxxWQpljGm9CHB
M1wSFY05FM2k0UpdDZWJjrB+J/4Vz7qEiQWm8ph0MZTpa7DX+SP5RtWaw2H/D7rNuNMwx6EwHmrr
zLSDLWSTh1+2AWbneSUGymNXnYhcfJlkiNqx0WrLf4ohsFDFiAZlx90Xt0yloIT6VMK3Kxb+gn4a
hOfFeKb9noY4t0+yWbLP2CaqpJ7OZCAO6pxysuISWUe5NjMUUf15CUu8whRwO2o6vXoSQIR5jL20
80+tpdZ0QWhBHNS88Cc19XhEUNMqoq5AiiZPYmF2Y6pQhLZPuzNrcm3xOnjDObPtr4Lfd+hHfWxF
MXKp8xnb6fnw/6ZZ0zsH8p9UPK/aehskt2lwNlh++UoPW1zj2ytkDiQF9rMYfxU5E8c+lBAXzdiF
NjYs6jaq+SKbJbeKidrBO72O2QdRPw5OKBx/PYOpcNbzMfPkYVAXLqug6MP38LqOrAG7P2c9k5tV
AG+chl67DpVm3mq3FB9gFouqKPY0GQ+0RkvpPuy0KdwyqHsv6H9nABmMn9twulmr1EQgOZoofIwu
hkxMPVTQtIi3bcfZxX3+6xuDgrvEyN/liz+cCW8PYYyAqGRduNDix0BsZH1cUZbHWptXUipmrJ4A
ydZ/s8Tm1FYw8cFJNl9llgmgJxjtu3T1wRtI51/DwZkbn4Sfa6JQAFG1dXWnAfDK9kjcFMMlPapd
jRpKZV6gdbg0d+mmiAYNEU6HRYoe/GM05RoOSv4ihHOpKt91iwtl4LRMCbAOLmW//J2kby35hwYj
mhZXv1Tvi6gpXQvosCY462p/wc+96/mW1nedHL3f4t82FTmVbkm21k8eI4so6N5SxofYW4qwQnq4
uDRmCK0Rqpj+3njeAR1ZVsYdyIl3uEqgV701FJbWic6x6HSIPYexHKlQosFBZxayH9mka8umTbGK
hPHWCvJCwyH09JDAB1ChdIVXcCF1sACBUvuc1JVJ+opvzlQ+APicQ1HZIRTlcgeznGvJg7nFfeXz
E5iyU6OOrqZK25f5hCDcGJ4AjM3F3kClA8Y58DpKkeBUBsa7QZmajg0YN3OrALZN9/gqrKh2eD9z
Y3SO0lFtHO+nHFpQer3ZAvpwcEkmehtDU9Z6L12CyL4BU6P9n6/ysWS7FXfzuMVw0bJNMRxoSEkq
e0E/BqGpLOm8OFlcSU7zft7G7bbwsFqm2JZpAchCHfu7TW++1QEE8YsN15oEBFyvcOqIqph3shD+
X+PfAyLW3yyVEANrWy1Iz/ANeyIp3RQ0bwcSe7rhO4t6HspiLUnsx/29lvoQanwc6Ka5rnPRtW7w
vRvuDqvANSs3fNSY4P8YHTffuFQsHF1MwJb9LbTXOEbgfww8aAR0blb9N/XWRuGETFaefi38iFDL
JJTC7nB/LupWTT2zuspMJJPVzu8HXsC+SvfirrJ1mlMgyIdy+jSF9PIQ/Xx9JRTu9YpAHdNbNoGs
5pp+jUwGRTAwcphECjzc64llSaiC8ytz6Ng7421eRT8KG2FHaCHDj7uUvch/orbaKiSt4pnlUOdY
8fwMcX9GoIAQ2++eFG+8NlhytGJ6ZdkHDVIoeSqaNDZGQAByynaoxbnGETDlWZqtMgGM4ypwM8lU
QH31NY5CqjIX5VqosqFVHgzyqqRdLGcC1yXgaum6vY0zoH24A7+Kh3bb9betyh0IVJLl+FAX6BPF
HJfDMDyVBcm2Q6itlkV0wE9oAJ6WvXQ7LG3kBBMUudm7Xniudc6e6OCNJmaY18esmSzjW5kWOeH2
qsEgrmtRbq+MHvz8+xo7ADYOdovu6D9t/c5n4CMaq0lsvXMvQABDJA39ZTeHtLzT8B0jNjjCwLT/
IVR5ry/9fQl/Yo1YKSvFsVRL0fxFlaaqIOcy5/WQV6j/rxJ1v4F0igrqH2AFDkzGxi1V0Qv0No6T
eoaKWQUeAPNzvVFKnH8kOEZwWz8H2wqfZ18Q6eN4tVt9u5E/766MSbbCEVxQzkSUJdAW1ootj7Gg
/MD6pNrxBYyLzFqCXJGYmgTgoirkzJpB28aQwlYfPuTysl4wZJGzx/g18lk8+53/c0JSngIE1smO
q9lIxCznyBxFjF72ynS/jlRpftYDFgOrK/CNsr9hIJRAi4BgIMk0BQEEUwwZMS9vHuq969Oo56WY
okolYpsTXUCDAjQIN6Wwz65J4WXBgby0PZyqVX6y9nbSNg69dWHU4Wq+oHA4FAQmWsNHRX8XOBqO
/58Urp/WgSKnxrR3qW991kow/jYtUJaixLh0jKkM6Bo6LJifqq+8//+T86uIHn3IwxFOsIn14sxL
g1bGIPfELL9QXhBKIy/g7Oi59Ev6mo3MRgtU0DUrE/oRINqLn9T/uqBNCz7P0zMNOHcydqJdGdy0
S8mmB2jthOefXMERzRUXN3020jUUowI02P/0ufMYdhhUxg8xmvtsdvdmwtpiHIXCxwam9xprPiVK
Zpbb84ngifnvK+teQS9P0RPUv3WJ/W6lm2rnRNw0uS8wK2pjTYDGewX8RcnRG2Q1extBncZlI69/
/8pWTqZKeSP6NSXDqMz+qvuWFUTodYTUZBAoSG4WJFNprOvCsyBB3q8QE3Dsf9SxTWl/2G2newBv
KoVSfknPeMRAhkz4y/Slm3Lthsjn86BujDFmvrPhA5ShT0cvKpN7lakckCoKlJnFaQ490rJ1SeWz
3Yd6PpKJx9GModqKFuOnqLZDOzBE7mnv99cEYgWrIi0D9Fd6Jv2IjuKRxcCbqAKcgnQj93A1xOQ0
xrk9RNP52VTg6c8plZadOseTI9Gn3NVqMKDTh3SJI2tPutC7mYzm6ffVHWnIXYs8vum6qDGgzNKO
sTxntqtytoNEP/3eC6qjMo1XT3WZmCzRmEcA6TgxeY7l9SvET1mtku8hmi8P0kukIbwaxB87Da5Y
35TVS66LA1WEq9kXINB5rr4eP0omVn5YrYZpq0mG9Rv6rlhIxVSSnsZfIu7nnto2NFc7jzp9P5LB
ZQSAmX/kZI0+n5jko6cPTCDogMJsWU59uSeU9GggA8ySZA4Yu7goJwSnr4LzchnEGHqobOaMFr1s
LmrJ9iLxgMyo7I9PAmL5CXVY7QopR8uHYP3Yw+X2npoex3IJZHFq+x4FVEPDBHq8/Gr+Awr3aEX/
zHk4/gEpcR0zy3HIup2CNt/eZau7raF0zMob0aWYhbMGjVA/3/TgsEwnTFlWdsa7Z9r3WzblRx1s
vZRZvTjxnU7TkJFCF636ovZzCOOGcThgtR3fHVc5l5JTpL3fR0gxG663yqD5T0a4ZDwjhGasIddG
IHBxhuEW1XRy+1spJK4FAn+9pY2M4hTNz3TYNIitOAHUABhvJd2UPl9fHIkv49ncZ1Fn1l6NwDsA
dvzLgzVVs+damkJsMkRBoK52Y0QzWAl/gB6iURDldPEoFYL5qtxrDCgBt4mu1J5ys0JS9pqN+sJQ
45FW5arAebwQII3UZRoDUz9UTehcOPYjrtfC+4znEjph3Du58GohhMvek9XbkUMo/+J3rhtvzEGK
eM93ygYS85d9Z9so3IXlVmVoBGO2flkpSY+wbYvyJdpSMErL5ToYy0Fo3MIrOeyT06wlZOce0sMU
koyHIydQvEwdh60escB6xJlQvjX/7xOPtGb4f3oFil7x1YbElSZKXgahLmG4UHvxTqHcoG+SWlcP
vKOmvK+A4pZfnwcPwyxfEt/paDubtXtkhj+cfZcLAHhpiSWNaF2Y/QBkY1iCyUimAWWnD2lAinqA
xE48Nk2yQ/Cz1wp9bwJqRIVeYqmedb2M2Mp4d9tXbqUrHO2ACpwgAHcEtVP2baquLLanY+sHOw9c
hYmOyn3Zvx7JEGPVpw64blzB88Mlo1N2D4XCLjNY4Hm5/QvPtvbEgFEtdH5vWkLfZgelyrmILBC+
EouQEqi/cxLjlSpGlmKxBZEMjTrNPxZRBSOW9tAbCbDNpTPrQtkdw0c0lv3Vb7a2v4PKuxgQdXYQ
9fjxMTQfj4rqOKOwhsuHauINBQMmM2ljXqG7shddHy6tKzeIPePAUOLCUOuMeuDRHFfi42YWV9O9
Zu/A0K5Y/RPEMRvZM97+3uTJei4zNRXnNelk1/1ZJptJgMeTJsi2DxOpB302+SJb0+ECkWgQzplK
CPdSKmmmdpuLAPRJu41vguUNBqZH9701GeNzb5FzSEXL8Gyc4+XuLCQmUeV+NYWAqyNXEP3Yg5x6
7ziy2Aa46u2v/A0fg0ICkO13L8177/3jNkSZ5QsUqYKwa0EB0UZMiGr1Uf695hsl16dOnoLVlpyP
gVVJDzq7fSLOY+nl0vVS4u8LZx2pI94mYtv+Qscaq7oBoUti/1DQig3e4ydkUQSkKbopwt+FXvr3
bkSRZXhitclEv15+/3MeHHpouF7rjke7dDpIoxcVpTbq1SLf57YWpcO0S/Isxd2kNHN9l613y9TT
BIukG+N0JdCgO5lBSzoQIiJpk5UKFybQatenMZWn9AgIB1xHO2ELG+LXLRTTdKnCrXyT0UoTXlyi
YdDz0D78JZ8SsnwOqU7d8Q3CUBXFV9Pnds6w20dfKmDm3EAlmwA8HfXI00UzGojxfgnXiZAhiLm9
FOcyJSrLtDU/MW4H6s0As8j+5j3TYTC0xx54cEQzeJvqNofXp6ANP/vnTP2R5xSO6cRDYuXDb7zX
DgcMr7z/HDbYRsURX9Gt8W0NOokj7XRYXluwB2T62A8Hs8E/ry/sckucGHv4exQckBtycal0l3ho
ZmZ8seHiD8FN3JtDZ1XyT/eCZnS74UxK9uC+9JWriruhVSmsRu6npa0pvw+CWpwZgmxmtruzleNJ
FEFskJPKobv7N8E0OtZmObXhCOiQJGX3+JRPCW9dlUuYpPlTEPc72bA+kdK7OQ1bVL3N4GmBRPSy
3D3a7IN916JO1TQoflg2KkLxP9Y6wfnKa65pbRH8vTDwcLuanPNpzUYa7JGWjzuH+0MhDsymLHBF
ftLy3o5Fs63gUr7HKWj/9nun1sXeN5Hi4pcCxJJZuzsP6D7QIU9CQU/lMVQDRiVN+RHPei4PVMxF
V7JTfKN9wayLrWK7l+boZ/wQHMGlz26ndxJJ1IPTG7GD922Rt/03s2zFhlOu86Y3F06fco+oP1JW
kW7fNc3L8chWq1Quj/b3o9fj8zQxL/LpgRhpzu19Y/Ieh2yk4QVH3vTv7BmtXWUPjsbR7INp4+C4
DusN9IgMA+DOEY+Gdx66nSIEWAg3bc/xhjrEk5rA8A/LEpbtCHRNVxOIHifdtBgNmlt2OPPshXVp
Qyh1Gkl8WDw6ZleGsxE/b6iBG+FY56xUjiqPPVJ8p3Oyb6WcQtnJfhwC2TY5UDy4owPLHq5ilTZZ
mht8MIih6KlhpcGYEDbZ9jv4oKPzLfhKzfOgcG7s26zSLrP2NS3w0OIeHyT0kSJA3Nw/mlgNzv8R
L4u9LnjqW1EJz5dFU2QgsVkI1bfX6TwZCODW2vw5Q+gArmcRwEtYW1IUJRn8/5VBiFc7/s9Opm9Q
uHr/nbwMZgPU/jSXG/kf6UUoNu0cBq142u2jFzAYw835SHS17r8nEz5sHlsbaC/MHj/LKOZCYsJ5
UqbUVB6GOuwHU5tOMXy59o4WueSzOvtdO33WcW7grtGc0ON8KGy5ASvbLig6MBDnhmzUZtzIMiyi
Q3WBxNlPQAKmACCjFaqLnZJUIsMiF5edmbRXUf9jmEISo7q2eZ4eD1qimq+6EcpfduJTVeEwXWRV
B3wxovaD1DU/VEP6ikTQDyUDsELGUdonUEBdI4isfeTVU9ZoM7YD6De1VZ7Q8wDWyOqlg6pu8txm
TZvQVDkv946duRcUB6K2idvdT+OQIXik23Bl9OUoiGgTwqg/Quh4CVtBM9dCJ9/LTsI4YoftxL4u
hclJme3xBIBVkMT22qakWkeDhkH6wEKftzJHoOkDY8CechmcgpJT1dE4QcW+AWADYWd4GcLU1zIY
NgJknupI2pclp5FwsyYonlk/sa6/2J3279ZYXZKLwceiNkBe3ffdZvF7MJzT293lMhgNwEOHhkv8
b4Jj2fMUREEv2blBBpcjdWF9hRPekip0oPjoQK+sNYOtmuI4H+1tCsx3l+a9bZKLdQMmXlqY3oEj
Vn1hg0G4vOTvfFnRaUj5USzFKq1hwRVf7lUBDJ+j5YZkMuA4BitbRUC6Vnz4bNd6nPHEsEDaWn3t
JcVTTFwBKNDinxI8IW3rCdFDpf1NbZEhr+ADPXKm61R5qxyiZQnZKJv3rriJjZzsvg2BshQmp4yC
wAM4wyoMf9Ag6H+TSOqn4iYH8ssTeFGz0xynFIQMFl0ioutY3an1bnBkEfvAnr7CBgVqjBaKXfhA
PV2YB9wvQOjtIrJkgg2gSgqvzMh10SaDCrnAJ9W6tcrjpTURzItyA2AOmfmDbra7ZW7MkMD/fDia
rxeosLeiPzscA8G9LxoShU8FLqU34yrpFVPmXJsljYNjaX5/Vw+V8+jAfmDmTii9LnrkrmNPUACS
ucQ01l/B4PS5ztUOc0Aw5w/4HdJIj07kVErIjN/IchkGQLC6Ig6nP8ebd18PS0TnlvfJ3EI2iJ8b
pgsKd5BJXXyrOhBnfTFNfQGaNhvlX8AjfbV7LdCXpaFf7uUq48FoyyJqfg2Yl1P88z4BP6CNmeg8
Ly/Vdo0PsXXIu2Elfm34MoMvJR2KykVev6k5dG5mitp8aOWjh2a8r/P+KByN3ZRxh9tbgaKA6dvv
VH7wHLYq1xWgzFZ8mKbNPW8K7T0XuxsGImeHr0JUZvHFymihKxTZpG7DopGX7hWE82QXQV8n18Fp
upFifEHN6nnO88+uvPpKcsHUy26YNzI8GhhYRi9TI1DuEbwo8h75LPIUSm6t3ejNxd7LwDDx1Vsa
GMyOv+AcRHc9E5Wp/PmFOmv7/d4fYzYLUBSGsSbmWGzy4vtYZ0bB84FsBLW9AL2psGcqOflV10oL
9wjn+2DqADbjsen4/KVpgGXW9iRpcKclwLagR4Oi6XqVRltOIEdSMBPOusmslI1/dmyg9PcxoNaa
8vkOXVNeKLFIMrlqnDjUEFk7fWEcfsg6wI/PcoO0AQ+K0hoG2xaAqPvrBN6H4mJazN6dsPjp2eJq
tCljKxchgpVaCenhDNydtHYfyw/6qlo15zoQWTxAdHwM+aaf6aF59Pc08nhi32y8WyBt5SiSnAh0
RBKsXtEUjKFsQugYS0E/5vfjY+EknFL13voRKCtWxAOJNneL6gtO2w0Ulnjjk6vlX67CUIznqd2l
gu6FExFzGHo0/b0x9sZ1mkrblV7KPkCACG+zzwL588hzOtT93axaj0tLl4MgJYRBxqLABQXe1M9i
lHzTk7A9L/QWTt21NuOdvMZfY1e0sctD7NuCOwVnr3q1DG5dkwufqPlnHsbfqDczTgmnB5gkQJDf
i/a96lDaooUap1z+LUzaewdPKeY/oufA/A7/s1Dr3ix18zyfpoz3Y/+7+bh5BO8THbTynKFz6frE
QOcDAi0CPu6XpmH8SQ9xLAUpyteU05CCyEkrBuXGpwSjxceoc1I0tFnQXsYNiwZyfl1+4NoE7tXO
rJ08H7AvzKihV9KERQl8gJSdyabiufw0BnluyWo/ay16TZ6qiB1n9d/N/2gxRAN3k6H8GY37roFC
rwV9PwvfsZDKNJmQoJqgzDjlUN2nthsQmVthNueZRXoNPegOX3tQnKU30OqHRgIhOl9yvd7OFu7V
509kbfb/mgaKk+urVzHHXrgN7Q5Wh6MST7Jg8iSX2sQ2Se3Yp+qPns02AN2Wu9uBSBnH1Um5V2vD
wpvJWdsnqpyVZnPVuyo3QAyYe9PMZBmcnsmfZH7hERYjYi1MgFh2n6a3LecHDSGopdoCvT/Sz2oX
iFfNsr7/sX8y0nJC0wHA2G1i1zauiOYk6XlAhfzudVMQJqtqRCLvs95R5neHCjYTC0DgLRGZ44ye
9LjoxNVIk0GuHfUCZC72rv6ane4GvAAbeVtnRFyRQtfLG4JO6qN4Fqt5fPdcq7Ij5Kdz7CC3yUS2
mvVgngOh5w2Y+Yhtz3SpG9vQBnVYFoLHuKSSEBZ7N/SKFtGbm0M03DVG79JhCOeBn7f2SaVFqboT
e2dSWiqvaXTdeAt+TRm77Nd+naUP3p8uoz+lNhwU0XmnySodg/EAtHMayextWuDT2VzNxt/TeS1R
uurSkRbtFi5AWfa3hv8sI/wG/FjxFOtAwE4LT4uWflg61HmtRji5UtCS+nsMmWk7cuOY4aVsDPlD
7bb81T/HpHYjHn6rdIhfAD3QloZj2KgNIizUYpetMSh3bEVMXT5UCl+8gxDP+nMaOoVaqx/eNRwh
f6vKXZM7D60rHeQV7uLCDQuHVEu4HTzbBEC0RWhHRu/AYvJ7t48jAwh84H/n0D1ERuGVkVqL1EQt
C4VpilFjxjUPsV9sioWPLXaaYV+bhd9vsHwwglTALLfWo3ZRAjlqYcZSrwmgQwR2S/jdxCZZJ2qK
Ef9MLE62/NxRWZ/1LrYc+BPV5miP6Z64XpTxHFikGrrP1h2ZQbmNrUSvuVZhVsyahLwBGLGeLQ/9
c1cwWG393Y6Ux7Ob+LZ0H0eyud57kWII+tVI9cra6Xl9RBtR3PYI84VDi5WTjhD5M91DlnxK4YR5
E+vitLJ3j2TVqpb49pDQtYy0CGcC0QZ6ZWOTmVqTYvOWVQoQbTUqc/K6FrzVVda8rBGttc4CEyCH
OpOFwGVY2rRT5kL/fOwnQ6PgdyYsBcz/wWQKtk8LT3xcHeIOWtzB11T7yG6beHSh33EDzyFu5E0X
jBkmK7joXq3tz5XIytiG2Kk1hqchLOmHhLKkz2YCzMFw5vSxTLocON+rB9ek046Y+O1Ebk7uTJjt
mZMwNFVvY6gmpiU18IJVQXnXVw+UkwtqmjrWbwSTJZVIqvqQuDzpeSLz6wRHx4m+hwUmC4IiRKJM
ykjZwU79KlFA7mDJKgM1lXVfNDFH/FRuWItAT/AqWGhgQs2pQA6NtiEpqW8eufl79B6ElM8HFLZG
xTBxXbR1Ae10VjYALYYOArmP0sa7sEGH5TADciPfDW5z1PnqM8gMEjR7EvAeo7DKoLAWLZ03G+TX
BVU743w9BOJ1iaodZqFqc23kgUAuWcJoV3Qnr5vn2Vy6+9IaPhVQYo6uxWOfQr3zsDsTrn7xnEsj
g7A0lKsGINQlof12Ee/BCasn+znfXSJs4G8if8hU+VwkDLBv0J0XjyukDXSmDyV0cw4TDttzwMhj
+Bv7xaRo1Sq8MUo5CQANOKZdjb6wU1e+URJN09gQVvv60ckw06KWgSp0SQAdAF4Pr6hLOZBauIoQ
MDnN8p03G3LIKVxGOsmEk7SC9WCA7OEUNWLJyE2yR+aKt/E+3yzRE8hfmp9umjJCkjTs0mHN1nn0
YZKojI5RXS0obcQGljIdOqRKmvoINj5Kck0wtRu+HV6QH+qq8RgFMV5xsbfhPUoVjTrdVJbhL0FY
N4A5RRbwiR1nyWg2piQADh4DLDKSpjwUho1QJDVjGneqxcycj0KU4ldQcrLkwV5rgFwrELSN8DQN
lFYv6ZTZxwudlHoQq5U13pW391xBnt30TqzH9WDKyTjBlBp99tryXNh2pCS1Q/peEq6MNThNVHua
bcNsYj6HOwHR4wkw4bDP46yTX3jK7WaZX6ljEQEgWtF8p5sFSBZBWwsVzezqQR7KRrTDk4Y58DTf
GnFxa9M5mTqrEqvc9TkgoZH4Kc5LKB4Xr9ZcjsVwCSsT6OKIJIag9S8yodTajDp6vm2YeqYdNPI3
Hlb0PO2xN3w0+azHgiGnQ3xyEZ8PKAWlPAWxq/KFv6g8K4Oqsndy6pThq+/4dosjx+m26b0wKh76
FcBA7TGp/L1ZiOFXuOIpcEPQtoOBR8g3YzBgOGHCZaPlcQxmds6K0ID5APkK+bzRiuVm1Uy6CJHI
RN5/1CizKNVM9nWBO1oBt7TxHPgjbTuDfFqcoYOfXtYA7EuhDlq3HycFlkHP6g/oL2IgH20Snoks
SpRCClYirOLcgyKWBsMDsPtp7zaBavdFMfi2K7ywRFUxv/gAHbOcRMReispc1wzC+2bXOzfSTYtx
TrSgWVeFIw+8Q3qS0lJ8mK70yMI/hQk11f66hEdoYd3uS6iWSPvMuHuqDm9vPISFIGoFUwqWtZfF
HLvGAEIEmwO+oP2O6d0oS60ke3gcVk5JEgm1ibzIE6S/198Jp0grSeecd90giqbGV/tdY8xC37HV
6kbpYRIN/6HUrPVRSpbFNpbdZgLRgmxmav2G1bbrL4wktc4iT1/QjYIffVXuh8O0IGI3O6BLixsq
KaNb65iCaoTecPFhD1wdchNfjJECjYQRbHKK3fhm/ajXC/FIZthDAeTONifA9gMM/OikikgmRfWr
ol0g4F3l7knmM3gLAirAQxmYs6Y+z5OrHANw4SWHLF4eLn/S+Whmtbpi9BHL2JO1qAAoLi0QvWHb
fMkOaMuXJO05/G2Ws4pQ3DnZnnFY98yItpUhco3RqTKSthH19+ghuRZY8xmbPIuv4ZpUHiaZ3I2h
52xSlT5PUFjQ2q+MMEaO52HnYxtMNaerC99yYl2lQ0BJrT7JC6B0dW+yfKvyxvEB/1auTpnrfdBL
GUPoJU1Hl5hC2vw1eGeudTw7wuFmSPv2vvUaOY/8M2Vl9Epgx1mWZyMIKccSoRRMsyJpNLlCOqtE
ZfNt9pi+OMgYb7BuqeLDHvyLwpLOY+15QgGE+1Sc3/LgXOkmZQoMZw9OxetQnCmM2boq/dx9AfMo
9a/VZoFzlAJ/pdjcHCEjsf2KIVDwZtDDOYVEYybbrU+YIzJYmsjAJw2JeQyOwhoHpeKlSPpp0J8s
wFZGu+JUAenzzBJKq1cySqDgr+aoG4RPt4SpbXDBR0G4KfY8Be9UXUxIWgH2UAVQQYjylA4bVDPl
o3LqWoTX5inMRyKGFzQfSy865QqkPiyviAuE9lW/GA05ICxT63pRBliV2sOkytpBJxDE+Uif7QsO
/Z1eAW6PpOdav9gnGt+V1jtUlo+tJl8XfC7cNr8eGyVG/CP5xgX35BeUruz/A1a9B8ClioqmDGCt
CWQRw0nXxwljlnwkCTLXs0s8CBP+EYx+nmyw0egtTpvFdgrbvGKteqh3G3It5BAzqxq/2Yz/86Q/
j8URKft35ju+zYvb5D8TubBz7xJXxjtjtgytT5RZGWd75p35ulD3Jzd+4kf3dyJqy3V6R/ww1SAU
bwU6yZDERa1Q8pAHf99qzVXFwfU8DXOXPsZ5nAbOwWuqZ2P8M+mhS0XVJ/hihVz7zdRoqgW7Jwy4
30fOOp3oBixPTeQRRp3vZkEB2sVvo93iO1V2339E/EVy007pZqLZf0Q9OjzzWEoJz48mM1CmYqdi
KzDFekQki/HFy+WvGk8TrFGm1GgB3/aCIzB8rV/FGjbhRKo8tBKE+J6eTyLgMXx4hdYBTV+iATbA
WvucvPltBbkQoHXNkVGfUvAnSwt1HUxCYlcE5R+aD52RoMwh1vjM02qWFetf6KVI71Bc0L8U41J0
kaBS+T5pkW1bGG6QT40c3+hdD58h+XcBZlV/VnRl3ffzo309K7xc1DeRImv8NfBS0SSgbjT52poI
ksneDTlNCerZLZs5RX0xUbACccA4da2qI8OeJAqavAcxjyGESnJ2qApTKYJrGtN3JsjgJ0ReGYxp
Gdz6+LjHvq4pn1D7EaaA/Zse3WWEfCbSbgA8rz+A0v1Epfegm5cd2LHEr8lrFdEt4QA7s5Zpelqt
O5Hn9c3eZK/w+FWNmtZIfP++2gbJ0XNOzALDeR/G19KnGI8sQfSbtngj7kGKnQM+l/ovw89Aijso
6b83lmf8lOLeE6G2WW3x9A2KJtZpQB/nmx0jUK3aYpf7A0p/kNwdYyIrHWPSIyDiTbQqu4YyTiUh
74Cj3GlofZ+wRPtBypJJZG0Krqggsk7mlugN6Lo8lie2rzk0X1u/vJ4WKegvrzX1LSro/VUI4rJG
wLRX2bKDxYURAbGipcSRexggDhX5FnBodMffgDkErLyMRXpfuRJ3RQrCZCDh00lSyrMVdO/7m+8l
qDRsUDcWt39GNSvedu0etvhEXbkuN3sDJA2ENkJt2woYtNmYsVe4RZ869U16j1nwlTpT7MKPtsuB
T131RNdafqpN/96CkyIil4m/wV9qFxWlxdCxCTa6uhCsIcIiv/5VPc8ERKePeoAy5E/G2QI61tcx
HRc9XCUcrzmYtT9vxbcst95ynBOKS8DDYr5m9r0rTPYQyPJzjuidRa9NJg/03fFANVgqDMDg3gO2
jIH23+KfgaLxuSLrlGD8I983Y3jLHWYIg+l4OwpR/lyY4/tacLcsQuaW2m1EMOEexX18n4iG9PBP
kuTdhOwqy68IOgf36LqiWfe1OhHv8NDYY0cl78vyFJXgWNSR4OnAzJagsxR3Ihi6/bb8Y1j/79Jz
ahSIrNBAHd7SgFZvJhI37AJhucmPkvFUG3BD/kzoN/icidPQ4lxJS/TUnFRMj2fP0nQZ1X0TxyKf
9GYTvNFaRHpYJUET1iowtEb7amf5xqptMcOKAsSHGg4UHZvofKML+WCWunWy6N92r1yccKAnSdPc
wXbH2lbsFR7flgZm8Hpwmsqnv0HBZwMnQOJhVqy6fBp8n6kC91QLglG0cMktoIFetpBsZydrDrn6
4F15SOMpzsi/S75DDPeGlT66/uyIHnetU26ZFIbScyLZKchJdlpydaYNl5JOPjl0NlieHBBoy0nz
WuavFwg4I2UFSCvbrau0vHCLBbodFzAFlqKbRePjFpnFsEnK5NQ2acZ8OSU4iVM2gdGwyFKuhibw
EKCM3+ATiojw21Qak+rblnqM48sSKidynDdMIHSd9cZSUnJCRKUWFQGLe/qo/t9bP/8+ODZYVtY3
GHB7snrqO7zy2nOpNNBPds+TBAA/aP4WhT/tmhAtmLT3Icd/QpuYRi1d0jTuCSXhrfQpTEzfLjJX
kTNR8fPJaKNVcplZDWJ1p04LOKaavk0FVkj40Pb/1hfVy16VBkT7MaunikKyL+lxWisvNhPlAGXQ
1ZQx2TdZOFWaCsQhZEYhhJ/h6k8g5L2BfMllEKl2VhAmrQOs0NBl+0JKQJ82zUYPqBK7QU8hcLyC
H4ZUEoylFZ7PmvCnnSCSCPS+Sfd0B2pSvWbWWlDER+eXHwkKHEIdARAYBm3A8jR6m1D0y81rmn4x
tx0R+tmBv99rVc0QZKwkzerya9pC+2Z9LRCriZshTHElMWLuzuiLL4M638sNBViEmGx7z1jY3jyJ
u7Yq6xvNFTg0J4bqLb2RebtXJqqxBgwKkLD5qTKD6voKlJ3IQip8SD+BF/csHvbDFGn2a5kT/ypp
1Qfa4ZPUZUBA4oKyPkeKWFtXLFbQKtqPhq2AEpd85tCNMfhO97aNWfISqeuWl7y61x0YkFV3vnRJ
eje7Q0YS0fo91b8ze+zxX3++Hi7UrUFtcTr8pTiveBy2h3poUNfXRFp4JfXHG0EwMuq7RCSwx+pY
8OPwPRthhGNKx/D0uF+jG5X4kQIgqTaU8m9+aWMAERJifNurxOe1Bwy2kJWcw7hTVjE8+z3GmHiO
AAdjpx9CzZS51lWSaCy7ISHUmX/+BrKVpoRISj4N5yh6ubTWw3g3roa7+cCQn38zkmXOIysZl08V
TnWTHiVyERBLvR9o2t4x3G6qqsjyfxFrvTqer9+8X0sPegPfNbPqQUtPN80GxtknXE22QqFobvIb
pk1sdcRVVEa8MURDv+lX38iUwaDnOh8MODyAqPkH2TgSgORhNb8UEkGGB+8PdfcxKoOl59ZNu2/y
wU4LMggt3vVxsr3H9T3gb1zIqQQ5HS7TVPYv6Y3ge3kNoluZc8r1n6fzRV19rSsZCxSiCFx4lJSo
ki9lUi1RxkeIzYREv2gG8ZxyuOg2BxNILVZgyRR6yncPRobqYPvqGwqEBl6LtyiLZJasJUSu60BV
VjKDsE0rH+9wnyTBUe4mrr+oSWbra6r1CM2jyOTTHH9WkYcgAh8dnJ8+I5laAqDbH8aWU1uNIudT
yhRzwedRpfbz2R6LzNRCqKnkERxrsPWLUMzbW3HbbSezK/nWW/ZIOH7UoaObI8d8r0beALVyDkNa
gMMEQF7AgWpZoIdMnKlQ7qOAW7riJ+DSZOR8YIUtIsNQgGIQ1fERz3dWRw85yJyKtcEGHb+1mM58
jV25IT1M2V4dCQ56VBjP0LlxvFP47XejdhVsG26oyWwRfLdk/Db2XtM0DYlcZPRDt9PxbgU1WmQV
AbGC3GeYvkaBC/Rblc7yeAxfc07uwxx+/3Ug64Tk9VJG7WSItScgtNMH178Jno88MV+nJecb954E
3wiuTrR22ZwlH33htYE51A6789DeeO2MNSLFS8hIECREVILEccx6eEpz/nI0MVZVrnVXYnACcasL
wBGDf80ZOLjACPLRfHmbfihOl2VmDS48W4I8xA5OUW4mRe8HYX9yC1A7N3Qe57VmDCshuB6s1Hqa
6BKJ72nsH6z/8CpL0UrGFHfM30Y+pBkoBgUtQja6WjUryo7ZlvKm85LrVCufsJz0NVOlV1fMrW5U
uj7POuabi7cfsH81tzbntuxaOo2cJuesrpuuBPDa81AVee2EEy6IDNRc9RncF4dmBnaO5GLU6giK
RyZcTPprrUgLDWJUJvebvUhXnV2U2pMDOLVrI+u2ay8SQod8PLgE8Q3Y6GvTyW1pC5ywgiNG3F4v
omH06EUPc38dlL+F2cJ0EZozMGvzAbmWnbJWZyAB8dxWOQi7c7LQfiVtIhipPtE4go9xCMOrdwgh
nlqKIMHe27YYi2ygnWZet6NR2GlCtJt7cEKa74xjp+O2JSfXtAV5IMlfpxKkWpp3pu/VZFmNjaFG
DaSEQGUIYO3I77nCU0LX5yL3mgeQ7i0hAiS1OeOKPY2DDD0yQ+kRCbv1hVpFlh+n8tRhHy2RfaqS
nmtG2084aLe3lX23YjnbuA+6UrOUOXka+MNkGLDLaEOdsHYrZmA3fMe0fOAESE8QrFv57SawYblV
NZZxK2a90ezrU+rsYuZBEWizZty8vqdcOzVX9/77b3PoN41/eMHG38Wd2AVBnjf+qFyagIY0SWl2
DVwKQAbId9lyx4cmP3vTlNmm2eq9IKHzJ5gmnUTBusNhvKlfoM+/2MN8iWtPpOMH2Mz18Busu+qd
Qcf5hf9ZjxfiIjjBlqBGIxExO+43JD1T+gEWPJRBViwyyjgyBoersIGCC45B0lmwEGXzff9spi65
ncUCbWKZBK+yaX/NGWfSD49vFE3VgXR9sn/6zsYAjYFG1CSw+R91vtYWtWTJ7F1fVyTMIX9ISpgF
XiJsUPbC64IhTOhU8qQN8MTolJtoW/2MBsv44+0yyj/L6/itBzVQ8fCiQCSZd23MOsdKRC4xhg8G
9yTrnHRmkLgPxdWOMowKaXsbKO//qKjTqBJTz3rIMiiQB0uMBy8vHp5y+FXEzPynYS5GGa3z/wRz
0O/RhUatKCYxjhXw2OQ1i4wDt3txxyYvpfFKm9fKHZj3MQRA6u0HEEgQ4j7l2OgohpoIbZLSQZUY
S+sd/aIXAiUappySw85oj5L4dUrtg2PCRTIpnJkUbFyxYLNn+VK+mzuUiW8CRSbFZhyi5D9oNxSA
yoAIYqTgZZkDYQUNGDvP0T1zzxY6NX17btpyZRlnezqo1yEs0IWDsbQoYiA6dtOxvoGUF1C1d8n/
Z+RE+QOEsVj5L1FIDI0m5rmdKyXjwAXP3Ni2ugOA8W2asG62r0s7xX2Lz372cpHkUqlIjR0jlgVa
t4ENkVscWxbT/2Ul4vWR6RJSiPXixu1NSL58YAU2MataJH4M0gKaAb45FahR+YA0ge1xuGM/DcvW
i3/19dGRK/Ntb+NRHCCGdyeUQ+KkPIN8ajnGH98wSk02N6kbNEjPE9ummX8NAIBjqa4s5c1LPMXO
NuGtfe4Kv0WRFT7DVxKB3OKZrgCUxL7UdcLZE7rNkeklWfokCsPmIxiVWqWxhZoqKyrYY5TcR//g
0pUu4EKmQoqXtcpHu2UvcOhVKAgYV9qUuFDotcbpFNwQCIhgdSEuYaNMDar/knCvHYl2+0LDCV3k
gO3cV5Fssm04qhc1wISO6y8mpF45yH/H6vfhvO9dRuohiU7uRgzbVZg9+SDifincCbs/TJj//Tn0
LKcU1S92VbTNomjsLG06vDdHj+VXJ9Of9R4PhuBaJWADMFnQdtYdfqBMaEz+yxPzFgCu/ytKAt70
9xcjHQ/37v5CL3w90QgXGzWtCcMHe9BdVHW23QhIU8Feg8xMb6lqGB0Lki3K0tSECz958b3WtWzZ
6H7ThqsOgSYc+fQ5l9dFP/xISVYCvgTUPMIWttLowF5kj1NxNhjLFt+pG8RqRpt1KSgiKtNJlDcy
XitWa3w3hP2NxEYW/29Z4H77CCKOuCIjga/yz6fdz6ZVH3Yosm9P8dI4TofWd6O9GAJzmCD0kTXV
M59xPAAqIijfkg/PWVwd4qFDk4UZwy/Ol6thciwqzR2r5lbBfdeiWFjg7dw9kAI8JCacl8mebLub
sD1o9mGQrG89i/pL5nR4TEor779mMru35rxN2nFSKzn4wttE7BnKxvUsAUH4Dclf8+ZpnYZsnQCC
dN8A4isCw6l0JpxNzvx+de/QuulDgZgcWdD6tUHVxiFQmW2gurT0TFSmyJzmwfq8HulLwDKxS2Xx
ljpBzrTyYJEfqUU0xs05glFxyjEDdvvwcexcp3zwKUDFSTcIC/DLQYrSDUEQMdLmeyR/iROJIsCy
mUPcjUkql6u0fGtZnFsXSXw45yUuwvssg6nP8J29SpxzEsmcUj2aG3dOj98qjj/1Bkb4fd9JuAB1
atxrGOIr+d+SdvhezUF7PglT1mVHub32/upfPAUX3oEiWw5WCXvRZ/Nr4jNwptkh8PpkvcKxBOkB
BcUHcl2dx1wmOEmu1sHqD3uynf2DPeL3AhfcDJQMyCjxnuwYoQLLu9aX+x7lL+x1L6qfcClrTZwt
SAXFsnyZWb4Xg4bxHWuUxP47ZO4ccM4iFy4VRpLsDKDO+SNfXh7TWTcwSoiP6Eodr6kzRwRLcAGK
im6rAM1/RYC6NgHV25i6q1++UfKSaYDXngzKqnOaIODw3qaorBbl0M544mtNXKMUwZusRlGaihw1
7mJ53BDDhUXBgAJIPelRt106d2h+qj54nQhSxjpur0+8rHaxlhHGjeeMkP54sHhgH24F0WCF7+tR
A6ej+21tExtAsysh4pmACudWfocJcqs4FJnGNkAjzd7ku8eYUwY02GpBdX8uUNIuoGhCLCrzEyaG
Itqe8SvyqVimFSAloHObVd56qSltka4fE3SspwyCcA8myaP6AqtQhdY8EiTAbEfwsdUFneA1v5CV
UmookUkamV5xNMm0IFRiTVga3M7yhMTbUhzoiYnaD0w/sfl5sdjhcN4iPxzF+znj3/oAROg/oo2a
QLz7ETANCPUm/JK5MnTSkCOV/ae77fZTGNix4jXsn2mXWXxYcuTRrZSbSz7Bq2yBRIhvtCa0MAKA
O7EUXjqDuuCbkMCFTLZDXJDlfJgDgjRyhviiDPvEfjHpht35VnM47P5FYp6bMQ4RqLxzRcsNs9zQ
Wftyn+fEZ2CloIPN49QNVjewF0pW7vaFf0s2+8bnbNZ5+QelL4f66THDxZMzABUjJ7tDnfhZ02IF
74W7EWjRa0rgxnQv2RyvCjgZYzSdm0pqEI56AshZT8TQdFORera6+zfkI1isebPW4omnCjnijzVG
6D1R5h1AmXtfm7FhJVU69bxhCjRRx82R2X5g7+lHNfG8Q+XxZoY/YvMAkjmFy5GUIwsS5Q+a3BUy
O6FfWyEBNdlqzsyyPNkRMsdzJRr1NDr8Wwl71m5lt6vKL9XEcySghK1mdRn36YHevVE8tqbGSeqt
xPztgImTT3jIcmiCjD1/4p+32gSK3j/F723YBlbg4Ewu06C13ldL+FQCyyk83d+VPlFxEYs1PY2i
PiYMZCjbPt62o9NLS1m6tS0eGLp6FhR1SD2zbuUMzI3E5dilWqrf4CrFR1fjnuOLUU6m0iP93kEt
6NSRzp1CrodSJHZ+OlrWj0tBnJYA1w7xQKr4ICtibClRxeYMEpaAPaVHkDzI14bydH/aIo0qLg43
OREn8lEQ0Df8Q9L9q21Bsa/eZw5hvq3/LfsLGVmI9dh1x6Tfwgri1Po/8yBALJL87+YOqy1ZgzGo
D6IsFt5l0MV4V7G9X1LcA8D7wWZJe67PuvWdQ89lbqToEg+YlWiXCZ9q6EelOXe3lYDvr08Scks+
9iaKpzxNjRqf4xHZq5tHfNFgo5SaQSwjgoRC5aak8eZeQuvMkr3EBSLoJsRAkcJL+ddZnRSxvnne
wlGbdKYxobxcjUd0w9WWfHXDjiEq/w9sppZ9YdDfzz5MHBORep6cT+JqL1idjym2ymBh+sWrdvbq
4XEHf1YEEnn7R4WzWXpmGf0gp2b8PJP781OtwaTMm4rFZ/M2fuubyEjWMzGVTzImTWaTod8gD3GM
Kw8Vp4MtrVSoaTTLLLmN8Doe2tMnw2Cv42CNGd+rj9XefudUs+MpOb81fGGHGKzvGyrDTR3z63r9
ukjRWioHzfSHvRFExQVwidxA97W8C2MYqF/APv4Xm+f56/Kz6NGue6imjOUAwTtMRMgb2W/RgWTs
dAnJJNXFfE9S/iNL/UXWMgspIZg1w0y2hmKkWFlYKk+gdqbfA7e4MsxRc9MD+DWgifDXCwaD2Fkr
zaTeRssaA8SDgwm04PwEA+y0HDvSK9qN2br0ktwYZyH16TGRvtiRU78LQcY/mZnR8T7iQch5LtSy
GA4gXco4G2BuNu27Iyek5WqpXzdiK0Rcf0zacs/PFzStPjqluOxuOKk3TEgo4JjrduBtYbgmsJsg
dSy0luD7qJ9Qi32gV85cKHtLbxw4aDTiE+e10eENQ4acTmLMFtpNp59eelv9S0b3Lbr8O6hA5kT6
VrqbOqI5ScHE+nbnNluQEU+949MU8eUj6QKBHH1wNIQMwgf5c+TqRMglRsQztxsp+8nP+Pd22fvE
thSAiqJlgdcJoDx4Oku5lvCPgZqRoxQ7ZL1lJX/mHwRcIyL8a+tNHvxMj75sivAS8w1zTNrYGB7R
n94UFfr1NoOFLWoXBdq8VTdDSv1zqe/+7bPxPEqJvYCeEn0U0+s1dON8M3oSMsbZKC5Yk2tlZdsE
bkoQW8VO5sl/tN5ax/GV8fDaY5eOWeAmiuNknB8ms3qD3QzlL8tV4kX7A/cMHKZPhNT/gLBbEq1W
ktWg9x9CC3Tcc9uHjMbspzC6gATlFJ6yKuzMYD+G+f3zqBNDlIOW1fQbzKBCSd4KE9cX0VN5+HWo
sZvCb/AQF5yWKSu1qDkiRfcjBs51cSU1YLmwKF3cbnzRlgw8Afau0MGvCMy6GZn83Mt1kJmvSRIl
LQYupVOnJuSuYRAFespKko0a8uG4H7wMhZf61ScUTdeXMHKB24Z+7vRpSSd2o/ZSsnaOD7u+HWdX
dAKj894alDe/MUDSYwp7yLnUELszlXxUEKorYcRG35gk8njt+NWjVdp509VSCJ9+dIPvlJHebtTt
glxUu/bqXkLabAGf5iZte6+C9cBxLyP7y3s7pWn8rx8ryCgGGCYTCa0Fn2EIhWUOQzccLGHvVRHC
KDd0f1TFp/venRWibSNOPopDxR256STv9GmyVB/TV7aILv6sDS0dnYSHFGDu4T0FPOypGZnVNqDl
sf59NB2NVixiSSxzjGgETgCMsx8CzV+tbDZ7Jra6RAF2EXb5GeRfHoqezh/f6EJnheWG8Epg2sPX
NQqDgWrpRzsHc98WIDd794AD7z5nXabS+wrGSFdeW0gBXdNhTUhnOkIvnHxCkWgKkpE4b7pD6wJm
dxO1t7fqfRbZy7EEVh9jAZx8FqmOvYwjGZ96Ei8qQPb7YcjeonGQcFAJa5xoN9hQN84cZBTJowg7
KZV7u1hkFGMtc5BNqYGiI2Zp7k/aJrOjS6+3iC19/cwnCFbkIjxND3juNeOLB6DzIGS80ouFD8Vv
/V0SZd8apXB/E3hElX+Td1UwqknzYiUxECIbeRWcfBC9km96zMBTVL1V8FjBIJKCdViqx+C4eNor
AxZff5roJ/xUc/PCeSmYCGeP/Si0bfQGSn2CjTY9C4dw0mwFjyrQYsjWyExhhGAIzse1FzrKxdkt
L2a7NmclumbQp2yB5Aa7kDjNpTz+kUuClfWKqCyxiZ/WKHuCNFYnUSZ+EHMvi/YAexKY4N0Uc/zH
Q+bOenMRZ2E0J111+QHAqAP75uAhqk/jmMJZ2vqWwmFqu/EzRbEwrAQXWIErZbB6DPBp5/Pzc8P3
7Ssko9xxvcsqTMp3JsOPIExf4At9WEqjDK/0wOIvYCpNmM5593gyPSGW2sRK2VumMTcg6wi+1+pn
KHvCoGffwgmZJyK2ndYPyJhLN7YXtsTvMp6e6r5FTATf6Ss2p/38Iv8pLe5U5g1ryV3d/57pwyxb
xvNGuudwiBX5kjyFAPT62eQ5Cin2Ic5DpUfR4azu1SgcNm57fWtpD9ig9i/H4ZraxAqc9EnS72+Y
N8ouF/k/doyZ4bGCcmNEcUxCAHfnKqvSTmTZmsSWXqEEuUGRTaVnX+CCDDBeLLN4qkp6kAnSiKL9
j8bc0alVLIVG7WVyhqwCjX0ePtSBVLM9a57d43D9Fpj+oU91v4zFW8CD/JS05wgrQVjkUtANd09w
qC/pHLU9zgCgjXGXKjD+pm2Dn5EaH/DF3S8bv25hxK5y+Ehc02M06dbmqEr8YmUlH3iglhWomh/l
7BqMbIMmD3fMJ794OCqhtemqugnOHrOaw7Ns1cQLdUlXdZXaAvmyRPfyS8jM4z3hkxqU8Vtt7FNs
6zqB7EXlWUdF4vpnmEg+IZXJp19zk4ezMjxAHdC5sA/O2xUMotCa9AOfipSPY9b7of7S9GNUKymi
8fpR1iruw7s0URLQwuiVBc2kZwkyPSgJeqNt/ZnE0KKYejGPABzYvQEfEtt03FMSaOrMldqBuT/R
lTkcCqrDpsUM5EwUAy7BD4Gsm5NAWdxf61JP5Qtyt+QAg7VvKqujQE/bhTmEWDNNO2bllOES8ykB
uw4F9OL3Sehc+wNgpNyR29IkW3qWZlsLNvo2neKW74HOpwu24orS9PEm0mT2M6IT5PPYDcTbxSXG
yUKHm8XZu4i8M+ciutp10tcqL5rE+7l0u7DG5dG4ORUYaV1670T6P747v/iBRhtFUOGb2P2vjPUQ
xc0qw5oZr/Izqh8cx+BChJdXoSlCSF5h1eiuPlJxgYHNoUiVZ1wG07YdGOzsh8+hu2/wx+bZQwjn
VEIcaU/E3HkZFVoKwRAaBqsFCpsGCVUEQcR6JElVIpFfLEbV8m8UputzoAjHCTXBIAauqMNH//gD
SAOVFLKpLKTgizhH5n5YdAauL96DyQWL5uMwl2x+4eaRJrlBE5/cmi7Z4hdvCsBmusetPIhyCxOt
oSkmZoQBxklnmlTfySKwvGI4KgViE/Mkaj/VbrAZdf4NqWRqD6ANbo+FPPqzgQFZzVmn4ncdB0N6
+8cPo0DnKRTuwJ50yWIVb9ACgy/xxVtt9Rohmm8+qRI9jeMlfMSr/71mBuiEie7sfxCuo6ZpKF3s
YMPFXl+amGyLL/hQ56bP8dDbvCCRaEuI0Ps4GM3VmpcyatwOGmcfJMYacBoOffVmC9tCN30nCrtY
3kQ1IcmJ3arx4tP3jOONZkGAYIMlszb4LJ60jHkHAslWLQwiBfBsbdZW3HlPkCW6WU3gVJMt0Typ
4M7k6VDTzk7ySpyUq4gqX8U8qZK80Y7Aq1ITA3HRm1kvai/njFsJxgaJOR+CQYSCXTN7MAzhyQN2
1FawViEZyxFZ8i3KlE3SHn0MS+VYwqUB/51Lm09v/+2GHr4BnFu8t0bDV6bwUIFxUYGzwfliIRu2
WjN+kD8JNiOdX4V3nBSga6zBD12hlwxW3Xlx3e2OJszUGc07Rn/WzITpskW6cKyaJIXuWgyEZHC4
UMYHVlQK9jBO72qu3gCa+nUXkP+S61pTYsdAT+9x7w307K0PooEbVE+yX0i8NHxQPp76Ngr/zw/m
Kmtt8bTZYFkeNdwk+nRNU4EvPXGHCpCnXE8nL0cVMMMtAytJJ2dbBBwPTJeiQc5dz8jHVAWkCuNF
BwPSY+XtDapJNa+0TxlM41JxiN2A8OlS7QqjCmSMewpxhOh647ul5DYczKR0fEx5SDuN7Liz/vcS
bUrlcsRh6dVtOKfoAoRT1GwTRPj8cK93xb6WWPp4OTYISCdPNnUcYAoS9O2oQAa6lobv04K+/FcY
LIklgrgpdxjiipwWjyVbbrXbj11zbEnK1t+98ZGzcKCFdAKswoxVsC3tH+3wIVgDoFR86klZe5Ew
f2d+vf5sUV6sxp4OPBCyPOKE7JK93YolMsMkY8O+k8cmQFIKC8IhzILU8wGpniUc1d849XJWVnmL
aAshklivarsZ8HCREuSL44WUggd3ahadMswr/K4ltUBKoVDlhvffbiyiQ/yHEvvsJDs9IEc/3CvW
GomZRcsBlTd7kJTqiCsMeQLzFMneL68l00Mrbzf14sWXaWYRXdfy44LDVBOTrtVJJClcSdncy2ZN
CkYf/6aFrVU5MDLgYsNk2EzObi+kxRhvlMa5nixl71a0WzN3hlIbq/mRf3O0veEOyeo/YBtdGR0h
8+b1hFUlQHh4cG6n1jSJwt7rpfGWdPKbpWRcMPlHYckgdcOLDlAwsrLpy2Xlywtu3LStgSB8JdrJ
RIAJPTqOsnJqgDJ2J821ym/qP9ECDjPucKpiTafwaorEd+72X0EimBqyPlVZgvpu2Cky67nIA6eY
ERHzdMqCVNqkxwWaK76FCr7OrA8ss1QPQxTY3QVT7TMQM1zYf6d1zvypT5M+iRKhiRAEj0lVhvFS
f9M4VCpMGH2siQPL8zTo6ond9VJzuNeLPbPdZ4MB5OJdHydBZb+s8JszWOO4yYr+dLFWJ7YRxBdf
Ow/XnDY5RElJBSecyTlB4+S1HrN1OA1hkkGsGvdAdnm61te4Jac0DaIRDEXxfhyQRnpfQ09EexAl
c4T4XeCbKrtDA4TTii8LSFUtRGzP7OuCvqJNMHTf22ATMER0icb653EuA7j1T+yKyWcDM12eNhjq
sXV2A13hOQEnMEme0DXZqKIUWy973l0Nitmf6Q8ODa+vOlKVNt+HUaKsTxsw9GHEbgBGN4WTYUuA
nao4wJnx6PVdWDgBn65elr1bPXOnPcf+/M7oBdLXLPE9X/XYU0SQUemV8kyKtN/DIi1LRGEbpJSF
CpInJqrwVlNYG3I+S4vYnD7yEUUKehz+PwBaBcXWeVn19DWCeziDVvD8uuTMKLS3BDOmK2fwqDs4
iJBCn+1S7dvIl8mX9sXfp3jnnaDfP5WGvvV75fwmn5cV2kphjK1zoKHOa6CdwH5yViDCbkwPm3Yf
Zo/myN4Dp/VSeL/Ktg/tq2JCPBBd9kXN3ZO0d8dqAcsuW4fWwgOWdjYN6uYwv2m5l4mZP1H7qNAx
BuHuszVXEtqKEx6czJvFopCab/4fIAIkB1ntnDnqV3VcMMOxYvxD53xnJfwU+xNT0u6i54KQDTov
ZtecMU/gHyaEs/hTIMtCBQ8PYXfelOCKh0+Yv34ik38Y4/8sAT/xoA0MQ5i+H84Newt1e54lf5mk
IG2zUE8oPVxFje6TlUv9XVTAOax6/uHoj9cc9vvTVihph9FB+JEkc3nJALoHbTEwptZYP3hMAkx2
fijgzmRA+Zqx2Mimm+U2826qV5MjIJZ3uRggRtWotTjKBsquaOf2d5OqIfUrn2Ofvh53r3cqRGm5
TsQSaPOtQT0ZZP7et2lafNLhbOkq/oL2UGeYgmXElcclNDUPpL6p1RxFHjALLu9iT9Kk6pxnOxyW
af/tsoR82Kz/6gv2UeH0EiFs2eeu6ULJzpn1L6Ygat3tOJTGWaUF5j/BgNUt6Q+pKkDt3wQdgk0K
dBVbPEPPz+gUkmCZVeb61p7L/DZeuNPna9O3ZTz7ZCBUz/bZmwW5h2znjQ6eHxKG3TRn0c4tiRFH
seZT5Q43YIOA48NHDEPIYVmG3Su8uSz5q+WtqrECGi69hE6TR2b/JVkZLZlW7Gkyg818RF5zTXIL
zS9Ibyx+KTLFvKVQ7ir9AEENDSjDQvHz4gEZeJx6Y1IKP8NzzjRS6hEAwl8gQWOgOU0abhax6Pxd
6JUJL86oX7iJpLcFZOV3G7nrToZf4EyygEjOKx2bSn7O8HdJ6BpjgIdcM03OqDa8HVrn6qot46GD
Xt8Sbq1rhCe2MJIlhqPtyTEKJb6POGCFhlnTM2ptTKsP9kP01Uj01ugs+rnGsJ6rzAzipfP3GQri
g31BFBV/wzUt5FHVnZSDPYUTt3xgSklOkVhieykbB5Y3l/GtUKZEcCUTYu/uvwQ8Ekdyh0EnJGvg
mQpuq1a7oj1OnuwmGwju6TRaJPvy6ZbgzlSitSZzbtVAFs47F5Y/z5vmw3whZcIsj12ulYvONk9r
ttDLXVNeT2/HRVuUWoZ4hNtJvTwy2RdAs8M3UappBsWirHvxy9czhWUxhuq5vhBZGdEgYh1sylk2
6lJutCIoNLczRIFwECExlz0exZQHc4E5DubF7L1YGF+0KhbtnGgvHYgERK162e9HMmYNBuVQVrVY
BSG6IN/6G2C3QSfkZfLZ4/cYlY3eWWFvu7X8FKq6lzs7fDCe21TGLEVLBvfrtAadc3ZMDB89YVBW
Vd6XJtEMCktRn/5EbFrcs9kRmCLwbXUwO9Z/ZVmuv0shvy+XhpnA7d9DcuE+ylpsZ6ojpFqpyvvD
xw0g2egwUd0gHbN9vT5HdiCWB3uV059D6MQcsRvHjZeLjxICq6PrZa4u8weyvOfy0Rm8ZFkm1teR
doSNy7HMMSFzZuE3lxmDrLGOQ1gbRLKUDcCVWCQ/qt8dKw8xqgQ06RoVlRyW1IwmTbd3evUC+rSo
yElOCBLx0L7M+oLmf0oYz2p3UmsHXg0RzZsXpp6C9Tk97LWnablAVMoByPhLPm5ODx3OGszhWKKV
vxPtON/GQwDDzB1glmXlU7LVL0nEbYa6cPHOq1fv/urAKHR1uxo7cwCUlaUibMUxvtWAwdqCscib
QHpEZoqR8DHlpFg6N41y5e4vDAGxWEp/6sF5+m22uOTMmXn2XsptiVB/N/K16kOEhHvE1h3GJKj1
Lxqp8oX/8a9Cdpfhomq2iyn/SoTEfLaQrwCKTY7NQJJTxIX28QBMQM0YbBpOO/XO8y+6G5F6CFj2
gsR8uuWKAFf9tyC1ImlgEYAwQD7x+wJ3yciQaxyu4t2Kt8cxT17EFy20NCoZ3Y0pRXdpVn8UpcS9
B/pf97DkcwucbYFHa5jkGtHHLb1SJLZJXEv9/HGQQYrYRhqFYtFUD/iiqFdAkf7qFBBPvLTFBicb
SPqiKk99ONgPfE/4Qt12YsepPLfFMEI574CZINjBwHn7Sr0kWUA2o0hjK/pBCQDCNzbZO/SfNrro
EdAOjppNpKNKgxB+PdBFvy7SIdmmd/FfOgQz9EaP/9yA0HybXivESlExfhiJtP76yT8CFPfNA7r7
trmdEaSCGa8YsVrwMze6VVsbo5U5lPrJiWlp4GldIli52VdaAEKmcbD/Kf2LKMdThPl7zrtmdrLD
9qGBTpN8AJ8b5p92wb2rDx6LQSMjIMMUA3XmTpLgUNRfpoNYIDrNO29I1kj7rZNErIt7cPhY0yKx
7UaUn/Siu2IpWbPxZHAHW4bc024/iNwJvisdE68qHoSQCEZL5lhsRmmr6zD9bj8jIMLdQsEVip85
kANonfvPdXL9cMCviU5e/1V1thXykAZLlHROvU6L/TpNnPUzYwzpBv7rqTj/UM9m+tEVDCo/xxkt
5pzYAFrJ5DESG2M0ksRME+v3AB4qe64TlB48Ag5Rulci7W7eny9OpwGXGH/Yw/ANujst+Nyyl1jg
lP2xFr3g1+3vUaGgQJQ9wEZMG+N4xsyvmaVpWgWc6FRq9Mbb/zO4Mq8pqxv6Eh013Kt1B3NKzM/U
MrnaigemL7AHD7gq59grUZYcyxSloRK2J4iVP8KUwyTFlXoG2cdI2buYqswdbk5mLxNCMtRY/xYt
0pv1eWKogeIABxvMRFs92bcJ7PNK+d1SRM8s0AESFxcMVec/UCGjFwoh8SAqL0WvIf4FHeeljImL
auGvPJqeeUPP0+MFOOVX/bD2lciG43iB/2g/Ol310v1RyV2VZfSjh2yLpak5N8+BlG0U7aztK4rl
IN3IcmohSBpBSbHUUD6RMoIK+wBU7o8mUu0AY15z9h9O8ymctiuEzIDc5sOhiKjcz+7f7HK5epnJ
/ANuE5Tm7rUZ9Gp3XS8i3FKlF9wGFMXzQtRr6ip8gDijgWi/tJltdaidsAob18frMwCbZ4NHexoQ
p15mKnwAru60H/IDGe7wEIgqC78LG/mX2DcL6aEeT/uFX8mH/j3dsPOd1WGjolfX60G+dQF9bXVd
JEhZTb0qw7asuuqzpryAYCSma3PlcaPxsOP1yx9wmtIKCsxaq98Qbkt4xJgdgJeeUA45wnd/nnt4
Cfz7XxlySXxGaAQtAaHqnl3HQNmg+602z40wuVR5jjMZuuNZL2dR2geZrKXYX1irj6iiI6LHC1+K
/KIL4+iL/0k8WtC8yp1SZnXrLosFwH8S3MlDFpQY8/G2bBPzx2kBpNxDOJJgYtiX3a67lO4hKSnu
s0bD5MOgoSGPcVktbaT5S3k5sbVKhYfh1l8PMOlk3Jg6cWaNyHRpS8j+hZ+IVRxyUC7v7L3akTfP
XcXtN7mBhKXGEXnBzHn4KduET8LNzOUMoTcIBHYv6cbcgvRVbSkPUYBvWAmz3qhxtfufmcxAUhSn
Gb2WHR7Fegb9/MfFGIE9/DT1jz5Kt6+zyePhL7Gr8GyU1/7vw35v1h2U1qsgJ0jvam1qDC9lXNen
zGh2rDoXbmxmP7yKaL4LKPLQZL1Bani7YXW0+6naJ4Ua4A08bl4x1imcBKJ+gkIwZYPKP6Hx0UQo
tlpsmTBnH3tFW3mPf5+M+JJ8k+PkMJIVQqJ5CLLTtS+iug9j9QyoZhefZFw0S3Uo1Ocf+e+6pFpm
3TOPCn49E7pZB6dFv9w+LOQlZi2DFDHmZLDJ0eL+oo5RCk1W/D0H3G/BHdL1ojBqMG2JVWq3FObY
db57Cmc6/418S+fyZPe92I46lc5TvcsqzcGP9Hfd79QJeOiVwh9gqiRBjAm+0+uPueZedbiPMd+s
/bbXEE4N2BBIJ+NRZGcJR/+b1Uynhru87dpmeMLz2ev6RKobPIdZFJgtVcqpxP50F3DontTsRwBo
L11Bml+a50xNgMoXR1xjbkZXxCuiNaqk3fWwTAeGJqvUMPQbWKhgGLxFlFThVjbsIg+q9d9jk0mj
lletjQtEmqmu7O0bbY0OJntU7BkCO+Swv68zOxZy7bFgsmYxA9+w5QBZM/Kg0QCY5Zf0s4FpznBQ
RfngCd5C0Bm6viGx4Rx7KEPhDrWR2wxki+tt87QBnTcEKBYM7oJ6oW8ag3s4awWnURz0Y8Gi89gm
QkubORhb8UFE8InS8MPwB+3rlh7kSkZITlQjttcdMdG17XAzZr6LPqS1I7AAOoJxHuGEHIgLdYmy
FE0BOJ5i3nSlbF1ouhCtmWKleGuUUXaroBZf65N+mvrZ0IeOyid8rFdQVyXsyYK4EXd9QSfKb6yk
gnrWar0JEf/iR8yjPfelNMfkvBN2yHuRCmyUIg7BtIvY/caGpkds7RPHAJkVXSmf2BVkQj4mOyoZ
iJyVCfvy8V11jtJOu8ZBxvasTKXvm5jVL8cG/ERfT7m4b95MFzXruu1Zw/R/xgmDWa5n6QO2tnye
3NyTBvpQjKMznhHQ5w0Dnwp0ZcFjt1Ny95VcG8HZdXZ/+E+mf02GMxY0DfgP18FeSyptzrCskcTq
+7NUkQ5p+yEqQmGsWm4i5Exjee51zKRwEMPSUC0hNg0mcly/qIVRLwzFSWiVFNXAcYZfGj4+VBj8
UhQ+mSr3esv1q7So6WuPBlhIsAnemkWGSnaJQx4dXu7j6HxzxoOVjxD5NHcbL9YprlTmEzCUtxkY
2KvXPogMsGFmi4uxB2bmjzoBjBIX8/VMi1YZRD6nqFZmvhUJxd8ioTzCDBamcLC0C9P0JJZ1rKGs
zPP8Lc9DePaNz1XkCSw0jNUEMyLXus1YCuff5pWALJXrlW/EAAM1nZvS/hUwtOvGRGup/pstyfLX
hp/yPDdefxQk7htsOAGBemYjsNvrMeJN+PxleQgGQ/aeWRnC8nQQk45uvFo5tmQIxomPhFBWFu6R
U1k5ZNHUnWB44e7BCC3QLTqaZs5uJWj+9NYJKqaDuoriKSky1XOeh7lmn6y+oqX8EI4SsKbTa7Ng
B1A5bPU6UCLLlBHZOylu9c9TqfMcLkiUdbn/NVoTywBci/22Z0xO2Agwjn3gDu5CAbOW4zHoE/e7
pvmcAzhYZ5YEHoV1LKZE9hNxb+o4/xpsbeg/QY6EVqWeFuTEeD5kf9rh0zvx1CPrp1k/KLdGBxHH
YZ82SMAK5+LB5C4MWJyGHhxQzcrBa+HtEVUHt4FnatCuNLJ1ftVTuma0+cQfJVyyF4Wc9qCLYJqF
e98rxaFCWb2FxVB93AkJYt+XErja26C43tS25iuz6CkrWUTv+DsLAFbwXzjGFIGRNrwgrHgUpCrb
GiojCiQB5VZp+twuY1eWkAta2uZPph6rtBwYtZpIkmvaEGe6/7KLtuX5miY9VnQo9C13vPg0Eb8Q
eT/WFifraIdQO6vT6wi/maPTOC+Myghlt3DkGxq7R1NTMeJRUX5Mv4rg+LF/gJ/9dnHCD9hfv5hX
NYC9kWQWx+/SnLTXUM2+uUzrwKZ8G0/a3Ulb7LAKgj4v0RHjxlPByRn48x8kCBZnv/3FsD3p6/+R
eG4IgeMVNUzr2hjvgqpaMYx0ynnyalPlJo4SgfeOvFkeNSNPysi0XK9vU50/fuTDhOTuq7tA4uAW
lYoGopSMYG7euOGd8u7jxswiK8/bGj23ITH5GdOqcSlaeXYr+NbW1loP1cCymdwUoatCUHvVHlWy
S9RnoJWKP23spMAqnJQqnYMDfnlSzvZ9DiIIu/DqgZjMxOFS5i2yx/K/dkoECLdh8QmKPVvda96z
q1DmzhxLo2YUQwJhwGgu+jLG3JiKBP/b2BhJzHirLGGVwqJ9+rH9CkvvK5taDpIQxNinwpbxO1Lq
O7cNmf0YKBQEBUrXLfZe8gZTZeTcYKhxUFn80aRAdODSk069QKkPGHQVn1FiBCT7xgHd1Y2UQbi1
HuDG5f8q1Hw+JTWBXNznQ54fIjE4mvWVAiyIhy4z/+zu+01KGVgi7rwLLKuMXzBeCV/KcyTAZiX9
wQn72TkOKt4IUOCYwAOp4lEZZoE8S09NxRhHKls7DT78MXePseZ9TdPc3t++Z1rpBz9TMufgd9pO
Au+qJEe3YIJb9yDXEKvYFoXN3qE2m8QyzLwKxVPFBuyzb6t77nYtTHYcyZFMYeZTncD2Olz8PFtL
6yeeP8C/d/VsSfihvbq8trBAl2AYFSc59wBQnpUi9yYPRc5jwIP+J2B6xS1+qMUA6Sg9tovfUOUB
QiibcNxUk0rqdmCN9rLcQtX16ndOLLDo6Ei8CwQ/G2Qhrmum+oR6wbAAnJMyeZdm4IjKSiYu0teS
WWySvHFmHkbqTib1S2YLQ6wdfc/NPboMnUDQIonjlW3BMoBA8KL8dJt9cAlkvpYhxMcB88Gh5ZV3
r/iVInt5mqPeSnMxVGe/+Aj4yGru4l2BoVJAf+njXa08OI7dcLKViWFSszGhmw4LUBwhGR8VJUAW
yXsd8pMs93s3smQjN/lmTLiwhnIgxtWZ/tthEJmJiQ4W4MD+m8PefHbYjcjYDruaMNpiLnTy+K+I
4Noyd8il4dbOCeImbHNmePTMWI26cMCXvgpxHfdBRkg4c6C/56T4plc8n3ArjqVcaPS76efXoVmz
ITy7V2sLYfj+FODjtMvm+PPm++1vai+B/YFV5CmAbLAuFJwI1TFbFtnIyoix50y4cXTPn/3kL82r
msPMiT4PV54hBnXwgPyTiNpQpfMMZWAwOxB8cPdnHlG2HhP6zZdwBE2plTydg1VPEq0tZYs4PEZt
Q3f4wJ72dN1xTxcmGykoRMgJ9hXGmlvfgllKvOSxNk+wW4uyFL1FCflcV1Dt/7b6ce9XaUbGwmYM
wvgkgSeWqgNPEJLtx3UM7VKT5hy5McG4AnHpuN3clzxtRUmwZ/Hrh9mzlA50DtAfk7ziiBqnOkc8
hS3IhQc1cvbbAKBj5SJCDoiKnUZ5jf6EI+8er4QRjaHSVr0heiDcTg9APekxhEl4PjTbw0kuFl+x
RyeseGyt9hIR0Ppri1gsZ072PpoHB8vxOg2l0IN615Jf/2ujpi8laa+1T0ISXrgEHQetN8pK0wIb
8aZlEJJM7UGZW2cUnezkroFEiJ11d/IawdYonaVn82VxCs4MakJc8D1Nog4q8IJOXjkb0uK6mR9w
fjDR5FmFlTtX+5Lr4VQxwi2J9u2PrTczm30rPcYRkBz1lSZf19U12Mv5VkWG5O/cXCE79uujZ+Ln
OMJ4XZYT2TxkuqR+oAAl1WFOxSexTRGEQ2gamTFNqV+JiJr5rRkL44oEbGHzJT75USo6+FBR+ovD
3Mm+5AwmCNjL1q6GADhdyCWfm+kfxXJtEMy68d/YIlifK5twyYuEbEQdaZM97O8emd129Q+paOdp
c6tSe8jypK1L1Eycy7A9YubDzY1kmgbQF315QCXmFo7yDfZGGMiA4NJ1Db79gzi47hCpXn5xwU2Q
jyGjH7KG+ZfsPHVru9/23dzcVYFOqmOmcZwMowyfMTa8kUj/hKU0kFdq4Y4dfxIxBansTtm9up9u
VzQeYWHx24BYR4q/BS6sX/d2+sYqiVu1Doi3LWReLSVOTjcf7yx814l1rXoBr4Frz5BtF7savoZe
xPwONmebWsj0osxgFWurAt3hsD7/kBkSNfrTCHqTFdfMcUJsRQMdPhDGiGSeMmtqsr3WT/2SfA2C
IZTNaUVxLDWd2USGS0bzCV9FTx4n2DNOiM84b6it/B9njnVgxh60sRPZbLkxpICK4y5OfqnJVYtW
jKz0M9v0dQZros1uOVCqI3K5p6y7j9QUiQPCJsMqRxH336egaZLe057pE7jdWMvSf417O7P3I/Rx
AtbPj7BApseQjK1AK5mrIsQ7Rah1MYx67SIA4tXEAxKvPZ+N84K3gUWaaUWE+oE/xL2QQRreyq29
6n6FHXBTrtinSpb2ekMmsOaepeZxzXJ/4YxMj/dbLanwEp9Cyha/J+PcMO36nE2TQYZ5J5cj31++
MP/fqDfh0tVpfZxwUookdOfJ5xByIsCc22c4j09VD06OaBEEX8ZV/ZUouM/ISxcF4hVHuekMikKR
EhLXXmokyHdvcbeWsYTrdOcx8C/Sb5aQI/sTyB3JEAwzMNjRzRsThbQ8PVVTL/qqJ6Jd1Pa8LoVV
H7NNtjTP18hO09tCAfAC11ZH5uN2GE9t7urp9bx21aa1cjrV6MV6TJ0rIyhL4+lw2YNX/rI8vx4R
e6NhS78CvKGftDPhYDm7QDShZl70qT+neKwZD6JsVzpJNIzNX5lTJGoZoSnZDV1yagG2coLEK6m1
h1jrWZse6Vdzt74dAcfI1z+rs8NuZIQtN599vUvGBGElmeFpfB3Pg0lOItdeSjFQ/ERaFJEAFawk
tdYcvm40tQtpbsuOXdidEHwEkJBN45+RGCa3Ll4ffz6kBL5Ek6DKrYlRd6PWepyLq2Ou9jtUvjfC
hcjgmizb/gH1FuvznCyoluIVdaeV6nAiOuL69P5wIQMTfXXpnh1wmBg8dY6IxD2ulz8JoD4LAP8+
OMI8hQoVmNuiLBoovwQx9QWdgSR9ZwCq+2bE/uyjymEHt1NrvWa5O04ErHIWpL7FkjUf5qHeBHfb
7nJOptaPN2OKdPZZyzxqw5Xj5O/UH4gDroHLBgTsdIWbA41Kf38droE9XMARwAfwUsedp66FcBM7
jQKxkTrOvFWkfnqKw02ULblQlF7d6Av0bhnlPpHhcFSOCObtZNjTP1GznslvxwmAaPI1YuA+l/XP
1uEIuh/LvPa6WbWBlMVJ+T21/dxz4hI0nitirUsjXMpnazK43jUjf7O0djCQ/KainZjXXiOrkBqW
r346vgetzgSWt8XAkjGlsrmUJT1tvoTG2hYkEE+S4lkECIQSRBQvaI4nzv/S1gEEWhZVkFnrM0x0
sDetI043Dy6tqIWkfy7LBGVvcXI0ncBDYwQbEyrib90UL+D4UEPQ4T8Ny6/QV0j4fRjwXO5KoGbF
g+qDoJTSmxXZGDBWNadnGeeoyBFXyn0TNKXWPljn+07I0qzeMKIy9PP+p3QnAn6ZagvngqfeUT3M
4UM1IQF518QAGcbbMlS+u8ig8hdvbnRhysXJr4dHBL9NMfirwqlrFRZY1BZDl458FaJuf3ZjeREp
/2lCr99vlhvH2RB+31z83/0jVjNKdEe0T1w7AtSlizxWsPyV9EHr+mNlGMhd0fAaaX5b9nVZp2zs
+tuHi/gDpqlUawyfI9Lok42Irsb0lcaKzE2FLN9TTFWtzkNPueObmisv2dOo1WtLN+Dgdegd/5g1
xzyTJ6Vr1c3JsTsFKasRGfX9K/L9BpSZ9HFfzpF3uJKZyF48PWp5TfumIK1f6Lr8kVxjo7uNRuLe
I7cHrjXTlMyU03hCVXyr9tWcI8kZanRxXGGPEpbg/qtZF00l5SDSzvGfFc93+x8esgurnslsyo8G
v4mlePajvdeciNfudsD0PYE/ez8kO0W6yucVsFac2umXAiSZZCH3uhP/YxpVPlYb6xh7T4bC0RsZ
1v2mXZvao2OpzSUhua4LcxzWAnVQjf/AAS+HXM/2rUFZrIqlBSbQZoUwQuirCJbgOOTihU3uuBA2
lEUumbPCxs/PL90+jv5+iBzRpFrGOrexaa0c91NuSrjDA0/9hgD0kjKh23NpgtilIaDk+Lmq1etq
G2WYXPDFpYD/DUSTnPA2/2QlW5DsT0YRV5WZM7ckIW4mA/uP9ChQZtUdja7nJPXRmC3L8WXuqvv5
ZI6tJSZGiUcceBDrObsDU1GQac5kCMR2jtKLk2pSR/nwIexluCDlldQvQUGHy2ue6Dqll+AVKlq/
GuhyXXtvlqd4b2koudEyIZml72Z+cJ8boQ+5bOulb11JZgKZrfzINZ6KbFESlguukuvTMN7Q7av6
UeONqBlsz4hvwWnMj4OeyFHlN0kCZEhshq0ZYGqEuNGND8LLM0gJjNf3AARSpgjDMxxwTIMKoGtd
ne98KUX6rx5H5ZgNzTL+RCLm4+Qy+Cycp2wFVRfU/+6wW5JXEKkigI3bxN2ye8Uq1I6gcu29jRlc
b57gSGc//pp1SAdXahn1E6RM+WML4fsMKZjcz5MGxiO19ZumjBt2PKIJHysYDq0MsK3O0VLpvbzN
tviMsPi2FtiAkqgbnQ8tD0b2KwTjj4v12EF6C/0QTKqWeyBwt6kqCBt8Z0dw17m/dQxmfPAzESNh
d/RSnT5ZfjSWlQjDJIEAO+Prhn+NbHgSZZw3dSXG3YXZ7qIHYdeEvo4bYO23fT6JluvSE5JCXk2q
2V+COxswN0CPGItnBCqlZ/d5uWgvk/jLeMIjbv8vdOtzuul2RQAP8L+bBXLHMaNkBTSv8hQkSH1c
md4V59h9I6HRoib/rIMSDQG5LV6s1pQmPHZYooJazVYgc8J+YHOaS+ttOD2A872swFapcj5SKUyb
u4dXI8OXq0zFl02gNwsKDwjq4T+ZB5k1d2if8gLdnrhlhYXWE4DkEVFhcBTVuLgHUL1BMvkNPbEF
6bqBAiOmTRvY01hyyipHxm/Ne0+iJ5BH1TMLJegCjqvhiRQ+vqqDnGawFzZgnf5uX0M6YtWEASR6
i4gz34FJroVTNxFn6uWVpr8/AJaKf/ToWtUybkwH3q1wB4jjElcOHxDejuZw1daYbTxtu7sI2taq
xl+glTW1tCYMppjhgEMOJfEgBhq7kYjstf13dzCdlAVYNI6Y4KtFAvKgQ8vDzpWkrDVWX9w9HGCq
2G5gzwh0vwdQOET0GbxpjJOvMpF+HDihRhU6HzTOPR4uyvxRUIDML60HpMOpoZmttcro+X0cTqJH
mi+JY0w+j8l/Q9vTNpMHzHJuun/+Nv1KAO3T/uCCEyBdnknxED00XzKC405YCWcy6i81qntEv1Vl
3vNkwrLm1nMi9zFF20jVKbp2Ej81yST43zS9a5R8QTyQuYM9oHaoD4Ep6w54/Fu6o1LzaZPWDO7N
utTUwFHfz2OyCx8JJ7y5ZTjw6yvwZioE/QcZkXXRAeFBWCUdmA45LLD83Q8ewebPyAIUMrKgC1v9
Zg/mzOZkzaPDjy/9TiC9V01TSJ9zCI8ePHyR/vwi+xDSR8uarVI32GvpnjrYHeEdGza13WQoQ4L3
spv6zmo38VRK6TmkciFREvnXkbRc+UPMZeukqLVTzabv9BSuNcM2R99sniMq7D7KiJ331c96ATLv
Kd5w6K8zlQQINLbzXJYs1gNubcKeuJpvQU5ol4Rk6G7NmlNZEhG5trs+lJKYiUHMtta4gkh+eKmT
QkKupICkOtcO2ifyjKPD3Ey66VMcBv50wIqTQLxDwHidi+KYbMCPXEzcaJKya/01mf4q8mxQj0kv
KJK2nXtMebMIxTt1APYD3mmTRJq89aNNSWe4h4ts/YpYf9Wnw8GO010CcQx6/YIF2s1GCahRs5sW
L5DfVxdk6oTeS8+xi1l/Wif64zThu8Cn+kTp7N2gAqNxZ9eC0hj1g7F+vLNllIVi4mjLJi/YttvE
zN4LHWCFbx5C8eniVG1PoiwX80Hwh+2coPoIRbPelACKjE4yrShctNByMdIBQ6QmlpzYwIj8DKo2
OwQu+v+Lsxh2MhBVbQ/Yqa+ZxtpaiXEfXB6GTMfcIyhAQpGg7WlaCSOE7iwLX9sMD00a3oeTnICT
CbV3p7mk2/Rd3wL4UpxCb7NhkKQ3itcZhFkL2oX4FrrW/TKB1rtZdQO4ukzSHO/ly+5H0QN1rF0D
EDxg1D+UTQiBeNRjN9X/FqV3k0cCAbjW75q7bvJcCsKP3GKKgJQewz3Du1kpcX3BbiwywjHl65rN
beM0r6YzjK3LCMib/NyzXnKolAbQABg/QWfRNhjOIePsfGDKcEzBX8zw1q6MtEV0dhqroyAqRsAu
ZiZQzQPHyjaxsB0VxU2UPEGcAwQnyk8R/kJa1escc+fDJRQM4U71obIbPwIru4yD96P5nTQI4sNY
hXcKLLECWxv562REDCvI2ame3dBwmzgOdtut65PwsFsyYgKOfCj+zOwNa0k8jVmsCg+01JS/le4q
H6c0Z5z+7qXpRCEypQ6VqCCZb0YHfKdg4BxfSPieI0QAJnjvkMZfJwVCVSZiwOAYR4gdrB5ZSsYK
PFgaYVjUgMKg0HjEmVTwyKAWT7Uk5X2yFtPn4ZheHfEbZob/mQIZppcMqoVGcWMRf+hooiiiYqTl
HBFeBl4MBy/tQMEmqdcGg+ZvnrI+wjGCvlDk03gTFM6WCwMGpv+Hc65T1w2paTit6Bs2H0XSASOC
ikHpy6NnZHkgnE/HPfSyh1FtSoGB3KfRtWMGKgHMkdtDZOvY7E8aPrXh3gU8HkH51VmU+Brk1wSf
FY1r2p6mNVpR1wqi5Qd/5dKlAR+005YK8rf0a4j8eaQlYORCUBEA9DbAWZ07oGbTVB8fupWlWtuO
k0K4fIrF3eftn0rE9+CUFFrMELAt7CfNInBS2wAch/jKszaYa4okqQtzpBWXtmbbHuKfhgLNW6Bu
J4pUaV1Qpnz77aF3UMWjaZ2w3tLw0CKdoBsPsWUxEgGPPMAIpCL2BZYKufT5aIubLVxaYxoxBP9u
VvK7fMW/xKZ7MdrU+YMnAlnhkZmLu1nG0VC3vqiPhx1G7b1TNwSAMlmArUnFF9iI8Vlge3HU5EoO
NxEtFl7THqGFGYNc++ctSVFv4MqcgK8HFrSMkokG+PUrYfVZPcUJsHxjdNTPC9BHc/5V2WpDB8R9
yKPQhJ5x3sPqumWnlO8/z4XhTF2wjYAP6b0kKVlK81+N8zZlJn8ixkIqNbi+C9nLL/CEFl2dumf0
CxhsjN5B24FDQb4qGtKI9QMVFedfbJxy562/LprIDVcvQrwUWKvC0sHRYBw6+mBR8F9Nh5YmJO3P
rgYc6idc0CmDlG1OVkdEdXvJZVB7M1+4pHPwK1fPI2vdjeL5dl29NCCX9H3ryM5AUZU3+SBvIvin
61lio4ZROiajD7uelfI6IUpaqYJMob4uutTlDgVTsKjzaiyI+5ozT3YmjrioAwatFj8w71jAK/IO
4SL3botW+aREvKO9KokAK606KXrCrpEgGOwOG+f9Z+bv+lWp6nnLzLvVtZNJa5E3zrfyx/vCR9Hn
AuDmBPFwINjRM62rOjK7XWV0AVqJmhFmZT7lprmq+cbiYR29YY6BNL4r5QdlUSCjmlWpVkUKCaFv
CpqJx5dQIERUcLaJ5OTqmIBmMQt2GOzgH+yMH5ZNfGqMvMJHwxNnN4cE71rIQGXBwCoAQAqVWq7I
WuBv5A+4S7uSOhtfow64+QiwZhGTTSQI3mrzrYZJauD+QLs/hp2EMluf7Blwf1BFY1m94RcB1tva
sSkY7vIfhzJ38aZN1fUwO7DXbJvbajg1NyCTULg0E4xB6QbVJOERoNfzgMP/lfdqYhBoMaVXr5ar
oPD8XRcWy4XhdeVpHBUbALJLv/oyq4Db5UUI+gXaEHC2icGDPJPJIcX8Os7sUqs1GMW37wZ8MP6r
BylPHlX3SqyfBKgC5dNhu/O3dtmUxrAV3sVTE8bOxEX7SgUuZ3V/5B2mTSlBHQ1UfhCwyQ0ouo8k
/Z1WecheVg6+hxj/4ARR86oVgG13ifDzEsRihKJalnzzQiLRWjyn5QyCgmwL0vf4XclsETLpCKYV
JV0VcmdV7isjOO9VnQ6bHseiGdkhHA8qj19mCl/UE1YQIyB2DxrdAgJ8IslcCiLBpm8QcYIVmxX4
1f2df8gtwEkt13yxIGiFaFzakFXZlPuLewSy/80H1XQV/pZ/JlHE4mhAepzPb3cbuGV6ysStdYCO
aynKpsGaRvx/F2gIEuyCpJZkE5EeanEr6lrQxDIEunbvOe2jb+qiBh3U/j3k5BReuEmSap1jbhuE
fa9aDtBUVLsHqJWPS1dRKIIm//bxZGKfLqSa5PLk5jxJP4Glpz1By7YybCetV1+ATB4szv21ZvB7
Rxo7eVowi+8+DyQyH6DBj01aYD/uhruUKKCOGfFla6uTUy9RlwLJLgeWBvwtseSlbyC1fKd727QB
hGHjzABhkOT9iq9D/LP6Rf7Kg6VXyIW1WreSTZ7BwTq9R6BPUY2XmARCwx//Vr9gnA5Q5/nZxzV5
UaLkDAAd/Wy0ipUwB2PZ+YypS5uzbt8Z1lchVJvXF5JMBeOfAysDUOChznd3tiFoVyUmwVZppAWU
ioxoxpVcJ4qBmpWkYplbII9ip/ir1TEN36rO/WxKu1OmiP0xl2h7zpfwc+CuI6QRoyoq6D5wfAmQ
UiVj9x1UTZic5OoJuUEt85pt2k7+WDqsxtsQu/MkZUIbBc/XK3lFKHlL58nHeC9D/Cg0neZd2M3t
XfSaWFPWAOztMCwr4rFY2zuM0f9MKYNoVz8ZpAbgoqzXvXOf+tfQacyaOVC0NjKiKm27y4InsXYc
Is4hoYdndGgPltb8zrI7xgsBA4GKp/b4p4KFaDOT/lViWZu9KEc+HauQ3PUrOgIHUKDGKQ3wijww
hvb8dl7xeiB6azw5bD2qMOF+34Qfw24a8PBuL2myYfYJlQq/+fj5ihBqywzpHgEDphJeE2pDEimX
Dyyk603jGFdaQl7Gz5p6xOK+4qN9GHu5soFLcSLjn818rjYy0IBYlGwKjAWWnjmcDUbtqMHDhR1O
SILlIMhNcpeKt0+QiFZQp6Pj3GDOb2Pln66Vao8UYKyQl2LEPM98trp1szOKYaFob0Jna94SKrr5
sehDRBD1FcRwA46tUqeOrrcGx0ceGgipt+iqieQaaNjhNi81SPGuJTkWrE1ZVxO3fBAioQg8Q9z4
EQ7JjQJ6CRE0rP7RERAL4hKvv44OJPOA0AzxgFvQg3EqRPJVyaPfVrAjFJ7vItg8VFRJ2Z4aLCnP
7FtxsQag9Ni+68v6YN2GjmSC3+WAhm/vm7/FJxlxgJaZAmKuqNqtrVocu9NOe3d98dSMW2i4qeRZ
JTwrqfb6ppW77V9brkLCfi0IYfb0wZMRXFfk9ia4DyvBvx5gAulH1j6sPAPudlzgQAs8RyvsTrsK
UpJJmtYelmHhrUsly1pnoIAJ9EnhRIFGZSn4Q2hblS4kOR33aZs6yQ/Lt/XkonfxDlkJBvw77uZR
l9nMPbS8saJs2Wf6bS6jdx/YUL1AeMKGCGabwD9skQMmXOR/uZyWy4zu2qqpTVRbed0fUPQLKEiq
4V2F84UBw4ixUiQmzpfVakY6A5Ee1Ugj9IWd9aYh/a+je7Iztp9jfg7C1TC2Dc5Uz5xS8OAHWzLc
C0NS4Ac2eILmGIbLfp37RFBxcHAHfORVV8rXvE8UI7N6+l7Ca3Iqx9Kj7a+W7vGS64SWWz4iQEie
e4aRWnvMS6RQ64J2SDsbzQgwUjRz4mel8rslbTSKauqqowjV9d4QgIpjlc4uXRkKzcC4o8uFGKjU
FGfHXj/Ijt4pPMzWE2mJaI836hkLwIcrrOny0D2Nw/qY/hNLzXI++ZnsTeJ1k34g5Lc2WbTl9zGN
xAloubWUP0UNW58L43hHcDRMGjsjZDQh6SdOwe2XxgqUYrBuw40nGnWc9BCPLvtKFtrDVTwrZYG4
mBW480BwYuEPPsH81JV+BC3w6ELo2A0A/aGfZf24gQMnLlgkqsjw5MoyEZ9gAYcqB1cyZw1PfHv6
emR/yqAovPfGpAWxLc47gF10XG8gLO81dl7WldluF5bgZL0Z/dUoKPRZ50JY/Oh+Zl0ukQDFwN54
DdjN6MMM/+sxT++BfiqngUceKik+LD2YuvqVmhpJSUrMv6Hwt1ao9YAiZYipYXfKsf0pdqlPk5ok
vPpInfC/PpBxSoA9JFAe4ufmbd0RnOT4tywnKNCwC08L5z2mEHBV3E582HY0+binUnxaoylZADfT
QzksM2rTB107qlcrRHlBrXJMIb0xPeR13ZzKC2YPmATEYVt2sBeb7BJjwQsEi2eh5Fdj0wmcKmZo
619cJaj2fXFwF1U5/7qaHInZ1mcyL7P5GpmPh3Y0AyqrUS7nVaCNJr3V0/Phu5KN8X3aArEmDXdp
a8TobLfW3WcUINl7oFpmUFFm98W4UvHN7l+28zpqCTOPRvLmOk1rJ4QaOD6E29eR6+kOCj47qVH3
zFItlIxNPJIkZUVLV68ZbQn6vlWFM3Ut+wM02Qg/tzT1fE7O8uTL2MHJtU+wj6iMi2eQXB8GxUMa
ShPvkYQNUy29ICDxEu/q/EeTIQx49tvBzV+soPYcNSaRmp9sDrwfZPWcdyRJBx2S51RdavL1WB5d
I1UCIaR3wh+HQN0eCp75QVQ7mPqH4N6zAHAsahk4Kl9Nq5WpICCK/Apag2jqbClbscVbA5yN3Qy6
rfQlvBUczXR9DUycHp9AywU6UJDT4G5JST3X8UuyKvSruV1e1WGdYq1hxZaJaXfRoufdo+wM5vit
7Neduql+PuSedhvmIeTwszaKw56cwKujjGeScCQmHs/WTQE3W3gfkwCVy3tCq/tbvVqPEkuKMTJk
HoLaGOZQAQmSerc7HXuX4wL9TasliBDLcXSDABzSVEsINV3C1x+m/lvi6eSkA1I/G9azYBsbjpvr
FWnfpvuoT0kqkY5ofMP5n9uh+s+zmePo+z5aLu1ppVq918p2yJDCcVWEgaj5PJQQU7+Ox0yMl5jB
9rgBNLBXqDyrpsy7IxX/3K4fM3XVOetYu5leXuboHJuI6eukr7TC9E4E6fjurtCMv+zFl7O7psK0
jE8qkMF0XMLTF3ybovgoaA5P90llaUL9XFcuo05qiqdQNF5tZ1JNLZj1eZadAg5xvmrc1gJ67M2w
3Cy/LqzDJID7eSw/lC0x/UO2mSC13g11ilQTf1h8Vbn4b6KB/IzklCszEKuJ8uvWr8erv1mJUWX9
NenWWD04ja+nwM/jOQqN0elfATTa9YNBnQYlBBqKR7ImK7MiGOa4OHG60CBmiUW4aejoI+F8RZ5r
wn179tQJqLhsdhbpeIB5ZT1+0gsoEjCGXj53lZczLWTe8jLD/IbDtCfz3+d9qOwdtfQwvxHYpn5Z
S1EIc0h0iCpqZjKPsxSmnoggSPwnQCaE6oIdsHIwbZfrC4xbfS1a8+AEibtiMICssL9m1NJVN/Vk
xObJur/o61NoURvPTkPhpDAu+EasSiTxNLcTCoi8+ENoIuAeb6JfVk8gzPz0KFgPoA8rdGUjad9a
U6qQK1dPNU3oRJELD890EO0ot5SZ4pCkRfoPy1DBzlogudgluvZami3c63nKFHbO8PEEqVL0xzrK
yV75yD4GtjTfnIX6qKZ9RNX5vRow6s35LC4pTxFYIS7R9Oc+FHnngPDHEFfVVVEgUuNPb6hkpe4g
/l9WoLRwnM2FfJ9xrc8oxOpBJNQO1VmcmhTgkslDJ6DNzQS+gzkuIVrQzc0OG02sVNszmBwzaxHH
JKYpzcGOKeRxM50gjPNPHEmleHG+dU0eKm40lhIvI5LCSssivWdM7RZ74y2QLA2Dr6nAgW91YzgM
9n6o/d3jx4MuRiRm1pGiLQpNgTvCuWAnoguRHwbarl8AxqgLU9yXPkNPe8FxH4UNqN18YnqwrLw9
07tB++yA1jrXiWbe3FuEWE3v7CPWucmrq8h682/+mredxt/+Y2G5QrHinoWyWPFr3GW7dfOFCWaH
GNiUCo4DUlS/AeDoqy0CiJL9vlthArZlrJS69n/sUrlSS93mn6gwDVU1BPdrFLiwYRsUdQTVsBux
E8DAAE/cwD792Tznnr45356ij7OlSCxyDCTzwE3zAh3uGpzzMdfOWwkd+GZ7JhHn5rTxpPpjVG8D
P+wUhbGacARu/S5jHNIcnA5kaLd74sHJw3Q5XBrf61wOZpHXd31a4GNH+bQ0Lgubft7QaWZFHkb7
3FYDVRi5OEb34G35okoZaRKGz2RmK4j968L7td34QQQIfZzv6jQ7UvoreiPIZPCFkwwjWmR4h4C7
xO429okE0COEDdorlhncESeXcgMPk/gaBMVM6BL/tjWS6gtHInO2HwmHKUKyKpX7r6dI2JVLOyjd
UGrp1wjxuiITrbqOqq5QNzeHqU7X1GxUgch0j5PmboDg8KtMDKYzty+RaE0pjwOLFfhQlwuoz+4T
rNhU8vMT3IQqn+/jv5pHwn/JqD38HoE6XP2xMz8Nh64ISveiFzbcGipIiTV/o5p6LwUlPbSFunWP
GLVCFT4Wt5c1I0uh6dc6Yb66XmIUkyefWZHfbTDbwwYpF71PMqzrElMnYwTQ54TbEHjjdQcOPbHg
5y8O5cRSkgP7PC6emh6DWjyvab7FGHHH0An40nPOMZTwLxc9hBD7H6DMGDc+equGzSMkRKeg8GAm
1ph7r96AeL17f4FR56RL8AXxfG86JDP7psysRDDnouIwMpxZb5ABihSGU4BvoWmbcf/M2HZdXaCE
zT4qhYKFMJInWsXt8zOwnQEPACrhaZgGIe5hDNrr/+aj2aZi6+c1uGxho7nZXYNW/bv8FarD7Qyf
DpTJ0Dikt9tXLGJ2ZVvs1BUC3IdrfyVeBKzQvmgcPApcSm0+khOjKp09fzdnx0Zqp6VqIayyzcc5
x98IAjbrcwIkL/m/CjbJ4za8JAVtMd099Nvlto+Fd0DB0Y1vmI4D3yoYGfi/FP7EEMVo8HoFamTT
epxTZ5K7vYTp1Zsiae16VorbLBJhIUYZx/qZyggOtmv7Ggg9v1ofUIZ9jNxTtgqT4/UcMgLKKFG7
cflUjLqiokk6pcpKRfpQR1hcq0mNjvHvNlUfbbdBzDbTjU+0i7plKMQ3mbJnGqt+5aqh64n06wzp
lAkr1LhZkB85bod30Ga4Gc1CiMvPpU1n+Fq8cHy05iyyOAt4FSaYrk9D75ArZqQfXvvhRLk9HQsT
rknHgLWo6oqdGLfdnwttWu2qhJGXY26KwKOyFTtLeOPUB/+9d93PYJ4MEIfmpOAEvUloPaR/dmm0
2yjZWktWzEYNXaVn+1ma1+/CZI1HzyndsSMa1JhhzKTs9VKN9hRmIfFDAOvl9PjsepTf/K79xKg6
Bt49UVoTwXyuvXZtMeMRcCu06czm/A3d5VnkBEvwPq+YurXeAzseESTJBBGktfGsWaknh/lKEtCr
wg6bgj6kn1pUbT5F3AJbkEqAnn9P/bOmOwLNLG+kVQOAhMcTWC2Qu028BFkt5QCx3d9wV9kbNc+g
hCrAQIvd/OVHws/bK1SMndYPnNQir0WP7at5viIgjInymJDFck+UJA25EG6Jw14TStRZQfTR6KnW
R+/IQpeqMeZ/KI+W7Y5iIl1DeLc9C7Ild51x022XyVw/9cQIusNNqthTf6IzAgMuu6ZMA1LH9w0h
dz1jb7R/h+LH0NQhK/h0rE0aPhoLKt9v7FAaFBW6WgQGRbCXgJ0kkKiwzapKiPwSfjcng5oIgwik
uy1OQxiX0EZz5MJKVDXGxRyROCkWR8skSPPFJAWGyRlmF42GPxCpdcpRpKqa9tBvjcYQTqDclfED
YPGx8uAQQ+61sPsw6NzMND/0CDHU7aZiKYu/aEOmz7vIw79G7s85yvmTHu6MqZK4mjamU/tsXsmT
oDeku0G1Zmv33/dbJtSTUvMX3GOP+mRhJd7AkHNIhL5l840Us2NUNLhuIb9g3OUeOr+n4c66DOd9
XFq6jYU9GSEy9CMnoeyaD6dLzA/jN5B0JASC1NcB/znwOOl9ImHqMVFxSZFVg28xZRG1RVPmUcW7
vjkZ+3mGTnleEvc8/hKBKhnDzdBu65GgM6REoi9bGSlhz8/VvbQZ17AX6i4NYDJqB88y9lv9yXjY
4n3XMIGG8nG5M0RAfLhePK0anZXsTqKd9KhgPe1hmPsbj49Xe78aE5TtjDvxb94qr4d1JVq2Errx
tXlAHL0BWXxppUaIqlzsHRxeQeAhnoaoEeFMvdi3p01xMXWWWiY2yRKdMpivs4/xHt1y89nAH4iG
zanoi18ucH+Nf+QI68NmStYKUomezUGuwMaoJLe3jUtnRNKzth0H5Xb6IT2w1wKoyRChSvvLeBcU
4m4goKb8rw3mJNpBgxbeDo1X6TkWKXsmSksKO3JPqeHSqvhzo6yJyGB/i2hTqyXNSvNXK/VIelLE
IwbwuNy4dhYj82PjDMOTBjCqAiejkwj/hDAaQdgou1ArwcSfCyJEbWoZZPN9yemu7RK0F0LBBTN9
5rAhenLh8ZS9SEYizj1xc6tnaLJPMYEQTFMUY2njUCEh2zFGe/OuHuoyFwryWMq+E/tG7hJDxZAQ
fjrmgL7ybKpPDPmP2ogQc0Al6n6jen9THGfRMFwD9gxvyTFhlo0RjmM6NWHRh1qN6gTYxWpVEiY9
I4MfxTM00OnUZJHsu2ZOou3hJBlW7C1CKfc7XQA29TiVOThARJH2ghYJNpwwXWfFKSXEeCNpIDPZ
SsuSVO+if+ucrbrrRG+AvMzA5gckxvtRUCRA4aBq4g3tdAlXpDskC4KsEt3PMttzymepGobBdzGh
pejJwma6idgX6Rv8z7r1QnnCQ9Ra7XNfavtWErgsoEZX02O3a9cyUNlSKbwa5a/kcs2s/EkydMsr
kvYnBqOoapx8KG1uGtAPL5SscyMBeJ2EPb/YoYJiwjCx8WkcaOUFjmi8r/sXcZMMgKRkX5yGWDTH
aQL6vlGiYsbDGvoqfukyRj5Xs3L166Kdb3dTCzNcD/1oF/pUVYau3oGhSHdjfSEmy/ijRFSZJF4H
ZrD2i95HoaPEsAsNopn8KGwAEs460xmMUB+12p1ABvVbF/9G/6cqkuP0zTBdOJNwU134MSCrPurG
QFAwLCDQUaJWxGoVS9NYCrF+r1ruhUBZWwFNENbecRc82/3c4sAYyLYc2qurfykn7CEo/cugpGgv
ThS+2Sm4jiR/1vqGdSIIVwRMKFrdPonQ4mYxvRlTobjVDVEvR1w0KrClkX8L8tTpzfwdr9y2yUx7
1cZxzuAhH+kwXmhCOaCm9h4uY84CfGii/YH1CchGH0mZ3tmKaAdYs9IRzyydx6/pjrriSo9Q6zmr
Yr74tqv1wtTp/4TpDUiwmiAoRkjUK5iw7YGKLoYVF7JZLuaSm5ae+Dq92HopvHaWaqeeLU3U6Pl2
/jcXu3Anl/PQvfn/rbaVGJlF/nGq5bxanGlwq0wAcZ0NhH7l/uWuofNjFHw575xKAoalZG+ogmUV
uiu1SAkEUN8s4IaPkA48zJkoZaySYwGfqr8Vou3ZVx8BJTOCrIXFSFtAKpr7MSGo4lijU+9mM7JX
2S/pH3bSv1JdrUJ9NCMX6sfLJhqXtYlI2OVpnTnvk73IXudR7o7MYNjnBvzw7Fxk3Iw7791T164N
dwUQ+57qRD6Jj3R1B2QWOLDqCvTgy+FsBnSSm4fK9EZw/sOusQhHdrVLpq/+hrLq3U213CZ1y2lF
UrDqq0b8RMYrJsl6V2F5MtYkanafaIdvDnUR7C1bFILirBjj6IQxFq4yYsNoDInfP03UxlwiejWW
cuIqgRLLtXbreEY1fW+Snebx6ntI2WPBl/pmfUPxiJK49FtULipOLiktz/Dxp2a5wVnNVwW0RAJg
H8b6dIT0MRZGr9my5bBVCt1a1+vRjnW0WbbmN+CyRJmrQUDm3J/L8o5wk8Fqpohh/D2ZLU8hC8XS
KoxARNGUR6Woo/PXNDobvLR1PNYhHvHvAjobB9NFbpsoLNIyHL4kUzlKHKH13aUQXp8iR0USqulg
fMpN8eYkMUL10T9Pead449RxNgBHEn+Z+/4BLiBg78B6pkBLfCOgJTHVvQcdjaZmpcCt+nBR2brm
tbgkvT3YIDhhqflgvVlVeMZRSFR515Gzde81d5mmd8bPDMT8R1Q8MpAQa/kOiasgFeKoaxkEABRv
J40e5Xx1kCey+O8aWPYfwmowfPDtGrr4wYqnGSu9z6MOJftxpKmmn3MGRFk5H0FiRmoLDppQmZhx
B+yimcgb92YN7jUdHpHZyy1zuedYa2mfV/8aL1V8TDYF5V3e/x02+kLVCa2Q3VIztVCfI3poGSxF
dHrcmBbbuUbWO0Nr6bcCJ78cj6qOVEulUbVzNQ7b3+ycRLevZTikt4j+4y0ls+1RNFMaNz3nBYdN
eRAcZqJXojT24EPJDX3wB6q/HWx+Wf5NSDkZMG+LbAjDgjlYQopeu+u6UjjET9dw6BrBVsIziins
djTmfDaLQhFo1sFK6UchKPGV/Tju/G4ReT7Icn8J/jPG7hpECQ6/3FB35M/YpR2+h4fL5Kx8X/ZX
xq3nD9CLU0gdIGOdcvZV9VLxTbhSTDSdghGxrcSHJEEkrQFMkgvClUFFwK+KyFoUFDMtAbjyHafe
feqcIBxxkuyjom6RnoKHcfx9zSJf+q04DG+VRidNbTLBR0cIcU0GCrjwbLqq0J/2e0ZQdaBo5U7k
MDij+PrMw/vhQQm2y4Ubv1s8NS3rB9UlCsILlnW9KmbvAehg77N014wWWmWLEsr3N25bHSi7bRbk
PK4l9t7KXrBPCjXDXfuPdUu41LHKlM9FPpl7KWV2dEuJLGCP/K3ARDYbHszRVqOaaEzZW22D+Veo
Xwz3V+1FkMsKT+3isu8ibOjiQxIllCcpIrekJXXC3P9Lln+hpryjDqFmqvE5PmAbX+cNjtgTOQSQ
+1fDecgX7Y2i9+PGwF1pbs6oRDV01h57KVJBeX2e9z0gKkvcW9EFL5n/JWZO98sTmTULOrvg1x+P
9nWU32OGs8c2sz+HnQEy0NMSQbgmqv1mDTHSYpIZSM72Hn/cYtkQvyxKkwSsO+w8CvkihgCK2C6Z
5TZL+4f1sAR9PIFrm4eDQizTHQhfDx4QV0u6rvSIvv1ZxXFiXP1+tpRwc69T6DMTFtT7e1zmALAt
6XG2aPqJvdn/4jxbFKqpp47AI5hzpdBtCgILG8+SZMgYw2fidEoRC/3jo0jG/gW/Z1k0e8lnQCMG
NQ4EVRLCNNJeWyIxADSmY4oxNJeWqU8uXE93NrSX0sAIWNv0czLAHJY20PhazccOpP50gObBUPh4
Q+jfKNRX5rOTsE4xzLQFLHsE4qPH35GUTVh8f1lA7hRbaQPI/NGXFcV1SSfnNJnnPswNL8i6MaQx
JQZBZe595vKny1aUbkjVjx66BJy/gXlD9mT7uCrJat3d2qq5Ktkh8skWgvPMimithTOe069DoHHh
wMwRRmKMfQrsG/v9SUYFmeAOeWkuv9oCIH0/8EFia0Qua3hPzgXqSkMhArgEQzlwkH0O8+ThZmk8
bG3BkUJilBR3znx0ECRXDOW+UnbjZvp1M04SP4OllHA1f9mb8+hbyaG4jWYgb1wWCcMuZIYCmqHJ
lUeOOldT8v0QWXitTnBbrsJuB0oUglldbO4FzjgeLaDjsEOq2rez6c9D+2/b0YHxVqgp3JddKZKt
s8oONm4UdunxdLaNLq0L2VNoUK/nOGH+SYJrlyVNOiGuYVXwjiGGjOJ9pFjFpDD8qFnLwVCnkqeB
B/Mb+Sg6DP5T16SW53CuFpLFvtaDWLeS499hJGgbNypGruKejqgWV7VCL1oI9roeFx2jZlUwI9ah
ndZTiA4DxyANtoVcNnOjiZWKUFL+UmWWJq5YGtkBR5oRuDWUAnz2DoBXuwna+fx3g3+dZBrdLz9Y
9e/og6t1QBcPYgCLm5/FJ2oRFzWMpEPCWgD99fDyZj0QUMnRqIs5oAwuQkcLLr70IlVJsuJ5W+1p
CA6WQ40M9+5QnGLkp4oSYMBnbNPi3A3nJ9lceqNpJC2TSPngxk73KXJ+i0PiBW17dvTBMmLKWkbm
rfhCwM/3we23ggdz0HAXE4ej6l48/DcSNBBl3VJsxEzelcrWRM/KZjouyQPpJl0ctiEMUCxhLC47
GvZgV1X02E0yxbcMD5Uqj6SN/hBGID3H2Epy/G51cSI2X8tB8avdrbQS0wOq0Au0cCx/FX8aTdB9
iVAuYjHOvdasOhA9sfD2hpNmOCCYaT6LdX9jy+genmbwCSykT7T9k8ZHgfP5fBWgv+DauUfT9mwV
+LLMIoLKvMYOFiua+ORwyLeJiS2HlMGMnii1Dvx84LwD+SvB4jPD5Z6+fPOBi/nIH62pcJkkbWg2
YXl20fB1NC6LWgmJtGcY4mrrtsLzW/ecCjqNz1sAE6PUMKvt1FYoNCaItmTPWyABBZndaTVfTlaA
KQVUeDZpvMWPlRqaqb8Cz7C76Ed63HMbry4ivS81PNOUaHOrqlua374qKsyvGM5lhpmHdo8Me/LE
ElD0gIijFvx655JYMark9I6ifhoS9m1EPJTcoVfoQg+bYrdh83G58x/ObFfdrIeKEUaqzyNLWo5B
MzuvWXWIX3/TSoin93CHeUVPh8kWEzw0SRsRSyM976zgRHFpXFQuOpwe4Dxj/wRzztfuauVT+w4E
xdEnjXbNycOpY7A1zfUigexBPeldpkC9zSXCU6nthsOpHGZLn4sAWGu5MoAshjDOeoGeKsqWJOtu
I+ziHx3WNqPcO7OT1xjjWEnFTbBvEIbPkjVujnpeev0ODqFFhkLgK1USk1qVf9XM8+rg0z3xSnGM
bRGozOCSur4ZYBUQCcxuRWPVFmaIJB92OAdpZ+l3z7w/BNvQ0yYnsC6Zxb4ey5IgUFa85ZdhL6JS
vd5CfvWL8WRLi7leIkHK91Z/I33YhFdWtxFOI0MezPNH5T3HyR9go3OCqs0mZbUzUmwAQ0QyVAMt
T7GCGt92i4TTFZhFIMLNRwGKfRbRBQRwC6PZs481yIKc5ZZC9wW2hTG01Q+oC+lMKCszuJTazu95
+E9CeaCKsDWLgT/NSckz6d0Gp0a1B7z040IMUB0Gt59MMZwHlOsCgWaRqMax8X55FfPlH6w1FpgG
JGuB2zJlnSpWUfEKAgZa0aFL+xyjv6u/tHKZGfeUJqAXhvQrJ1b/nkTDJfrQ2Y21Vq1b1ol1sA9D
yBJ5F5MyfHq2J7LH5VsRrMfMUCiy5JPjhH8eGR6sErthTvLJ3GmwUCdmEO2n3LHpVT9RhJb7AhQ2
G7deNhXyy0hdZjUGsAW1xl+4OzevNIaCmtiDAcwXzAntMk8FkkCJnouRwmW2XsZIc/ApU4ENuisq
CR9QKoBsaqqa+43jdqQiwp0tNmmL31uisDQq1+7+/WswpKyFDD7AGtauzR0yorrkAdolsTc/gkyq
KdWBVeUlB890SolJFlQ5nFDh5Vn86hLN4txZhSdHya905Xl67nIgvVJGLhZMXhQBfGnjFBOsh8o4
JiEQC/37F3vmi52EUwmlJIDk00gYmNDMoiNx98lEhWuVE+AccivTlh1vaOPJ4P/RgOLwKiN7KEwc
ZHItMDPHY7Ncm+gWRG1RSaXeVW/KQRKo5WD4f1imhklGHEeVbVdOyFW2ElEVj4ogsKPTRXumwj6O
nkFFmT61/0c0n9G/i59Xc4aMk0/4QSuB/8GzF5XiDBq+9JvjfFclp/FdH+3RUkgIqaLjqSMNE3X9
RFzmZUxIsZROO0vfSmCmgbzuRvhKYKsMgciaBCAOtsTbjsd4aOpF90wTNntNxFUhc+r8ASdyWk/H
CArLzUwgFUorKNb4Gly5/9mu8GKUDpch2BtNH9CeX3fD9BFah4gsNpZ4zwhmah7i329AOYgkDSz0
z2MG28Bc5xW5r+pCU5arYlGc/OK84He3/WU2zgSlWjqSwkldMpX+hzzrAqYhddEN36nPBSVDg44b
l6wgR0aZCHdw447Req8iRk4CDmwTifxJnSttLR1MX7MilKg6mcCGZ3KND+vIzBE9JJUKblqWJpnQ
BZ/fClBF4UZNLOXtak0ixwmdtvwlXC9fQIk/N6kVGYX69jLJCZIB1Yb1+5AXieXx7eyXJex1WCSH
rgQ8hJDbsK9n15a6ai72LZcb3c7AlJPa4E+XKxF/Aj3oaJiKYDMfQ83WvT4WswvieJX2x+gMcVA4
Dx6j6Y+v32aWa3+3mc/TIIZE7hQFJebZm3KlO6KwalBfpi3x23g9k6iPjVHE1uzNjYBfKSFBrDlB
TmDhiFx+v+9vFX58CoZ1KysZOxIDTh3HVYT0p3JfryoXNo6UeeOgDgsEYPt1JbulTILd6jxgQWVT
ilXG5tb98Y5Irdp7obRPOwB9SBJN2QMv61znwR1jUEZ47pO3M7rJCKqvW973mx/XnPO6rwd61iDU
7fNBke0BM1i/RUvdAgxTWxPGDLdUGRsqyDoTzfJsFZuf8t6PaOiQPFL5ArIVMTauMQ6EK8Qnjl70
nt/ARBHF93xDJRwBqOtGilts1h0xrnZg69qqHCIU6VJr8wsGZ1sx8b6qR7AAvjHLm76yhC7jwviv
neb+8HoBtTpbCnfLIJRW/+b16DOaPHL38sxbJpV0UTpreKsWGOM2kj0QiSbgyGaphbp/NRwml3hF
pxvcSb6rJzSXnyLFFKEJmisd+U36iXy6YxhaJBUBzGNDrAXvVLngrvgalAjm/ncbdHss2I34Qe0S
CJDbf3nuvPAeR3qJH+tiN14bf3SvnCHb4u74znpj7RKW4OI++uHSbqBfL1cL3C7zauuVR8vsbERb
DtMYrkNzzg7gM0hH/c3XfIoaow2hWhNEAmDmWKcnBX3Mg7WDfhh7iXlYDxWBnSuM/9bhKBiyvICH
+Y+HNmLDwegKvzgZBCcWYRyZf3UruwnN4Kd65+/AdUelMyHlijnF+IcyOknvztArgA75qzBDmc2s
mgJYkkABNdhmOoiXzkUCgGMcBeAuDYkVPA5xwqyS39Q+2QWLTES8bAWydpMMuEWFWGNH8wcr8gM4
2PzU1FxX1ENETqEBEJw5JJp3G4AoiM0CQPCgkIKfGgnM+TdJxwtqffRwNgvkvqz5PcoUz8mUixhr
2kpbjeJJ/ehj4CkNmOn0Sr5xuGUdLGXa9Ldq+T1fAqygjvSdv2MdWjdyszthgWSoGhr5sE+J1FxI
JPKgOqX2Wt1+yKt67dp+rtYgurEzF6Ol5qxatooQpoHKGLn+CnjrlgvKjA+Om3+xBzVI7UWQm07s
0mT8inrgqj8U19slBGwQfREGwMDFQ1CJdfgzjtf2+4/y1/Xb9fb+XA73uao4ApeSZaXSwnAYzGh6
3/vDyHy4IJVo6ZHLJXbZXpGQPHAyxHVENN6wTve/DtlhUNOr7f22kgmjfzNBZt9BsiUEVSpuzFlK
hr4nBXBWmgP4j5o9bkzeft6BqPTjtK+n8wGo/sKkOBLUtImWBQz2KxmLf7uTdVddOQ8YwXsypKyv
Y5v0iwczQgwNvnULjJRLUVQb954sCqB/q+19JBnZUpCy7xwwiU1Bi3Ha9qZXsJd8dbKPagsn35PN
1JFlFhBXPbjXe+YQ/TwIsjFMrwv5VyxDmOlysN+mx2C9/Sf8VXha1x3/PWz5jv/4j/ZJVYyajFHT
CJSom4epnZ9grSUUIvzER6G+XDw4w2JXjxmNKjw41hvShAgkm37fjhQC3fLPpCjti5pXCdPz4U5l
eUh/RPgdVCB1qml0SG/op8QgL7Nt6VQUcIkP/9nmlHmGtu4EvOpMhUj8XwMgAXU11O3rWM+KymWl
UXObS1CtrErDCrA4gKbKoWhVX5ZJC2L8I4gvoKbEWItcFuU2T7iJCG1XlLQ34beyMSPEwyoLL6Kd
kjgWBZInA5mAAXQWupLTS2QV+xsge15HFg3HVHNBDUGtEue1HlmeF5HLZRA2RGLI6xZfFGe/QqX6
wzx6cvdqUPdvoRZX2Ai+D8MeBaz1BjoJU8E4VmkWo4NF/tWTMAiP0zLzzcobD3UPvsEDpspGTMfc
CJqEEVVnuwjf0e8U/LeA/4+vcUpurhSdHGJtwNcf3fXNLqO7JdeWroo9sAuARsJQiQUmt2OAK8Yn
oULFd2oMoK/9vcEuOovxv9eoT2hG4dpVgxnfd35ESdR5dHli1DYqisSBdOM7SBOLYE5b/1Qnv/Q7
jBcTAIfaVh5VM48etc3J9tDNKCkUM7pILGn/yz9ovz953FSjMJXuV+Kymjh40iTdLYKrHN+WNGOu
r8uEXaSaiwMpv/lD7HnUButX3lz7jikXaRlghqfZdg8XO2oCKcbWJXzpKAdhtdNHJ0FQpRE2FX28
AihWuUJXa4F7BpHz+6rnEADHQGsQXo5MWn5+NbCSfa56Uzj/HebSlIaFz3gdwg6slE0yYFZG1l0P
xm49F5Kh0uFvrQqO1gxufVUaroYf9yC4nmq09PXG8X7h5x0wG8iYem4h5RyIc0gIYRzQs3gFL6Dj
npVxhY1f9dIYjxsplzTowdahrw95jAs6mBOdSABRKhV34W2IVwyWXUM8Cu7yhfXa/f5y0M2x4noB
bFX4EtFJc7uXiK3V4lbMMFaZDhVMvuDgq/9HECon9jvGmOv1cT+Q7cseLJh7Jnv56k8Ebfcg3uiO
Ce2BaYqa4wcBSe0eHjaQZX2zx8DJcrMxKR3aSs1bUzNMnNpuWQW7iCFVcBVHcSvvfkfoIrQ1kmwr
XKGc3ENddvNoBRMU3csmHi3vWKB+IELav5oE+/4cU02liqYFKtWdVOw5b5e3oCmeP+aFTLpRKAXU
BK532TFwnshHFXCu66RcyosDVZbps3waWbZWp05W8/hkPf4G61TVhzUyxb4TLCpuk0CnOdafwscc
bPobVsgXnTJUbXSBZczyxmZUq5nyQTf/4DH/9ifjEo8OBkU1BsRAj+MAERU8wB9NlGQ2rf85y8Ur
mRodwcOpySMDzYcihwzt9xWhlxuya8XKVMDswrpiSEIY95C5VW5GhU+F+wkBT0yEJOQP56K+wJAA
eMM2XPT/HZ4zA4c+arOMpV0gIN8z6TV/Rka8a1sJjvaUgKSntsPy+UcoygSC8C1VxQ0OKFPoJXtW
AGAviD5TvjmrwuoHyLoAXcUgceO1D1wJ/IVGjdLXtL/02pHjswnR5EaUEoPx3oX72zoc7ZGR4aIO
RG4+U/vSzRzpKyOUYQP/H8S9hadSbKGZTLRAxHqrozh8jfYYFB8GG6/OhOaz1uPLbHhet+MVp/pZ
0/Ciws/hYGnoIUUJ4M14uAi4sc+deCAByQzdTM7/J64f7M1LdedEK+4L214PXK8lzHM7vTq/Rnpw
ePDHBtvOtb2dx6LALcCZgyu2HhXM8YeptrARYydyXzXHNetpKn2Py2OlLf9saPoFv73AK01v6ywx
OQVxHcivpX0mKiFHv9rRe6bLvVSdKrX4mLOan8NyGPEk13yrGnf95swhoL1dUWsEkJEAK4ROQz0u
Jrvy7bKHrnex3M/URFBPHOukk/Ro8kNDJH30FjQsQx5Czg19IftfHLs4CFhBrHHL2w1jlVF5W9Oc
Cm71+lMWlYT3uIIgtbzKa6bffajgAZtZRJn+1jbmI/7TRXZJXR+TifsM6GcN7R+WsND6LxeMr8Wr
qlreRWqYqyT8OMOJqyfPyzXwJQIDvGZY4Ee02NEPLMGr48pDt55PrxKB3GYM/q+9pQ9su1kyzFE2
4ZeUFEF+54h+H+fA2x4/WOvlGb9iA4AvAvnKRF2+adrg9BWuAYi7hyLQMbvz70NDGDyzev+uRZXN
9dqsVA2coZIQQQGeQRLNszfSwxVaqSjInnwyiIBLsy6+bNFOC3keRJdVddfriSOkr7f333hPAx+k
Zy+Y20G2QqSGXvkdzpemL/W2g1IxLvNZMq/BQuyxIwON51y67x4UVaUK2p9L65dWhQZilKhSdM6K
Cpo+SI7vtYRNM3mb+p6N8qtKWgMD5c+hLV71eJNt+b6hwKvc+IVSXEUdiInqjtysY+8hPqgrRlGr
ASUb5AzV7gYoeElhncNuruhcvaMFcAc/RhFceB3x9nywRBAQklVdRfcG8wnw1zqslow6ti6cbTBa
JL9DONDgb95irr96Xu0nXf6WDZyF2P80ZyI36PEi/bmwXYysYhb7fDXRtqf/G1UpB3DOiOPugrqe
BfGX0f0KAv89LV4WIfu/SQB/c1zmVxDMuF+M0K5UBXGjqdvQdGxn4tygSOlp6cGewZQWeyAlCM8/
6DF/aeOC0ul5At7Alh3VU8p3AWLSOit5+9GHsJqRoD/mmueIx4iqt7+8MORWeEZWgy0tww6Gvk8A
XNmTUDU7EcyJtWiQqZdZR3pil6yE8TyYLs0fTE4wivxJIIiF/zudzb2tCUNXsz6PClbVzbDaDqqz
+t5nnggQ9lH8Z+Ahc1jqsm49COp1do60bJVT1+3Lcy4hfxgcS8n6zjdDvskPTCNypo2PGCfNgYtI
22R8iGkX2oVn89rMYJZSJHJ8HfrPwOdmQ+KJL62FRJj58M7lR1EiHJKjqbQFBkKZJmC8IOJxL7yz
nUF1jBgl8kgIIONYLcd0mYOsmdFCmUo0HRj0+GHby1VtJV2ADqQNqrt0CQxBbXCzFJx56VfpxQDl
q4N13FiTi98dXPPU2tBG/zRvyGynYTBgS2bSJL5colugLtsPO+2DlkQmFMkC4p2mep4ZwtSNiZGq
k+/gVu/YvCNVBEMxbe12KLoVAYvL23FdUXpttxTmBf5fJ1WHDKnChxsM5ZHzYRkLG+5LKBrebgF0
OiJTRL9NbFDSveXuWziD6E44e1h9YVhB7gktDaT6p0nATUaobOLSEvreYmMVk7PF2JyttbDArYVE
67h/6sHuqFExg1WTJWLa507SLqFVvBcfEzIfIhhsTDxLuhRV2oVhyMIXkl+16xDaWrLNCyW9jBzl
LLwHFWg3XOahcxRmY6LBEeivSJ2TWK+3QdYTan4S0UW5yH7zFo8C5SO/SkARAqvqqdTIAOh+XUvj
GeJG9RI6/c4R4jF1vUf+jEx+lcTj5594zcF61hEsyd8eWV5sM++0NPhe0Hn8Cvz9u7cRChpuFK33
KBWTqO8pZdlCD9XoT84PqGH7jqGHG4OyMlxwbzp5LmI1GqDUYa+l7HvNm/nBJkugqzLPKGQQbaa+
mlsyVZW43o4TzcBseLSPYoYqJTFw3YZzONH7UAGu+2bPw7nc94EDFvsqZfmQU2OFZ4/UAHWsKWMF
IgVLK/BJ+hM2ie+6L/giyiFNqZAimiiH7PxbuN8SMb4B+VIiXnGbPUfFCLKxFdVgoqmP95t634uk
j7EvW+g6Vrg5R42meJFcXj3y12jU8P1XzmgglUcMZat4cLGePNcHtdmnv1/vb+Z7mMyK70NGBZU/
iWcVdlQIJgJyUNytTbFbRfUjwES380L9JnzfMwF0UnIZ8nqqVXNnBoaB9Vpg6avdGRaeIqUM4TLr
X7rx2wPn7xQQkFnUFF4H/Dw265zcyuUd484M6pilGUNQRqpJNJPziUgpNJxcBl/oZoTEcZkRn2vN
t6k595Mr+ja5uPTz3hcQ+xzl0J9VhPDniS58K4/XisbHs0crS+Ead1JEaEKjwC82cWxHSyPR6wMY
dUClPOU2GXd1yBGQa/rumguzZe6ZHsSt+t22ImRhBs5faKtpk6OMbtaixk/wtGtXHS7vRzcoBHb9
mPZt/rpwV/Acu621FhGYebAgqXPrz5pOciQi6KyWj2jlRc6HYRenOSqIITdxIiQwFpi8fxh6TW1c
vWiXiD7Ito2hze8jrrWsLZWeEEOhby732gvIP4dslSNxB5nZfhVuwaLV5LakDkV2wm1gOytPh8An
HqejR92XDPmH77UlRHB9WXNf8CAY2yaY6RD0v2qqrau3bbuQ22R0i2KG4OdcGEReAi6KbMVTSxzo
IGVZswUWsACXr/oexz+rQ13MRzYDmlfFfBqqxJ7xS8JDnJIsGzYjgTVoRg1+OlV8Wuu0nEINm39A
x0/N9uR5CW5ewaY80O20novhMHuCDZiMbIguEmL2VKKJKIT5XeQ6WQFRasohsL8HX2lx/KRj3ycs
8NNCb/oIG2nlj4sk+DTFGjnj1V/SGSVLFxJ06wryInImcS0W4jv+bs5kqO4xSCFKqXtfk9EZ8Llp
vnorUQm+k8MUc+OdPHVwkVVGZM/cc8bWFMIcMVi5BGfn3oajAJbAWA8AkV1yWX9p/IE67CfIoHEU
ZlFbvIb736Kk0TAN65aVC13t8fzxkfAounqXLpfT67hFEF559jpy65PJs0pwSDPNs5wsjOFULOHA
OwJeCDYNhAIljvi0+wLBuWhEyR1+Ur5dX5ZH+dy9rek/BBb+P+OlRz2oE/msZCoZdOH/yw5Y/lCJ
GTLPl/nIqeQYbOz44UrzD5GNsHykRTBg+IpwWvs4MX6IwYg3rimFJ8PIUujX238fGhmeDveIyMwA
cGq8igGHXcFb9EEbefz3Uib42npm/csXtqBgz63Jn4y8l9oz2nBADYTrStRh/A6HX5KjcqIJFTnN
GGx5KXYMUGF5H8qzWKwjCPXq8/xILz1SZfdFRrHSt1aTBwOYa4Aot1I24L247We6S9vZ0c2JMWlY
1hyGu1POCBTropDuAnE47A2qNq0G1dRNsO1CD8P3cPoYGO0ZuFzpY0CC5cSaz7jwxYuUaFaSriES
O2xEMT1WtX1LzmYHNjA72j/JYe0qClwIDjlreBzhneXui7/MV+OFAS1LsHKll4QZ6NFi/BtXX6RM
jjTSw/6+v/l3RkVCFdcFYYAKkBgHW8d0YOu4HmaeLkWjXYii+/5oAxXLyzgbt/tXC6pSh9pHIbri
OOk0m1hK3dYMVdY5Jt1EItMW+BpLMRNKhHXeEoV9XsdjKvHWjLTFAmipWmb3Bih4jGOAClNpTFfU
Ah9jYm4tTnKqHMLSG8gqiXkjRUDtQjW1opgDbk99Z4EbJOCDHLoJYKJUQ1j5O7bmKwgwBwXBUCx4
RV1Is8cD1PSJIW3gCxrFKrJG7hKYjc+jzV0TURa2IdiVpkh89hTWRUHyfIeCRs9R/LoMUNQ+9+dJ
/b+qJfCG7c54Q8cDcDWmbButCYQnfNGMhKrorbCny7jbIu0QDTJu2Ek8IBM6CX8kyFZsrkDxYhYT
SUhVdzicSWcfN0+ahsiGFK+v8iANlNtULJdX2ZfkaDisXNB489jJQGDccNdmAc3rULSGaLzFzA8Q
/yvbBPfHL0zF++ak5TwepRfkuP5b3bH/znQLTdUkgeMMvS0c1HLiW697xkL9p+/x8TboEVCn/SWz
eliprX1Il8ZlI2yx59B6qdgsPWp16uQ1mjZzGWZFPfZKUEtcWDZPqxT6AaF8ahPQ09HWoOQPrD3j
NlAnR5HeHeGj6A1OpcB49lemv1Byn4r4op0S8MT2QW0njRzH69mn1qXnQG4OTfFEH0FMUGL0lU5J
J4ojBjAiAg2Zzol2BpNXnz9vWLwT0EQVZsoss1wrJW8v+5xSAA+DI9EH5X3sje2BjFAzv1iCMjpB
mq+6BHMOH+eQjtWm916qL/qcHLhIuNaaciPbSP63tXRr45Nqc/qlgZDSUtSkv8CpBqcc0eH74rnf
OiLy6ubch70oGT/DmD2UcuG/0zBOrgbxfNi0uBDvfDopBmqgydOtRi7/dlsoskPmy2egcf0SF530
vXNOcft90KSVCETpRJpsFkbWhfmp8AukXNZyvE86dXvQphiWNZQn+0X5ClPZxuz0qygGddNUqpEs
4yfSnin967AwA3s5l4nKWDbY0pvCssqVYw4Ta3uXxnBI/BagFpVureyPLHEIsA44nwqCSsQlFNJr
YVOrrZyaIzAXPxEhqM0uTRiGOTBGZiJMVmS1/0chIbFtETDQ1KgQjJYN4ufPu+cjWEdrSMG/UHGQ
n7YKQox9R0uVQ9UH+Icjr+x98ZFtuKy/0Py2LK2bTqRvt9oSumtenbhvGCZ7B7LoiAKVPdfzPUEW
9T/7wCH6uzJliJ/XoeQKzb3N+yI4kVgP1APdkxDAqauko0dCjZKE9BxRtQsibn+BR/0szWXEFISx
jUxwSnqfo5SCkwRFdUAWRIy9ykuzcocD4zJOq8IVlnHhyAYyqZcWd4MVB+xC30TesjI+wGXaNLa7
khJxMxNlMljB9cfUZvF5au6lAfCaF+/IeJjE1YXE3RYsHFJ/jxbERBn/2TUud8L6VM03HceQABlp
hXIqX2YSZxZTkeYW1k4b7bYPYkcZH9TnjQN++573pLRrmw2oa4aFcrwcNH+QCodj5Rw+qgGYgP9R
3N9+Sj5YCFQPq1ef2qOwc4ueTnXBGt6Qq+F04C8/4EXv+XCE6g2HNLyfUvTD3uEe8i6zIIK1Oqo3
9DBsigs7Cz2MwPNx2639e0lK07pLALq2i60mZ9YC/br7MA9jaMyhsI4QjTeTwWNDc+/nmMdEs1js
HU66Bd6VAvuqcSK35j5OdY75MvxXMsiQY2D83aPjlf97Cvyd8sWaHMbt5LZw9RCO+3HObIiGInn8
jRn4DXxwPjxPqWSerB7aUJqqh3o+RBdUi519kiMoSoFWvS/j2xF96OL4N9VAt2/LgXRJZfkKEQbJ
kE0iLiqPzJXU7X9JNZlq7Oyoxas9eB3a0xnpdztzZjyxvKsbKfeNRQQQN/rcve1Z3KPVtPO4EWmm
qSNq4Zn/KkZE99LvGLMg5mr40oih8u8BPRKv/mAzF5U/8qeipd0J6uvtn/mqOVjqepZGl+umAMiF
bvk2w2mofV6PGDleNWnUCEESFMNQIleoPMpktCLCI8EQNTDCaEYgR/RRaQneEJEe8WrQ8KxDSH6F
qULhZG3GnLrxMff6xBx0E+jb9JiyXiyMjufj5g8OgWiHE7DxmqQPhZQO/2CpY7A59M7qIRRbQS/i
xChKEhariGnraNwJQhuwoU6EBFigxPlW/zKA5XacRulU731WBAF1bLdNOjeRYyyQklzfXp4aXN4a
f3ggTi2X8pnnGWrP5COH9Rua1aSjRzORkJwDQrg+ZiiIfZA/DiSiheIdU85Nc8XAyd5/jRdoLI1G
i4xbd8jalvUPiiHt8GTF3N0QmXQNBnzJfIWSZbpERaRNm/wn7VBmOYtsgwH+To7lHzeCfAwXFp9C
kTzQHZhRaiaY6sgOFfbP4JP83VoeU443Bd8D7KkcSo+4AzK3GWF6YV2wFksmNZK9FzCdzF3Wn2V4
PsAooDp5bedSAcTuViH5CvW7mcaUUj8R2VshYxDp7cX7nfMZ2ryIB8vz8HKk4nVy9EnhaYy2VmdS
b8JwB4TWUGupi0DmZtJ03uFa9hPhAzJMejLNPx6ZIV7OLrIZ7e1NuHI7yBsKSOUtr9jnNsGb44js
qqwTRVaFlh19resfeU9J/5yNOYX0Oe+yQyoPNWlC8NTkTxpc4r4DOCSwfeIceg25NuxlAG1pHWWI
qryYhH+JF/iNfCtvuN5ksjnMiIMQ4Lb1UagF9E7Heo1xGO8m+D6J2L9C87dfqKz8Evb7onywYtU6
hF/t+47BSOY5iaERhkY93RoTAOSRTqOO5ldwfaVoYeP4UThVDUKc7FZYkFKC/rPLcWspX4cDAMnj
XLtuC+qUa252mfqATgKBEdvjWyTC3VHYU/sc/VX5DNpPCH7bV66V5t1/LZXTObSxgeYpKnm4JgAs
+MAlF1BaEMN0ZG/RlH9NSiwvRiAx6j1f3vmRrDY66hih3+U59m37cwrGZz4KSe1YZ7lG+fCaX8lo
nHaPHhLmQ+Tyrb3msBcDhVGKNHalMwftr8CWazCFSaW26WdoJf3/YRuWNHFVzMgaiWF5xdcQ5eZ4
1+/9r43szvWv9WoNFNuTv+HdolEyc9L6Uk/UZ7BeoljsWO1B5FRgUztD4hKMPaPm0860s4NYX+Mu
AMO+mqMYHzM40OntJPAtbO5hDOt5Quh+6ixlMyphoxTrQv5nGoVcW2wKholnFZ8NU7xF1lMTvUHx
ZU/C/StuWDUvmig5V0XH7pHJgKxh0t09EFWhrds/aqKCnYpIWbWlNatjBnzugQfD2BQNlVenYSWt
kL2vvi8CssOc+6lKlYtjFj7xEDb2YoSbdtowJGGPeV6y5S5vmVLIMtPCl6vriiVkkM7byASkCY3f
jNkoeTH8MC4noMf48NWPjrUc9vhM1vqJ0Ky9wXp7WGgFeI4W5Br66L3W4Egn+x9vEXckA8TBxjeD
UqMMFqx+EkVn0FETc4R1w1ThRZdsAfd/8auuuFhvNwLN5Y43ppmdOt2J3DVBWpTXp+Vg4+u90U/F
A2vOMHedJW0aDf66O5Bxli97LKQ7dMuejxG9dnqwBYe6ogXfDEuRVnWj977nkhm4Gj64geCCTE8J
RhoppHddo8or9AnXhrpZ5uDCRxd/UUzKtTTyzlJVe8h+RyPU6RSSdYd7tLAdDsDjv5svLr8O29v0
b/+0LbSdGnN/mjT6GIkGOkZ2owUKTmte4nspg8bfK1sNaXyKHJSkpl1MgShUxgdIXL+HpQRJCE+G
FeyIdpsliQasb+c3v0R3q2UuT7FXYOBUoQK4luy5b7BHQwApOyhKEmwMW3aEhuzaKHtrakBEjcmO
hwsekphAPV6OgpjaeeoO1PFjcf0ru8X29u8zVWXKOXvmaqIc+BnCFmTux7LAGAOr2XRDpahfYqk1
k0GEhiVgeUusuhkZlyPi222ge/4w7NhrjMu7s6yH88yy5KFhMejinU5e3Kwqy3lvcUO6RzpGNpS2
MMxIHivw3hrNh+QyhqVACgajrpWYUbFBTRu3RLMA7pfTdcgvheE9DD4RRXtipvCruOJ/8sssaNfh
mEv66UIHbcb8cEC44UKqXaN0UdQrvQd1fM3HPMXx/GkqMhcF4T7RjRqsiXnz+GQ2WF8pbO9hvYqD
8zPx2YVREBlK7Wm9WjPR3nYJgR+q6uxw6u2gaX2QkYL1MOSGvj2qyV5+835rM6chh2Cel5eE/VRZ
bqSrhZOovj3+xoptq8NwnEJjPbVha+LlbU10m+ghNN2nD6MtoAYryOcNFSwJ4UEIbA8H4D4ULjWM
1PZSVlhipeY5YfcygnOGztTGOqP6LCBU3HE6N+wrUXw7qo3ePlXjyvs/r8uIs9cPOKzTBgNZGuVy
OK6CGMDZCSPpkI4Zj5VPDt9lIUTfw1E4ma9pGD24pA3ExfsVuBPgT80TtN/yXKtx0CPGWo4q9g/U
ce/DNQ/CAisoLUtZn9DGOiRrJwwDCx5N1IXK6IC3Lg1py8Fm/W5Rg+lRLHe2hS9dDKCmLySQCiVJ
0L5gH1wLoCYgBEpHm2a+yhZ4AhRbM6wxBFY1UkJebGuy6HCKYSskgC2TFuDrI2iVS0KvMlc/4Vjn
tX7wlTyquqiQ8IT3JzxWT1B35yJuEIrO++x9V8Cq36qBjlybIVMXRDluAOHXPRuBmnQGEbFW1jB+
wjyiWE2yYLwUAqJ7YNL2VSRbXxOeu8KWAbJ2H6sDdNtdX5QTNUkXd2k1uyWoIs2f5bMgWl3EZ2ML
mE/BgG9xcLugpxkH35N7dCJ0SdnbSQLpsaM+1Kkeu8lftb3UZGQxPQeHHJAdc/pt1ARUj0IQSUFs
2oC9+B97ur7Me2kphTzt8Rvj7dGM5nZpKu49730DnQTBYaxxwL5QDsCT6AWTb9lfOVAFYJh/FRLa
i5Q7imTP6TJv1q2EHXHSSogf24h1vA38D1yDEdLfJzKJP5paQ/zWnSWx3vuxESQnUDpxK+1naf6n
goam0+7hBDqvBL3OHenLkTnApM1KbmzI0ZpEMhmdhC59QOj0iD9dtukz/rlKRR8ar6KrEbkt5lwi
kt7nRdYRn1mwtVhsM9F2iTTAPMOF80mvM0sftJdvqrnDqIymQz2YPv/Ry4Bf9CoIoErdRqnJsZNz
NtbgDXdZLEnjGByvyJgN59iVv52LPEclwzIaPTnwKl//+HwmY5vArf3DvVsM+CjWFWDn/U+w65jn
vT0ACbx+y4EvAJ0dCNzgwP5c0V3Rsbu5pGK3WQ5c87dSpDtHIfVVUp6+MCmSK0kzuqr1xLqvKm1Z
sbb7+NT9cr1iBiFjlRedxd0FG0ZPyNE9wBfnmW85/mURTeHLgZQki36Gpoc8ZqQPHkI7/v9BfIm7
5ZQT2wimKIMH+4xOIAi2yfVRkPSds22mOhtOcWvTzCxdoeRpV+hY/Lgipbu5+XnwowT03xYRuRmB
xaAfrb8POp539THFQhqVuzshGre1BbzxQoO+6TMzw7smqmn50BnEnZtvBBLkdRZ1gvNKSAaxFqS/
oTPsH9ODjoShn19rjAziakk1Uh0IsjqIUBl+/aokNEzlXJzBQNjZ/3rVy6Z9Dqq/iBwmik3OxVPg
xVgJdwI9QqCtrpj4Hj4JgWNa1lgfM+aYesdOxhutHCWgYUZwubBODdER49PmPC81ltxZMEeKRATv
4sCi7UkkhpUKUTI+QfJTPpshVKY5nyj+JfAzfAiq8MoAuKfHb0ufEa5LYGpZ+z1zsRaxvZo6mcw9
mBXpH+UCTg9iA7vmcHCcUkNhXqLHaMzzqPdYhIaQxG3VMAVF1AEXvWUlq2FfvmgjvhTbMs1lC7Ne
PS2NQpMroHFp090oAek/lhxV6i3QrLFijkubIAlAMsYT03mKYAtmq7ERBG6PTLdDZ/Q+ECwaSYIY
xSjAQNmdLwPTSfwOhCt7dAcAZ7DWxvDzi0pAaXl8sZ3w/JknxLtWJjgH7CtXni4DFfwZtHMlwbfI
P6g+91rP7um6w9Wde6m+L6LwdqnjxWMp8RhOsf48k5SP23gQoqoLSg3X9bKiy2pnAroSYnY1VyWa
Ft2F4C/aM4akyjsdoJhqAla73DTP9f4d7jzo842uZY1AGO0C2ulVusL52Vg4BT6c3yIvYBwlouWz
zmF7/t01HxTzkPxevSiW8SBPEGRcSkL1ARpdUaHSfxP/DOkJwOHV6UtZLS+3jNevOaaIksDjBsW/
6jCBdMO/76+64QGoBztj9iKc+uPeU66pxAoxnJNe6Cmv0XXgQ1MxHCv43D0ZG6P7ABS/qcA/+UdT
WJwE/IcL5Od5HUkzK2W6RKyd5WgvdV0osNgviVcIaZaYKoIHBp6Hv2yE/VndRM/f573ggFzSynDc
J6X06YpPhQdVeXOCx6UxwrrSca4UxLbqCDmnoOIeigpwUl+vchH9aRhCfbwmeU1hYAjbsoluiQQy
eHdAsBEXz/Fcaady7WNn0nTFUv3d2z33l5cOgeO0De2/Eodzq/Xcf+Qbi0qFtiewwVebwSOI/A0T
HDo7MVxhe91sqBMcANcTtP7GL7pV4tF1uZcU5uAr8xiXEmrH/6PAj3dzmUo8gBTJL5fwaTHJ0C03
UxLXYcMKBuFTvXVr3C1gEEPaltyHMsnkq0pIas4aKguZPPfyJ5QahtFWtfCm0ltPDTxZKlWW/WEh
ZtQd31iHPyh1voqoxVUeawfQ/KIOPfrsL7kR+advWCICfckdiuFdp8PxouMLlDO3eH/6h12a9vJr
dVlTO5vYw1Rjn1y4IOa5ga1EyDKjcc4+fQMProb2dX2inkm4vh71ZcjQMEpKuSuNDxX1wxCJL/Bq
fRSfQxAvfnwMWIJYiRuxjZqUVNIA73nroTuhnAx7LAIUsDSCu6DgYI1Pcv21w9oye+OHZx1g8+hJ
aJMZBMNX39tRh9NjGUI6nuw/CcqIO66h77dLkds8rpRGW9/hQG4FfELDUdNt4Q0r1AYzSkiVaFsn
zU7dq9toi58BO6Cov7R54MqiTF6Uo/bfGipLQ5zik6uU7plIRiMoweVZrdcQ9QnTTE/3qT3m1pKr
CoTa6UJI0yWx7Ibyg3YgH9aGp1B0/likhkM//muFLjKukQc6+zDomYAbcjQPoC8jDzDRU9y+ftm0
FBcQpXwt4EcYUSvdPAlyn78nXg/WRCsgPQfABbetv9hJtAgmyiWBkyFqicqOerFX5N57dNkHjYaH
mlQfOOt1vC0EQz/2z5ACI28d1OElrZkuIuMYFzaUYB8QtQjwIqzzGL0ZHkj4tSMZVcprXEruNQZz
mF63Ng1DmHybqjI4lgvyQLsHZREfTjVRcehK45r/I5VRSz/lj+4UPc1uEHcDN1wwFA7AKGLwaf7K
nheZXcbOEn1PcGe0E/wbJUBQO7fdR+QfMKikX9fudI12iG6YjJODv/Q8izrkdq8DVxvPw6734ayx
iWTWna6pDoIuBdQXE0WmcGwK9FNg/avWIhMqCPRsZmawboAKWmU7b9icIQOcKQXRjkCJMsUZSEEf
uuo25+L0sW3BgII6vpyxxQCPs+zLA2CQWDYQWZAGdYZVy2B7Ie5A0NRRsNuB54YZt3kb2AGvA3wk
9RYHF4w3KUEVyd3UTHRSMrlAlFCRDl6l89d/3eQAU85FERMnPyyn6Aol6k83HG2Tcc+XKXteXTJN
vBqa5Gz3lpC+MkkBA1cNLyFGll3SFAhJ5D1LF6SM/mGKqWNbiZWsBfuI5rKXs0XysnCodoJRHswy
IF5qj8IU3QC+pC0/1aRijfkVoW7+HLsNmGMFcjMFPC5mmp2P2vMN9f9oZDcDhntq7+hExBjV80Cm
XQYfbAP3YmMylj0NMyRNI4yz8El8yu6tjQvdhmvS1HGVgEe/3e+QhUdkufzGgRPGz16DfrfnbL2j
X1qajjmRt+PGsJw+UB+HjMt1ZKAz20DdWAcqNSgRxwMvlDtCeaEi5Kzmaj0H4UwRWveM1TolBS3W
Wn3DAbxt0ezldpeSdDNnVOmt0wcxUB9qu3foFtz8JgMvqlKVoquO4ODiRed77PX7aMqbYJFqcQ+p
2DsladkcqYgejZoQfwdfLEI0zddOBjKJs8qAmfBIkGHvAzkHLSSTzxB1n+OkXiipGnRAAaf/JwLS
J7iK6wO5pmocbJZEm9vvnD0JtQuKJgmu59zpcRmLOg5tF+4mBEcW/3HXbnMb/B+HsSB+TSKv2Mpi
UMTCr/z+NGHuEqephJ400ooy9VZkoBNYYSndr0hOIPAzUXtfU8fFLOy92g0cP/kx5PAJ8HkAOrv+
OSF6JaPl4MVOgHEkPldNB0dPXF76LbP5vMRBVzGbMBo3tCe9Vf2F0G045AVlP8bwJNATSt5MQsQS
DCRgjXp51Vb+6kLwmP/r/L9IbuYewVSLFZH/zQiMymGkljq383XKXkMok+q4RxbcjVmZuMSrLSx/
lxv++gMOPNonHyl8EcpGfcWvPx9rLWh7NlVwUyrJQSlpFskPrHsQSCmezXw/zKynKhfWRuoJK4RU
iRwr0QvkcP1Fm1E2vd3v1bVCa6U4IeW1gaaqd7kXNA/fgUyssYj+U5Lqxr/eJkGyrYrszXdEu5y2
CcyngC4wFRhYvf1owk8n8v20zVYceU0tQs9o9K3G9Zd4NaHbgoyLN6RpWHv6MiNHKguSOWo29Nt2
cPn8BjX9M7u7QPATjnzN/IaYxuaUciacOUUH2vwN3Rc7MMiWA9JysYmwxZv2a5iTb7MEkiWnO1XE
OMeZ2A+caZ4Ec4x1wtTrsdf1i+5J2/n2mJUpqNiPl4XgLI2TGsOJV5/tzEcsOqEkVIbq66V/AIem
5IgIpcw0m5oipZmsjXsLS9K0zUSutbF39LVIrFTHRF56buNGnjClf2m6YDsk/BhXtyJehSVAbKcA
7AmIpOZEYp3cJvaCpdu9NXUJvmuNCkAdghxocqPesozNvmcKjkfpfFqVm/iMUbyC3vgooRamLMOh
IT07G0XPhaTk9CeBh3IN2wAslqQfmtE5puP06NESWzy1lcvNkh9LSONLDEcQCfRV2kKZu85QIT47
ZNbcJSs5xGQ5VOhZEajDibweGZzkX8cZG5udtt8eKAwz5vdkRpMG6hRNY043+AEgz+WWqm+dhFTJ
BMc+i+uzRVhfUXuZBfwqVx5VyD2O/DOm8l0TGPtE9ooaFE+uS90k2fafRjvr7G0r4q2wy7T7n134
Bey8plPqdZ7dY/uNQGcRVtJf85YgdJBRMkxtfLQfRFRDC7WXZ0gQVrimy6q6mXGHULv1wMU6d4N8
24//2nmIYUSDtX9nFj9axFB1ACTgxjeuPirVYK54r97XBecFz2fQQBhxbH9jm3TM6/u5FMrOGvRK
GCvd9qvsLIEbVXsLDQTJh9kTkEoK0L5Y+EoW9A4DiD5rgEnO0orebff+5ebw/KSjxVQ9Y8FpnSs9
BdGqCMR5i1rt6Sw+JhVLW6e4jpkfGn4eDMWasLfHvcvA/hi1+l2jtdY0EBRIegzii90ZL3gedmYh
Cz7Fd3UGnV5TCjb0u5KR2EJuiz3akfF/6k3M7w42D+W0no32Ll4ywjqcZedJ3Jf9nyBYLflg/Jq3
xHVNymNYD/RhezwjGc80dOcL80/kZKZEGIZ9cDbpbmI3enAggSwJFENN5gB6QMyHtqfKh9gZMCsN
ZpkLg57olq9JmI22ZzEeQ3gcajpZjICMFOzi27dn6d1R4Kb1ymYOZBOZL4Q9PVbtIGO9jQN3+oE2
1om3aHcOCi0JTZqAL8TFuJ8USboOqkyMnJdaVKAhm6DfjpZj2dlNNq+x0eW7c2CP+UWHlSgcyz3u
1z15uv5CxOvJUJ5qPYJGxTqB2ejf41oWlbHjcNRUz4dAUrc2MqUx43rarogACwty8nD37mkI15yf
5nyZD/BRt+liFkIACmmxeeejD8G8F5roQohiv/DlCHQQTLXHiwPo912yX6Ov14J256+iIHq5ZOni
bLkab5AC8iTxIgTMWPycrmCjxyjOhZjkt06PpYSK8RQ8YTw2dIXsesGBrBWHofhtPS4xP+b5apRt
ukTqKuxxpO8R7ZgLdLMKSH2ubTP3p2O4XwjpeLNjAFtd3qNPKGfSmn5Vd6ksbFfCNPtp6wqBPPf1
dQ/hcUfmN6vYInSFgu1Lfhg0LgeKRFiUeMe4HNaZYq8XLXWUyo9iT1DB9oH29rmhKqqM+Sk+8oR9
/Ly7HEH4L/dRueiJdzONygFwTUh5E1UKUFvDmL1OKwkgeagk6eIc/yhhfXZtBQ0GqLeeh77DyoeO
O0Oty4IJNrX7/sthno6zpXfSOH4cxltw3JbRN20sxH9+wLDBwZslNZ+AEpET7mXMF0RgfrMKjd4o
rFSc9dOBLMhxfJVoYXaBlezdqU3HEsgdCaXHaTTEIRuEBT2OilYl/3dm4jDkoBxBn0zJCHaBO0cj
A9zdXb767UPwdgcjh1zFv/6m/FR4GBx0NQdS0ltLFW0rhBpd4L/yE5eXmmrl7cexirPbWtDySMXI
xMCbSKHS24IfNw+uM+ojl6cPsAyqLRkBbW5WKjzMW9xxYe8cmNenDFtdu8sZRossY3O9dddUuqfA
iB9UbLZQYJ5J5O9QlCEH5/M3rkDJQATfDFtmq7+hqkYs65md784Yg6ryom7wev6SQHSYonbUBXdM
q8o8P/SuZNmcRw6gMJU+XtjW+tcrJMfX1SNY5OxGTfTkNGPQ4IkGnb3eHJDDOvkEvDp22i3Uy2Di
3KcSPmT7mDekORI+6Lw5Hw0U8+DlV0GZpFNmPgQE28O5JJ0enCe/6pftm0Ed14yAt2ELQhx0nbST
SRlysLOBUd7xiCUZnbAwjDU41QQ5aizQIp8xlz0gt5krCSAbNE6CwNmLqxkE0620s0kmPng7uW0O
goB9UZvUUYtd0liE3rMgNugBDLxKob8eTLxmFXyBTv69wP5Rpp1DEkxaz+8rh4U28pyWk06KNduK
W9rG5O1kLsVhc4zD2dIYzi1RjVQRLahA4mRrtrY56OJkYbsBdaVQMlyGgud2z8keEE2yI2DRNxpT
Man9AZT2QiYDfUjfVH/IG8KpBTh3gJ1AGloAoe1Jri8pmC5xY4gRWPC8QzDFe81vjF1oodnxkDbu
1kWIkGYaEqaTmq/BxVtR3h7GILVaEZEQK5jzkY96sQAmf7CItmA2MSfumQ9QXAoqQp3tr3O5YKfz
vL346TMUGzUn/Yu7gmG9igPwLth8Q/yqFDHqr1sQpdMeaDdEZUDmxc45fOgImCbFBKClgj/0dg2e
NkWmfKnMuNX7CNfntLDyekBte6E7U2QXaP8dN0QRU88GifY1FubWqWlfOUUkxAnFRGy3Rd0hfTH1
YHPLlZLBxxxXfldKWoLHg+3k5gUOLmZvqmRPUWJCLV9j2B8qwGSaGIPOeeHd5w7mR1P/MxlgoNvI
n/hqFPASTjYYvHBGU4qNeHrW0Ok/BCs5jZ6frsGKbkKgsWZZqXaT3s9yiCVBDu1NWiNl6gKn1zPC
3KstX7tUH5C6PUPLDsrWdaAdp0HZuFSpXJStxaBwVSmUpptGeoPxzEHQVXcoySQ9nziG3/wVlHBF
i9PwqpKBnP8ih0Z+/Oa+7SoX6jal/18V2lTaiC92O9i2jPMLpqIVfQVsw/tG4Gpugcb43PmxF7XP
bCwgz7p2j/PGLIOHThEvh7AzraR622mD6nnKH7FbIQG1XjUTlAwjTcDntqUJfCvGmciqovQ04gyq
Fjk68flZaCozTvUl3U6Jfi0OF3F7ykZrQGXGA0Rfv1LGTMxsS3uoPodRW4u9Mv17SQRx6i+Jx0Xv
D6L04eeIQw5iUFU9zrlP3zsi9oFzYI8M5JIeqrw991lR/5FyRZjR+vFZHJtahTzcgHGGRTe/oC5J
kOc/VUng7NcahCEbZsRbJVSIt4WhvaoAhgubKUZG06Ey7hDbgTqz2Qazm5eRvqUiT+GqXuTwmRAd
3rBZOuo+Oqn3YyiQMOyAP2he/543WxDi053aZKJ1tohnefC21KbR4EwtXNTIrqwmIFRU/+Lmmj75
D9IdsfC8GpGoPzUzu9CRy7/ieEQBBiCb7YlLzTm3z+km3EbMLIhDph53XKpcBKvWhGczGLmSu4YF
ExdtwJdbCMUHO6AeutN8s/RrXU8jUpgL7gShwe2MFZGA3BTo5uDnGwI/TPLHvm+XUvDOMOFKC1xC
VbWvNSheSAlTsXDkHBcvs2SWZnCCzW0ZYAiJFLqyWHKHts68vld+qFH7qPqqi+PJWQQuYkqcP5Jh
Vvf0+UyyqpBNlO0LYZwHVVmtDAed6QdY4YLw3RO5pe8zjST9Y4MI+nny4Ni1OB/P2j6wQoPr/qiF
cXjYPs+dRtNHfCvu+fl6fXAfUCMgpt+0kcgXMkVVas4OIst0BgS7obN7NOZ3rKKdJc/QQ4RTIOVq
ROFagC3PSTe8s3s43s03L4T826X5UdfYqVgrXovSUoH36oU5U2i8YmQdAnE9XWkGETeuur646F03
77A6vIzjhKGfBlOizmNLmE5M5ozZ+x0w1pgC8xvvp6mwx5f9o4NmVw3+OGSVHm5EBcsgkvaVce39
kwQUAveQsnNMR75SUa3YqIMvWWlYuoQWKD+dC42lV0ArLuf9Fh0QWq8/vksYJWuk2EIjnrB7Ois/
KcKLfXLPJX9E+L88yTP1a65084wTOOzf9eN2Ozy7+qjZ5CzJeIkoDZjI0qmme857mkAvtm+VW5/u
dljvg9bb5EWWbBa6/fIDh3Hh/DDzWniGSWxFXy3KleLo1Rb8KKDWkpv1mjhsgACoP0IIWVlQczOK
kajFa3Q5YeWtyFIxyvlrSaN+MtyVoufPxzFo48JmEDpy9IrsUZvVOhclmShcbWQ3FQtO2FcShYVF
DvHHri/5rMKeAzw1trj3gFVH03ekO26Y6idALAeyn+0OT6TLjSxODKT1n5KJeVXkO5H4KXC0EMi5
n9dUdyVqPmPy7/0sJEx75VbBtBFxYHudJkR0Xy7itiM6SZXnlXFfKFvCLOcFyCTX9+mwlfkAW+sW
bqXg2j8RAiYf8Tf0+kBA7QGg6soe0Bsdr9+/bR8ERrYq5J9EKGqMT9saXWhvcjS++kYTBhv2p5ZP
bZ+fmAAfoov4+/1KK5U2Uw5y8h+OulWsxRmPfpFoxThswHzFQKnp7SnWzUMOCM/YCDICuuqtyEva
cA27gV3rOnfUDZY0DEwen6pXz56WiUL6iK8ybe0DmSTQvSyuTMAdkGUkh5td6cnB2ujQbs3iTtkd
W9XhXjBxzYAalvJI/ofWzoFcJ32cuTRXR3jdrMduWcFIpQ/982mpl+tr+GWC/pQiIqnCyOwKp6qJ
AR+IAmbK3UzDrM6dApJNZG2fpYPWm/TsaRt+dh2hkQ3W1+Kt1vbU4GLFXcKp/hbiQ/G8DTt0ILp7
CMXPJSpRgHGQLURbXvYKZRymthAGxiI1qjMZFwG2RuP65wRhamdJQrM6j7ygjHrGZoTS5iy+rGYG
sSqRnZ6kUkrmx96aUwZf/El0BeEWX9s4ezSytVZI+n+fD77Ub0tHNtJo8zDg9zTvBzj2WBAuUnzd
+yEW2JoYPMS1UbMAqx+tt2+OhzZp8bqBzOdGMMMfe3haQVVCM18IriFeIo6eQIO7OIYKBhX+STvj
2ex29G+lFd7LmOQ2MszcLR5Y6Ru8c2xzUES+6UnPJlZT6YHs17khz/TvErhMTJm6HcsWswcH2ZXO
FkRL4+5xQTG8z/i18A45ENJ7ieUg1QpUnfCteb9VRmPZkeczEN3JzGIHmeFJBXbzRfMtnPc9ufD3
XNILC2fWLpz1xYietOubwMSKtW6PjQ18YX/f1wVh3I4hqIwF7N+Lf5Rc8g3bVlclp2qgvDBANHXv
YL7XZ6U/TuVfuXPBfR3YysGyqRZEdUOrMw/FTx1h/7YbvkpCZCO6loUSCbzAIJLJEUhQw9bkBe1b
GGR031AUJ9UgTjqUkPYMTId9K4SlZIMwCnD7zuOfhjxJTEq5vgb+AlOkh57Q4xGMeltXTaC9yM/s
Zm4ZNqGA+M00SpqWm0Y3yGR+4oJ0YcC5R7rOfp4TZ9mTinykyQQlJ5bXJDcVIOlq+gGUmTfhLxYo
YdGwcQP+Qqxj7i3tHUQphSJfcKoLZr0tJlJhzrQsvv+ylfILuVecUEkxKcam1Fv5hggfLFJ4Vp3F
HQry0Z3FDBgOKlhIWRmrY4BhNZoiWRfc4JJkucYm6YVwZMtvJdJzc3cPE6XuvyV8rf6x0LwEUl4V
EWYYWWiR+un9HOYBPQ5l8+1+HXgjMLhbDnjBHsGIVmgIDsrnIYOlP9rmKDuYAbRpabT+McC1nf5o
WF69COQ1NRSV8fTHMDLhFhib8HR1Nv7fUZ93ONBYWf2VKZn13dU0nGpR3vYIg59TeDum8Stg/qSl
XtSvM9jTePivsSegFR1X02S3JRLRjf6bJLqgYfYBWOjQPn5jHUrstzap8+H3tmhbulXA+81T43dO
dm377MxAuk3elbC62EoSnNLUMCjQhQI4mhDlARsuIZlu288mJcB3nVDBtbC+xLM4D+29X7gYbkDh
YRSZ/EjveBTH4Ui+fqKUzKeuIF7Ncf5UEUZ9vSNxOd0MwdiepjGLpZ7T2c5xgdIItyyAzQ0lzZwe
1ImQWktz2dsmBay5UsD5MeMD3zssaTUu/ZsLEborTQ5WkRAj9D+MocFBNR0qDP/cnGOhFUCM8GOa
vUcXkqG6JEuDYsVLIqJBkXsCwhwxbn3k8G+0V/fiRAVawjNgzddjviLKatndGmW5JcPn2HDiE/34
KjTYWR8C9c+L3nFyv1zxWAuQ2UcQ7pCOe23CzNVtUElTNEz4uz/qp/ts6HspEU0ADcUVhafXiwFD
SXoTFWr9iefa8SAlR5gA7dFJQiyuHDeyKn65U8GF3M2mhb+K77Smz9bOWKY6vTKJfkhGicNt6266
M28gK0+KtDS+kihO9DGZzwc3N2uRKKCOA5Ga6RknZUnbvlXkxknrzpNbFQSYBkD0k5nd7V8MnXJb
WK6CPH88v1Q6PzdJ5eVVdWe6VTK45VV75GMMU6S7lBbDRJsQvZITV8xH4FIkUhAE2H9xcXmrnHK1
OLjmoVVg/IqovBmpAopddyI4dTDnOWiInc3O0QFg+iQS4U+JD97CCZ/f2ebfyJfSRZRf45iSL9SR
LILaFPxXHLZO3BNQcyaaQoKULnrQrgn4JdXfF+3jjuO1IFT/FpivRHOGpIONocO6lhwNJVGje2u4
NldZa8XbII8+ePhcIShsH0XRV11Wf1f7zanq8Btb31CpKVlzztAXQQx5K5WePcEwzQTP892n1CTy
OIb8hVasS07IYUklCXtRy9W/i495w+Rg/xYbSGKpdYaFQhAL4WVa3Whhj7YYicNhzrVblB/DhRRj
3jKdjbuI3hg+opD+o8zl5HxwTiKcsksGRlqhfT2Sv9keRYfU6Rny/36BdgmrZ56JVUIEF6u7b3k7
A9UWHy5N/vbQKBV3ei2tGxfbeBbpoPUc/lwrGmGdsh0QsSJsvT/aeVYeGQXkTNLzi75THsyhJt0j
f4Ce0GFsE6LeJFieFkn4sBkV1fTxVpM250mxVaYuX+Xi4QX8FTzmIDnsMQWLDvaAbXU0exU2dCno
J4UfSy9yXsq+NWTT7biYpi4hc8WCTP8pYwtDEehkTEwMW9IWaRZqdINWYVojHzB0GNmnYEcuqMHX
ow01pyTlldQfy3YOoNNYaZfYgHR3aPDyjdkv53vdbOKf0vEQUnwHJCnlEOj5GoJv/1X/sC+sdTfs
ATlHjazH2OWXmsQox9bQk8Z3AOtlRiS/TL01E1K1y8emOolaqk03m0eJMIB1GdekCkFW+z7pIoql
GY3hL/ccW2j91W20LQNWQL5TR2qcNoabsMPNsj68E0+XVmarlqZESE1y1Bv8ppZf1bAQ74ZXRydr
PXJZ2MMuWauSAaH3o0EmEGDyh/T2MnVGmOX5uHZkhmb2gTmrOdBFQQaLtWZMwsNZZIJODFfvslmz
TlQPomy4DbFSkG/DEB1ysSLQ2+MLEdhmO2C3jktclu2iYPQbdjGsA7rZJFn4Ib3DeqN0ygU2Yzif
n9uTiQsMnKL8brJ67fjx0vU0VbZKJe/rndc/6QYt6pEIuYh/bLdMIUqteZPzYI3taeTTKs7llNsN
onoLznyJbfDTVQwQS4F8NkrONwVOSG8s/qFnYMDaVBOVvK7BhI8myR10DSkqSH5Oi/J8GuOvUP1S
7JTol2szFBaQVGGvkIXO/24obR5zYfs6sDmcBQZVO4j33xg1Ojv0LNkp6FoVb8fqUyoQUo8k0AJt
ocsIGCaHRwaD6/KVwKwoDVzMcW2JfXfH3PSgSMSxttbOrDQ8nWeBpalL0turXQFzJS8PGsEb4xwN
ejx9i/9iKymyzAUBmuwdJXbt35xpG8TFNUaXJ0xa2hS8iuZPQ/P1pobKyN6xzuWevPMz2uqwlssr
edRWiiqo1x1cyE6YQFm0UYryqw21v2y6WfQtCV0DZE4jN35RDTdHs1Y5RWC37ufhjNgfMVKFWYyb
xbLb8Aaa+FnOvotWVpI6MIndeY8EFijO+z5zsc2qmGBLMV2yjnYPNSiXBQGhArkP8KUunFdONLWc
cLULtd23idFLXr2qd7ugVAPU1y9bSdq2OUMOchVLeHMBYVIBe2tf7MGBzJHHJjwZGNkyCcj8GGDV
Aj1j9GU5jf6j3FUNYtxC8gQqt/NPYix1wU1TL8ndTD8d5bsEN96f7r0fzZDYI4uSqrqjB9AQ75oO
dUql0cQFjddfFOO+d2eQVMThAq/XEQwTZLtX7olFL98CxEr3zQZyA1Hnlx4KfA+RkAMIThZOwCW1
8ZamS8IDJdEu/gYJYtQDe6McoWyqaLPQUcBLX1Mql3wh5BBmgZdFoMlNlgi69jbS+B70bERzpuq3
b16iHFikFE3gzsjl+ePwRqbQDdjKd9qDb4kuSIy4LDUZCcvsz6xn8OGoUB05yyE85YSnAGQqjvGu
IsvtzRfVCAYX3WnEy7BaM3nwg1hOXgl0/5jn7A6pxZFAANTJBgvz3ECrUnYweGpBMptaHwvUpZoN
qdh3P10Kc/XOxfA5BgltJX6pfIDQMGUyec8EhTlrDJrT0EoHjOaSvjGNVqvqKzzz0F4qjgi/maeH
Qtwx+l8/zMks4oPqITHnBB1NPhTTQufLmYL88hgSpQGj17UhUmivOpJNLYZPLBzAdG3ZvtmMS+2B
eEaiT5jkeQ/q4ZdLbRKfWbieq1x3e5D2U1gR2HBGSHqlLzy1feZoZMEQCyIRTuaocQ8o9YtoQHoA
iIXj+uqom3/LT6BD1gw7arHGGMVGq+L+y7pfBk5KdnDqzKweEhjOJvDq9uWl7fE4e8d7RyuaVa/J
CdjlQfaXjWKBtKqjRoUNRJieQ6Zu/8Q829lEkMq4DwzePoeMylP9wWGn7I/zaGHcDMzk7fGSMknT
y5jKTpvXGoK2oNtwMMKV7/5jnHOXvU2Yu/7Z/QXJ+sATdbC9/7DyAT1DG9cedrw5SmXvhQ6uJUUv
kgkg/Qdho4c7bs0nmpUFdhuM61awp1lqZ27/Gj5TdNAPN23AhjITG9RV1mLvCQmas7nm/mGnLi4O
QOkzQ5xFtsOtiQIe6a5e730xNuTPdkF/yaHSPpCC70xVonPnozjiRYVCiSr5Y817eRnY2GWSfVzf
7vkn+Nc5GPOiIOF86/AlN/YTDOvCIOSSzSS9ZgD7/r/fNbPD2S/uQWXEFQ1sWwrAY2zNLQN354Sa
G4B8TNsoStWG3gLwERUVGDbVAVXbXAMIZKJbOZeTJY0rRPjxXeK8M0iclzaoCOPxMGVV90OaCYm9
DytykNpZyWGaXhFSl4opMoSBR90qGDKRTEVwQ3tFucEHPu79LN+ugsxEbG+UXNc7wYZ2Wq0tYYcc
dfTgiu8bjp1p3FDyyq3hcYfPrbwqq3Rr9eMe0A1pFEQ5FI2UoyuVFKFQfdIRNvk2GZbZNL0z1ljc
B52gAscPt74r/uNOgivZ+6McZ8GIyLBHIOcFX49d4cjbTniOQcxQoAnQAC5nqxhdOKuAa4UZoSN1
b8zytAeMsk9MJiRalUbUnlYRCvsdLmF9AlSaX19ktwX3AOgT4F7Mv1POdsavDYZE176BlYWA/wbs
x82FEYAbbjXi2A/qBt6FlNc/mu6r8SLOFMhk3Z51J2aAICi8PflC9/T+ThijceZW4h9pTUxqW1Iy
LBQP+k8uo73knYLmMjXPfJTJYzpd+Fc6WM7oQ1K0/b65FLiO29Q+dBODUdeKw31nyS3GclUp95ql
JUzNuRQGufGdI0dgSbwmNhGE5TijDwTvO5/5oNy59GZbaJulsiC1yOgOt7Lg2t2fQ4etwtGcsqGS
631eCErc8PnlmtM62b8RoL5yw+tOIdY070pmvXlajaURpqYhLQ/SR9WCLl9seF/JIx5KdxzVc7eA
5WQZrOaoq//4QD1F6jTDMP7jCjNkXxcWblSoH+6yzZGw+u4pNX2k5623o194nicwGq8Afa/MXBdB
8qmiqSiescN36gNDC5vHntvXLdziepLpQaqmqDCodfSGk+rWFe6BrWgAuoGF5vh4L/2ZX8f4+IEV
onX3zbWlF8dH6ICpNEz/8pZ/hxhS2Fzqbgb0aZZUz9Gh7p2ew/3iu0/x+wLrn0SnJ83JPZj20LkH
qof3KoF+xRiSpEaV6R6zf7ZZNQtTXln0bbk37Xtce3TH4OeDxjrBlybyyKIo7au/MFG7Y7DWU8IM
a6xGQ5QFcO5u3NGD8Yo78SA7bnTRSSKKJKlevL9YA0AaRooj8N2YpRboY70HgHguX6X2M2gYXJnc
BlR7zCZfE/YxxGEQi5IgGj/R7gEvtvV/F5y+47jaMRrnwxTVnu7dgibGLxLkjhnNLVy3a8u3m6js
Sz8P+jfarYmqctotfEdlkHPO01SEMiFQljl+uqY6yD10bfKXhKYyAHG1bsgTohN4bjpxTxHcOQHT
Xao26+i2Dh5/Qb73ccrDhVPAK/fxgZB3RfeiRPkDeDBOKLNjPDL1dQ3RM4Q5LJB3b8NXI2t0yy68
+iu7l8k5yWhL52Ctnn063LT0P9VU3IR0KwVNRYkTWaNmLJhvNuAzrs9xi/J5rj2ZulGyIupkVtjQ
0whdxZtX8/FOH5aJqgr43wDa99oCXxRl4X3mXn4rURKhJWTaYPC5N7UPuyGd6Kj94AF9BtyP0KmS
lXXoFdIM7hvEvziSgMfy/NWtTdFzOJZdvrWqrhiHzYPxSlMkyLK8QDj9Rh0AAED0+HVmIxXMKFHq
Vkp3lXJDgtCgk4GNxjm5Eo2cvw48RqlmddskEPNW6XgxBu9QM1ZvANLMCEYQICI0KP19o3vQKF//
wia/blNhX8WvMc0uMVGIumvXbLjeX3eiGJ2IQ8QdR5JKnsovyAJNwQWVVYrmE3VnJXCFGnZY/OBG
VkLyGInvF+CuyzbVTH+h3H71cKSrNMwmvWWJyhQqMYpFVlGzYRBUtjn0QoZkoLEfCG6SToSLpMqt
ZcFV4ba++v0K+9eRrkATc3PWBtBWbo2xQvm9oKNJMRfESxPxiNAjEo2/aJqiV3bJgRrbMGgRZ3oU
cwbzFskMCmDWG68r1IAvgeTQHYvF499xasNsvbNj79TPInoY8HeqcKX95aW+MmR4Arx7AftrU3QB
adcSGdTg0ZGIXTr8BpQLj6yTo0xUiaYRy7AUu4GQ4mN8EBK/HvJ7RtP0/MOwQk7WitN+MX3SnmZ5
VqEcsP1WPMj8v+RfTo9y/kt0PRqpNF26ADq7KEEHV8V8PLG04LeaqBgp2pcbrfhPMxGFnpFGI8Xi
MipafG+x787Whv6T/Eng9QhRbgDmvYrjMiHcv3onWm3fYV12Use1zYVVEHu0I1FJKlZhx4d5wEVw
7Wg7AwrdjqLrSTTRDpGTJbJYwhX9TxKp+UzSz+TUm2Mg/sQyc7vqBB6MWAIcjWfR7/XI+ZcMKacx
LRuit0XgWNQ+U2LxVuUjVwb1CMQm/fagFIsuqKhhZRHR8tJulTQBYsQEmpSzJKfFfY36oFXa4VA8
EGgkG+pheNPFopykImHy8pnXIak3RFPUDo+fSwsodIj4yQydIZSLOXOaM6rmR8GimEGnc/hCS7x9
YmC1D0mvn1Kbi7lEUdEeeF9KDs7wBeIO2aAtsCeZfhhun5lrU8cC6cxxeRdPtxj+VxYQpqmPij2u
nVqW4i56bmDCTCu701o2iKiyVnpnRv1pKYN6MVeWjyHcqRerdYMtiZDNSbcvwMV/futUMwz+RZnN
D8D+X7Em2TSeRnu3NskIAEPB6BVRllLr4vJJWTtrjtVbAc3m2I0U2evUsJT4HZbUyANcyl2u142g
gLHXB9FT5To8d3Byho1v7XjphQybq00eiezOQNZnll0grgJvdNOXUKSwUraWRuAAy5agOrKH24UB
8lFFPCuaMidO1Qt1VSD4gJF8SVKtQ8vWAl5PzmN43OCwqKkvH00uRlqfaKFO51+OVKC9IxLOMGpA
8VSFzcklA+MTyVgY6UuuQrSIEo8pV4QSbpuTjOHigtcFG9yPWcDlDOVZROAd4dJYdSIMIp7fhtxv
ESINCMQg4rw4ovROwiAYd0fy3yNy7oeJG/nZ6ufipIj91nWBKCrVtGXSIUE/t9f4h/9WkAxZ4jpk
qLMOuzgEfYvtBwPLVs1mLi1bz/vM/wQLYA6BmTriRJro65o5x2vv2EaEQeb1qJwBRWwsd5jfdZiw
sARiF3XQnk0X1DflZ0BR0sBs4Egq1Zj//IlVcMT+5lnB/MloaiNUOeRHJxlli3mW/bDyFumehRl4
SuQti0PEU7rzXxeoPJXHl6KWlsKzJRQOWK1+GHSZ0z2b6auwAldBu9BClFUOdXIF38fCOPPEvab1
kDV58po68QrpxyZJAXXP4BqNf6113HtgpDKuEtvY3mueZ/K/lS6kD2D2LI/Dh+yw1yqOkeF0jRb6
wwh6XE51UlYWEwk3ukI85PWoUfiMQbonju64K3p7QmzP0GuuOuORyyD64HoCGnEh1nbDoBc4FHa3
Ds9MRAhWAnnu04eXFVIo5l5Ci30+mP2FQahmr1uqmzZ+JJIdNRmOLBVph3Tju0jhxC7Ir/k1iQ17
VdQ+8OvnyFs0bG0RIM4ldxqXEPF/g+49/YiQ4dEOns/iBLN8/23IZkDhc1Sl0trDKvOg5Qqkut0O
biqxPjY0WG3dMGFst/mHYqsb+2bKoJFzADaBC1vzmc7bxmAEliLniNgVheh8MvT8exGA3ASwbpMg
rjpxi/UIQKsGaiDTDSU9EsX05wvqN1MKmMcIhJzfO0t4X/K421B0XgnJc6Vn2ZERovi76t4uiXb+
6QB/NEVNDST4E66+aPTHBSfhJEejmz/q2GxEh3gpDUhhQ/EODsfNugx7re7teZyEMOm9B2fZ3lj3
KmsEcvKa73PKKFXUXBkU92rEog20KOmn6fmG88y7WkpHx6FZf8D1LsKtc84fIks0b9fSFds/uAaX
YexgOMXFG82AlMU6Sqj3C+KLu5pp7yT4fSW0v/LQ2QRBJoCWXiYvTGvgpNvC/8sJ4Ydu1ZtYDokn
ykSBHryZDLiB6lOZSDZqh98udmJFa+Svd9V1VxzJyXdiPCytruYPp1kWh0kWWLUFmW7e2LU0hLEl
NbYzzbxmT9kOW6Ywu+QMhqJrOInT7su4FfFjf44Wm0hpTnQJy/BXs+/8L4e/xqkMNF1z90uu3sIG
1pNWfaFTKAUeBbCL99ZRryu613FdOhuqz6oHV7kdUC/45icx4iiQzBOckCOGtpluSEbw/rNclVAN
b4ARgUaNfM83W+TtvuonleUYjuupyAcrJBPP99Fr0cEN0wVDl0NLGoaNX3HQ7Aj5drpUeTTOkbY5
YTqAOFxto5VqT7lSCV1tUb9i246sDIetxNKA+rDnbX0XWbxsAr7Y0xp4KKocEjbXehDv70avuyaX
SOvk0yp4ua9bGvlumk22U1Ca+HxX9Ow3UirFvm+cxsBswjKJgM0IiVO849AaGo5ozdJ/nzX2UOet
q5l7JGVNWAOvABYNvNGJ2hkY8VSoF6IwqDutDLbqbaKIMTYrtWDC8MUm/sdhgHJb4PC8mW20JtNP
lg/zOwY5xArOPjLZ1Dze9yMrkwHNL8GPZzPxwFr+FJT5ANaO4s8TyPabcanBD4NOyn88zdi678WD
68TlfAUhu4cVWdenBStjoOIpBGHOCyydwKf4MbRyDuVFWNyJF9v8ajCmIdlTU/fNneXJ0zNBUBtn
HGOKMD6XqfvFk6kUEXAa92Du8qa1UxJilorDSI5T3App2ket1O7IgqI5YQB7C/7E5k33Xqw+dn2K
+xVBQT1q6hNINjLRg3p2v5y573sbwqTVR8UCcuFv559cW8I0VFUwqYEZFniOkY88ngSFvsa9BLOm
bofMjyAQNvGedlC8MHzwO052wc4HBRmBTKBIbbYYZD7St4qBzaaYpsFfQX44AjbKkZRi0DibzoTO
CU4vmTodC7zxGHSzDPQ0HGftzSsLkBDONw9+I+x/0EwC+a2Vg+OsxC4l5R8QXTKE/t5QSGV0asdq
oolNJ3tTf9CRk+ppcDVoUwg2WhWZMobvb+sAhcj4x4WrVlz8cRuZm661XsQvjf+GT+2Qe4bOq16+
+bWrs7AebM+fUJ3/ciiyUg5Oxx3QEqSEMOn/x3VPtA/I0Vix5tUht7D7SBVMF9GzPhiRsoO1o6wl
ENrpgkpM3UgzFnrzKhYZpvaePNB50PB3IsxNbea7cSpr5oMcT8eGOo4NH246P2CsSTv4JW8gZfwh
MWchzXxzBnpWJc6Ot9q22rMOMzpDePJf48K66Fn13zN2hjy2HukwVMmZmNdLMHbB+2iRqgXmbdbc
kD79uDHyyn5diz1P6SM3FUoCv78srKwI+JxYGmOBLGLaSnAAk1mo08auU9kRZRMvsrwByYFJHzGU
ewkAE73a79neEpRBpYQsh075fvXQdrEoel6C8xDME7Opq0cqCTLgAYjvYI8PqhYrvF0KlIl8JxzM
vJIrf1e9yCkYeTI4nVyUPBe7hf4yV58iHyVwlgIpONtoKwgmIcS7N/jqTvKok4G+DRFYOXzxQOi/
cuq+T7hN9j1jIuR90JEG+BLUcim+pY0E+/7nlbxdNE0vqay6pialdHz8TPYAFt5wDcuZw9NAhCH2
PiAn5aD1Ww+DRQQGirDoBFBIv/AXMVtD1rm9xzUngRVt3UBL0vLQX6Fzf78e2/xbuJY2PjAoAPos
tGA33Zty4vsvPggHePDZmAK2v3Q5Fe90utJMPVL4zx7KM8wQKeXHX1L4lInMyRudvmEnFVf/+cqt
gX8oQSWQ5wlkrJitKBpeb3zM+qgObIic4gKbjaH2SIay3ZS6vaVWEsqxbGJTHAQycqKVrC87vLOR
4W66wKUZYpN7f769TY3HgAZkBzQoGuIbTDnkmuanXecPW+fON79X3TReqFTofpMpBfNyMkAc82F4
sB8nQDXMxUyCTPa2uA4Aku/VZ44SVaLdp9BGiTuQAyFZnf2irG5DqLMgwSyVXxlOGgI99atLDtnX
mlbdq0gydRfwBP8XZ03BMI/FwtpCUxbEYeIri4o0ZmS+tdIq6K0sYC3SSqwiHY+KiCHEE1DywexU
Fo0EkURhqhLtQFp5AaWeuMlYckI8P1YfnfgQt+C4h7Cs7ICQ/EulPVNGbozJ1ADybMmc7RmfFEKK
QC8/edSut6B6bwh6d3YdhHt8E37plnnTbe8WJ3lEp6w1JF54xiebSADO+/rTyJWT1J3pfRFIACrn
COUMEE2Rhcz20KgsJJX/mlTTwuaYX0+rB9NSf/K6qz+fHkopE8+dtPB3bM+zHyprDA7kzubtsSDx
zFy0GUL4vsQVOZsWR2LD9nl06aF7BsTxgy6nkj3Hb7yWoX9U6HxSLgHuUxEdGtGSIErGm40f3QY/
jxRhZZ+j7MSCWHEsXmkzbp4CM1wTKw9/CrpTDp/1BxSevpn1Rymftg6L1OEnqFykykJKHaxzeByd
fGnIqBSeEJsN2aMtZXzSPI4t2+FBd5JYZznh3uLRcs0M46Xp//yDy2bsV2sBPL/jftH5vvoLCkSM
AJ9r/scboolUr3Wftp1abHdSkMOxcS0lT9MQfR5obMh2SMw43zn7KQtv11+7uTdCgooihaVPYaRq
Lvu7bTbDcHn82y0DS5XCU3TtVyDvBZwNiRJS3dIZDr9bIFhLWcPtXZuBynXSOIT7y+Vzpfm8LLDU
wmlj48AeEhI2utcZcH1JPO46Avh29avW5w5uImS+X+NXNxc7tpCGw3P4mpDrFOmQjZe83zO0W629
E+gbKJplrCHPF338esGfNeMSWimG/hLyRrb8StxaZgBg6tDqKOOwtaKgFchvpU2k1HSZSiAQtJkX
HzjkVJ29nJrmvIYctKRiMEZn5fK2O8mCxYKfeitTsCWWR7dwHnmndaY2aD67BEb/Zb4xmsQocnxo
tUX+W5p0LwU7oEX/bCNsoolURfeWm2h95jzjp3DGxZWvOSp76jLe6pWGN16VRf0hICQXPenO8Yo/
30XnVAR2h9XOhcYgjtrMD+DDFKU6IL37pTzb3fpbX2sjbwVIcwRdo5kLQVm4oBDrARSH1aGU56lp
e1i/VqqhqZ0KFgdIDpHdJvqPmfuGsod0dZZgHwgB8hpfBOoGVIUvKSpR4cWm4Q85+hsPCUOEaKNB
SegK3EyVxxaP4UnadD0MoKvpupTY61wj6DEI7ixNnRI/GntUMPAYdzj9lQyQ+JDUAF6T54H8oB2F
EPNJj4u6V/FT41M3PHokYjinMDVxeZ0wFjnY1gsxoLf3qJEWmRCERmYGYucX37mqieecutpT2b2p
vqOIwjsZmmSwfoCBcoWVTMRKRuB8WoBrshgO3oDUSd+m9cRSufgbFyul1nsaAR9TYE3WO6UFFePp
lwqnpoWWrHitbydnYXqSTYSIbzsCSwc+ONrqNp7MwYte1SgvnJ8iyEmNC8CAQv1Z6I4n/RGNB9a8
w6LEb3AFLBGhn1aNWKwQIcZFHdBnF8MkrpoezRu2WccQso/JyuJRWsUcISZ6BIIX5no6MWWBHonm
vA3GrCvLF/pDU1q5OK7Q8k3UmnuuHWg6QYe7dXmpMYHdT/VbU6fW/SUTe5tTk8LfMq47CCHZUgTn
WJDBEx0HZuv4GjCNphnDYFH+PFbDC6BAtBtVqt5SDXvTR4HlSH521KOstYNAae4bc9WBZ4Z+eTi2
Q4JfRP0HnuE8tf5h5PyZVfPqnuFY850onuDmW4hGO/OS6XxOAa4XANw4adeP2NW38wFAeZfAV5OB
cbp937DV1IxHubTn4KGkMUIWxoqNJAuC7XXVblf2PSgyYyH8IhLDcWt+/MJuYZBUSLmhjCtvqEkn
h1n5r1OshWofSjb9/itWReAK+U+MMii0LDzoCSNb6Ue7LcfeR+u3yRFbaahEhPG2N7wW+nrY5KWi
2BV/icyj8Iyho7qNCu3QPREz9TvSPTL82/5NjYrhYkSTiwueJLDT3IsfX4onwc64vp4hq/mdBVa4
WqT5vA/AUC5mz/0S8f8t855jX9GcZ3+e2tR+TQFwxN5jwp75m4IozBs4hpQc9eL5GqrvVJf0MvDk
FuJvt6BZfGSHWB0Np015wm/tZdmjfOpyTsi5SoA8SfqrbJ6D8ZMbhJTu4Np4+piJgjhTju1zbnSH
7aKsh1/vWvLSfC3WqKxsJ+M37aEP8z6CCOwmA6cVX/yWNIFfC5yzm+4mLkgQRQVl0bOgn3xPkhUw
wSU8dUlPbh3aqRkWTSomLjezz6ppQnuyGQhuWSqBiEXUHWGd/ZKZEnPYMYv2Eilb7qwU/CDKGYcS
AWx+XZH9WHbmXefpZfZxiJzBRnHxhgWAjZUdoGsF0pB3k5UFraAYSPtWCkFeOSONJ4l8LQvxtdcZ
oNPfbAa8nyLCzBeKZZXmVel3FrT0q73iOjf9hdOTnO25gcy+QCKxAc+lMXFzA4w6Lw89oRYf6UZO
vaO1wqF267JCW19Dn1MxJWm9QnZzGyPqkcx2VNgAuQxywpyYXCcFadLYP8DnyOBBceJmbwN6YDXW
fhw5kpiAJq5QfhDpcpjVpu3l+pEQGhIT3R1hwEW+W0tmuALhgiKQCRJ5PKH5FplG7+L2OXzFOliD
ZNKcNyrvOv8QYbG9nnXLc3WxRGvEob4oikgn84N247ideVlGz7OwB3XSSbu9Kpw1sKGSdCL/ti0J
SM/Pu1GJiXann2sAlSVXOVWyBNvdjODxVJSJUgNpfDb7cOBytkLaheypnsJ3KVcy5H558Ttarrqa
0iaReQr38uT8uoImIHdFH9FZQq71boHGKTa7aWCn84rIREdNy3Sps/swjIHo4vwTtJCRLcbS37RI
YmmH6SjymHwkv4n0M7OZvWRKHsCxYZ3krAKMjYP7ZYInpcGfK4O172mjDU4YWNbAXJnXiuEXnuKm
w9ozFilIQc6XgFu19clvTII0z+4/plsH0Zemos8P8PAf5yhkUwEYD8JbBvIHzANHzcsOYJLZNHy7
MQeTk4Po3vwMf0PLof3O2OxZi/DtY3tbhye7s/dj/qv5uQ6yZE+D9Y/vL12XVoErUeDu0uNVS3FO
3DtheNoDKt8SqUVNjoMNzXDDJCT5HjNuiVSfcS7cP3QCNkAKfzWVGZZ5N2g1TIBXWgttx7cezhgR
MjH3wG05un7kf+8J1LcFwwc9/BXPuP7ipP1psXzqC0V74CC2MLUDUyvR4aMQiE4U7W18u/wdzxnP
ZTMLnq3jvYx9z7r9AmB8p/3lVg6qaUshdTV4wHH87G2l07evRPtzoLm2wjSzFwDCRvRg3Oz1gk+s
E2KiwdObhn+qtDbSRe0httoRlZGekOQqiIFYZgWIh5xQDpkxf2q83q6lpyDfd1T/wihM+CIkFWDz
0D5uUoT4rS38MY8tSGSjiAplVRjnr714YgLOKGAJKyq/I9dRYAmT6TSAHsrSss8ZRen/erx/V7FW
2ImwvySClrbyVhurz46BpCGLKsGxc2H93PdN25OgG8lG/BbdAEa9fPeeMVIVi0OnRXvGqC6Nfged
FiI+Yy3DWdbZxTofcqjxCcg9cyr7mXyf8tncgrzLqPFncpr9gZoYZOB+Fb/5wbRRm9t2LFefBpBc
OebwH/TbAIzbUJJb6Y+NXcIDqAxlQF6W6gzTnXw9gX0x1eZIrY13MEQEmguNnyi2/2amsbAxq5x4
lGiZwEkBprgZ3fZN1k3H9eNNVBGgrO8219PpmvqD3+iG50udOmCPs72nIhx7CZdI0zw5JOvTAX4t
s9Eh2X5yLkb8uYJU4ajMlBkMVkhd48OK+F5RU0vBQ0tarx2AU9f2rTQc0CMSDJvqZmbWVAJkW7Bt
KL6xFvO2z9e8b8j6ma3VZ/X/D3u6ahhO8TA494R+GVqzOPlL3HHPyKc1mWHrLn+ro/hH5SXE5BIg
OK8NtX5ZKEthppPNqbjzvV/SpS2CE1faVA7YVkwh0512+bU0pZIhAAVMxj/1M/u0u+CuLEtzLrn2
qJiMfRLJBcl4ZUor2sfxN6NkVEBxgI/WWtCJJIiQE8rJu0vo8M1bdmuv4sVp4BWU7CGVAt6MqKEF
DuDb8xe7yGsIw23yIDq3xzLxkCFQVbD0uZajAgxpG7Nw1SYVZ2KssvIHi/oVeU83hgTY/D/zyCTf
OfRdoQtvnIR08rnB1HxS7hXtB3nfOqyZKllqRebSanysOLS/9Xvkj2u1xEoQd70aAbKMskZQHGS4
qjp2V7zwEMa8gB9ul+/ZGJScoHXvDRYCXaA6zkn+sY+fH7mhT0/O951tMNXcMMfIOCoWCxeaaEFc
q5rAbi7bBroQCXwc2hZDqRLw8Rs377fUJBqtHmMydDiGl65zc3wLq9q1O5UYEnzAvYyT30+cMRhq
jT+SyeIW2i5Nm1JqdwjKzuaeJnwEd1yQcv0L8u4KitJBtsoHwX/8GrTX/vFHkf+nNhEbyUsVVY6V
EHYgLVekb1LsECckV0mYOqGt/1W8rGbX0EOeGfxVjFjrF5gns4pkvL3+MEkaCy+0ZLyH0n2x0v0+
H013X/NmE7KPmNPlitQntPZ6EsrYt7Qu6dE9O78Y8MUqNRJawVAFeYzYPXomisxgRbzpJH6cA+oG
7Am1XZD/WifOgRqbXfueC7rTASFo4gRqByM+x44ObzLpwHKi7fKxa9TyregA/ylSmQpgNY1XsH2n
tzztQIoKtcH0r6RrYOQl8QP/Je/pq/8bPF/uRI2DCP8NbcGf8szhM9bDBCb5TlerB9kR4jOMhJE6
a3cH9FxUq584n/PgmhLN4TVezjMY4h5uCakkRn9Dypdja2CCLfQYJWGPLcgJXryAhL4fZYVLLWrn
uXdltj4z4mmm5TQfX8OULfdWhvs8u7mCq7W7grCY0enpvX5bQAzZMzzBS3JSLYxfc8uViZI8JgHY
7LGuRGkSfqm4pYnbEdvss3FiGYqbJFUdrXr+JCJn8uimrD/sCOt/vQsKw4pJR10T5bQGxy2E6y6Z
6DslsRrz9huenIeZWu95XoVI0sYeEHtgqWPtOLEtLGEpUwEZl4WGY2GsV+hrLMNDWHAmPRYU5BOe
Wfii1m4Z4FW4NXQ6jld3Kp5NDDpflrFTL8j0oVOzxKt5cLJXbJ0rUevTjPyEhAANBf6oz99MQorU
LJVf7HhO7vXwh1rtVWeKT7prgfn9Cgr23hj+pqgCMFhNlrdBU36clmpkR9sXQ5DDMbRCYBnmXgzm
c3QomJjwDbYfyngNrGdjowhPyzesvGJbtk8Z7rNdJt8K1vLbWuJz4IqWsW1iLZDUIWQWO91DaQc+
vNfNwXl0S822Jlo12KqtYhNLHWTIqtHoyzJYDODD+okFu0Y+c+1BrBQjkFTo0fn9kTVGxL50KipD
4Z2eUlHbLsakMAVOW+moQPA5Al7yWpEM3R7JL9vvHMezhmQfu9OW9v7hyvnJQvdiO8f8SM4iF98T
36cwTH9ZuHqSjflaqADEqOfbf4lZgVRySXVqZP3OezDNu7x7d5YhcQyHASl5qH0BLSjbQWkCQrfl
vHQwPU6JzR4yxHCMIBHtr+KP+uT7SlFWue7JsyZPsH74D62cLeELQmy/hFPubQRJARLZMe+tiBTk
ZgbiNqLtyRIg4gdTeHMCUKiz2bOueVGBXyrQltVdefOxPLqtARoKp5SjLoYlKD1syxxKfzSV2VbJ
Zep/YzdO9DLaGC8zYMZrhhDR6O8yWpyifZR0WA6fJTM9cJuUcp2ys8FNo+1fA2Zhp/kt3h8w/XQ6
Z0batyvDKpaq+hV4hWSUTLCbHNu4YhcqZiann6/yXZDD4ywNub84CdXZa1wjV3KNUVjZ7PoGwsVs
tdz+htxwmPBLSTqRS+0ttBi3pVXCHK7bxV0TYyF6oTMPfNHlOU8JCfqNOsFN+xM6i5EYjNPvMHWt
ggVIFS/QUOBSpWSgmNCCML3LgR22jGzcyDykqr5PkF3UI8dtiGsXX67HwF3BMz9fzXVrgxbpvZh9
Ta4CGDW9OJaxWy/1I1wRZST5sDzaaAalZnl4GLhZlKNI7+SgeNUrUauyRIECivcrj1LVb9j1VyBJ
8R3cy6MASbxNMVuLRKDHru41XMlauPHcyI8NkI8pzda7g0JRLh7vd7loNsR61qzkqMzaeMAchzKt
yZh6lC/Oq9Euej5CoclZAsqVoHzSaHfue0qO56ZpDS0nf2uBv1fVLEYByt41YbKnylvhF2u6R2rG
P/PjW58h8I3YuTGtKBPx1oyKmeHMWxxlFhIgtY7JJCayGiY5kIecrCE1NYaFml1uETH+pNG0fqrO
AzqgwHOBZQ8A1DuvyoznCITWfQQCjeLqaP6b2f8C1ZeJn8e1W5k/c+nkh+OJN26RBqIKBet8Zcod
6tTy5qycDk/5FJoX9w2kwINk09Tc9ZSdrwLHgK0j6G5r5p2JihO78zXHE5cXRngNhRjO6FQW2oV3
jAEvFABqkNk/vesLBUmRZIyEwUotzhWXJfIgry1ATBoGzxHc9F/cgF1BlgmuWHooU3qhOGGPQQ7n
qgk5pnh5pnlBlvC3mDsmovb4T2sgGutsc3gCwfTMxkJ35X9bt2vspOUxX6MebG6CckKzeRy5WmST
UqusUfqYMDD32kSjNagPGT2xAI3aQhPi+OPV2LTQrZo1DcALF8/1pDUBakGHvmW9k3M+iXt5IBAO
v3rthJ+38rgYGfc1E16f2ML3vOtDyxXbJUuFA0h4/ol3Tfas/WREhm8yV6/VoufHX2H65Q6teAmQ
I3U1cchIk1XofuLBXKPcLa4tokkupHiq9XSHKN8sHz3G+g0cOkpA/D0Pp96Pol2i2zZ0OPj0heQz
2kZfY+pTO5G88B/iLGzmKRCSmf1VHvkohdyQsH3M4dohbxarXFkW06kblRR1RF9bCVx/x7DVYW8U
2gzDOvEA5ht/24l8g1zsk0Tp52mBBkaSPRgaaLtVlv1rthuA/udS+TlqPcsxcoQePAcCHxLDJyz4
UxxPWE4rrms5JcmxCcv8voGhOAbpzJHRPhxYZ2/apc5NCtKhhpnjwZtBqvzGzYpTdM9z14nPoWIb
CQX6JOkbe06X/nqjsvNisTmc1YUqRghc8lmLhRDwkUR+2uOqNnueOopMYf5nqCzpge2M0QYEiJGw
eR/som2SDC9v13ZZfew9+TVgFzdBSlTdA2eh7Fi56Ee+1L6a+zaWigjdWtW7aMLMmZ1us3XaptQU
6096xIMgUI2uUdMLzG1Gq6d0vnFn6Ax68HNzQQBdDJ4zZm3axAO9iKMLar+Ay/nOWTqj6UOtHHiP
X2ojh00/dPyQ3qMf1N/e6P+UhPoFTDL8n1CJYV1xDFTO5AH+TyMagmNdInsptn180uqD8hAndKGB
6sKu/sGXmD01DInenbdieYonh5AQe2VhF0SaJNmW9bQKvSxYfqhBofQimYepIUb5Qwd50Zhk/n1r
ATeC0LKUpjbTrU04UKqmJwrcTsvzctJe0k5FYaNDOMaQsq/UJIj7tKyK11Cf3sb9CAMCpBV6Bhf4
7I30Q6lTBsMi7CyFgyKvpFZ+5d9xm0CPQ6mqajRsw/AbGjdCAWRWZhygVJm9v2J/0UKJp9geNtL/
ma97iWqJjIGdqxAfHosraEk219XyEJlZNfwRrs+VX9eKSQWi7Odu5xgsxKkqid8oE+SgW1ZF8BTd
Paa/y9UIR2OKlNDg6C4urc/0ijQ5T9KWQpE/jD5ZC9x8WNGFkB7JvSIoGVjseSzhyfytnPuWrY12
a6HmbDAIX8o3IrtJSbD8NPYaqpRHL1MDORl1XvOC9ud/yi5wDyfCIaYcbhgVJVKOnPbW4XfNPp50
pqGruyAA3csBaYmKpGeeGSgYR4IrnIJU89yeQA8U3vChEBrc+IhJMTjEm8lw42679NMmbZRTQsoB
fnP/czQHSGD/B7vdalCp0kfzcYG+M3O2TU6JZAVrdS1c/6XbhajT5LHQu42OtxAlunN84CSFx4mb
P7t5hqMjiw3pbbqbWRdzudZPMdP0JAWz2uDMRWgL0tpsagxhatQgyAXrR7nLr/TSm8qXQje3oBeG
e1csCsBlQUS7lvzpO8/iW52EfdG3my7mmCwCq8p0oJiYNAeUOKNgRPY1C0APCZZyVO1uTiyJenTm
MG542lEnwRdsyFQ/mx+Bil/a4YoYS8eupeempxVi5slD1A7j7JrHLpbLxabq7IspL99A1SomnAVg
AsHnoumNBgBgfIV+k5QyFo8HZ/Y62D0tCgMqoXjpQzzio0MS3VOA3Tjdd1Xa/VXeQTUqjBJQEbYL
yh7cLy9nTx714yn23ofb5gdM0ccI9eGF365ZQfkfCdmS5fQAlvHRj7cwanhYa3LiO5Gjaa6J9Ddv
Q/UwYYtrLIqfpc6FxuFPS6OzSLJt2ZI+ahquM/vxNT1uGunWvrDJjj88XW43G/K+k6m+nYgZUIpP
uUyiPW4iNB7G76PD9k4rGw/oJdnSVTKPlavmz5mK5DnU4DjNgph1O7X0Oj6pw3Qf2+cYqbalQP6b
utSRwTlToZOtI2ojWYZiINGSWSvJl8hqq3owbdOaS/aFhdY+gHwuxpna1f2XWnbaijvV0jA4LlRf
2PODCpiYIAQP2sXljvmnPxT0tdmLf03G6NQboRcXHyf2tlrJp6CRiJfYjTez4FqKpj/xSysg4faU
Fw+YvvBlhSuG4+ziHlFi5t5C6jgV86DVGW9gm0AOctbjHvF1o/O/cRlfueonCUBE/uZ1aLvYKHKE
4a7LDR+WybJv9qsoyyVRFGd5LXkk/sKuFpZeQOL96+GZMmVOMVXsVO0JllD1u3zt4ji2Fgr76tpQ
ctKT7SXz9g7fEkBJeg22mj4iQVg14b8KPgLqrWNVcVOgqodR/wcRGtgx+Hw1q9eOfL4la35VMo7l
t7mwoNE2gXIfigzWArUy5ZCz1+FesdOSZcOmsPoYnVDCxh9cQ36Pd3IbW2/CRpRGcql3gYhktD8T
PEWFycUQD1OtgW7G8OmBe7xzXl9yIBYgikD/esW8lvT+UtPlkyoWAOwERi7kthT6ii9YuQVZNgDm
dKqHuMoK4sg5Qr7Hu53Zlq63YnpXJKKwsA+6XBWT+FuRwcOP9e8hdqbFJbaUuQ6TPzzW+klKa01N
INmbgzVfp4Q3Bj/SGsN64Kzx0Yz+6NPuAKJOQYvGCYr5dwhIJH4nWD5GveunRsYYm9SXuVSQMVjf
2CrOkIqGrRA24V//grGznaaNgNAlw0xAxDz1yE+58btMRsHW9g+Vv4vo4AMwbMLyRjJTNCCQ2hsB
tcY/5opXzMj3V6lAnswP7p+4Xv/RQzSmMGF9vbfON6xgl19j0fq94otttygroL/r2DLgXLzsEmvF
8JorscWEDdWCmtTNLzm6Mtpys24fjvsptFlgjR0PTEe4tqfOceZh+8y/KoaLHvbITzJirWlvx+w8
TUIPlumT+RH8Wb19RLq4I4vx+pCAgs1H4G6fygBDkHCH6iDzaMpQugh/9Nx4KMD+Y/GX6iJ/1E6U
Fc/Bo0gA0Xa+93Ldu3bsOe7rcO5JxtkRSyU1BXmtdQLhArwOkIwqEPxR0LDZ5rLFtO4ArmqD0jzF
iOSBXI/zburz9aD7cSDyNiAt4n4wf0gMeLGkF8yPOpICxGunetq0dmcCx0ZHEZ8nkwSiEwIuXXKS
jND6uQuHGgvi0B9GQs3KhpCpQsmnyv9CKaVfXm98Y8nsRbyvetGRCpacdCmuD3Xe+JEbpmgX/IIq
3ZW/cBL+BcHFIsiQ874rO7zYexRobm+B3Jl1J5eBODdZkyfCCPc8YEtwkhegG/Pr63x/PVb5AM7e
dRAeFS5LxCkl21GZ2fDxJS1gGC2wyHV58SNwxyKwOew3XWu4XaPz/FdmIK/UXVG43OCJg4CyyZRf
ZFpU8AO21pR7YyFM0DYjaIg8KS6JoEu1J8W1b6NyoJmJ2L5lyhGfZcXYbzNnx/2QfsJoEGV7UdCL
KiV07ng8BQOdfjcw/0ooGRc/seCIRgbXcF+ubzmIe7h9BtjJOdl7/xS/U7+L4oIdi4wVlNSzxxbi
BhRTjaiZi0TTuiw96qzIZAPpEEGt3FTOK5Opnht9nceiErEhYXIDSNQeO+fE2GI376wYh3WcburC
RFVRVHQ51SJNs4mSZa1pyD5E3HG4sXKtWWW8mSZCMVcY20GgBsEQCi8gf+n8k5MGBbgyqX5ZmYPE
L7cauG1kwRqHb014DCN2xzBm5MuwWWjnbJ5kds0p9ZXwWSUguRjSbmC0JB19gNQsF0W2b8xr6QX8
Fj2N9T5Vpw6NMiAL77+5Y4FdMazSOloEnibRSTjfCPd2n35n0NBxA+GAcPS2yZbltORCNlbRXEVX
+ulKBsYXXapo85ErmUHLFcpQMNKnEABD8JOYG4LXyQ7rKHfPw9B19tmM1Ds+VM6WVsEES1fOQIo/
GTiGmn5RI7JFu8zN3+XJ5M6lkgfwE1hwCscbaezuwccafiU167WwYlt9huOx6i+WKLKFKZSUsWD0
MDFu2hlM94SVg18pMSk9z+Rw19yoiVw3kAtYeGvgF9s5UV1aSTIXcCUzQEgyYEuwkRuD+6XpBLbJ
1I94qvRIimFuEC/CTgigBMAta7ORU/44fJcveVcRnj4HAZQvtI//YEs/rfeISOHvcOJEpxA1FNkZ
IhlN1zqBfRHK4HaLLAb1TzOVRq5U/U/W3f/mKB6J16tK18hrs6SFLsJDnGjiwqtusQ9J3RvgG6cA
luRfd45MKaaJL7YPfjfQOsUwE3XIJMZhR12OSWjXtygvFY4c5jOtuMft4kIJlVEFa2AmQ3a9pJ6i
sC8B2Gn+vz19grFQW5ko8tmfR1sqVYs4raUY4I7nKQvVNlh1Z1v2uR1GZxpCfjYtoDGjV5klvcsk
c/htPJPsmljAyY6ipLOxoKWzSq7lh9mqADsRnLBU/sNm/oLyTokyA3fGwclxzaY8+a60nye5hWIa
fKSLL6OtFRpTzPJNKopRewhEuKT70WI96l8EZDamZz7Xge8DY3B7uF84E6n1WUbnwYHuNOfawmml
zTXqbwDZBEUy3gLJR6+Bf8B1QzdOGrSYHaAfYKUxzCn+nfvdpF85oQxlfrjeJgFwXV+5Z8aRXCbE
JX3nCDkWF6R5V4Kehzx9QHQJaOH5aPaNX2cxVFTUsOljE0y2QIvSy5fcylLgBHgkHkM4jXuYsgil
IcdU9XpK+7fhSo+fAbBup24VOR/F6WJFK6hbykY8EHRgvp6TEVoY1OeLMShj2WmvqdQE1lG8L6Vc
rafMlaTwkokgwGTyFvzqYFPKzBcPxO3Y2+rMA39U1gLo/RejER2bZGIoFocfkduCzRiX3knula60
1zcW4c0q79GKnIPlZ49a1mrHXyFwyS7OrDUwYuYtOIgvdhC23KpSJB0WSbAPfjmexasjOaMNPZ2/
AojXjpDap2y5pmu1WKQsAoNjDWVjEKOJazmlSnYfKhC4rwh0VL+8mL5A7mPJU1Lw4vFwTQUTMFxF
9rGbetHeBBEGXvJVoGrZq+uf+l1z8P5viK06c6HNh7a+IhOD4mc/Gvw0WDkBo5cYvErNgJQXzcgZ
QwPIY4a+OltRvKLfZedl/BmSmGaqNZt/XvSfslS9of4Hzb7+LBZqwISBpuorY8oGDcyhRYrzjzDS
z4fKp4NYxe2d4AEJ92vNw1430EjzhLsbmW8w9/4bhGWX2iamb/joB2VXTRjCoLJZ9ywNGImeQW2g
ZGKDy0P1OH1jT4rS8rt6xT2lWaKFDh6qL0YooJLoH9tX+faz/wRceS+CJk2oh/UM/Y9FihyXpj9G
0uyb7nuORYuEyF7fcTrNWpwxQhwmsQoaF8Mu/+1mQmHv8RMooGk8LsPJC71i+CglNAykeZdqtPpU
FHkna77ddUcFttzhhkixai08Gy7k2Zoj4tQW9KRMQFR2PLpzQSlMsus3nH/QkIA+aXNRuBtjwr3U
RmGGOXaamqN3T5Wy5OPad9iUhTU+go0A3u1Fpt4WK4xbjAT9eku1Ieg+7Mo8WsZ1gfo0yfG64pnp
XWyKx9jvFc53Btz77+PMoyKG/I1D1e1v0YLXgrsyPVs5zTUC/4bXc4K//Rfg7iHS6KDXZV23ugdu
/LpNI3/sK8TtORFfaLaEs5IbfEuINivBS++I948Qf4jAVrQEd2fq0tp73nGCXQvNWU0leiEvwo6j
PLI4BB0izb3Uv4A7KicQ+kR5C3R3J0c8lCy6+UaG8/O5c9fIn8M7lK//z91GU17Q/XuTQv8w7Na9
pq8bJg2YPwZjbZhAeuGiVpPRelb858ABc8kJhrTldhprL/hTMv4ezPhskCRhYUuMNHldlG3+8D0r
0UeBNKzL8sdjaAgooEAqVJEBAiMZFmokN3Phf6yXbVD3k2zsiD+dQHVQSNh7sc9m5fq1xBvSUHAd
pO1jIE1/gYNxaxks0LnlLhAt904+WvdWtwdBrQjMXUyGvWjLKq3loCQbL5saHptd8z/T/t7mSYw7
dUqPaDM3dwrg588oNgTxQa39E7ql9CTUjUZIN8Yn12FaPYypFV15S/cjv3ROu29ex7PRvQq7lKRJ
6mCbfxlMo6cPTf+xqkw6EGASTQYQQyd0DlkNrnM8ilbvPGnH+ptNFpwbr+vPwlcG1ogagvfNP7Kg
rhtgRtxpAXM3vbdRVqUWlsk/k8pYnihnZ6n9cOXhIWIstLYIpDcBJ2pcKYm9b4JB0KB1GZRpm2Du
kIyuqiaXNDN9MW7zoHuZMHJPqVADktwSFqfk7TGKzUawT/7oA/x3kba4X8CV7vR9hSn/AeR+FKTd
RVwCYbwVM147/LXtYRt0KP2H6lSqEMhqyNAWRibV6TwabIdcf5aEoJPBFmQjdrXPg3o2KIhsfsM5
xM8b7DBVMn9+k1gGKVQMkkrOHRNhlYyADF+yGOEgluzgOFPAi3TOY2tGdukOEuUqeI+QMk9hM5Fc
2tE6zdO6717hfr8Pzt9HrxWgDNeu533kuNXmfA6Ar8tCTplxrSxbqqQNtrMFTlFE6B1twAuk+pWl
S75ADli9fD+AAMvw9dmqnJubaGSBm6JAG6yNU/WRnSNV1p+e4OthSdJcSF/Q8hlV+8E3EQHMn5l5
VQVRRB4s0vd4BsJ+4fTaSUyDi1s1Z6qCEl9YvBOmVyH9gnoYK/tEad3L2O7QyC0oZ7/q0Wnh1AJj
yEYGRHYIy4+FMGe7GZA4jQ9h6Wwq9USgu2DbwtwsfHMSodbEM+E8fh5kDZBOpnpYKhydA3H1dP3l
wNjf45D7iXPvo16alW11pXgjvJOugia+RDTP/S/i8AH3bAaJyM8m59gX6xLmvRJuFtVBtO3LqrWf
VfZndoqd2fk21yAwZLhsimir0Z9OnRkZM5AZ09NwGirwlD0LqhfNcYK7c6bZaNuoGGAE3Zdqn0BU
D1plwZHve0rnqhzT/1MgA1lsEtlzIJLPUbVet6oXD+hxzDVZjj+o8da+b2TOOWg4NNi2RaQszv5Y
uPvRXatAgKPMV+FelU29qBs32Bdw8AnjXAZRS+RoGezKpuF1M/XwFjnWoBjNc72ZQmAP+/+Q7wxY
ez52ehZNVLgCgW3gpVz2FuxUMctBiXIMbSXuYJBtk7OzhFg0lqwwYJ+eUQsuWYEnJqSqaP+4m2aF
huVIi2ogGPNPVsOVDjS5EziiXcgZG2XXKGQTwSEwn0W0r2dQpqq6btxIsYr9bO6JzGvmNcUCY/yq
SY93G6TxJz3Dli5RNtwX4g2CyHQTat29sTMIwqaEf6c0DMw70kMGdFRzfFOqfdfRSqRmVFB9rtAp
7WX3gHpmeDu4ErMWSN423sVulvH30Hg1VfOefFkqXAHKjPot0CSOspe0DvxOdK07g+9B8xJHeVGh
4UZNpDZe6jcnDpoglr50mrv3w6y1pqeCb/mozM06VtHedaytux+ULZNGnmtHbHZ+5U3lSsJYzVax
obFlfaF6Np4SfpXM1GtrYrUu0kPJd/k50JaVrdtAaMljg3M6sLudQp4a8tWDLC8qe86Tux6sBIK7
oldqiHEjiS9Z69zTK3trQiSdB5Sky00LJKMkMmKQ4hqNp97T63fIn8YGvaF9MqYfiuCwrHWVN+ov
DeV01AS+0oEx6LhHSn5MVrfdzjgZPzQY+IBQVsqm1/vLeoL2n3GKmcGEPBBVtBwrtYxzQVk4W/Cn
VEj/pijRebK6uai4YAHkvKyHsjDHm++rEsMNVh5aepmvB6RlYps+NsLWQFK4CIOZQKdDlNDdtunb
M81GbziWz0TPgCYaTrh+3zE3DdK0q4DDXHTQY/S0UW4H2RIqpG4/gGIxRrdNJz+bBR66krImPcd+
p5Tip5Ji9WwYUUEurH/A4q71fjwGHeQBYH3BMo1nBzIYyBitGEAsAPK5QebSjzf68qoXSRgX3ZdK
w/qD7kPMsET9HuTbxX+N4W94/w1OJk+g4krB3Jckx5LnBoE7nkD2Zdkg9OhGP3b0Sc4NUi1cF1bM
25xZQlgPMppierzClqmwdpHAH8/T8ueCWd3OTojz3BxT0emDdPOW0kbivzBliGQ/dpuWSJkWTisr
idM6NkvqqgJU0l0wfaKpbNZQMBUele3cN83oBLOO3ZENyvOlEHQsJe4bGVau/Kvti2/jGBGRpKQk
gg3P58DcIgx+VZl+oEBY+dFhDwOWwBqDXATrvf8uG7ZcS1tstMJe7hhW9G1upzdx6KcNGqbe8B5F
JlKBMozm1McLyp/jdDpCFCAZicglXVT3XoYYqk0b2rcAkGWPz/T4RltF3VYFhf0R18phEnObCKxg
NZgizl4QZAjpu6Fha0qXMtdJYhMEZmHwQxtAY3OsS+Sgz8pkuZ6mXUctXPkv+RMbKfSM3g+sLjLa
rbkxG6udTKm8I5idaU9xTvkaj0X9OLhpJ5dJ6VFdotQrDtSbD7O/UOsnYOV6uCnBusc/GpAHgCWh
Xa+1X1KsH/FktYCYqmgthd+rW4+NNLkCpV8EMxrvUtz/lT65OZotYkD/7JezRh94bnaxZ7hlLIYE
PvhCeDEIr8C3GYFM7s84A9MW29MipvN98vgCQm6SKCNhN6fYIWaerd6hXetCstCv5VuBK/Vi3ryz
qYYv9XMIoIDRJQYN69pnaq6sriJA//56eV82PTQIPH+S41r3ZgvdYboPUdNNNYrP6UYIeMDGl9V5
BAQKN0897kbZKPFyiJdqCZWJutVkSb48KUz6/m9RRGN7TYuFjwNsBCeQmEs67w76OdpKwD9a6zAH
bDUmBi3hJDbZ1rQ4Ui/2cIFEW80zm2YvoYlKqxtU8jFP9bFYQe1TjGqdcoonKPZQ+/88guzY89/j
cn1wk8oR2G9QB61tjTucydD/B8S1fiXYflOdUULYVQu4+YzO0cMMVB2G7vbbJZzYoWvYOz3GSFQ1
nvB+wue8k1ww28qr3PxhPNMoycB12P61/I1tBuFLSvdXFtWGD6hdgLBK+RSD388QNB4pp2jsQaL8
LjcN5wIuLAQjjOYC8cyerrREaZxijdFT/k/3JXKT2RYyp9op7wYALmPs9NQGh2+I5m8N8KQiB+6P
QSxiG69s0y79pfQvjpcArwCU8xUIF06UNMyyh6b4uHwOKrAJzj5597JIDfYekWHJ9vDUbitfzGgp
0No3/SeZy52Gp2s7ree5hzeePYusXAKSgsmX3ffp3Ko6SP1wFQXbUnWLyp94Lf5zejscg4jjq3Y/
tLNewReswCcC038jcEOLWAjxnZ7t0KJ/t91QdOShj7pOrnudh3p/eI4JeqbhJPFGjv+228YTZYHA
lsp0aPN6BYCXpy81r75BpkLboxPDpvjjHL7sp8LGnTuXZ4+Dc2CWDYkwk/okkx/qDzdgOtIiiq0w
WIK/LrpNnwYyqjai6U65zpwp9dRiqHp85FeRVgoqcyMsffDYY/d+m78MN9B+vu8UteUSPwcFbuGP
eqFL3/v0GikszR/9wpSs0X8W4k3U/luMxnB4wSIsu8OGLbGxIdbYawSZi6DaEoRE5zL1iXJgvmmW
e0XPGzxuOYVOQKbgD2B6jpGAXdRonGuyhOKbbIT0/ZuJvM0mg0+gGQB4Jwy9oyHZtvhkbe0P+15m
SV0G2YJLJdTdI4UWPXK6F+5w3ibmDjtHiQbEZne+52VDs9WHcQbAZeTtP5U8whF5QM2dxvXYyo1L
u2mJzNbkaPFYRCrz4MwavTeaElC7IFLObr0ww4SUlCMrFm/wvzgvJjt+Fzv9dcwNTV0K5FMo3aJ5
bW9LGJO9ajwm9eTiTkFUP2maAmwnS5HkZ5/Ug7L/knSyF8fH9hGqBgzk3OtOS7RWUbnSe/M1xVfS
creEYDt7kZgNelKcdM+sGBRhBf5jCs8IlNa0vTk7hfjfV6KZVOTn7d2jVw/oWDBC1Euch0jKYJyz
5U7/Slgf32g4yzqCrGf4QXeGJfE9kQuFjY/TwFfwYdB9MrX8707Vj1lHvYA0oNVh0UiJhR9hdbr8
IgxLhiYMgShp/5CEUlGPVqN+AfFnGm539eOQ9M/yB1+YCAgm1wCD/4nnCCfln8oHqUaowmJJDWaK
GjfzUX0AF5YZieje22A+1vqRPRDK7ULv1Ejmj2jCDtt8+ug73NPxmj+36nWocodLgOD5mxPXa6gp
h7dEIS68l06EFly/rccqblJgWQwwfLA2uYUm9c/uTZtAoX1hgyUQ4WsdGf19OjUxRXGoQ+z/Y20H
25rp1K0f3OK3UmTd9MLB+24GiNKuJRFyIR4U8sbd4D3JdOyjwJ/WNWb0+hMI3463K7ZVZsUDz0kc
hnl2cICEWRdc28GF8uBpNakjRbVMQhPCTGh1ACh+JlXwg3myUZJj9UmKUkQrHoSzxdL3C6R4di5d
4vO6iIey327fa2fdoDx2pL1oMjG/BPuoluz3eoQi9PpD4UKjfOXA6UNoJkzKP/rOjeLwBuVinS9A
ZKKT5VJVMba244y04LqiX7Hj6v5JIpmap12uwA6sRM0/E2ZpYFx9sSvTEBhy2D4jxYlO/qF7v3Kd
17TUFJaX2ZGPUsVScOIHtkuCkR04ZQSmIDY1EBXsE9oHyxDpkHORGaw5hwC+SaRIn0FQ6L54GJVS
i5mbkAsxmy/HUp+B0JT0xwkAmfKvwuGVS5dhH0FKUaTsses1/shfSvW8qZeLXs0y3wiCah6FP75+
UYkHdy2YIJydmkN7ORUayqRW6VjwlNzVmCxxdAl6r9sKuSzywq5hbi+9dcOpJWgZxhUVyz8AXQtR
BRNDk1TX/3ta9uAv+XxYxrFzM8NiKptOY0oEtfQvNO6G+MiM33DQ/yIxS/s0XpuevP4jAeI1BvjO
ZrQ8Z01MAqzpIr75TZq7mjBwyHZl9AWS2S1/XKwwoVEr3mFOHyrcVldzUZfNF05MPddeUhRrc5t3
3LCQ4uXsLPqs2/c92VAdWCLZQ34tUxLGPV2OyJkecJHt0+ELUwphRfzOWCdDAAJWNOa2DaJWh7pH
6UVSUFaUOy7uKzJ8BCWn2J7GkokdIjnNH9aJR6cV+22972cIVCmH9hsHownQWk8z4dnzvq2cNYmG
8BLhu/zTyzNTZElnbZr9OEe6n1bRfO3Vmw0fuYIC0ZohlbiwphtewHnLj2lC/9FcB5qyqMUXMvYa
PXhW8DOim5o5aqWDLdHdoY/aQNmtF1gMlogw8mKV19eNCO4aOXTE86lQB6e5WqCBJ+jifBqHvQFh
VjdoLMlGelxuLf01uX44pj9y0d+sAHLh04/TUBDh90Sveca5X0UFXQSy4LLQDFpuhdJDnfEvaJ4M
1FqOJ9rLsrJx9zM6+orNLJ1CiXdbn1X02hmnn6oSO6Ei3cdLW1Qq0MCBW6drx5sJzeFVrktOFd+b
4wl1t7y4liFesxSjJKpfnJj01zI8GQjJOlZKBwUAR144CYanrTXPVycPjUv3B4IF1vKljDO2Q71c
Wd+n0G64DJhDCprH6AuYAeWjEWVJQf+C9y4tbx2CSURI4G4XzzdfH+w8R+8U3Ed+BazfNXhA6RnE
ATuUPOxHtv13bAtjdTWtZ39v+Endd7uhg0KbXiZw34sUIj8htIccWuLlQNTGdIQaDrlX01Qf4K9Q
e97lutMWfPTypa0prpTwpmB3dF04zqEAjOd9SA7Gt/DyP5gw9E8OpJuOaiFIcVxiA9tZ60ZqRrwM
YMqD74r1/UyaAu1qVEj5fsSEkUuSd4yDf3iCsMYgMgmMwi3JkOOOli6X39+rYYBz+p7Mm7CORHTD
IFJns36iLWmaKSxKhBuBpGQjHL3Uch9lyBSsD97F2Y2kgfLZddzN3+FZXgKSfnCRU95FrBXR1M5h
7lj9RKbkvePctUhjxervRbakPxWfUmAkX9iPfgtjK1+JtnM69TjLz2gxV430DB/ygFWEs6yFyQ8M
EQCAGxGyHKHsE1WKSMAeTlzRumRQuTSF5dCWjKxCpJbVGLfKBavgTw7K9ZlYOXqKFR52xLM+1cXc
pQAo6eaJdKzRpOuxucvElAAmZ+fSqn2Er0jt3MpnVBAzW4b3ab0ksKwWEg1Buy8SSDA+qNr9h5kq
S6zAEtIvUbKnPnV1MSZBGc9gDYvoKfOt4q0sGG/nnV1VYkRjjUdjcyjhj0O4V6w9M7W4gt3cSBqV
Rme79m24u4+Mvr0uHHVWSH7GmdoNig/oYco7wKd4a6xcm+AznlcdoGcDnS7KOXo1qjuKooXiYWq5
D3IIDt91psg0B5p49QoYCd2CIenTzMi7d2wJ0hna5NH+B1LJxR6ubdNUeAkD3rXXP/awQKRH5S1Q
XFqCyqZ0cRUBiQDWu7KyYXOB1vVoAZsHdkaYlFfUpTMndGiWAT76A3Skar3t6qR1SXwVzaKCP00I
r11wvNl/XV6ke9cbu24RBOGLjSo4h5fbkyWei2j1SZtK8/O4mYxGD5Kgnvx3LfqtcMeXwWXlegXt
upcUJ0FrJdWmBI0z8jS58t+vFSCVp4Xq70kg92JwpRLB08876wvxDc1Oe/K+ykhBBl8ztn7Vt49v
AiMAn22UjKtaSrl+mbQYEdxsfgCoSECiOlOUwcBE9WxZ/XNfvX7b7Ibq+4eJ82aeYwCPkim5A81l
5kXNh/++yvoedeHD78QuChNKjAzVJymNAGA4Aagf1y+vcFdoaximkdkryOZ/3tLiJu4TUmlXMbJQ
Znb9at0Jt9FKtLY59YoxR0VPPVNDyk77FZZgSe+WXEuUfmrvSThwnKjGeaPDhCaRPK5g/od7thbD
7tdge1KilCNP/anEbLQWMsc8ZY/8lY35HI31BNOT6FB+YyxxrtJSM0C/s0i0Ijon7iADyHUME5hR
kjpKKtP7oZYwlkC4ZuNFX6c7fRYVefgSpp0nIsBl2ynAxQlyMYE/qJbHDoVyWHKWdQ+AZLXSR1GX
KCPv250QyBVtOfdBFCREZlafyk7LhU6n83e+cO+5vTuRmUvHrG/F6gBsQ52dvoMBLLtzvJ9FgeXN
d/MCXKSgGGWzIacvXmroeoAHnZeQ270Lhf9IWNEDh8HFdFtNqoOo5vPLpZzaHAl9E0kGxXEqRauW
+95zXFJ0z73TTOCgvEb6VK7lt/OTBANHNlvDcU1V34hKZ3QRm5SQC0W5/52QdeMIVK0JsQZEJypi
ybz4nkcs8TIaxV1GZTWxKqBniCHVBFujuIjymXlcSW/nluQW076Jpz9zAyOnSrWbh4gM3X0YgK4M
FwoZxWNZPnPs8K+cA3WUEdStld9C8MDEByLYhAc8T9vHdO3crDMi9lwegNWcSE5LHg8y4jS3rtwJ
UsLmQpQvr/m/eBNoXQ+6CybIvHdC5EvRuRST4HmJ6g5CysVvvdUIVac6wgo7rqi4c85Ppy3DLUfD
U7Y8o7R2kE35N78RLPnXD8xGkNyJBu1AiwXxneIxOkVAm0KhoMjK41HmVRgHuVBZ2wDpKB7lcWWE
scA8mOEHdGT3KWq3y7kMINc9N1rO9m5UGvxwazItqX/2OwZ9zLK83hapuFyD5/XA8H7x08QlzHeQ
RlNCVqbnHRSur4fdmtmHSRuKdc61D6MSa+6kf3gOIHo4/e0Kpc5woFJhGau+lT+22cDK+AnawmA+
8ikeFvIdxE1zysWcoK+bjO2uhxePbBJ5Nq49vdM3oFbW2ka1EV3xQQ4jeTyTBtCbx3gxdRawQBCu
Glyi+yieHA7rCMgXmq5LvgO5MjgQhcajn9WepuvMwmTXsMu2f0cBUd2pMpCAGOSXrQPVCGyYvV7O
0W9hF9cJXg30SSTN8C0vkQnFjNPdnZjC0mjge2G20U1vHcsMhltWpV+0TS7VK0MnVQi/j1kxtV9T
kI5PjfvMFCGlHFgS84Q3UdSxBIl7AsfwzbwLwJe18EjCE4xI9qbD/RyTiR8FjNUdwfAmzNtw/5yx
FFyaRcV6DKty8KA8bIXZn3vIelJ5DJoc99Cnt1s2FoAzvAKBPqYeYdKJj19oaAe3zQ6VyAzJmE4H
6gWjePm9ubnWzZSO9KXya8rFbrItfTcEm8xVfz3/1sDmMpVLonyAKoQh4tDUyZ2DfI39LKpPqOto
1sWShICsFo1XI5UH3lL4mcrGrm/jywuO9MMEwQP+Fva3Rdg6jOUv0dLnvq+UQVjIc9HYIrQDsXhM
2scezEMZ1uAqNrjk34aWU/7E5FXEZFHJ8ma+7QMGaXViJPGd5vqLDzzSpsd4IyckauhzwHIN4WcC
WjStgOxo9j4lyYlZ10GTYzrfAvLRudDMrO/W+1QFugAzDgr27QsaD7vEJ/FPjUKfA539JNWg3Z05
o5vlD0euzFIwbJGVk2jGVYI+4eofo3oqNuYEYIGhnUXwInpCh68YXaEy/DvL6Eud1GRvCe10ghLW
XPaQ/weGzXoo5ADdzKTFa4n/AuW5AiN71g+eLLNz9IW6oPGrVi3ojZhQ1S4jFZZ7gs5X+HD5bBck
5z2pV9yyGK15BCMcjYr201kbwETK/73J1pyVzAYvsC1K5140MIlMFDGW9m1PEGOJgnSor/nGlWFd
PllAi8PNNPp+dz1KzhYmtCd5Z5EzJzCod+vtDOnN+7nCEdty58jpJ1LvECHu/MyqTTA3W/UFgPfm
fu032O6w5RKEiPA0KhQ2z19KPcNTBPfRio8iBF4QJdqdgiv2fnqOu08BuCEJvHLNtzjEjGV8v6wL
+oH6ZmJU7TBOaPHaB/anvfWUtDk2jcICkJEXgZgAwqBpoS4qUksZI+yt/VfP60EI43ULZ40hQStK
qW5/+8gdPxqzmVQzvTYWHG626dejNCrN2YbBk9PSiwsiooEK+Xpla/T9dwKS3wRkXRYaPA4ucRW5
1LOLypEPm+IDNNFD7lUMqSVQ33ly/9NArFrQDetmGPnfQ5j8CNj2kkBqshKX/hvo4qLwcN8CRj9k
wDi51sVLXxuYjFqiJZaqV2nKX6I46mLk3seGcdHnMMqkcxsAXlto4MmoOy7kHE6JDAuQSDbAKCME
7ArzO0ZyK2SJ2JeGBmA6OYyqtZLFfhRCwm+Sfsl5c7HM7gxqaQVwVVrx/ZgV+S4oT201KXhbMy19
2ue/Kcn3NR7Yc/6iUk3g6DZk5E8/Hk6S1IA4gWAkik9z5k8cWf0pX11kf/lsO9KH7+jivEQ2+P8N
0pWuEd9ABet/8KbBTd2T6XV/58VEi9/p29FI/EBJkKvhAZn7yt/JB0+UomqlTjItlKvwp/kjxUy5
Jp31PlDeJN1htI5m5m6wrMmw27VJGjBWVjoNupONmZMkOEFKpTqVBjmXgg0zKbL0mNaQKMaFOSZB
Ypf1uPGwxM4z+kDdwYP7N1xyV65pkWn1LarhoZI6b14Z36w2PD2SmX4R2ljcPVb0VKh1kWQWkCcL
fOKKudPxKSdp+NV113x1qqGA5Q4IrdEKhdKBMZJ1XP3d0qmWGYLsZK/wP0LHtxkix78zeTLgMaqw
WWGTftxs6KP4i02Y+L05Jzj2tOBWov9oBRpePx2xq5r+TYqFFDrUooRtaXn6O8ITMbLKRni5VqMS
MMDGbIk1TZPJpA/gAtpEzBvP5GKDB/UXL5kpvRXtgZdM+lLnT1HF0TXDViuvzoZr+uJp5Y0WPd3W
bEPmVBtdtMwWk61yij+6DZ9YinYMkN07+LtPJseB2/h4kiF98vkgNaUqAczyac2JEggf3M1w9MGp
U/JqzjNFiPhVzyLnHJ768FFR0ucnasX9Spnm8wNPjo6h7t50vEMWr300zljpm5k47B1vi2LhYW5n
1kwW51+JRoXWCUv64e0OQSaI3k8JKo/0ssBypcgb3KK4R/2lSOvjOPPJ6BmIAWlv4OtfVLhtvHNS
VQzLX/Z96TQPUlMhpscLfMz/IhrgepJm3XkouWaF3fBG1wmuztjnfWa9OTLWT51eF9ais2qVzv4r
PKk5+uyasd8/YUZag5Qp1lYsE3vQvKC2DOYVSqNzLnxWxTzm0soQF018jFlpLqN/6FSx2Lgxyh+Z
G2WQN2FP5x+osnv/XHm6ZRQRQBFyr8xLfsv9BGG5K1sowtTuqi6kAJiI7e0GTEFROPybQxZc6lLU
f0Oj0OUd6e0wRYl9CxQhWUyTJGy1QCu3t7fnxf+eH7CX18GW+iSyN+hv1P3aGBXjCnq4si1MDcR8
9hTeq/K2U23toNj1S+6TlgbZ3AhMHbjhUrSt8knUtLp9o8fkebXfzM60o8mtOZdCnwf4GUQ8zaz6
7L41H/CZ4qC2pd/ei7u3NKuBNtmlye9T2UzGmnK4UImUrQpCxYJqKX3uoEmo3LtFlBUpsJV3+rDF
yKxkpFWmuGQaRX9y8z/pX+w3SaIzlr6UJkjlxm0EbfftElRwJVFXR7ccAF71zegI/IM4QxNnW9f7
CWHWLVg9U9ROIztM9Ikgj+jAKv8vYivmVn96Bnsx8SPkP1zxmCtT58W/u2V265ZFnNDWdz/yG4cN
b7Zo3oIyNBEAyidSX7QS1hTNy601Gj+V5C0kKjYJaeFDnmAch5bNfGIIBv2mzjQzwHF455lTukfn
iLz1icBCwygi/FMK8BeZZ+WEZuj6is079NWTPTjx2HXNNedl/y/+4U5zzDsCxRTrW+zwQP9GqYMq
yYlwtDzSe5JTHALilX+UpxDXzPidlUlmd+lwfpq6tDFaXzQdOWr6hrOyC3Q+RcYdnuwlRUA3LWn7
wab+c4Ne3r880kajRJwV3rRezZtxFzd80Z/DN9JUibfEUniagu+wJ5mkXPVgWsL4ly1LWovbCSc4
vUV1JcKlWegW0Ld7Lkf7FX8SpJH/zc9xT48ijr2750Efc9odFjFv6g5qsP7y5LxF9CFmQ6VNF3Rr
4vh1J2UEbGjGSENuxYM9AKXfel/+x/8T4B3BVpNRtnCVUYwp7UkC75MTiiQnrHoDWcprTPW/gOBi
hIH/PlgAIF7itG0Tb5qs/N04h69uoMpc4TdZI3ACR+YmoH6cdhk3YGd79Q2koA5DMy2OutykbCyb
NPftnM2GjMmj1XxFqQQ4lHYK3SpDFUUbvRD3wvEzumA0I52pWoR4DEDMddCCQjXOn8h4mNf+MJmZ
Aa62AV/crg1gfZoNaRFmOIhwnXaFzWQJtXWGPl/yo1qlahb8qPQEoYk24EwigeAzHkIDQsFFFYtD
1FibZu7DyZJWAWCCW4bggFF1RLSfSrzZYHr5rbftr46ltP9Zw+gHSsdw8pvS/1hb0Uc6McY1TjKM
e9ZryN0q+LYqae1+nV2/9VUjn9wUIbtVA49yDSrq4BbiwrQVZ+Dd/bEzrHkeWonZbQnReAoGpr5n
8SBtpVzEzr9+GeuFhd/REUbIWGw1T5eSltbmQ0nLLkHzj6kzIOEiXajSeAUWVABpFstXZOzs9vCC
k+U9XbngJwuxCBTYVNLQFvXitmyqQl7+lzNBuIdnspdIQAEXtvqh1bd5l4aEhPhp6STt4lZu2KLE
bF9xYupEmU9IXD6H266r2AeGOoJEwnRT41sN+83Re/oyjemO1wcluLXW3cjfnSAWPwDWu492zeLt
1sTkMEU34kdIy3s4RzhLhYIjtsHx3cJxpnCfHla1qQGimzLZpK/HHDJn+Afv5Z9/sonDixXwjt8d
y7PZ2B+7oyaY9T2Tjy8BZR0N4nJdGaT6xAjrM7xqwu+UmkI1QRW+IsQX0QMLqDJBf8bOej+9FeGD
d0d4P2quQU+d1l0kmewuc9K8GIaxhQrVA9UqBSy0kbIx1npz4cUWvaWMuyVpt9LhtyL9isFxr4ji
oAn0jiy8iJoDi2cW/TiWVpuN052vbfQhQ/5A05OcU5gmlkg3WA9GSwCchNIbVLBDwR9p20eJjOmh
0W5pbUhmbzy+/CS+MsjiVcKN6GxN1dw1ZwxsUK04ZIqmYGRuknEWXdAmB2GYSMyyXK8y/dVojrBA
EAw0nDnFgFL0S45YMp/4uZ0CuiAMFCqZHo+mXrnrhP9mYTlVL0roY7cuG9/ZBFukdajtQs8OAIM7
7JQ3jiN/spi/tBCR7gtXFCD7ybXfUmCWEy6Jb+4IShdEztHFhzwdhXEHaDWKu/eoBzIyWsgm/9E/
k/kBR9yBpIjyPLLL+bWT9Hqu4/aS8k3V6aDOCCdUsKTfAlSce/am1O/6Ur/R5d6oXZOWtVErzA1r
CtPFm5sBG4rYJaPWKn/ksNuCsMbWp+4wi8KKf8fbIR6pCPb+xJFro1tN7ksRz7Wfm84W7WqOTlJG
dUg20uMCKonxCxQxDaTjMbNUPKJ3HzdOA0qv5uDLJHBnXM8Jy1zaxO0Hdh8CYmOWKxBNt3S1kxdh
83MIKgAMVbSug7zdS5L6OCbvcwepiLb7GcUK+a9Sm4tdsocw7o5crFu69WwQeFMBVJ0dCvd7hJhf
n2vKA29izpq0X38ZnEJmf5i0VEAN0KDMAZytMxXvZRnq6OPIC2rEpjRdKeiapElITcw5TrTqUExV
+Llgl8hxqkcsuCSnJXqhbWZdI5LD3hjO5PFHAVhopJz26NTsrxvoBmYfdtevTiLhMA0QhdMK+Qax
LgOsDg63fRVBEy1DdE8EaaOQyq0pthZfNDMRePaybha+trsKTeoOsfWtFDJVTqZxVw69W5do5264
WfiyCD0v9RDMONx5tCOSgzWrnTntOCCADcI6hkF75tjS6hC8VS9KUUbkNpWuo6veRaKksG8xN+B7
opAJNr36gXHHbmVyJsD9RPXNHMY8zXzYQ204ihbquKQX/99V+csvCe86/VrUhr2LcX5edNgAsNw8
FsosopWuJApNS11K5FYbCVNEI9psd01TKN2ZXUsq5UbIAhBhQI4GZqyYMMTt8cAnj2QOMuC5PW7K
kdDHaycr9CBCKyoCUSYxXeVRMk444U2AyMf0ijYhddqnx3oFoYv3sXBYdwhsCLXhGHRbb9zFeRSB
QQiYBtMLaNDXqdafFBhcxy8o7XeJf61jGgq9sQ3FkyjuUGw6r4zugvrsVxz4Tdes8qA811tSGUJT
EQhMJrlzFZtSUkt3Aqcc5Afnx3a2iW5eiCOFkH+oPhpKz9F5//OqIkbqejipIe528J8vVHoWWBX/
m8B5uY7M0mHRz/0meH8ENRBCCp1Pogd3ZJYE0z0KKpZt1F09jQ2K+IKiPdE7q3PY/3imI0gGsV/N
xZFQlSvjy2S7LawzwoueVhcr3JMBJITNafWi3GSLWwS+MrXQ7xP2TUCEJnD+9CO54ZHR8nqGb25j
2acwy5IOwXRwts4GFeFhhfAgA/+H7rXhR+Nk49uVDS1z8zNTIl6b3j70MyiQE+LWS2lmDVoe5vjO
glLKQ9I+s3q0YUUs/z5BIWs8FXetJEF8bmsJO1zCECjQPDO0wKCOzcsyxIf22oqTdnw1NkmguQmf
vdFf6qkbSIP7k/WIsthVGm2hQGqrk+FW/bkRJ5apSu1WRmcl76gN6dSfVmg2Kle/ABw/xNGfctE5
yzF1o4MUfFXiWrb2b8BDGNv3WqiHn53pERjRgZ8MN6YwBlfa4iAzO2APpek4JH4+OHoj7NcMFV0K
BoduAwZP9ONH84RFlnC+f6QbLjXMpgvglWVBE/1hoHEKxUMl7GsJEmnYrRSJIzIIQK9D7JrtlC0R
k3gELhcg0ju08LuYJmDpQr4afqzkNan8fFUnLqIkKE5v1+aVurJBpT2TjpK6qOqyty7Fn6QHkDnq
OFOjeKniNHkt7JKA1WwHoE9MID1WFZZU6+LFjYEUg+aRqxZxyEg3OWxBf+P8dkN2Fw4pMurl4uXh
LZwQPBab4lGlL5wHTJAVKgb/sV6wPgPGghNL/arVqxo4WWeXSV6f2uRyFLGVzrVnPoSL65D6BHSb
a5CcbsqQJtyELlPYia8U/nNB2/UTs+soaGCrGrp53vW2ADaZsfDFJYkEux1LQB9aFHszzut38MAh
0FURCzGWSzkwqhyg2YhKzxxMHYDEJuXjaj7/3ai2Q4wgmCnTLqgDgRO1mbwLguWYj5QzzM1ot2oz
t581E21nX+0SDIznyLjinxbpg2KUjXgrpYTl6BfqoVb7F6DcbSyxRP9rgNlzLNwkXFYt1YHa/hCS
imVBrLQe4bDBnbTHYJiAdbKXZn483cfIGV2mqnauq85RU7uC6vCmRfPDPHD2K7jhLlJmZiMpgFGD
sELLGec+ZUYaoSh0iRP2bemwChGzme32mh2zfzqkbLsrBNuhTaiFwz0BiNO71Gn7Ya4HN6l3/Zue
eipOskrX1TJufLk7Iz378sLyRhd4FXsolq7JODcqJ4rIJQw8qBbKCtq79AuG0e6Z/92xuC7DTGmM
2J1Oz73T+swC8ujYxPfCZkO9AOg1YHzAXdT28Mlrt2I3b5TYST01/IRm5Qx58cJvxb0+otAlZIJ1
zAcLvf3QD4ruEPjJXMtpISG2Eg8fP4FWe7G8/TFYn+zFl+VL5mvBehHQKOZj1ZH7sy/I7xKUfbsY
lLq2vE1PL+k7AjceM8DzYe/0KT1Ns7PvTlM48lNSLaEiH37zj1Hfqxg2R+C4He6w7a6j9akqY7w7
/WGX/y8kAVVQ9tFEx7Dk61kQj5eSMOCeqneWKIlT7e4xTC6o0MymbhDQIEcKSKFRkFHXZP7kOgE7
svCSYwHzLAjBN3Ne0peFTbDAN1ZpmLRcOUF7GyTmCPTxjwV4owS/M1pf3kI8fgNkLQXU+NPpsMdI
io1f3Q+PISB/LVKdmwA7bBwawKsqu7tgfKDvfw+nvOupYp8mZhMNbphnzMso6GlW1FA0MwedLnSI
wCZMVacEfz/BOrDB5amTArbkKm5RoYD+HIdCeMFnpvb8V9gJ2omnFCXHP9uCNeVLq+AN2DfQgo27
DyAjxrZcf+sxUX9vaBQAt/0+l8CjIAzMmtC/oVO2QR/wU3lj9Af/oUoVPnwgA9j5IY/KI3M9a5va
kCx2cD/qfRGJePUI40hz/+85xUmxdFidGMkHX8Cd+L4AfHGoGs57jyjARPl6x+W5XHy5tEQ1zZ49
0G3coTEojITl81Ki9BafenHRUe4eH8L2NRE7xQmeSZa/NhzxPwE6JyQN+6DvAFZ8tcODTK0x6i3G
BvBWQ4F48iEZvI8rSSZlygNaXKrDfLhvPPOBA0ISMmI9d9NsJOFgO3WsDPs5xn3LzSDhTLXYoYOV
Mrr/SnqlwgSFT6RD8O5NNKcgJt/hiQVQbt2F7gY4EakLtXPPaKaa57SzmUMoTalq6ZNATh9v0Nn2
GvnuQCm1K/PG9xIDXouzV8a0wpFXRbCyj44gtIWZ73MOx4ESqEKvVOvJLjlEFcA70uQSXi3kX8Oo
49kmSUv1xo0Ll95F965qttvkIsAt4iMLhzZFgS5p38CjaB+xTT2oKlMQSR+q7h4T2AMpVxdaVk7b
E9+4OKigj/32WyLfv60RQnC3EnBQwqykNsQZoAfYJ7L0U8/sJclihdF84pvdeelf/0mYE3vXgfDX
U/VRCTfkLcn98CSzgZp7hALkX0MulKRmuxFdJlg/fQhaJfbOaknmnwhnixDngVhrXst7JRFjkpv/
/2yJBYetOIRKmymJBtzHeEab1GEEkS/nvNhZnyRXXZGx+ilQiAZ5JyfNNssazXAahb4tOCBMz8Bl
jpcN475DozS3HNVs1Uak/M4wlX2yGXg+uUTACY/2InHOto2Zl+T+C0WcekKlxTgj6JixrmDRAk2q
YxtmraDGv9LyDLqpGCSt7wh0qqPx7nFwWi212bgCZptHiJKQFnwfSScpULXf2lQE4faVE/dxGf39
D1dV4TzkFeNyIYUDmMsT69yS7JRVEswqgyegkCrY+GXc7qo028R3WNRV3h/6sLXd50clN0NnU0eh
vRo3/Roc8gbYJrSGv9zr2Ose5zhxi2oT8jneX7YsctHrElQK3gLDn8x2TwVhFkdqlsdKsYo7D1HG
jrCqsfzw+HByn5tR1KWQgdUOMrC0xOLn4UXPDk3n96D1Lm/pX9wAZ6n9ILwdYDmvnbbAFU4mjN4E
89qYnhaahAakNoz3fLOoMhrQp5ofetSStk61HGqb27gWld3xQJ94SkhG6hnAuqa41HGviqzFZ+u+
6QNT8lT9EUvq/Zfzcan8vESybHi33nVonmNMVhCqkg/ptp/k7LNGBBmPrsJuJCu3n+zjVUr88+kE
ig9IqIL0SIlaFrlue2/A5L+JP/pagjf6w1WlDj+zhXQoTaKP/59QF6XUHnSlDeWDr5jtgBybjWh9
8sKsrbAldFBgG/I12Y9OBeZhUQeRRVAnx852lBU6oIofYuSqRkRpOC3GuGBvpA5uiBV7M42eXmfk
ShKHqMP+2pf7JPLLDJtEON7IFYDjXW3rP/OwTe6myKSvR8E1Uz6JeWkpVQRIJg+ssjmR49Mpeg3C
lOxbCvVEhRGroqJCnQH9b1m2nft/oI+EfPTEjhHZ3al9+jxZP/J4gAvLyDtFMEnI2Q2Sp/8ALTTa
tAC6W4RvDW4SenJ8kT6eZTrZmrggK63IfJ03XmherhCK70R6lY39iXziQl8Eg/rQcn7LhipPO7u5
eOUbh6/aM5DwnsrDw5P+HQSAPoHRboLV2qc2L/DCsVIpz8wQaxyrrwoC3d8R1KMM9wcFQXeLHY5F
+Vy1vuo1GOo6XGDV8nPMa+nEhluuy8/HczWdS0tlRllXKWTCVaHQ770BgXjvY51iBlxMYK174cR6
TQYwwnXZylCUz157Inn7R9bP4hDcN442boWizwLAvnR+co0sv72EAF8D3e5zwWWxyVD9YddIDola
9iD+KDRmoLm5qhj6FtmXdJOUF3USBjajp8dgeQLqBNR7U4YlUdisu78cyca0pbkGjKYdCBmIeC3h
sLlPraNFu0BLw180cz/B6laQ8ZuPEDMwsrvArIN8yWmXyJt+EBZSkvRP9iTUTV/xfnX+v6fnh5ua
dpkcnviLlWXphCzw7xVJs9zzk6s2p2eqtFyM53n/Z5Tms60mywj9I9Zaq5hiTynm/+w3kZmrpMCf
87KzK2Zcx6w3EyHk/myl+zaCupv1aS7oLAOppkLkol2amxddybIms091F3uOSTX+kkn0ON4yLqAl
PAEOOs6m76BNynv6ZDA2l34QZJKg3ttnnLvazQ/pr+JzpbXCu285+1bMOpJEqLc6/EUwuQ8sw1p1
GCk3/79zv35gRoG7cpGsDJk3et060pcPw7Kv/P3ZTPtN+4OZXqMmL1HGaSSHTDRacAgRUGdNGXMc
Cuq0lOfZQfkhL7AhtzxBICUtEl1Xyhzf33ayXzJU+J9EFQAqPk24wO8LhDgYivAT6SoZ9ODaqyhw
r/YIudG8xJsqFAAmHX8fGFRSRTraEPGDcU9BBuCa+BFki3DKTPnB/E47GilhNBxKHk6E6Ez/MPAQ
ngElmlTxqW8jsAuI0tnWzY3qsoUol8IXvBrFlx7eaGIkUKcW7iOYZEOhJ46WdXtcNRFwpiKdF6K7
jYC/10hHQDHah+RGQzmOeZ+Wyicv73d66wJ+Bf13VtGMzKQuNPPedTgDaiDe/xEkiJW1iG8hiS2G
54G9hl8lmEn2ZnBh922oMI/uvZkduZeMNVurvpn+4da2TQ5EF97SXDhRudzU9Qj+vj02mHAB0XtU
ak1S7XvEeOBr0A8Ot/5oXr4pOy5rvVbvbCaQ/RmEN/fczphyv0l5FoUrF5zxF7P5bdrPkwkI5W9R
/WHxtCmj+24DB48lBsQ+/nhCWx0P2IBZSqW6AsbtPZphDTj0I3VGF+HiGJTDqlXylgMNeXPAW3Wg
rLKGernPUdV13yRggAGEO7XCMuXeYY9X18nWlS+Nc56CiOW29G/pgze4D/PZJnonihXaC1gZWSvr
z1e7+q24vvxVm9CQAzFZdMHWkkbKP/XSvrJ1cewd3tr9F8DTLF81JidGVpTW5LhzPELrmp+HRLXt
8TgBAGQLpwvziGhdkP/lJ7c6mdqSUp2BuZbL3Wtkj5CDO6wATGIj0sxwBykrk4KpVnFSmOrRtY2N
TvFSkyYt/ey2ogEaezbbOna2N9mU/27j5iwuMQIOJKZcbVMymYnkio+nKsBsPzdmdkPmGMUnazfj
hKahgkQdeJOh6Pr6EihnGtcDyT2vvOMQLhWDU11xa2G+fREybChn6xNuYXGm1JglbssriZFaF+Yc
0QK/XjkUPr7X+CWGUQ1305vGzSWGo5ptK1CnbCzf6LZcj1AK416bYdoHiTYfXmIc358O4dWJojl3
jN0RW2g3ebk/aPl2Z72gXgnbzouEmHYG4T7+Ndank6rJNwEfHyVGHbg4xPyqPtTYktEBXfTngGzS
iS9MEUbHuezhQ7zcOlz6HICeaYqC+nBo+ZoMQbZFmWwK2z1MuFkVa9RlIU5SrsjSuFXoJbFTjZ5x
8X5yXubtXGSFSfZ2VZStorxXVO4iI3Pa+04oESLI/nwQUGMsC9AtORggMdwSQaqrIo5ntEb0xdcG
wqRQfgY4SEWGO9k5heV1Djgq4f96Q3Hv5uoJa0eeyiizMZV6C7dQOFCbGAqgCRB/6IYyi6jIucKy
lu9Ji4fy50NgeFEWtkNg2xMfA6SqjnQHAhW7Wy2VHvZSpoK/H97cL9WttflUAYYL4VxPkNeETZnF
FJwFoL/RpkKMqw/tFgewaOHVJvsPmEjFEmk9+Q/Ymc+xk5oNDsusPWA/IX5lsEHVGuSno7HOwYxH
ROc8wmpoxj75XEGxgiDRr3C28+WIPaH+33Uq3LLAnQt2K/Re6BwooIC3Rx1k9kRbZHHkekyArwKX
HdKtfYEG4xOr2JzE21YguEmQHCWpZAd9shCRz9X4tFeCQx/vkr1VyUqmmXA0Aikp+NAkOeJlUcCB
FLT3zsTvvzgxMzmqEI/zsorU1cX0Z0Y/aDNU7APgTWSu4MgXueKSvoknWialU5TtFaO1phjpPj6a
+N1GHDddFbH2QbaMDfXh98GwYOYYqh6g9hc4LHYCHnyFzoEqbsS6klV4qQe+gm0scR2coui1uoHm
68OtBLvhFGZibSPQEZPWykba66FKoF6Mwjnj2n90kPIvKVJ+KlFjD61+NmdGreTgIaadMW0TgT99
C3WuaWdJyOSCjgHWpQATAN/AVLLogkNP7P8XKoDekfOggUuGe/oalgnDhgujJvC0ZCmsUVuFeQmm
qCWnJGDTBHzFEN6VhqX6rN1bXroE4e0TOCktLPmYXq85YFNP0pupMNCIt/u1AMTlpTR+z6zvqqzk
24GpQqXmNrR2FjZdQv651e5msD0HMAo1VZdhddv8gROXZu61OnzJt8OkC2qBjQig0QQkW2UNP82n
iZjd1OfCvbMRO5+YodwKT4sFaNl+nNACifOj4Sk89MAJ9BvZ7nrVdk8rQCZEzqBByQHBW9teMnu0
lifIgPO2yIQP4cyFd4LgjWZ0ek0goS16mTtIj4tbo5GSJmdRoCW7qrMqd/t2IdFtaJldMPi3IuwY
00qKocYoFVx9Ls6noNj1Z0ypEUjtrk8JljO2ButwoRlpHG5qWaPWQnvwx6AORVBcANZyE6JdHweY
Bqy8LtvcAisuZxQAHhTGV0t5C9x8OmimNv0e3FQBUiGPwhncqzliM4sOlgXErKHYlhpB3N21Y4He
FvPtYDa2Jn+1441uyZxVPDpCF+n05jzb9kYZ9n/1WekimEX4eoo4vkLgh2ieuOPbj34t/OHCxm5Q
4Mg6JMvP+WuJ9AGrQvCaXEjEsAurt69sp9cav7WMjwWvvBhkyQGsJh6JcI6Kwbd7qgpYcYKy0J/t
SspsRm+ygIu6Mpe8S9IZRQH579bdtmB5aMUhFmxTQgApMxylc8he3joTX0c6HheILvCrP8Coz/As
2A45wfCr6zfi+PY5yTbDUTN5xLWnYldfIfQ4WnDPRYdXrdCcHR5Z3tMvB5WZmStiFHkqAvdnQHuT
zheFWthyqY5VPI6bQb0YaHif/K5aCyhDC4FxXPQxqu2Bdo6FQSfJ7vRvMlPNnN3OKsTSoCoG9+c6
F837RwtmFMgKIMp+fXYKcynRqjEAvDrkLtMWdOtaZKKFmvvnCXkwD5J+to+/vc50ItkJBd8oTUdv
2SeW4VczcIGKJTY0LM9I9bzdrly/MPtpjKvRKZK1QENj9gdwkmuZ1ryscYGLOEb3SqzArGLtrUER
IaLbk4x2OR2Mn85U0MRnszKN44Cb0q9807EtPl0s9nQRzcgwT2rEshsoNbRIMXBTeQfJ3ffyLOHg
5aUp8pF0M6Mm7nlQoMZq0XSqF1trlG5s1YYOWdUvemM7GzKBAvxiQHqjPNnVVn82Xqgkky221QhC
R/M900eUWUYEfaLuj1X5U9T05/wKJ8dVQ1Pyl2ZSQDy+9PpK9PnQun1HSGWTl9fA3zrGpdJfEtIv
ClKA15DS1Na9peO+0YUtaNWpaE9kWZHC+lmX+LP7R5fhlX/fExxnsjFMhWTkh0NqFKi+o6g6d0Yw
bT2cCmCZWpBNjmc92GeM9MPiwBHaU77gMh3WnWczF0hNzRPbEMoA9K2OjwAPjHKzM1G5zn3wagTR
0cvmBO1HoM6tdCqt+1Ytyv9SLvRdy1zL4L4Vx7h5Q/BEPyceSoaUBKuQ/bUsYom4l6l5yLD382Mh
FZZNmzljSUkBCOc98KIcPkKMIMpMRycjHqxIT4G0yKqFwWDlpDnaOn3da/6+VLeZNAXHQNCtnxRf
gy06GASwdD8AKfXVClEqgKmvJfN6b8m7ZGCIL5zubgxwYz4HUC5eEmZ29gPsZ95ruwlr4En3bWWa
OmqlQvnjNl09SFVpBuad6s9OEqKHXb19I4jJwFyJkYrS8EiC058kRuYEW5rBef9Fzswgx8uOu8AU
tI10mdRGX0t+M3sSt2mDzpY4tBdmWDmlWdryuX9qCsGrX8ur2VXr6OLDr/Ey4AQvXg4c76erPNWD
HY3Fr8Rav92XHbeCdLVd2HZv1HNWO1nChXCO5gn0hOLOIPWpAR+d5Bzc8YvcHSlPohZbL/3Kg3JT
hH6hj2+Qe6SP78MCYOqQZ6rj6t5sxQ4UxD4VPL2x+SfKw7Na7lIVdSP0stxvO8tBfLzgkKogR3Zd
nalGapWdc3cLV+SUJAI1jOz9gcgJdFSXxACWIJ+WmUgfOhhjjdcYM7PmC3Uorvpz46xHmoL5MesD
OMit3HOMf/w9sJA+rkUbLICXDqeE8D+n9r0VJHIdf74DPJwn4er3Vu2uYv8ZGhE3DcJdxPmf1ojD
DLM5QyR2C7DMu26z4e8LZcDH4BX9Jiy7qAQueS1zoUOkyc0IWRFCQ9AW/aDKU83eBtBY0iS4LdKk
2BCzQl+2U6f9b8ndarr1BYIHCPR1pYk1/oNKe+xlKu8PlJLMkd6V9blNyVYD7w+RW+0rRbqH+Y10
ZiArdoN3jY+eE5sQG6BJjXHTcGHCmVb1Vz++ZH3AEDoYgUcKOBBs40oMVQlqyXmenMBeO7wVa8xb
gIFlYpCaBg18jBP0oNsypO9fOUVvQiCeE2UUrMJR5YJ78fsL0zVv8JPs4XHM2+DxCh5SJdeK8+gM
LUW5Lnj6F8GhudDeBq8gLK8Aqmek/B6tz+Xqt1gHFD9aboPXQvZrYL8G+emdWCLkJWa8fQogPSAi
F0lpH7mZYY8wyr6gXY5aY86kHSO+zFP6ToNLDn4B/iOH45d+fu0EE/Cm0BY6ITyG/l7vHzQli0UM
HKzH2VzJanAgcT9cTGddrwo+u+Fn+tGS48TCWbCr9mdPoYVk5TJBfJxn8ZW5uW5adYJh2/YJHZe+
9Mwb9k5eZaUVXaY01TQXod879JAQUMXKEBmReU5sG4epYiaOC/EZyO4GxBdjYw/qm8pBgVolBsdG
g2FF/qvkvAlpO3N8k0DUYKcaQQteNLtkgxNirmTYrHNKvhrGbYcb/88ay/OOCixYsJIXHLBl4U+i
qrifqtIf1sgWv3lNLdccp90rQOQPTBqpLFN6aewf8rihbaVDTNfw3fvEJdvkV7xXja5b2drsUGuI
hL7f7PyWIKse+nhPXz0Wg3bP7k7wjf3pVx9d97FexiB4HkyFoRqK9W5lSq+3VpspxCopisFSLsso
e7WJmxD9Ijt2LbL2Ol9sNf+FOJX8oAKwenQ29YSfp7f2o1X3Q+SXg2BUl29SJeJTPQM+7bGRm0WB
YxHy9tKP39/V2niFdn+6HlE2q+CeaoE8kkVbdIAZZ9uICrVEqaKSAU9We9MHTcvPuKsq1i6OUjt8
FcSZYxbVk1XO4nOZ74M2O9YCX8Adr5jtxstBx/T8z1YjHipIZrpkfMEe4apQBUlzUfJkIV9+pOgv
nbEqnLIpFbJOcPYrcKjr88afGemseICldwmjEGTrpPs1cHnAyPOBJHva3yswhl+D1/6Zah8BcjU3
HaudLtrw+CM92I6jREA+z3KRLnd+VC4hQXqqFyTHpZDtIPV/mbGkS03y7P/I/xtwwwvImAIF9ymf
x06D/Vn0KRRzB2TIE4p1UsbIK0oGFgiJCK/hGleA/W2fIOBxXtipirHUSCPknbh6oLOfMCMwRoiq
vm5+DsPIP4Bew040sUssOWjcx1wZK7VYkGMW1EafkM7XN5KvEgKoZHQykhA6TSOFVg6AdETXZKev
pqKSakHzsCqldAl9L3+LtP3m/YfKST5uX5WKcfscTNHq75loxm1K2giDg/A0m4sEVtBt8UiclZqh
XeEv5LufRNwBco0lXLVKrTlWZQuYfkqFfsytEufiSfkmghzpCCD/qRfD7Rq5jQKzy4mvDQeo0P6P
ESXGUMfDZNWnUL7dBGic1Cmdsalhg6gPPjMGv0Tz3EezrkJwt6ur0o9hpX67SHPJS/hrbNKN/mC+
F8hDIKSVU+kqkPX+nnoCtB/EJEBIx/PnbyqmSekZr+DT1/EH6PR44dbjBpYr0RkkaxD0067fBn/k
Zr8/DhtVMT+saAsjJJvwWznfIPWDas04Q0aZoUHYT/4RU4tzVgLLkku6llX4EXHSs3tDpmXm5lot
J0E9zWTyG78CtgL2+TfAUXpv5bVdFsi5kRZHYK0xj7/Bo2GkdPM0YlTLidnyckU0YrXZRfuWKird
K6MzncUvQ7FMmghPbojhAkCdei99SPxYkewvYnZK4Kt3pnuDALM5zWPo7iRWMMDEVEAYWkuTeYm+
Hh0KzgwS3jNNj/xllcZDOMkhh/bQc38BD2xYJo3thdjl2+j0+oRGR7+Fm9zwJcQdW3pWneN38qah
flaszTpvsG/uR3apvLkGKt9sVs+A1xvaS68FHyLp3Uex8ss6uxVrjvSwo7ky7fnwHMtTDp47a8Zo
88AKS0jT8I89rBDRTQOOSvqAxgpvtBFyaHs4NY+Bh+Y4ut+g2NsfrGl0okiHyPAJQcIL5qBkEkeL
x0XkLEKxhRgVGY01wpftkKUtfNT7UoJYmn3bIFi0mT/c/zGe17GnK49sM2Ih2H09RS+uhBHzljRt
y2ZkMvjBK2/fPOUPYfj1ZZqFrCD3AicsQ+k+U5m+pQ4qLOINeB5b/QsRHqKLKQXyvpBM0TvDyzRC
CtSvxYXgzK/uTQJ14kPDoPMGZM+FlJLsguYdrR2PFUyMzlEYc+sBLHB8ckYN15uLq5Y4yPZO5dLj
FcopRahLkVptdz2kybkugViZgsVS4mzVl4iuark0koERvWZCenNyZYNO97tiZyHKp7J88H95Sr8i
Ge3HcgYaNyeOjCd0wSVzPuL9XUJXj1PmVuj4oXZ7d50vPuPU0CMmR7tktz1HIKZvf5Beu30+TNfo
W8HvOG8G7mfA1hKN8+c/eYIs/mQqw/MQ9vL5f6nyqg3QVkyerUwH9c5Uuscr/Uki77kq/AAHpzRy
GFSE5/upeajYOQkYykWfMjMx7OUMiOFfXvEBgeSJfE3cTF8nnjWhaEEQTHKAel7FrP7Ao/mhnWiw
ZmaT/yuv9YRAOC5We0yKOG1EAfuZ6yBLUzeHVDpnh/j3/9u7o7AIVQ+hFXw69Ar/1/LKlq/++KfS
tdVdqRjb5IDJf8slHwRSyLGvLGKTq81hQtzoy1M7jnTOQnXcETVr+HbBEhsona8mruILJ9ADWvg0
64sAwcDno1/1XPlrZN9FFSetPq219G0JAkOYMEw1CIiGK2JLOGiL/GhqWg92pQa7QtfW/TSK0TvR
RnpKxxRKHRjcmg2eTkLb5S9PNPnakuJo4BejKnSTd6nYLryV/QipUjiSMpGDQYRhtPBsyNqJm7Gg
4sN1XOPLXipuOCnQwInMwiepnk7rhmT/iUJ6nUXCYn/pUaAMGXxvIUR2awvXeKluPEOsw7vzaRZo
nF2vMs6nSy+H44MYkxd52kQTp3hWix0xZI7rbDQybf0oxroF0MhpSCxj8NoYvgY8MTgL94O9Oh64
bGv9i2ElOgbxqG/MzLQz+8N9Ld3EKXruW5USyQRxG/LxstRmZ5PbWzR5Og2z/kPYtcBGBGTCa8MN
8G4C9VL8VE46mOEDTdZomUblg7UcXFi5Zp9iu6q7pAW3ElUMFrYiwmO4Th7I7YEM/pgVcT3jCUtX
2VmeBj+UuDqrVY78bD+3YeeYy58HAIm/YkPT0cgTqivtMa+b+sEi5K0D5MqaFib2Idb/QUffzjQt
uvsw4C2VSYZ5rcC/vNHHaINl9m4Q4EMa4MniNnLV3khCaECEbQKds1tMW7/VvMbr1X7MchCBaDxt
cfXYSm1xcDyEatY1EaKAI9qV+ySeBAfBEcWWEmnX1WKEo7yq1zjX09eBPGSi61ocGWsFsKxAMfON
vQt2SFyF9qTQfyhPH7iF7NBEDtbfRK+zAeG1fSORoIWTTeIutmuVGJQP4zDta58Kn8DIfWuSDRHE
tQBA/6LKn0FQ2OgwS+flGoccf5bwFUf8Lm5ubJe5oLH+Kj2vW1HCBamci/4Vy7R4vqXDJwS1kQ9f
F+QZjz6Vzrrgzoi4naYtAyZ4OdmGS88ctrn0JGrNMWRBHvgZXC4hQ24VPhE9DyhFlSS34QqxeLFS
Oj4+P3gtgPEA3TvNn+H1DG9eFuJuYJSDXnlEWKykouM2I+0KR6XxxbJ8ZsB/bzkHKP/mXHeWlU1A
uGt4x1RTFO+YWxvysjGxLO9XGifuUufRsi5xqIkH4HyGd/WTaxFZq8MRtKw64SZeHPk0iOmdgck4
dlg5h55SGdnQteKzvlY3WuWP3nyzOVa2heAwUwfr0E2T6sgZ1v+Mu29Wzba2oK7F7dXkEPmOHgDI
JEw3F+f3id1ijHuNr6do+vhE2tGaA6EFfbrl4ZjNDivIQ7gGABd5P/ynp3ioHGFqBVMvtPMLuVfU
guXzUPGpjcv0AvBTF4c6dZ6qP9CXE7+wMQWX3gtS+NNCUHivLFLyWqW6KGbdrZOCDcwk4Kp8iaSa
0XbPaBpcMUFQAtdVBd92SimweSo8h4WYCe49I15vDvs9Se9w0ZLnWSuZlQl3fUTBppbI1zeQOSbj
rwFlhRw13aukWAPzmQRzSh400BKlKJRFhHIT3GDIhOVG0rJrfvOnrYrBK91SVEP94kJ+g7SIwkhX
56sx414YRWwkZLcoi1IJ74FoAnPIBvdNW7F0pyJhSFJkXNo2p43QuP7tiyaadCmQwjpH/A5AUch/
DDPa2GQ5J59x+8tXz3vxjdwCQb45uq1uKenqu+K/yrH+BdlwAGDh9++WGn+/5UqDXBncfTqz6t2S
TkEN1oBn1D1EVIkOTFCBqFPyrogtFO5jf5MW6ckAczDkvk9+HHI1v3mzZb7UxhkwGjfeW4QZ/S8v
NripIN/vNsPmj25+O3zyqzEX87ygiCCzOIOskSVymwWbmgBAo4sxwtGLK5I5XSmoOKa5hAoC/DSV
BMHhcLvlO3W0LH8WPRT1mkD2bJ/6RgbVAYzz37XxNpHHeZaatq1+FJPtwteFtepvWb0Pc2N9zKVG
G/SkY3m2Iig3/viX6S1xbgfkFz1VwqhRIFS7yX4Mdd6Y00HVeP9R189q18i1q/rCckUcQk076v/2
DsQSjcFa8/8dvOfSRhf1Hp1qPOE7AH25wkwRo8budHBjiaifH6rxJd9o+RXHOkxn1S9Bnc0WPGFk
viXm3h5lbs8MdfgLwWjUPkCaCBEmAPpkwN0p2DtuaE4VRcBzU1ytpWaeZiNoSLAgHL7Ug7OBjweV
EKLDHl0kb8586JVbleNBudtfC1BV1tRk7lRo6P1MOoMQgY8F9xs8rwmBYh44QxH7ldI7V+p2aoba
ebtYC65BbBIkUSIIHoI6LcWW4W0U1LA2TiD2TEWsWN0tTc7+agM25c9omfuxX8w+0+vlqBygWEdo
XsyFQ+jOsr+5ekM5V+8U9st6R8ILWUMIiLidwo1wazLYKyBm9S3WZoDZre9dRFpaGDqHQ2DwpHwD
uSiLs4ScA0WvuL2E2m3UMqqbArV6IeqHzQzySg+sNfinulVuNx7eTMpssNC8kfWbR2dihJ8dkqkx
7Ihw55bn8Ycu31YIsn2j3zvxeNeVUQAk5lS0Yyld114+ihUrWHpRXB/LlQUskobqVAmivBCcVNhO
hd0biA4fcjaH8BFPNKKT0q004UtFehm9uwZWINgDVlr0flpKOLY6m69QU63oUuWrF4fP4Rxhzcpm
YZn37/Nk3RF6Hxafoua5hXqvSfqAzn/Sw9PbdRqN6zvZQFC3b37Fj8EF2B5MAyHB/fcnAgvb5lrZ
iV2fNl7CNlhKmYy7YchV9WYKwcyu2M+Apl5PJ9m90PSAwCSzWSivAAUIWs9pSGue5ST2zrcM/vVF
vlHTdGyKFUlNDb5/Hp1Nhp9ixPY6BKrW/UsKb+knn0eOeXXcv5xh0yLug2YW8/iZPs1h/mraTpEh
RAuqtknP84YrGUN7+0WrFhdSZewm7UIYc03Zfm1CoVio+FVfpNjCKW1dGXk118YrdZdjpaQ4LyHs
wQ1N9eVrjHGTYBeKZykG3WK7XLa96DkWEjjmfzUiSbv7424PWInCZ8j/eIjsIFn/faj5uyHgJ3+I
ufAmpLYnU+pBwG4GM3aA4lF7oYG8mJ9JHA/P2Ri9yb0Whef/K5lm16C2W1qrZ3OTLmeehsqDBPXv
oQjFl8AYQ5Le/Qh5n4kuiGpBVL4NbSbqs2Zq/dGXsTHxJ2mFd/rzW8C7N/q3g3fctuQLG7LTAHoj
YsW1H1JCCI9qI4w9AeJm2Z6qI/8XLZbiy+sft1lLzAuU+CtIoe4sii60EL89olLBVK3i36O5+gHL
9VaNw7BIpNVbN/P3OrBcC693lcr3vTLNabqGQh78t+eB22j1L0owX85NfU+9rXKoPe/dxpT2GkH+
O/1dcRH8X5nCcMD5BKT7J/LdMFAyRYl66MHlz/IhWtjG6brQWADMi5JUDTkisXiFIctmi8iQO343
MZNyInHJMqXDVbc2U469UORPHq8mERCyb554V33fyTx2PpiHP9UI0lAY/ZVYdRcJeE9MsxOTd0v9
gMHrgwzVhwAGTonniYwlJlldtuKrPJpBsjOiR3Wmg0oAByjIknC+qYUj1dKq5XFV8vD0quge2C/v
26PIynUSJext2xXS2bEeY1HIcqtsn3ZDRwwE5U3C7410nlnHYI/LVMbyP2VK43b7H2VaW4M7H+00
SmTqbKvv4aQYTm/2H0c0/+AZb8i2epC4CI01+2y00DmXClv4+H0+irBuGz33HHioUD6q2fPtGTfz
Kpch8l5+f3wD7I/E0UQ8QsPYnGX9ybZqR0hXfP2ZPxyHTjFyeIGGw1lP5MXZg7Heq9QTEb/KIH3n
AQEjGelXjJekHM36zAnabu57LdyHC/Z4Ncv/868K7iwuRAO8V1i+TqmpYNWp1PRHVAEeO2DPV1Cn
umNXd+qwQXYpogiyBo/6foJVuTwoZ8GsECmZoUQv7YAXEiX1ARCQTasqel+cJtWCDMHX8jZuEI2V
VJYYVLb4b0/1eAWDsVJ3yOe/Y37oa5iqMCA4MOz/9bpBFpWiXfGOKkdm/jIxZvEQDNn7gf8pICaB
+Lg5HTsCiArjnsIRt7Nu+BVo9d5afEqoGUlJWdzQhuTl83/YmDsONL4tHLK5gulcZhoQEkUuK/RG
9TQOERa6+ch+69dZoS34v0DovVF+ex0fHL74+LOkJQ800NbU80h+GwWorLPqsdm0OOnJZI9riwl2
rNSqVAgBD50lOMyV+fBv8d45AbOJEEzjdWrqTW+qx4OY+DzLiF0HWGhfMAjzMh0Y+qJ9xhNiL+sm
zzB/nTDZv4ZtF/ekbyBOALuzCj/gFUXm2mBqTcPyalWs9sTqXUfKzT5PNLvcunD9p/xSe23IOQ9m
k6FKvFc9+mED+Q5+OUCKtVMuPba+B9vmxLagTfY+cZIc41ti3czUDwRgXIt2F7P0xdXgzVFFKW47
7qfxSi7keWLgh6kOHmyvgW6f0KkvvQUYi5NqnblCXGKqqR2uaFOlXslp2KXS8BO8NUQAliOuhsX2
XPmajq5JLjF2AnaQE3BqM1erdAWg62z2JgcXbxrauAUF9qUyUZENsvqZDv0oQTmFzS0HCwphSuSb
XcVWQ3eH8zPGQEYwWUPsVTBLTMp0F4odiKnBPs04SqGLK3v+uJfxWgXsXgewtnvg5nK+h0rjp/Bm
IOmDv9TwcoKJUuilwsWH2uqp/7TppaPybXHt+kQcqfOBsroY1QbSkiCUIVb7ujtKrjqnlI9s4YjU
rDI7gfzeU8vemUwwSlkMUcpFh7uHcbiJpRwlfBnwCt9LKeeGB7xpdR8tMxF3TdCj+5yjCnS+4zhp
2g7gXSOjI5O3TsJgU6mjTJPa7N6U1eOSZ4bCzGgPipekeYMcQ2642GwNUiyY55DTPFVeNTe+OIdb
lFcjLK2gHpN24UAQs1rt6BDPCPwGqZkEbpOE9bCHjzESHDbMq2WCwJX+8C7sA+OzeL3glMDaXd2Y
lfmrxGtIIF+qlZ0NuKoyZHRuYb9j78qmaEmdKomoJfu+Fh31ckKJSqGVi8jBGMGgHQlH5hVnZxjr
m15PDuZSJikRU2rUbv/7y2uXZlns69eXXX+hR0u771lTQOl6zfGZiqj6lVgEns9f6TBYxdgGaXHT
2zOjN4hUwB/phz26OFDLxd2UlKhfyHxizy/7qXjGmDmb+oBknS3kHAcIxelE1o3RxHPfIBmuxUe9
+6ZsRhNn88/vviKUkx1qtu+FlgP4WwuUqarJdVzRa1G0k9V2pdz/+2S1AzgBpEGZHo3LbZg1PaHG
rb3pmeawxJMuJzoFq0XBMtmoRYfQeEbbDLxrmmq+eMDLqtschTMzZih1/P1NkeZjCYC2CoK+/XKH
OqEtI1of3strppyYrgDGqR2x86FmfiTEjUWgqai+GuIR1XShcn8kXXC/cFMAwi37DnWJAsmj1WPR
k++CAV1bc+63go88O1TIapygYug96zYnDaM89j/T+MuFiiCnWK0Gm3rPYCf09y3MIzhEtP/F7vdy
WHsoJY8PJDSCzCz814LutDzG/yNd/H1muzsIDiVh3kWrIgaC3mamAwfvCkd6MGZTIikdXcuflOGs
GrKObVekcJjwuC7NvZxsyavvbl5AEGAm79N42X+Um/p1/domj7ZHcbixIArpOG2+MreU3nDPuLnR
ZT2jgCExOVPURZRESUEtQu9wrsSd5fNWX6UF95Lb4jht1C1B01P8bfkj+1mupKlbpa9QJgRfAJC/
C58r43RRZZthqjSTuStybhKKeuHjxZ7FbuoZT+3TiOs5S1PJ65TQcKZxdTpbENkBPZogvBrMa3v1
wJ5pR8VSrpn45Fv6LjelIf7C4MqZgc8C3djZ6XckjL9pgHM52InEkmYHWS6+eGW+qmhsncd7Oy4w
ufdUNfUZkxp6gms19tvSATv8SeLWJ1UtI/i+ltQhNbD5XQPyr4WpjeSvp0PVAjELbD2UKgyCCnMH
A5/04JtmbIOqYDvy8g+jIslhlXpgrcABGEYUPXoFSoUGakyGshf46ng+iFVrKD1+fmSITGBnUsmM
EVHsVFlKMJZ2zeDvgmgAFOlbpzn8XrYZfp3sHhqZjiuefn54KU94Tu7sZyvzOXV3d0oZq2UcFfKZ
rAW7cCDTiRfUR/rfxuEKjWtJaQSZrpiJgzD5Y20vY5wH2CK0Oy3kL7XPEU+5KaNDXZqaCiPOQhRO
FVWOVQIAgjIrkUUAgvUn5+LSOW0mmLHe5P1BH8yWC7oLIvrjVAjZJWvLl/ppLjEtJYIS1+Sf4G0h
tUpMwlCKmBMCbDpjcDKGRAq7N01ZdCWwzkHxiMS8hLmRqD7eZjsxxSBy9lABujvbnaMcVLZT2l1p
BB5kK02TAouBhgi4TM3RA/ugLkp8pSuv6acjpDHD4l9SdVcUNJwCEbvCUGZFkCEsFQ4IYr6YS+P9
yWFIDUglJluxEoVz6uYMETFZd34LCnEkjZzMbrTMQb/ubiuCWww1g1Bfih81otZtNWmzVG7+fWqc
QqfvCAI2sDVg8pxgU7fu9AKHj9o4vTZimZLXs69GdbmX3xUk8r+iK3PpAY1Zl6f3AoYMieOCqyzq
u5DfrpYZC/MTDoWSAA+aWtYbQ71LnDodk8q54R6kCidavC/TKIKBGYZn+wa6ZoUSYWUnOz/LAq2/
72UVJYltPqRyfZbA7iIvaQkyeD/3yg4RFoStFuQik4WBrquqrT6fYyC3G7cuHcHVyutP38RaLAq2
E3YBjqkvtjKeCpEgcQzNswTYPNKrNitqxO7v3CBLLnQVCLs3Zf3JB4U5N7qxXMT8hR0jMCQzLJVX
oiTgG5xLN1F9wEh3nP+KpuY9YN0PP9nNHghjkhPZPh8uJedcr3p12VjvyXXoQl79FYvZxOVhyeE1
HRiq3pSe3/HlQUM6Ro+U2lAUdCI85z3n1Jnd91LmjETEv9n2BabBTD4a/Fdi5cbUcQjPTomWIDgQ
+b8c3GXhT8o9GHyq8+iUmwmQbvP0FKn38DDcTts0w9lE6Om88FAcZl8lpKlL9RaADI1tmtPhcCZh
AH0s4gwQivbJD6BFS4R7qamUIjjjveC/pQLWW1DSA0SPSXprGQxDyzyAIn9OkslbiKWWB62X+8yi
IDXCCWhkabKSiITQOFqsWMbDeZ46mNcLaM6rYujpnZJ/oyf2TqCCNKn/imNzXhnAPvt71KgTDtsC
RPRIbEvf2s3OM2OXTYxwAWJf7igqzNsRipaQa2muJ+TLm1hZeaokqFotEFktyc3+hueDvCcWmCMm
lLvUEujT/r5kSy+R4hF1hM7qGOeBqRUv901OS9cED8wI+c4OejKmRyAMu1I5YDt7WqbeD3HTDQtR
d/MOhW/x4I+XQgQ32QGse2oe4UBAP7NelRrc7pnlInqowZucKTDAzrj922+EgfqGyvCrkghT+NBs
iOW8d65fvlIJOKROFO/Vk0FTH/yniSJ0LaoenOSypbUgahbykYOeMBd7mmrhWS520iyNNa/KyKzX
cKCMbrVXCvE6QwRqyhvQ1KcfAJKpG3bgguslavJ0O3G7IYI0LzpSQonFG4wNSnK55efDOFfRne/2
8i0TU7JJHeoqTQU8YZ41laacfqJ0towBEO29f6IEHm9lVpVdmv0fDmGpgCs5KHJfshhhOCVnwRT5
r5Fq2fDQ0QO88X60n1tV6RIEqsDtUYeGDUVS4FZNjHYhl59A+B4whaDFbtnGWJs2lje5xnLDApqY
Txcr4J3SMsKX25bPANCRxmhrh+07fZ7D/RQARjoEaKsEG4FJBayxnuQzRAJnh65VSdT9tf6ATZyO
1ryZD/QZJS2+G2FqRm5n55A/sMFKCZ386cVjWb6rbmzisICZQNhZLuIcAV0Lar7eUHAMkhYcCSGt
L4hNh6QWZopyySsQduv36CoB1hyyOZSZOlUhzSQod7lLZKzoa6yR6CnMMERhSB8x5iF1MMwD5fh6
dXekgAaUlHhbzqI6JHCv3D4vxK9e+P16N/AZxL8GTnByJreKs/ANsyC7zT8ceuCMC2JSLTAEFyFK
S3/U9354HGxa7hM0TTvlzoqmJZpg0FQ8UZFkkHugNISIZUIZX7NBbh8hCv7a5UPeECOPihwmUbhA
UyQaSltX7dYEGVCSWNLDDa6VOQooEEMI19afdPPGCSLtBPSPQA7b2Tafpbm7HYaTQpRz/JP378Jw
dd2J5wI2dYATB3a5FSftL7Ft29p8EhnXcLiCsE6I4OSPPTDrMYAv/g9fkIx3P2YwpwBkO592pOaK
ufHZkYzgM4SDARh5E7UCniemockZyjk0qFGT/hj8aYqwDBtYMKTkOcKwkJdDhtQZfiMJFxa1oMAP
MqJlp7tsTSjWS3z40gD7byH6+R25X2qPBjoUIQPbmkS8NWFlQinORvcmgvSfX+0fhsgAktICO+Fz
Ma1uC4657WaByYFjz11mryO6MUPLqLqj/7uFTlNCogYJstMI62oqziveunRcr1KE1v75Galj1qgG
utdAs2TJVp+JdegxwGi4c7Lo9yiUwWXtOxW3mUcZ+CF4asCuuusxvxGjkevmK3ENDNE9PioOAP69
pTUseBMCI8mA3Psjib4terad/GhoDXwKDQOGipW5dyQBkjTWfdKawHSsUyd3RuV21gEYxi+sxfQe
+HTq9kzuCFkx6GSDnqm21Hab4RmiZcI164vohvc4jYW3FQTG71oczVaj9+pQJyeVDMIzJP16dvHw
vE29RrN5KKhhFW+SjHmGkCqyU8CFVdVbGOKwIRgEC5PcZqSmSVyk1pTryb68VCyNN7Hi5VzvP40a
ZJU6wy3Vcnx0ZYy3Xd9Qn6E5ROItoVUr+yi7TOP8//dgSdoLuCQD3NPiKPEYjm5QMA6htHAa1uDM
ZMw9KGjYED/pjgMECSiu7lbRywKUTMVq6mWmAqFw8JY8VCPqijiwyWZB/J7ycF/HAC0NEr3bpWgu
kUeXzudhjvlon+rokwGMyOv7EKYPt5aPjTx5SF6RBdFIhsruehZd5iLtv5Wwf0EF8h1gbLDgT/N7
A+GnFksefPqF/+BPHbvSh4kR5WchIfJrqNMxEB44pY6CbP3gQrPyXoZNe/TDtc/U9mB1+s9eWMI5
N+o6D1l7OMJSF2v+qzEJrnOHc/nwWITBgKN+KkOxwsBOnMYNYMpOChopBCwD3U1LdJRp5urGYuOa
rSJ5AqABWTl73K8GPI5DFfoLOnnDD/Vuo/yv78ilbbmEIsUV70EAJFjEPiRNtRou97wQxtmvlsRL
gm7dwg47lBOTbR/XdX/h54PcRM19GY9z333fVd7MC4sLBfSvqOsnWcF17hnJ/LD/R1cyGM9ip1KA
LM7+n7iQtT9tZKAujmushiEovbm/3thoskJJP0Ae++X83sN8pwwuR1ZxeMW59+L3oZL9lWxONrtp
1UqZ4Fx9C6/Br4o6Pcz5XiemJkn+m8A2GslGfFdC8H0C+L2V9Ykr/bkw5rHFun2K7phMUwS2k8E7
igJ/vGTYqyoQ4NV94ZSpDLgpp6nuBzZHoUoJ8S3cXtX8QBIht4ygLT9yWU5regsVzE7S2qbFAEMe
wXfV+HM2XCBJVu89pK6FQnzDbaI6Kcm9ruDLNT88b1Rb2ake6GhQYfoc3YJ6ODZWz2/FpAgNEDOs
DDLzJQonwAdfwUUlh/B/NaqEawGKJ6b07c+uVZ6YGuQqCdzJMMWrh01l50xBe1mJVk8E0NxKwzlm
KggQ8y/EVW4sSAPtP0KQQn+84Jrs3qT2SxoAM6n54njVdbQrjBlJvzzBM3Gu4WPtehCFkjoJFo6q
sXayELr9dsHKHqYXOmcW0jj8JX1n7c8GsIrylLb4XG6aOlxKmdxbbql0ZiEU0EL7rY6x+MV4z5R9
kNSVnhWGR68DLDD4OcBEV090xVA+lK/yw05GxJMRP7O6NRv187a6/hu9h+Rw6+TEfirUkxtMFduZ
79lJEsg0RWqD726QMM6a2fTaH5UgvATYraJr4NEUf+OqMEatir446UW8ZPLyUcSRsbYsIJnsda2+
p3BlLfhKrx70MU+gSwR0p20o5heRUm4hpOp+vuNJTgEeI8b4F1mwB/gf2GS9uWoTEYZArQ3bUtgP
7AgaWvyCyvT1flnk3NlUUCpcuUJaia1HZ9VTDviad26ZJRnrcVbgaY+Z/IS0GeHo3R5ifPYFWZsD
nwicS3XRHFNsgmXf4kjXYxg3SfZ1rtZeeQKHRxgC5kOShs8OSENgxldCLUa/4LWAFGn+a1srA4fX
I1HQFbCsWLalgowCO3+RAZfmUddwuWjdbxxgYi4IU+6JpR7hgV4S95wptZh8sUEmDwWZzBJIzeGK
u+TqY4nk7t4DTkch9e38/nWS6OUFfvjAIzClZJ7ZIf2nWrchPu/JSgTpWErw+rIVDye6GWRWC++W
57+8csEd/qyEmJGLBa9iCQyX4fnKH3l8yXdyL15PrzHp/u/j4wRN0ITShCwEVxTatbDSiP89nXIz
Lx8NyA9Nmv/5ilMxBRGgpN8zfyVu/hX7lC+7aLUtBSZzN4p2YBLYHPsNcp8Cc5+v4ZBji7aS6ZKW
8G1jUa0hqeQzaiFnW+/yaakNHVw2Zvm350a/wpvYYue+SeoIVfUp6nD5SL3YcVV61GAUThyCY1UY
XGg9HGFWilgvj1BHAiCIZOpMiNgs12V/+k1h0CnAHPX6X6khGJacL2wK1pyIL42EvYb20d5rvP6z
gSLE/+12hBJutpZrg3DxjgDRBH2+Jv8Rtt6eusd94UXDU5oE8BZNoQDcj63y4R9OBYkhX1S1wFeT
W/CHeHSTECZxixjvdX0FVQ9gBP7e0ysQvhuDGR+vi+/54oK/T8xsj8tuwns9/gf3y6wPBfs/jTg6
+FG3ex7rzl8uRbWY2Fc8OroGwNHQvg2AHeuwuERhCPA1Q8LSBA5N0m0r6YoNivAqAkEx5ZKChdD1
6ozNeU1l0FglPvc28oPS7CBnOtuo3m/eklk97PS8EMFUG8OAeImil3IlG9jIalFmVlI05HAmgx6I
vGx4CTpmOKVUqWKofxvy1VXUDjnUCVVPivOFCVx4jvPQW+L2bhfvsZreLLhKh4A7sqsxWvQU++lC
gQTCfCHfMdTnlDFtEDDls0RWux4TFIdEo8lHY9p2ZZpqrcHRNvTBGW+6OL2xRNQhi5DATzcUiHMU
kPtSpLTu2OluoaO5vt4RMudr3vupSal3capBXJzV6m9CSJqNSGwZIBxFvwJw+MYp+bu1Vl2oLVjN
VnJ8q5sib9ipx0LsD0GBCWdD98w/p5GF2GAJR/ThzkHv2u3UIPf4pkukazuMAGlQAsHy9/WRExzN
5hJpb6wBgyRMUhHBgIpuHbIPMnrIH77dmkJGjlwx/rnxs41ObEAYRQXy1BqTED1GmL3T+A2pHSVJ
msIyb+0UpWReVwBq8IBL+QkQC/ydFmG8LEYMTLkZIX923Zup7IloF11tAnBg7tROG3Lypzv+GTpv
hjTHBAWurq3m676FoTxONRo154bbkn3zA5MhKIuwdQhfKanI42/tWjKJVagX2YcXflkFtmzfGBv0
IgScZVAKNaBoQ5v4wHtVtocJIfxA9yA2TAQ/F47Zhe+fors+afSSxFLdux1Ll1YH8jcKxzFpKxuP
IW+vQgs/d/lGF843FII7SQ8P6P33KOFA2ZLhCvADQSid6ddtN7AS6f7N7VgjYN5HFw33E/Jbw/+f
zo2JZzOV4vnkz0IpwcUjVuVBDGyIibW1c55yi9mRdYrNoyUpzCKBTI/PQaeDEnkJwFH42UCdCSXz
UZ5nfZXDhafWjN17s/mLsXFrAaC64UuST5l5/bnaQV/Hp0KTxxmruArsF95f3gEJE/dK/+TC2TdE
k3cPc+DoSlnJ7Y5vWQjLvN7xKVUPtiBCOBc92/h18fM8gsdmJIQqcbY8jIVV4hJV6rpEFGhcwfw/
y8nuZ1d1lmfs8qZInSY/iLLiMrT7zL6fnB+jy2bM6jwnSc58Lr9SDpkZ8zD/8RDVJHvD4Cej8vWL
P6fskLDUlW6Gd9xeukGpQDw21Keco+Dwty49E3DhMQzTfyXg7lL/uI9qdeyaJLQAWveKSJRlJHgy
hCVGeBavtn+HEOPV8XMhjUxofz/NB2ZNM9xHCdELspyMUrUIRgPEgQPrIGQrux1p/nQ1lK9WcArE
FTEbQhXrYF87tTaAbz5GPn9H6ul0aVZu+WNqnEXq6o7JcJWnPWGyh7gT33OeS7JTe+qK6DV564DC
AZ/ipheETuFAWRP1/GOS6cFkIWNCWfzIUUUcTqVAaz5xSXameh8auZyx+KWrOr6yNexYm6yVWt2I
n4P+6efc4h5+fBvPwyTqpnN6hd6nZ8ws7lHR+/m5s7fHqsQbeh0wtPpdV7ILA/yLe3m7UNJzuorU
tM30rElZkUWvj0LyTqPgho8eUFmYt7mTBWzlz3gkslosGkkbnxkDIpEL7fmDXzsnwUE4o7BerV0E
McAFgl/HymvbGKAhfeZ2qGlsbpwY+PHvj/v10zxYcDiB66V29vhqAJZ8oDLDNwBrSxcbz89bzKtp
cAy0sHygYMTeiju7n3pKlRYQfRClx1RZvsbmMwT3Evrd7khoNT24UbQ7o9UrVRNNn581undM8fGV
i4cB51MBnodEBWauRgrWDLGyaIKHMqclu6PyYfVf0FRYBh60M4TwwptYaARhCR5FNVUvKGe6iXAD
q312kq20nbQuoM8sGBavG3pHuAT2VPLJclKbTn3OgLcXMwEa/vM7zeL+81WrEuwxJkDKdzuvHUsw
Cj4QzBqT5cwSz5THb8UHH3JgVoPu0tNVsz6GreUY/6+es6kvxzNf8NfwX+6WfAgThLCErS0yP71h
CfQroWqog67ppfNT2Mz2ACwwKpyPZR2eRxPdpxiKbcSOr0S+42IEkehqWgLdDS7FrZu6ymFcxGFS
vOcXMAaoRLzMzmA73IPRmb8DGm3fa/9d52uK3aaoXxfQQT5QsIQbx/0pLIwJnIiY2q5+gDGtDwla
IIyVfmOXnAhZjz3PQqW6fGD0Qi0TfDbHeyNlEWBHdPZNlYR2RyyY3xo7PJqy6oXZAGHgl8azmGVc
fmAECeTql7dGoR2OmLf3Sq4gkCYT+5EIQypZ3vTktWvNKx3iBLJAwGrjexA8e616Ze/8OdkAYnHE
5p/V2gllgW2MrJvU67lyi0BxCb+layMi7kK68DgPYZaKVciIZRdw75My26BnxyG91+9miJiAmUQk
NBNsPv1woY42KnFEY7O/38rO/3EInC5SbrwXsOcHwGLM9/NkcHFdkEI7dMKUi2CAjxGltrAwY3UX
BFCHL8MiQykYYwVwHK9i/kqX1Ibf8kaysZDUMwMBrkIgqCvhY1Cgp8OHLc3eeLsjC4n2gUQmRy4R
8NTEaxcF1y7EgICRph2rkiChGPSeFiLiDG/FiRjNmfONFET+11cX6wv1mtKmBEKpCvDSGf0Oa5UP
2m1LUAWKpdkSF7wxgtCCS62t0RGJ75lK+Aqr4J8s55lhcmD9HH/MS2p8IcP9Uhw2X/Lpdx9eNSb2
RflpaSjCc92l0r67i+4ai66TBs5shPcMVtcCw6ITCYOS3CW8Io37lMcqWZxXrFlfrkBCbHqPoTH0
MxE4FfBeNNmxMBsjWvxr7oIjqKPRfYcLq6Kq+58JDDmv6RSVJj9QH0ZUxfzuxVrgTsRUQWFHAyFA
gb/V1Iou1Dd7/y+3Tm/EfDeYqy0wJla48OxSEZYaOeK8GisjzRAvXVYUHOlqqTqkpa03sRh0Ti7v
FceJNiJ+XJrKibrMaejoGAclirVInx+XwTAtVGxw4A92Y1jEu4pNVqzo3B6xfDpTvFVMymdmILR+
y6qlbiTkR+txffcbPJ/CQgosyOwRWx1DOZETfmkU7H2XK38xEdtvLyYbP4xb4D0XJ8cUN7TWQ6mY
JRDHFwLMA1grptaZByYTV0TBJYFcEIBaScUbMvGg3FLS8c3Ve0/xPRwHYbyDsnGoBKaOqbFB8DPS
VLbHVZjJZ2YpnY78x9nRGjTUVzkfJ31N8gNG84xWExIBX1aXXA9CcE7Ax3dcGm9eJUS4RRQdt2Na
+e492Z6XRcRD3aK3D84LW5AQFjZOfwGwh1GWM5vF14IYautne4yiGG7eXu8PXUEwfnfI4UNf9Vj3
EpyjAHlWgQL9fqTGPDizvoHr8mdFHgMFjMdUArRqwkhdQNBzIAfxmEKh9gSsQcE7lgt3ZoEmEVor
sa9AF4om6vJVK/0gRHPBwPxsb23Yf27q98AP9gziZzT2cNd9FiBGwqh3XTSKzeUBB3u7+bvi1CK9
cPNQEELoSeFSu8DrOKydAzl5arP/gf3xdga+afjPy0Vcb5kFIcqeutT7ov2ivmR7wKJa5LUEf1QA
0SrMA1SEIDomGZqrw3bMLb1O9tm/nr9mbN4BKYQLrkWGvm5Ppu3pryBz1Jvf2MJkKIWsYp8+FwV7
2ErC28iCS1JTY75YaxCw1d65ySE6UxmVc8Txtxt+3cW+uRyXAf5//uTyc4oVHOOpWxjC79BLFAnd
xafgt0dLek/EM4kBIhzSD/hRW4wu6ka8PPbB8RgBP3hr/yVBxatx2IF3bDjTfeXXC7hwasWF1KnK
ng2Ns6V04SoXyXgfHBDu2tCDkAHwNZGkx+dUVDHlX8VWWHLN3XSNH5EXs1KCbr1X7dP07qz5a6ux
fx5aUQ+5Hb2D+4uzdLWBueBW/Ho2xsYmmiKl/69JdwTE+WnkxodpjgwMixOzVoOH9AqSpjAk1EGY
lnP2iVb3jFHYRp69e/zS4sWb5oJJWcWAX38wD+rSe95iazluxF/kzQZuXJ0/V8fUO/Jf3Q88focQ
ZArIs8vzJuEjxcu+kYeB3GQxrIM9uyiutlDnwcGYW1JV/3VJ35O974pqAs0xhLI2eTT9FH8txbTr
ydXn0MXmizcv0Aa/+UT0UIv0GVXnauUudWUQWsSTrv5xsZTs2qFIIrSE9KrntzgzAQ0hlFlFXU1U
JPYFu9If+4wjHIPcwiQsDhW3wNWKVxNbPkT3KxB5wx5ReBNorB4/Fyu99oS1LTGqrALqzjnJ6rlJ
tvrMC6AVJX+BKT4i7P/fKydlhUMSmfSrd5hG/Lt+3MbHfGYOnTq0lUnpHiF0NCGYVWuSMWMtESrG
clh4iXl+uFEOH1QaErSB+5Vz6kOQlwOYGn5qIfaG0EZDjCF1MU5iaZ1Ap4XSSfPyMBNlXpT+n3DO
frBs6HSENqSCmQ7ZBXUBW9u5FshTmS4KpwFLxCDqkzyZnticjetDAARNgjPeH5NaH3cWsk10NhjZ
8cuA6nAV3BMuq+i5zU0AILOYHYyDFAVVLk9da2Bie1IF0QLoKR4JgjlLMmevWdAid9pPDNo783XR
8jn8HVSIEsb57LYdJH2FjhwWnun3edT6vvC9lpCK2fkARw+jspuphjmBPmLKawTcJ5zJS6x+CvSB
wjpRdhRsEjNiVDzpI+d/MLTF+fbRuWm429F/10C9C1V08l2C5bqL2+OraS+P1kkb/WJW5EUBH8z9
qBgG3ofdxYSYuHDYUmvP10TcGv+rOitCksetgUCZENvHy0ApMxC1sgD0LrPy6FS9zR45NvHTCJaP
CdN+NtrwcACbXlts0aHqVSRnjPU6q3m+3/Y5+C1uS4PtTONX2Rut9Vs+zLlOt6bSaB2wzXnnW8bn
lOTLZQHtwotewi33ZvAX4Vl9woYHuofbKYEI4qogIjpJeXWQohuSzk3ZGhlnIIFCFrqojF3h5sKR
vYDwmT663/vQFabCl8RCJjsWE4HsP6etL7v08djtG0TIbSfXnF5axRhJ5zutzG/e2/uDBnPzmTCo
81yvF3U9SQLbkHj1aLSDXZhrfjBvgl4CcutpWx9Kj8ihh2NgbsAiYs++zytN8b4K4Za/F4cGhYvX
VmkfcSq4Mi+4JcdnQeYI4JNzQA0GrJeyKardkXfJdPKMQa7XDQ45DBb+QXXQ75lw02hW1j5niO3Q
H4djnvBPEc7LF24OpnAvocVKDV7M1Ef0Lkofvr8fxVMGU63z+Zq2a88EDbG22dDO7HBNXH4/QXyQ
aBYvuh9hPTr2HgoOtOK/ltqs46OqOpgFvMd51z3S7w2yLkpCESAK+4w+73iNeZRJ60fzNq4jI5qH
LScKg+vtGLgiwvs0Sw5/wSzTiy2WQnw7K6LjqkyKRI8gywgas4qU5uBcR/KDCak6Yo0hulC95MuZ
eEQ1Wn9uvx4D9SjyXA2/yt34vDA0hzA2WqACcI/uOnqC2B8OGFPa2HxFgC9IjTvNUmC/l5bx/S6r
yk2aXf1oSHEF59MQqpSwfbNErEHuYmDi5hnprUYOuayrp4wNQydB4igNyCCs7ASL0cgZljTCso1l
lDuQ37Gtl3JyiYyBaq4eTif/SfQiKEyfXSJzkU+u1HMdD+q7T2OirU9shXc++f8jjmJDOMtP7kUb
7F8bcOLM662j2YnqoDKSgOnEWuz0vNiT0E/pmbcZQ7mbx2IT9RKwPnVxP6kwYT1fkZA3pFPVjEam
k6hZgwmAWsNP052cW5ZU9bXlCm8pSNiSws9gaZIoaakcp6Kdz1pU8d0zn7JGIf7xgKYlsIJkzDma
f+zecrC6vqVuAACThcT6YbXJHqT43oq7g83QvgVu0FvffAKP7dzGuBehqG3NS7pK4ekOwfwld7W8
uFLBT6sgCHCl3qfaid7/DVLGGtO/UBzxqnFLOhXekpNFxH34HRUnw/QUy54YmW8UoPBTn650owCg
hFR1S+RcheuNvuaQ9MiZF1DJ6Ny7psFQhSGyfpE7cIsMlukA4iTov2VOalJrB8mKchtMqUkip2ku
OcC9kuAxnhE7+7glx6Cqb9MyHZDSVZLzPNJfozRn+/dSd5Ic34WRDzTb3EqXJ/kIWfEHICim6AN1
H3NphyKuNPCGl1aQ3Y+or7hmFt/oOBrd+en3KPkclO46HC/UqS+XuhDM6zUv1YFbncS76X9xJUhL
Ppivv084O853YwRzoIWLbdU9qIWjCsHjGN5rTYUYJxVVdUrPPf+RI7H8DsC1/aTWlutjLUjv2O9e
92nSg1hFDDb3DzyY0nZ6zZ/C+/Y76GEWY5WIM5h09X/fudrF3pnaZE48huKUkAr8MXJGAL3Rf6XT
pIYQz9lfh8BqRl72GnGfTb1A4wiAoGHXk6jsRpZ0PkbqTB9THge9QXOhgXGl4816AEgQeJvQBbwG
dDssu1x19cmJ5s5DwiI3q7dFteZdvOeEKq1ziQskWsGuin2orX4UQsJIVaxlNzgm3YrLvWqsIa85
pp9UagzIoL6N4HPJDLQ/TaGrf3gIPSJRP730dSKsNsFme4GX8jdl4ajUwdeIfy2Gr+BnvgiwIavw
3ABN3YDFEWww1psImHB1tZX0+T8M56lbObPyGH84IPLQmbAq8/rj4ZAClt9ZuIVjmpu9coc23+Zp
Ch/evdlvbOjn5A4JzIOcHvnDoMvNF/MCckYrVL5e8dB3AUgpJzlxP46JO5Oz1WpcNvGmyostTQpc
B4MZniZSsrZSIklFd8J/X5qEAygI/387C4mpt9+Svko03Z1i2TvNC6P5vsevUcn922muEjp5UrzZ
msu3xQi3uKcPgsIivYKj0A48jD9yBM6aFcFgGyMdXOQluGxlbjFK5akm3dSUK5FWU3A7uSDP4VWY
OX4qWtXMskIwpq6aixCqlVYNECf36qk+A1jUglrRWR+qFERLpjgM0owYtijybM19ZkuDMtjQwG9E
KUQSPxWFOtUxjJZ1d+sE0udc4QTYif5ny914GprNQvdf8yrrI8xtUsAl4C0700kDjDi3992cQcL+
eq9jb2DFsfxHYMkGN7ffy8zpfCdKVUGu8zAlbvIBaNx52jN1pOJ1ae6hSvqi7EaYvO5wmxLdY4pM
Ze6UHhInUvsDA5mBTNHUAYmN5b1VFTVFeQADwUchlPlyyRMMbvVnXIy9ks5QzntWfNRyb2LNOTNP
tr5U3IJwkEe9AgJTBu87Q2jpEmq+eGJxeKMZZW0G2yakl0KWQhgaSZfWldkRP7ZCag1rvZBuhTnO
+KoxNBEnUb31ZEXWxem+lrfrmQ9gxULiA1i/HG4ntLYmPpYtJAdfge1wMg1TJoAaF0JJus25neDe
HHbKiE687YTblpKPqtmLmU5VyFWJRDHTQ79l82TzBO89l1tsqkxYCE9EoyvU2Xz3yEk9tPf82POT
M9eygXrFET9PRNRhiaAj8GkqH+cQ773oN1wI/UtmcSvkukTzZlxkdBjdF40k0UYshb7+Wl1G4/H0
vPyy9lYLmM6t24QZkGPqF2hErHgpnfuxKJVcx4xnsvXph/99OdU5MeoYMIlnSfrduzvy4BCeal0s
/iwy26HDREwTxqzVukWZSEa3iOAWsCrtXJgtzMulM6LljY0PXn5YaPneSeAlwHl3wR3iB59zEwNx
eqy2MwXjYZcW9gGqvsmu2vIz6vC1lRL44lEqjhjNFVSdatVjI/IlUTkISjQ002Zbb/p66rHabVzs
mNr1s3oa+EWoe+X1dp5WGZmB0NXYzm+cSZoltJb4rV4Nk7drJh1RxLk69QhLuXeuE6byfl/smN5w
xszaIGkr/QA9pIoGyI3CquEj7TliHT+ZzmUH7VS234Hq4J4jkmGdYjw1YskifiUE5LbiPsaCpAAE
5YANsWigWb1XBB+cmv51uHesm8lrmomEbTk3aEl0LWwmM7klbVY//JZON/geuiWEFnW/a0tE3Ac5
Mt2YopdrHJEohhFbHBw3Kabi2iE8zRRSzq7ovnnf4BOe6W9OP5/6Rsj85vSk3Y/ug/GEYMsrJ9TR
zLr6UzNO7JG0791iNGTbmS4lWTGX7m4Py3hzSbp2gk7aMWid+6sa15Qw1Fr6gTgEfiJNZ2wgQ0Qj
WBkNxAZy5DfTHen+mw/xYNMoM7NVp9bnOoskium2fuXJcXF+D2H9XLB1ulH0PYCQGFsHYs6CeDYB
/0P8miFLtYdl7lxsZoRIRPMLP6QKE+5KdF2TAXMvFOSlYxFzAr6tW00NL/HWDZS+n87jpTL/cKsR
9w+as5c9dvKvhoOSdBvnaIQf08EvAcFkxXbBB0zC9fs2ZSmaZLnS7D6eSCIy52kftsNHcQf3fH5E
Dh+NanlO/PyBm6Zf+6NOe3IK/iojCJYvWz5ZJApS/guACcRXk8PaFR7V9wxvDhNDB6Qzi4/UCqGA
4LykBkqh7jmDmCdtBwacfijqZN2trqdUzcij41MzhJwVc3qVkke0Q2uCg5KpW3ilJq2Y/+KOf6KU
MwjHoznZ2BPAnfyhoUd+sUJbyW3BxkkYMwlgzDNqxymdj/ZcbLOed24xKMEa3KBQf0OrAuE5/shi
QD5cJf8yIKUH7j0yqP4AaMgcgx73BExHmDc+O+TKzXa8QI+ueKO1tj/y2a/v5rCiddXRX9MvWX8Y
H7R6SxELL0Y/joPS0exDv3a55NTf13n4oOzY+1mxNWKqA+v86A3w4S8bs9tbyruCZVzjfS15d0qY
kucIbEXNaNM6PHpY/WxRJvCDT7g7LpriAQZq5I6IOy22RNwm8bKql30ax3S1gSAZL8OBZczRCRC6
TosSNteO27y88OrAK/yGL8XlTgd3Eqf/bAdBUXVtAPOCu8HLdNAcphdNm/FDDrfozvC6tAsFzN6T
m0Up1a/hQkZEAOvtVC2s2+ZSny8bdD/7fcYMg09sFh9x72xu+69q6VeOrYRGsLHqN9tTgkJRsJAf
znpARa44yZRQPiYPwvNs0cQgMEoNI/ehZpuyEcjjxmpsbL+qunUZT5VUKC6BsM05+u7+IdEUqddx
THKLyE8W+HFaXOCrBBNq4KHuKnd4yqto0XwJ5nqbYEbdLTW9rHNC77vXBvf7qoPAHYwjkfKDZen1
8OHUj/StgP7/kdspFZh9SWNbSyC8KUB8dJvhD6xAQh+RjBB/l5f1iuVK1Too6T79n+HompcnZd5X
mvXda6xQY5JmjN3PnyhIb38Z1H61CwX6jN2l6EFc1Wu+CDvQ1ojFLxgtn1HgTdJP04y2oVjKz2vS
2CfwfzZKuu4Ys6yTfB8gqP5FLZ/c2kcgYSvoXVzbp27ySYgJPIxpHNcjjqM+bQG5K1L1ziQqpb2k
/mg7wLFRs2ozX/6SRVxIRs1ybB75ZeaCF4I8jbqgi8jjCcquuRhTVvyrt5PsOHLSAqnIYV7oGx+R
D8u+KipxsdXVdT8PVGBj+bN4lZ58RtZh/jl2FVB7pghEA65uERGjElCvIU4caZxaVqyql2D8w3dK
QvsOMXj7eobf0zQ8HvJgpNS7ElHePXwkcZ79XY9Cbej0yert71TFuZ5cxOVxWMm951JGHoxCLGO0
mn058UgKhAOOrTLmP+TOpYCtuwYIoQdhcUwM2cqqc4NB+10w1cWJ/lxeAXshz1JCP7/jP4kFtmOL
ZZYuPB3RKrABN64PtJMrHn9a85ZwXoq1ol9X1IfCYDzehma43PvDfZjx+MX37p5gStMUKkOW6HdM
YG64VOYeetJCG1U6Hn+TQRthMGbLtOiar7mIuO/uaLFcsvyfRBF8MJXFcDpRNuPXQVVZ/HAZJsOX
YUzKBUY67+igQbMmBX06QSHd3BCmuFTUv7TJvhNEZHAphTygz/LhkwmKNudYO7mlzWa+5rhzHhs6
BC5b2RqS2gTD11V5gxX35elH3664FuXfEjqdotfGUCjoocQp1nUS8s/TEPrdjORzIbXM5hzJ7RsV
uC3B9WjbbCNOI+HMi924x+21VSwHe2XK+Q/HpEgJRUcHGVSdy3GTC2u85drxji3qtk9k/mDhvnEP
oy6s6eCPL+j4u7INXHskvwXuwMBx0E0I/FGJ+JqOwMscwlqFG2dKVrtBluDgsltYFQQiF1xYNwKZ
5wQH4lh5Tr9h58HIoOKPFPa8WdKLoUAx10bplTLnpAJZy0NMv8QShD6iE7nxXDcTht8Ny+3K+Lzf
ZJLmpsJBSfhFzcfc20caeEuHHayNPJast/i0zsbrw+QwSsN72exDmJtelHKxpNosTLWQ0L/RkH4D
uIa2VxdgcYHA+OnJWhY6vAsSrvIkjZMwwpHIkc+gIiDyO2xUXZxmmkJ6WxFCER6+Ad8wzL+umQuX
OTlmU7rbP1jL1m1uqLKDPgvaN9pcfw4FqjFtZjUuusIPx9ILwp43KXNXM0ONn6ecWPuCDtgZgxBA
0m/YLZq0myM5FEJIEtHxgM+efoa0KPyooDdzuSFqpdWHAfCeEoTI36bUsaxc5JXLICV0jeFoDh2o
37YtMYkcQS3ZeykNpFWJK50mUxSd3eBsV81HTn2FMj/hsvLtqwo9Ru0c+VdVuTyzcIpOiEBQd3TF
Q+GnaeFVLJWorB8U3P7qERxzT+6BIA8ilIzltBtCAOc4v1MPAEnITUJHJnbmCUul8el3Uj++0pdV
Sf5dcOpouLXkyVSN0cRZr41QKynFNRB3+GOqGzpEspJ0nEai4jltBbq01vBP2NlEd89KX6WIIRoL
hbr9mVpMJK0fKHTUeq7wKpO6D+zfqQ5yKsyASVcRb/KkfQgnlhVosArJQWrnHlyI1Mi3yk1bjvHa
arcs/2zTJTcI5IBxVQXJgBKUvUhVVi7W3Wg48tuBIZ/JnE3rBzHmUW8my2J+iSU4cGOBIyrLBtR+
SlHXjoQ+EJjb9YWACMpbY0iruMCgiD3wpIZQ8sqhWfLlCpCyzDkQJM5/ZgdhnxWRp5Ylnb+Dqm7N
55IbnMPbqILoMfvOQ0l556hawesaL8bLbcEZcGxyGLR+mFlaieoA+fzqR/rKiK5J6TtVU74Qk94M
pWLF35jgPOHr0S1oQsCvpHRGDl4VRia0xRt7oSL+YrtOz0gv2AU4yKHSXrwJ2AyZVKuIuqEeuLls
z3c0Ejw4GathcpWR9fE1IXIKCPzbUhovOcE/XNDKC/C4hKiV3BKZkvwVTUrL1ZKMcM11ILeN8DYj
kKXf1kSkzEZsPebJVpZIP0xfymCNONAwwJAibVllX4eiIYzvjUbzVJnWyYRjB5QpGfTNGfl24j+5
HQTH7thc390AlXDgL1zybHD/32knFOx7vmaMhm69RRkNCUn7iABks2qOIqm0G0uvX/1qKGf6E8Wf
8ns/epkavdu6emiLR3mKJ8FJVrzYhoJjyXwV/yu7VIq/d71bhgb39qgxlosexz80dQ0owExB0zht
FPd/zrCDNQ8EORmc4ElI+N2b3y6dktrXvkBh3aL2gMLh4sFnuP1YRA9dkLta0tzCzmREpAJzMCB+
94VEDXFD376KNaevEVxY+J3CqzgzAnJyRTgBLpT1NF93J//Qv2DIfxiFRcIwnEEmTADfmneFVrKM
nD15XZOEVvXGk2oVO7CGzAG/yrxTadvrrHNcaI2yxTbH3BqgYUfpNHcUimGhi/xZ3ucdspGUGIMZ
f7QMnw+Y1NX8o2JnB6PwOeuLq3LTHY74CWZh1jxyxB6yV2md9W9FgEN1YHnLwYIx3itffb3C2F16
tTwQ3VslScDG2QfYfW7zkHjMLjbRKqjnw4sr38KZHwT0JQcAmm+CwGUqcfJ2QX0ypccgBuP/XhGW
Y0qawlQcGQKLPqwBPzNIi0cVRzgJhlzePP4M/U+A6uu3SBw5jRqxhIG9oBreJMZIN3Bw1m3DKDbf
7ju4pAOOYAkiGT4izjigsrV8QyRk2+B/Ik2Xe5QsdYjwXljK7Ye9qhSwncnLDc8lw/U0YFwjZ8au
BUppgU8WtUQXESNdZR9fKyhJkT3+HBcLrE7HWr1kQfMKNFgT5P6/Qpc/M8A4QyIaAz3KIpcgTw+k
t0zBDgkFEa45yj8h0iA3dmyq+jMcx+18M5eT7Dm+j/gEC5b9UEEd7qTqzkGqP5rUSQpdrvT0fL1g
vcf+xsX5R083un0PF68r8LpP+xC9Sjwx8TDMKP8aPLaS21oy9HkknNjxqND1FsUnyqb4vb61scPx
AjpD8hkRckQ4xgTI71tWWCS4aNz9sEK5S88FviMvBaIArhOWl1ZUnAJkNo5SC6jPKr1vOlxLD7n2
AAHrmg+fWIbrjCjeYciGBNaHiGX3qmsV6uv0XB7JzV/5YDkApnpaZYL3hpxZGxYZfMVgdJqwaWb4
FyVml59CuaH8KaE4NUIJcg9I5/rv9xbvH0QGeZYSCVixQZMA5hDLXo+SMXVPCqa6p8ztCobq7rei
C38+glsoHYEJjGhINO8sfK/hZzriFv1HE8HiKGqBWIQMZCsC8FbEDXTHJjEn6zf/wMOa/P2MP/ew
dzW8mWfFovHQbOj0luGqufcv/bNbsqVi2fmZ2lI+zylcoZCzw0g+Mqxq3dkX1y8d7rYBnm0YEWb/
rGZOWPfs+0JTyiOc+1ZKfNmBc0KcM3V38KkqwTACuQibt6Zpds7fBSbPCmV/wAerOqBwYuwbxTSs
eLDgcvNil3Zlt3IQ5WnagZd6YitF6lFm2N1ZPjo1Z1UfTrqZAg16JB3/yk06sCHS+MYGpR556i1j
7N7hRktOjdGyyFghhVtBAvgSq/rOhsu7LK9XnA97GBfTRB0+4+cj4TF83D8YrDd+2r6owY3Mo4mF
QYFw6zmUtOpfcalHQOtwnUlUXbvo0P5YGZHBsRSpcEUl6wAf++Z7jNrx7VhGJFQz5KSkKHkVl7aB
c+Dt6nndVs2nrmiPU/4+Eg/EBF1wCsZHCOvmVwEjJBFwghL+ULDj2TyX05Hdo1Ypaf02HK9H7cQq
NkTr/E5QTNI5BmbzS0WeIi/9fgFmfoF///ND2TP7FqWucNupXUvhL1+0gfnjcTHdAzOqkcJpOzqr
N7RfdlyGN6r/mxr6eZBThJu9S0jBOQdZhl1fMCGCgTmym5lVS5jZxNeysZfoJI3xHlebbBfFzk40
Y2PonROmEQ2XlGcaEwLUDUhysXxrtqGWeTWZ5bm0+sZmnN84fcOLwarzrekIE5CmAscQWFDO6mHC
nh1KYx/ptkbK8/WNW8WCB6+bLvAbouCmfnEaK8hlefWc1Ld1f46QDTkQ0EH593hCn/tXbhiShy+v
xnVcI7hGY2w/lNgoMTkiUYon9SI7jieH+hI5jcMY/HRyK1XMAMaZ/lTCbx8HH810IZtJsB14XCEw
2GqJ04mWf+3U21lkQN4ebQJ/93AP8cM8SVZKvBX2SWAF3rqpN8KOOo2YnZiGmBbOnd6TQ/KG8uAJ
M2zYUb2/DaaGLvsc81wArFzSCMT78gGkuHJAa7JXGl+nN666icIOH9Hbh/YcfzgpQh95FMISKM/7
RP9xkwnW/LAHmQmfeHKrcDbJnu+B4iIUxjOCI7mo9BFnhyxtaMsSU12IsD9WIfdoxqKUZnYYymtf
ob/rRcy631gKNuYbot/JrQDlqNHQctBx1/JDgQygZlkEuv7XjUde1x+eahZxJDNUKOcpxSpQAUTA
ZxBlQNMw0S8hLt3AxygODqXtvBsK2wZmuGUijkeNzu6NYwQU2Vy6bh91mQpK1UfmzLCs8CLhSpaG
jPlQ0WvGGeYB+66J940cpkQyXnZX9aM75uSipd32qO3eLcU469M84EJkhKiNk5DHQ0wHKQw34og1
QIMQmz/dIOPzjzq2wkMnBlPCw2zfeh/qAJApctKe0hbHRDA6eTuG5RiGqazGgzls1o6m18fn1hTI
CKpRlFzy55H2bwQ4ftmW5MbwwV4dhgcfPfEUmXtzJdg+gr9egLasZ7V6lPXSfmhjtJUUMBKuOygR
SMw9hTrRKHxqNeqy1+BAiooh3uEB3y7GwwQz5kWCStW8CHwK7VqPoldwK6qGclcX4/Xx7zS4rKR0
47m3g9ARBn26F7jQ9CcKNQPnG2Y/brnHmE3BLmDOgVvpnoN//mdiOFhlvk7mDoNRx7vRv/rj7ks2
jZNg0vg+x0lyi40+UTMcqKuSVx9HPq3rU2RpHN63KcN6GPP9yX+IMh04+vGeqpSR5txcitVvyan1
k6t8XuWGEdvTKSqY904GSvLeIuFyvXkGQdSs/Zc1dVp7Yi47stVFRAM24iA6RDVTtj/hbIdloayG
eZoJ3fltc3YB/ZF78L1UYfTtwx5axo5q/lY97xjCYTNDBc2Y3VKAi4XwFXkEGXMfsGuzz6i1hHnx
MNk33Jw+uzu/mnb5Gcb0GM8CM7YEv3lDPmRZ1vge9Lz/Cu7LY2jk9g4cM300M7hFCrZAhF2wjqjV
yT4wFhTHLDlp6o3LwXtcyfRy3IfrNZn7g5rkMxvbJgJGWrwp6ZPhrkhDxXUbvGg7TezmyLgsiZcw
UJM3qXOZ3HGouFA4C5z9Ct2C0IjtRfzROTEv3dUCnuBY5k2BLUgyGq9LYaefQeGZVsaIWoxL52UO
xS9UUF+ClAp79YDlDn9pha4pAfBAYtuXT/AWTUlZEJ5aTb00Auk0pR49HiStar8Gf7ZIUN/uMFDP
xsjUCAU7dHKrzJInOHlFedT4fhWs4OnDUPAs0hzP6VJKHwckWr4VWDTJzrZQw2QJTSLbPCkMBCIH
LG3v6drpdbGWuKhL/NLrzXzy7Hch0BTer3BJzbySVv93Rj+PL6GV+XJYiSHgZ6+9rqe0srdyU9JI
vMdianLbyl5PEJw6fkAhjYYhbaudgEfqSem64o52pIVHs8Ikss6l8j85N4zaql3buL0lW9p2Yc3/
Fk3ZJ5YnWVMHlDw7R1PTNY8laXAwKGUHgLZwUO7pTC9Z07FVPyci147Z+Rr2L3MkUv7DQc9vvg2x
RyfHf56D4cAR+IpfAhOzJTsuz1muidmCG8FliWKAhUEXzV5vk+/JZGZJqAltAjn8TGc384gjwdZk
aNr/QBMVhOCO8wwqZosPWBl9kwsOKHelkneMXV4OA98QjgiDzoxFEvVQ4PAS2m5s+hJtF4DVSlTQ
EEiaC1m+lwihHco+8cjUxEqe7vCcAe525RFVaHP8bT6uRNw9KuZUMNl+349CIc8yC++NcLueVKwY
prLkM7NcvEcMuZIFZuQXsTw3qA157tXFjk/cXVZU/plnquh93rn5KrxPCGPHh6ItecUWQGtS16Zj
0tqWzEQS+ZN2v2T5auyngt1Kroy7Lek09x5HPdp+POtvN79J74NNcZ/UQTjgl68dx9Ik9kyeow8A
hAvcj1mXhdwNWOLD7uN/hy3PQOxDLT0OoeXaCwl3W50CUkwSYYtoPylZHwn4w4wOTUCnd+y5lWGB
iO0T8LKyNbkHkM1EfCJnROaZc5ZV7SjaeiBGPwi/Gs11gscJ2CsRCmBkxfaUbBGIfhSUHv1EHK8E
xQ9R91ZQ5hLGf+4ZjpgKrQ6a+byndYxxl561U+Em6/z5+6OScJSdlhZUt9aX4/XY8fYljcfMudSs
7zV0r5pXcnyv3U03MEaJQJRC/3RcgeHLJRuq0g209qe5XN5Xei/PFMJaLFYn4lgbkxXWGR/Qx3ej
J4tRBe0ULMzZjYRdUiJ+g2BSLIhby6kwTxdRFA/osyVh5j+KWgxvwZW6rMjPVpfz6R/R5S533WRS
UpSUlFvw/YEk2iwzn4D5lTzGssTelOLn2bn/iNe44Txpps/yLt7lCr0PLMqQT9ZDOB9rwjZep1l+
dTGGvIf2JEVHVJ5ekRwGFhFsrcDWp6eXkJlUpB/61vh/vFMCdXZhpkdxJ0m3dqcOAX/QFLM22jJ5
gb8E/9TzseYiWG+8c6YeeqeNq9greBi2TDGkb1Cgj0UFEbKOc8VbvNXLbdxkhRw/dW/ngn4g+r7Q
nTWPnpXBcnyK+nucL7IFBWc7GkWJld7jx6hzrCUD+oY+BmS98IanKxSW+GT3x/2V8hMf/lCZ5vNw
sg37VE1ixqBtWZ/FY0tdlZrP6HGdFGMXn3ctcLkAuwDSx9NTGW0D/yZvSpvaIW9Z0yvcKQNholng
ccdeQLZoSSwwLzVGbiJe2+9jcTsojOd8aD69NHo8zf/7HddHD2Rpn3+lKxfPI1+ZMHDRxfWj/lCC
zng4EnM9NLPJh+viyIuQx5DCYaeu/9OVfqg7y2jdbHCthg0QfDtfhNNFxcBlEYPMA5ratNykr9dS
JwgKnLZlUADMDVC7g2u6uZ3jwy0mT7FjcMnK9A4xoMwr1ohfHvmLn9QC+NsntRPznG9UPyB/Z3mw
S9deWpQmjtGDpfK2tNupSLH89xN49L13m2sX04jju3mfWuKs+ZKXOyHo+5RAwqfmXRL1RQaXe1iJ
VQTcFEZK8xb2JS90AcHAzgyxno4r9QU0NiK4tFtbF9vcHZt05ktvyv4RTpPgs/2eVjFpSQY/k3d+
BmrjCqCmIvuUyy/sgu0sni8WfsGyAt63ydIDYTa7VRNaby65K07/guwwPLXbOiTqxZ3+s0K673kO
J5xsIoPCrxLNz0tma4gKMZDNvQcd07k6xUtHkn3jlwwjgq201xyMhYbtAY1+UFBWKOWymaW9H6Eg
RdMr6yE/3/owWwPq/bzlBYRqTJX+O4gr5FNxN8xmm0RG3hxB3cYwI+1ajwbRMbDwhaEdyvLIWM2r
rLeB21sCG1MYjVRqpEXVIDbwAMAenjPhSk6TRCdxSQvHlAjKf5JQn2mdPFCm9E7OOT8naqQzgM94
rF/DlhaZTChx0LJvb3tFZKJNDjrZYVk9MzCF5BxLzLhzF7+QoA0d7jBv391CV786VlMC6UVxxQ37
L4c0ZRXAQUj4AVhyyNJ5nj7PJWFv5OPF0TBV7OsmHy77Toep91tRj4XBIJqWineObt8Fx0Tc1tqC
Hicqui6uDYEhBHKLDO2IQ+Z0/FcLN1NtOJ1NLeOcvOOCMgGX8MswxdUNF7rK9ko20YiY+zMlNuS/
wQvWiD+RucvHIJ5g4hw29pp5rMJxYlx0Q8yo78k19+vrUIf+lJV/yKKRJp94w54m6KZn2nOXiVwW
4p9Wy7XGwSupGjcmb3mVwxoeFvkLcAUVKxvdmWFf5bniLx15vOAytvmrkIDzsw8NlQQiO7XZ2Bc1
vKNT+RdDS/fyQV6CruitptHcwXGqloBR0Vkpr2CFa2aauWnRjtY+SE69iRp/y/xk1mOiql3+u98j
WBLE8q3C7Wgy4PZdu97GT796hMAOgjrp3NoeTAj9xXX4VFXLOz3eKISbpTEUhEKLlL+v1CogV+T8
aNwUx5WP5nBqoHmYdIT3yvVgk7Gn5Ik3Iq9+c0cHgeQcW5rx5R9oeXpbaH6f/1jv1zxEO3jTe2oL
sHnECx97m2O2waoGXLMY+nqpLQT/s8avBsIIARySttDtBgNFiZAtL5cxFT7ZoycK7p+iV/hgXrN6
hHPaUZds+NS6x22E+0jXGj07eYAeayEV3BP1wDNmJJ28Ow67xYmWZ9VeRMTCzk5TPEfJGfxeDQkk
BgwI/OupnpvsXF0wxUk3FA1CDCRqSyiaGDxt1tQT2lyDtKmxp6DMYRLtfH5WxKjTwzbNh7nhLl8n
P2ErxZxazeMOQsaptl9MNQGZ3X1Iw4oplB13WfgqzJNUr44PH+jz8xp3oTEEA1C59o5iNx8JR+Ju
PdFDYK8E5kxSLXws2WMMqUGx49r0JDLXe/JovhHhabpP9stMqCOcpQn44l8F8NBj1cs1UUB998ec
3ovZW1FAfGFLWFsqaJbkxHazaY2sm/H9av+DdhhlSegqpp/GLBqfBGe+/qMMFPHp7s2OqQUt/vKA
dc//ztpjpF7tAIN/nxOKcvqKZ8IjQaKKEY0hZGJ1od1fqIXta/zqiVHtZ/UEoG6fpoxj4kD72EHz
gkKGbwKqGDo0ExEY3SYUVrgN/nIbEAdaucC2Gp0rOs1I/JHv/QkgYxeEnTu954Ce0Y89DR8O2b5E
p6XzQJ/6Tu0P4Q+uXHV7yBfP+VyC8wTzEMay3KsldixEEUD0TU2vai0uqsFpGWxbfwpdIPrVMwuu
QuS/pkinNstjyu8J/McZ3P2HyuSe931UaT3sTj9S2DJUPMVpzB+sI7SORXmfJsCk+I8tFbgATFwP
a3aJpkCoxmUgg1gTtjjGSs5nt9E4Ag+fsC+cvBASOwF/5WbBA9Ji/FiXcfRGmhVjmL6WsGFVtJ4v
XTeg8ZgNu17Z90AxglF4jF+2ZDXwliDImiqLd2g6xp/gSRsWq0dIKRhYIogNxpY9cMuiW0+fRyYy
dn7QouX3ZmON/U8x12/hAdLRor90bjtraYejgETaKNmN3Axy+YdsrMBVZsnD/NQ3O5Z6xN1mchMa
dRb2eHcJTlNOKND9hxla8TKdmdk77v3pfYOpIZckIIUyzNnSZyNX5LpSG7lnDHv0ggm5zaYvg8Pg
t213SrUKZZG5QjN5MqqxXVarphdhwkRplM0Sr1ZXs4k7RKpr+wEwGbJ02mAQbb7mcJ0ceT9Wem49
A8bGJERCoDnZsBzTAn6tcTcJZQcV7j3PbGP6UaxoD8xc3oDsiAi6ED6sbiQAjoECUjKbi7TU3o/U
ahycr0SsjHvInWV2U5ljGBrgmC/fAFhunsJmDapYxidngAj8Ie7gy03sj74xcrcTWkqQ05GmacZa
FfkOfkDeSjw4kNY87j3HrOzLNC1x8j4AfKtTGsbV/lPq9QOheD3SrQhT/5zZgO7QD83Wc6Q5PpVf
VeYW/K4fuIP0roa9KsuL+A4PHviFAw1SHsyEj2ASWZD6XiL2XyNAKrUjkJiu2UAEP1d0j/XexvQj
yulv4syGWvi8fKB0RVCUGR56RA40J8nu8g6B+Oso0E4i1AmGAh57uA9acuoPko+Rl0ro9idEuP3l
vJ7WhAWr71Wnvpva3wq4Pu9WLMYtwiO6JcS5ztSjCVLsVAEDQSZKxRIMzkkx9ZN2R11Ko+Uf/0Mv
9IL3u1Wnfn7uNAEno5WAtlmRCIoUADhMLw5NFShMEO7cfiTvXymNQ4tynM4zXu8a1NpzZ9F4W9f8
0vXdGpADWCS8XF2c5G4sqoE0AuS+t7999F1ASY22mAAkQFdTbzECg3k5XTat7MGWmxdhxHrtjyws
FCaKdmlG9XRI9mi/fNQv/jL7AwuafRWgqOWhTry+REKLny76CpI46xljcqvcsu1B1VCl7SvUWBJC
0FSYpA9KVLSvP6+gNq2mO/oFq18lxgPokj87W4jCdfUharh6yeRYrIAqFGMzo8RNP039T8LwV7u4
0h3qga1lxwlXnRl8N97v9uWDcwK0iKKiYb2oQvLYDcQuXfQuEsiyby3uAunGFeYAP3fT0jUiHvmQ
TC26E/FPQv/AgppdRX/CSGb0a+1gjNGGsOjFsoJWzban1PvcZ+duoewTrhi1KoN8xafFEK0jE2z8
4LMpXIdxaS3Qp9t33Rc61i9MKcO0b/sC+aRe3iyJZCPHqcqgVts8aHHiEYqHxt7Z4kD7ubeibxyB
zz6TpFVf/d/fDQ3agKQ0TixMjJmNXP5urt0gozns9Gn9orppoezUeSP/OT607pqNiG9Y7T65LU/G
yOiwderVe8QkprGaaGMSS4lqvKY4Lu/CxswesCo1ii1plE7Tx1voZGTTpmi4O363vkLf2bvESEzC
e25hWP4w4R/ZosqBpSMMmyjzLnxOG2WZRja4vy7bdIf5hjoab7ts8yn++D6I8xa4S0eiXZYPgIPq
PNeHkrdi+bAWGHJz7AKDzqNCi4e/Jp/hEWWap59Q7K+SF4pVbIq+QGxiWp9SOpBh0tjxXMWv6jaf
lmHYW/tB+2JHo8tmGG+FMR4fob7aAuUI5KXPu8ljWiJk03EA0/y7XYh7LwO1+XvNcMdQXcQD3djV
a8Ogjnjr6zFnqUJE45aQNABHWzjhj+cfy2R5lZxKy7fRTEt9g6albwEuHei0smfaV+SGzqzE2J1h
PYxk3gT9P4Y4MC2EYsqCCysleaF7mHmuxG9Fhflrcg7RM/Kj6381/6bQySEHHdfzkHE6xceeBnAe
fFXAhUk12iFpyhTu/y7GD6FyTImEpQ0UNYb1WopMxlzXD7RG2nWpsN2t/Lxs/Wf4VHbzqRAWfJHt
+3lnTAA3TzKCk6R3ngd5rhwhnNZa490+mfXo2vS11Dd8npfT6QbwMik8h2HVIHv0eyp/z2fjgfeq
cvHE/ti3sD9mQhZFPDta0X1SLLA+80zMmSkpTJAdVD2VW7mbcUPMbsDfIVaooJUNvVweWmGVztbF
wF0ktJq41mAbPGiwHSkH/z8WE4NtMzDTHiu5jZFY/Xu38E0B9u53gqHyyR7nVdOkz4XJs1P324Ju
W9hGSLh0wcv0BGLBTCdaDAjcfIcoSDz5WtBs5cKTjE9OGa1jt6CYegIy4hQBfoK4FDcxHCPVVLxe
3nqopF6Y6Rp7iLIVptt7Rb8Y50M10OgFUZY7aPhFQLf0zUrmeQQBSIu+Kpb7MspvwWEopdBWV0M2
CTda35Vkj44mm2CGH3kvOwr0JqLpLpYHWrL/aXVh9r1dSkoZxhKXjlo8ArDnnjL9cYEZWO2ZgfWK
vCzaypGNcGOltuaEyHML6N2ZkxomCVhR4AFsOnHd3Ry16RTK8X2/T22ka6oeRliawJyDl2jOoRjb
EXHViCGBzwwxq2wUSEaC9Adokg/WYV53oYM6gzNNWECABLTfbM5318z/DpAQ/IED1omgfug8j7TU
yxQ+N/4bFtXGNPp7S87VukMX1lsVcn5AYlsEl6oGbBiDWX3aVDwCYmJMve67oemi8rOzCWqiY1I/
eCUq8gPxCKViLNMF10NWtVS0LlbYiGwWyzxAonIOJ5czumKD1yV5x/eV25sNvVj0GDyF1bTh4aA9
zI8nYJCBk9y4SB050XO77bRlErVLpGrUxQOyGlTO9pyggkcGyFdJy9tznKRpmMX9YQ24HZ//SFS2
PgPKAXrmxjSILS5zd+d42oNJM3sF9hjXPseAxf0dz81Py14X4NaF/szVsc4N+cfwr3CZcCPmVupU
49hp34SZfruZJ/9Nmx8EcgGvybgZpmbMZvY1y8FDYWEPxifRyl7QjPVjaz+ZwKWm79A+44MLyG+w
E10w5xzwZ6mONIZHtn+CRWPLyoGVad5GIrWELyEZYJRZin8bbrFuudZCkTfQ5PMDkwBj/Hhxm/NU
R4ALbUtYllK444FdqPeDCd28ypRUI+U/ga2ggK9aerUkTzd7mtwEmlEdS7PLHJ4cFyUnf/0Wiyhc
XrHFSeQw3Um7TALk3M9x3XE2Rm5owA3CxKVUv8yOgtu5dJM6a/nEabiwun8BSahF+elExBlJd+Km
zJ+4aSi9SB4769myHKYbtutDNKq8Nj+pwX00e+QBf//g4yPwGr7fdrghlWFOyKTOu+SG5Az45LqW
MjwN3IWqg4yrxboeoJiBI9TS7CbVE6D8QIEKv49yCPaMer6ybMRwv2CZNW7AbsWS/zSzXUNzx9sl
R8lRP81H7aEX3eddAnxJHavRvtABLC2yszPSAxWVpAR5bJvxmOYaCNvZKtcnxC6J6SpYgOvS1mt7
h7UVI+HclCEam8ljctS0yPoSXZ+wnOP7EUqen84HaE82aXfJawfLKXUnb1Dvk9olyuyjoNNhPewe
k5XXn+Gq21JeI0TXHNZ0vWoeqiWeijjjtRuj8rZAEx0/8W8qXV4513/o440UjIrMq/0C43NUljkG
Ohe/we3rmJxIddbqhOABXrPTuY2pUgGBD5djVW0hqT07IwS4iNwTzo0fP4bV02FG4IRQIsgyCrvQ
mbVpGo/e2DvY1myU8rcXkfANcamUBZ0HNFOCeaqYytwtqS8nPP4pr4BXiVQT0vKMIwF4wvkRhOIQ
EX3Bq322PjVaQl/GsMlIFQlOcfyk6mRIwdaKf1RnRaPyC6an7qrzDVaTeg/QT+iaqT1sD8hHb9cH
7r5IfwMliqrv/To4qPIeEwn1Kx8FUtphawZQZ3EMFRDf8fM8ivVcSoYrCO8EX5ToTRD5dbDDliaq
8J4KxhAY42FQ51xPYVPzA8g7eoUX/GA410VApHtoIuLoAeGSwymtCfn5uJumlWFfxDtBwxoyh1Si
h0qFj8poQj87rufYzYtlaBat/Oy4hljvnAIlji7jj358zVzWipfwzwm3LAy03Yh6yDoLF0CNFZ3b
z8mzLN2s5SzVQFV5iGqI2oP1S3mXNaYyRDnB3vJnBh22RASFUpeUa0CPZpOTt0R3U/Yo90DHo5H9
qs7HKFhZoJpqZ772tRXrRkYeAmgZ4ZEK1ZI4QrgUszKbrK/HgN+NqnlFaEtdjVzA9idmSWeOmgr8
CdIxpU4m+lrHO9UV6BB1PrWt7XK4bp7cMwTIrQmHzSshk5tr9NwvfQp8IThiusXOjZnsoIyg13vo
yhd83citdoh0hek8fSp2jPBHTJMlYA5yATf7g0y0tNT9WOTg96hH5RXMgp7JCY5PgwHeEGTddwDf
zfmuvpQv1mphScWeC/ZYyfR6jb9B3My1RQ72zw19CnvTEzYxYrX6Bo9Kiqb8bCTnFA0KUQbrOYHx
lmPQ0re4BGrYZOE7AASPI2WWloB5lb2YcsOHhZOIF53ljIaPJoUJUHgcuH7FZg/8Hn263RzNGVsW
MQvblNuRGWDF3zAfwCD4mrXUsSJLmnCbzuVX2SP5Y4s2fM7y4P3Z6vIWLP2KWhBJxExskYEGELBP
dQf5RHlvyGSj/qLEDmEqroNXCzWg1qviRZcreJgSGlJvYZAaaRKtTDbu+nPBaaiJdhyHUJCMkTcF
RneGYHvXDQDaf3J11l5Fv4A0pKoLnOft7zfS8BEwArTWBEO/haH0DXK7JFr1Y3Rb2idOZCQFVIkO
2vV6sWt+7UWTVOPqMBw55tYTuhgv7HDFtwcrrPU9J/7XlNC9keThcoP9TKz77WnOs3ianv7A5p1u
Aitv8ueUvySwyvOo0v65DlSxzf8TUY5PCSGtZnCDIDgPpozW+6vJj59kJ7qPxoQDCbIKUfxMWg8X
2Byx1t65Tku27a/f0yb1rsbF07RMW4IlerMPqL5Meoclg+/ss4RuHAtnS7LzLDi3cWmGLSZXB5qW
SSMIlySYY/hNF+4QqcjTSDksAhUCjOGNgkDoOoOITPwEZOr9ez1MCBPvDlQs7XB1vu5MlHOW3doL
BPrhK6h8AeuTOS4J9aGb4PUhr6CzLMF+LLXrdJVM9XPM0GJDMriucpFo1OzcXnTMBOp3tH7c9+hM
/uPEJJ1aRLhWzw2fRiZ1zoCcMlQPVqymLRP8EI57yvJ9BvtXHS0r2pMf/mYo3zP2YezcisFvcMiU
l98GR+5cZr8i7hutLX+SCosGlADboYznFXn/bvBTbAJQW2ep+DGdglGLRZkR3FIVWQK40uMITtGx
05wjRB4LOTHFpaNedJTrOQXEpJxWuCpIs9mSSqwqLX4ZTMFDWTLqZNx4KvKtNfXHSlivrj3x22+k
0D4LPWZDRGY/QN3Sp78z9ijrYKaHJP2wqaNsrW+UDUHBnuuVwCLeH1epPOlelnDlUWJPAhUK3m/h
SGEG08JHpVszowcG/C2NJqys1YipztoT8DEs78f0ETt+4+rWCSie6IT3jKcXEJDwrOnlXRj9Bn4j
epxjmnrxakZXG7qounmqnuluUGD4NESab8Y3PrSc8iZxXBp3IN10uhqVS+8fiVq2kQydVK8wEJ7j
UngcHZaJr+VM0we9Uy2TxWBKNJcfE6Gu3u0gLG++2BePmAbvMdti5dZPtCAnUw57MteM0KFwNOba
O8KigzN9AsoyWgFlE7HkEXoqrGbwS4+t3LwojpLUPe1LQqUy820/ei0up7e7hOP9cT8P8fnN9lTA
PiS4XFiPrWodMsi2yhr0VZXaH09adVZ7GhloweQP6cSyZWzqTmfWzmBsYD8mDicexImjW6KIzjjz
lFAtkYlk3DvM0bsmDpJMIXDpwAED5zzPtF1rreHqXSAi1DnrksAPDB4d6nBfdI/HIB9yb++EwnfZ
1z6BbB2Dlb9UNw0KwEu5FtgGfB7+bnPEpE8DivTlnUyAWHfdqBL7JInGmcr+yvdh5D+wp+18F2xq
n6qggPEaaH9VLf2ZLkspmBHmt9LIF0f4EC0bdc2aVJHZgXu4AGOhJQc8p+BGNzOyDNEHdh5/1FWB
h0BSKzl47TcuypQYhC1T2Um0JljQFvpfSHKjDPYOMs5oC4+cZNCOC1nABHGJJOJ71kjXM/NHSV1x
KDRD2AeCsRjIBBsrNi/YWy2cOQk8eWKSRqYNbLuycEbpgWS5lNOtOTVJIzLwlORgU/SOUKoIj1AM
G5Xe4kVOrOEnTm5RQV9MO8UJcta0Fh3dYVb8WJw/8YnBDHba1OwszHX3xmTiLJCUQNLuJ1QECzAW
nOEonR0eZH1BaaHC0Un0YndRk7JM4MMbM/UKWGekcgrbxTA/r3IfhpqREiQ8nm/vPQbUGjsXTxR2
fhDDewgdMftx2d5FmMrWvQZ3VV+4EJZYLCACvhCfTMUbDjHU9Pk/b1exIsh5doTU+ozLrsNusXHM
jybaPYFfSROg4WfZxO4wrWaGBoYwGDBrqijSmK7xgE5Khxo67VmqMsfXf6um2N1qf6Up7xtsQohU
JCUVAE5PdnhAi4OIp0jEI1X5kxMun0hFd2zv1PYX0EjJDiSdiYe2OURDYH+l5A36AreHqpu4XTog
u4fmGzLzDWSb7ROh8ruBlawhaCAwEzU8oUyufWpffyQhIOOqHgixBn/XObRzHs5QpixYZJUXQgRJ
BsN9b4/+YRljCl+UrcHIoHH+1kvRSgvyaNChun1G72bXzyEKHVowKHN4o+1Fwl7NhfmeM+HB5qG/
8PT6ViLjzOavVGHyLRHUhaSVYCD2bGR1SzubvrPd/x4QHuFTe1ZdbWsVU2hZtBY02flcK+5zw7YF
qHiTllo5qvIeZh8frQKaGs8OD0GizEyW0hCcdzXGbLQJ8WGXFjKu6r9m/jUTbcRJgSyaYE24hseW
yEiQK7KRs/097cLI/ZHZ2knJwlKHpRv102Odmq0kKsqu8h82ZgnvXVNa9iBV6XBCpsnvA+IyrivY
QomZP7tkQxW5L7aysYfRr+9sSqP0F9Ebs56nBYK4NkI/Y8wfr59MjNkLaOyzvdL01YiLDMLCBGY2
T4wIMjrB1MeP3wGt3VOipolsR4bA2FRvQ8mm0ETfGU+1FaItroN96bVlLtld+NzwWrTk82HNsYWJ
HnN3PEp28DGQXhKlkHgLHCxwm4v7734UI3GV+uf2r95YtZlaNryAYnMEvXQcfEGPb1YUB7Jnfa1r
8iQvhG9RbOHbGJTX3f9s5WMHuvPse+NYSH2DJtrKdkuBe01dUjiMV+DH6X6wR2teTK5rhrnngghH
2k6hzmQNLFqJXfM/n40GL07egrqQPCkvbaUH3BeLOnxlDgaGuW95xs3g4UyQmFP5YQZOVVpRJw+5
EQo4NwabhsQBINmHaNnA/AZlgQpQOYnABZfhdqnihGxg1CSh0GCs8eMjs8OTaqkE5K2bpe9kSf+h
Kl35FL6eYCXDNbkb1oksxwZ5UOo8Nom2dthJ4fd2KNpXVrJFOJFUPIXulOI/TTKbfm37nruvYUjB
ZChDzBxaXvDx/nRqnzp8eb4AhwjopS3Nk5lZPH34tyO2suKLCO7sCUNDUQcUWeSJxEO3uJqTmyiA
81530XcjKuMj71QTbQIIV0PTa00MKxkH7TTSfFJQiTBcA6nsUdVp/K9k7NK4UiBmM/YgcuKWA2RZ
V+jpmnGdJZQ8bLgJWR5TinTs2Q045Nx/RCCToKsGn/dYzNDYf5OneCILGvn469i/k5M2Te0dDkGE
3mhBdJDHMWjQ9mRz0hgJrWJwNUecaVqYV/4ITI+MK2i+Jj+iXr9HEzzJPBMyuE/YslTX09mDtrFW
U23DrTN/bgbNNCm7Bdb49hhvLgOgzDIURuWXyZVmX7VbONU7aOyHeHJBFP7JD1RFm7afFX0nU7Dw
FgEfb/t0Vnew83HfoeDrTb4e0fV0F7xdNxqJEpwIL87bBW9MBWKDh7GaJhQwoHR95ieuMpLcxepP
rHDqTZoyjTwhTz1GFoRhksJjhbI3NkEtkF0IfJrwUF4j+wAPzzLh39no+Atc9DgPYjYqG380KcgQ
d2AL/tYQOnn0iWlL4xJOXHYJNFMTdPVG49v3ORI4vo50ZltspYhmX7xKcySsbX+bv+6A2krY/58r
u26P6jDE/9Whyb03LrQ9472BRpk9Cs8mOidMTWk/J256VsBt3QL+tHIQoxoF7mXKaQdMd7l4/ieA
LzQPUW8v65u0LrYWP/8TeDJoaeUaxAZ+96S6pJ4B9btr8ylLDjuPpgoQwPDvwRukgPFwcNe3hb3n
15/A+EnVgbBp2ph+cJuSw981U3HTZ27qBUlcRVx0B2QDoqjEyYZAlK3epFGsq1LR91/CnI1CzhDM
6Ck4tucWdyZcX/vQV4/+EavFy88kp6c3dDn4YKBB73TV/IBBhKGWV1NJzcXzt4QW7gL+TgDWGwMh
xzw7lgxG+XrvQr2lN/vazUDKksxhr9ocI2ElpVOGoR9egdon6+E5316POrUSzoIVcI/a4ZjgEIC9
C8VshKWslK/QQT2pPMfSXdkWueQKGQ8+hW9tr2C8Fpm5mkWcaPxawd/12cWeojlo5VCHlXYF2oMc
f6ifkw+pQiMkcQ/Sf8FbqfNX5mGVsdGQf+IfSNlfcQzk1OQHMA+R2O9G5C9CGmcZljiXpueya+zv
oDJCX7qGfLAVGxFN5k4KYoWKIW+Qg8V96rG5iHmta/F0xvm1k7YZJhRtQAAJAaz5ZDSn9remhEP9
cd7j4JD9XtX0RFVlN5O1Vg8IzUdCSwCM8HZSx0sAnnm/afoSGiKIITH30kYRI6i90KaTUOgMb1GA
1DxdrVGZVCPZUXsMELPORMo1B98ocUBaX/BuNaeS+Hs4iFIT++9pUzjFtm5HfBn49j6JLY8Q/6Hh
U0GAceu65DVlQ2Tad7jPK1gLUCFdDvLLz14UBfJUMnOfy990RohLLppoIeX82Ic6th2nek+vtcw5
KddHE5dTtitRih8rbDqGlIahSHB+q0mloJR0bzL7cE59+wvz+7Y0grPcOBFqb880+tsEnMtfVsyb
YmYa+YXo+mCWatViWlB+yH4EsNb/ALIHyQgPKw+2exXKlOR+AA6/6EWd293yaWGKmPZOgzZ5HwI4
T/xybvh93Tg8hZ1ulp0vRy++/FRJ1NDvphSI+477tj6iOLQCqm6Adctav4n4sgIl/9536KzFadFv
r/Y8W9K7/Wjr199QqX0Mge5gpPYdHXV3cupkR6pD2yN+WJ/bl7KqyfGiyUPRI7a8/rKtjyPxb+OQ
wb+EbYBjDrNriEAU2fpb5dNpa0YpTv65vh5ZJyMiGSeq+i0i+pMz8XG2pF4F3d15v2kHn67IBDRg
OuB/txs20blJosddKYYojyFvE3/xIwKnQKCLgBDdbakLBqB7HYHVXzrONAn5eXvVx3czPH9fCBJn
yvehcXtzniS7kEejy26xkZ1PhGIThX31G/OcbzeOZXut3slRE39kpqkqW83jid4d1GfTfGX2Xuej
arYPmvoRfIBFHFKuNIlqOdZdKvwUYHN6jm9BH1l6J+nRHeRC8bBTrpfcnVktTwNPdSEnc2dJSzlT
YKSRD5DZ7RPfgfL8/lMbgr4651i/Zkjn25YU62vGR+6Kg6YumfFW6YQq4X39NFfq2vczXlu0MWT8
5DINWLKLA7hOSp2veM4EN7X62KYr7fJU2/ev/iGXBmFjnUSQvASA/QORxfBgkugA3ExdkUYmYC+Z
ivcoYzEuGTFwIbynIjgQ1F9fgJvQxNazyXjkS0tOfGO5/HJOUC7Lx0K4/7Y3u30a+jN2Ox9ZhEyk
MgU68GKUqcLWq/Ltj7C35eANdvczb8Se/SxK274I/Yq6xzNMjgC1DXtB94rlZXBneiPdFRrkH99g
y9PAfeU70RhyvIS3ZF4LAI17VhW+V1CkX47dwmJLJmL+qWpTt/duhTMy6CQoPD2TRnt+82bnbuuj
CozFGV2IQ81X9n0GX9jS2SSpx1XCzyiOua3GN9uKihXl85xvRRnxijAMOredyrj4UlFM7WQtiWsm
8n0RsBW+/3dNvcfNu4qrjQuvXu5Ni/nHTlwv4SspYS5y+66KJo2VMlWYm5opWTfGD0wJrwSZdtZ8
qsuJtMwjrhYbzXmxJ59t9NR43C73J9tp68kXnKCzBZOuJ0Yi5KaYwMDkLO1daT19OiJ7PkJKqaPA
c87u3QvDEVWZ8fcPXSqITWkWznnODAD+REv34DE8+PPLWc/ePDmYSuEJLLW8fiJL2p/9JrEerci5
Rw844XzV+M6ELwXO6c5fBUIJMRLslknZjonKvimg6cPBvH5JnOMUvjDQhT9kM/uzDOtaf2KyXEpb
2Aw1qhJwl8q/TLhIg8l9SG6kRIEZCsNHcFHHG57aley3E0+oPl/Tn+oJB3PLoJLTTXtgKJJ53zqY
9oM6NqyNx4mYYVOAeqwLrpWQ0jo6vYVbXVh6kAics12zMCu3+vjYd5wZ5fUopBKrp3gAxTzJvUcQ
0/j22Xppskkl7QkKg8dGS8NjhU62WiL70RD1/ox5qQhUPcTfAeDNUM0NxLUFj0YsJdK6Tm4HPZZq
j6QJaAaIHGYnRpGosa0alDu1FV6ei729hna3+Ppz/JGFSqN9u6tbXOv+hVYQZvU/QwoyTgAMiLe8
sbYOh9QDW728OzM56lHWKqTCgTn8Ae27XS++e/8BHIOccRoBZ+gj77E8BkBtNP/IAYxi9JR2bkUR
gCY/G3QnX2HDfbe/VqaMDGWY3JHZtu5QI2pGZ5jbS4oci7eJs46bwNhD1VQe7Tbno3xUP7ZCS7XF
3wCXa9jKl3f0FhXoThOo5PumPBu4mZ6/ucJ3Vl2vt0+ENPU/bkDTcbkY+r0iQNrtCy4arxX10ACp
2f7DdiJEOaVIElCcBvdDd7k5ZZw8lDjkJRl1yEsbV9EWGsyM/5xtX2H5mTxiyiygboI5bTO3gt/n
dtHqA37+8v9KcfLVenfvx7uHhUDx3jXkZ3IJ3TkcKjEWu7qf63N3RO2Fdg8y3MLPBBlk/RhtayiT
qbFobZYGGHkxSjLfEC53O0Tx7T3gZ+Mojlriy+d3nvYY3gdV+Z8wAkv11twc79Wo08n5zPk5wa5S
cgb3WLZJ8riWb2tu8mFs+nfgXcRln7HMAyAWh6l5O0w9Kyqbzga4tLdqnMP8tYAxFnIMUuHvyy6U
ePB2+YdTBjSpV7u6u3gL2qCs+jbOTrS5zLbpYuGluzppZgUJMv4QvGELUHc8T7tgvGqf/TK9JK46
aW2H4QAJiKtVatOY7cyP/JlSyc8vLzhmkm6/0jPE7hQuTtOwMA3vuEfPZ524UrBktSEjlGHlMOQZ
fKAu/Q0NV2ms5DDUy8SLxKuVy6Gq2FSRxcDAtMYmJtGikB9HELJstO3NTkDKyq68utMFRPTnRIUg
anqhR8qmVU36MungrooLJyY1Xq7EScJ/ViyAK+lCZAANFpBXP/4DJKor7Mw/SsUZGoDO+sRDoxue
UInDs/zlMTam1XmlEZu4jNfpr27DVGwmH4Q1+tnurBfVVCY2MuZ5/HMVTlgzYtx5Tye4f08F5tlY
VEa+MmENxpcCNP2v78TMDNQR5U0k6i4MspI2J48Zr1/w1Vj6Imm4lYlS75SvJWkGHqiFL0zaHY9G
Yea5tprz4/4zBawoAHvTD3dEHkYLD+YQ4Yph90tJvx0qeMj8oX4Wr7LfFcu/xqNC0KjZtg/UphnR
6cHqxygsZoQpBc2WhR0e7Aj6rCPRS4XOTaOAqv70h8+z0LNEnZMeUf0G5YQZCZD+fuCyntJdNEoc
uQ57tEo8kJnITCqL0vtXkTogOBa0LD6GIKkQO9tn2PCXWGJMjudTFIMvynnKIplfapB1CAM4mvBB
bJ12wIMy5aznxyCyfMdG/lw3uJRr/j6wSycxrK0QVcchDOK7LOnZAeGc0/48JEJYewO09fAsROZB
UZbmVcpAh4Lezn8No+w0y73/QVZpC1bpKYAMZ6Ee5iZJ38M1a/EMfp7M/GOoIfB6bdbAMtONm3X4
ds1iGBtNirLLcbiSbuNT4BRq5lJb1tIGH6MeSDKoJLwpna1I2a5bteBuERY6AnJVfDQ3VEKV+IVS
ksJqqhNVBrTYM2RcWyN78txUv72KstBh3nGWw5zsYH73ivL6x6amBX/HtwtB8roYjdn0njZHrWEG
NR9JWrKy2aW4ov7LZwTQ0sf335MnqJrGXb6q0HvIqNKUhOTEc9+CNDQzbv+BYF3vfDG3b0Vq4ibU
C50ib3Vk5RVGGvWir0xBERiPDK7tS/BKWqrPeFUJS9bmJrPIfeAkfUKHatnPUJM+VRraLAUh5b8M
ktqSFHr9hfMYwCm0I5yAByP3aIGEQV7o8OgWE96zzj6CBOA6bLewYrgJzRj0Bcsk+WUgyMyvmfT3
rBk3/V0ZkVa1PGzm9YkqLbyQ7Kmf1ofCX8Zuzy6+cyOcECsEVFrFDUwp6rs3Dnq5pl4uUIGdDY+k
wQIg1cHoHMN8rYV3rDrQzYBvtiSga+BpAEdmZ2y2CYpNoY8ryT4iFL9jWeXjQU2U+6ROFUBJThct
2WDOjGlx9Nndkh1J9hUGYpEUFmciOfaH31igRigtUppK1jjYGXsUgf+hotBSvSYTlW0R6wqc2SFL
eL4fjn4zOP2LcDqLNScNub176zQZXJ3DFA7Kylm3TcdnV4Agt0kaaQds/FLDVo4F1H6qboFDQ+vn
9Nf4SePdoGV4C811fF9tYoOznnpXLekn12ETUg442k2uWkI6cSAoDq44Mwx7JxsPvmM3pPFT6xkA
rr9kc8LGPZU6tLwNEwvm9txxXTaGkrp8wgvUFSRD7dOzM5DW6XvZGm76bWQjj1DyUivyJ4xr8QWn
DuF5/wsLzIBa8ryLTgW0GcNwL0rBOqfMZTaY/nxVcfYuSbTmWfBEcN3nO61luSWVIu/P9Je2E8TF
iK3unHAgUq7uJSFjbQem5kfbumgMjDC9QPuT6nyJF9HX7hYq9h6UM7hq2rVO8JwHtg262N6Gbsqx
94d3E8B0fM5xkMvAo4WKMUGRucP3A3UmffA+cfw1dd0muooLYOWWa+GJ8lhynQKhJ93pnHpkvMB3
NgRs1Lj0rOJVxBb4RIjReuRaNBF3MltFGaki2/jt2PdzaGfAHKOTLhZJ2Avv/JSbrUzXiqj2EVtX
llaKzyHDPtloHLjkRIU5vaEaHb275df1k9Kf2AUD6brrajw8eEU9eO4Sb9Cnslp9R5wBWbc9v3eB
6Bwz58TFon6PX2D3W4Y6SR8X3DX61puvkwG7+4HcnN58pLZ1VB9aP3rVlvmXS3g7mW/ZPSstrAev
nyEy6S3naoNJEds2xYAq4zyzKf1oBAyO1ADaAphY/9zJ7xjg13d5OJbk5HM2DsLGafSsab2zwDHq
DtsV7j/1Wi0dFAq1QcOp5wFO9RDHGMU03s7kig9vANIeD/XEHhuFzanf3paYZTRnGz1XpgMkP7dJ
2KIkvGMcZuyYzkrjFzb/U0bbwqngxM8ES39tluJUS+zDyEHeNk0uFnxHA6FTHFulnuSnohkXIvwr
9bwcoaT8ya6CvamHhe/cVn47IuHc0h9TohzXA+a7cjI0A8iqsf7r6bHN4YAekunhnNHw+v7M1n0/
dGw2/hm3xSi5a20dZCDifoBS8YIxmE3Up85+pEPh2C4BdsH0EQfme1txDMg3xE1l9oBNMj/T+WzL
cVR41eqlAvCxyQLuf8GjR4Xr73m4etjEvnmkOrB4H4AUUBuwkJnDwcE4SbbV1fDY8Il5OWsW2wsE
qXYjRwzkvhY53fVky+d0QWQQJju60n/wAaEGUIXtZ04EyphdGYkN7lrph9vgCmGOfv5FNGP1nTj9
JI/DXYr0yC7E693p/h09UD7fx35BXebnYMw8Ua+cl2qiVJYZt/DiXfz/f7X61pmghVgScEukop79
Ep3Y8vukuqYIYVFWHDMeAH2uUHzflfwDi25C1Qv2eZ/95n4cgQK4GMp6dcSSLtJ6T+eihOvoA1zG
GUq0NWfOnG7azlH5qU07RJIYyC9NkElcGBsrHTMEWbt+Ib81hsAfOrfngbAIXo5g0KiMwmQO/3uk
m2M2hILNcbe2/1SuNydDEBS6uI7sj9S/YtgISJacjt3buBXzMHELgMsIZKdBgLgUzHioxuVctuTZ
iNGo/BXhGU1X6XAYG1pHdeO3mZ4Nf19CpSElDXFdadGKPa7hk8d06axFPb2EYGz3VNLQbuDtBHuZ
B9Y3PBxHZ0l7YnDvSJ0K1B6yS/e98l4gt6RFnm8+q4aBCIAQBIkUdffXHCcEn3+ktFk3+7T5gywc
wtd1PfUhcxN5HzNZidMEIua5lIIs0KJL0l5UenwcLEJ1/+jijHBvDmCjEWcF6QBAElOTiIj9XoUM
zEV9wScqCVkmkSRxng6FSs2SYIadyLqaYTbObFUK31ZpZ+Bx/LrBp8/yEGfU3Fsn7a4Ay6Vb4OMD
NE6CsBAKhfkItKoGPr0AFTE3OWv2C1IzpOPKuGuGBr5ubLptTFua5e219GhHMXdDwjU2OdcZnXeW
YE8K+6DZWcVvD5BylSjbOH6PpBqFpkPvQrd70ZZaiiqly75kWSU7HA0MqDnC5UtreeyEldEKzq+i
7fOthxvAT+jxfKd4Ga933xtScA25CitfwZ+NGcVXZF1/KHetyGAHVtpMqIMEIcROHdiqgOaFWuw4
8cu94Q2HkeZ67rsJzMsJNMgWMs7MH+WPWA9kridUiJedpRI3t+C/rJ9VdFUJvdJjtJmmIPyzL5oG
5vcYqEu35KHMGij/7wa7I+Y10dXYkS80KjBYsFLfzFWPEdVg7h5q1XszSKV/oYJHRou/wlSHCwHu
N52kNGvEZP2uYaRIYP2CLb0TjYJBJgmdMVvBNQred7JXNqfbtjnxMbQap767tIfsWXaaznj4JV+W
fNiu1Rn5v9V/M+Bi5iT0emAK1A47YuY5jd0urPI5SXjNMlSwW+VbYQcUJCQpBxKQzZEDTb+wcLD2
ngW5BJO4mSpDqrZFmyAVW+F6kcj4+zTdRrOypMPHf1B8TMaJB0PhwI7GoK7WkDvLVm1lrFHM3mzr
AlTzA/8hw2F4O5106solXoF1Ot22cVu02pyhNorldLQi6r6QC/sOUiJnGzKSlE148TSQsBffD/8Y
L+baG5heQC+4Ns5m1LF2hGKxW2ZWLSrHC2eKsmppcCiMJ2dbJvydEJtGaMNdDkea1zt9eR0QLUZv
e1Bu5CtTLG5JEve2H4K1Nkk73V6qVlL983mRprIy7oFEA1a4f+mVH/cWOJuCf0zrVp30Th2SOzHD
aVEDu/p3ZiZ1JT0+pFwVmZjJXZD3R12kQ06w6XXV8SB+gt9FeFg83k0ttOA+Awsv11HK6R5g0622
i2r1HoTXv8GcygJx6UjCytSJKMOtVe9fdnsCwEoz7axClP6UylAJpEd+iqQ7InCRRhQnvxyuR6D8
C25RMSw75r8ThMNUIw1UlG2aH+aG9GKZNszzmhMFN5v8e5QmpdpO6XmHldjiLuzCxXSzrOjeeDi8
UzU8I2Hai1nwKbjkqdFHJBaXMuI2vsN99fFmlunti8T3yPCYE6yyIKmI0hBdOdwJixUfyqY1L+Yc
2pktVQqJ++oglj2sZE6MiGoxlP6otbnirwpmkrXnfamQpK0iXTHzj+01y7wT3XiGhPSPy3GcY3ft
WF7zMFDAA2XtHQiHlSNLrWy7PxAWKPOi5ItWr/TpINPqHsbgLhyl7D8Kp2bVKTLK6q+iKrIiV71B
ZbediSJ+iFAAQLEJBIgRiyfG8gqrbLCXM0IV8dpTf+J0NnSC8lFG5TyAvGSB6dJR1I06pYi7y02f
c4DESb4Pg6OkYOxL8d40bFugKJXUbIveFEE+BOzucO5ZK+ny1mMWOkkNLXWci2BicqkGWM3SpMO8
ZZJKnOZKfGyyDr/EC8OPTlueZ+Pjcvw+jGGvNcwR13MTx+FJs7Gc9BNOGR0Xnl6ExTRG/qqp7noy
QdxvhZ0PGF50+7E4btiEtvanuZLEP5LYaJGbqvcmCkE/U2kUjHY9jRFqEmAdsh1vi9xOiSesofMM
8xpGU439f0MGOxENhIXnZlHViXnzehfhifOy03QHQoY9FS15K//L+eQ8VxIXfUwj8m3XvZfwSQlF
UCd5UGY8tmvB2eqN31Gk4eWWtmGi9WZFDWSpvQLG5x6LVOebf/5/g3DGk/h/9V0UTua1Bsq9X5/H
+j6E673MkhUN2xq070g/ljKLD5/ZOYFI+Pn8F+eGeMMbDnePm9lgMFSfSKKIWhUST4c3h0Fbm52n
LOcpBrXG/utEYjZrepAmJRTGUsC4ah65+01nxyPPMr+SF/tUn4DutiCO2w8taw3p1Ga2h7JQvtyI
JztxNr02L6c7TJsaNrp6/xXWPpj/K67QscBVkLJLGBjc/goosOxrWl+ou5r2b3rQ8d2XXKr/HjSj
UWX0TNtGwPVKQpVelJo0Jiv9vUGB1r0W2M/3k1/Jcko0GhSFQ7571X1WWq0gsX6v24M52b9FsN2f
2PWy/YukRTrbTDMcdp6y10HtPF6wLwn/Vs+VfuTqeWfmbp0L1X92XUINzsSGxf9a0u5hyYAFFf8+
0AbbyRfa4FTx/P+3xEclHX7fqm22rWBdxvtS9Gti9CpzU0oV0Y8/tWb+L3s3BX3SArVLyaxlafkj
0rZxiVqjqxAfQDS+Mz/MfV96jasW61WtU+nfSw2a2uYAFrYCNTBLXxACUrO89pKYXeRWBFmOLbaA
qjJowbD0F17u+VthddRpAIZ753MZL/0AEH8kZ8WdO3mNtn5bYDEwi0SFhcCYrIsGxhIzbLd7zLTD
ONfn9MBWtrii/0W6R3Be2Wq0Bn6RP7XOQHR9PceFMdrAADSPSrs8FgPh/lfzkN5BdxKWmFaUQ7S4
m1GDOolE6mYJLxmdVX4wxcnCPYUN37Ox+PlPMeszJG65jBRsN1y81EjP/KbLcqfEo+KHgzc3zFRn
GybYz/uMXgBr//v0kazftXdaGkHV8FMWwd3TUk8EKG22gguPixIa3yP1M5+YqQ9kuHcMf1tTO3qZ
JQZ0QGiNkUjLxb4bPrm10JUzNivk5LgbtvgQslSkhuReLc7rp0xs88gpq7qSA32db6+yQX5eIEZZ
VMemw52qCBl4TTv4m/ZL9Q6VY9rJBFbSHEGc/u6wlCcMaHAGWfmLvmMZNd5vQCDt/HKT1MiCaQ2x
9RIFs1GLwzM7h7gREbGVkRln/wE9WPFXaz8PWN22wPWZ7V5XC4PpZ7MpDQQ5SnvWf29LpYieYjp7
LR2hjfrmiyf86Z5vBmHU3cMhRqwRNJtB7SnuAGSocmEeJURHd76Es9Su3i2Y46fEofKHSw7fR+bn
SgY8BV2OAD0YWst/xlEm7I1ssHYkDRs2aVtxvWHpAR6kV5o+Ejbx0DZE5+CKFWxq1omogP9jzip0
O/TiF4+BbuPwXlT3qohSNwdJ31W/G8AS0pq9xrK5vNTwKo6dGbeoSrIESZpMNJv+x/oy26CnW1as
vYEgIq6MHA55TiesYaJJqub2ExmnqDfxbSpARH4ijavjctBgyo2Tth4v6dTMD61IwAbZcTfWlFJ2
mbqN6p98QyBGburo/gsbagtzN1YWtmpU1g255q24BBgvo0c+MkxLb27TS//4SEbUED7r0BmpDfpA
VraHguRuFYlUfwp+ngGoe4J16qFm1GPtCrO8feEQPMf9tRN78ZnS7j8SG15jxgb4QEdACoWo3MYc
tHc1IdQMVOcqAL8057igEayBOInXeuglRMJ9Qs08DOh0gyqRVD6xrGxa62NM7S/7Ih++DNfS+Vi0
oD0Z24JcWasl2a3BsTmu86jRvAStY1wMmwmDYfZejiSqGItHr0Bjpi0evPtOfGCe2V7dRQ/b0qgG
TsfTL4XC+KhZeVZ6/bzJ9/dMmmIGu2xvVE1ek4cSKERZWQwIYvOeEGTJVjsqMYXIoz87Ki3BACGo
98VAYeoRku1i+cBJ9OYx6fNWrZZX46xY+flpfwx2qiRRrroj8EFzd4RZGdB2lKLJ5WfK09YKSOK4
meM830/4Z39Y5gBzme1zz+IqMLJaeSoSZfzSXmlkEToaOCcweUBH71OdKUd/OrRk5QU8JNQiPu8U
56j2c143A1GzIHp5egpb4scajCr2XCzZMSM0jUUWnhTz7COZB5L14YAM10tI/qD3nBZZL555XFoa
HaHtdJVBm6lBjCNhRmvRG7vbSIA3sSKZRwEGOudm1No6iSrBB7bq4ZwjgAEptfBWVszt4FY3hQ0H
MP2PcggzrA2WMw5yXCN2zIrhcDhvyJlQV5NNfSbThpnXiMA1MR94AVWu+hQdORxKJsdaiDHDVeAI
O2O4e1TQdv/tEHgNdAR/GmSFy7zCYfGYGPXZ3c/Bwp6ZvNM3ZYZET7v/33cPs/0Z+k9aDUbrfaMO
95Rsvbi6mWannXM64m9DwVIQ9N8TwF3XDG93i6BuQWT6heuwBloRDqg5qx4fmcMMS0wOfcpe9Ser
MS9aJBPUH6lfKkkne+5zk3lOPzWfrwHhHK4BRPFCbGzRrQt++hBnKEOHEVdV1yd4XDSh8zdY8Nhx
gezHaN2IDDlKmLdE4I6J5Wff/M+NzSN41XzDnInBLdU1hNV5RQP185wdKzmxU6El9PoYj/iqnCU2
YS/bHCPw2NKxFrSynanlSzZ7mZIsm1zlLiXc0KwlsNl6cRMQeHZ7L/lUw/s8kCAC4JImIZDbnvFH
IejXwbAh9OJYa/hJNaMm4qU1WCM7T0K0FsW2Wl7sPhmdNwF3Ne5vBto/ZkQINenLBothdcbCYW8A
RO2/szBnW6uTQB1VKx/EJLmRCEJCnYt5D335NIWZxmsGfclKNnFVbZIKvcdQdl22T9aG9/g2cxaw
jjWtXRD4/8U1S91WXcYoyV/x+BUGZz+637GZT5Rwk24bPHJQHX1r8PMeHM2ve6ZLotDpAbNV6Yhf
1Lottux857EK/0D859Mda2qw5TWN63YkC/0aUDiCU58gYS3XU7ecoTOhYaRj/18C8W+ZlGwQTVl6
ltBTt5zng1TK+LO6OC7xnzj74RDwUVzi2Y0sHpazklqYz+t/Qn3iBreO8gR2rTPD3EqMnwueBbEu
HqeOXehAHnIZHsRHUC7ul7pU8TPyQwmheHyV20FCb9uvsQpVUEwYtmGLsgJC2FIO0YotxNMwd92e
qotstwtvG/57W6L3SMfUEc0L+FTTaDmDi3FdiCqXmakvbdGsO66ilBf/qqvh8YC2Ey2Kuo5BXA8M
it5HQemlwgJeCVs7JQzxGIqquvbUMeFIwCZmB7msuh5dxiBLSNvv3g6q444he1mNXcbhzyVmw5tr
5Fq+i5ZGKsqV93x6ydCjDZxaeazVjVJq4o4a6Neul3hU95k1eFKBLPjv0un66BxXcJbA0y9BIWKA
PitvTEhd5X8JQOD5zNYePUvd+DI2ze8tAl94sov3QNSge8XvmYqC1YMlmLLTIPFUviZLxZMEx0/s
f50JjLzhkvh8dykmW7UqUUuorYjJmVpaklE4tBoKz3VNQkwn8ShunuKqZVIgxHamvOMTA9MJLf49
srK9X45gy0/MHvsBOvPhW/NmiaotSp2rgv1M3roTTRvJwn6xvjmtiQtaXd4hRt5+SRgJRo6W0OKc
GOH4sN84FHarmX2s1PzaOZ/Cla5+CZAb3v9YAtWuswUbZ/pG/KKw/2jkB88JmaSB1Pi7TO+ctXX0
A1X7BnuoZ5ftu6YTk3nDs7PmBpLzO0/0Kc7ZLAmN0/K9nyUnPJqgYbCaAVp4Xmnvlcma/91o4yjX
df3KUX9WPXHZKpxbFimM3YSr50DwSIl5XaU6hqMCUsd40KDyqs7zEn66agJVi+7AK8tDuWOx2+EP
z+3f4T+cU8odV0NbBuJlRZucOxzuJ4ZfJ10i0kTsfRLpmcAFwwNqSD8d4Lan0SzmyHjrlln9OXV/
/vt3q+xLLHMN8XMdVk/kDEa6N14Sjt/MZ8zXIho9U95cvuu0k2CMAaCHOZg50Q3B3FJZaN5YHylC
jjggTP+W6Y9daHaUtStd+zxzRwOAjT8IhDDqQkndEnJE93PQFa19PcpY/q175yGZRIVvFh3XBvOC
OeS4HjNNYZ+vbPWyskupJMIzeHx/FuEWiQOsmmDG365zIZXUVlFmH3GsQKlZ7tIfh6PdTABngH29
Co3Dok/qJET/M1wjHNAy+h7gHb2+81iYCMGhtbxC9aoa2xn4/dWs41pEtRnjWkSAHTjxonkP8WCJ
tXUuaPLYwkI9i7Ia4LA4qy9/PNMPsuEK0u0qZoDOxkfkN3DZ/B0sXgslQFTyRZsTiVlrg+ps8k8J
tVn40PHl7xJlLI9rY2j5g78NJjZkvwtt5b0uowqf/5AQR1dZGQDbUqdR+chRPLlLMtyLMPp/T/SB
CBtOpBjp6digg8/8boAj2Yhi1JstY5d3vitxekn1maQUYU3zHU2hexzlRlNfjFs4FoQ3vN1urF66
5EIrb4Op6j86NP6vrqD4TyvJciKXpCBMu1a/uFXcPAHz3UjSUmMq9e28Q1M62vq2PJZpKd+EyJYz
7BhSoPv/rMh0yI0YU3dXZz9rxYTSbg1oadak6hfhYCMz/lGlQsG2jBbpEUegqV71DDWf9uAtNhBw
+426BcMS48Swx52Yu/32jd2QhFH4GO0lavBw1CDecpHn5UkO2W+cU7/5AgocoaqFoMp0sYDnw1Wu
cv0RfSPKGe2kTTRQYp2Z/MwAmjl4/17QiwVmkdc2iygb4aXN8k7P7x4/AnOOwAfag7kbB3oprWcV
/qCsUcw3WZ95kk+1E5Xi9grv8E97yrBBjZHi2BfuDfJpry6WQl7VHKVACsd2/jtS+DYyWeKTLQS1
9uQb4b4c6yRQcjmBbzkhFeg2ML4u/14iYY12nk7DzQ/S5tcIy7EbRT+LFwS6VmYx8e+zErIgKVSO
SA5iNTaGi2x8ZHr+FhlWyfVddWbdXRsh6bsUd2hncEsdDs1cHtvWItnoPCsawHWSVdkq0fcZ4tOV
CH38G1hQ+rV/a6gGfcsORx7VzPl3UR9jIqZ33Gzy5uoYCX+k4+WhKzPKs8H+Js8SD5XEpVbm+0v5
uOdNtTC7sICv4yPyTMA1lh169bckBo3vTMEYAmvbRates14YJTbqJjzdVdOKbQiq0cZ7q6613Vq3
Z3omfl3yC0YAvLtB/w3nYhBQ9Hj7WaWZVxLw+cDExJ/I1az1qjPETdbIFR7sLREtvlF62EMeVYmm
SmysdrIZj5wCbouno2BnszasuKAolI1eFS6Awx64aCMskEopND60gBdL0kLo6HwFv3giFK9l77wK
CvKjauxMumhSXAxtgMOtlfhd920tuQhbK5F45v8iSrss1TvPcdHeeEWgc1/rHE699JHjWTDXlmpn
vF1WeZ3nE0XdWjfBBbRo3o9qBGrWmt0QZS0cAj158vyE8d6aTPtRVne/5o2C0DoJxKVXwEIJOKes
1sNC0x08rRpqYJ6sQ7/yJY/kFgk+gdKgFrTiNWft8HT7Hm0JXpbYZlgcdlxCEMCJf6SoHcdFlCl1
xKe00xwcB7MNDHjDl3w+2c3VhAW4qkaFLzg7tA3+1AM/XfeARyNyjid9Ktf79nwZRlzF0RMyV0p3
1vnRUwL3Du7j98OdFCGaAodSI7nPMtKVZlDF3DmjwZgTyeXF786bjVLvmZ1Jy8qUhCkmIU91eo6z
D+F4DCEtytjOoSrsSBcuBcuoTfnTCn9lBwtmf5w5chZTgkGqJ/X6p+U0ZKrdHlIcy3++XdQcLUHt
qMHaFxhzhGfoRtQDaXpyxw36YUElgyWEsM9E+MTFxfYfJDyiTCyO8GgFTbfS+Xdx0XGWTwngCvzP
T+VYxxjm3xoVn+3inSFcIOJXONjBl3kN+6UgQsMsxFqviWBIQsn9qiBn4mIkN9w87drtTfnlYJca
cZXzkyPXhFcVKMWqtJg/S75DYd6U+DCcIy31LJ3w8womdUJ/k6wOPJeOD+83XbOqwDYt5WWmNBKR
Wf2pN2welRgUTbDAVlFwtuqRYU+gauvuRFFFZQyWoWv/DdLebDMIMNsdYHwzmj8opP7+52YlVoTj
jF/DNxRCrFZNrQFnGB4SYMe+wpz+Ybz/yxMqCKX/6zCpnSKX+1SdDGf53WeJHEOFaBsb/vu1vZWC
cnJvG1Z67j9R4Z7rWf5G4hUSijRyyeON+JxP+2KbhVfjSDJ77yjoPqIhbzPr3FiOZiYAd0vRmfPO
gkKTa0EaYg9WYkzLXxiR2kugI5El8eR904eRwzCbM0oT0Qu3Tf1JdZyfkZWRTtVk0OyxfcuvtMf7
mQPQyoFnx6QhEQgX0fl52GwUUkMC1B08p3SOol4ZuPCVQLduw81UZE0og4g6K75uq4pof9WLF1kF
zu+fnTfKFyydNR297EAJ0fJVVCdRoW5ZpYyaULHWtAKJnT+kfmMXCCdU/SO43x5F+9a+FLm33QZR
jNeOEAvJ5tbmywAUi9SQ6uT8/Uc9gtbJONfRYyj3yLlHAyHkK6RMQKap5Yyhb/FSnRZibwka6EFx
ahWPKlRHf/k0fr5mpqewwf+lPQIR3PUgPCCePDuQy4bx8qs9Lb/mmjRE8qb3eCsvgps8pE4EwCau
A2/XGW6pfEQb4Jk73iTPJ3ph6xu1YzA/GdXtOMYILKEi25z3g3pf001G0RHbeL3Q4ou1u0tRvOtA
B1nkB2zyfNqNp+WorPaNJkUkV08GmtSbLpueAI4iQni0U1GQxWmf5gJeu1dA7NRs/S2UQ+mlxK+e
VzLctV69ZOY9N42sTytU1RtMRgrdX/4SqxkSUoJxylMNBixpqQDCWPVF0t3gh2HAv8+65KovtoWy
fnEQGtGuXaNEsWkVsAFK1YYSlL3Hy2gBSiaTsmqZ9Sp15btb1MjRQiIY8jKI8ttgt2dotIT613rY
lKzr8gia4Pk1utu9E3xObaTNqkU+nivOYSIrJ3KuS8uhEECZR4OE6gxOaVy4kLiDiFGZoXSqvJIG
BAbe3SJh+1wuY2UWajyFhnPxNLgd0NnnEQzKbrNAVI850eofMGE1UM0/EEszEQD+YgcG1abvM5SD
ctjaa1tZ44gnjiK+zE/4xQCq/xFME39ikTgNtBDH5ygBTCtwtlh6Sn3FY2XqZfV1xVYLrBzg1EHd
pGlZXvbp1V54+UN+/N7aB9X31H9+aVdfHEJ9Hwot3g3ZTw28JGkq+cDBRFjQCawz71PzGxbRR+my
QDc0nqDQvrlhrRL++uqSONtJAHUWPyTXT1IVa/jq/xmrVBmjtxoBiuEucsSEVtwhmrfw7Ly/CnhU
RYT4slLj4WcEtCgIdKlhhhypMAjn+tAGXP4yD8hso394GbchEzMEhcMZLainQXxXkki3jbmxqYNv
12K3pIFxWwAc40U1fiz66UvM8Bk3gsEXhFumYQ3OuXL2rb/VeZ/2NurwO8qU4yGpYN/fNhWVmeqj
2hvvsyR5Cv2G5s0/ZHmxOcul2tIKZ3L9RRkpPfyBF++hs2vuLcwCnbGJMRV6JFVIZ6uhMIG1gDkl
1vVs9h5BrbPn/XimCzItRDcbWp4UnoEQTh4E1Nn22Q9hEaVNt6yTs1ASkRxqGOgbXhnNKP9RE9ti
plAqkDnJvgpvXSC4o5oSNO9MQmtKn1ZIQfui+pQsHRHrY2LUHeup4/cvfxSljdg1EHBpSUhb1/wg
nws2ZxBw/HfpztmNR5Nxcvh2wPmsqQ6pDSRW06gCcUnKJgkRgsUbBLx8bgfnK0RHxjParRHwgLWR
o8uLgwsGHVf9kqg8R/NPf0hWNG54YgVagrjw0cPmR9q6qFCmhr7pH6bbSfnaJoic1js0beIFdKOy
dC5AxTs6RZojgMSoD7cIAy7ckoRRlRo4c7Zs+6BL/1SPDXcoJxZJhO4qQ+g38/RD2pBAepil3fE0
xGqs0RWGGUvk7MDKFfqaXLJSRO50uHju/Xg/L3UPtmTeOBpkC0SJHh6YQx0vl1aW94G5Rektmzlm
JQMd2dvtqKQtD+fqdKoTITNfi6YJUPpYRqQZ+Bu+pmxjqjFFnGmQl2ib+L2Ux2XgWhOHtNo3TE9r
RPDIoMmZtjX4GJyO1l0EEDkgFXrs0m+bfQKhU/CPm5HdOTKKTWHYf5g3F1SCrHfWjUndJ89d9ubE
AsS9fC2ayLN7EOKb/XnwVWxIMDBrrC0oiPFohPPkjOrQNKlfiOPDgLYia4XjZ4l3O1SkWLoTlKMZ
tkrPM53yRrAbgnzTHePUjwiR7tyf/aFXZASTqj2pdxr6F3pMJBkLWTGnR7kyhZ9Dkqze1b2SkGMR
HcSJ+0w8CPf0gDYf4rpFuvEIhtQzcYFMBsMdRCQAXmNvUL95ze0Jo8OcEhGNzOc+EGNrmKe9p9l3
xXaBn9mybAiBYDytH6iBYt6QY3/w1ZeXqWZVKPa8yxGXm6Laz187gMNJ464Nz+LcsZmwptHspsOx
Eeac+Ndp5UAqhlFV/WRD1wKHEWs2LAZfnclZadFAmrItNzNq2+Bm74jRItQHNGtgz017BfKsnhnN
cxjnq3Edir/7znpUjPmBVfQipNtsV8M+AV2GovuV6L6lDNrTUV3RVw6zK/yufiaD/oxY5iDyEqFQ
ga94CsATzAAlZBJco93lQ9X2rzXrOETa0jdweGVfF7G36ROM11QFuzwSWi+uwe4GiEbIdT0mT9XU
CKEZNtncB7Uymzwblmb2XpOpTVw1xQJTaUu+ZVkP4GsowQs1gw1udFXPQI8xuN/YHEUVtOV2pjUu
/u3aHZHioArB9FFWraU+UgdrOBG3oxz31aHTzHFPO69SmB95JQ0vm0LzrZUX/PMfHQ4pMu0mRyJJ
vGjUKAuqMGk5nyJaoW85HMwU1VnROOFlo0iSy1GeLV/KBGFIcIu7VYteqKRCe4KaU7vdiPKedKm+
RaYGXKQKB7mkGkcf4OHov5cRo9azvUbAoucKaAi1e9VfscmcsVwYf4h2jH1LcqcMvvBbix5ysLWA
r0tbdSJcZmnvKoONemPgN6TL3drShtmqSd5poh9x09/FX7bTcJCJFR09FM3SUPweOdRGabcHWred
5Tj8YSx1OAQauLZ6cqgy9qjhKi7eGHRaxleEjlsKd53B1RoHlDnwLGCTiHUPgM8mv+CGkVbOdmtL
qCIOQjCcQyLJ6sR3uPePI1dm9xfh1gRAysr0Nm73ocCjfS1nafoOm9yTds2D9jbpbXFaHzz300lE
zzU6l/QJ6YC0Ik5a6adaD6Y3OXhNlv1fPwB0OqdmDSYBoQ4XNVr1op5AU3tnkVJ+ELjIdK/8nQpt
L7TRjIz2xnBUVNDclsE7FaYeOKlV3LNWx6OXi3rWJBIx2FqIy7fp0XsE4mn9chfQhqtWWC9YsKNt
GGFtjH1+ITbk8Zq7rLo9WYbZb2CMw2eD8GCfE6z/rs3hI3FCDRoQBfoB54rgeBokgvWA9tm8yLaE
hrXFoZiLgGAqBxK3gM/EMQjeDOSiENuFy1KUBW7UGdY6G6ockNnnj7Vk4JHQCSPlDMeyu+PJKCy/
yFeuhC/QY5ZNaDnDfUKcvB/HXPOwa8ycszjBGwja4tABtDn0HvysioG8sJwXl9JEJeQvJRGAnkTq
/wNasw8Vak0w7wFQssRDRcy3iYoBGyr8tMt2YCMVTfF+MUwqsmbTD+Ftn9stKrZNV2mNPpFt/jH9
p8QRNFo8XSUr0rYDhB9GmXBI6fe219lS3L8KbwoNj6pbiZn2qZGY3dWywSE/is6sXs51C/d12bjw
BbM79sJS7gvE4LXXdEdB1Xu3sjRzbA0CM/+tzRt/SwZvJzJ66vLXFrcq3Mxh9hG5vsIly6cjj5Qh
9c4s+so4cDmivjFJ6CJoK8GQJ3pU9y40jcq88etLiXdDd42gQmyaNHzhcuBOoDtSXfbE/OYlxLKL
MJLDan3LKPrkDiQGPIjVc25P2Fa0Vhv5h23AAgeNLpA/nYbqVpPE579zxwP0AhTZ4hwmvacxXGi0
6KH0e8nrixTMuIYA2dgQgFeGlmf0MrpZxlWljYbjNs7h3JnNnRd/6mmZUTUz7uTSzoUdRgtjLkBY
vF1tHZzORo0i78x28vmmOHYTbN0KbNukaJF1yas0IfCHpE3N3SIF9x0E/XjjOV2JCw0EjuR7JQam
mXEZ5+jfxcnVI/1q06kjLIC3mtyBDmOxbH6PyOuGjDVvyhlHAJQB5p6SU/5MW9dxpbBadDNtOOIc
+GrtYQHuYTxE1ZrxZ9ZE1nx9pzUWPtOU9hMLaKu8sZAPnwP2kvQRWxgIAiCyqL6zdq1kNO+FFUk7
YnG5GK56C4j3jsIlfFE/tB/QwA7pXayrG7FrkWhp5lQf8UpungFWJB/YOLCDL/+KTBd1j+sislM3
7HHCIBvSjCf8EkN0nAhtznKCBHt8wAkmPNHoC5+rlFJ133kSB6RP/ZmKqOD9kLipY7tapFtuUvnW
TXGr60LewxLLtqa9fDLlaUw7Xz5hlgxH4njablLtR4EvHTBGVcs7fuFLXY2fwO4GlMcXdUY1o66q
rWmJu8af0mtDkLBi2MGQ7+kICguQgYhfybTkV8UvGxeM7a/+P7BGjb28TJcjuVcrcWrWb1Vi76By
0PzgYoKXPDuFAmn2yxkZU3icWJVheYzafAMyc8XwDZ5kuzTTOkd8/iJB9fo52QMQ6qMpASlYkOBu
TkpVY6HDmkWbFfOVIOhPn7r7X619cQThC94/cKmb9tmEv7ud2KOgAxK+HbQF/ejBKwggSh9z0lqP
i8dkC4N4ppvM2/PHOpdUe9+maHcZDFJxcGGYgjozgSx1hQ9hmVFpUhxVtNJVxAx6719WXxeuBlOf
Z7Pd+rjAtNEqJSyos0uWMAMtAYEGOX2SCkfGtvPtFyYcgRPetWzyvyml55ltfCMH6Yw9s7BS8s8i
iB+CBHUsqIe0IZNYNKNI/928uFmOGgYO8GdTcKtyzF7SeA8ETraiv0gfuCghhw6CcrMo6V7unFQJ
4GUK2le7KzbdlLI1hkXueVkGyyJzH/MjymkifLkNWWXNiu5C9AFQcaeXWe+UY40jSB+b1wpBYCxS
nuaG55OkdOMqejF5RSHwx0Rs/v8tno0cs8pVUElzL7C6wbKC7nlP1ZB9JIUisJoSxa4bht1KQDtZ
L8vx3eu4WN7rBf7wITQvYGQ6vkj34kPcGfeOH2X5OduAOb9lHPGjO/oJqGnkH4CpzLsCrbo/9Rkc
8+1arGWLBHTmvQ4pGjrsMPb4BkQHKeEqaKYZTzs+6o7YfDt/8C9JF73F3eYyLmT4ljVJZ0SttKb8
KzKAT+OE2BccgQdTmr9RNSpFun1DqCXdX4UhcoeVq6cwEx6PjCCh6F/tifnb8IB7T7ipuOrqphiR
1sgN6S+65ROxXTguBH8O0mD2O+PYbU0ssUZHpyexRSOkL+0d0P3mXjuM4ZKkndkvAyIqGW0L89sD
2Y9KCnINIVX3iaKKroQMaoWbnwCM8dGiesQ1sI+t4MHEqa0kUw+b3dFT+zRAfBUnrRcz5uVaBCw+
3Yg3AOzUAgAnit0XkZNEyVWgdJ6TFjjtEk4zLJEjU5QDfXTLkpB1E4Z8sAHYwhVxtwObOk8+AMNJ
XqjL5RsgQvHs5aqq8aTnoCb9JPOHE5Clly6F6IeEWbdnGIfP9o1PlrGHkHXJ7b52ySmtaRJQMlXB
rP7C6WWNHjl/TH5JbPOjipP8brFvwmPmP1tFbPcUCvnzViB2ixnRBG8VmxYhw3jtfnr8fHqmpujB
C35vlHMTPnkI1Vhsbs2OUnDmS4Wo6cvWDp9eyDRzX8wMX60VBBfZXvBt1iM+lRQ5/aZxDFr8ncFt
Qk6+G6jFh/O8XXdMiXircWLtEL8vRRPgrjkFdL4mhWVx3WJhx/Nevx4fC34pT/PDvc0L6DQeBGFx
FUlJ56jPdM66wVEN1stZcyVhrSoFoIqxaAcoT6uTxsEYUaFI0dZhx9n8P4jItf79DK6lhLRNXwu9
ZRsSi3MSfUekT2nIHUrFeiWzCzPPjTEN7sU3ehgqrqVn7V1kkzpu5nzp0w8fQ4pQPBlS0TcNU/DD
h1S8rZRE/+EEtIvHPEzgH+rWgqsW4ZLLq92Wl3uzogJr4lQ2KsghUhBSk/SsD13dYKlQxolaoSwP
swiYkMBVKVk/fTIqpBWVkoyeh1LrBRCnNZbGVU9aRVxXVGYxzBxDvWVWV6MxxHUxZzu6mmS4ww1R
W7sb0OPqkjKjmOt8FN18clG1418T0I6QOX+7Klp1/vB+d6/YHU6BN3BTNKJJQ+s7GZQoLaRR6JHp
voM/ej8x6HWLLre2tyFCg/uJ41eTwNIwK060KBxHk0t6FLbNRtZ0NexwXe2FKGg2DZvteAjQXpzC
8sfCT+nd4t2xFOXZxLCCiPgHtb1xLNnUHOMT5GU/yasJv0NDyyf64GUM2qa1sdRNszVSAlaSvwov
c5P1d0p1fTFC4sOGgSXGICok4ediiVjM9/SDZYoRkhXNV+gqNVmAoUF4zARnI6Fl4CUo5FFKIO8U
j9lFYfhMkPNPbPqygtI9ZbMdBuveoaHLQ2Y0vZ2M3RDk35mUrPucVQKTJBKexFhMhvu9t0X+BVc7
W1QyNs5QQPFZn2KyucZgXHCm0fu2sbSLY/pTS4uvf8MFsdsJIVPu4tYbRhB7QfrXTMf9DRAviQTE
Y9YhVYOlIHqmL5pnAJWs3a/aXfm2/txSvzC+vVtxhrFsnnZimKVs9B5vgn9FwpSv0z6ksor9VsSY
J+kFfoQQ4IROBDrhuzgD+mtV6WHFbgcdEU9DVJKHK/XgGPvFtwMtqEoRqjVLDlB4aNco+AcYnigX
T95KmFW/jCKPACCmKzn8iLGs3T3atozuGd0iMXj614FDOX2teGk4KiVEk5LT+YU27MrDiZAo0PAw
9Q6EkDBdqd1gJVzP7LH7bSvF2aq5BcUD/Pog0vyhvjCh9Mo78rvoeyVqB3VY/Di+fU7Tn6ffu2iA
9BD+iCJkbMZDooZTJRWFhdq9LedLwkA7sZL2SAJueI26F8b0Wfo7u3UCBVus6Jo7dx9y8LVqfY8t
bi7XZwNFPaWni4Eii8ggw2Pwq9uieFgvVgk283iVUsEhk6wLeQZafiGoZbV4H3tdMRwePglToowP
o3c59b/EMbF3KgvocnLlePGAx4S+J0VL9Z2mJk7DPXZkfTBBgvLyT10mX9c8YsrKoUTRpvVkDN9u
FaHoWr/IV5FPlsGhDgb5Cl6Bkgy8GELCqWrXBt0T/tqTKDjhoCFX29YpKFuaQkXSIfuO7OiR4U95
Btjl4bSU7PNNInsJgwFhpbZ+u5oiygjmBgR6mVszMM4LSDEtxD52K9iYX23sIjxy/GJnEB/HozFG
EgyNHzC6r243tufYVN5RHZ+8O63J4U0cRAFosPyNtHh8OUBRYHvekbUv9jUqjYfgCKAkMlswd7W3
Pjdcj5xJ4+UzLw6vpCykmY1EVgivEZko7jv8IbLjxoAnH6kSjAtDOg4rEsxf1eXqww3aKgZeCEOm
Gqs/DSjuUvvT3kI2AYWTGO6v+1t0vakSqBnbFZTw2nTyamTEWazgplNdpOn3BUPTgyKWGYl0S4FJ
FZdhm/ztHYHPOvY6atCGwYOu68xp3EL1OXv83+Qp2Ej9ZvHfAtHSKVPWb15YWIOJUrUCdtN8OGx4
m6J2ouMf8bBwmY1/h4HolWr2F7sr2VA9h2Db4jklY8p1xauqN8xoQ1EqnzG7QmHct6/TrNidNaEn
Fw5hFFy5j5RDwvVp2lYlmrcW19Bbx+gwXGlL/9vmUCXXKauR43SC6+1MjWVSVvrI3lrPBaVW8EH7
qqXLXXr1z3ir3Bei+4W2XWCkV9ft7MUFiJF75UhuvFK6aw/WlkyrLEnVh4GJZXwAuPz85F+ZXyIS
gP8ZCRyT8fa14d12q7WWZEC2XoZucuU89WO36ozLnYtYpgEGC4XtBsqT0ozNITovzqTPl1+/RtUc
GZ7PjHK9NP60QxnXFP2nGny5o/xdX1rWn+POBqmipBW4qrogA9U7/F0g9FATQTArePc358b1+u1b
0M3m+o+yIZMaG92GN+ZqWfkUgifG+zSg01kMF4yEoQG73rZvRkD/HqZxETL8QtyGhUtgwsDWJVaq
UWEsJB7nGV9mPkO+DiEloq77yoqamtAHrZzScKrB4i0b0KbjpiRPGzJBts4yxcxoDevA4riot6cX
hKT4TVjT0r6GilZR6DSr/GdyMutP/zAR4v3g1sfp9TWP+B55GGzy9LTyLOOEd+iq5C9fOkHypoPT
BIr4sOB7Uc/SrcTPK2JiprNZbQSxtJVmj4pi7OMjJCC/jD6T0PtpPXDimJxgf0lzvFRZF6F3Sleo
+QcDiH0Eik5SriXjZudfhZCoFl7B2PFKswQp1srZlO4sLp84EAP6RleXpiOuNSvdNUpQCXb94TI2
n+ckTgo1c91BAwhV0e8NYy/xdlSSF+Ls0m6AsQOmnCDmNfG6sRR52H+oQ05HUpfC5xLSz9P+fCQW
tD3zsSpXeJtQRU3HWzYDwmP6QfdVMkFVcjrawGtK+HhD7K94DNK0KXYDRQ35wzg9Mt5zkaIACHol
MJHq2Cw14Cxsjc9kyWDecF8Al3Snqd54loMOppHfmbA6a5fIaE2FVf4kDTmOHj6ZTooKIQJEAOP4
/XpxT2TK/stQ//nL24ZzGy5ImQVIwaNK5mYOfDk2py7g8IKn95DyFn0kc3uoxrEpaNVq3ALVQ1mO
4ZS660wEVobJED0uqSh4nFjmLiXv4SLXRZrA2BtdHHODUDBVVeRd/yAqULhrGXkOoF/P5uD5ikvM
HkhS4HQddkP7GDOWa43nxqws8hTFZhUHl0o6TZOIXuEmMq2SGpmAnaAVeIYePYDDhwCCviex4V0/
lz2rAFLiyTpQ2bT2a5Cbcyz4+Ko+PPP0gCaXlj5MfMPlREqCc9+IE0lWZ3tmslmVLpKEeRHdWc43
GGPMEbDjk6v6WCmzygC+keX93FsIQfy1hzbaJluQMfD/wtLoiS6Hp3kP+Amhg2SMQxa1JXiiVJvV
fcS1l1f1QRj776T6WPExhXbmCBClMO42OuSueEjKaiOY4NeK4VL/TU39WdHwvGaHkVrQndk3RtaX
Q0jqysYHYJCD0s9SG2qWTDUITe+3rH9niIsW557qKwq9yXVj/UcGV9mNrykYIAW/son2V8Mqmc0d
nvLfaQ23DJ4GkkGHNa77Ydk3RmfZdcZkGN8BqX4zH0irptZL8qKIA/eIpf8CLtULIPtrP1vtYRZw
vB255s7h3x2bP4DUOf1j8OAtN0nvzhrL7Y55RSj9RcEuJSorudvLkhgqs+g2d3Fwl2rTtm5urJH1
dTFzcYJfIrFjr5oaIB0m08wD1IhZ+uKsYkyUon6nbhSP+P4th0VCwuOtS3OEJKp4J9mEcLmntpDX
hfaNOTdKnwdslK0yBQOBqmZ9dxwb4z97jeZpD54qUhA3rM4GEin6gcTGGR4sGnFSrExk8yJ3IbK/
OpeJ3Gl8dRNkNaien6DTNO3RuOjL9hAQu8JBQyOIePEnfZI+jH/kvRHmu1xLuPlvd9V/s4KKQets
WSTfnEOJMqltYyjrYTPiREvLDJJ8k3ZgijiK4GsZGwtuKO5ggyMV/H0ZqK/n4ysux75/qhdgbAcg
OxlhbiQ/Zeaxj7UvLtYb/WEoVJiWKM3f+QX3dmgC0BxGBUu9guthdb+Ra3W9PBs8l/ebjNr1Tvf/
eF6NN1T+li/FseLUZn6E1M3b9reMXN5QhzuJlBM7Sc22oceLlMaUsXp90c9hW/PuLwdpVzkL19tE
rrVK3o0u10VmGnFIXrRyPvQ2Xpc3rUTnF7Hyb8KoGRXm8M3Yl9TkyAgfk1hs+GB/1RoTsXIwFrXg
jGia4XeT4Td3QsdiZ3sToXXUvRtlFPLJ2+JSwnCShjfDerT9f/SxQoV6DfLxMiw3PMknQQ7sTH+r
ocUWXbU7cFws2cfapcu99yaZ3DD6KeN7wUdsFMGOcqNbG/PgOruD7dT73mN+PHA1CtJyaq6NZ+CM
YfswC9gk4sVALeOa8gqZrPOmoOjKpTKWpfFQyb/soOUcne4cMS9XL8QWESZj/WrvQq+eDJuVLTbp
tJNFJPR0dTRmGzcyYFOabeO/oT4sss83nARTjG5qbPmJLfjcfXInr9b2h4TeFn+T7rDda5XqbCza
dG/hPgPLmZgsaeoS7uXU4AWFS3kXA/xTDKlYD/4kGnxifTRtjo9EHpIRc7hlB20rd7pyZSH0D9Eg
R4gqHQITjWSWvKFeoQa0YLL5VGcqnEZtmXpeu2sn8WHEC8DWGvWN+Ypq0jdUB3/+DE9aUXBwKakj
+zeDnizHtXbDKQBh9D0fO7opTzYpbIGFQ+5hN0A3wbwkREn0KIcco6QBq5G18ak6FFniZlZ+OXFH
sEOKjbbFCDGjF5Fe7IwnVhcHGtpAQsfwetQJzplZCKO6Z8ogS7MuhgH6YfNbahwj3GZAT/jCCXkJ
+pRONCrcYuCUn1Np+3qp8lfKSr9auB4YfRbA7EQFIWglGTdfiDy6k+9rtPbq5gHwk2zKE4af1rez
XIxsGYTI/BDGbrxThhNuEtauB5jUeVXc5iH7yC2IGwyi9W38xzhbksDScibyfcMDbv2lU2onFrNs
vuaRM3xnnnV/6Vm3vVNAMlLna1NMkod6ktyyHNer2YN+d0jdeaO/IKHvw/qEbyKRhFuJOu5Uslca
b0urPpUHEU/0+6zrDr8f+O98o08q5nUU8VC4sUnsnP3kqH5362kMrGLQ6QalYsZ3rBS6gda8vq3v
9W/g5k6NLYT75Z2ZG/u3jLV66mKAbYMyosxbYZJOuCBlEgHGTIAGXSi34CQleIcUeCDxLJguxM3P
dSWtSJik+kyv8ieA7xuvS7dXxN16MRt9qAI9ZgJ7kzKL6qBopaRGGUqB9cPA+uDo61ikE5V5S8YB
KTrGU9rXLvB6ENwHW50So7Z9Zwpz5l5Supr255lZXEJ1AiUye4F+Eq5AkRqiCd+cK+ey53+nwOYy
GzllPE9u40js2NUsyFsomkq1rxPFmXdrOf1xvdXsWMDXYUUr+714RqjZZU8Z/WTdro02WmY4suJE
BJrbFlXUdjXZoyFtTx8h2lklR7RZUKBzku3B+9skVou2xXtA0+Cau947Wvc6KESs5aCcNFEHIC4D
uoek1GvRTj9xkraz0MqqzH2Yr3IjrkpsMKbaE1FdIJZCxG7Fs+BWVDRLKvmonLdI4ey+hCKG+Awg
y7xeJHvluT0z447ipIh0zizWzP1ib2nRKir+WVeTPRDpzNOJat4MA5CcUiQXmYqIXJl6EmnSUA1w
hhH/MkZwfbvDiaZbXgPqxRHIPcg+AVVPfM965ulVKeWwnSowSDia2EGYXOH9xH02TH/DXlno6J9b
5Up9L883WIGz4kqhVDJU2TMpBZC867afAcin16XawRqylakKIRkznl9eHiGs+780BpTghwBpdKut
IioKCOTX/Qa1+UcRMGXKgTMvWOLUfeEtUUg+qvAd9yalV+YGc4yIgZ+XPrsNYaAK1TyY+/nxaM9l
//zeOlNkkMwm4V95cPUtmYy/zX/7wIngtAbvMOZ8NspBfyzhaFxiqgYC/OUIp45eAyx4vbyYIDWu
GVmP8ao6HhVzyIOC5Fi7WfTaneOm6jzV4zOweAaKv2VHHUOspRJxaKQjus7DZM9r6aZ5sZukEjU7
92h1S5XEK7U8LtQEroY92JsypQgwbi5BMf7BJ9iWVYx8uVex4BKWZOIqlqsPUzVWUuByAs3MGO5y
uDpNl5UvB1f2L50yyccGkzDzK5UogK+nmctnTHWhH+bpECP1iDCu0Jf9XKp/3WX0GzprxRgqlh2X
KVReE+jgO9Pa1ZWhN8kvlDTardbt0hhSoHrW8hnz3CwI5erLyVzmP7O2sJUv8TSgUdBIVSXoZQ2+
il8tlyxfL+uGRLQoJQ1NuTZZ1fmpOlG98sThvZ+GkVxtV0pRd6pvs/RFBb1BYPQJwR/C4iyHM/W5
PJMKbMoZf38bmgGh+2Eep9sb5xOlpDNlb6E9de5VRrPtR2su0Lg/UB/i3XeemCDVNHKLWC1Izcz2
ZoDvhE0NpMw/3ugp/QrEyOYCEHJ1iB/2u26j6Q2O0iJsYRFbUeGyKpOvfEDdVPS/k6YPXE/PCBQp
+wrwxjxc/O4gZGTbzYf8G79LzUC7BfLEAg6gDWF+U7sXzNj7C/KtZPL7liztJFo9pgZSP0bJv6Tx
cOJx9es5tLL0rsiXFVwTH/R88/5oaRg4NVXTe06lKsGlybobVHHZI9d1mFxrrRD7AYgIuD3NhLVF
WOX2MpRoR8C3RwaI45QOAoEJB4DZIl8HoH7m6nTA/ARRfgregH95p8x/W3hsY4mTEdg7PVV+37HW
MmfANTe6uPhAhmcZ6xOwr/w0JwlCMMYX3/VApa+1XWfcye4CqZYkmQ9+9YMVrY3QZqfiTiptAMMb
cJg/R8/xeLpZETac+jJrPMikXLDok7sNFX5ClEFXICEJbLB+HDS0VtHENCd+ZmpapsfiFNVQx9Uu
t2nRR+BKvix2MFLrhmbwsnMAdBO4CO/yY1EjT/C20SNjfA8epACHRJOq/69nTfexRoZyFLLbsU0i
XV2nJNU0POelIKBA7cWt7SHXHw6B3R7Iw2p5rA2t5H7Qrp0BURvnLAykXzM5Jzn4IpSnEnPbJoX+
cgxNyRaKLgXLfKRnpbEVCQS/JYEsp6+sec84dcp4fewvmzU18qq465+MivKYw9xJGMzIRabOum12
eyITJsq9Xgrkl1znElwNKgZVW6Do/4Dt5Z0TLQf9aOo6A/ZZgVQDdAT2u1PQW+hy+mJCh7BT26wh
rIDDIVDvsrUn51ydClbiA7/BIM9bmoI59mvpBFrQrNS7L96vrhe2W7wuwxsGw0ezLdJYIVMKSPKJ
9w7JfNMAVWKFtiiMdT6BNdeKxzmy8jNh993ez23Rdj4qDa2CGHPojnrEVOPHWtmwfy4xYX2IliG1
3iC0iE4SJO0SHPxgSZvF1uja2ltR/FI0YM7yaW6uSLkek+3nY4Bdrt0ZJf+vCYb1DX/mcd4flNCY
QHANcqpntTexDkPwxsUMpPmTRVWlLRAPPfOCVs1WtQlvNlDw3icwASGT9pQMM0s8bxzDX8csikZ1
TQ/k/bLess0UcZWEebk0hcK4MQNu28iAUurgFWn1sYPYhgadLdyReSZ4988UR2E2wlAk4ilM7W04
Nn0wvS3kCpIur/nweKQU+zMLZ2GryV3iA/mJ9+xiiodpas78uUOrmTmUzvdo1Q6YGf1xsTXiCXOF
H+KXS/xrMi/YT9ii2pBaDicVI6TwfKWnuoTJEONJsT9bE8FASkcv2DDG4xoHkyYR82Pn8M0bx5jT
LZ/4HLW8PISZ7JQhm4q+XKWrJsSsy3SOagdPUZtrT2tLquf9125lY7uSXywSurR/SnXyY7GT1Cr5
8jSpUnh8IEOZSe7dJ6Te6G9OzIadlu+8PkU9ysYzvK6iWsbvke8qCy9LZTolGUBJkFpayOpaRlKx
rNTsviyp74oi7efJ5O6gtYTZnWAzrTgxS9IlXvviWPQ8MKSNtyyYMVnA3wZSS0YiSwAGtJc8NGp+
4KXDGJnlq/6oHDFyAK+tuFGNxVCtKHqoxzlfpdCoLZUZDnMZnpuae9CvXw5gLV1k58P2uN2dYIdd
PrIu9220wptO1XnbGFvaL6na45HSkRZ6CQs/uzSSLnTHkgPKd/dW0OY75Lmct+p+NRIJ45jVuZKZ
gVtEm1k3SJnOT7fVud49+A4OlwIV2obdyTWdcxWOxYJSfDolwhl5arD8jaykXKuAakMlsdBcZONB
P0UUTqJH/MY+xx8MvdsNCdUhy0TZhkarww0HhEinfaj0o2FLh2Ksqn27Dz3bzOrCNND1HA/GsqYQ
z2DZGDftJ34ukRpeG+bZiEDOMDg9H5wy/3nGo/gYk5yliNKNJM8EZepo9aXNMWq9XV8phXNrLibp
mQn4fro+O+xOaWeVlRv5Wtl3hE+VvP0j4nrO1uMRfzcxHKX+IbrKXGKJs58j3Ij19lFyZ5vyI0S+
ZTUqrymDiXKxyr8qk7MfwZE2UmL9ROtSeF9EJMqlgOKbkJChL7se36BlAsOWdMX04wxO4kyFZtHW
vh+gDHCl+R1IXYC11ozK6TdEzVrjp5CJx6pCD9q6OfwmRiWkD7Z+431TgSFgwgsn4btiS5eF6GDB
SM1rM2V5qj9bFqKHYsQ9rWC1kjdaSPUkyUASEIgnHY+nKMGe4brJi62/p+ek4j6Ttibxbhj3mGLP
TxDhrhKn9KT6vuqZS1us7sFyoUq15T2niqopz/QkpFgH7l8N1dt/iSgxoK+rkM7wFcn/+dTE1F+R
51G6UCW/3joe6Av9vgPYxXWxklAy4AAsaXQr+Q9xp0E+TNWG/TYCSgGDan7fwkkIJPO9KGGGe3qy
yT1F/+tIAEhRpKIwMXqD9SWifofsZC0OPjbGteGVg9SBERnnMm+MlgLcUTptt2UpQOJNduZChnr5
wIDujiEKILSYMTe0y3LUr4EfQQ5HBrkEP03HCkV1wpUu3mthC72H0PmXjAtsdnJpMazPZV48GnI7
OoWhVQFAwu1Ev9nVBjSfKgqruxmAJCdJnEplvp9BunFOQw2SIq/4kPekcMkINxeM+pPxvpLXnr3W
PQs/9cN1H0yMIYxLxMBSypiL1lqIqxaSGY/RiY7c0X5JdfpSOVi5zR31kkEG7Ag7ECTZM+hTm4WU
eCD+QWzbGv0esB2ujlieaLoVSRZeydO+pnpnDW/cqp7jFWLKC9rVQUj/tVXEmcIk9MTgKJieqAjv
pCbzz+g5yxzWeZIUBcmmfND57gru8qdmXtQtnARvngyZfVBeimReq1QMve9t8Vr22s65njaMhtcy
CtseAbzkqG4d1gfaR3keCWgvxc/l6QIm9slc/6lEO7RCRs6tiWL/XucAaxqnhIT6ljJ153uv9Cvo
4NZyzonS4GlBUm33xeMMSk++qUUfP97J4wFXYNX8qgfTCksDbXO6bboKnVcn8ok2MF+xGGj5/jqy
d1OUUFCkGeccfwQ9GpUx4zr01mef7/z2x+8/XSSGiZktik9k8f4PiD+44Lwh2Hm5LIYM38lWBNIc
9eXNref/Q0msLYLuH6LC6IF3RriSFMdfDunZ5jGkTuMwWEMQD0AfVHOiq0H96cIGkq6nGTpudEPp
cWTWGV+wG/Vk+liNCDAC4UJLNBmuX+a3iXUcOjTdgnFbSpRkZjo3jHIKy5Ay1SFIpi0eWCJe40f+
fB/Lo7iKDO8Sh/VAS8ZZDkRQcVrTkt4KKsYQecXQfDUgEWsWsMtQTnAObYhAFfHXJ+54ttKSRJip
7IuxRR7be6jPxrRyaWyY1K92ve3FSsdeN2p5qDhHqF94IrueTgcTyyPNH9OEpto7eZiMIBoKC8KI
T/PFIYiEpsAl6holabHa7/3K13tU0FM18DHuIPBYEfnUJibD25Fgnkjy/fx6YOw409mxE64OP63+
zvFN6r7FwHFd4fb1Gj+1rsw1+1OMt3iCKFurpjneJIjsUoUZwWx2RYoVDn66JH+BUWOamOPe1ASO
16NzIVbDCkycKca+wna0F3np016sMrzGH8xcI+8TTRJWL9IMVAEX9E03kNmplVEq3onKFizstIfi
AlHUgUe6t5MCPTQHFVitR1Wlea3HYkKxLO/uKK07u56UB2/r1tE0gSkmA2RC49Kd0pqsTHal80dI
ser5B4tV/1hk+JNgLN74pz/z++R+sP0fiiNlg58nz0PEBAJeh/alwZQ20Vp0ZLryLv0mW5RLZicI
IgR5bF8poVyyBsT/jBChYL2a0zzCOYTT4abxxLUJJMBKPOiBbClcryvwCvRF5SSTuNaermGKtReo
5NvtPalQ2iMWtjBSQSz8Rc3kWZBSM13Ae3ikn96OA4AU+3N76GyINdqpcKMij5U4HljimaoE+obW
9KB5G3Hc7WDYldI/fvyVKFzGTvALgiOeoCKbYV4hHEj8gaIzX+m4rxbZLV4ih5nLah0oqD6BlW3r
eydQegAb1VSGz2A0P6V/2x55SGEyQMED2FpKpwqLDdSfShkDeoktkQk0FHl+vNZoHMzYMMNmobNX
sYlkzjcTdk9SJM7WX9ih8bivBstPrSKUwFUO1D7TW2S8M8zwUtPnP8C1ABalhaqwu83TKGKH+jlI
jxJGjbW2uspnbSTvlWoFNc6CE4VwUjoVBQi30WA8ckSsdEv5UpAi1dFsTD0GgBmp2iqpcSeuOvV6
9i7aN6uocoRjFMz0uXL9Yq/jIbZuURAjMRMx2pzj6kfd9MuluyU/fjqVM/ElTAJIcwaZ/YB0soHh
4+POScQ6mgtt7GWejBsBoBs1fQotOggENruEq8Gu3DLbnoI3rG0FWjOY9iNLNNKjnbIGifwQv6Dw
1Vb1MdnxSVL+uk1lO/6tyedByF4IP1zq/Avectz0flxX6S+d/Cdg7cLB/GbB8wimxYIzxIv42BNI
rBcIGBCpzT4UnMreLqVRzSFVVwmXgRD+/KMYeYPAQn0wi+ysZbc6w6cpCvkaijfoj10t7lrWS2SM
pEhVYojydZwRWsL4Jf95gbGXDlt/bPWGsjUHqdm9I9V54vUDLwSbQurFMTW3l4TZZET7yUxACUle
x2AAVaO2gYEA+AGvzArEMZrQfPfrhGtxPunumlf3Pk6h+AIA6rJTD3P6iVIZM3cuM+9284rH0ThB
bC5G4RMew7aFamV5c70YqL5oR4BYy8bvFuJeuIuEmTof2MGUxLgWF786lJ6wR+xRIoEVmGbJijZ3
r48xa7whiOPS67BEFhGApaAfuIDi+BJjjqMZgJJW0AUuDlM2QhGEzUX+puzfFNhe6wEQnPab4EeI
G3ymhQVbzok/BeSPJXxLzrzfkjt0mzbM/gLnHisQrnT7dNj3ftkozDqNjxQBAZ7NaOIvI25/H5Ay
ohtoKi0RpaVOP7fqn/J2yK2X0B06EWHhVqcTIut+k6OhobnMzdzrUWuwHKj89vfRfQ++xPgo43HC
l2Un37dCeIxkZjVAmTqVw/hPcBPAQz0qr3qYMwuJfZlBONfWfHHWfstJYldj7oLaioiVjLsqDrQZ
gttjuSUeOuck4jZVr74bBa+bkHkwZfaf8RAgmTqMXp4BO5xC42Uuge4H3VqYl+QUNIYjsLEk+5QM
1HO5Bkn6U8MHpww9p0WS6Ytey9jNYaQeYe+kJwP8tGCIfjgF6fMKOGIhZBV8nM49gJYl1X4roVR8
NwkKqeKruGZ+mER6vUi930LIVKmir0hP/rY2en8Rt2wlSsJyQWJuD5x2yjuBQDrxcPHRsq8VqNgD
sS3wVo/r9S6Igi6+J0VMUqWLFG83MYFpB4RbjHxe2x/kEKc9ByjJS8TLuLRS1T/pScFMGcJxn2fG
bcs2AGXgVvbOp5PszsjvDdKkYsG+JqnZpNYmmk/I08OEBBcjfCzJAkuvMp5qfwOW0wbt7JP91s5D
NNaVdKuNDcxCg1yM/waU0mmZax9vloCC2Q7Jka022s8AgCGOcBVb/XEvlc2vxK7EXkPf40fFV5LO
ZVphge3v39OQXvqJ5xtiHReoYr5Nt5AN0S5kD0ew63pu8nTbobPx/fJ1E1fKsq18T+zo5xf5+2dv
E1d1l7sh39eyjPxfMGtsJXajOkJG8HEjxJ5h5WrbRKvta0Xov8hxPB9vP4qTFiN/+VztDJqIy/Ud
f6uZ+80Ya2uSzU6iepPUznmpRem0HggfwtyikR1Bj06XFTJw5ZUDT0fpBfw+UVKqVK180JMROr0k
dTzXNrBcHcdnn26LFuzn30fN8tT4x5eSj9jis/R2Y9kS4m1IF1Qm8ya/MergW1yRt+NJ2KkAt2Zh
Kj967x+nfsmoWUt4EWLNZQzQ6gCC5lKJzXyBHmy+avRSFHKJwuHswhCz4r16G3ovoc4vluuJG0f/
VkWzj6ZBT5tIYFTLxdy9prKfbFDO5S611fEVKet0Er2M7xMqhBHq/RHcC2yishXNbdbETQVNzl70
YoMoPUtk9XuI3NMLdlPB3R5Tv90RVtTDOgOx7aJ1mVXrKsEzuPQnCPfcMtA1SoJoz2cYJzGkkjW0
4ekgLJVzdyCHNLT/5gUtbW60kdWK0ILIunyfRFIOHIcm+k9zdJFCdEfVrBfHtaOeVprq64CTxsXV
Hy3/pV4bbDoF4rVRk61dAJaCY77hdrW/KvzsFGhfpis043T6zHYYxg9qFhdFgFuxeOq/Jo6uiXJ8
8hGD5j8MXQvHEs5KbzuNv+DRIhUMq7LQ4lfDrbIdo1mKX5phWMSI5sMxAqlO4neeB0rvdsqgvO2j
GqJYBb7IiyddIDY8c8jo4zpPJCzyJL/Kz4YlqqVaJB703QdkkZlnqRA2PBAF+lXMXVEC/3DQCnSw
ALiEQoBFb+WGJ7U40PqT//ZfV2z/87CItPYbfednEoqv26ZujOWeBlaiVODe40NJudETJ/s6ojy5
bl4IO4/VGDybMX56eo0o7wbWdtZetZfZCVYPI+rrellIxnaJTtqlAy4Yac0H5yNYgp24dMO9F4P2
XZ00+MnDYXWjFcCa4gxoCekwR4SP+LtcazVQrSfHev7znzJPFlAFP2sodoU4jbDXGfwnJuYD6Zj2
HTxXizUOXtQFerWd5DFBprdDgLzfWJ6w+odb5wXtBvTCtBPd+P3Ulp9dbFJnAmlYN/N0Xn871TKS
4N7kujUfuKyZQYjGAaS+rR4bUkCPknKtCXohvz7e+c+MthO4XRz6tQWKUKks0mYc7tt9FVf6/v6F
LqvkP+KzFUT1p8LnaNLXiMOyyCLZ3uioLiemzkwgkPIApLV0Bl2YfZSgMT4sLfv7RVkuyqDDVMLM
7POr1h3/iY07I+lxAv6h0xiDVlIk5g4opsuMHaFYP7kTH623sVBkY4rCPUx8WLQGinEEJ+gClYjg
toUKxqcEro+JImbicVFu+6/Ly/f6QO5suKvcNwk/SkIgngzEbikOgIdZof03yzDheDdh9PBegrfd
2cyz71MYmQdEnGQ1AMVztGtFHYyvkVSgMkGHLgLF9rmCAOYez8TGketBSINadMSkIESn8+VlkYP4
WNcZAXYNPoi3fD2fA/VbdD7i3lgr1TmC4gR5yUQBj1y55nNfBGdf6sLUgIity/6VCLgwzdqyBO4p
oFN24doAnYwwnO6TDhjmVDY0GFl6tGYkoKqB78O1NFWHeeBTlul5TB2u+ebFaqWhyvBuDFLRKID2
96jFkCMJd3Milyzvc4yLASXWXYwTvKLSFeCXJ3QtDiEWmYq4h+6wIqMXbJL8iXy57AxT+Uns+CBs
6KFcHDWKGZHinSFI9ageEjRTOD2N3njswgQck8XqST/smuhEa0meK5HhVVZupr6HQmXfaKo2VnTr
5DDmIMqIRsMgjGq3PJZDY/otWcpW7v5qSiTj2UWBLSgAoNzVZiF2vVORF0jCRiuO5wKd8WPmYI+C
ht9rzWEtGI6Bs10mKwWU2GhLSJ62Ht0J1Ou1Qr61+tQ7YOu7WCtR91IGm6OKLADdXUzltPiwELSW
D3NvG2sKExqhheSUmgKmYGBtwhxCe3eGGrD6jf1XMAlZwUfFUytV7BrQG/zc6WPntcrgZPFC+k2a
c1m3/pan/imw42XrAgUshgxHFok6bQdWb+A2yhOmljd/YkUdC7sCMW89cvV7l/H76pfX7fss1qOM
Z7Mn4OtDZ1q3NSIyqpvgSKq89xNfYCQPXA9H77aSvLzdiLg5GzqisIv5xXKtfy0pyZHbYh153wGG
m7iycAFv49vl1oDS5ZyclemMHQImwTEzQo9UWHBhkomPEDfm4YVYlMCNGPi7/7t3kO/EGd0PS1Cd
YQPAfuRWWDW1oFeCWtlfpnhKPB9q8qaiEkCYNruFP7tqlwPfNvXZoY7mzdyepHtCzX3VJ8w7h0Eu
P1lYPIEYUzr48iw86oGzV0bzvtaELNK+0wbl89TBPySud0Fbw8HKiV1705AgNnXes2lFjZcqs8JS
9TKVPzAe6+EQFgf0/8G32OXvhLFf04xEp7mqRkn9EQVAL0BbmwTlUjIwj6uXdIb+Eez6gbP53Eby
7MvDhH5apVO+h0CAN9uNiRV1kX4Z1IwE+sGHhnFWNFwrec0TgidjcGnewANZ1Gg7vZCQ06MMYzSr
EjWGw0fUiyTz0d7zbFTvSRx4TyBP7z2X4Kf40usQChLQq/CxweXlF7sFev4eczTh3GsfBiglbNSU
2ylGHAmlJ0/uTRKFabb0Z8E++MjiiC4t73OzboG3kJ+7tCJjze4ne1X5O8HaNchNQRSZZrRLB5m6
7TSo6I3WYGTpTkRHFtcfWB5PK1zd8uOKsEgndGKLJB0r33njDa903NJCUVn1sgrCLWND8UINQ4OB
/WY0AovCPAjHEYqg5r9jRbxB5PLwnKQhS8zVxxC1C1mrdaC4f3pVYrI22WqqfVBi8GxZ1F1s6m+D
w+1NVANraUVngTAtaU7OzfeisBCaQxJtOQjtspVbPtOAaQ2WNtLb9vEIodkvPZzxpIG2n+U6Kp6L
DSrZqYRztWWGtEI/f91kmUr1YkZv1MXqsElU+jzlqGoP+HdCgtKwr9cOfcjP1Dx3rz3RxHbh8K2V
gJ20FqGq94/1PIB3OwZZLeD0XGvtgYC6wA28dvW2XcLnAutZnTTH8hl5oR2rpVEI4jO1P5wVT3CQ
8QArhkgj6/xnXvIX1X0bh2MxJ9AKPQkCmt8h8glHMuLcQAzN8IbcDemc1tMVG+cYvU8omT9Oqib2
iTniB3tWtfqZYjeI4wkeOvRsn8O1ff4MNtUXOgeGagKBA7zb5agHN4bLF8ZKFmvux/+aakRSKQ1c
OdJp9VkEKXElGpoSQDJCw8yRYKro6IsUq9s7GbchBUFeALWePmo7HkA63FPlVY7Gf0ATboQpoWBl
iepEvf+rHLT7nEy3nIf/axJLNeeJrsbDD72NU3K7Njm0xZL6biMeM4Q+uFsVmCP5J6QKC+NkjWoN
cPKw3GFYZeH91LT6Ypv4Ks+ap1/y0yq2okAhXztWFNVGsW4DfkmByoAHdpboL6hFOJdj51PRNIkH
Oi4K1JLMJ5ZXoqwyjsqR9PFMs1wVmVeAZ0R3ZA8slWN5AnNyv9jfRrIA9K6dGc609746rd7/2Mnb
PIZDHI0yqgj1ZKuTfEDNkzmQJCFDd+rFlA/F2ntk8HwlEWU0YgCGH8KtJa9VrwsH0J2/SShO4ZlR
8tdma7470Qk872kTw6FIm8Qfq75d0kq5xXl/J8g1wcK5YFjVyvLVwDsDxnt1rDkQuFDwTcos6q2p
CBbw26471SEDhcxIe+IUYBlAbFBQMO31Sa0v0ptgqkJSP6hGyJNlfSmTi/fIWVX2n43qxNovqV7Z
axqwQj3iccOeFxisT1wwPnvyE21FmwXHNj1VpNhdakjCRJ54sE3xC4R7FUKTiFqJ2xOjtaMh7JFI
VdLJPrSEE7m3cGbNs5H/4XeKlG6sKqisCCYvPs01PqBGKvnoVIzQTXemB4erzH4FcKAI0ageLFon
L44qG2Kn+lgRAnh45xGuJbnzhsstwMwz3QPXK/n06H9xcT2tpi1McZ0Uf0X7zWwjra5W1weUxdG6
99evSikkvUdmmjDyL+x9klR9BLjjjlftmbUUJv9jWEWNDQ9Qsxm99HpMxlspNu8oihm4lA+HytbM
vPhfv09ZjinGqrkgDwf2mmJ885mnEYhq3JLufPPqbDpVxszlE3G1j9scRuAYGEJ62bUEb+FGDoT9
hI9lRDOTcfYv2+A9Zfz/wpuc3IS9M8kC6467SjtppNMRaENaKWQ8FQvgsOHDUjXZ6L+4/xHBASEX
TH1SQVtEZwRc6VSXEFZ9L6F4le3gn6oxriZc/JrtcUlXH28zdeXFm/WW0BLDA3T2IbGE8HXLqiQI
N9Rx4XQMoBEk/UIANELNSZyehJYrfw2sd0Lg42zyLNvHQlSYScQLX1+IfhYHSvKLDCuksFELvLoD
WZBduxxx7nBxrocjtgidzxkgTLOSS/KGZvpogW78bRQb4mAJA+FacP2c4q3qvXV6ORSoEwZSLLIz
qHYnP8YtWt5hWG4vdkGmO3yByDatbsXhoSrZpQdiZiWef4VLGzScVgtqmJ7j3Lwt4bkAIrRnysUB
DtDVEQdIyJ3fVFtOS1YTD1ltCVATuBEkcqGQZ+PJeEWmnfLe5/1NkLxBCKOnA/ci+TVgfjszbf7U
p2ek14Jsz6UotyUBtedYXUIUjhLucjB/59hh8tZg55ROuxvvEgG0dJ4vnjxRZqNc3GRHmIBbrB+3
DQ7qUSUFdz8ACwkEYbYRtQBcDn2b5SWsIjMO+X4cqrsU08BlQd4o4X7jf2geEXB62rYZ0EANtXcX
ROEuzjJwmqjr0zocyOiU76Jy/oOp3YY2IGsTEHlLGKQnggIniz1RsgRExWiH1l0JKwichS6lCQ49
aXrSOcRj0z+XQUpwxo5QO8h6qoUaFbCUZOFAqTSmcHYb+waDt67+7+LbKPcyvKPRTSF9xL4w6awD
CbvuVJcg/Td4lWS3VCeXw+aW4FP1sysHpMiEIUW6ed2bgAawk/lPZxJ1JNsOCnuV0/gO2SPwsnni
TbKu3gcNGESdEgEcxWuz+AimPAYKKdiWYevtG7ZhAQT2kpZwX+cPbOXzc45EJKe5+SOo5R0hS7Ie
JOvfDNyRapYRcymdfU0QtJ83hv4RRfo1hEsZ3QYLc5qwnBF/voGDy5IDX3scbCCTGEpNEAGg7zgS
eQt2OjczLKxazcxgqH+CthVRm4n2fmedyqnDTF35Wf7rA13WyzP7TwFma0/GHEuFE+5ATwEzKjf5
B5kZTl/5i4hHzdeE83AeQN0x8e4QhSiGCspLt10+7v/bxEeR2sn4KFs1RTBJFRuk6599HmMDTDbs
95cSDezrxyU1hXR+y39kulTYOCsrUQJeOmuKjXuYTco/ihObHOCqlcRECEXvGAcERAJ/p/MZMyWj
TvAAI9Birvsfo/N8KcBeC0fWoaMjWhUL9jpyqFBuPDWngRcDVd2h2FHHlW97SiPtXFpRgBaENWzv
CE3HSKOuGHaniM5LocpR6IoTBHY1FjbP+G31OttfipXEB/8JZApCk6Cui0Wl0+BzqsFWGP6vEP5o
XkUyTxQM2eYu5fa9U+7jFvtGJpg79Ov08MbpTX5AEGxecqqrD3UWoPNbvW/QrjB1lpqSPqeDt2Lg
HCVfjFR9ZfH3LvAZajykQ+P0laPcNbXjQ3i3etGwR8H8YE9CVAVXY2yVjbEbK0hfw5BiQjNi0CvG
EXj/ulTS/cpzwYKAxHsXVCxWRN9S67Ri8gh4AZA6Gb5gygwpdJ4uPUAXcG+ihubrVj6V+EfBfxLD
deZlyQb6CowA4NFAMmjVXWr/feTyvQHE8KVXmgUfQ+9UsMH2NtjcgRqXJzMRvqZRSQ5HxzAUBDZD
lpYWqOb1iwMXgJpEM7Hgt/wn9BIf3B9f3j0VqMH+7M81x6sMwglsTf3HFKMhiFMz6AUbWgcIfSFb
UYq8SIDz7N6Wswn1nmUZrNtQMTK4jCRrr+S04lTaln+c7BMTOM6YIKWM7rJEwfWk7OouE4qKPw88
n1evQU/BegEQ+iLJ7x3ivyZCdTH/CUsJDLvAi5fmcv03xd0i3+qL3z+zfbgBHFA4hcQ8uWf+TNsc
9U3X4aMkZhNYWqW/6cGB/iElxKRXHnrwnQEKexlmi/CNk2R0cXppxCt/yg6fqVXFKo/rZ7QBZxag
zVMAzH+TUqgw+Ujls8S1pY6sIQshTmzvkVXiLnLUH9Oszs53L0mkOmYomDreLtvAt89PithjvQ42
RhWteDsH+SKCn5Tq3TULvmfEW1i8gtAocNsgeB172XOFbSiqVG0gK2UKg904k95VA5skPmEXk9gB
OvvyPrxykRQ6DrQkAJCFIwa2o70bBGoGMSLj/Hf/0i+G/GGvdQgnfPNQHpfzU3O/Hb1Fy6qjEClm
woJ8t0l3GNn1w6ztLM0iJOOLDtUYi8YuzxbJRElOPWfVtYc7YflB7VUriQGVsgpv2L0s/TbP+HED
dhQam+kUICgfm30ge+xJXBvzjuNRI9pyh/pVHNZ0x6uXnVWxIxZa3/V5Jx89eBpLv0pbp0De0MXo
ZhItXzluMqqtQpH26iVsr0zCkBgZK+h/gihV5gHi5VKwn46E9oDr8wySvL4vJlunrnS2NPs8r4gR
zrtHSqghSjdrVOXdeAJxt0d5Wuqe4hq02MRRMmAG+qUEqCB4G0T75eMuCVb2ybayrJTZuQaAR7Dc
5mgFg+OprRmINjlU32PG0IhPEB5bRSCv2H/mPb3N9iA/QObvpnH/CxqCEFjMjT9590MW2xF85Vnv
aOmDKazyWKcxEqg4lGyxJWYaHLacZdyBBWYRobNP3xqRYNo1eiADGxO7M5l/uu9QlzjttryO8ppp
4vbWr+Rg9gb+ig7pev0v6hnaLEBLc+EkHdhmnQicvROPkn3r6znjGWYJIqYFdrBQDO4jD228G01X
59JGP386h6IAChxu/uF/4k5C6HJTtr51hHsGHLf3aPONwzwpf4lr1G8zU6dnAt7hq3+f8NjLRwXO
peiAHuYgW3l2EOGAII1mZ0STyKT8jk+Ep1FE9ZzLxNVmDWFmqbn7La5d1pQhwkB7IYbV3q6N+YzR
cBpVWsUxzLHwy1Z04Z9KbgSkDKU1VOeEmy3fA3JIc8YPunQZoVRKqiWNARigDXzIwBkrWla1vCMw
ENAxqd6ARGha96/3LmCrFOueQi7QnWT8tgBHZglBjElteDwjdeMwtsx8kjLNosGmbjdes+7/gOsH
cCiPSpR3MVKVKznCNaxruaqApoE5xPBb4D4H2wV8SC8OWdQXN4SpX64K0LoCyvZEqZ50Oyabbsyd
Bs/FRam2y3yrQyjebTjZKGWPZHm0Xkm5vp6F/NUaMOZyhWbJHjF5HjU8MclHzmiQC0+6bx7LUA+T
2qGrl8Z/uutVDvtFoti+9tTaYRnwcHq/H+N2Sa0QEcDfbwN9nMaithhRC+IJkVFdPYFt+iDfuCCo
59qw2Nl1wItRxGppXY8OHWMFNvzLSXdBWu1WA6WIgrIa6lrsOc1JMp5Hc9laoRssqkCijhaVBYMG
L6VaFsCCgpiYEdeTzmCp7oSRVGkWGpeEb3pa/XlHcyTbu1gXAaix882iNRn8bNLSSVI+WtU0po0u
z2oC0hiUOPe0jXSexvNGNEysqwlD9AR0DE9gDIyAmZz+6mXWoipRqwE3aAjkX0j2heewdZn0m1JO
dCR0MoocfI1hMIoBDyVsGgA54S0Q8ItUeHyLmdAdLuBsYUV75/7tz0d8aXUn8NbLormKMUz4fLPb
tKHwCTdo9S+8x1iZ+g8Hzmof1+bFrb0T46jXPT/rf8jKL996wTsHBElksCT8+Tonuj8W8uWG+vSL
z4P0RUTi7JWkS1VdVYhWC5vx/k6yZOvgufWeyFv0UQ4TvmUHx6iIxQuob1841+sCu345Ohv0vrSh
lwmINoJz/NleKdOhaBchXfUykduv9C+y12ugXR+v3XZMOtczIkgkOxkRMUN3AObSBd4GgHPQQ9wy
OcHNGGIA6boyaSxVnNR2JAFDnypoa9DXkSOzWCRfLlTlPXxovLblSfAnSF40rKJAACNF+fN6BIWH
Tt6o5Srk48buLasH7k3NyV+X+4vVW2IDGOIudlBB5pn1hEc2xOy+G1vePtn5G9uERQagtUGfsN0t
S1xragDxPuzvxtDuduKIXoMNh9J0XQhRBKbOJrYvOiuDSQ945MTqD6vsSB59pF2fWEDGyCljwXT+
IVK1NV3qIRSKII97YidpDXqorowul8q381VLM4o9GUrudiSf2DBud219Mfrr9A9X0cgYXEsHmEn1
/FlSUV4uAjJkE0IhvpmGSlZSUCCr7A+SWuAIb8GJQkAnagfB2PkucGESeVcprCGn7hU9lf1fNrIX
bJJYeVsVHsEd/FMw7qsOZRSqh/RpKPG/263iJdr2vNnHeR5t0T6fNLNRVKbCkIg0fHZqcGdnl9Un
HYuv2xVMACqtjBtZwUVC+uTHk2q1m8bwkKAomXl8FfKO6kA5YVF5c2nget4O8DEJoTTmrGZbrT90
KZBYN9tVyIFNs9pGJgwhVJNablykvIbIp1Y6fyxVqVXjwdgK2+cySq+3kB3hH7Jd6SpxDlzCBqrk
+SE6wuSLGDEp71SO7JQMDeI87ocC4jnv8PHWn47Wn/tfyP59GU5KREgM02A7B65d5/ioOUq0FUua
0nNJ8exrdE2OQtkILZPenMQ2/LQgpfuf59Nz9UsZQoCdlI4h1CZThzSap5xRIO2KMumoUCkE3SaK
dmzIEaa77tQ0bjmFITk6wtjme+F0GctpDYTfn4+8h1BLkO4Oj0JHlkd3TqJgp+ICKqCr84S73En4
afmFtdelux4k3GprwWu6AT3SdEHwf+kCEXlSxZig2Micmw5GJVt1fSd+GEQ+Ri1q6I53jJqeH4TN
WLAe5ubFRtiAnpECRXxFitJr4bvpuVkZUxoneu9T+u93FbPmR985J662/eoiSiuEIdOuwr08NADB
/w4sVmguECUh8WlON6lY53iIo7J2Mwo9q09UK53cfyiJE/SGUUiXwvRlLtjvpScxb2iInmetCXi9
1iB5TM554zJ4gzM7dZ6ykDgeIpSBdDFvqVGafGVQWs95Mt3XGknZz8YmlFkarzCPaKcKQwJkBkXd
T19KPMz79/eyLyk7PRXfOnikHV5JF+fiC7/JIujkHSWlxaJwF1rhdALQTNRvVX8Nr47qFne1e8ay
zzQ5F5Wr7H8GslZxyfJzcbCFQcYq3pql1vNLmozqhCzTPmo3TYt+e43Ku1RaNoPIPywANBWOd5AB
CH/kGBvc7kTKTXyZ2CddV+oD9n62iB48lzxNYgY8owjaT/wqw3t+EAt6CFryyHB1g9meSCBFajPX
vYcM7tn7iwd0NywfwtrlZGcw8JcQDRvTMHUK2IAHk7IeickdxRsOFjhpYuivRW15PvCFJ40ydtpW
wr902e2Q7Kfx252ICw8oFqNgXo+P+koPLkD8gZza/43pUpQh78fCv4V8nQwLM7T5SfRQt6GwcG/W
mqV9RRHMaD+NiFQcyj+KZUNavgbz+SAz+LCSKssgG+py3S7+Uy+Ows21EmQvSmsTfSCEqhLwE7jM
l/HSsJVDBJF1CzZZlqdJVzoeIFmYjJe3tFglP+586D+p+5EJ2tn4ApLpBULLDqOERhuKBfH9lZU0
rG/dvDEP8tVLEbmd4qqr12F1D+nkt5rAx+90sP5B8ReOSwO3QmMGS3MJB9SZwWkQR6ftSVE9jIXT
lMpiFhg4SunjMk+BD4Dvf2n3Gs45+qeao/pecyDN4p3YYAoL0/iCFFacal3VM+lgPpKNL7MQVP6T
gQsGTV60LSFQsw48jf+oU6CB5Un4Kj7MYhPTTUH2cWaV51f6/DaGx+nMEKH9idv3TAnKNj36OFSF
act2ypgHNTCeYNNO3DXlDgT31ioqzuIcSZvTdg/bI5oxcU/G/N9dZG5tq/PsQPIS/dCpMuc705k1
L8u+BhUIa29p9Dhl3Nh3CN1TQVf/Kwi1fU9MJ2EZCe6N+adbwMuPoCG89sVgBwhMyOP3kPJjz6Ue
qbxMqqdocINDqWDhZo/HlMygPwQsDqLnLUenZJzoNuM+wOhjPl/i9nGJe+MoTRd3Br8k5v6KO3K0
z1Xc3Y5S6tRw+YR/gYWT9izY+qpmERI3OsplDTGa16TBCpK5tZ/QcK5CI1HefDHPxZ+szAnkrpdS
ok732iRSQNDMbgRHKpaYRYtkPotYTivhaKDd6rfICUvtkuHL6U9RpiOgiTsQkpN2b8ohpWKsPw+F
Qnm/BQ2pUnGer9Yy5X1/iAGABAlQoaPMb5wOhEVJ4yt6dLeVXe9cgOpW0JZlp5M+GSoU568vFuOM
V4+0lmV+8bDPN57P2CZ9iP7OreJGUXGddEVrOhlpn1Hy+D2CE2ImCY/NK808fxaGOXaq1n4L/1Tq
/XuYy33Fk7HGKWqhrDXKWeSa8+4idZenvE7S68KPzJra0ae/5JTfs2NqmZ1xrNG86cvyfOsfXpEb
aDAAyvdQWL7tzgPZSeIQsxeHssHk9BAG2wlNXG3dNQEa23/uYFp//o6E/dM2w21Vhg2+DC+t0hDB
bNUSt6u+at/UkPeMyF2Rxc0/7nafr9kBlwgzDUvoXSp2Pwe9Ewzwlx1NpTaQ+OGsLaM85F3CDwe3
Ub8b1imcCC1LkrOx8NMVfaYPD4WIfd07Idl9Xrpg5u2tBRcSC7eyRILbf1eTpmHpRhZrhTC+8yDM
UB6SBFxzN7nPbgzJ17LPpXmXPTF/wFUdMh4b0XrwFiDgL68TpkQZV1gQ1cCgJBY7JrJ4DYtS9FxV
rFUIAJyg+PMLSZpX2MVKR7q+BCXZZcy4z6o9IrPygqKqc9JUV4RK6NF8Kp6UiHAHdSOWUGW/oNIK
FcmcRO0m6K1pmXHxu1XBKY9QTvBts1hBHBOmFBQADuxQTHyyk1wKEwIxZU334odXENGkWDO+7L4K
1X3gtPR2MkHlvmKXfBUuUaNYkDY/xbwgu9kK/3ed8gDQRJjrYH5l/bHZdXmAAYifGbGoux/dFfba
IqtKUe7xda0g+V7SZbNSBYeP3aLGm1CVsA+2JfhJjHWwe/+qXuGbPQwAr3BDwJ9nt14QSl0IwGhA
vA0nYqj1+a/8/K3FgK9IqyHaSFpt++1lwXQU8lFmvRHZ+nQpimNpOzRlMpcxMuMo8xhSjDukHEMB
fp2Figr9aafg1Aad8TDFQjI0LatCxLA6GVnALVPHmGvMarkJ0vUdqMMFm/yjtih3vbQxRS6kJVgF
jdf/cpRQLvKfwzu0Omx+DfBDuYQLKhXuqH0BlDPvdZUDLHqnpW2XDbpcR+i/kiOpemT7AynzjjBl
O0QRbuyRSVCEPG2JbHPudlMKm2SO9/14WSXondaz3iezCUrZIIoHoNolFqC1H6xfBYhDfw0nvAUR
x0OOVxDpiRo+EiEfFhotDbCNv6CHGErr+7QH9eudl2qH22omvINk3bzUPfqXLL0tFohFEFekyywP
ifK4F4+mjoF3sD7HbGA0Y+eB3gDJ2so5LewT4K41oURYJXHFYANou39Y7ihzBmmKFjhjzWvxn34D
bUVZhYGBbTkRUHawUnjyrvYDFrk4xRaGqCrUyoQNnpezyBT6iWTCfmN5SfFdLbzSpid38kT2FOtw
O+7BKTEf8zQSUOvwK2d8TiBLZbdtsk4pC5DLvGOubulE9x3ZC2TFzxNOSYoUZHE94ExF39IvjwI9
CZK25lW5GYvbSbvdhPUEm3l3Z2e0JuGtRTeTUxrr37aIEBSVmjMsDbziiMYVSo4TRa4fXbYGGCtv
vLvdU3kVNjjXjgVYCabeIPUnLxAuLNXUkhveOOFwDquR767V6QB91t345qyWCb2MeOGVgdDKTFBW
CqmBnvpAjUIY3NKtyHc+7+Bnpz8QSVby14OSr8OM97zWCScLWrdPKR+5uZE0PRPHKPQY6aXPKFi3
1xUN3fIqmzC6gEwrtECCptu6BGsRQwH/bm1rCvEmBpUIOGiEeh5gKJPpfqoulb2TsR5F+N5oNPT2
3TbsCYima5J3ib0VxCar4uKbdDrOFN5p2xGK8rI9YgsTW0SsuJ5bC38TaP/3KL+u9amtHXFvBTVA
bsgrjYEC0Z6YINc8UVqMAnXSmiYeAtcXZRgZo/A8pQeAaXhNnxbxK+Macrqgjfa7Vf5gS/CIEYs0
J7dQR7Pxjkmn+fl9sXoULsZ8a7bOVaHiodXBpY4II5CC8rMFdC4/fkZ6tDOxmDF3HQu3pfKrm4UY
7pq2DtDeaO7y1ekWFIneAv95qXKpcSho6BF2wXNF20C0hEPXIvuCIWTO9ur56IFAdaHWXXA/lU8Y
ujqZdbkTMrkFhUGMbvdzhUTmla96omplO4IPCcY327KPb4Q4UbQGMIjbeaAKSCvIX15pVxSHjj+w
Afj2WtQjiLCiGccTKwu0EJjspe3MLfBLSLLf4EohjR3tA8J7492N+JYsbSzPLE9JS2KP5OYwswtC
0qP2eFsO7VwdvdBqSicLhWRETBMz8NEW+7JSG44dA8sySA9CGB4G6P28tzrcHTxS6PLGeZ83BQM8
rUt1eMQFfGMDoRbNZRj+svkk+G5OfG4ufL4F9H7hJ0VczqWCLCQc0kPplWQTzWZqswyTERaD8ex9
ojcAS502gQvFnLEas/rNLYzmFoX8ax2Lv7XteedH+DYucIOYZpDSzk5e7Me3Z6VtdnX54Sd1kdS+
UTTBkZOmcbo/YOM5PNsQDcUTp1WhK5hS9fmgDJd8uCz++CoYJtFCI17ENSFwqR6rKIDa1sARBobE
EzEwE97SelCyfKmiO3Ly9Chpv4eeq1n+cZgAyoYwYBS6ys0ANbmAOcT0qjl1AbiOCXJIweIzEYvo
ooG4hFdOHknGoEdA9UZib5YSNZJ44MmaClxk/72B9ys/JZRe4H+fqEwYp6V1eMvIMyL+Ywxv6hE+
eG7cV2vSgUxGBeuWeBCAIg/ok0JAxAAbPiO8QmEGS69xpD31y4DP/FTaPlZVVlm2NN1ZnklZIyNB
RXDRAPIKT82n5TAvG1M7JD1BCWJ7Iyq8iL0LWWHTuczw9rDNLYL9WGe8JgAW65W+6sMjHtwqa+ok
b5wpD30eCfMvXOx1ZPkh+evLQgyE/99eXHEwyad2IepFNfBg7deUSGWE+jYUiA2l0akMCQQC0PpW
Z/b/BBKZPMhgko8BN4RUmMHwlWsqtjpdg3toYPty94P85sV6ghOnpTd0L2EBn4ESD2PeCuXM8JtQ
G8Smn7vdKsOUIzq0VXaejKlIXB9XgQPFf6RjOmZkxcA/i0NUpwZZJALm49d6e9L1eTh67GUFBNdl
6BGTQdZTfteeOZO5ThUrLxcpU1iIXq7Mv5KlCpURbVskxlvFFywlyp2144OuvTvMW2D1PkSd7d5Z
W+/pBEKM3OrmGcHekLOJTQK+1jP6tYbioGat53O2YAXESXEdaw2T5A+XzdL8Fqf3XRcwRu3FMOz7
4iTIELs1JZcfVtpGPr9puWqtm3r6OBxPSAGxFkt8KvbCsKcQnVw+92BWDNiD7VMcXDEeYKhBKRko
/sxk1MfpKAt6hkU2PU3gm6x64vJmYkBekO796uPn0VB98jK/G60NyhZ5bI1hfMUNTK28v4SoUNdJ
EZUK4j8fpUlx9p7zBzHm6MiMiV+2Z0H/Zx6sEgRa3SS6A4qRzOqqUDL/sLuNnW6kudlEwJHjKsY5
26kGZtVGvqw7OMnqx07mUuVx/XXdNUHQCGcWHhkhMpX5GG/9IL0/yMoDY/UK5wn75WCR6CY65rC8
AIJUJZ424ERErm2zqwyC+tS6uIvBXGi01U2AdCPQq/Hbb1dX2jZepiRhSAlNjrT3TUqWgkI+wXPw
sTybPpAI79kU6G1ZHDfjfKSWfGuUSj+jSG4Xjz8T6PtrrfnC+Wx0VxI9/ZEBDn/AJuvGXvBoG1Bb
Fwv9bm7H1vYSOS07/3az7sXhAm9KO6yyQu6HlsniG6Nrc9+MBNtXG0wC4O5nsOQsW8D6uduvHdwR
/n0XBgavHJLpPX4tqANW0ykUuA9XJATCIqpB8u8bKNv0XeWphaRE3Utp2CPJWLrOWSbMhS5PXxx5
l4DmeI+P8Mj4sCdvuSnGPooS9EaHmX1py2WjpIglz4MxzIxKLRUnH5gpBteim9YZurMQ6l1Wr6Pg
RuxXDc5OYH6rPLgRLHuoujBcleuRXK7NMRFqdfS5p5lyee/Z1kDluQoCLTFmv32coRf6NQg7mAD3
8SXrv06+T3rCQ2yNuLidOIOTciIBhvZtyC5gr0bNvpTEr3XAn2GTid8weU2nHvQhhYv+hl1iaWvd
CO5zdlXgjz4CXzNy7LlILmtxTgLp+/OZ/0HwoXNPi8kodWthZ71ENLvpcQYQo9lIp4XCOv9eqHJY
jrKB9mVm+ZlRrZeU4gXzoSNJ/DRU0IMQL+cm7kyXaOzzX5kDO6lN6xNUasDuGn+IMK34uvy7V9qG
VHEs4FCRXepdgHFsUNGM8FZ0oPJZnXicZbkda+JvUXH3+1B7W4nZ71g/rrc9/PoGMoAh8E5bf2Le
OZr1yei3OTx98xS0eV6/SJklfhUiK4EO/9gD9nbMIVXtJyLg9QZHy9WJdMvTWxniMo5XwOz9xbwR
RUl8tfuXbA+mR5ORumgrXtnODqx2h4xZ95pLd7whjBXL86z04SULF03muUS2qjnir8N4EViL2xzE
yPHe29Jp6rRLcXXTyYq2D0LHv/vLzn/UAS2CZljfAwCeNIXgJ9Dstps6Uge+QQOO7GJDA71ESqDw
mg/lY1GkwlAMM1bDNkPQwhkRtih06SKbhRZbDeADZgXsj0ooAIV0WBC9SAD0GjdaA0obX6pDJVVL
7b9WDrDI5b2qDeXlZ7TvWCntQJ+WPF5cReyyiDCS2smWDsuE5N3kUscvsaZAJblcu8FAI1ZnsvsX
czLyvtsJWu/y9nL4IYwdBjsou4720B8hoFW7sy3Rf3nLgWNAXjNbEhaxylDQEh8KUzk86j90vqxA
BR/lO4v9IylRBeeDuxVH79DOmMVY5BQr04GF2OdcjhqurTbKbzB+2zkWSpuiNRCMkSsLid3L/PFR
ES8tR43jMICj1qD7W+nRv0cuGXlXZWGrVnKJyCS8OA+jT5pTWuVy+PYasvToogXqomqmHANqVSJ6
xzK0MDh2m4AVR3XkR5b2t4BQYNydlIS9a/vobNtRTW4/cnp/5dI5aue+yddVT/J5lqeDZH2Zo68n
dlISlY5mJmNl8Rte/U/Uh4bFQfePiZkycTHN5uXGn/Jkv6wY69t0vWNG2uBpL9OKAJd5OfwB7wl3
Xe2x+Xk0eQRarymboYDkOCbsbIFAJU9eGI0KP4/At86qhKZocS5snCw1Ui1a/2JRstc5T42dBwOb
gxSm6loEby8QythMAG/pUvvt16z8PxprJEBbQTZlKoFAOcORxfQsdPqlRHmveabyUjun8c1f64ef
WzFUiy4D8CWU86eWG5Qye0sOTUrJWWyt+4/rjcZA7IPiBxl9apnfeQ27Kx89MWAhqXmCBMz/lmvB
MFKc3GwBFm0K5iqxGW7wuOVnNszlb4g0fA5CLY+QaHoTfzzW4DuC4YYUjBiC2duzREeRuFCn3ZlY
+AbRKRwfZPzzk/sjOUi4nPPa6VLNPptLP0e3Oe8An8FnpSrZATflkv6hf1wACE6+co/xNDsZ9P54
PWKG9oUoVXvSx1aKxxzY1WWfKboPhBhejsDjLa4ggE7rVoJfELr3/qByRwGPucIX2XS4Yo73Th7e
HqoViVW3X9Lf6vgavSvuApNlrbs2TO/ciyjGBvu7LmLXCXQNaei0dXnNKqW9gVW386w97vYkhFUu
+IwtNfO2u4rNLTMAE1WeOvqzR17T26vOLPQ2kvIvEQTjIdZsRJ9Me5PWl6yHyhKTP11nBgxpxVTz
OCdXA3+6kA5E/rQbLabAFIAZWyukbhuY/VOVpCyOwMqgA9Vkbv7TtTOLmkF6RkPd9Bkrmq7Mdtff
2lDqTKDQRlsfO7QIeyT7CbKqsSi1YejGT+9dRd+wqCnpn1v68ZTRU/EILWtfvKqo+Ie/RWwEL0Ua
J1QGjokVR7sROIOs2nmX0q7rx5ZLBfa4ByUsbV+wwMtxvD7Jp8tOj1WxBmAFiIJ4oRz4XYscyf1k
eZOMyBK+en7aqsXhYcTHSvk9/Fbo/A49D4Z4+0sSODZPSWtPrVl7KonwXCfLix5tCNrNLcvFtsp9
MZTsrleVtdOSu4v+vdb5++S/uPDKI2QECE39Ey/Ahrg9gewsoyQ4PX7R93xVFbxbnzGyrctU/X/j
leTJVLIUneKtcsSMu3l4bJN+XwhyCbwqWetq8SNUYNNLYm5hmDb523NJSgMiUNFUCBRr+laBz8es
/Wbldy5LExFjwi0OCUBQjJrxEG2j+uYA7Ndsa4oTLESa6C1Jt+roDu4QcNL/x+t5LrU3gC4hMe71
TgwB8dsdCTCht0ynXJ0ItR8ZFg/SW8ufP+azuXM8RVk2MQqBFTmR91mH8IdeoS9PuroiyLHf5ZrY
ef1M7cUfhSkaW6xSKqMOMNOchnRvp+8cZolJZ4QfRf7zj8OR10Z+1Lk++VFMTZjcIgzqub9vGXPY
+DzDOPva/uhatkmZPWRV8BY0JHBQdxhkpSMzRBi+Lz4gfeUVUYaYVdPl1LjMK85Ns+HW3eH4OWtU
8GB0nH5Hru/FP7XHgIiC8DowaMHUqWc1y+JNUD8ONHmiTCTpOQtPhtmloDFSGFZEb3upbFnUcif9
VhDxsYy7TKnR8VBLVmR/kgnMxD4wSAHklKWT3m4A5NeL5EM/vvRRHT+syV4qBAVw/Yk2Pqs3QhsV
bGqIqEM5Q8WISvRpv5O9FKzBzXXrJaYIDhuBYlbjmzjrDNHVrkTHFeKBXuKSntpkOw8f+Hp9IJXa
mJsGP/6hqEHodrRZt4c7X64Axq5qAeWRcWspjH/uNQ6on4PavVLO3lRZZhmRUmnEPDd3LXRXBMUO
X1HFGBewgyh2a+Hodx1plUPM6JNGpqCzPNElwZr7ZG0kPfWKQqw7MTmTVmsQJtQVnMMLHw/CSgUG
7m4gYU+GZvoJnApoJ0GIG1sB0fazGAlguX3CG3WAeScdX4t7WXUWxS7gKbWaGAEiSrCshIN1umQt
TkpuO1tKFTpdCG39eTNwZQYi7q6jKFIzyA6MAuubQBS0rFG5i+GyLYcc4bEc9k7hAg1CoSqxYPq7
9WqS9+1w2LUiHl6fIzPd1nxFgABTrQU5wGZTbm+eS8rE6jqUzwREJBX20PCZyk/2zMrmUAv2O8ig
Mm2lu5ZzCsRi+IVH3YcbzePnHIz/QDGX1/6q66Tu7e9YklDHnX6jKR2jm83b2IyzaJbtwskMwsD7
4/EQKJLOn+LaVIzX7e6gmZAbblhPOG6o4d4Rwy4iu9mBklMVw309EZ82qHggS62PiOp962IeIJW+
svEsW/LURqo8MsZVMQPLbomdS/W7+/yytuBKILPIr8MBM1yY8ynuYP+c33454dAZRmrf5RuBX6C2
HGI3g3bK5zAkvortfwof8CIwvMCZiAgBNDfJ6m9kLa+yMJA5G+Uq2hMVH1z5egl/fhoSHUS0PDbw
bF6123i/lbOGw9jsNiPE/AYqG53SwCySMyzg/1DUubBxB35WmprFArHKkw3yJVHjK7gzGs9II3Js
ANPocnce3NSW7L3J10h+1C82Iw3xWuD7U5/5AIgZCNJQL870UYXIj/xmH3ktXaz+QX365vl3GD09
TML9yqoJ1TkY5MliEEG+OzFw+VLdFUIs3IxPpKkS4K7/FUWEZFaKy9OpCfjV/J62YFUIAFC4FZgy
Cw+gWqsWAWtIbm7s0qs21cVp0B1ZBtCTeSr5S79T21yP7yxahm4FjXdt4BjBMRLna8RmqCWAFSas
oZVf7fuQBsSWpZp/OhOOrdBt8J36UuxRBA4XRlzhH+Z6tQhVQufJFphMDeB46qC2oL6igq7DFBiK
f6VINk7WEtSNYbJz20s7q6Y04T0SdU/TF7qxYADGRTkg7zs3oso8eWS16lK/s4cBAQifOkjbl0vb
DR7zysYGcy0JEqPgSdWpS3ozw9jgusE/mjfTgWTQDOL+DTzL3Ou8W8z5bQDoQFs4NF1A3iVwo0P1
rybV9+ayB2mD9saB5ELTAw6Q6V10Q+WrgWocZPgTjb6QvoanBkr2RDzzW9+4VKOMNAf9xHxWwadU
N6KiHeCFPi0n1UxaQKIajl4GXb1i63Xv6/P0GG3Aksh7x1Er3Ynq9gOx1UDTKKWGVxOrRCrP9WBm
Q20QgrCPFVV+492FSSzMHQcsq8OdUXXcRNPghcmdmedif/Vsc/1sr8uKp5v/OZm2fuyBg3/8jd/q
BsvWOD2+5mFoy9CBeuzdKpRS0E2f4IkxKGgXeuJhKe29sgghre5nD0rD62KCUmxOT/QxQ1TXoA2W
yBL/MENseyLcSLyH0mG9wC7yFHfJaNFY2c3vwDu+GS1ml0yw3MBFXz16uzmlNlovMcnFsQxJoL/N
1nl7W979C4NHbcBvsopfYIFGl5npPv7NsS1t86BxYfpVKQB8MNgBfCWA0ft0o4HbAVPZka9/Cmyo
MJWBPL69MkKB1kKO726cbHvKdOsFrxCcRol52JRkfhJe03g5YG0IivsUrmYrYt12+Z3TeU7De/xO
LYuykSfGJz0VSplS1OcXG+fflPxQazzAucUWH2gMscenm+WQlw2m5Vt8ntcGnSCoic18p2tAfwJs
l2sTfqXFqrQg7pSIDRXg3X3vSD6o9+6ds1VWzXx9J4cJgfBnnScd9sYIO8+er/ZP76F0eommN07/
p4rlAxoGixeF1EHtB/gIrZmZzV+pe8hdJuX/aJPyDtGjzqK9zID8K1cI2c0lYZAvSbgjatcLr8oM
8QYrHt0FjSO3Xh/jAU58SKJEQzUV6yxFrjR/PfjDIonPA0slKEg8Vz8X3oD5hvlOKn75ckUmzVFR
bRKwSUAl7fiawct4TzfRnL00KwGFH5PyYcgU3eV1j/AyB3uyiXS5NeqYKjySbQkNzSkJnnYCM+j2
m1YhETyPUq0zX641i0aWhPmeYlq7Mlt9PbTmdDgMOZ8YtCbl/KBvkJ0U+qlguoxMIk7IY+MR++JD
WFQQNpAriu3lDfyBvr5MZHuqn5dUAqamGCPJZeLRXhG1d3oBQLxRSvbGd04XVGYdJ2kWrQYjF8il
2Wi+TkUQndYpe4Lg5XwfXi6OIP7T+XyKyb9sL0lUx8pfBX/jzr+YTDxQVKX+Oh79k5EiH84ZlRm7
AIECX7IfAR0Sxw8w26At7JvNWY0b+L9XU4Iu7QhZotkxNjlPCBOYmc2gdro34Jmk+BWRhI1SFhVA
lKMHAZBEK23d2oIPpIn3JlptWYouNbiOHwWfMoU8NAc4+6KVy235Q7rUZk9T8fJTvmsMCTMPoCgB
iCPh3GdY9sYFZtunCIBt/8KidPeOof9clvV4dEAC+FUqglv1wC7QroknItccw5pb/7AVgWS4njdU
XQ6F4Oebb47c1pPVkarf7DfLXO4/NnH/8vPQAcO/cqDSQ0TztFAufx09f26vdPpRCxGp355jnd3M
H9ncaE1b4J6CJE+4t+M0zGuQQjbk4AkPBy3WERqLufllbbCJi9TXX8hAYBr9vQobGei12F+gPCO9
zw8OPE3+eYzaPcRH/X8/m/By/Uj2tzYhVo64MijZQp/hXEK1owgCCgEWmKzyeGbxqB+s2zttidad
cOJQuqGOevM2Y914LQNx3RWZbnEKaudpIu61QhlkphKN0rnNqRdYJ47ER+ig5NY5DeFLToZLa4TK
MdMj4dCo0EKg0G0/2mpnnYtI2EW3eqPTpwm/XG+88FUD+G2VeNUsul2u18cGNjZTlSc7FKfND6nT
uoL3dwkKgpxPoJU6drJTxp4NTpvkaVzNw3DaoRfnFOT3/c1DL2s9j/cgtlv6icLlQ7fDUty69dhQ
unchoqn8dB3ZsdPj7FI5qbqDNX7LwNiP+jce7z69Ynj/yyFDAuWjkLrfaE7pmKNMfT15zvqV3B1d
5ssIO7GUWgVqWWc1Y2XlY0c0+cJLQexZoTy4UwsEjbtBqE6wgHrdF19Cr/a7Ibxz/AsZBXQHyWMX
CrS5OPQM7yWqTrlcRYCgSBfygTo5/RF66qjbAaVro2k7+V4JkbiEc39NuIkAmbqYyMaRqjhtcW5i
8EP0oGHDTfg6Z2nng3Vij4GI6Gb/wdmNPL+zIfXcmVFofqOCOMb8cVkQluj2aUw8YVBTKRPrKGVM
b6f37FTZ+/OWRB97C0HpsC1IUsduAf9S3og+9LkW+gsERNGBeecBhgFwT2QRLtkbs0HxUb6oaU9u
jDpiHK6op3f36JQ9+QktAtx2u6+bqsojC6YKF7SHvJ8j+34WVeabsVZFNHYFxdPrfDdyLIyHUsKU
HA9K1EdUiF1cnWTX64lXA/sFpzZNxuYus0HwcfejJZ8PXKa6nh7CZq2sNBSvpJf7G1iy2JMGSA5d
f0f3ph9ZcoSXRubdbiaFS3CMqN36huSsUYSnAaLrRRHN73V1SfoLsGSwCc7ywJML5Ut5B11HLS9N
z3pazj0iH6J+C/c4rXJnf+MOQQg0fFIVcGDip4NO0Fp+J1efud62MFeh8yfalZ5fU9P6VOb0Qvem
OXDy86/uU4CiYeVczvs9zF5c4X2urobM4nXgMNeNaVxcyIz8nSvhdSZWKXPJDgSzIXsDaAag5Bja
F/P7yayK2Meqz4nfPAUExh7b8A88MQr75atDFDih16HOknwKSeUix8QW0HgOj0plB+mQOmU56tQ3
08jleNkAmxFQo9/YLZVjYqCUkXH3X3y6U+7y8Ds/k2ZjRL4J2mIZnV9V5thju6bzYkIhtxSOgS2E
swOzL32shVyiG3/omxpfIViGppoPKiCODI49cG8LSP4o9qGBpf0wT+lZVUdnL+abcD0GJaiN2DZW
rH6ldXBO+HXZA7FPpRWbh1Bl+50w9uQ5QODgHvAnp+qwWVy84Lj5U6kz5xCMbYXwRylo6ve9jVg6
xlzwS46/qKS7yXTFBKsSg+06g5D/RA53RctTFVeObOQ6Qzs2WJBQb0Nl+xbKYL9EvniSj6Nx1Wd1
8HQpNbNwNxP5JORydm9uoWnNDxnffkSPXfbq/3bE0paC5E6LfaPONVJA8S9TTv+HFjS1q8Wgfioj
Lbi7PatFXNZyby4QZBQy27skIApVAgSOgYu11wwLx0kuRddE7A0MiN2HsM4+229LF5cQbzoecikY
jKzvIF3LT/Aoj/5ZnE2TtbXBUHlRqVhu8LxRmK442AM4h3ETByfb2jJcepFbt+Oqr5zLy/Tc+rQt
5NKL7T9qnv1We8O+kwrIGR0z/XRp2TUvjCZ6kyNCZqEjqZ2E722DRYv9ipVHFTNvlqhXfF/kZCbI
z0xyHMmw/p6fgT3IOzCA5uIMUOZmvtC8seAGI0BNbdd8qtCxbplT46fTBc8UZUqHKu7hsVllSiT2
sAsApBouRhtnwTeaibHXwGAQMwaNyIiaEp00ycPJIroo21B4Z/UVe8MbeK7MssXh2eMTqlR/Ttca
ixEyEv6ZNU0WjnK/m6h12Z+e9XHCXZhGDWu5xwJJ7lhHE4qcaMFuBfK4QpcJI8Z3+02/YdbynP3N
czteMMnQ8BZiQNWECuj2nMFEKRmzg8d2PrNuV6J9byIBsNvFyOR0weZ9XAtTtxK415ATjikQjImj
FemzNoDnCqCnWKooogJzCAIQI7Asr4Fkq68cBVblT2a6HzEN4dzDDbGlqxiDa/nF7Zl9Cm8ftbtE
gXrXK2xo9n223yydD3zocXXdIuc9aON9wRNTcy+bJ5eDGVDJzI/3cczZOQNGO0WbWLF49f4fc0te
veEPFCJPIAC5y/r+RjzAYbujMvalD0wvCOZrLKLa7HB7AHYx8tIyqeuXQBZiu1AboFvP9AD3YfHA
lisD9nZlYIVSmMtGoH1MiXs318uWD6q5/34i9Q49Hh09Fp/8nrrbvrev1LhanlA/M4PdJcgho9J+
ILLlEvoejbQeAH/M1B6a1W5vO2Bam8Wey3iYEF/SwFGmestCyAHlWMXeFz04QUg7wnMCp3gnW2jS
1ewtIGP/lwNcPvCIDMK4iMUm+/mQVdKEFpbNRTVP6zMl0z8fnQdsR92g9yVxFOfXJnub1Mc3t0jz
s2fPDE77gefMedc3oFC2/tQ+tqUC/hU3ihKIyoAUfU8dprL3Z2DY4CYHzSpar3QkUH7JwRk0LYxO
lBq5ray2gZO23VF/LCDMxv68YVQpkxrB6+pK8gK8TREloUo0Epra5cqiXooEo+nwR7H7vpGR6xSb
tW3erXTI3vNY8cFz7+D9f2Qq79MUCJsPAY3TyBkijVJu0SW7lV6B0wbgzJoBKMzjUGfwEAn7ol1p
2TSuPliwHoiz3ZPp8j8yFJHtj0rJLKh/PIeu3dSf0ZzWBfNYDJZgLNq7IkeARm7ekrRCF+5zwZ+w
1EOwRgGYx6O/gr/lXkf5kHek2q0IJExeuKaiW8PFh8LibcuceERtjLDEfGnoa6Qq04POjJRi+95a
eI4w3e4t/u9A2Pzce7qxx7BoNGF7DAJWAepLHoUAYw8LBfmTtn7CsU4ssU/gh4NE+eu91tvVJQGZ
2F6r9/xg0iMdBAkBnfINdf01JQipD2hC8i+2voRxAO5WE9JLNGrzCyZNIofQg1JOEoib+Mtb6kTC
/IfSBBRATFt7Dt3vlENr0LWbtXu7xP6c/LUfClzo/RFBmndxgYQG1+theqAZy04INZlbyUAerNP9
DOSgpyV+SXpMo5oHu73N9yQEsuiuag/3g36o43CROiUJcwuJRFiZQZEtMo2il/qiT61g0QiyJJxH
wR8zb6mILD5AXhUlyFTqB4KUNft0p4KYB1QqFx+rnWohm6sfqPMdadHbDklPoU1mWcd0bsGlXHo6
n4Z3PL38MSObHzdWqTbAJ+oKDO07U10i7OueGNcQ0WIB2iQUh9gfJtpn2wS3RP01bZNdXqHVjcB9
1t6k8Opx/FvOudAgztATmirC0s51YOWzhtRYkRqVGpNFhTTbAdBgL7XfPpmp4HbYlM6PlwwM1aHp
bgx70IxE+DTfnYW4ZeWPqmtG19QIIdmSNRHbvhupX14fl0svK5M6hViBy1r50SJifMKhHZHswa+q
4q24LJ7NJTPDI551sm85CILv4Itp+7q8u4GxWE8aGq4WM0oBp1KohBrG/yBl/nWhZVtRrITbAykH
rmFOpgGYIPfocEP7PfXcvncQZ6x6UA0UxIOwbSRKXjIL5OkGHlVBF76xbYN11/O3DXl+rIKSPoDv
N2UgnCy8ABTanLoaeS6oAr2kdquxj9pmowewtCbHJQcaJJIeYeD8TjrpQnWxpf/KOjoS1ikHrp3j
zfMYtm+EeiQwVLdZs3Zy/onVKs1oiBWlzoUnehm1H2iCcw0louNHPthaLW1exarDDsyIk1/xwRcI
WutM/OuLmAaEF8YqROz5A8fSnCGKbesrpyxRBlvjb2uYABwZDmik64yh3qmi3NIVswIbMejg2/H/
VNkpDJXhTSKkB5qdqnYaQ1Rx1Q649hl2BVpcEN8ERo/c+kb2ZvVEo79U10zfRMhJQYuhiYHH1u4q
JNVS4mV47lxPyQmIWusti0kPNW4fJZCWFqHq2wAmtHBMmUJCcsRsN37Q1iZKf6YYEOkffPK8b6xG
GnmEHGyBFgoANiAA3nm50SpfklF72FI+qzpYgJHgIh2dzS2BJqtqfcG9l8zhVqIaKrYarLJgya1H
3uFkoDQy0uQWYlowhieJl0wqdl5lBOLt7gJI+5FhhBJExDF7HSNQ6A8Vb0e6F7wg32ecMdlMLAx/
s9zdjgKhR87XWYAKAnsdwaqa/lMAAVU9DN4j1vDbo4HtgyzA/RL3qfOcBFSFtISK3PZBBb9TWcaX
MdF6zCeV0+v2JDOH/lAS077cSyuUwW0xPiYLt11oLNWHmoPl3UyWWDIms895uZmCIQ8JWOYXTVZM
DPO56RI/UcNdJ+3GUEidXxui/V9/cTSkaHXpwZhBiC/Sysv8Yq7HKu9LhlP3VHQW8FUo3mCc/bRp
R02P/Gfh+VDlZSmDPRKm0hDcNVQww88js0N48GBTn7nDyUgwplrpRo5NDH6KEq5FgDjnFTL+ByRJ
FBkxcNZ7c5DAthkkn6OvyHQ4RO4W3HG+exUT+E7BoRV2oqY3Zlh/0orCmMuarEhl6JuABwPQkdgi
w84fXigXZRYnaMXaTPpwqsMaJ5s/uanPojPldwzKQ0txdB2d28IYCB3C4k3/302UJ9tReRWNna5M
O96lmW8eqsz2oaIvy8Xujy5x87/AOaW/OFx2lPyg49IikXzD6Wgt4VlH7IngRrdUIMQUi44tkATc
dkLmJLz1cf2fVHLYuKaWrK/YvLMW9DsUo7ZJGZxIotuNGT2d+5mYqcfkm4KQ0c1hphm1HVwrP9du
/DzrZ4rQTW7YBC5e2mfl8UQ+Mp/jeuHVjIIGikVEeV7ZKO74xC7X94V1UNy9300WXVMqw8kQoJhM
Tq/6xlps9CXjQ/RLz7RIpwtn70ZeuYamjum/rm1ZvZx/zoVsb73srfrSdU/SWWCKBADF1GX3dxRJ
4JkGvPrY5SiZsVGQoG6Gb1qKttOyDyyBzGJ17vjPOeYVsatW7WfE9L4FMpe5cKQBT8NPCMaKzDJ5
9FVoeZdqVnZUSQ1SeTAsXyyJVn///afbIM7UcaEDwTf9IIXAzwqTdEqI3NVMLRxhtaIE1MYhNVtQ
+IbYtpjKruUOwneSx6Z8ZVTnI3MwMc26jFh0gWhRh97li5VPe+Wt1tU2bTaRdebWKRtMTBYUWS1P
BLwmC1pwG1nofFWMcWSQjKbqsafD3czsPZt36Z7JI/gm8Xg6S2DZzD0AIkAg8Bc/mgDWi/kNcDX5
+KxngzxhBkAj/wB/fOAcr02srME8SL/rioCiXTWrVkXuc7aIb6ko5WDh4uqG6JfdeaTtSmXjhzZU
ugfnH0cIgrHtPIWqzkj+8yg8yrZFe8BUsTdEIaZgk56L0F2yW+iYI0nebeDdIuYVGdb3bXWOWXGh
nXxNNDdlQQ4Rt+mCjym9ILQqmES/ci5wkfQcGwObdxvtoG6gvSAYFbZj/kN7xc1npIs8YZeyEGTc
zGYNyi4dmbvjnqPRYUVx6XQBL4QZGZgFUjp1Kilmj1beAKWDaRia7FH8gLUl/X+oCCT6BM09kRxE
6sZvgFqDpnuFdEekZ0ALAvVR/W9KpPpb/mDm26ExErJHn0N00E7LiZoXDAR8504SCoxnUPQ84OE1
akFGxuimLUQOJ58VFEMuqR+sJWB6l2ee2k5FkmhdglGuyvv6K8hxHTDHepJHXcutzDkaa8JAUMZv
woLt/1Vk6701bF8a0oz1ir9r9tNHOIzMDTnV/34twM6zFCXNC2kjARt8A0pJ2ckxIi/8Z0YVVVvg
PM5s4/NdhGCG6GriL5UlnyLR7i8JYg39+22V+T9fkXnRXMEJRsOcd724DIm3ducdDIYqtNJVv/mR
ykn9F5tNZ68HbDURhiog0x3+NVQIA/r2UsWb0rXExvLeeaVnIKCiT697ajoIve5B+LEMyAdnPESP
wbihzREejVqkzfxpdYZURD14EfKkORFXNTI51RkOtgHqIjs78h4lzYvp2nLLzQiR1CQxTLtJFHwU
QzhVILXqHibFcw9G24knTVBS8nIWyzurHkBFLJDazv/OP63YjnjN0VeSy0LYGHC80pwK7hNCECMS
EHyvvPY/B+Bp8TQzT7yqxV/8aFRqQ64OUk5bjlxpJrZ/wteTkmPmf55MpAj0ux0NLHqi21lGwkLs
L39QBqai5SswwewnU5P5Ecw+GI+VzWgjdSZqRs0OzJiZlkTpxVXnSN97LxGmc2BYd92CVHXxc4sj
lw4J0NCRTFjbjw0ZuUYX+Ge3cVTpMq2AjGM9Ae81qyJULkQs6eyV9D7PhA192pyzNeHgWkgxvHgc
W3BUFCt+/PIrvVfMuO8iEiD6UPm0h4JfkXO8S/7XQz5MO7lTpGlWByvavQ0TCEiUUno9IBbSii14
DuYWd49ZhUO7eoXDpnHvrKmA016A3sE3bw8dt8HZburlKzuFtFt4XmYMcXe3M/42NHAmpv5VI7pC
3ClvtjKcNESkeBOt/oIsXa9gVwJyyVjhKIZ56j/LHH+mVjZg9rOOw0H4l3/mLblYIUUvvX0UiV6i
qFE+h+v6DibJNK2gMEDjpXJQbgnEp+PaZZpbCQHM3PINsppYrNOiq93QM/6J+FoFnn8dhpR/s5/5
QYmNJ4AcK2tLgqX8MkwwlCLoTX0SMW1BfApSdTZmMK6aTgyIZDIjcN7qqo9N8Er2V/3d2be/NN1p
4r8TaUQ+GP0WW10VokpDJ8kfEiwgqeKBRVkejjUbZwgxHH19WhV7tCApkZTfky/KwCrv892YAOK2
d+Sv5dqSkclRaRgnbxl2GuJ8cFoRMIM45wxIdMyasd0g2m2IN7AIfn+jB7NKAyHOGAEjeuJXd81U
JL+0Xf6FwPdpqrWPA6RwKjE6EdrJ6ydf1S7V6MNezIt4WN7uU5uSrldfnS6kU5IxO2gj0UDdfuZ0
rxqnZvlvbdGZiAPqU2Z3P9eOAbOHpfyLmzTazgvStEq8V8eaCBl/bzObMoZSjuwsgoAhPDGt6kSA
9gdMVJ1C2N0vhZdXaDuty5ZH03VDSm7ZhFnJculixd7ToQAdc21jQdyI31W/sRtFtsLMe7L1Ia3Y
XYvXsQ1sHpd+Kc0QBvc9a004G9Ek/e9b3G/Gee6X4dwzaAXPr44L3S+p7x6cTRmEyA8d72eA0k2b
0sryNxynx+33QO3ySTppKEdR0dKeMU+OYmi3Y9iLQ09dplr5euef1S54KAjxFBPT42YTvjE/BAH+
1uswHCxLpNX2alSW8Qwv65GQJEhO1oZiQ8Ut6mHMHstf5/aziHfGwhjmTHJTBx7w2TN7PhqNYq10
f5CWbQX2UqxUH5XftKAEFYZcnm3iG/v4l4B/KniWpHgE4Z91J1pEqcX/JsMyN5jS/woA0dvyY161
3hDttQsgRgy0td3c9C2xWHUnl45Dnobh/ANkVoDKq+/0dk2uVtjO3hMoU3gzX9x4ffGvK1w7pvOk
51gJdphe2lb15ZhPmetYfNYFlgGqeP7JnD3SaHG3SLzNoJDnYWIHSmmqICMMObDDts79pVdy6DoZ
KTrKmAztNLsT6qgYAzvSOkF3xulQJktjkDvJKLxXYP+tMQOFf9QswpnhZK50bDTWgqRcuIopDK81
mMqXyLMPJo/YOmScBcDAmAecnYZMW02QzQNcuopedeQ98/goSDjYvl4yWxHaeYT70MSrxhlt62K8
UrrJUXGaHdCRpkilSuFS5jWb5kBSzBghwsshMfXMlQHlGSkq0OyVciwPpBRMds5erRO+5IpLM/qI
OLfftKCccgIAGELsBYdj4IBnBiKB8qpul/3RDSoOwqasSDGGgnwbXUAsjLiYV+CaA7GVIXJiuIyj
Vx3D0zlc+Ku9ttSBiF5i8bLeKFaS4KSRuz787+e4vlCyHaEsdEYG0AWIo869Gg9it6o1n4ilt2he
x7TeESt9OlvHFXCfl/T7B71afzDJ+CEhWl1AxIaRrpWdX1D1kMzjz58rbAVPg3IHyXvGpg38yVFA
KIJmS0S7xhgJU5FJA7SxnPecsWJKbaXrkniOOkLS1HOblQ2B5TleaYz0ih0NQIesD31YQYH+K46F
mp/x4uiTdwKG0YXKwyeBj4ulIBMqq0xxjzV45VWAK2Uj4y2brLsr0soVSnDVy3/1OwNuEJC/gimR
LrxCw6y8U7MLpArukXAzALy3n1bcdSynfUVeLgrqP3Sv1ikNLQ/3q50VYTnGIaYbdrbpmhO6unZM
Xz43nkb1AhELOHtRCzPuZB+E7d1uFvdUEm0jhrRQfoui5F+Hm3SeFGWeqhuZyYgI7yRJ8bJKrN3h
jJh3mC6BY47n/GqN3GlAh3J7qgcnO3SFZZ8QhFCfhTo9aTQWmfFdOYBR0GO4yEOpfLIneQhVldrG
14Qnmuexj4MDAt3GLGNuo/ZP7rr7M0F+FzLWZZVga9MEUm4T+0Q3LPi04RkQMr1trQ+Th/v+XQHL
f6nV16INdSN9o6kHBpjbTpwrL7Nsl7QVtJFRic+78LQlakWzOUO4DutYwqX1m6A9gakzmOsAldvY
z8zQefnYbG/4Lh6Pc/qO/EdsTcRxQC9QzNjVp8vxjNBF3EZsfvkCWOMoIMJoO3YzwAjzHYU8FBvU
j0kXr/65cyP1EjUtda87xZ4X7lTrhAWbOIiTdPun6BlU+DiBS0YlVZvCgmjOjXniKnR2N1gNSQLe
/QR52AYWLyX9iM9VSKtBGSemOH6iEllfpYHbMTq+n2T3+IWwRZzEzLAPC6TS59cCDj93pncxucDz
f20uI/7siwOtnh8rOcvq6O2h8PpxpsV47Mg2vXDE0PgOjy3wJ3ToejszGutJmfMsVTc0b5cor2Px
JmPgUJW4S8J67mtgsXB6guU9K8zdd4E83E6bKaYxoRgewgJCBhn6z17EMs34O8W+f8NCblwdlurk
AHP8gpG/TpCBM4b+Ned4Lj+kwN9oFv6uKTrB7T0sFK0VZhxTHSUpqKyKAye2NfhTycMVImgmbIr3
UObst0hfwoNRMxR+af1nt/8xRNgVNHa6f5siGmbyXgLyiO86vvvKyXHAi61z81+yCwxamy4joj+9
pa2ZezV2dfbOQqMUhN5fRVmIQnJAiLBQBB6JUwHJT8bIqlj3ucHxQLx5knTWJ0ynfLWyMd7E+rgW
K+0ypo1UhkObaBDwdgsd0r3MaIxXh88AzMwayGjw+nym6OrXdIxTZJ1+TTg8i8fFYtYrbzZYZcIt
bscdP8QDCTQxq8BDKkxi1kRJ0/KchOO8fcNuV42L7qw7eZwwwxdnWGWp3najmDwcFy7bm1OtAEd6
xlZIBJU2sQivEejOnBev7WqZYU/nITpG7QTUyDRHkj2CH+GgCKS4SsX5oPMQe2x/kkR8CZX/Eg3s
tkGVPorRcSaYwNNbbQjjGWj5JzG3hj9xcfyozCA2OzJAPVnclB2YzaJAYlQtP4TexVQoMSTP4Ybs
SxpI1DvXBk4yYu3Qhs7Ltuxe3n+TSXiJgnweWuOSjsgWdAUonhDFj4q+BJV/Apj/d3sylPaMobVq
fOBKcvI2g5X2bY65eBQPJS/BNASogDJ8liteR9tIT82UlIvwjdOtjw7sn2nToBTVb1rFWvQjyx65
7Ir3XE/NS9CXiccRqJHxLNZ5bQtZFNIHx970yj8CsD6mXYlUYW0RHwCDtkvccMqs+ay2ar23mEgK
tT8Gaywr7xIgvjPBT0BhiR8qWTTf00VE8pLqDbH5TcKMjd6Hb6RbEmySu17SRD4r7C5jgd8+YCZ+
g7SnaK08DjxYWLnHcJhKjfSWNjhmqxa9e69ETV3ag2ALw9VdZPlf1/RVnabAWTjkxlDG801EZo4W
4huJ72N0wd8kYzEmZNukBXnGLyKUFpHzYFlp3JFH2AwSttho/ok+i02azIRKKtoDtVN3IeLo54pW
3eAmhT0S4cEtaP6ZzRcGj42skhtAproFVoMKY0I4abADEOeNpPnSN51cPlb+LIVTzdkf72rSYJp8
w+fYfSg2u1htC6mejiLjAw8PhAJBBZdV9q66AroKFaGC28vzfV6RBo2xmu+DOAQwHNjwj2gr1oqp
3DfcZDnTDM0ce1YEZtP5KV3KAgCHacv+7VruXkp9vdibbUktOOHkJTo7x+tmJ4GXGmRhnGeacRo6
+zJkpoREJXKrL6xcOJq77VfzooJ0iNOb1g3Ea/gXaypmhZh0QSDrQDbARYj+a6XNrae21E4UWKlb
V2Y8x1mZQtVTM11LRLPkivReKlrE8UbhQoeHNYPXOJal70s4oZh5ToVf3EaSlYrTaGXhWDByJAzi
JHKLMrpmIW+HsEm0oI7zpyDLGWmMIPNuB2f1p16nBo4iqb1DDxLRCSykXIt4ZCWptiGclsCKbxV2
cchRBXoFKQP8lkMeY1p7gn0OFRIgVUV7OO1XzwUcrwqvbDlZ4e9vCh2q1ATynMgfe3mxqhu3vIE7
v8STEHP3VttBvClVTWtOybUGtM9bduLvytso7BPcHKdnAJPO11IyBbPdggCY8S2b2LzM9h9ley7T
2ami+fSfejJvqNGZES5nkRn8OiuQAc3VN6FHh+V7tgd3fWKpHpEcskha90YcgHnSpnA2tIjNcTAd
d6DIYyvsCw3bGA5cCuURi+0S7pa9GsEBxYQUDCCVtX6R8DPujUhBAXJfLCRKQ3SHaQ/oRMooigJK
/BVILEq4ahWaVeEBmQqgaBAxSyg6U69HqVBjjfWap7FVQZ5XYvr5ewTz1Zme9eKb3MiDAydQ+YNM
xfc7ppHWblduudQoMk8MhoJkPa8BtU4jO6APGXq+xEY2BMX3ctLrkWkdjWqHa95cdJ7bc8fRVr6O
MqPHDVieRxEKFCq4XgSRdu/F2FcyylXbr47i8W0F8/Ot4ahUBN1WIxAvzjUHl6CZI23eWXnMmMuc
g8Af7wNgpMgMu3j94An/tDDJprX7Hb8u+0FLpSwE5T85VAgxhE4jQmuk5CDL/DSodXQBBBprFofJ
YOokLQzFUvglOIEcp7FEv1BeJOZNp7sZrLgBBT+udxnCWEcmnG5Zia5zHEl09JPTzihONF+Opa+r
f+NE2swovtB8P4dpnavWGvQiS5a4Qrv/hbeJE0uRbrEEE6w3F3XkgJHwNdTu/1o7Antqmwp5xIAG
8CWFIVFi7kqhWuo2m6eAVYB7c+b8fWUaCryOakgM/RGYAvHI4AFb/Ghfqox1TluZGD/jdA1VzFOf
7k9xpjkiHNJQPxZhm8t5BwHfFBPbzhCMg/wo6JbaSj7heuJb4zzDHODxFUJWTAsC0my5LVSn+0GA
SpVnaWYaGYVwwUohXZk4I6p+pFjSS3VBjEA14vVDd5+5C/6TVK5khqf/xdKmY4zvlo2UqvIRmLxO
FOLt9MkvcjTPxiu7tqqwtnG5r43gniBULZDuHYCQbwmG8+n3NDOrYpGBroe5JQPfSMHd/ROMUBaP
ZNauAreKU3ZPLMiCm1IBmRPdwe1n0rEwBlGEcMwFelhgYqPmAa4j2T+VHmxse4wXhXa2zLdA1NRa
/GDqec++76BodT9UH/xwF9HyDimwEiIKrb+r3wYMy7Z+rFHtFIMwriSJChvjRARn+6Zu9OAvkUdB
RSlIvMMS9hykMFBSPrlWOYe7i5jDN63Rd45fr5kJAWJH+3gjE+IFoqWwEj6/j77gWiA+xnfuXfMr
ESmV6VrlTXlF2bCgQvX862Cxaql6U6aCSjkgGYR2scbOikePO5WDWYhUOYRyBuOoGmIrFf+HzyLL
9cUdNjfOBlq2jiykqCP8iCrkdv3fWDvdqITqyAkqTz63DBV1fkMmZVyJsV0gpzgJieQu5VEDPM81
yD3naksZPYX2UantQlheK3NFP9Ruva4qzY2oMMJ/v4HZF/VmZsTPUPsOyx3TaaUM8AKp/Y60HCGK
hxLw/X70qDVpdvg673TCtVl3+Q/OGbsGYdRfdOTxIh4Tk9kbzx+9sR/up1Gav5MQcEDASFzf8pBv
UhjHqVhX1H2Q+QOIRe6l4z3Hladv3eyLB88FTq3fXqT+XN5BzIxUKkB1cBFl7StS8FOAxMNHEeXJ
SeZTIp3b5p/UfWb+3fhFIY83aA37Jz0ayIr+OSxhZ7WAonu4ST0lO0Fl4110UEOAFNMMIyuqFAOZ
kYsnz33VMqiSixNMnM1eMpcaArq1/b9UKqJKt9sPILFrUOH3I7cZPcgrQmMd5EnlfD1TWLLoIabN
waLz0upxET3A3Ru1EqrjQYRrLrXwn7eUO/VLIFlkpVdZI8eo80aPE9+apva5GCbHMIkaSqXBdC72
QHQD/ckwgixgkPS8Gv7qhw/w49WJFMIvPauvhBYPr6cm3a7J29zgl327DLPromqEWHHsrDTpwcsa
gKWZ2kjiE0jD3mAcWstwWw3OTsV9AuhSTu+6VaGQQ8Ci9sSumjw71QfoufBqttJTnncBRYq4aJSs
jEtzjBJjPqpTA3ps036iLFXSt2e8mrjEkR0Xo336O5+Rr4PieJjq9UPCMLrQ7JPNKl+oROeN6Kdr
Ma9KWZzOX7N5AzURxOPSYnm4JVdCQc+45T+KWbK0U5Jp9pHScBo/pkk6aRA3NrdGsDmdtZRs0nzk
1llzq6ft6xbT9PA3q2vel110uIDlbW9kxrcWGDpGzv2TeUtbgSPmHp5aW92Q/ylxoXo9gxlcgSYQ
nrWEUm+ciAhCErP0EzSqXG9c1pctSbaRr/IowdIvdL/IYx+Xpxt6AFAvXfxR3zGzWOP+949L0GCr
RuaXFG6p59tmT4N7ZoYJ6PAgsDbnXKV8+uJjpPLuq+GZ1g/m/qBVDMN2PkbEdBFIteqwxs8YlS3K
q3Fm6ZU7po89BPq/QfO+8Q9utwD0z4NnpFbPVr3ZLi/I6B0EiV8NbNpWDYpYE9uyOmQJCqzb3zuG
Z4CfMijobeJEYrp7Y7p1G3s/oz9wuD9ZncwnLLmJDlfRrs+o0Y7tjiKdFnhUTEgjgIL4vSHQhvwt
EOnovnoW8FQ4pAplYOi3dBdJSxkNlW7yAgPiUUJj/UgSku2rTA7CC4iUGE/etCautr2Vvol5nc5W
HC+WBbi2YustXRtMMUzD31+t3CKNacxC94djqIYGLheUC0huO3gcII116GopVnrSCzNXcmB9bkYo
xLLzgHXRTiHrXHv1VJRZEMQhBQ+vd4hKzjcSyaRX/EtbWK+GiVEB6SqVv1A7iZdwbRI9RgGWuXip
sekntv3Pm2+AWL0HnNPDvsKeRFk9+LLakUYiIfAoKkbUxLB6CzPqevd2sgwxcwqgWJwaS2Z6nTrS
zmHdL4ywoIXdWbungVBPvqDUVfkjjk77n1WLTMK2OeixEb72/FhRias2Jb4nJu0x/8VqvoJQTVCu
zdU/E61Q/zu1eONCxR4l5MzjUOkoNiRLw2eJnRbW2USIsMlEv8ifKab1fOA3JK0NLnB+rsDoB7no
fQ3UZ4EdMWMv0zSdN7xD0SoqDDF3nxvLR9LCy85VVxyTUOcbFdmK+EOwZtzwu8b3oK6i10bv9SoU
+C3HFMspqcFYT7LQl/5LNCJZIbY9GekCKgpEgjcc0ga2c/L5G2AKjlMPVIiBjJ4WQyL3JNkf3Mq5
PL2lcsg0mni8R3epN+iHstx0HmNuvY+oGIuHxZsKBN5aVaSB1w1bzfCzUsxp1B6AHePjSyT25wxV
c4SMYbhpRMlvm0rtf4yDGVKix8QgnXSUPKPLTCaEN4vnljWuU3khPsB3uPkUMfnl+O1hc/fDc070
sAjqqFH/gWOjEqAKNxAQ/+XWjiKWMySZVullLV+kfrtrwaFqerR9EBat2gs9Vgnhen2HLWYjyQVx
p25CRvVJ0FfRZDc8WRTHDkD2S10JaiMbcpVZAw64dIskboDujdQTjGm/stcfAJ2LhnYtGwV1ajPF
BtDwdHEVuNP0xGR9/ksK8jsbDTYheeS0vVYMh91FYjHLrssjrKbNZDfjOWBm1x9Bz3MnPOnAmqkj
Bi7a9kwVJnxZReS0BaWT4cJ6Yfy+ToLsjG23p3K9Ygg+Db70m3+4j/Gyi/9gGD/0x5orcsR69W1D
lotioFFfRHRrOCOIP9hBH9tSKASp/vle029xVVzYcGpA0yfve6scw5gu4ewL9hMNezoVMyMURQAs
DZHIWmRFUOeDQWWknoDY/ws4kgu0oLZSKGi40jIZSeuSTkZdiFn2C+LdEReTffPvMKHaj/abjrZN
QAtVky2gttgTfoSFWMxRu4QZh67PgyYmCX9RE9KtspWY6nDCNO2gV2YJ7nKZz9P5adDPsqPKquth
r5y5dB16GCnO1d8ZKaFAu2ZVUKtTw9NtfjLz71In0edLP/NdwXGfGOZa78Pe4ikNbdvkQmtIdKT1
38NOj2yDOL/xujKD8toBcGDoCZTJsztTWEHOHaqU9Z27GdHzt7MdYU/tKojJwIrGY+AO191YsRmQ
DBys4Ykqz7PHXRbgVM0oKm1o/yiYY7saQqtx4uYoFi6Yc6QU3NOWGq21L5HjvxE7+3s3HbKy6Equ
lcEk5beaKVLB9AumfrRz4sbTVFyFk/MKGiz/Vi1aJzfZIieqJZ0C0Tt4LIDo8R5eqO91QJIIMKNh
JeGGTlmmxRi/2BnmdJeXUVgWPNXNLQf0emfI2/iKXQ3KDgROlcBuKFeLYVRpP/8Oo6FzF+yIG8iJ
oOoYGATbE3NcZNnrURlhs6jdn2RXRWHRvbEZRsH7cYKYINkjFPfqjM8/yOlb1zhZBubklKXdN3rZ
C/GqK5oFPxvlT3eQnXfP1VTcgxwkm+zhlS2Lts7rRn+VCsj3ms7/Y78zLiwwCSQmoy4u4lmIdyM9
CEq4E36VlysIypH0aOCNMpvlKz8XfTWEZQEW2hTiiC8vZ11tslwKxNxEXlz4w87IreeHl4rzRUho
kRnhCPOh1T2ASN0XSv6BW3xFY/XEdB6jAjMvgWEhq6ewssSIjB5ylbmv0ptg6ajzY5EeX5s5cxw4
s+m+xSJFB/GY5+u9ItQrlqxEU7JQkKNfWDMzJiSpzMRwKBxWUaJX4Un80hAvTUEyiDnRsvwcqU9G
T6Gf/T+XF3MWL2rLz7B6Vmg4ebuVYpRMBnZyeHgwajzQxrveXie7B8tGYxRK02OnpKPSUZCTc7nd
Bi2iVazkq5iBibzbl+KJufX+mjTxUNQJpl+0UrOe2mdvoWXB0B1zbSfFeJXrWhfB2sgOwY14XiS4
Qqi3mCSXhDCQz1Y5eGkuMgqMFUwLqvEXZdRD0NISTg454WF0pCAm7Ng9xj5/Mj8H+f9fZKL/LGwS
ZQZsLqpQ8Bq/zE/GQAfovQvPC0e+MFo7feFW8Q4A+9M81I6T/J5vAN3EapOgVTBqLyjqxl2pfMH3
cjoB02WHhGmRlJDLwvEtP7mHiWK86g0p8aiTzSb6AVDJN+ggMxnaDolHi+a2S9u8PlFr1j4T8BTn
exOBia10dnB9sugbU6mEBlXvxSIMLTsnRxR4kO9mrl0cZ15H8yayjXuvPlOLRgWDjMuiac+1+WDs
tCvmYjC23pBY9tD/Ga44ml8usYJcwjZRVClqgnGTantofcdPGDzwGd4zQsR0rBDoZrzyt21kb1Qd
qEfRGF4lOG3M4wpdTuBhmVWkDHM3cwP/oqlsiSvjPMx8W1TJcpzSrShzpYcHDwXDy2Lrh9xsmV9s
QbFZZAqhPCRkumG3NS1yIAgOC5L+UX73S33GEWAx0RvG1iXnbI48Rja6oR6SJM8k6x/JVApb/brT
myXS4PZoNmN7BN2kv51+YySl2qQXEIQSHpNXmgHxq9rGXVenV3SFw/h7RNLifQH3PTtFUwmCRT8g
lQun/cnNSRbQmciMypWyXS5Zg1SXm4sKNcV0C1TL10oEEwY20qgSKWhN2CdyIyRyzHhtNJYpQhTQ
Awk6XGZfbn6DjGHM8m0HapIdTXLxEw9iBKhU7P1iMQmNqWhxlZPhHCsVMCej+UnXGURyIVKXcnmq
DuADnA+FX/7U1K5xF7stl2O0KzO0Y+pFQScBe2EVlDaqCINVVrig28hq46ylCwPGKEc+4uq/B1Vu
iNwparllNfmy7h24osG/HL3fB5CdGIztqCGAI4BTOhxGsq9nm42Vyr1gS2Iux6wfpj0WKZouyQGs
8qlOY36e9hhpVUuOvajvdQbxdHGkmt9DKShbjSDxTEAeAvo8NDHaZyUsvK3isYzj6rTyhNXqqwwx
WRElBAmfY2WvW5k5sGewWmOZHM08rnMrpLT1fg/vckI5W13clKjc3h13MBNLgDU9NsIaEPhj3WjQ
6k7k+KJoZI6Invw5ZMfD4FWaocUnJzJK9G/zAPnPA4LiOGp9nI+7GhJLWMW2uB3iTgjAsLgZr4RC
PIzteheOgum1GchlbM5M9s1se92fae1WdwMZ2l/52Ep8TCRpJIKHDgmJtxUzCSfMDKFEfwTZBEZO
opTtVvQTQaP7CN2XK97wMxso82HF8OfsHBbixdAhK10aCXIPv6n+CngGVapFf15MbKs9E7tLeo1K
2BFwS8GxuU+Jz8BJ2Xsp7mDy3VqXbaLddHdGsFlOZlSG/mUfVKxXTIPvipfThWE6wyyFLLJiiKy/
MPmzfzOLRsxotkQJENeu5Er8MjJmcrL2lKU4AJ0gBcRnEnIrqfWo5zGGSQvTe6RKXZH++AcnW3Rp
ZKsaYs2yRqWZT7FAp9bgE40VB8PINC1JLh+l2i0EC62DSbdJUS6qnX2wjc/loCip8hJ7WC6VNJuA
U+USp/VgJ2j3sCFVLnLwKNmmBmjd9Kz14T9BxLBLSPmy2LG3pagPOMeDYAUu28YSYgs1UWouqT7c
EebgaiTMOd/MmL3IbwX5DUf5WZlZz+08iVuMTB4YQvZNl+mO5Zr2Rvf0JQ7CTvwC1qv1moWs8uSc
xoR5KpS3BA/kZ3R7+Y2nbT3yW7jVj1BB4j1nIhYN0yEzUlPobphAy29o55iSlRBK7BdYw5r0T9mI
Tz270xCp98ianWqNakJiv1pprO7tNXHaG9tw0pvfMEvLENx8UKHbG8XOEpM8i2nAIXD09ceTj8PU
dP8bxxAFYi2LmTjgp6W/lFiVP9Z9wFTz1zsTDRtB+ZZGf3I5iO/voAUi5vzf4MNzDrCvp0hsKW32
cidtjaAzqN9qTOLHtxCc8910qq7fo8xwskcK7HjjLCGuOeJ70mjdd9jr+RrjD1M7SRIjCvObrX01
5KV1TnNbiVtLZvPJUT7LcPqlvyCODrrBaet/ami0ko/Ok2G6HxY3/3GATzHfU9jR0+hcWAHTwy3f
p2VawGotHQnnwfqKO5PEbx6suQl72jAHAJTtxI7nEFv2nky074dCvXxGLX6+rivliV4Po9DVSSP7
Gfwt1RcK41Sapc+5C4ttcqw57rlCYHHjFQemgMjQ9A0VlOSMzoJPiNB7cwhaRmR5Hu/PaGlT9rvy
pVmj8O9hXNa1G6ooh08fmNGrkqPRWRb2DrVm2YXC+5WrBvONdZeGZu4/9F8xwv5HNvoJV+/SwiAW
w+WpIbpmrYCSj2iOrOGwvTlhFsJ3RIwYRNKfB31jS6IuvPI9oYTXcYElxK3AeQk3fVLZ+f+AzNO7
JX+qC0kRVRnGstKR+omYXjYKi+fSOwbxYNeKEtIx4m7gER16rKDbOCmW5OCfAR5+S++FWHZ9bl8w
IlBUDpK8ws+THup5qX4LXrXcEU2nluHfpTTVlkuK2Chj2kXDfAVg/bsHCF9+ASGhj+PA1J9lI/WH
eR0NiaEOUEtAgJW2enOI6Prd23hbLt4SbbbpFOsdeZspFS9qb9oAthx/7co30fKTG2XedRoIU/ve
mzQ5lcN69djmfa0f0bie5xzNf4mHibaVRF/ShzBSyCWicnouWmnqNNlm898yd4pV0Gv9wBN+h683
nMOfqglXCtR5vHv2EjdvkRSIwp8BglZiRNWiZBfVQqAlFy7isCYfGhL3n1BjmD2kyP+PPkLYXhOR
YXujQOXer+9ESLQndWaOU9MNLIN5MHPlfbmWCQU7ytyMm3Lw7LA+QoR+fieduFYIwr68J1lc6xPc
EExKdW91echt1/WstCDn23xVgLdMVo0i3nkUbwel3cRaQ6eerAkbYprNwA+Qcg3H3Ce3yLBzL5aB
VHmWBxN0OOspjVEFfbf7GuwIW1leFX/FKEe04vKZk8RiObwDF60vkm6BhdW9aHZoYrSFC0+wYt+c
5SDXd4CMZ8I5ew02nfC8ksnWG9cY0zL/XmEKs7B6N+BMhlTG0NvWhreGAS93yt6L/+5u/KXta0ZG
WMI8DGngQ8MmIXltUnp1+LtfRZnwWydONDMZ86Hgam3GsGMqSXa5cI/Lja0Zp00BOvpQvdV8hQfG
TzWCXJH4RDCiXq+WzqufAL/Rw1ZAMqzx7CnYVSzxRV8d2Po2cxnPv7rbEEOXEmUuYA/irtU69qIK
ZegGON8pMQcYNpDS9EOR/aqgJW6ERPhUmyqNV89e0jL71eZwLBwX+efcjtns72x1LUtCRBw1F6KB
VCUkNBMm8YYmmBzoyFLC1nzBT9DP/TgvlKYKx7YidMvoNDZ2Cx9Ogy8JxSqnf3arb/1cRcJ1K7EM
Qwu/MvHL8SPKrA/6rNv9+B7h+tdluX6oK0XeLJgcELRC7rj2sBHRpyGsj8k6bgEjyshbSq2Z58Gd
q/mJo0Qpr7+hgrOm39tyLHkRnGbTZaLF87RlO4Os6EiOTR+TwoucdME11VqznqYSCiSPFYBqNArn
WPVAzeiRSb62CgJiOMksA6AFtfqZSoQ+ecBIWQv/RdXSs5qQj7O6nCKImf8e5RFJgzEv9BiQ4s/Z
8QPbC9/ppa3r2gPgm8pHQuLWfS5CAQY2DCkRBz+O8jWjjGMW/EIyEyAFUE5lG4Ufpyx14JRVvwlC
suP20Bfl+6kbqu5nUaHRw0JtEKeM+dN4Sg06Tish1d0jeT1FfulPGVyQsQ7ZivrAnTPtV9Xx5O+3
RCSV6n0K8Hk/eMkMArFX3yFRkoLH5ObWHJ1R1W+C+mUR/96L/ygWArMd9E4xUWxgn1BQvhLqq4Ka
sIKpudpJVylykElc1V6gNuZZ7d26iJpaLrNDa4ZtW2chulECL6rTRl44Z4RFl5aqLITrGZob8wbY
tYWmh+L6zNPsPd4SsQyZYu2guGKJ7IT3T97Z3/qLn77yJ7ZLJHhfr9KoAzq4NsS33TLVCpxtU8wl
8+0p2ctulfsSeaOBxayw7+mGrU7TwUErwvZEIOzW3IEyAKACLghPEHg+ckiOsiaXI2QtDnKKxFfM
vUdrSytB549L3sPFn+0WqmV0xGU44gSe5uMhTIMABPzcFoJqbRwIwUhGUSPTPV/2nqZ82rTT2M93
O4IDgbGRkeCGYyy7fV4BKxuUXXAbIcUNsr2NONS15/mPtrTQG+cyWYpGrhgG27xRPEcx5qida2P1
FII8+os2+QfMzpixG5S2wCwC3ytk+0J4Ue3IYKQBJZzJMyS+7Uu7Osy+Pc/+lyVayjqdqqNCpY4E
6Nl9kp+OUzKLrw24MMaQR6Ku34Yv1vV1vaAX703fy9HmWqRWgUfj+5Jk3mdD9H/l1sAbhK/xJE9m
Wjuhq2/Nd8ykaxwUxDHlf1yQ1mMEkSrmGD+rxjfK4graz1mtyl+7Wu6ayP/P5yZYbti51j6iKlld
rQ+Gi9vpcK08X2P9WM2ZeyC/vEdYRCHg88+x0bhhRB96VgpEO9l4rIG6LMRGjZajWUS83chX4dCv
Amm0elF29Wx5UaqXaDEmBsD2ITz/huNzcI/B13dfQ1JXyHK2cslLFuk8oO0g6gNkpWEmvpawN3BV
XjVpVGH+Kfx/eEzLKo/LyYH5jx3pZxkq9/ot1ivSjfVuMtgXj0zc1L1MNfwERd+SS9hUbnWkQYz0
R7ocL/gl41TOsFw1wtvh6yT85Zc7o+M96uyV72ncmjBU+DVKkOl7dgm6B3FaywmQQxU5BZTK3rJ+
eZIycbA7Jj6Fp5dTcfNZ/tps/Qs2Hj14mlsFzBtXgt8v52+J5+TbuDzpGnlfriJIdvYw0fQbqoFS
BZp5kPSeMODovosdtXcSbuF5cANr+b/OcrEB58d9GQBo+L8ce1dVdfd7OmX9wZ+XPJrWLih50EOv
YmEOtjxZ4s7Uq+x07gpGBLbLzJ4SeBzVnswE0fez+4JbW+78+vs7Grz3HqYNX6UhNtv1YPd1IgDW
SYzmfNmrNvxrQkJiYMgeg7NbIJTt9tURgQmeswvCJiNVaJwJWfzn45I7VKY247RAhqCdHogh92cp
qc9pLuvcFvajLkGwSgd3EEMh4/eKcKHWrYDspx9SILv9Yzbjc+5/Nn9oolKkTbdkI+vGuEHkkElU
POaxQKbfV1CL7xJI/D0/apuk+DRSfKK9VvctfDuMz8DAKCOX8BoJKQtNmo6V4jpTLnA70cs6H7bY
9mseNv3hN3Swoz/ugATh7/3JB/4xUauZfy3wuRd6i+xrUNBrG0n1fXvp6wQo0Kfxo5+ymFwPxzck
/eHOp4t9PmAAJZN/4lWOsR/IAb10R52UQIPPGcwcphfs6Jwj2r53ZottX7SJ0WLz0mVniCTLdnin
Rib9IRvYVRdpzIWydH7eXY7kVEsKjkiknR8Gz2pyDeDTREUs9FIh2Nm/jYJIxu36kpebLKSzYK48
rjZk0t/JGUQe7HhduNfa8ncxD0AEAf/n3VWipDUzuOClAkb4TgM7lUWEsGJsXmrdY4Xo0Dda86RO
tRHd3OxyBFye9sZeQd07un/fskuaoGAPzORoNpZviSn12ROkP8/jGzihPswl0mbW3uRgurYG9jpC
EoYWBUiEWuhxlr5toMbpkpgkUpI9Whi+I+zSIoONsENv+C39Y3lXu0qeU61BjZ9firUS6DBKXnmt
l8xY2OniDCGtp33INH447ibJOoJ+TfXNGOCl046jWII4JGZwsu+cnt7SFJVxr6k6zsO+9sPJfY6F
vwTKSz6QYLou5q+QMnvdzvaddETRyN5DZ+FTW4o5S1OBOxRpinf+2RQvHJoccp1stQD7wfhMOQ6E
Mq5Lv/DS95dIuUKhWX7E4BPTRKSjeC5z6FAo32RGlWQe8gGABBcBVo9iQ5qfe3r4fzKNHTHAOM+h
aYjUB/xdqdwvMfha+S03rS8Xy6OYoHTqmuD4PHrS/w9HLNFUyIEYmXB4XEJ8jXEhPJIZXzRF7Gyn
dbicEm/jHBKR/rhFK/iazMRgU3OFUZKIwyASNTT0/ZLvFOjhbHcBQB9aibJbnT+ciTFXtzOlEuzW
uHLH863qAuTfdBF8aHF2laeiCZyvYNj4ypQTLbU9bA6uM4qfBR0bPJCcG6nU6HjS1HR5dUiViH8R
iSZfzzLfFVXZIhV3GlcRP/ztQxgochPKIJl77yLlzD3pkWkU7oUvBJSP+3BNEq1K1QM5xzdzLo9N
TuCaSZe/barv0ey2WiE41r0OkD/zqwVzwmmAbNj8UtvY6v5nW/9iVBCgvZoAYJFygDDv26+NQHRM
nqTe9Kd5K92UdZOBOseka+GV7FOky1pszMtWQG+zMA+lFK7eJXq6EvYtFWQ+TQVlqMoCEnBdHt11
qaj3geWx2xzbecVxsemTSn083BQe6SSs0zcXOqxnrLW7CyqLTepIDpbzQR3OxrQWw55Wp8EgLvUb
3pzmi80G7+Ciwk3jVZxpAw7Pw+VIqmU5BDTyw7OX6ATkWUAQlpKdC0La4nqYdqkP19HzGpbbee+8
wTQvQbIeTz3goY6jtIGrZ8W3eK/bWAJWLV+J3hQ1OkPalOCgEXJghmdfMREBPS6IoNIqQVUUGiNJ
K5SKds/r7vurnV7GIR0ED3mmySlo7YA09TCw5fQnYFW0SG9NK43B9LD8bGpLJxdn5x+SCha6daH5
KL57uANy+YMF1WZi1h1Glrx4HiqDpoN1g6drIFigKVj4fx8PX0ojYPXDyF1jVHuStVc/q0lRER4k
+SIU7THVSkYeR+5dQqADp9jFGPOeh+FG/xJ0x88DoFk1i0cNY3us7UMf83UEIHDW9CDrJ0Tx0/1I
egzYhkfHX3u7vQ3Ysdls2rjywA/gtcb+RXNevRfW/Z744dPfxl987JDPbzXg+kxezelKHH6WgZrx
3w1vH9xeXcZTq4McNv8AMsMf9R4hADYHbypoX53Xkx7+s2i7Bu8hRQIztowb1UN9/4CRzOYcYveP
TZo5GiZ5AfHpxBdP3l0o+xVBU5ptxoenOOpZ5YbiK+gpEG5N3ufshgrFLzFPZXQVGiQHQu0ZjwYq
bNJEz4EipbwVPgnkNkzKbwLug8kT4smJCRdaMshiLqASmQWeV2i/wlzT+pdjX+oVRROep2XVTXuc
fETvXSoCaoZw8kHhsezvBMGyR7Y2eM/Mvz9ECqRl6XEnadcauGngQPo/i+8nMHeEw71hjOKQgrXG
fhjXg15DrgFoW6k3BoBWnoEQKBhIlukF36PEPyHXOyfSJgR5JBWSJeQ6LUkdRY9z7gbNfjkUWSUt
b4JXnWQc9Q3uHVfE1U6YGwqJrJfgSjcRThrobzZBnrxulunyXxKx3sMMRhuxHyDINtW59OIp8kOi
4R63YnJdX5Jh32f9QeZwh45rgwpgWKZW/lUWVZqeF2/P7rieQrEi8+MD/gkg/c3DCgqLjPejNx7i
wT+9cljBz0DnvbO1MTKFBmabh8ApGYaqqnbRiXmCOujhSzMzWf+820OplyJ+VTcaH2Fuirop4CIL
uqRVDPaIMeTLGLDPbY22+wdYRDFZwfRFZIfFuxY8+QgVEdP2igo0Y73utZA/ZcJx6Km7GzZidbBM
dt9+jsCFT10Kk5RJoc//ol55s6wrEfu/prXQ/ZBRb5A7cFqgbFYx5YY9hn7cIUXaMltrqulRkRWx
vhWZpRTaMV/2+prMX1iO5q6f2uSIGEhZ/bZT+mAQQaSZ8SJHeEvVBA/i4mK8wOb2WtgY7Sc+lz3y
voPuqPv7PXf8/PjZzHDMX8tJmEknnnCm06X0LM+eGBlrdxg+3ucOHvFRnJ33/usbgSCnHb3C3F7Y
a8DGjgwNiJJgdZDpj6xn1VU74TVK6thrS6VDfzyKi7xM6QKnaI1SlnEVtMm9mG6Abf74jW01ix9x
GWFZtfNpC3feix6ocObt668KrwMDxAoGPy428G2W0I47HlKPRnX2TpcvskdTTT8V7h6BqUAl4Cw5
urR/PlH4oP09xAnZYh/23fakyzG7HAdojdvAPImUMuLeD75T9orMmQLvFl91ySGhocMT23IsXZrs
nejIOt2iE43hpX9SvnW33z2EndIjdgVrlnzwQDnQE8/fY66ZuSS3+IuEtrb0SARkcefOcdU/+IKN
NTBGM9v8rYtWdRY8vOtbN7PxOf6xCwgReyJ75Yh4K0AbeKxDO/zmKHoZ9Gd00q2l6PFkAzSGOCw7
NGk9DEYNyZqgvrk+3FK0z0qVZDQDzVT+++eoK9q9g6vqEN98pfuxTGmrvh8tmlXNpRX8kmCUmXDG
y1/29yQYkGbSMN1HykTbtA8s+gJ5h9SsSnT6SOlgNo1htjjGm11frIs1tfdfBkTOMVIInNr3yXfI
Fae2GEFEiN1oimQzwDTXs30C20J2u4hBo1ElX5/0GVzZdnzkdpnES8Fe5sbELhMtQzAu452/N5I0
MkplOLwhABsPm/lAml5bf6Vo53zWPF0zdrXAmXph2i2HrVsZpTI0DuIIGJamDawH0JE7+zy5cRcm
6mIeRUWyQ3jf1MfwGrL5EuR53Eo3jXDUY9DmJUhI6IiEu3c67tGdadMkTTKuaXCgmtQi3I97wthr
+Zjr+GFRdW1oXUS7qUodkPjTkUmwPi8Ov5V3lJ0+cdkCf9EEJcFCAu26UMPXZeciqSxyNpee1/4O
2qzkpJdErYZrN4czn0/IP2WU7O30M9YU3SYlUGRpew+4FaxEntwTBR0jO+4giKLlloIMNa6aCk8Q
UI0cTD5xMVJmnzh57V+17zB9nHUAN6cLeXXkqONDSuY+ZwT2EnhRA1YKMyPfmpA+U9jp4f0rFqXn
1YnYtpi69HMbBqhZQcURyBfaBuaIGG10rfDufdGo7uDFYCJCx6/pMNQiL5G/CZ8ePZHrj019jAR7
GVAzOQgJGfhGppNc8c9R7brfbN3PhbxQpTEbGMu3NOYjcmONl1xzvdO656ltvMW8ZoIgnLPSE1Yg
8J7KTtRz+CLIQD7Tu/Vbn5MuhEgIl9ZTHOper0zqLm+cm8pjKX9uIgSdvoB6h1bD1ve1EeBnkjfR
P3y1SZa9MfHNxMVA/oVAzPqXv9v14TFImz9fk3gwYn/KmCwHL/DY99b2VxZyuz27ZmcpoUe35IeT
8fFU+gpX+NZJdn7v9UFyxxQ5EYMXF5szC8jgdRoBW8kn6NDpr0UUNiJ+wZICMCeUdvrBs2Qz7mXc
YSKD1cic85Infa+A2gNXClRIQx/Pih0l2UfntgPphIAkjipkGIDI5sWKy5CzCdp4f5jUWOF/rIze
bM+YSM1IBOlxry2euw9xM+iD9pS9cVFW2AfX2ZC29J3d1O0u7pN54oFEYyDrw/03B5UzVLAsRTnY
c3MZqvhcc0+W3n6mXFPu1jduYUBIn5iuXvCi0kTst3eFlzjt2ktoqHCqx897dpPzI6/djOuCM12B
ztEOqErmhKjWaVYeyMRR3Iah+wal55EITpP5BcO7gQgZ69vGEVWAwPqoQhTQCrKZrHy9K2UTTGx7
Sc9dHFKXhxUi9oT8PUcogdymY6j9aNApnaclCLq8pCXOxVIbNUJnI3oWhkthuYuR/q0nRkDc+ba8
klk1GfOh2jJgfGaaWKvavUTqNIGebLdR3WjSs5YItEm4Gb2mcCKizs3qIPmpbQgWdGfFirtYMZJF
bamxKr/liMNFbkq+yWCLkRq6B8FPRtUEr2ThGBa1cK33+CVbbrkwz1n0+1i12c2KBZ3h56NUKfOY
GQTLe1F66fqHceV3HKBkfeUkIAecgW58bdT4UnE3koNB0QXhTFfRfuKquiy2mOV6UnYZozTJrS/V
YeQydqVA+A0qw2yhgHohGUPxRjz6qBY9x9GoxZAufCKOZE+MMbDyZh90QIkuYiwcK+bfgjuImBzM
y3lCxz57FD+jIoWvsQzyoUV1OLhzuNzqlY8Sk9KYLy0CjITKRutfTfKNGeagPsFtQUeLOhe3Woul
ToyMrFu8AxanA8kMG9/0/fCZqkn8486VbPQdkrLtpLsiFRFUbiPoC88E6RgQ8aupta3hjAUpDLLo
RYZ53oBSoZsZQkzIeKeq8c8RobPwjKbP9qa+rm/5zi0slHjelJDbTP3kqJqL082Pke+XwlwfleaU
BMbtT1lskCKDttXBZWPKIbYOMaX5UYFx6fOAuojpMEwQXCLyENfvY9wBi+ucB8NLJ3RWuxuO1HsM
a1xJIAiAliGkIcurNZsy8PyjjxczjALC8Vkp128U7wR8ZbLjX7EuNha0kVM7vkdpAeuyPofYJwJl
1AQgdhjZP/6KDBVfGD5LwuXAZmeyFqofSgyx/hehsYQUUUlWp8DF8G+LoUuX9zIUy5fUGuuXXk7A
h/BgfSno4IIMf1bCA3OvA28Y3gnMrZ6H4ZZY4PROBXbe9qWoOOIEdvUC6/cMLHzZKz83zCEoLGub
gE6c3Fj+tUPHRBl9q84L+ooQjhiHrtv6p6Xcj++C8THcGTgO0TI6Ra7JGuh/gEqPPvEOpUX3ZD4i
F6Gcp84/on4BF/PVOEYwzMXbynXPEgVjYPjHMMtUKhed4ahPlCrJt7i38ThVUVdXKKRt63OrH1Ft
I5ZHeEbeVJOQGAAKqxwl10xPg1+prJr9xIu8KwKIlklfiXpJd4Vu8TuD84+K6XYssrv3alSIDwxN
ywgj5QPPjoJyLjodPdDxl8hyVobmvj4nhzBz2RyTIKOMUWIC4PBABRL6YaXfP84QB34KkBybio+t
PNJpZ9/6BS27p9yv9pBcDsRkF1JPX75ahyIyOD2MreaP/z9clPiqErjDLvCVaMGFNL7brF/WsqEp
Gs3Ef4lCm4pf1YFiiDXZW0lDsMCAssMO3eJ3KGAUQxg7UyydYgZr9pm/2C5YQFJ0bw04DNpEgaCO
sOWXVKPiQiv99hMjRQYMAg6TuIV90EZEufE+gUUV3XO9KXnpEeOGLadCCd+3r96ivOpGqK5bF8/1
N29KJqiOxGtuqC5DjtttQ52uxOYbF+fp0VsX0SVeolJWCb4GotpD5KArQ70hmSQB06s5Ozfzs3Q1
iMH1U4d+x36fY4rYxGtVOfRosndc7Ca9+N2zc+iefUthExnO8FYDpTmrF+8tDuC9lbd7Le09VsrC
Qi8/J+UfX4w0MN9am7NMv5ED8bowinku12cjYl+0XuDd6gGMhmo+SMI7/rfrSTRmUUqkuAgZb7M5
ZnTyHkVQ136tRf58HIw24gfv9S+ef9wQIi8fMfWbYE9SbfIIrvxbz5DBTitmp5T8B6y1MUb/GU8h
nQ6U55PV3zfWfc9C5qXbQh+JozQ38eOzwHt1xkw9b8420EknvETFjlC9rxTkqTIgDyytzKtrxpsr
UGZ1zUrmWyi5YDXcIbn3qWLA4sNOPl5BgOr11jB6BxTX0J12fpcGv7ZHCn7ksJSNYmtYupmnbEAl
wOlMNk5NMptPFzlfhzwDnU9lLAxOaWlJucP9iuw9tQ7SHNoEZTu7MiSlH9BT+R1Rl6ds5AzWoR41
of3rHz2Skvh5hI2Eq049U/O2PnT2/qUZhpRqyEiUEyE/s63tLU8K+K1cQkr49rq8YKwLubTLKaPI
Qhut/P7cF+kBC8UWodMk1dCEiK7+4Dj+Y78Y+YC5tB2ZERfZOImfLM3o9pBIKMk4Ls42QJ1PUFM/
PKeox6RvVyMOJLalPBVjFoL32l/+Ao4yFRQWuQIfEHXNStWFfl1iy2UU+46Wt3aIftozwrsUYSkW
keAvsDnmLhgnhJ+uLmtvrDv2dSy5v81P87mfMFTqu2QEhkw5e7CCS0OOmTyib60Zq/ZvL1G+6WUJ
NxnLVMzQwoUQxDP4zTI+R4IMh5S6EufB34YXS7go9ZUr2B6uVwhkIpWEcv+kjxQJVndNLSiGyrwJ
56rqDKZmFeDk7DHDc4wpeuWeb8eGjaMXVtSIZcTVt4ZxfkHWfgQ2RN3V1Wz2ppMIwk6FtCKGEl9k
rgra1zDLjyOQgosZ4TopVfNGWO0Xgv9YHLYmfVr4ikB1M/rhixNBnhiRHgZXK6ZYOV+zNYQ9wj+2
QfoH0ctKach2PRhw2DR/m0iU3AqaxSsA69dfs5FCEsEHT+rH0luAL9MtdtCAUqiSbhRrB19nzZNF
SYDEkbhyTKcnzRMh9O7iaNHfrLBwsYODn0PwcIORxLMirWxRkLrwfM2aZHSWamK3N/e7YTcBZpfU
Af1gN4vlHUjo7b6YM0lZVBKnEZM5QQWqUNRa82ytbvr++LpR/uSJZQa1SdP+dQt2IEOVhUTb3UDz
7Pm7qye8w+KdeDzvw5Pwu030XmAQ85wykqvghZhEB04i98rEOxYoCr1qhCego/FeObqf2EzkLcmI
hPmKbS8CpBvDqCB9OqgafGfBzblbxgrzFabN3j2/bc9nSKVxN/xeeAwd7qNd87NA2ZG4bgVcaeDn
uQdYZIXRY1cTK4tiP4eYi3Z1RgVdvxyipykAMKpy5YI3Q7SFT8zVofM6opFmCx6G34egcEgNCaAX
UQ463tpJCq0lQ+p7dyZAeLcarYKPyNkp0kWHN+Xe9kj1RubtC+qEGFHIcxNTqcdRJAsfm/cqwUX4
W41z/2clAeEzv0p31/j5MGXLm100clu5bjEFzsrwRvm3C6663Z9j+kqEjwYEV91ru21z9FG334tl
EfBH9jUsZiVtnw0XCd3IQ6FMwzT51jKnZzg4vBbOM95KMGHGA1eCueZk+5CTg2Yz2TmD7zC7xnUj
v0iaZQTX5vdeDSHNH7ChhBqqVZE+Nsv5PsZ6uZnGjMsQO+m6FRF2CZFpLpiELrgyr06Q6uzpwsa7
+GASCEgn+X/iOtshMy6RAVvTv5+CJ6n0oLxVowWo7ZthNbYZvssyFCvO+Upoj95PFHD9JnaO727U
KivAkKZYpi76bXE/J/lDQ6JRPxOodx/ucnH6yGOuYqdgf8J2uXEtyvGE7a3wdt1NaWSdhZ+HWdAq
3X3zpoTrDQRWAdvz3e8HtC2CLleFGBUd+EsHi+1Ku6zbBUi6qyOgEsmDKNbn/oXmo366bLPhwvBf
6dwOJZME78OkUUGM4yOcvTIGgDzi3J60RzYTSvxCnVudgNsyGgaFv0eYfCwtTLRnbtVWaWRdw70E
e0QRQ+/3Hrwo6mE/RAZ+K52/Vo3ToQH2LHoYQKMgJauNFuM8brFAyxrGY4eS+ZpW5nIdSHfHYxYl
/Tpgap1JtRJx6t5bFv7wZ6AqAk1LcIg1r/3M/VHS2diks51qfsircmLWyZ5Ju38YCvV8qAqg3bbL
7oBQQJG3S5I5hoHhEu5vchF0f0iUe0uZJ6skbo/YAtt+eldb2qlF74ZteEnE8FAYAgiLc1trjVXV
RuxqDCZobacjfH8JtseYFm5vFaYC+FBOYmXAuKcU8RmuUbY9ZeJlGIZVg6Vm8DdiTUTPBNiuVh1M
4LGeGcgXWzU5ddyUzuftzHo76w35JJcVi6PuitjS0d+kVt6wQoGAWUmy3usxYntY76o+Gsd09uYh
xv7O8GSJeenAbHpo+EVgiWOPyDByUAfak0ty6Wwy7GAPS1OxnrZtztBjdKzXzCmoTd4aq3w8JKm/
0H8M9tBZ9ETEO2uU9LHbTx/vE8prAgoC2vsQ/vYcqluTL+1SpctM152iQrWVpVSeY1LujeFN5egZ
hYozUSRi0yhH8vfH7LFoiql9NxB7URr0EQu48hHS5gbT32UAIk26uCwUdxVfAE5h3IJJKFfSpXY0
7UD6IHIx3XERFNLlheF+vuGHaJRpQeEn3yiZHv7bDJh56a0+14JqwnDtL9SpoaVRg2aRF2T7DbOX
u7PwfhPclXYQWtj0MsYY3KBM+/c+IY1LmEZi2reI42Q1zHXyzghCHuh8eqzi2/icHi6xRWJ13nTS
lU/5hTzBj1+Jo40aUzbRANzLeiTOwxwa4GyWiM191mOkf/MOIg54CV+SP+0sv9lie3zLdXfe9H47
jtd0naDsL3ZrxGtbr3g/NNvVzTvtKRqQtNakZdBPpxNPJRpC8isg1pYgvIgc8JMc/g8ENPOa+X+Y
AP/p3xDVXi5Ci135A69XJ+EtE+oF12kFlROj2IixWZgB86v8/AKoeNLfDM894vHjeSkVNAnuwZNK
H6CP1U57P4ryeUG0nDAkbcYTqbCgaSzTqwwtKDEEJD68BJBYtV48sqMJvoeGMAlOM5S6PzIG/qfu
ssVjB7oa0JegVYt++X4dcNUpj+KehoJG4KEZm0mbvTCTtHeX1uEsZlsmTkm8ySmzbrhCK5pXowKS
RRiO2X5o38E+OUwOdyci6X+UFCR9pCsiq6KBqX1SA2nTDy7Q03hgNsTgCv1jrNHi4J+/4vjHMdYy
+4EiEb3wcyJ6BcXDoa6bsl+osD6h2/78tnxXIaB8/OScygJ2he7jEpli+M8gWTkhdih+xlxyCxVm
+ErJ/lu4Ios+cT5G2R9FGroNiXywDRR3XVGLjwsit894IZ9li0OkHPCC2s+QUr11Jfq4iGp9XxSw
2Phma7oww89VbM0B0zbPxHmXPaeNbXXKdppszHhgDSl8Jz+sGnO1+yLAj8jaYGl1ifINFSlZ2uka
r3pv0H48P/trs32i9gam8Z5epZTFqHE3v9BAzO4lSSXWlNEwS4d5a+Iht8Ccc4BshN5OQLVglzFO
xKYYrq+4v2DalNdir/1Rv5UkNeVDoB/dJZ+6Aw8DdNeZhVkOK1HEOO7I4fZ0kzm+CQWbtWSL3MEK
aXJTluqf6I9cVl3nJBrMd+iTIn8nhteWZ3VvRj/apJImn6Stc5isOnUnXhzbJClq4WYP+xtTFFxX
6LHIC0XuPrywYpclZDTki8Hb5p+QMqXFmyf6SXRLjjrTwq9IYpTHlbqtWy7LNqkZVFs1LxMyZptM
N6J9qf17U3ev+5TXqKBsjV/HH8QtEU1xytnqQ5+lWBWskUWEZxRfzsxhWOrvYYrw78yNLsDbBk3i
gP8rOD7wfUCNJO6SdYe33IKBjAX/H8Veu+1vHrhBn+1aBHo04iASfDeCVUj3f2qNaxXGErEhXzsv
ajgIS99teqQtq42nieU4621JeVuyqv+CEuYX3F1/G/gLqoI+Sa7K25ntPkxx4fNS1e2QO649hTdB
RwyUm5epaIxPwTlmMzeDTtZKzJoaV0Cwej36AxWTlaNknK6RQbu3qzlE8DaVwId39EFnjfBomAm4
8joedlHIRqwUGyL5Edvi8GmEuj3+E2Z/TlcT6uNpJNevKOIUj59wsGsn4vzfZwhlNNtkkZb6Awex
CjQf9tS5OpHbqqvknGWfN1xfPco5vEEeHoZVgX9uljd1Iv7FAlQ8lVg5nXFrGIVRT5ZyUv5T++A0
5zPfBVW1B82AJlzFH9QS5WTXw1snPefkx18INDHAfHrAJgLpa06OYkcaqTuudbUjSKF/VVH7Soo/
RYj4I25hgbhUVqVjzLG3xtS2F0fepsA+2LL6F0FTtGKBnHbZ6uD6F4Qer2fFj1gZekjLSc4L7BJu
ChWyBBf//dUqlbd03k3W4v4a7bUHZCm5mSTOURJfrv1sGIE3ihFpHm2qskjUsgyDrVPPtZDKmett
ZkkYcXxlBGYh5SlDnuGahQcjopP+ujn+UMK4FVkrayJ7TaQgIG8rs+3qtCMjmSpWlNRZb7JL9i4r
j52xFfiZc/RmxR8kQ6g6DzADFtL6AItg0qLXltMV8KGG9fBgiq+lqpg2MSG+jWtd8lBE+zwnSTWR
iD+Bmk0k+UPVAMjXsN2EJ+bN418KEN7BhQgMQryUIhOWDLbe1Ydnt2+HY4oRdEcbZCq/74KQgrlN
tEH3eS32XIGsX8DcGZqsARSaDI06Mb9dX7XSo91Avu8JMwqwNZK0UIMUEexn+7TpTsXAwfOlKtMN
jYYQp456tT0O71UDY/CywBGqPzaXMH6v0bkvUNZmccrn+rhQMQXv5d91XN7Z/mYVxzENias4dJS5
zZ+3yBHF66j075DrbALb4TqWEcNZM7yN7einKTxdXh8D4+lYZhdiOOYehOMFqG5Zu4ddbmxjZdJt
wgxbUrw86S9jfsTnQCUPYgXG2iSeQOcORQ9OnCDGAjI7eoGYc5RjPqtjMxKeQb2ShGe9ex0u3U15
SUwgDzEqXyhtlAoyqAZ7Rqpg9C0Fd7/D9MO69c6ceZKmdTswY0y2UjtV2S43u2QjbU1MrgWC+Ynk
l4lnkb8EjlgVXwGmMx2NJs42nLaRPi2TRnsKWiShSQAH+CpmWFpF8bIRSBiAQQk6IKqy8u6hfSbS
cxN/BI7gXa3DmRo9YB/tKDkTxXglQ7cxNLF+9ccnu5FDKImQo7Gu/B6OdgIrEN93pQOalsLhBHXG
Iim/WkFKS7ej1q5ZKq97B7L7le1BXuS7IrhBYHML+4TCQIoa/h4QvXZmtDQ3LjnigGF4p+MsfirN
sz5Hn3lkm2hZBSeLG0e3rahz1yLLxJDVmgkEV+4hjxY4vbLZtPOcXDePOs47MlnRXdf8B7EnUAVf
SN1jwMevlwUmHrwYtwbOentGaAAvuV+nVys5eUN0v7/DwjYa9r9DnRmypEUWqbHUjo3g2KQVxOPF
sa+vcn+BVmbAUXxgDBClZbXRarqw+ygZyvPvAN+2UBSatEwAaZqJgDrTMg5HNahKtEp0kXL/6Jed
CyAvyP5OCicbZGWei7YU1rJADi42wb+w9yCHbqP/DkDPlrGFnN7SWE0Ffx3rf6HMVUcpBjf8EzJM
wSaPGA5XL5orNHQS1Ex/VlGZZCKLQSj8K+xRZdKn5jD2Ulf7HhvBTBqsG/cuEaA9bsfarfv7TblN
M0mDd02QOBvOPiXsqLrLa9b3G35pbNdz/CYTqiRMpIWXugpLJf4uYtOqDc9UpctX1sGVxldC3gw4
+8BUe7eyxW4TsPVpJWNwLMk9kCOpAx7zsHSj9RYb+tAt05Z4gaGNgejqty9AH0Y7Y8Z5LGOpiQcf
R80LpEm6/sTy7sXazXizosaR7H2WnUDFjbVFFWZ2QU/b9hCpyK6Y5gcNp+gunU5R4J3As6yP4X9u
1TqF1RxrSeP2L6EXqTzvlyedIobK14KKWCdJFVs7tFnQDBsuwNJy6RriB+jnyZP8SS1o6sEQPCbN
mEbAFSrBecXAipY4j6v1wzn5eV9BuVWtXXqHMt0VzTfIr3uOL9tijGaxAfdwxsS7CCRfMrnnuD+3
2ktWcA1xHRvwKO7SXpiEo8a7qDuRT7CGFqBd4oVdRPYHF1xwu8fythg3y31CKkUQQkLu+FCfiPkg
r8aNzV33eKG4PzWz1+DpJYKWRndVxtBpggsZUYrjNFv8IOijOB7X/PfXXRUO+JMI6LtL3K+uv317
Te9aPO+12xjpEn+dJBHFQfbl+gPLqspSzbD/FynSXGTkObn4odk9uBFefE+rkas49HNQFj5zR29d
7AzoXAQE/5Ioo5NQetjUgj+8XBmU7py80NSGVn4bqKlA+XoIMStMvawG1y3cEU82/1nO41EYLu2h
PhAiS7GNGP3e/57GK7MxFDmpwM06+0/vMLcCubEvOo+IVHi41tzl63ilB+Mfz5pdxNcV2E+wy8UA
Ds+g02sgKnvU31XTUTbXsgiTMzRD2P/4LXnHJaqApBUlQx7nxSZ7T1xuTbNBbdwKXoNzcxUciJqh
CUvQySUKQMUogphd39msieMHVg6cBvqkjUOj5cVYYKpm6Mvsc+p2nyhO0sgv4zc6Ok5ezZsbXB/z
hV+cXX4IpH/0O3FxrhExb+yVsNpVE0KAvEJHSE8l7CkUl7kp9UsEHc+L8ZfToaRmqh2tWWaBXMaT
hpRP7fb96EIwKrJop6PbDH+fF9oJ5cGZAB0r5CEXwjd6NzvM5wvCDtumnpnIyHOyim0Ocr1UdS4v
P3+hBVcX5GsNONPTEPg4S4dJBQaXpVoPSwDnfnPVcn7PYupD4WXjuc3DAN+ZBpjKrjkwLzhq7ZrG
K4QD/mQO2jC8o5ng+OhPGVZSch0V9O770fb/+jKF8aqhhNJ8mR5Zhcbt59kogCK5FY4L6RBWS4Jb
ahVErwtIXnhXnvdZeLNXiPcIDhmIHVsLSBA6RRHvz4ybKOlqF8ACXG78tcfR1x5ig7YJbC3ac5NY
MqIDBM7qrycN9tJoJek70i7wx325o8Qj12cwFOUeZ4or3QbY+s2D0VQpZy2raVRPwL5EsMUX6hXR
H+rOPZSzCy6FnLtiKpHmie0J6QoBhuW/1uEfZTLM0tWAxTanYBwCb9FyOOz/ND4FEDl9HX0HNvrG
h1AFdMmUXvFd8i9yVbPjj5fxdUJzQK9Rw/mlBiAIJ5WbBEvUWWgvKi3f/7IO6Dz8pr32FdBhSk1K
ZmoI4FfXWMZbc91Pgt9MhEf+/e1DBd9iDJfvPOvOfZM0FrXvfoqa9xn4tsbPuUCrmliOkCMdD2/r
MV1DgtoMzRd5usESbiecETlUuWKrRcf2zYgcHidCfZ/H4FYMocSNg1A3vXdlfDYnLge6K4NVFD2A
ZY7/fz9A05DTjK4QZcGG3I7uL/GzqnaL9T2Br0kjCVaugIo4roTwfPszxOSRqlXS+r9T1wdC1XMH
3H1Ry1MEts6yLd4i2aPHcMm67COV5jPlsDR5nqHQ/xhnkSswIF9W9H2yTGxt2fQsKwX3mTdw/f3P
HO2C4m0qwkeMIGVMM7OghqxDrWzRpbQTjFz/AUPt31TlmfGD8cvoNg6EwpZN093Ho5Ewvnorbthk
voYguf7HMYdg0L4/jTRdxho8Gct2THfjDl7jgD2zq0MybMfZfsIRWH9BkLG7+BN222O3N5OJiL5j
fGo04VaOcRQNCwDHp+t6tdo2HiyA+vcJY99W8p49pmFCkwH6cXG4AyhfUPf04lGcoCuQQ0fP4avb
HKsK/lUoeVE0eOqXxLcnOJIIEM/wXxMLLQHRnMlf+4tMbEQbSHsw58aj1x/FF9KTCWFAvOfU6QmQ
y/APFqwkPll8bcmKh2wX+izhuuTmtMdqT0LV2UQYO2Cub2PUuWHMq0yQ+KTxNNYx2iY0ICd405NF
v1wVRM2pMrrCJBIN65yhOMePY+9reypO7hD5egOjSzPAWI5A7I0aGMzOPYfkEuOQL9ZkLl0W7eWT
NZ9K7oxNmp6PUfybDdiD4qz32y8UoVjaWsiK5+eZJaL79bCoujzT/0P7bHOnCL7APDsYqSfjP7AS
+rCLJxov8cddRv6IhmuGPPe8vFP69gCznHzYbPx6CsrAcfUwOjHAIa7ojA7FlJwPTsUPV8YMFoHb
jU3sSRmVixuG8l0P438ysJ1pdr0c9P1OLyvuju2j8kd+fiGnljSSX2fORGx7eBqfdE0sna7E84uS
riXyCQfI5edBK3L9sTRzcItNFFJi2f3LpFsTWo7yxX0/RB4RXlsvFWCeYognjfOQK0o9eDmwYd83
/4adn14FcOOzRRvdFzQxrwQYBP3fEu4sdw2kKT/2s8BxZH+kYRfY4elrhX4dBceH2rKCETkbRXET
697YaRMMPwDBw8Tsg2qz2AHYALrJQcIVdTQpelJjidu6DvnB/+Yf/LPcXo6KwC064FGq2l5lUtRC
kOU/v5BUxb7o7WdLez75rcJ3EVfHttkgQUEdgZgfHRox16eiqJ1gcSBRK5QZQyr99XPJoiR5vedW
6BOpPbFBv8g+AvJfaUjR/R18WcPF3njzavc0rWNITQ1ClZHJWnLElepzihZNO/rzR1FKIhGx8GN3
x5fG1ZBYJRgXSzhEWIyyh5areTNO2ARz6Vb+K3hZOF6WwQ9X7C2aeN1pN+l5Jj1o8mslNY1fOb17
g8G3HLt9yr1Ggb0parS8OYqCZH1rho/HE699eGdcQXeoPRq7Feas9Hsaz16VhrTr63EEmUEox7bP
ywC796UvLFHJEZTcqmvWSv8cxcVR/T0HCaUFb2JnokqUblTJ7/o4k5lw6uVTWvEyeZDe1t3vrfx8
dqp2vDl0ZocPhbXrVtWpTle534rO821f/nqn+ykRkAR9ffT9sDo0LITTaG6PjmBWINJORk6dqhBk
1rEpu5tOwGr6co4BZFg1ly+QtmEuGueh/6HPDdn2xLEJ0HfOkabNb11TiP90BLQc+Qt2YWcYz6U6
cXM2bhciiiz9lX2z5JHCLc4vgGS2LbrkhRlhCK5iF8byEMhvBCvvDjv/B7BWw3E2KJRsipgfuM64
jb2ji4Ddo2Fxm4o11Cbff7DRDUcjRvtZaaJfd4Cv/vICdzaR6XxbS6x3o0FVtEJ6UgYZBi3GKJ1y
WCzAYjk6dWZHe+hb0PcXICbjDK3rHMkNYAmdHCwOCoKjw1SN/DxzLWqEsPzbKznOGJ+UN1SEr5j8
cMofESHfREEegqAcYirsGMOADr3guH95H49dUJYaSBOSqXREh8aRnGMXpsrV+r1w86VcNLedXJ/9
GxOsyjUQF3MYrHSikEjmdxkUGGM/OeQXMpoHI5yyxF7JoZoYI0zTjRbH/7QyA3yNiEciGXCzyhRK
wdHvSD4H0ssoNMiEh5GV0i6HjVUL5/h8vMJ+12jfb42nMHDdP2xHWALDFRlOvt27q/UweLAXVsGc
4soc1RdWEfGmbBrdNzotPj9qpynA/Pl63wL6ab85uJ4tXbYPkgMulK5h2OCw6/JwJ4mXX0GHgPMe
i6MGJEhmopciACHvEUHudwqjhLFxVw6ds/T24Pr2tgGYC8J/C9IqnIvtFUwzmTKyK8uDTeqMtWJ+
eLqpQP/RLkyoMpXQ59tJz/waDhi9IhyAFdJXSGtJH/u3lMZQe3mc2RLUHeU8lB2+oFJ0gScswxzz
/Adb/uASS13PZAyg0G4z3xBDiU4jZ1Qqxk3wGMwkFzuTXdY3hP8FEcx58X70GSRZGFFQRx19ib6t
8qTMPD7z+u5+LeXdKhSW0fDgAqXymcD9wrCwHVtGkeuw4S9z1TTDP2u8k3GN6KzWBhgpVU99cWak
tW5Tc3zadIUnoAMAXieKzKuIqRBznpqvWTQjcUMX5WwlzukadH6vLqNwE7yVw4BQuEpTe1rnTM3m
c5R3VIdRO7di7FLMwEiqG6Yy/381SMc3EbGd6L4/FsOvVy4yzUiGAdxuE7of3ODwNfCdnPnIH4T1
s1E7RJf0X1YNHKguWzSWfi3eBLBkpc125+GOHtPpqRZ9mjzOxxOtCMGT/MQc5rVOt1xu/3N4rMuZ
dvEJ+DXxhUw514am90ETaLvu7tPY6uCNEs6uQ1mKYwFCgVQ/c3wuIXp0iDdCh/tiaoIFlqnvGu3d
Cfo/lFN7W4w3bxa/l502u/zdIdkVdahPVp+6ZSzDtModUCSTIF0YcAYUHi74VP12311tlELeXYwN
63K+lonhB/TFx8s9Yo5A36ICg6T/5PHtG2WjJ/OYIlFniGlCpMFF/F+SQJsko6SXLjyOBf+C/hCX
9MBuDFo7LfhRj6/Q8qIPuZk/z7MWPPo/97+Ubb1LkccALlpfYc7UuAx3eMabTxq7s5DkOgAfu1VP
yKWGE4ynhs2ycw7K0p/ppI+K/VziaR+l8PpTHMb+oK852KOSJWkiTIW7XNx7ebtbkhGNEuMT+J9i
2s3S+GNOlN4UbwUkhQQtWJxdi741++XVS/iexSH0KuVQBjzArExvLRqs8PU1BU2FvelR3MSGsH/V
QhCJ4VZ02Y2dS2+NcVbDL1Nk/OlR/JG2BN0CKb8cGu2aCile6bNxqHJL0+pH563+7hF96b3x1jK9
r/7NjERsGZpyY8YubV2H5UACCB5Wo6zog3vg8b+eVEDp3ie4nSLsQaKDfV3sfjHwuKVhkFPnjSMP
z+0NBUwF+H+/QfAV0P7UsKdReOpbQ8Hj/Eu1rtJTr8kNjle1XT+yHvBuxHRiETdxlAF043ZuJnNZ
FOXtN+rB0VokTbucOi+TwPTC+JNILAkwTAHjCW4RVjlrjbY1+PfQyI7S5DMZNYpbLVPjAd4RxCQY
WpsDI8QW/wEw8+Tf2kqS34lCVV9dqheqeKW9DSdYAk/8k9wSusyksHsFjrh1ba6jQM2CLfTeO8No
0SespQLG4odla4LA7H8p0K/0CNwuFZppym4Bz92pup1yWn6w776h9UTiPxsnPR3Q5Y6kNcIsN05O
Hbx2HalANSwdjH6/CdLeMZUiMqamVvHo4vn7V9tg7JueMTYmaEHXLj1TGDyKLwJZCwXToOeNRTFd
mqKbUZHSz0OIM/gJSiY5BjgwaVa73DjhBgZRMfjorEj4W73w9/3fu8kDkTzDImx5uh7DdY3UrWE7
CVgHJlbOpJt3/JcnY1daTvWEYuwdmO0/Z6Ks3OKo2ykza5GMzxd3tlL5v5Rc7PpJPwPl4xfiYD8O
vWHz4oK660xF9Sr8rxX/bYODUIvx4wnsKRQOJt7mGNvtYSxockEc+/SvXYnay/pdaUYFBbKabXix
AqVEf0ZyI++HLc4rYv81Oq5jtdB4Kc0RZrJzXmRC7fq63C85p7n3sccFyQgA+jgSQaFPSfQSg6gE
Uaev+N/uuNNh/sKn9Gfbz27nDsuB18DvowivWakT/GUsIaxEUKd9VCe2BYHzTq3G6mLZmS3ikOIK
JtJj8jLxBi0J+htzTAF4Dfjev2gLUTsmY+j2VAmzt9d8Poc200Ue0MwIoHqdsv8WQUCl1XX/cXGn
O3RajM2IOViq4Omw8YkO4OB4Ie11f1O0BnLb2Aya5hzftvRzMOQzmHPL9J6M+iifr+0F3jmJstRS
eQUQbcHCCbmlFd224ij/XI8UyhKp0FXr8sJDYRHkY3GMKEieFYk8ukogQbTINUBUZHwPkgHlVCOk
QwVh+TjTBj0P411rIBK011J+Lu7Sx49nDjEESpou/yCN2O/Yinacyxq5fx1oemDAMH1adASZiyut
7Zv0W6LSwqVZ+0NsXANUOq3til/C46YOM1V+asgrzuIwiSxVstQmGGUvMFFSJFn+QRu+pD7Ds/K6
ULAI7AnYn/FesQ/wnVuz79S8seXFsVb1JtbdzaF/TVMqUX4+tDK5bn2BErjsRXw0DiTlaIcw/ccW
QVWQNA9hYw3nVyp4uVUocNTwLpPtvm7Jz6zcFQDhar8uCWGkXA5KBk4edevDLypIDGb+bhW4FqFF
OonWA7qTxWH6JlbzFmg/2k28u8ZaKgcSpe0bZwdq3DgQHfTeljaVGOthNiKgQJhHICkL9v5viDvR
g4UuA2PigNysCYHlSfktvxpuGAlS8eyFf4coErH5m0iqEBTIUmTyPYyv314aDd9oIsuQGjT7OfcU
EOwJy5oecpJeIbcyPyHqb5eWxLbyk84gZLDb2T/OwjGZTa4lDRtT6eCKPsIIT/cCv5r8/9tjmsLO
UjZA/URzAWar1ZGNXR2LqMiQqE5R4k6KXbU0NC4Nzqa9DYNmJMHczDoz4vQpJ6DdMIkVQ6GwxNGc
bFlsdtAifL7ls7TTutG+gczS8Z+Cf0Od0lbplTqJi48DCeqfSFsvi6LBZfNhQ4JK4g7jYstt5KBC
8QxcYySjQmN8aw2YRk9kcEqtea7nvNnktE8muh+0VKNTlzC+U0QBzzRa2m6Qafxuz+0inSMyV5/Y
Ci0wEjG73E5eO1JqVBrtF+zUIb6Uj5IeYtEQDNpLq4lqNZObwVcGL5ZLOSSpNemb+b/MBjM6/Ve1
1fPawaNqsfexS7qOheC8IDNdluylqwNfw15A8yIVtKCeaYfxO/jtSuTV9MriJ8ztEHucVG3A7IeA
GsffyFQWTBAsHzpp6LUoc8Y4W0N79grqckvm9N++z38IQAeUk8Oc7GXaZrg3CVQQaAvnkvO8LOYN
mcaJ282UmcZmeKGvufBInGo2KwAcU6+Zq1aOfuOKc2HsYFZTGx/YpGyY0RfBQZ27sal5/4X43kt/
09tiFkXOBayEHqwVob/18AfASMKIxZ3my3S09cRM2vDLb6v7+oWWC+ZU4XBr+FX/O6VDGb3GPF3P
Tua806hUtS8Bl0R4v1589pTekJUUUp7f3lPDy9nJYx8d/v+jyyFQ7v0DxIVCwFblCqtf4YrKvyJc
9ahGzUyXbCe0oBx7CTIhxt0aSU9VYAGfe7KyrIqc1x4U/p5PMhiezKNUlNwF2rMWCktDY5CMOuei
neGRDLGHwkLeYm56SHUCqO4usWcxQOklbhJ6Sj8I81YvzJBYJjaLgQHgbujsnbFJ3HcM66E90aRf
hVSQO+dDyuaBfF5bPKwADOlIvj4IU/JUfyxB6ns8PQ5/6aC1MVhMGTXfkEBQWCtoBBhql7A0aHNI
3p96DzKJ11G3oo5vkIQqswfqddykba9/LQz3Yj9xwK4dK7F88xiNDT9eaJHTnB0b3XjndLKznX9a
c6SIjhyLb0tfRlt6JBIaB2mkElZ1664SOxExxY1R8SiLBHNeG7NTFQ4r8yI8smsaDNZnQwdFj1um
hZt4pjhVekgsvr2wCH7DnXfwSgY3i4wGPmMv/MqMifs/soLHEXTmAaxLqc57UGb406Z3DwhiLsQ/
ytjFyaP0nTnv7NUbWOTTOx11VkEQB8jRgtzt/NdLXXaVJKO+gpBGjxhC+Js8dckMl8nP3+ZqAlbd
EAhjNlJ83HxQytAUSc8CW7P5sXIzHBHF3vjumXEulMf5/a3dd2Jr/5CuGP1PBvqRFZ2EU8AdPvnL
xzxLKM5pJagTS4B/m5hHP3kYp72UcVhPzWkt/yaJoOSm48HAmzITOZT9G76k0OkqLNmClL+S5Raj
Z1ZSLhYTTwrHyfFCHs5Z6qQrsfPURptB9hnBIZOU/cJghkT7GAGhuliKza0jnd2Grsq8SQNUKmaM
TfX12LLveXL5ECmHaTkEyWvkvDv8LAfQozhHL8xLHOB479C5ae6kEj/hFd+IDIFTSA27cletUGAv
LHBDhfTkNiSBry1QmedlmKvTWoFn21b5CvLgfoOZ/pOcGFLcJaUFruSvxyCodVUHWSu6p5Xnxjvx
Qyj308sRpixhBGlaxnOs5LHipHlr7mby7JSz+Kx3OthTcqbvXc3baxyyjR5ZCJGUVyTXOZX8NgB3
f443fD9OlM8IeiN7Q46GBrN0xD/2V3n3unBwWIO2JEhu/MeUvvDWKvdl1SimIHChc15laBAyPoZm
82JkAMun11rSpuDM/qqDXCjig4tYXfWlAMl8Iy4sBkgw+drlUcBK7SM18S6Rp6p7VG29a3SwebcC
cmqQzEC83Z6lZKu4istwoYn6gCLVVpf4t3RwbKxyY2U3EkaxwE9XXmibggS5UrJc2mSyFeFbQZ21
fVpvGpoMwKWDZtHbzrLYDT1EjXL40sQ2WaANlDcPZ7eZAwYf4+WxJhr1iEEtZfMHzlgx8OX/Pawl
gdTN7bPHQQaVAgS9o/VE/l502d1eYfYkZkNWiCEis5q0inO43XBM1ih/V+JX7F94ieg5VrEl6Avw
ukHeaAXfva8GYlwfGTECptUJCeJfWwRl8vVvf3gw+Uw+Rn4gpmm6Um2bMYCgSr/LWNIDs8sZ/Shc
lUUnr60mXRktAkBVxG2Dugam2OWFcVpEXUYQynEX/ng5h9NrY5TigqwED1PpVGksBabezSXXmqIb
0fXklhG1HjHD8o0VQITF9VfeQANX2FFN67L+Sz23AQRxFEcm/bdWllghOGtFu9/yCTd8VACBt9Ha
2JdBFv8zJcq3w/pRFL1G960xc3OZ5hWs6y5CrcjOpGHlTKmUUaXzKSp912OTvOLRerZBqw+Yx8MO
B/o6JaGuCVY365LC+kEU4LNObALGz/9r9MC3htURQoBf7vXpVWpvQfYFEBZNlZP7coV+EV7yUChA
G+KsDGy2VwLzNwRFXTZRypF3TFjYH2o0f1MDTY5ZEllq4ajShC4Dbi2c6h8BNwv6LBTjweri6ZDY
U0Qj6nKVLBk6PKqyjzksceRV0a61TliyFQTtglnfHNpUdNwJTSd1+UGPvOwyx6DLAwyyvKq7Ghx5
YWOifvPdvs61GHYUdvHrIbcXAQD5VZOFehddML4hhB58evHF14DUz6MkUz8T43gsCehEj0X+9zxJ
YdRbz1OM25jWfcXB1wNNs1HiRGKpk0txHGb1jItBwAGuES1seVkA/xReGkSmJNUimCIaSkMkGazm
LBHYSe8ZJ83A7PNUeHfhoimdIZd674ra1iFFrt3+DYq0z6GVi+qsbknLVmHTWoD9f7Zs54PizEN4
K6MB6jdV9JgjIqnzqKfbhyXm1xQL/mTDeYKzXyua1JXTnNFDA8ySKMKkjJAvs0pJKSXvnS03ylB0
B6F2m8J0kh3pSoWnbuRGWhQxIpZMAI2nLxmHEx+QbJKBy99iX+9r91H5kE7mQpT9TaCno0WRUR3v
bFBjOgNLyCHVkTgD4TQBpL0LxzWyrSc26vw9QI3pyAI0MZ+zwpAhE0I14RH+03x+9pzydYX5s8IP
k24zQQMijxS78s9AladlUZZDqG+5PI3mc6e3iAFQrAVvoD+/wZ1kR4NVzq5f3lZjVYKqtj+hqEH0
QTXtHnJ3dQrNT97jW2SYmn2/5CG7dv/UUKXdCtR/7QfuRYF6o1K+7Su83Msi4KB8HmYHI3PmLffJ
CwY4iuJ87ltu/vXbTkXe6+u4aWQu8XaQitPEhy5LuvYCOcM5hn0HJNdkduM3mI1pAL0rO/eEdEOl
vtoz0ioUa8Vtsfof7Qmxf/Gpc5PL+s1qzsbl6M9I27TSAW0XQ5eF6ibDeoGUHbAQ6zU74JGwdI5g
3I0CS8EtToDSAfgsk1jKEriDthcsm2i45kZhgDAgv/wy6QYljzDXCKhL8uN8CLY7N6ZPkmVTR1qK
Ehc3KRCAOLF8WkGR2G6K/75eQ5p3FdO4VPYLA2Gmxx1LvZFZ6uyzVuSaG0O/HLib5qaMGWxM/7L9
dR5ttphpNBIMdysJbsxym/Blwi8zILEGhNMLCDyIjUidU44qjQE0IpS/CtzM8de94dMndTSk7uJk
aZzuGcYj1IcHn4Jv2Su0nhCPcsK9mdOihLI8az2A0FDK7PjHU6cmzwa8V1nh/kek2Ldq+VZM3qfZ
DH+ebg6+DLSixtqf2YTYh/51YaT+AsUdcM86h7u/WBYKQzJsw2chb421d4PhvLiwDuk5yovKLm8l
6ySPM6QupsGmM74S5+zKXopqxH3JSA0xubY+ujYwq+MjoKnZgTVnBMBf8qI7DUOvXhrcD84Uhcfd
ugBsylKbyWyRs8R/qPrYq3y+gHQP4iZ3c3L5SJ82LxiAKDlSZY/Qu7HBt5PsQhYTtvsvX3WP20Ea
y7bc6o4WnTYvExdifbnRDhXvQRer7iw3D3keHsk9cpaoEeN3XPYBLJENaX5WKH9NmLYHaJN+zdDx
9iNrDcQy0hgyg9nJed+o7rjt22YFBLZr9UN+PVFtWumsqpc8HIt/jFtqTQbIRnQ1yh18/b3/lwir
EgDND4KnBB5VRRG83XkKQRSspM94Jwj1WccRHKKqinE9o7AUSNQ38VenUvt7MU8QOq9wFiWc2eAv
TrL2IXsl20DwWUNUrt6//VqVwErXCPqkGxltHkEnvSAnezv5WjcsHFspkG0j2JxTqFH30/gxiQrL
/+pbT1B4OXmvtifRCubxlhbbTiNlGUUmA/x1MxqmYBb8aAzgaaqwMgxsnnmtk6hkluS7yzZA7L3R
fm7ZMBExadZkYzWKW4bJhAJ2VfknnecAfYDVUISq8Ey8SVY4k9NJMquDnWGHj1EAbYoiUD5wHkNw
c/WDznrEK9PmRvcM80g7DbaNehRfVo6Me07Ne7USg7laIuoWhJNhFIpNUsUOrSY0GUYc0YyyWui4
7xXxe+uuIHb123/yVAs6Ua82iUNbRtElRkFlKtSgsoFE9v5B97M6+68cBfbD0qM5GsrVxhA2QN/P
Y3C+xAikV+sAvR13EZxeVY6TgqIINJEsY8l1mBy9EKwFlyz7FoHCO2dnz1g2k5ijxi7iz+lZP/xX
BL++gwxMiVZkLrpqrXhH0LnCP3Ik18yozc8IzrcZ4/nNPc25iaCAiByISUONeGQLiWckT1oa5W/1
G5nyaJOcOsEV/h6ug/OD3f8qfbw0ygDiddS2LVKCo24jlw9QjOdf4DxkscS4nLRGgPQwuEdcLOyo
pdDRGEJUiFMBrFGwT4C+STcbj9VKXiIQLGN/Qe0milBHBsSH6DONADflsuwzzTRKFNWRM6+sC9/1
1OxI1nCWNFY4rGbJdtaAGDGRgPEcLzklS55CoZoIHwLX3rblFnreSJyjKLUAbEMI8vwqZkdwuudp
yX1lVIfEaXxMNXlzYuqiAldkppYJ0R6Cco3WAtseNGmUITasbsF9sIIsG1F/P0cGMDBrtqFDQ5nn
ljsnN3QE3yiOuLr5EwUkwotFaRNK43LCRHjCUnSP9RGKgRebZdgHE4bwb/YSMfZYWcJUa4T4zOSk
GUwu56D6Wr4g8AWxGmlBo40hrNvPFa1hIBql8sziqDa1b0ivjqWnENn+nOsRES0aqdFj4ua1h5+N
1Qr8G/jluaM+u2MtZD1LDaIXReJaYTzE+77BiWfHVKyDojA5wGseYBlTSl2UAtWcpG7Tuj2upv9u
1FbhsuQa3HVSXN9XFoVqfLsqlCDTvBAlddV4CE/4Rk1kUg2eybhrJ3mM8dMA+zdOad1xTZhFyXgW
A/iCqfnzFK5JW8ye/YbkuXBkcg3I2XXM9AoH99HIJJdkdR2R9ZZm9tkEtVRKeWrippogpPNuMrUL
T87hEyAn8jSD2XC1yNkro//lX0gSGhheGHVDiNxNCa4ONBhc2TGzVHJtDqM1ogIPzWXIorqPqu12
Gx6TxAaaKJrzUtZyrCa0ydi/eVaWOvuH1Dn5HgJZU5x1ow4DN30n4JHAvSVZMJlwdfBCyRTICdFw
lClk9JVJfH6IlX2ST39jV0fuLKmhviBCZASDzsQVHTIJxomjveYnzfoBUuD51Z9RWEuNo0mNuJ/8
l6WL1/k090lOLQINkQIym6hvKUGGY+MFwTGdJQRNsrXXs2tR0FTnvTrTCS/R2wX6HZFux0ttLhv8
eLw17juswj0DD/hs2hbIwU972JeUWsWoXAJv823Vtu1AG3xsvpjw3nlHk2+sJDAnzL7oR6XRpb6i
/2tz9p8mC2pKWD+7qsIlY4liPgWroI4/8YULZvCf6ws/T78jiqmsTnVyGofoKfaZirievdwwDrgv
RnCSpjCbZa7XpKyGdnUuI8MSTwU9+23CrprQBfbc2lPrBDUDsVyDLt9VQRKvyRSs05uRU/vmhGj3
yLWJWC38mxCjc3+u82DfmxxqiqvagH8nJxjQA/UlKhXdlFMq/OHwFZvZ+F/rD0OyYpkGmqSiQ5p3
9uAs1GIH4qe1loNdxllTFNY7Gtf75nwOgwQCSWYid6nKW7vM6oVqMrg7NaOlMh8qcO4XrM5LvEyZ
UxT0gE6nToFDKK+6jiB3cJ2kNahPGAJptRs8bT4TVcsb61RyErutLNIzOTw3ff40cufNIdV5ZrM6
p5EFi6EmL4hrr07vDlWW0zaMn64zuoqIjPXMfJCvoTk05O/aP3Y/z+MiGnpnOVl2F2GAN517zUbi
ZGTfeYmlVfj+ZfzpaLCtlq9rlompk6yWc7tBQDF5+98ys9Zn9s2f9hvtaawsN2QBaRXE4nVu+BGa
hJeSA1NkrvNIFLESQhG4n6GJkJ8eOMr/iUpAyDmPRMyIUsIQGf5XBt/7qwwfGmG8aQskdQSh3Q7D
fw5ipfGSrcW0+/vjM9jqfs3xaVPBCNyhd95LkwmrYrDgneneGJQZE1QOe1ArPyhcJkcZgEmtLVgl
Rv2iOyphJumfk0Ppr/m+FVP5zwrHOUjB2ZqCFsHGEmXObrElR9Hv2WxpagxOR8FuzZY08KtbODAL
46Sw1KlHsKhJPxO9W+1Z6pFWWFrIic3surFQheLtwvFlhdpuwfASTmmoFP0vuUbaZiz/NPLUQALg
/JSIK6bJyu2T1HuNiDNL0Z3zNcafcfv3HHFFS3GslppaKyat9C9aGylIZwKTQmJNSzyr09NWycwQ
yzc/XSPxiaDeOZkocmdvCUVNlvc6sTUgtrCS84BfZvqZP/aXfWcCAWF2X/C+JzEwSMUxfC8WFvT1
fkxfH5JoYRbR/63Dy5HtAgELbMRI+GxlRVml3GU6mFz1h82rdDT8NETrI12Hd97NUMw/jdFhHCp4
ZRLG18QhG+0/u0rRJbJZFV6+iWDxCjqqauTP7JaXYzhaCNPHXYtpI2XUkCmZ4BVheLIqbuTYiGAc
lO4nsFzkjfK4COsFi7Uws/iEEJF31YIm9pwN8mBhhOvBF6fGmi9POOFx9N/a3TrSmmTeDkSoxcyE
HpQ4BsmvQL8UvRoYOoumphrmFnJGMDtbTzsmIEudGUeXSUh6jmAWSw0CCubUomkb+B+ZH71r3xk2
ncSUPwkuBjMyTYJ1dG5r4Ao7S4R80RsIAvNSLJEhG5Riy3J3pnBPA5ZGd5ZK6JPbwyYe960T/A/T
G03R4I3iXADxJasp9RVhZgHy5Tv7l2trHfZANBki98SBeXBsfTUHBYSRFsCZdv0mLfVZlzlfSYNF
Y1mcXJy8kUuLDltKwkL+DX1elqOMYOgnIlzD2+gXXUZDWo5NG0oZUxe8FSd/zDg2gcN7K2ddMnWb
QpypXvCu3vfnwMD/WQG2TjmCChw6eGYVvJWxzFhX6nFRSUVp568TEoz69eiAYouy8dFnGfLMD7sD
za/zOdRouxjOMq3MTdPP0vI+xKRwTpMZaS6WUnJgs/ohWUKqRutQbwwIuRYgz47GjhOrcpnZvaOo
Ld5KqilLq/pjpjzl/ipG004LW/cDZBKOJ3MUNbjmCqEF4HiNl4NT920U0RNT37425XP6ORMuqnRf
hXHTU2ngRwzzql8e4JQ/0A7YJQzYIjeWqJLes89GHQs2uiJOUQe0DozyqSBNJxfylpvdb7Gr6u2t
mwKsNe+Mn1BVGN/jGaSHRF4gFydzapHTE+H2TRdK4yTmydaEfEvWUqJmJmlIcdWmaejpAT/uXtq5
cfObs0O4iI9j51o/KMBKyUYnlavAxg78qLtI/4gzd8gNbs2uejKHUg4MOh5A7VLDfdkHtssHh3WE
DQ28n0QqWeiODJ1zPTEStNG+fRV82HnNcEK/zwe5B5Umgs+h+ATxyBhOeEWytubXBJdhMQd28trq
QVJ9vwNJr9i8Pggtibb2YaYsCSq88ElY5MbyVRP34reTDIWxIaZM9ayD0+YFFGA8Ygi4rAYv0CB9
TvWRjzARpEGYQ9ff9rZg6MjknMWkRoa4jEX6Mns29YrkNOR0o/t9d5m7EbIttCABcIRW9gWc8Aw2
lqlrVyTLIP0sWAIROLebTJAMFk+NhqmrDX5EgeG1Y/Sb6mx0PdYJQJ2oM0j+fv8IfUML3HQEUCqa
/vV5lwK75mOuxCJNjn69flwXbDwmEfaz0AepgYwx+KADngYhG1ifQbUjbZ3ay/4MuamrskiX4G7Z
/Zo4oUNpHGTQuSRbNeHIVFzo6C1hvHLluBQv8eOREt+BAN8XJUzRhXmZY9tYfZO7TB+zjBRmsbo3
Nh54JaKXgEQRLtY8wV+rHHu4I9GdpyWcWZqgezhfb7VPXqOTjxz0kkqSagM7ZC0O+u3nI1cEyexB
YQkWZRRFBLBRcxpFqw6i49vJ1lWip6kvTlborNKQUGJ/DjUCqexLwq7oaGk0ZsQr8LC412m0nGxh
ngySuvdVRb8Gr+NC+U9QRLRdkKlWdA+7M53EFiAaxGf8f+z8y4lbG3AzfwMgIwDIW6a/EQcumyiy
yhh0smg8rzACh4CWpjTpg7RY9lGtjitrM9uUZAPK/agQ5Dzqi4u5XFB7ujtQzPhIDdoUt88WKKVX
OEsvYAZP6pacLCFdL9/gn2FUZYMPWVLWiE/YFYwR1Ie471DxOuvSuvlq/YTR4u1sCx0eA+fzdURX
kYI3y3LcPGzt5rtzwGojWsx0Fo9kxmrdGJzb6hWR/xeut6CK2gkxFXqOtd3/XberZe+PBKwzmJer
5Ikx+n3u6Ba0LAOgpetsEKx3T4bsW2pdaLheT08aI8Eg7C8CoIE/XVRI7qMOIrxtRtkp5ax3Cs8s
127TTUL8UI12qb5V2MkorwSkZuLlVIcvGlxZzcefFBcLacBexffvRHfOC2ihWnW2u/RyHFiM36rD
X3y0mi2HAKR1BxYdq2lenIcH/P3/ZytF1RXJIK38dxVS2lS4DNq5kODtzw0MCuWHG/kkCHasnaWS
7LbGfBvhaedf5Z2ucmGw9C9Gq7aeUZ/vs+gT/l9M4nadrU/mmq+N1QWhQsRZV8S57TigVofb0nPb
WdUWSWHUvL5PjVW4SyPFtXR8wfKN+/HBqs64HEi086ZoB7QY4O23WGgXRgUhOpCLsT11MzjqF8Xw
HeYnE53KHkNcySiy0r8fsjEyr58Jk/gjnsb4CYgI8WYLbRMTPwhRdoniv1G+zemR1466NxASkzPM
aNIJncQyO9wvW/frkwpr4MJUvpjWKlZHUJYIGj2TivySjGVVdnfs4+K6Y0Sr+bGEBOvzWMRhj8Fv
vCg6jDVLktpcfocJ2PbdAC4Df+Z96tmZ6d2skvNa73BXozNKuBecTOCPwaWGgoyTVQxIJ1j961cz
q/ZTQ+CtPQvNX1bESiG4RKD+3t+Ch7XM59v1VFRQeGvUUUZcp3MjwyIFhhcSQ9xdc2gCciZU3RyG
fBzH/IGABEZf5u+znYfRh6nlHanmSJDr+emdaNWDqMhanTTPVMm7CnnnaN0j/EHNr8WD36C+ByZ8
LhVa/86HKCV/peoHlpwOKiGWfU4dgC7sITFpX2jK+kxuVl8AAZ6lKcvTt0p34nfKNqLIvrMvCa64
oO/B/QSNyLIyYq+TtYnKCES671P9CCI0OI4jnEOr3eVXFk+LdRLBtdZoGsdyYh3Y/wihfT2KX4T4
zcUh28Up5/EcjzwPGTZOXjWfh+NeQq2m9QYwjuvf8+HYPRuoPxKQotK8/kOdSAZ0Ygxpugy04ZkO
CXP9Ilbxy4ehxoLsAT7aHgC72Hng7Cf8voCdY0STcUxW2VMsAO9bizd8Ej+IuAVGdM3k0v9kbhqm
1soILDS/BQ9ChEeRwm8ed1RUSF6mHkjt2VjdvgacOWeQnhReeoSgjemHlD/rNySWN5555FWaGZab
Ixq5h42B/DLNyOA21M/An9hWUpSSBX38dF81rpuePY1aQgHHnCysGkZA+xCJJhnNC0rODt3KRqXl
ee1REJUy0VWrk3eNlZcG/2t77q7UL6ZUpJvc+OPP5BgyS012NMvtZvMnLa4RxsMUggeo8wYPEZ8t
EIpwDKotLnrZotL+rt292BhH54fH2XVYrfpueE4Ypxh5+m/5+R7MRgdjmb6QhN4bMHJcQe4KCXes
0aLG0dzrqxeP/ohB0xBz1wmqcxlXYDpw1K8WoOWl8ccLlYfwxWdvrM16SfC/KZPbS2zCXNKhX/3O
fDfuSlyht4G5uhmn6bltj1Iqy4YICrroGtOrLeHJEmG2fUnT1zr1itlnAnGIZ4N9MAoP7cEKyFr/
ndVOOfIjnjVFjkIpiV8v2FEDTk4q+KspWM3WiP9FIZmTqESeUboE8pTpsKovF2SVKY6ZqAi2sseD
P75BziM+cuWY1mRa2rw3r65tKxHPATgAf9l69eeoVYZdNdzdeRrOFuuu8eTYudyzMb5BJ+PWELuW
GyaPPIxB9sMmUOHFPoXOEIPnRw8jAtupeOHCjWETVWn4xNFd6i7jP5REF+818cFo7s9i1BQO1es7
ya9OKAopc4Y0MyTSlgFNNCQK38UcI7Ol0wfTz/TGykmzFTSE7ri5aRDw3eJAgj/06wNrIqnXdIGE
/6OxmBHcOs+6xTHndlRdZv8jSbLPTpkI2HJWQjmyHR/VkUvtiKwXF7Lf23/cfcuPdvaTtpLYb25n
hqykFC7wSzfK6zBzVDVC0HGLkjcJrORtibEftHDoZpTlpp+v5o75WWcpmT1L59cg4+mBZN0UV/Cs
l3Q7C98j4vyAOhA7t/qVKGuzMTXKCEmb7ZCUlJucG+SxgZu4byT9sacpkt7d+zK+PvUR5CDcUG65
jDw3A0BkN6jwUt1plzZ3jc1IEKzx7010/XToN8j0qkSvoy18WtSv25zWP+PbpHVFmVJjubN2Tav7
kSqOFVlDLK4/maXBsZKpn3kHNTQf6PYMYtTOokfE2mTI/XbpjGohBytC6zKeNTirOr1O9d1wEMcI
JifyqpUVX76Eml6sopfVcw0a/4Gnv9YQ5j4XJvdi0NvC2PZR7pB0OCSYu5sy9Xbtw66R7qqaNOYF
zix5bc2J6xyGHn2Xjwzjf3gLZaNU9KpyXUc2ugE0Ii6aJv/BXo9YjKeTtrEOd8aqsMx/5o/bZBfv
zUYmvoSmKk7sq/9W7zST4wWyldfuzlYbK07sPc+clh803lY+x+ph8tNqsxoBH5/yBaWoytx/w09s
9dU5ujr8ZmvH5x3OIyY9zvsHwQxpm0xddLHPP/EanumUCZZ/awVh7TV1i3i3Xd0I5Rm+i9f2ulJK
JB/HXVxgtyBG8KQV7DnrjbsknToRCRDdiprQxQpXEZ0ljBVj+4dH1/bYpTvQBR09mP+MBax6EdoP
PaQ5pCT/LacnNjQv8scRovRBUVkEJ7IF0qDjOPAjYaObBhqLWdDP0Z58cIJTKg9afKca7MfuupTq
bNpnsRLVzodwa3yaLyjgmpiq5rAcnrt6PRqcwyXP7ZbUhLmzQ7SYEsa4qfb5VBusUSJPHQJMkEBx
HohlLYwf1LI3p+KHPidrdTusEz8jPM6qeZrI71bb2Vl5QaVCPE0YiP9DFmXN7slgZAigYLIBV+RG
NityjWfY+D3NX1eeboamnf2hsm1MTI2QUZeHcXDcBrMf6p+sTQlcJ6JgmBkJa2B9U3v587ZGo8Qv
yK23J3bwGH5zU/RJvmcHInftPp39774pO1mbe9JRr/mxyCaBtR63X6XFimPxtcfUnlA5xiYTzAly
582cp9yA7l/2UHiAMTEu0URLR8WuY1bxWOkXB+I6WJ/TSUt8QhQoNjTPxRp2F98hcjjF/0XNzdil
USCfNyLijkMeC3J15iM8eU4zRPe3NFjz+OOhEiePJFQS/oCjwR5o5OwjruA+To8KCtmQGqarm7ut
1ne0ygZ3MykGp3BehsBoLlHsO+jW/05OUzEVQSuJ70DYo7q++5qUEbdEQrjxwtvCy4QGca/loTlL
qnCyn31H9QAB7Y7i/v9VmDx97fx4gCAk9sZhBDhv2QuNoEdoez8NSDiCVXos47fN9bV5oasjVUMQ
wYuIvGwFdkiUDQIUQf/hOpN88bAd/iBTlw2W39ihh/dkygiT8T2PCTKonVPcu509K/+EKTAk9xlm
mgexNE/MJ2FXLz2OJFXB4bNYACGX+CTx4Y+MAOsa/eJjCPRw0Y6HT2yLbckrUK82NAU0tMGhSNwK
DJS8DVWjzyaO+VOOuyeRWeSXQks4SzRkByQin1mFCx9wulo9v6xXTm+qTB/WPrsL2i4j+nf6AuCv
R13VPmaYzjNiDRF3Y4k/I6H+H/VxHi+8BRocyN8PTfsoLi2/1AVd5ru7ABa8ztu9P8AY7WFJnbeB
gWxJ6xXRvgMrpEifQANk6ObUYLBcgQxsdVV4CmNTnMCU+LBCg4fXqh8y+JTR6MbP3Na8M1Bb1Wvo
sb6nTvXQ+I73tzQcRp3s5dDsywIncH2aIoYVr9ID83fPp7HlX9RvlGnAgciyhlGSd48zp/jv3lYj
8D1HJwlONntM01wc8EH4Ef2QQpzR7Y9Kau2eKRSQ8MlkJG8NndgYO44/QyqMzveGnReVmQfMJn5b
TB9rUtS2PaFkwIsU4leWe9QGNaTGrXAr2uCNjxLMSk0J2+0pbkZWyGUn0fFXMic7kjdIU0Pi6XhB
cb2H+cXIqFrOu8OVZ4Ram4qp66rnpkblK9tR3t6AjLUUoJdq+uQPMshLh61s93a5cdf80RzpaRe4
66r+CvDiHR5T0PJSrAAtn44O4Qi0S3bKxkt5PPjchC5GozoRwV5blh3l2i6W5sztcPAjmxSWuO1I
ttGtQhYn40Slelf5CG5D/KAQdMvhA5ArCNnnEspGEMrOR0OQ52psEz9iRMeuMZohOK7wQPyBDJLZ
F0XECoz3CtVH4k3XcfMqyCVpFJLVBpK76VHoKNJ1ev439zGSn/Tu0RPwsMji7+gFjn1u+Na6jEUy
eNUzNz4fNA+DzKn2UeRY3RJYWZzNF9L5c1v6NFfRIEL69aHf+3BWmRwFyRZBfG443auR/eKkksB+
xWJ0YdTT3Le3W1Dr1xlJHBEN0WcpJpV+c7JT1MXkthkvj8D7MTmoEXEEVhG34lw0yeHd6dC1ZFVD
Fn2cDmB6e6xP4W8wyxsQ9FWFlto+HZlLR3V4P7P3UleSfx0X9GI0BsSNAl1x/aA5MGy6Ig9ct3JQ
diTswDXjcg9dr9Ff62AR32hdGfKgVlFwJlQnysKdkrWDhVXbuMktih2gWTTeVXERAZoUrq5cVAK0
pk9hZ2JF+Ri9KcYpFUVoUWGt8vw90yKcUq9gqcdScdNC2aOcjzI01Sg1vSIrmB4haEwYrsrY9Ijy
GeUUJQ9LqaSSlO7ETKNCYJVINDI4SYvlrBuEhKXhP8tGeSiD3an7xi9uniNSJ7t/X4oA+7wakG+L
m5gM+Nkms33ELXUJtGyQzTIFtxDUSwNCd2AWk+EbyZatkCk7iy4xT4wb9YlBXf3m+OPgMCUPprrc
QRxintsLR4M6wL/HxK0NH6CLrlGZ01YR/spStS/IFL/X2ZPJNFSqnLiZSIavHIUUUur7k+e5qhtz
kaYQASeO9NusuuWSMI3wplGOOYMQmT385AV9ht9TE3a8bgiprPn0R2rcWeaNqh44hZxcq16hiRSE
8YvMlJj70rA4Zv6MhcSkLB2UBRoMyWoUJyKUYP/9IsNESjHeKJVVsGeHijUMLoEomFiX7hphTH0J
dC+TJ66q7ad/x5/fxGBJ9gKOJrAGL3ebrpL5bp0o8WgZqyZ3XNVvZO1ZQWm0Uy0bAguDM6MIpQKd
YOGFSVaaLA9zmD5NLyh1WYC4QJMf4iZFG4GJ7bysTGFXXdF662zbMDb4wi0gXG62RfKzhDi5MSP3
X1gNu0abT4P1GgXY82aS/dW1doXRgRBgsru1xZW8bWsvHoDDnbDS1BvNkWIkMdj/UmQl9xiP0gPK
bB1A4W3EnuRN/Lqul/++KH1Pslkw+I0AAqaxWRPyDc4v9JLe46BQjQ2BB3WyyTEpBT5QI9fmjBJg
3StUhYw2Kn1R9/qvNnP+xTaqJ8JMcBmdnvyCO6XOYmoD0hiRC0FRU7iYSzTlVKy1MI712BBrQt4Z
gGdxQV2wQf2Ime3y37JePinIi585X7vBNzJZwiyu3eP+SYRbrrOopC4TaEls40QGp+trKB6F4vFR
1aYYnwFSBdRKQTl61L6t481DF4nMZkqBaVh0eC4gt1BuvO8Q5Z7HzbttEAfxgTx2YiL0bqAzbY/y
qyO2QHNMbFIBJ05DxImkMujxVwhA5DstfUvBws41mI6HP9fdX42d462Is/nWWnhEGuVejecas/HF
D0Jcn64nB9T9BsBEtmb/4zU1zANATjyjQk561Ifs/CwXox1NhUTL+FnhsxyYB49KohtN1QWe06jq
QpDO9h8rECuq2aHfwkyGtHB0gNW/1AXH3ezJihpIOqMSsB6MRs3BfTjjJPOXOI+NVyQ+TBc0Fb3V
kS1n8XRj+om9MXmFsJVyQpGw1Nx2iihfFmvMORXkw8Oi/V+LtCBCVEboFJyD84U1LU3iOYohVcza
8NCEVkCxBfhvhaRa2CONavhdLiJTetz7IOxolvhJ+qsf/zmNGg7qdYWF5Sz8Kf586SV4izTuPOzB
1oeqvSJCVbqce2m76E1q9K/kYmLD3CZ1KU+sZRJHts6MZGGIbMvxtJAovELCCbSSEVNW3kg8S7+a
25UujxHjLXaGBnaTYCmoygAUNYhqcYqMqd4c3G1YaTCdOIfZ9Z7oEQ7ezuO1me1yp4SpRyACFQrF
fGKNlXpTnBd6xqGK+oqoeDzkKgP3vve9tkWEvB6PacZhobzvKniXnviqdaeT37rNDcgec7tLFBtS
sNdJ4S7/60ppU8f3gqmYR/DRcQIByDquuoIlpMvCeieNeN8zkFFstH5Q3vEiAyOU1Wr5eTghW5O1
QPHM6sjJMM1lsp19rRqStxKJXHNPWvmwH9vgNqW+pDM27uZmrt7OAx0B5/xEifkzJiT4Vu76zPff
4UtAPGwRjLlOAIOh37yqibiNs4yCppuY6Bha92QfeEkRqdd6VWEIK7YORa198J5fP/Dp3FmU6z6X
OIJu6PeZz0vU2lF4BA/f5F9JvMo1xxxwSsnqXw3YQu1bqE8mBXOGU7n7YHp/qrBdzOlU4oKzx2cy
CzHjaWbFBEtXngP59oTvaVDDf/HLPjFK41NCXG9K1w/HZOzOhvQViUn9Emc0ToRSIdKJRFOmyA4n
fzPtPimOGIZsWrQ7DWPL6+mPziPuYFQ0kMxyH9HWX63n0gMtuqdhUF1vz2PfcMgG8/d2OuHXC7ma
V7308WKxa8OdnJuwQx8VE+6jYtmWa43oI7bxRR2WvC2QQo3ez++9D3VqHcot6riJC8DU+0Lp11Sg
MxGN5xwqxa58oYzr/0GWBm1GnEI3FTjbhgdR80BElF5mU0FitbKkK5SZhLlv9H1hJEFb7giVx11u
twsUVB7VU11xk3+hk1OFBRgUia2733U7ZL1YRMDfunRamelQE+j/TvTtUrXMgLDPMQGMQ2YIW+XH
/XkrlcydehwHpLIJQMfXFFvQvdmyoRIJtRSkfs4Z6LjAONeKbRjxv3IalcNG95lvFmnhAU+ku/bB
aVNM/9RKRJndx6e4Kg3mjDv+5vewCLs/2B9PfOD/yotMv/aSHiBVRCVZlEuyb/TU8pkCUbN0KmjH
kHW7Kq86RJc7VIBvrUUp5kcHGpebqwFaIDgH7XKrsRWF9yWdNc7xcOVfQmxeR3DSAdbavE2jEmLJ
JeeaDi4DQizsqrQ7GkatNfMEHWx3xAiu9jy2rbGOtXRHFnBwS5kMdK5yYS6OaftjLXJCboNLRqBq
TSKkyU9xZ/UU1eck8PbkvpAvIy8qD77Rs1xS+lOtzyMFhU+7lCx+Wfmv0dDs+yr3M0Dhii+Kg4MR
Gdwf4wcnYdrT53jHVaoOOs7yQyegrGJjdRILEUY+7Dq/AsoWPOEgKQwlUtOP7lyrhfh5qfrRnw1S
yeKsESC9B8or+HF/sdk+eCq8noQKizP1d4woWbsSyNPNVmU3AfENi2KTdxaIJr8QdjC8x/UVHsb1
S6a1Vo9wgMy07ve3pJbBjSTTfiYzTeTtKsegDdAfzIEmKTALXEtapz8fzBrPdhivSoVM7O9IIwfN
VaVo7WVvZ3BHC99BlxMc/WaFH2NBnVQbe4AExBLTXT/HMriGaolSLM3EnKWCmPoc3perpsdQAXj8
38y+DI78fQZyNEfgwV3gb/29vot/4iQjo3GUVOeQvjim3GQTAiXXfsN+1ME5HJcnsZrajNb3VZHO
VwyMSz1/rX7EDDy7Ya4xakWx5JH59M/kIezHKqM6EvCZeZDZcq3uqDLu8Y8RJ/ZhKJe0X4pX8GHr
g36Iml9zbKzU9gmqBC/Ha78sjOm0G26jD1xEf5Db1GZExvVwa/c/W0a3g4IYdiSo0ZXZ+u0hDCH/
LGz+csZiUrQ72tw6pKBco8qWxle/r76rNETpGFO6Q8vsO6FQ9Y6eLTws2i4UvB4qQ0j5ArkkETo2
+3Ewsbf8EaXAEnkqSUUoHOXSqPZ093iYKBJdkB/XGhdfymaBpSbXuqizyn3hbO4ACPrjRt7p/tRS
EcgIUn2ZBpCkCUj9vMIoAbSOJBxBi1qK9MHOD4XvwMmDf86+92E5GPKr1XQ4mpWO2xHMowMlm2To
cKPjsEUifjzzc1eOHnJmylcgDx/EBvFOC7/y+tzvrH0XQthY0Y+8exM5ts0JcGgGPHt6/EEfilG+
SOcvFFHRsUgWdXghap7ok4PHLXufTDt/JXQmTXcergWcFATjyiAjw8e4Wv9y9xiac0UUavhHwVzc
bHDkRzRnYr0HVgF1ykFi1wG4LM6NGlB6HQRg95iPulw876mk9ZRBizmv5kclxuo/kYhGCyDjETUz
YDuvlueD6XcZtSfPyilDY6fuoJYZgS6UhUHm/UaTfRqKbA1s5qXRyADES55buWnMsiBWSmtXKJnv
sHHSRGsjo/i5ZsnVjI4l3JV97H28n1u5wde5r7b8Gu6Oq2E1aOTpF+Bt4agbQErLD7PJyOrdMaHe
dVXItNnZ4XHbWl67KsMX3KrHbkn9WyiWaqOY5UmZkUwyL/UyemjFhNoRky+qNtMxna0IQ4i/1sCf
2jWrUdgsCls3HhIlx0LPWiKVvf+Wphoit+A0bezhJRRNAgV9w3piZkk6G9Gpug1CEESj5d9G5AP3
l7N1t6vEzcpOaq9Wck+srr4/jbH5JPzvoGg1I7gmyJrVbYdFl20heOWC4b/gH6EQRmUUY5jXn36Q
HxUVtna2Kel/6Ewmhu97m8lpW0U5RVqzv23D4ihG81ZwJdSU2YKD33dckERGI4ob+nY8aQR3U16F
kdanTUhDqzILpIp0KCx8jspJTjxake4Ytn21uGYPQGbbcN52gh0kbjj6dRkS6evo2mviYWkKEnOl
MHEYb2kxHsownVjRtIye/0doZCNoPZHz6N9FIFYO/X2UMH5jwaTngGjmEt3uYhqqgoqAfLts3whx
wZRPk9iVx1psdWoBgjs0/c1+MJatcT8iOKbH/Ke57vHj0nKD6fWCmLEKOe4jo9Jojp2AGvPJOyQY
iOe2eRFPNSv3MFMBHvgIoY/JoSE6Y0np0FLs0Ib8Qgz0y7LFcWV1Zjblxl5FKvI/uv7JvuF8bpBJ
0j4rzdUzJexx6fdZ6SAkMSFpIsUQNby+FC59eT7b8qTDrllpCznLH0Xyn+HoxFWedSSCSF9uYrOm
GCZwfdd/M/cre1AY8lt9de5MhRtkalWkPrbqkhv/deT+tQW9mjeSNg6kgIHjlAPynu7VxoFXHGXi
HxPsW4iu1kzhfKZNq1tC/yFiHa5HjnPGkpqJttnpAqqM3ohltdW9CQ6s6ZiaKSX2W+L2EWl57ODJ
ksbjQkwPQ7SLBCJ8lftxaEImLxEqh46AP6WoaGDsJ7jCwMbUc2/isP67yvqt9ZlMlQDGiEd/WN2B
hNtGsgV48FZGlHojPMd71PtJdNNG1f39scHRlnKo2kVmYC5yg0w4oJpXE4AYcTjsEOTXAUjIv1ju
0TEUUlL26XaDp+CLI+xTif/d2NqGmiWAL4ZKF0jUQrDryiiesNoJH4ZZywyQ8qcX4HxDMf7yYMQc
lrd5nPIOH+NGI3Ad3U577SwrrHhT4CG+ujl5a3WLSHp1RfCjEH5ZFasWY6j/gkxQnLyygL81Mqtl
iv/XIK74dezcpjnRhVFw1FxGfi3bOr0ZpQ22qmINMYSdsGBDTwyQZ2xvSDpZRTypJo1Q8MU8UxeD
pMk267wvLkSYlm4FDsAGPk4c/r2y5wcDGvMoa3X0ytlEZhjGIEeqfOaBtGrUs3ihZF0q3DWUtY1X
fNXGvgG1QyapWCD0rCCba2015jYoHQ+2Pg3kqsMKL2AyyuQYFncW5RjYR4lfKVQEM0/v34y98kot
OverYuxpY5p7wti6uQtcv1ItU1HWzZ2opD9HvZ8W9yGo2FD0tNwuu/PVLvAgTruwM4NYn6C0/Pkh
abyNicWD/mlPexszxM/mxO/1R8kOdTLkT+ce/53vleyVfyIM4Rtbtnx9WE3ZIJzXHcuO5vKKhusw
d+aHXJ6AFNBHS57OL+XfIiMAIh3iWiB9vnAe4Fm2M2nsMWrv1qESqxlSmcjEOmvJp6TlATWjc0R6
FlAJgXtEaPkpvEtA43Cqln+mXfCXhzK5Zrzi5zv1dQ8dNzRz2wBFYJQ74wj0Jj5ooX8thgk2Cw5x
RqcKIgFZmLfH1h83BxuNM4kBFEKlfc2q6HLuosE1qFFnCn2K8Du1N6doE8QcLJoDp4cPGXZATKlf
KdV2DQYg88MAwqGQSOzUATSWxg24i9Bc+logfNgb8zSrZenrmgVejMGzCSdtp2+18HpPXIB6oSxP
Ub9OVeB/ktdVR/kgR4cG4DH0wObxSoZVK1IWgUH9ZC4N097pkaPg0f+GFLPMYSgN5N/9aHH1kSld
lEFyqcbenIyiNZLCOjER8Y3Oij+pG6q4EJGLXT+icRkLiTyQ+W4cCpiMpvk/jHmoqQaUB6InAyjN
bkepxAN1z6GkIdxorzWehddYhUtKZ0CKPLTw2aktNUEqbr6f6qAJ3K094ixsGgbesyCBl1JdFc4K
/hvI5L9u3QUC20AtLwDiEroEwTVr9J1WMkxxHb7VwX6p6LKsR8I0JWDrXMNLCovHTT4XPIO5/4z/
hyFgyzRguDMuUZ5nzokm7lBZosyM8F9MpuToZNPp4yJ9CvqVcLnaggzvldipr86qBDn7aiQP3wCG
iRc16fqVdj3CogDQGlIHtxxGifwflhi9ew347nk2g4ynIRtBF5Q4d8uE0oW2rbMBb9rDp76j0o92
jT5hTCH7KXsKeCuyG9CMHmHEgw29ddBHlG31/cwFEitzgjiw20jFxLEoCouoiczltRDR+gwlT0M7
hQvJ/1qEpD65+im0fqCwz3/POREJEUAe6RionfBBN0NDjlZW3ekHzSpi9NUrvCLGNMLOJWmyhZH0
05fEz3/7fe3QtolFlWxkLLDAElOq174aAxNGmChaDBtkQCUUfIq4scK3Sbk4gav7q1i7sNS84m8f
yLvlgKhxkor2P4ywybiZ+hJvmkRZXOYnYfZyyTZYAiIJSC/omxnckovrvs6Q3tPoYhKzru8owHjE
JTEHA+rf8kphTTkwD9+e8VrpsZXPukvvll4DrpL8PCf5+pIMWjdmmlzoz8antW5hFfv/UFHN0efi
9Mb4T/X7vmwXvqHxSQntynqCQ7VwVjaIa3dkrCxKS9JDa4oPkvQ+r7KWnggd6j7Mqtg5QAWCOc9u
0l2OOIHw6RBPiZ2HsqOwWL+91wWYWFVuGMsUexPC00IntQh1nS5WLsVrt3MXYFsrDmu1whyUKjhv
h2Fcj8Ld71W04eOOOLW8mRyf47fHshiRrHTyD4zGqu7i4ncTEA58i0Kf430YY+TWbeFh3QctxogS
QSrzc+EA8pwczp/y8o/NeyuzUTPsk/qxcsZxxd1h/Y/4yqZ5gnvMAuY+mtKWNwhTGYh0qEQy7N9S
dl09Z/4fxNOyct/28QN6qmZw0JKcDXZhn0ONPqbxS1YxPNqW9F24PzGvIofD0VbidEPVfjGJ52Ig
eK47zW/0h/Ywg/svDlmcLRI01tOzPVTUxZNV7XfnpFzGJd4uHYyO71jAU6rsAwInUYt8/UUIy/nU
Bgkmzex4xDwD8C893kMd650bjqmUrlesu+tfnmmX3492dEY8HjcKQkzOAFseqoZa8X5BLcxaNX2K
lXt762oWw59Vp0e7fM13dsOU5edbfrs+2KYV2oR2DxQ2bLrXNaLuEBVO8UPfDTa0eHMNQQqibQ0i
Hp2VQZ+pumVaxbhGE/94AOFmGv+E3edgW9olo/zRw6jgn5gzvHsOM3bSTH0FXookiHyILMyO5h1M
CeQR+TDQQnxlfWqxMV0qVXsDAboDB6hcfGegs3Yd/16jFd6LlL/Xht8O8RZq+5CaBw0ePqRNWXVi
cU9uMiUwO6BWRyfQ8KG+61BT/1uRw8SNKsrfJzvcKQSXh1WCwLwZUkNc40VJu5EAKiRUerJGLcIh
wOFEeE60yemp3VOGdMObIquLwla/ul0O2jlPJr+wouNNgg5b8GP+yrEqiLO8Uks1CM7hxgzn02fz
aSTIF2S/sq+hRb3Ep0p+eWu4pgXevQGbq3lLJAczOnPg0ATJtn1RMgEZz2z2KT1YC8y5iOzBeRmF
2fRUt3N3qkaRDbum+iZVWfM/YiVbGeNz92hOpa+cTqI9Wf6wLdtNfib2Q5q3Nn6DhJJ4Rn2T4/kz
Z3EI2ICcMph/f/FKaZus743MaJKsrI/AFYBEsNTyuhHSgTeMqWX3F22ioPtIxwr4aqfZavJ/McCK
QaX9wG2TghUDRrhtyZFuFISjxrCg9Iqjw/SNUdoiahLHd+bo9uwdMm2qH0wiVg3xdUDCKpYCPkpN
je6GpHIoySm8KHe2NPzS2yMCso37+n+PlFqgKVMhw92hYzmvo75G3o3ZEyKM+iok2TNRhTPBgVOf
uIqhfYdS2YEFiY3A6KwZowyD9QvZHPLiTLUH/ulE8hZhu8OSsdhnkb84qaUUNv4frQsaoHbPbMYX
GuhrapqiMlB0yhb/Lc/vzgpZuXeOc2wzTCaJWeTp04X1RsKyoi7+OxNmfAE3ZLsvNTGEcoC9RkIp
Tx9JrLEQy45qmXmXenq4ovNaaiyO5UN0TdzVZg+xFCZLgcJ9u46k6AL0Oiyvjtt2pPVCYhWypKae
O2LPF6X+N1ukH01e8MgBQ3fdSBfkLJuNCcr8Hd0eqsCMXBmokDla22DZPXhNcgOCzE1GKZ9g23m/
AIn44/sApzU1bNKqBwghOjOb+g3P2JaXqeyISVlk2zUW/AueYcfzCNHXiExoElpf9kG+jGHtkfwO
knuRFaUn/B2bQ2BM4NVtUrrLhYIxSKzo55Ec3V5rz74NH3ZDNBFxqLHJOY0Eh5aLcIpd8RlGfrXv
F5d0ADshF2bFTaDxez/bWtaM0NNqbB1uBALwrxYJAKBWayHHY+qAq48U1lD1cRIF/tCFd3MdUYRZ
YTwwIsaiXRs7qTIkAWsu3H0O9kDpP8+Hyf9zRYn49jAcdxld4MEt6iTOQy+okj+uNwjQ1I4sS0ke
38B3BreniXjrDQYZyPTZTSWS4pJGtgb5YLeUhgy5P5+XUac2oYcBV8qjKLFBjeFRPoZpzfLV6dkd
EvrOUJ3ZNnCeS1oiYI2h8jljEIJU5k86LhKpv82DBI0CiaxQ5FR+9OGatHahObw5dOX+6igsuwhU
X0pxr96jjvVUh+wjhiNoirn95BAhTSzf4yKihjvCQzkY/SH70q42Ue9KwPLr6fPKrYhcu3el53hF
zfoD3NwK2Z8VgW2BHAhEXT2cdNGqIh1swtWAzHzC6OwSR0cu1wO7q6RjOWp518qyEKBtDzzBIkyD
GQBfzzgSb5Kri5PTzNTLwIl6Xip4b5ei5Som20f+HsaHTYYV2eMBdYwmaSp7Qh5wTjko9ijLJc8u
0z1aJ2ZjSf4+DMtBpkxyMz7UsPHimr8lbB//062frOdglyKjcoSb4nFkrmeKtb4rpzRGlAsXpUbu
QVfjogFg9CNTsQ1ymCXuC2p9lzkPsEkixsvMWa80ioveQ0lGIsQXLK+zV3Fvj4IFqb9yG2qf6ATv
+Gl2nbslILN6vWTZjEqF9FP5Z+c3FONKG/RVz5OiOklLLUCQOmWVdxQ0/G5Ch8+rEkOweyu1H4p5
eyvjMxE7wBfmAYmSK7tTgZ83RoWfPfcTuF1UOL6kLis01eAlX+G+aQc1zXWs710IevUN8zaI8vDs
5PV9AGEFjoZyb4NCR1bezcPdQHkw5wmygNONy6V2tay9UC348q63Njc+tLDqg1A9Gt2KbCtvOUy7
cHVzdOPBOuDpUfF+tOfA3JhU6h9FTNhTajJhlkMLTxhsO4KnAo72MNiRVM0FF9RAUvKxDxzSbMq2
y6UGgiNjmVQrS+AQBzbOo1u5pROhd522tOB4jy4kiBE7Z+UVya1UwgdtW3FKN5qbQ1cB7ZDmmGsD
BjMCjLn+2PY7HXyVhHGugubqjHJq8LYuG++wVvZxldtmEM+iZc2U1AggBSfNYekmVQO0wiDJ04ol
4IMpjq5K/u+zSYsN3yhUQb06OjLGZc7SRp1U8GSje936Ip8/yHf4C/2HCMJlPIFf3bPCHLng9RCG
/1tPNRxEZS3nqTo+HSeh21mPFFljcD4vhMEiXAjN6Iux6la+rzF2dWt2Mx09VrwmpEg2Cp6OSkiO
QWNnnpEDJcilA3+VtQ5UWKqV5IAiLXsbeTGDPBO4J6+X7IUi9shr2iAgejXcsRNJDnvQcpiWCNBy
ULQMWOqfMv1Fy7AaGP0UmmoO+t5FTK8T6DDx3COeyh+PHxPgYFXGOpNQrXpzPUGFVe+HUflgORpw
oLwCv/ENgOJdTdwN/PdmC2oRXRzcIHpYcEDM9wvV/lssS2DN8HMvSl+HtZ2LIyCOlvXm+ELKeYZI
2MaOL0eUbidsW8OosXduhfDWNe3v3V6yMOrnHizJwZkSm28Zp7mdNU2iwrrPpSshnj4yOX8n1D57
qirlSh3j2/dOOVyXT5BX5/PBtAmUpuygNKlGUmSTvuy232ccdjPhAwcgbO/W3fP5XPHCdhKQ+PFu
B7oapTjF5QjlsQlM+DV0MeiOM+UCmeE5c8qdig+eqRkjek93ouB/hfblkAeDcX4EuZFowsoXoJIo
4bindQTpNl0/+YiqM2CeWfrgRD1gNzeUgtjztHrgfRdUzH+SnP/6LgKViBlreg9qj24svEGx0fQk
Lnfs3W6nR+sBsrrpNzMCOqzWnUDdV56APq67613eCL0i7Epgt5ttweENzvv370hacGhsApIMTO+g
akqt8bKejGdxHW8JS18bwAThc7fW31MntWrySEcIQVT2tln72hAB275kVYriH4xmpoQWLfQK8TWe
2K75rlWLUL02v/MZowClY9Dk21HgLVrKIqHq4Ykm7FMz015xjqDSLOswBBC+jP9E3yVZQSxNCzCE
wKyXCxjEpI0/wswwXENNLLKnypqlzwYsrfmBY2JbAAXFCKWfQg2LleGsYlqLS5rYD4Snvzq1KZdp
9IHIz2bGPu2yXnFxaCNOZvomMAT9mtNLh6dTwoEnE8PcWZUcGN5eL4AV/tiMPe9R1gQeTbBlb6pR
oxGmFbCftz3nG7IyGj64hrsWLNrNmeAuZLtT4ZEYOVChaqnPgRvYN9fG+/L/NTCL+8bZIDkcOWv1
3d6LRSp1zR8D3wJA2OvBrnVHKMWLTJF11IRhZgT8wQvrGc98sug0XeDXKE3mz4fu3KeZP3sAV731
9WXrkakq9QV3bUGxwnIPP/QQ1SrxMSRPvqGEIQTHwI5Z6djxeTSk/6lpfw49YOI4psjdvEUvK+J9
gwiRh2KvJVjGTOtICiCTvhmswM7Ak7iXGV538Kcp9llgxd/ZEDQL1qTgapNQPksP4wh2/2KbkNzS
XrGXsMHBL1cGDQgonOEq4gtutpbei2hKUMJ++/o+iqQLpweSWIy8HDv1VsisjlbuScJQxxsSibI2
v4rojN2m5CrnnjKITh7l3mhNOxBKIu/9eSsXWPzDipda3yglIIYpdSE7sLU1uSt6rwA1pHl75IOQ
TO/vgS5fvZKSz9zRXwR1a/WutgWg+Tik5vMS8L6zUS4O/+yUF7rvXZYKJSf1PvEZsXo/t8VmvasZ
taLcftBAsQ6xKD+igOSiirLSam1iAabB6amW5kFuD/K00ZZlJuchER9iMu+fdIaQaF721W/oPixh
zmY/b/7SW0mm2c6/r4AmM19C8iHPHmWpV0o6qPyP190hSCAvkA6oWNYxhKhtizmpMaFXZtjecKIg
yoZoFt5oM3LB97Um234n7sx+ZAlgPiNXnS/PvGPwuur07GmGKbVE44WkQpyTSk7qplgMOjn2VzrZ
XS/mc6rqwoze1Bss3FXS9WrVUxXuCLONIlKY5NKhy3CILs9mGsWSALwBnsDyOVjyeyt5iJon7nBq
9O53CvlTHawvDpZTx/kWq+2lyK8Jif0o0o6ii0htK+yK6tn49Pgav1ePH1ThhMCF4/KGxFegdx4Y
AvyPDv92tzoQH/8gvtL4r40TMPErm4SS0aSINAqe2gbsCCbmBYnxSjJWBrmpgRUAaAGxwYdp5I7Y
2VlsFM6Bi1NfthjwABf7+X/ZZgR2TQveUsDlPY8kp/r/IDl9cTLGen829lttkjD158yhP1YZFwBj
hZyIymz6KqomOEobRe7BO5aaL0UKYsz+GokkY/uNoCQ+mLeyB9yd4Yez8d9ABFcmmN+Wn7mPmr3f
Wtn2DqvVqc8Vudwb1nwljrDCEpGdmiUJIIN79Zd42iZXmYlsfSx0A41ILzOKCxupaGRxRGzAZtpE
LFitwXnkYaiym5m/FJhsB16rXzf3yoiQ3j0i1oxf54lnCTnrndQVxD+BnQR5k20O/wKjEC9hZAV0
2gJ+gMlkQ3yYJ4mBCOxOaJ51B3JRerXWcWbblgD6qDLm5bjlisWyVPAja0lFB6Imi+jtlLyJdTOe
SWzJyfJb3eaEAjnXRYwBFslSGcLyUh+/yIcnLKIrjT1kbxf+M53noAoZpB4zu5mzRzA0n9KT1M5h
rEl8rH7hvFgaP8eYq/eNSeF4Dz0cOC9lDwRgRhuWbXvWd9j0baln4TYnV8+gV121zENjcMfSiKhD
E1gG779o73j5xNaFuSY/GejrRAMm3NbeT0adF0z5Tw89YpSg2acuXUEf7xVf4JINRh+YAbG/7guk
EjeIGkQe2tNXOJslLbwQRgP+5PvCSby9PewcLP055OUlKl3E50Xts64pbp44e6nRJLhUVPbw3e7M
pYu9tfKc+WfN1jJX6C8QTApflQvRvcU5Z0vZzeMZpLph44V/wgkewAg7/9jPvfua2yRjDCvY0ULk
WXRadRTC9qxpZJiTj9QlfHF0j0qTlcplYDxWiSPVzWrFw4yyRgExZyZMsUDDd7jIiYh3ZSVZ22hm
IJmDgr5kwOyfiNTEYORb7egpRe6+utG1vz783V3PDz7L9L5TwaugFjgHO4xmGtaISbVbZD0J+wq7
7hXOATpbMUqNfegEHSV0WP20FBQ8Cs/hIIt/GAQ8yzcv/rnPQ5YQHjFFoP843F2MKML2c2L3pqpD
P8g0isTRyk3I0AkFk+SdaqOGuzxBZ4WDGMikuVrNUd8NcGEHNEdOI+5a7SaFA2J9KYNmkZwbqmWp
XPz/GdWncLuwZo8OxcwIBu7SE9dU952LVRJzO2gjfhmQscblqx4uPqpAiV2NL2X+MmlH4CZ25lY+
XUv5yDF+MOfPsVTQBjR3k2xh2DtgKwEOeuXnNKULCWVtLGDAkVpWg0K17ISGJd5Dy8XaGN0rBaFw
ltI+WXCwq3g0peiGR08WYQHPkA4qDFhmaFVO70CBDBoTcRRJKmmcUGOrvd8j4khx6oHEPKLMMZ3U
IomGv9H2PNy+0Fx82XcxBadOqgtPDJElteQMFExPhlcrVYiyMsk3zbeRE4yoyPb8jeDbx9Rxr4zd
4a2QQBZynC+HT1DZMvepOqLY0xaUK7i+jcm12/cuoIuESimz52OIYuFsgPM1SR2Zyv5gY88FungR
eb99MQe6wpiqBIAYCVBB27Lk5Kv6mFYHU/5Tb8YW4wnoootg10oql1Q+L4LjgSgKSQEE9iJtu8Mi
7MBXOrqgQVe6mdGwtZhfPFqDvIUKqKxkRHM/hoLa6DB7AjSgd6Oj3P/m2/0U/uw+YzIPEVzf4grr
W0q8TQeB6IZhUiTIUCvVZjMLhXaNcC9eqY2ZnkgJlVr/EoAlpf4Klm2QobCV6pUuQTKys3tUquX5
3crUQcPtJN9P4jqb+bwJuUSO6iEVDHtmFHdJ2bw7qsJxjtPSQpb+d89zwtd162vTFCNtueZSo+ZS
FQuY+Yp+OafGf973j5C9ZmXXXpOvPh+9Nw/Brb3Nzfh3rzPe5Xf9mj/yZRExdYhnPtIHzxg6ZgxW
d4jXp4khzhMQ+qCVBg+JcISp7zUK7sGuBCRZH8n60GrZN4VPWpu5ktqH8Ygw0GgIDqFZzO19RJri
naYKVnI08wdJITA6LFjBECEdfIPPyiYiAnUy5aP1kqtucEZTbBHGRb8uRyJMCZZJaiyexmXyMt+1
VAvn8ap81BKbCTdDalQ+PK5IaT8iS3l6oa326jrUipecv40MJ0veZOn6MOQ64bc2tQ2AAfcrujA5
Nsmu0dOwcbOZRiAEnDNvNzro1osSclzAMZMWy0AsPxzARV5NnbTNdafovaRydj7D8ZQaSV+ubdu1
VG/tW9zPv0oqJfMOg9xtKt7lozHM6GX1sOw9xoC/nFwKpHRZew8UeqBJF3ljN/Eb+Z65sCmPnrTC
JhMXy3JVkXS6kQKEJYSeUNaB63dpobxH+VrZloW6w1fbDQTYLX0Gy01oI9JteAgCF1+yOeaYtGSG
WEd5auxo06nuh691bUMLFjBrGHypOGIPzwF3sXKmwdWuWBiEo9/sVm+XaklJRZACHlE2LnDsWsYG
Ph8FN8yMohWPSkhECsNEP+82IzIN5y2Y3oDI1sPJV2rwn1096vQhnk9BwJgbFcsv81bfUohmeKmF
yVQ9KJJpaT3jDpScppJKuIrGi3mlHpChIphPi+xD9WAiKeJHHS3J8M7PXXXSINkirM2VxqeIz0JA
68kKIj6TVZw/443bvUA7GTo7CpjHtCXVFVozB3hG8+yUOqfcg2xjW2RNXxIG6dVa1nqhikH6RBS6
0b5u2gxFgoAvE8fQjmg8KnIMVXtkDiwz3y9pTM2UyPml+iHIxfWAEjquHAcjQrPLDcNM/tSqQ+j3
MlrDtGlK5EnurWtLuGy0M5mbFT59wOs/vuWR6baUg0VuFjxZgLB/9g8zUXZvxcTAJSoq4xK7rigG
A+nb0LOK1JfVUtXJUWb6KbiiheB7jy0+tNaqKmbY8UI9BSLLb4VSG+i16jYDfn9Q8t5H0/JTOmWd
LvVKsxNMl26EMPnpPFmysCVsyliikn4N5CABiCcaa93f/uC/04kEsmDjAW+KCKZqOit5K6kD+Wus
p/18rzMF/yw4paq46gqp3mvnzmQJgjkauJW2YJvLO89YOYnk7tMW2A/N/+c/XTd4m/x/xPvnWmht
PIq+hXDo2cXtnQVllZECgiSlyVmb1AYrKAqmWKq7mlGLrUUlmHhgXz+RizLwRsacteL6PGPIuYHT
sB6JfyQyU4C7E87qaG0OYklT5MlKWYANAwFuqp4nkozTxLcjQWdfCzX/+uotCmJG+orKFIbyiS1X
BVuC7wpqelm5vlDomLkyFvgrPzmiJJpKrgeLC4qflb4l5+t5xxYYZ/73+aGzAsvpxKPfSlTlDwaU
l20fDS1R1/aCcRsKi3ZGnHYuXweYixNqGGQurUzeN+I01iFeSWBybglI3cgCKBubTc/DDUEx6iYQ
2ygj5vG5DFDC51MeTuf9xY5yseaFYsvVC+6MHMiUeQVM1Bz15KB4QMlr1QM6PjSlbkotXgQtiBQp
wOfYrs1O/KZqBLin09ZuvtyUQYRIFGTcu8F8+5yTzX54ctz3W3ps2v5iOZQIVOMjFFrX2/3tiM2T
ez2/6LUf4TTZh2ibP8SxsKI3hTGpTWf4fzISoqmJ+HNKlBRJaa0+q3HtwpV6yndZCY9WLldCbcy6
6T4+A+t6k/cO6phXy+SSzpDOEr0pI9aW9a88oPFfH8yYO2RayhmRkKzM/pq89PbKFl3vM/Ww6Nxo
cVM+f/kEw+Lh32/QX2qadC6urwioMJ4TGv3j6T0JaeHbxcalmDkGGvAAn6ink1y6ynAyuCR2idzb
A/KRMbrTSvDTtgoDCanep0vIH5jPFwVgtcXqt3N8ExTK8ohXhQDn0sE5Akl1G4wFbBTwrFf9Kid0
oYKsusFZokzZBKFJIZCJJIzDEq9V4dKvJ0GX1fJ1TuRkuESdJZzZT/LqAm/7j0d7bnujVVAj5T1q
iAgGDcUwHwyZIBkV2h/5qJ5cuqQPtjkArEDkC2UimuF12IyhzA06ClfpzH/VU0iwBpf8hiiUpJsQ
swLXd84Zqi7L+9I6MHp+VYjTk/hQilkWoq0gI/hUAhDhvaPeCQxY3NcQPdgR6svTbp0mxV6ICef+
qw0iSAUtJ7ZVj98SEIADdQzxaPOEgLTGx3bGKk9drP1iMHIIAkRwdB1i4KrdcqEO5VND9cw9Evp5
Iat0yzFxWXeMAx1SEzi3ej7Lcuc6vwuYhhZK3H14Dyy1RHftEJJzaDcVuew78PnVT7blQ3YdvLyj
QCgVCr4FqmNFkVWd0qzSageo/P3KxE4OoCWLjkgYMV7QyFORniYGxyUqvoKTjVXCSnQBZ8ltzrnc
nfoYez3Ahxzff/SkrTzJ+3ywbYD7eGDdLgTe+8U6uKSADgwOwGF7H4+hULCFyKRPRY1l9N10i9qB
5q5b/XEQShZpFwAccYOySKMfnp3zVebXFfqyBQVF8J2PW/lYfgdZxE3pVC5GsGLy0rJwqDL+cPva
zraV6fDhNXhzBmbxD/Op1qULGmtrjlERPKPJCQZu5Vqk7aKaqiaf2aWV7X171uBR+nPiurCrehJA
z5IpXrw2AshnoClmZQmlpzNRfY1RmfgFn1SepmIC+NEkbsPW0yETYuh10GD1kPEu2vVZAAO+ras/
D0ImnO666h9GG1VDOR4cPy+qPoQG03y6w4ztRbLYQgF72k6NFXb6VGO5P3fQQkBTJg+F4XP9VgWC
v2RgeX22JJ91wEuadZk4X8eSZ4Yn05XmywLkTMiOtsCOytxjAi5ejptyd/VQzoLbUXki4KZECIDd
s1m5Git7vygxWrV9n9ng9Lnd+XEEcUZg44icwPlUFcV3/RZPQWvydqPwqEsrcfJF3tC0fBW+1eqm
A/2Nj5fvpM2DBGRBPSmFdBAje+KmCHetlQaNcl0JDqB4dgifyrRaXnz+ca7vO+AGJcsupWLsoGTR
J8suwfnubc8YlMcxWPWP52AVfDUXSs0A0kmmtVbNm8njyaM3IzOjf0ecXk7IWjlEFHTWkpd0DNtt
CNsWmbZeqOqzuKadS40k6aGPOai/W/swGYBhqkvBksg24SvfRl3tP7QlNDDjXvboPZ3erHAGuxJW
TN+DnkEQmVbH1bE5TfPL0bQn1Tjo2HvhqydaqHo4h3qc109AQTctEJI7+9F2dH8sldxNmmgVbBO4
tnNwW6SZmfufuC0s5L972K4ya6lLjlBJ+nio+u13h7dZlK3wUXBF3uJ45XNnyu7zMu00GW/wFpAr
irz3e1WqszjxSguGwVU9zHncRgsyj+t11Ki8Tb4/blZdNgPmy1kiC4bXi0uY7Q2XPNmsnblM/mF8
eCsMarVgbUSusVa1WgFeTW9Ba8ED/Y/MZnoBjBQwrzxLdykN7SNrx+qmiyGTqtaedEwLad118ruY
SzAlnv9+rUCnc6aOgrV1OtjkVE+llEL9TWonnnjTFrvqpN1CMgYBzgykSE6Fj0inMIHbH2l7B6JC
Cl5MUIjn7ARZ+Eq1DJ5vU8mY/eOTdj4UH2djXsHtYfNkC6GWgxGMSpi66FO8kT6jcQCMJbhVx851
73fiiMBkq/gpcpwFhj3H49CrKks1AijZuM/1/aswr+ANNFRMGXOAchl/3vc3xiDj5iI92ywjfZx3
UijfK4SyA9t3RJHB8Yh8OjubFDrPAVT/ZUPhQ5UxINHpG9gMplnFOEPXuRKpjxrhmwrNx4DwvWcy
EM+gdeVS9KXj7DNuh2lVs+cO0614tVc96gmhYLB4ais5HSb57X8sh3gxYpix7s56CptVPa5Z01ks
n4oQMz/jLlQTENftZTt0vlsZ2aBjxKkIme+HBZzWXVduiRB1Q7QyYHqErk6wQ72w67NK7hhk2C65
ZONtLL0DVM87448WNOm47d0PRE676VpCkuj0RNmJUoi+IZfTL8ik+Fc287gUp2+0jai7Z5r8uxqr
xBVnkFYKzfhPoKgUKkUEJfNcK8tKM0NPbJkfH73dfsUD/8NR5NfvVgkMh4Na+PQvwx5vYfHTi1fj
Yyi305yGcxmZ344J6jvVfFVWF26VmfYQrbZQEirCvNi+3BNmIVhzhz5sHfBGmXKpz0CN3DSSMvqi
ZT6Ti7//5JF9UeNYgLiAp4v1LZuhQwhRCreaCevbMxsl/FfLEDZUq5oWE/lYUDQiTKoHPHHamN0G
oqDEjxJL+ElIEvddd6lOi5VUziRN04l13UBi1i2KD+ZLesf0/XgslcLbNXnNvG2+ptNbKwpxXkeB
DUe6QhYQ6V8FpPQUfA39qfGztoJm8kayuXtJ9udDdBZq7W/dKKp2gii14s3mUXOtiU+6SIJM+n0w
14Wz+15NyW6okAuJkuQc4GnvOvWps2O8AIXdRTtfhofdVA2gBK6IYoHhjo/PpzK5tXn9JD9mWivS
OUtflDmsdxkImSyGB55QmNjK7BzAUC81GgdhKO+YT9CTqVZhic4laHw/cie5jX7l4PzBdRB2k0lV
iXEzOO3diOf0wsvpaTFYx+X4dfg1YqYpv33PIyfw4g2IkLVjwkNc3Gn22MGnGpMyFNp13T0Mtrl+
Uk6zR3p+6xdfOaaMHCv1gb5s2KMIhrU9KsdHNotxL0irW1KqpYIGP2/XW/BXeyScwPOzCggCug0b
rbEgHa8MnAdCncnAvQCdLh1Y43QlMFppWf0l0j/Fu2XWd0gbgCK3HiI8TPFqzCJmuZW6niQfGIEF
+pZHn2D8Ih8BX8R+EsGNv3BSN2fvkjI3eTAhIKhAaOu50Gi6hVkLbI1T8CtHjdIoWLuUXw3/GEGO
Q9FM1JTGXKCJ2g1nmmNYkO8Ch8rrH/t6m+N5LyFyv+/D/1baOSkH4ovdCb929JqvFZPUhUnJIQDB
YThjcw/walmhF7FstUA9VaiS9dvAKa2ZODmL0uWY6yHoBDVXhPiZblXcrkXFJOM/kE8yr4UGbU7o
rfuCQuZWViiCUZxc8I5sbIaZ+gsxcD9qFEz8XE77Ad0DzcxXwvAoiu5xLpisLWzKhZIT7nmj7O89
ywUoMDkZup7FhZ3Hr/UWFgavhGB4fTvFdu1odkQXvSZQSubR5mnGb+I5HJcKmytqsi34QNIdST/C
TB/xa+o+RUA1mxuzXrzCHSm+sCYAjzRouIulkTb6TnUVUw4Fr7cfFek3e+uocZPijWOrXMlMK1zp
5bIsCh0goG+Pb0IBtcoC2kzyIMqM1Fk/b9u61aCKAeyF1xivTNHEYIE1sMoQhTefdZIy3kIRGHAS
Dy/Ph3axMwMnWc7WLUWeGB3xuFNQV9zDrqQFAzQnPb2l4Sut9VJX6gQ3phCGaFAg8xd0kJY1IP4J
p6JvHieD+PDM5YYJtnR2PjNoTQhmCH4qtHb3MsVftQwtphPLMpRSSP7u1iPadtsjDoF5HLnLOhEy
lBHo6jCTNRQKhk5R0v+yYxUESaY/L+/sG0/IPCbDmIo5OP+9Rhm4T8AFgdQ3dQF8fyjrDfuu0LzM
756Z2NG9NYDKEFyT1fjecWkx5WWahfWku4MunI56WwaP0I1vZk0ZmAfRlAjVxxrGcdktBo5p1rI0
wuTKJhqcXDGdkMK6YygdkWYb/ARbsWTwCTVaBulACweAz2GRzxWmRLR0L0xh93Q01wBoTClEPN+M
YSdeXvH9JQzQL/LHtJRTfpeyNWbtESts9Qjf5v6wShLDbEqvjZBdIuRHQTnydLSP2T0rNnb1Zn93
O65PHv37UCLIVjkaiRzjjcqK9WhJn0XAUf/jw3mnJ5qDsABhpuCQfMRYx+blAv/WTyLesJRLg8+y
JQuN7VuPups0nEymCQTtcDcDs+jxgMi3IdgiPSYPGQ7zKDO0pnkbiqysTZkqIH8OxZN+sm4Wzpm0
lmUVWV/GOLjrUec9mRKd3xuTJFtnFGY3mqs8ZNmo7ck3tHt8hu3Dy86zPNyMym7puirySySKWL+m
wSL14FJMgYWoCr8n1dYnC4T3LBCSXvllEo9IWnEtAt3iYC7TSQwJnp6tLtNOqcbpD1KZDr2RgPmn
i/CkmcUSsdNSsGlgoz9t14xluoCjATF+iUvwDpOHrqNiT9pcnaxHlKnJvRdoGXmooZhAalgAuL57
+4lo+D4eMoew+mOAaprTVU9zTqaVjpMLPoK47K+82E9ZN3bIvgWyAyloqnbe/WDYVogWgeefQVSc
Mh5FAYUQhUYScOMcobcyoCyku3q0BAIL43GMj6noBcSksOEC2XFC2XKLAoYPMIsFtrjZopXhoIXh
C3E5c4HFKPyXyyLT4MoM//EpRwV6HFyT/am6Fbbl3SjGgk61we/5FJehczt3p/kssKc0Y5gxWKa3
2pLnydBYdJfi3HyRMfEwN3iZeRchSCraGWgXv1hN73d6zIVrsTFoIl9mPHghD/A68u7A4YSwP3/m
2vqrcZDh0qgFi0tPq2Jr82MDBxX5bWCJSNSOrGJIhPizoNs16ngRu/CVm7veyXZupThY9xX+eNT4
Q7UkbdnmYZrg1uMzCr7oD64oJ5E4nWt5rsR6yZqqYYG+nBps9qobFth8U2dJsoi8TdyrB0u2X+5B
eTAra1SVeq/1v2VmsB2dMP3Rs2JTdLJVZGrTW9MSK7I4FA0Tg2zL5ZDyolP++tPX/VyCTTbOWg39
6vxvp6MQtnvIMvcStgFgakzEu4FG12J45WxMqw/cxL8lTD/EiTBh7jQdF3GlFPlmHnalf424KU17
0DosgNFZu2oHJmQLbf20fzXoKjGWSpRVDXhSnBz5ziGO2ycFIydfpT8177vchw8hTkIPDcGCPU8g
pUuPfwHB0VbTfKskbUt2TpzZDG+c4lqzg0WK/P9A0sOoVQDp170DfcU7b7NhGaFrpYJHMWZfhe2R
0gkr3ZtkDzWXhs0GiulLxM0V8jLK4pSc/eb0nG3GqihRBaTPAUaxCBNYSBhqa8NKnmLOPxPSLdvC
PaRYqYszoQ23HekRngBi9f9wxZV4mV5AemdxNwkrlvxRFBMURajCJTLxwmnEjWemIKfNPfX5Ut23
CJzketqkPRdYoLfNa+NjsAf0E/p6JHM27sTjpIvViqLpsfvZ62X3bbmtft37znVlvSsEjw6MQxya
CcFz51rtMGmWJKQ/tA6JcFWbRStQhVaYsPniuJWnsNUwIMcWVYR24WW54I8YaFVxMjHB5DJFoe0x
Q4EmkSW27Tw8zT7c4VLEq6NT0/94I/3wTLHoYoYiTr5B0KkwhEuJdaxll34lRe2T/8EUMbAgKDf+
OBV/ODwALzFzanK/un6mfQFZkf0L4xP20K0FIKbJRtJ3ckAf7qQCNGgXPZZgJOzX4cJ84VioeYIs
T2QB3G5bXAb7FRBlCFs8g7Bl9InC/YLAbeaaQuFpFUpKVYkkhgQTHA4B1q0SE0hJuI05JhAlBoaL
wvHc7jPblj55eehSk2rUMc/fBtklasfQraFp2+gRm5LqOOXviatTFxPciQ0rW6UhBY+upsAb7OFN
4T6rWJXZ2seW9LRrfgUcxcFGh7EbOJynwUZ+kh9fW01eBg0zbwGyQRKLHe6fELeIwET5vSr2lZWm
NS25XkgbA2s6DdrekfRUJTdraIDlMZDovwl9CJoNt7aZtUgBM7clamFAGdtqfZTkRYC8vjlMg2pw
Q+UbCHmd5MCTsF7G3nfhNolQwQiRlY6NtC6Zw1MCoB7w47FrXfMRcSYcFqWmr5eYuYKpiQKyw4IT
UpgGCPvvxRchKWuVCB/TdtJdCDnNj4KGr0jF5DujJhlQ8AHvHSvJUy/oQzpH0L+Bze7zREG9LwZz
mvYdVcbfoCE8noibk9Ftuj62TvTZVQ0k+P5mHVU9g00MVCYdJ8r1wn+NUMUnRXSXpGr3jdqTzrzK
uTcBZHlFnNkq1RAE7Ju0C2ujBuHreskXS8KNWJmqUecu01Nc5Yz/kNPegtV8fkro+zAJkB//9a64
1q5llA82+EbkKXzffUSkYSgL1ZejD7TKP7K1oTQKdb1j2LqP4YoP2SbsCk10/3OEd45qeFz5KIuZ
KADrCeocAAmMbZtfmWcHHHyTqw4NyCEjaJfwgEhJDCQpVxDCS1k/iQq0I7yBlZeP7SfnwX63ZFII
WSAPLrd2wpHuTqd83bLHLBUrDN5x9CroFSAkQxMgAwlvZ0YzjFQXJs8/BfEPdPh9BGUkkTt4jUch
pzLSewg5EbLHZB8meyXQqZ/xsMG/GtfMzYtFEcBMMe60qHsjS24ZMwpGkTbtn36cx83J3Hlff8Tq
+Q1ikKYpBSY1rCYMqc4herUVCMDMzlxYPKuNMsPMkvjj4+GzKrGlqRyzF5S9GmMbx+hw+eb1+nWo
GfrjKo4DEsOUJwA+impGsOMFAsCDwU/atXCQ36jSLA3Z+lSqtLI6aQzs4SaXRtIOvhD3q06hOqKN
v5q3wHaDDzqQ5XtAsquitRSOOQgIhVWfoA4Qn0VFQoU401OEcJ1WrrpcNwA6CZF01iWrl6xuggf5
bkE8vu+P91fM8ZvQfNTt90wWAHFQ+AApXBN6quckN/xeLuvpuj6w8UvRP18YO52/uA8sTNV+Q0za
99Q/wqW+j00smrl98kU64kHM1ilBnqUbRdtGVtU+Qp2jFG1vIKV8LMeIOFN4Gapv04r6nv3cv78K
a97kn1tPPaQ3WlnGy3oQillEANOpsy4zhQ5shAUDkZxNGAgXFVWdshlbGeuXY23KGIpgWcHmdRcQ
22e7ut64E8inApOY2nCFwavKOKFtR+dON+cC1sOGHzUWQaYBQL3dVH5hNYm09heMGlLa6aKFp2d0
yvOhV5ASOqdFHTHWVBHfc1LLCeWNGPwxwxa+/x+5kY0T1clRVcifuUcj217P+p+b7fy/O8e3k+gc
b3NltW7FB6QWzXwtPZNCv4S4jmGYi9FKARORow3eXyYpwFQSpxhKsg3gKDlV5vO1Sd9tFcyl13Bl
aS16/FIKla+IRcCNJM0BMdqzLjYHLgAN8VLbcxVnSS/XhqdGtvPu08Py1h2XjUHU0tS01OweRqLo
N5lI0E31/RV02LLk35f4V/yO5y9rXcBURuizd+9TTpzombqUP68iqjJFsFJGokfmICWIH/OQO4Wz
BUDiF2SBo2UTwCcWDY2Ngz/Lukd+85vxRyVsZ7lHFLDd1J99bNt9HJnTeJOl78sMlOzL+BOs/TMv
43uXyZu9cfAC/R7NSh/AO5wN6gcX5LzWyX7iRoPiJPXvK/+N8I7TIuJQVrsZXb7m3r9z3p61jfl4
XC0f1HwfeDk2hJbZSXF+hwwxr5GGF9i2ATOHmm8vIY31ysC8jU5ExIZxVT+C4MYJ9EcMpC1VqPsg
hboU0l9zX9+kvKpbDj19jRxwvOO+MVXBw5ycr1l2yFLM+sbfpVaW46dOOyvthSDKWX/Y14P6tlhZ
n+v9aaYmWP05+DswS/E4h4ppEAdVe4H7DUipiQMQvVurmu8P8v7Mq9RpRVgudJ0hzzqPlTnBNsA5
Zdu73QLMYvTP57zBjMekoXe/Um2Vc6P/PckK1mQL7GN0tjzDzzfjeQVcqxCzOT0Y5oWKtJJa4T7H
aYqMCtFUgQOjnkco6o3na/ClKD0fawd8x8i2wCKcmxjINIK7r10iVHlbfo78R181FfsvHtTI8Xge
+z+5LhF0mqGNtF1mYts2V8QUCZ0a0wH0XgKVbRpfr9Jm8jIIfZtefgi502SHRyITjzJSaoE+oZfq
JhLIiyAWvJWAcbnqu1j+ED1NF2S3cYONy6Ha2xKOevDYhGXww77FYwWQ3qTAYpDKZbnw5iRlhPAh
9paUGqXLum7D/y5DYYDwDCncW1T2Bk6ewEE6RhIT0cNj/bXIkI1uyjzTkYHVKe9dGuWuwtjrdVkU
480gM9uawrR2I45+nMKWEjedpuJRI59CSJVd2KUuG6P4cVyu5iT4naCoWHdfvcoDKVJgKtGFAcKW
8Fq9elXcqBRHYcy3/xBNRhCr3eVrpdHmzMW8reDK/u0I3j7vFmHo6rvXHffvFWow7cjxbaoFGrB8
nueFEcBGp5Nno447Jnal4PhkJcB4GZfqKH1VGOGv5MPAin1rokjRGr2w/DHhAScvy1fw8zT6IJGb
qkPaYgY2xKFwbn/Sqx20pKYPK9o2Fe2HimF0Ug14yZHb4qjqrkHwcATAkCt/Qa5v+X3jcL7dtqsp
DrXtaoVOt5yVyBKRJlRzZx3K/3XPdlN/ixBSMBPxa8llroSGMVCAEPjlJyuqb++H5CCCkxkJTNWe
MFA64davAKTyxMLfxto5vgVXMQ5MHZEk+Ec8sAf80jD72esGdauMLF86ARcDiEx/6ylFk1X7ifcl
GHJXfJmmk25Mn1zeOPmJkMCBlKNmeq9C0qxCZhP3LSN9uxEOvVZ2Qp9eIwvtq2XQpt+vxFA6wBxz
QaAVQdp0XxXoJ1vcd7dvgctHHDaLB6n/F3FTSRrLOS/eTekU4airplNNnMZ8rUjO7Sa5gUPrciJD
d0px/GBz9eYVy9y1pW6o6QDuplU4JmDgQsXP1+yTAXWbVmkyBXD3uMxhO20YN5OcC6gVKp7+m4vx
E9L9UoZeYhPP4ejdFuyzdwF6M0bqODjfpPm7Fi4ZCKPIyHm9TVxwZg0S8PQBotyy/9qifz+QjNNS
/f+K1McRpDI0YWUH/VuJAWfll4X1tuE6qQ4uhfSRnb913261QaX8+xdE/nynh7+oDynb0W2etWkG
6gZzUykw97Wt2AuSFDtQg+kCTi8i0U1BKCgMF6xh+mFpAO5DwETQE0ZavDjoMAqqC0T06DSZki28
iQqM+fyC0vHb01gXBTddOFku5apG/VODnLBeKH8r+jie1G5ATzPgoCjAZ/xXjKBxzbwVOOdIq701
ZHiFvqUTMm9VxL+fvs3jiwfGq5qIUmvVsy/PaDT26EEmNUB7IrGvgMz39waL9aXKVisoAbpdhuCi
2Izb2u4KttMMDnaU+gt0lpCCeiJs78J3SqqaavufrxW7zYPo73r8jUAiWKpybgJwmuZza7DSxLR8
oozGeOZkcnkBHWfkq7oSoTm4F0cUFoA0MLnEZCUHHyRc9tVflqP+j1yyp8AqWTgDA84L04Jc2ZCd
kAk0uo6/FCis4vZXod1cS7dfRS4PjbVEv8Zp7L81knkzO7tGPhc4hyw5A6eeoX11DqOo+qdRVB7t
E4ufPx2TtW1wx4855YQY8f9RN3cb/Vx150/G7S58nFIXN3Y8Mh+Ger8c0aSc9NBQrpbCnfi4J79x
tAXsjTBo+NCwYU6x6TDegqQ29rW24lCP7SUL9ixrclVnHJU/1Rlf+1mgGbOnzn4W2VzyGuW2BOai
TsqZohN7q/gJyvgLOyzPUmI5Cnh6poF+8+Ihli1Xp3ptM4e9/7uJHJuekEPIryz44FEL1rF6Q6sF
x7Uqp7HwZFlxYxW9VNwAertlFR9ZI1Sek2uGTmCncoJJ93oCEJBpdC2ktgihV8XbOwuXg8raN9Xo
LLIYyh9ygberHuMqfxGcYZuwyc6+hS8OM+bz28tM5cUt2kifIZG7hZ2maIAv94SRLVQ713h8G03L
9Hz3W1AoIX37BXgKpZmuzBP8vWuzTYzcPFNh82vD0iSpZ8wwdFTbcH0/H/+YLDgkU+cLe2ippXPE
8QJa5EWlJ0bsqosRt0Wjc+XOZAD9zgJwwBU0KJoWJuUXo2Af9LoQ5fACGuOh61oyhMG1t+bIn7ZP
YeSMKt1AHXFHDHJjNEj+b1etUbAMo0Yz+uTj9jOr1F6jV4MFafFz1Uk8xsV0RmwLgsdYuvVyUYwE
mXtQiaCZrGx5ikL77Gm3rdturQxEhelU/J7naw0dhB00BleE+STUtQCcpXxS8K3m1MsjfTHrSZPr
svE4dG35RUtCv/bDtvC15s45l6TEJAnI6eKGnSBOvfpcAB2nrdrU5s9/+q8zVxU/CbLw1QSsM3op
bgtxli0pkf/QE3KZyYRhldc4GR4lGp8rRRlu40OKorrbDo6snQ+C5YBJO5SG/dWtovG76PNkzWKs
8wXTr+5q9OF77wjl9Rkh9ENZuUtaRPvBIq9D7xhYtbYV1c+VtJNspApPgNay/TdD0zukMDSIhv8U
8cDPIMRl9F5JsYQHBaF4goJI8sYTCBsZlDo98jtB2M1BptvPb7/rdTczOCqd5Zx21h2i/qlSMoZY
NDh9YNxLmpY1eDmUBhXFg99Q3QKFV1Dw5Og5eTFHocFIs2kmVzbLcgLCw+rwYKC7MtwSa+8Ee2tr
RELsEVCQO699JwhFriMht+PxAv1p/oUJX5KJZj+mf1hULkziS9sJSqDXpLSwHg7HAgQSC/M0Iqa3
ZtdRcM9MbomnF6w78ash0qlE1m7QLmWaovCIQb2GxBFyE2UZ1xaaJehIQ3+3sS78R//aIPmtyfUH
zn/eblJNZEZ7KT7lfdwDBlxq4QKggxcaCoL5daAdRm9OF40EBOaBFb21eW+iJtKj/Hte+9KkoEwH
fRn1CmrixrZslJLD24AtRvU4NOFdcuhUp0bpqYsxpxwQC5czDuPtHSgmvnQE8wGmAHypypPrS7Bz
5De6MMmvSWQ+FfwU6Pif8lyHKBIRGiQpvZ1DcmgnQdhLewc5snGbwL1knvjZvw74Lxx+FWFiYZsk
Xq7FM4LA/2KG6gTztAUXVdOESU0bIz60roF0KUDUTOfoUPSeZs/X9uy+4+vCyQqCg/kkONvrGGqK
/VSu8D6F8J/zCg/Pnb5weq+/rjYSCoR/b+l0HklZRcCbQfxmHiCl46t7OsbmZoge5guMuk7cwwa2
UpdQVFspmwbjAIub2JR7C0u9qf008iYakb/KqaCwVGM5EoQ2/EPIF3vpz8kBYjqYOjtkHPimRJlP
GdaU1EifQM5DDvK82B6LaWblT8qbYLrbtfSFULnzlj2hVLinwEfjsO1/sNdHJ/RYGJ+xzitJCakH
71lH2BFSVs1BwELlg+W5Jq8HwO7ScOcgUnL1NSrM/ZF8FObpTfSV6+m9EsTEsnebxkbleNW2D6WW
m2+i8CZgoqkZW8uFz1w4evUiIq+hRXNCViA8zFPKrJzkyLYMyqvyW7hKmnr8jtfPcS/sf3jk8a/w
tDU7L3xU8qcjbyLucwEs2w4gfhrISn8LHrMHu1XafiRwrvTWov3mu9OrHwJNNrHsdyK0ytNcT3S+
pgoU0BKT+rqOiCL7tIowLzhppxsEZ7ZNiTLefXiKNqPiteIvonA09hsNTLRHB1bE7oRPPrIN6KT8
9NhN8+yc1dG5fenMhNzk+aK/qaZoaYxBhNMTYY7ssb53ZmohsN44AGFiFgLDq/fZ9fUTjYCvfTB5
mio2TpvPaaCAS3QCwWAJkcQH18E6l8R0cvajtJ3ISnkun8eOV92qXWOrqsJlJv8nQSS7Nli1hJUQ
I6Xxzd+uCM93FGHe1d9ioeEFHHEFrQ7/Ssh0G1yf/r7zFfSuMYdR/jirJxheePlkPsnDzfMgHa4M
T9Zl56Mp66Ou9pZVFTAl7Wc27qzmV9ZaW85vmmNnXHNoS4DdlWYusj+il42Q/uDlDMCqZ1awhnOH
RfWvjCHsToidgIwwh00bGLARnBFTYzLNPjfSOrpr53GkxlbQOIW8r4x3bHTIh0UvDDmwZxmWxg8d
Oc3hy1cmsFZqarzZRdzwm0P/iomp7zMntDCh5qXR0BY7pjiZAO+UxlMTg/AgPEV27NiuCRJcvazR
1PNOLUVGG3d6a2HI3Yw7S6XtkCvWcerjU8+S2K9BsFnvIayfXskfzB5d99Dn6ri5IaG7GapPNz5y
j8Qx5qaIwpKJx4eAxhqux8pz6rUnEcv8hgDfbI4aDFcz60s2WC3jvU7dyxKv81k1/sF0Iafaecdt
kwwQBWpIfd2xN8u00XYi16rqVUecN0sPnzSWQqDsQ0shTR+PaBivSJMiIJFN6S3ujarAG/6lVxuu
IT7OfG8uR9zhw+STIBLSFCByl7chFbnW54d97EYBbJ+RSpntvhb4+1mpgp/0l5KfkF3PV9S82eNd
D5cUT/7PAhp0unLQqEFxAYLiJ4G02lxNEr1N0U6f4TDlkOHM1WpQOaBy99Ixpa2FHPO8Qi1gCT8E
5IUJJGzCMaxbZgpDzjYb+hGxfVTPIdBww5Tz/qt+S/YjbxNpuBP6eCB8RPeLbml571/A1RNfpm0c
s/UwCwFAet4zJl3QjKuUz58gQle97QEpGI+qTO3wEX+U31P3Y1o/JzWIyV1zRnYBvFKTYUI3rJVH
MuPWuhvj7Ss912SDK4wDAC2BzPPXvhVn+2a3cNoSgnzVv9CdOTeM3Qq8OaN0/UQF2OwcG/UPwn9P
MguLDjiFR/fpX9pzcZ54PFqrRIDL9tiD824BuPPxGgrbfKVYL+YzOwRw14rsFGVU04NxGyuw2my3
sWJIuPy1b2Xmbq6txaaS8PdLJiw8+3s6LR0yZiiGTVDg16O2Rz21rIh9REMlFwSr3Qz5NgopBpXZ
vv5AgsfEWzEwuyTGoUvfQvduOE53+9slR9Sbzrkb7lFVwlWaY6Lc62afXzf128xcRlCYungiiEsH
gITURKE0XtlNxP1ueIlvqJGRw8HvZ3kB1F7Z9tpOJhPQk9v5aUTWKBmBT541/mYI9rvgcjYNY/AR
JGSisE+hMnK/CXCuiMGU5UhxLvHfhJH/PGHzwdEAI+6j77U/nAhyb+Lm0xYgfULNbPBY4xeCkoBc
QrgNgIVoyPvzM/2A3A1xxtApXeDfa1LpSKuY+tRULCVNzLB7rq9m/4mk+7g2qGFdkhD8UuBlHL1I
JOg1X+lzj/aiwttGE9MvxFY5tCbqFHgavk+aDqQ6WhcaTtV6LbhSv4mxgmi68LecPxcgnkHud1o/
nwcWSgr1eohsT7evNlHEb1tFFS4iow+l49pJf1Sb9OrRIGF38vXvbDPzNBUknvYYhZ6ZysgyQ7jE
ze57i2G0LpUpGxQQ7QNhYuIOQNlTTm1QtVFVbkGmNdj2JSpZm6rbE5awQnxX/5GJfye1lagxMrNK
oaZ3j4RvYgjYcKv/Hsvitu71TjRPzbQO34XcKzhBWGcHq0pOYIcqNYfg8P7v17a4wJnPh6Ih3kZr
bCiH8asqqM1707ojAk/fLE6jhmqxhV8II5WOVr6p1ASTVj3+00yajUTYkh0EE95zAaYSLWoOfMYy
40q0w8FIZOTu7xxGfHa1MTa/mlizD8d6vN9kT7LqMgjL6cZlzrKHejhqCF+O9C/KJ+O3m8GH9qey
4QPCXmcf7BwE2jYuk/BE/AI4R4ARO2MzS3tRWoILAIKplgmJRbb7nOxBOK0SjcjwlxctQZrQlCMO
lrZD/Ll6BxfJs5j91JRiElOT3IH2nS5DFGV2w6G6E/TqmlWZDKBHv24syQa79a9jSfVDkmLSmTaT
BwySnHADUAWshkPhqwGyT/Gl0pU47Ssf8VoHP6nwLfAfsuBY7eFbiVp3rnU0omDbapMC/Id2B2hy
UThEg6LBKHlkxJdM5gj/2uLsCaW33FqGSIfvwgdRnO+8EewsDqmw5pyOrTPz4JJK5oCfIevP8C8Q
7hZEq9uguyR8k9up1xXBVb+CjflJufFRg84dI9pePABogDcI+kLTSUOkS5IEHVKtFrfxLTeJz5vB
f/LuwhR8lhk9m5cQ38I5zs+LisE6vw7d+2FcqWKb6deD6Q6uAPimuFJYXtgS9QZoHQMwqAzIAG0R
1nDA+hUrrXyQMkp9Ph9Xzfj3mgxXMGOmWMG974DxrJaS4c0n73hF6lVdl0LorxqMhlTykPtii/Ja
oPDJUJqCciHfauT+PKScVBl4ccl0L8stW3vQC8Hs5fzEUIG9ml63TWAx2B2SS8L/SD2oyEw9oGcA
ZkQ2FiWAAawboSsjojv8Egr9zMoKwGwk5J4/gwy5TqALq8ZAGjU07n0OATMhWdqJR/3nIkLbv2Gr
bCSsUTQB1sgzLADREGcm8JxIOMK859/HfUs1/u+a8gNiVm1LTayZcQT8du58TpS5uMfu9sj2EJX+
DU/e7YSMoIikZdBFE4giAuIoDxFeMSlEb+hI2whyKrPdlEbtM6O/UkksX+wrzpNS4fm0o1GK5XoP
jm8Fa+QlvSPt7Lk3Lc8C44vo7IhG8cMRViaInoLi6SFs58FPIxDBwyyJun+BBfkwSHaAe5nRWL4q
fQ37ZVpJt+27G25sdDGS0hfz/tOgB9+0nJr9TauCfkefgun/SvfR6S1WcEgOeHA+9kByp4d55Cc7
Hjq6z/mJYWSGfmT0uu3fBc0gG6/kzXxzH0y4ynSh98JZhp2wsmdKheI1Fh/Q0qstxAWM0ysLnhSB
w/0wtiU+1HPLdeN31QVGMyr9LvMw0a4SEGt5uDguhPiQCFEaH6CZzevrnyT0VKZKxvC/+ypOofpE
lxBbWvGizHgrujIiinB8I1Bb+tPHsAvvaISvCXE5FnrNtxc8goTTWwHWNC/U/jBwM9Lm7qd4hxkf
vgDv/petowOUpj7AIemFTd7bOrM9t79+dlRCMfpSbV6MSY7oZ4cFtCYz/Lwf9Qa3VceGq1bIkIjb
Uy9KcCanQAmyY+/WwljFEc0lRq0QZ93uXijK/BmJ39CW6BYifXk5PMJXMTXDS3HnZbtRBL1SJDiu
tpjeK/j+AVCLLab7gs9p19MQLaHXiJwccU4+0jIP/kTle/Vnqbs3JCxjMPoNfxqc0ZwvYmz6KGob
r+HxwBILX5YBZrA8k3l6RT+1QwDCln9PY0Km7IGXLivAztEDEW8Mzff9hWfF17FrIYzhRTiZadTg
T4RH9ytx/ZIAIe3cOtQYMBTIRtix01Ub00z7jaiDNUrRW9rgJP/dUc7DeaGXp7o7ukBrCXEwMQcX
UL2UXUEhaN9r5eBcAy/VqVncTwrFvFijPWS16VAsusQnesQG/LLKyoSF1pHxfqaRNqRjdAI+JQeM
rWkvr+YTQlLDXjvhlgWDkdlv7hKI1cN/VaKvX6rPoADBIdcURn5hlaNKp7y8zj4lqXs0tPoB9vbW
GUdF7EONoT9yaXlcxVLbqwklr3Qpn3RRN0lj2jV/Cb42qITM/sFrIUke6NylO9P8sxpMBWHeJAqd
sdACpl/Q2FM+YTmAYPyFeQS37pQKS2f7tVf6l9Qiz7NM6u1vk4sRTHbiFQ6xvdqv2FWjRvIhzlS3
8zpnUe1fL30dbrwDyZ5wNbDOKAbBlCHxWAj27li4aaRTeT6PG53unnYN8VpO8198+hIAfdiz8mVa
hlpMYsAW/GsJ9lH841Nr/n4KM2CIJvwqz2Ayi/wlxRtW7SWbURkvEsmmiasO2IjOKPnyfi7xTnIp
LI767Kr6WXt7FVBpzIK3WrGBS3UcgmGGs41HimmGC71R8LmitZ0sHBiHYj9b///gJjnhdgSBcKVj
S8eYK9+pQqQwAnHhEi1RXW+oBgIUCPGPLXrt+D/G4AU4LHgC5A4ZMwY9vqhJV6J7mwme/uTRpl6v
75Vo2I8gQzfjgA+IN9sb3JLF5uRFbq4UlRZ+rY4bXMy2jZwHSzEDBjgCFtxczuQNmojvd2MIxvIL
I2DAJZfsLuDIGvBqmM6QOrvaX9grHurDuE9Tk6grzk81DMqK/nbDub8aVyuzEnA0vP47pwjc8U7F
fje8WKBQr5XsipEsjIa3MPKR7T0OzvBWcEAdaDz9eOexRNLjuqsyIts5uTRHxQ01viTAhznsUTjK
mbIZMdtMgbeogaU9c8m9ji/0RrRJMfODJHRMKWiSV5vWFwTp5zrNnLmZiv821df+4ljtQ7cfA2EN
JkHcu9yJ1wsk2+tUBX1hjvPSRYs26dE9OlrAVIKBsnSPxSeCh86kUGdex+cTFRCyYhvxx7+rgKUh
2uFUIaf/mTzSvf/vpvJcP63lKfewPbKO7WEraUDRBM5p5X0k+HiNqfD8SgPChiz/njIsMGCx9Gqp
ACIv677ANP6pUoomyVe6fggN3+SNZb8Qq01Vdf8u5ZxB4S7KqMjzjhcFlNsisEC2La0AB57TRM0K
SzJDioX/R9gp9xlOMdBfx7wkS0aM01TNYo+jF980lx4Tm2UrktesGh8b7PmfZryU6QN24yB1Kfym
Qe5YAYm9/Sv33NwIJGi4gPs0Vrf66CjTd5DB8aQZGWnLO+PgqrADv1gY6YV0IEL54Zlu9DyxaWOa
mlmpWUsc67YaYn6Vl5wVx2a5BNZ0cp3qd/dAt8btN8WBFxLi1kqwaqZ0p8cBUgSAPcWO7a5XKgTe
//bOnUDUx8OScvqSnLqGzaHiLe7NgZEDTzPFhRfjwny6YcfcrFjgIIj2cGkbXX7Kdgu4aBKppKLw
FX2m5uhjdxZwAc05retfDV11c7hu02ZBw/cMn75sQFW6lUjvSSRMwzZ76V4SvjO/jcd9uHbljElQ
mAVhoN2SOl5fxvKaHI7bHFfNxKGYudzH23uKyMWQ2ICdx/aAJkbacDnptppVmGU6CyF5N3od8DBX
0HGXwnk9HZdC2dtuVPoLXArFEwo7ZPNzE3Oi7LjCJd8O0VcVvy61xPjNSTxZTBEdS/kbQAC/agdT
PvOKwpa1QbyH5y5eGlFa9IwqU0llv9f7KczcgRzeZQnlctVB+HxW1B/qOPxnLHzCp3Hou51/nD0/
pqU2letC2gAqu8SftUeB3lN1BmWZpPjpPZUZZ3rq2MtLTgodlF+WxDnSamwzdYQfLCLTNJxaxDBx
U/8ubyuQOz+nlR3RMTkN6OId4q0LNO877+AIhgFc3hiykKOO2LgrCicDxz3khW84o02JZT4VXLet
vzapQx/jGUYXN1n3a0PW/DwTIMyy8itAQbzOGCzk1bwPMW2er0FoVcLm05RiYkkN9Pr657qJf6ox
ut1Ox1RQ3fgz1TIhqMA5LGEFpqXuBGiqbtA5XD/AznOH975GJKEC4EfsAaomFX8cWDIdUaQnxjmj
iWNR3VfRcz+cJAt72ICFFV3Wz9RCrwgfThho9oJudYjZbC961r5YNhunpXI2eMnCKm2HAA6WwyY7
FTYjkCO61Vt153yN0jowVvTWOZNIqf1JhCvUws00zj9qqItYP3+AX6CpGSAGnSPNMCkT9iirHXbQ
2gmE4t+ptPq1a20PJ9COg7dnzSQmFHRjbH23su/xJT9LqJkdlIQk2zRWuXCX8PaVKXplkD2lquoK
as2MemLoy7MZ+HB9WJNqbtBlAUrnMrBMjGAamByN6tgUtoetlPBwJX43Gc/IX965WAXqN+Fp8xP+
43Q8i7dsTYyvg2QvG4Ui8tpPDyzthQCPpw55lZlycGwGeRYJmqqzuod4yVbSXhMMBahB6jUEDwXF
XQkKbSpcwl+zqe0CMAeElakl0i6VXoRYmBRQMSJhDc8Kt3QAEeI1YOAs+2zEcHuHVqE9ouEudNYG
1eAkOeAaBMvh6bzQIs9MVlpCpCFKngsGymcMYYNIK9tXdNSWZmvfevdt96kPFJ8vT1SOXCHSQZeb
/8RptT+nvFt6LVeqOaRD3eR3kdl3Dsx2Tj76cmzdGrZUW0zcofh+O8M/LS9lOWE0eXN95yt0ULww
7EooJWsHiKoE+GHFcCFMIWQXzEy9vDU6nS9LqJSYSHkWSh7c1smKSXyKjcN+T1Qxk1Vw2gtdUwFO
DTpuxvBXwIZem0LZysMbgEkfQu30BoQ78COrNCNcYlsuxJUtLd9c81lNEXVCXoVeDcSxIKS4ouQU
poQeRIFt4UnRa0fLyt79+PcaPjoESB+Y2PE3ENccpZzoqrkomVYY6rLC4nOZbApod+cV6Eh67pmI
T+BZEzO3QCJl4S4go7OKZAiJpD/ZzFpj7gOigexwG88GLAmSI5nEqZPdINIAQhkVUr2LAruZc86Y
cYzeTLp2/e87gsurQBTYp8u4dB5DDKxqixMsRJ0WxZXo8X41GJ8Y+5oZTqu7EiOzpJFhYoeQij5a
woVqiGG3XLTQEmJUjmNR5eHtLZqRmbbVIprNyN9UHJhp2eiCtAo9CUcjdSD+YV1+LAk8A4JXZxVo
GtYV4DSRZ1CSjMNuN0ztG8CcnfxSwdI5rezPr3v045Z1TiydnKP2c+7XLyVnf1JxTewQVEm65aKJ
RaC9wnntcGwUT6X3pZUgy4RVsWQmEfaewZXdojlziJZYDGy8kI5y5nM+ReeyxHlYY/aeJjAAMkuk
fRVTICi5t/DK+dE0kaiFTbwcOWw2dL700yuULxUXtrDUP5mcAIIXIXILGEI5e5JfuVaAjCASZurM
v4dU3S0B3AG+F4FCKLxV6uM4Djdrmvv/DaArxQEEj2INbJwmyaF8Iset0+U5uFW6kH0UNyHL/1mP
ZbMP9qUmoA1tvlAMFLorMZUKBxYWu5nHPNDp48v4jAiNR38JFXWj+TnGlsuafyRt0pMF6CZN5taB
Qq7+ROaQc8SzMSY7AWu+pLjfKQ0opz1xLKVUxObR9CTxzNA2POJIOKtd/FVjEaUVD9l1lHeXvDpI
GqA3u+G2cWa2IEkLokFMRfvdKdhlE4BEnsyYr2i6/AdqArtkE/vWlKLgpFziQlu/r/peO6aiZV2O
8bDMTUxp/6sGmbACjFGvc7fsaD46iDvbuxlgScd1LaCyrGb2rkf5sSKoBFT1VLsJt3FKxwik4Bgc
8kZPip/sqP3Kihu0v0pCUTXS6T2Sy02553fifZ9snO2/HbY/TXEZ+xMbbXVjw2iHt1KMOspyw8uS
wIQ9pMOQ1MpNMLcP8bAVyF6wqhcZ7x7p1FcbHAUEcP74uFCJalwUPBTKz6Z38QgnlT0DDM0yZMHz
/Lyp3S+8QTrndRz6YqM1FO/8lz+D8B0U8jg9Z4+aP3oAO3obz4UQ5MLLgHdo/qsbOlZUOvPgl/Lu
SdrWtCHv86vVelv5YZioDpSZa/C959vWt8dY5FzJ62++ZQYUwpJsXf40+bJPqxUf+kVClb01dYHY
hmh5zoXLo+12IFvOnrZ/FeoMrmW0zH7nLwOm7lJRDJcvnpxKyGjko5DYr7TPlWSnBcxgY24iCiid
Vjsdq0HoMn7goJZbZWDHqAeRgOkujKfIHS773gmZ+b7u0xEwq7KYA64KbRD2I835lv26h0Lux0Xh
g7P1tV7loVe9yeBIZOl+ghtcQfya8xQNy+CR3c+DyUhBkqyTSr8X6If3+lJFfG+qEePvs43byBDn
z0JRfKrZTZRFxBWxFQ3QXLhxk3n4xrFBQs5j0erCaeoQLvdD+PlXoZZsXk5fT1MQFn+2prSc9I7K
rCsWDABO0nq7jBkBeDHy0w0LhZlZZWKFiJRmUAOm0XgX6ZIGfkj+64CUNlOj2fxmTIYt6VOII19Z
DqPoTWBEZy4QEwzR8dU67rukIEjOl080cGcbWWINMkiiEWlCSFShF63pNFxJvlZd/OZveZa3hgXg
Pr6urPI9otJDGDv9iEtEFqHKt7U8Z4ZODmPb6q8FaxWJuBxaUOo+MMhUEi/SEqU9kRN3dr0oc/lp
Fteng4BL49llA+a/MuPs1Ck2S0ksZK1161WN6q/o/KHTWo1wtAwy9/ldFQHYVjsfnXmRp4d6ABVD
4WHyrF3laqRH9qdjrVnhPRaM7kkZMV37dcBRW5d67tn627t7qPW1i/luL9V1G2z/KTobf+9Egfk8
dKotneAkexQT5qrfAHUfGi8GWSh3dCEVitVcWK/GZDnmtEumv+Sno/Z//w2LhcIQzjjulaIcOU8p
6PbQVdPSrzt0km80/T8POsJxRgeCz9aA7j5QBa9pp/mcqX0o6aUIV0ZWG2GX+G4VWkMwkJl/u8qz
FWSn7aRtMG3QOLZCO3QLPr13cpg+M+qS0V+D2bEUTRmZGYrPOV+YUJiC+sDb523JCc7WfA+1J5xd
quuUzPgCAMdO4kIorPUDLKLEkOc9SW8NhGfXZonmmwoJbgK2BUGzj77LVushsuvk1Quybeyt3j81
7nrIEZbTURm++g0t1+HoFUV8Hfbju4rzpHvhU4vfPDOpSS1srWgyKAPb0OGlLEYRM5o8FjAg6aLL
nIj8Igt0Ll9c1WmD5f+zjHWlv+FrqZwrwmBVXQO/Yj3aSJFBIRKjPGPPLJXnIgIekL9rxWXmi1V1
vl8J1+j9WIfoOy35IY+jacIrS4oWustb/pb3F4ob+V5fK8rOnaPOG/Qc7/LrkDepTU8eL/T+0oTw
76JcxHvwv8qUPHTWBQn4uDMmOMvpkDdncMVJH0m897psB+0nxFkkTjYCR0rNDfvl6lZKrv0Uq5QK
W+MFEjMwTulvduOuN8IilUKIHVl5IH7DdGKXz/v+/l96OVtzQCAlkBpGK2QTy3c6ESe26HVG2oSm
o7oBHg8czmMqGdbMlV/cXwB7KqW71b+RkRczj5Htzp/gXyVM+OkXh5PpwtofsbDyp7JYGXlFUOSf
cFU9uCyQ6di3qdPxMlIo4mXN+YlzFpo+TcOr7m5PiDZZn72N1BH/tlrQOTyWu9S9BMTh3qtWhkEl
UehXNbyTtVjtBbBd0JvudoojaYXsAsdErs7vzH9T5nuXXWJ5MVbtrSc56E+88kFju/+xVuWbwCda
WBs6sqryP2UGv17Bh71h1k6bRxOmSl50JiX9eCli4s68UPNyCFLfcX//yZ2x3Btlp8qHBBA49+TP
vxg1DJwZ0TZXDUc3iAL+Ze2UG00IDdZZzi9GkOVjfMb8OtZ9YUv/NQwHLmZwWZ1tXTsjfTUzT8iv
zcbldOxCTDCbuGJSfTAZ13QSSt9gGviXgqrIH2HJBgtkDRytyyt3s0Gf0Ag+bMVZgdyVVLtW5wFM
Nck2ieOVgk88njDbatlHV1O7QY2+fVoelULwMzEkF3HVg3cO8zMIfgbvIS7RDy0Ct6iKfmS7xtvd
ESMbsCBEfmS6RS3P02EeG06qnszUyeeM3Y8tl2QGce33pbwiV/QpUsRufOS5PPqSBCmfGWOmCNUL
r4a/o+a2wxgkcY1RrAq6uudBJa3JJ1szMNstRlXS3xfbDHozKAsMDbReKthxgxc8AdU2nhEM9Jex
KC60/Jxb9bTmU0zBtA7KL9hXlDK3owzHha807RhBg2p0WWNXByn1U+gaKtm1J00D3NxWLsVSnmra
5nQ20mY6TXC0tL+8w1dPv6Wnc4N3W9SYzAg6w1nqaZxv7c+8RgyalKa+VTMvd1L0qFrUio7Eo2LX
KQFLZupojn5bYBv9K6pKGPFrhCJXM1V9k1xq/IH8sBFRDXTAi/eURSKk6SBtW+u4f1KE6+JbAUNr
EEudDBoEY8i1jeQ0kHo1z1tE+6e9vnsHLF7BMqWWDQq8AjNBlOlyNqIL8fmNZwO0i6rbo201cVNM
iurSHJ91dUOQ5qHMYrNDj21vbzGP4FYw0i6R8Y6AepAVYA5+sd0gg7suDGKoic9fzrNofh/whGH7
/U8iukABl8ogMYT8N4VVu9tE34KWQcqX3Xy7ox3tYOUBShLzk66EPMsw5c6USISWgA9j4NesQ2TK
PAvdgTiGSERCUGkRWcXIxTnXn4C23znVK1OfWbF8i8cgJPfU8g/uPyn5ytFlvhkCm+A8MSdhMTxG
pdykNIwJMa65am2dpQmbiZR5bvBqjZ3rNNJ/Ez0E0kKJB2NC4kbPcGBEbApaqf7y0JEoTIHi7cKG
YnjXP2XiAQDgr6gNH/+P3G7r1Be3Kn9UtJ/gTWKSvUaDwl/XmtAqtvhrR1voU2GKmheGuSlBIwLD
/1tD2kjA3koXj6e4nzRTFU4wWxsH8ob+ud0WPHd1XLDDaPJ0TgzA4pEdJAWGtzI83VoAXoYnNJwv
2BA+GDPqrMgl9uhMZjZ+SrX9X0VooEI7RqBV+OViLivuR+RUgkPnIh7jz+Y9UuofugNQi+EkPEil
vLBTWDSLIvYMWBeZadmQwvR428luHZJahTreyNxuK5EFC5DlYE7XSX6WIxwPUJ6dlX/B7ZsWoq80
Aldbx3Z31EN1hIjpigYeYSdPyO8VQK7NsvK0vURTCj9wHdqTvoRH92H9R+cqP4vdPLQXwNoIUlMg
h/xrl61Tq/x58y2lDe6b2uS5bk0RusRMApbogkOvNyNStBYEJQ1fCoWHT7K2ToADLoY9BRKF8Zpn
Tejqng0REBY1v3HnApICxYu3uaAgQi6GmVTKyKF59DrDNi0PbtO1YwkzERWqUkdHqV+Sq4pEXog2
j0SssEBxG+ru0gHQdpHJdafVC+yfNrJPchRjeCVr0KD+RRGocefaMsjJq4NIIosleWOfGvvTw1OH
69ESttXcoNAUhU6WbCSrz9WV3bqgAE29vxkVYfZXqNpwC2eDcLkEbj2NzqIaw5kPMsZ0y/+hBVK9
iiTZXxvvvdpRJd79sa8LftPMaqipEvWjPyXKCFsIH+GZg3VsiaS4NlcC+IsOYznKM7sYzOza9hnE
tKQs3vmWhrzai7/k3pcSlbVSVDmdQlFJa6eo8uGMUrW41njILxCgUrMiq1dc/zDITU9XbLrJgcrI
b/ZsNoZ6taUKncKjuI8IL1XNo0hoK+kwb113/Eu485FnviNZ5WRTsU24wsRfHeqwhq7zNpJX4yYq
dChC60n3IVZ3pDzoH9Pk5L5FsJ9fkYluGjy0hYafJxxuk5qIYOW8OIYZZpovorYAL7LsKqVasG+1
IBX/9aTP922gV1OnyO9m3xZFd3BYX07yIgp2T1HC7k6a3jhdPsHilUsW0ZqBOD1g5JwYUVF1DH+N
bVRXOhaIqinN9kkyDVL6ysr30SCYSRhOYa1m1jV8Rrpub0OHyqwl9jy6+U2+lVuNFEwzRC/RTElT
2p4IcA5KkwZrKMDL6PyiRPdkMvbeZoCMVTsTD1o/fYKWFeW5O04swwbaNxFLZuwwrWEJyR7umNkj
cybJl5LI1hzN+3zV6+7Tnmg49PkvmxLt1SC/RB2ekE1DM5h6ac7/B9CKWef06I5dqiJ17BmslAOX
+TBi5p2J24usYAm+6IgqfWgC2SHictyIwc2DoUyt1oodxxv8IAYy8tiCYOp3qyVUVtXWr4ngsQPf
6vptRyLFyCE0s69U5bShpsOP3HnbBO1D7z2VKoqlBhXdcKzu6aMjhdcBWRSRfkr8anBYNEQYHWzo
BzsMssQKaAspEKdRlNpqocxMihFgnIHiXcx4d4C26VJ7IVfyblduVq9Reri3rMPxtyHmTVS1DR6r
GjtL//ZIRRrYbF+eo+9NXQO8COTU9gOLTUU3wvV/18Vn2Pwq2oqgjCFyLSj+rBjDTZnpKMTZC4++
Z4yfa34y+jnggoMU9fLw50sSBRpNpkPZrBNUPrC3BkK0aMkG8UqHYbvRUNOyxfOghO8jzEINi0tN
vhiLzfiHAgrl/YoNObPbvNP/cE5HBzXyaj9vjoVhX44RQxb5PBpxP0hg62YNtq/uEOIq1XRDXvVN
Tw0njUi6ps7YGL5Ffm4y0X5gyO1r9Kn4CS9g9F/q2FKouMRd5OBoUZZBjJoKdGDc7ighh5nlvHOq
wloFreb/VG57cwt0oEt9QF6+16daRskWiZZXrFvEHMA0WTx/ZlDDig5meD9y7e1PEaUnRRb6yTGM
776tJFob1fnuZjHWzzlq0ldjecIXvajgtWtG0hcUJWRLKC/zCxOmw9lRdNpTTUeFWS8SZqDwjrYs
nXIuwktSfQ/nUBThSUWUv7fCPrrX6x/9qwcSUHftJ9hXsCsXq3PDDL9B3ACxudQAFP5VdCUaNZTF
jAYOsZ4yEPvf03UrgwGV5F00tPmICYZNhG1GBv4OE/+jrg4HI+YZRj95QIQYWZZAXnvTfi3g7TxO
dDJ3dVOTK4HceZ5ZcYdk4KwuONCFVB0JqNBweSb7WNE5O8Iz8zjBl84B+I+LwGW5h+JrwO2FXyBH
vDTBALlWk4YnPe3PhfFQrIzcKm/OjKbVxusWRPWrDvzqdU/HE4wqfPkzVY6TgduYpVxA0d4n1LgM
6cKloZZhK2HODCz2A2cJgmhknW/TuQt0/BqFEqROX+nHeRxrudEO1Mt+xWTXjB/1th+x0SNZLd2L
LBVPm51ii2S5v5wvCl2vKOvNxdo6QiZglcBABroq6FSXaahIZfDcnyFI0YF6RaWKU3XutsRt7Zy0
FRMmiSl17iUxzhJG0kK80Lz/JCuAqNZ98Z+z5chVk3xLmtQ/OVRfZ2YDF7TqrP+DU8HxWx5aJFPp
OqkCRTxc3uXtM4xpQizdY8odzy5Qg3YzBjC9xQ1J2142632Gpn9ehS8dmc/jq2An4l2EaeyHSWH7
Ab8qndfY4hSpuR2Rn+k71rib5EXLLx4qllfXCAjZacjHnRVDc+l/D7r9l5l4j3+E+3sxAEAhu/9r
EUQFap0j3F1EJS1lFZy4Z9HBm27lMX4EGLaPCA8aQsMHX/Jijx2klvmLxPu9tUZuBNQtOQdpVa4N
7AvLg16NANn1UGt5d3MoA2XJsjDEcsOJE0ntk8Jr5VXUZ7c3+5Wdy1yraEn+ZwgZrVY77uprw7C2
IKjZadg0Z+iV6eWFgMGrEzxnSpVFpfaTqdz9XCQSwCNWJH5S562f2dCXr1EsfyXHcBbjN3oqvzzR
arO9gPTrTHLZtaLwrVbFNVOTh4GMOCwOq1j6lxdHFSKiVadZ4suZuKT+sPxqQXR5kptzwnfdCTly
FEQI/Pf7uEFLn2klomh7hBugu3JPK9uYLTkPobOyNddsZIOmEteay/WQ34LzdxP8mhEx4oIcj4c1
+l3A7LnYPfKBOm3GlvqFQlqh9Qrf4gwgua5Ab4Pt0r8lyfpEzRZRa3CuwsEJWkcp4cuPWFCm0yaZ
5ITgVcQJaUr4FN4+Mh3K3B+8AddU51a3itA6RU56uhtRn1jsWGxfUe2GQOrcTVTua8bjZ/cL+CXr
VQeyqssfnS3mOklkxHnbKFw51fi9NbFC7EnIunDwJBZ1evuzFfKaVt6cirf5A3+LrmG+5KkWcixB
mm5QkjoatYsNNu8aU0Y9n1i6mkQYpUk+ac2Ep55UuJHAyLduBw+4ala8pOeOTUT0GLJFdmzDPtdX
iFCfN8BA25sYFIt3j3buvePAuGwEoyjCns/zde+Vcuy7c4V1wP3MQq6//aUTPOwRTLFSIYtfxM0G
8sNEpUbREGO0ucnE9yuPm14V5KsF/QawN6O6DId9aLYBr0RMlBjm3M7T0rOb9kEPrs97lhVT7QhS
gRyJqsSHlpakDnKWEYnzwtOj94pwNg2c8h44VAnXQ3mlKXOhuYPXd7sm4s9VA7MKs1PdZA/8hwUH
EgJ8mGE8ro8H5JYZK7EV8/IX6VD/BxXHo25JXtfhe2REx4+S6dE6KA5P6RoL75bgDiQWuRH71asb
CyAMyktlw0Zex9y9oqAV03jT3twsxmjwJ4UYh0+xqFmxlUB2vOACUkBtAbnOHN8azr0qTh9oyaR5
hSC9ktCiAAOJHTyw+S37Y5HBdSRnK1GG9oqMW1cjUvWpWxHQnlQbpCyU0HLTDWJhK4eAkBnrvOZw
6PFoLmIBTL1eJ1hliQqE87hIJZbBjapBviNEosZFlblMqnUOjSn9sF4YJTjG6lwoxyIPF04pkr9x
SEpwz1RBdQoe10Xd9a+p5mu9VClQPOf5BqsjpcOcQq3JZJ4ZMuN4QhNDGa6KuMEvG1L3H01RrLDp
E04ACz/aUmUKnJV0KdYVo8PCeIRqM2/hhseM1CV+X4m4qD0Ib7mN0xKMTVDFnKzGKsxKzjibaPLw
GOBzH20664ac0d5+ocpv454qTBz6fw66AF4dkvNGXO1nakOpvA93IagPVqljSSGQL57GZy58mlD0
ndVRqNNnCeruXhpz/yYN8xSEDQUaQyrssysw6rTboEcDID52AoBSK1zQDKj86UyFteKiHf7Utb1c
qMZu40jBESKwPVCXkIpcfIrj+3elIHEBCAgnLl01x6V+Ink9AygNmnxHqPiqyhr3Ry2XmWC+yrkw
kzXNNS7ksXxq0KnFKLmYeOKNy3QQJfPsW9kiLxrw92UnP9xO1cVdFc8dgBi3C7Ulhdhm0FCt2dtv
UVnSWhx7Sr+5nqRKavw2jRN5ZeYy5NPvq5U6SnW6R94dCpZ0PofQyaPRgfwVq4a/mkKxWPibDjMS
rto0hHBB24x6ct67ZRKgpNxuAKBHhxk4/RP0RoGnTitHpppL1xPgnCyIoQoPL33nNroZY/z729Lp
1aM2nzA02GwAH3kIUBF1JS/wA/tT48tUgc3Db7Y1X7XnSuQYzZwJYTHklXtrt3T2KfUVhmwJGMU/
mUDUJiuFPe2d+YwD0DzsGuM5kweVjOlCfbBm1yn5HxMuV3Weln0a97+MIOJQltDTWZiwhl0Zhjo7
s8Lh53zNsxWWbb5ttGdd9DYcxxp8a3+eRUfSFlcpcx+ShURXe8LYjWyQFLtAvgDvlVdG28DXWVGa
ztZhKPAoLgLY3cTRTIv+sXZwq7njGcRbMBv+lW0OBWF6lKibjS0XqZFolyrLbqYFMFuz43JB8O0F
2KuAiEELgRfeanpl28omwq69dooMw/nxdy1Gw3uigYbJV5A0T+klt25tuSCV5EF2AzkAe7zKLl77
7ccsUG7jYP/ygqZMjhuo6uhHV3VT36OgLxNs9otnH/L0Y0Bzlmtrca7Q3wWZNu63qMtlv4jNj+B3
aME6Xf9a41wyOXz2bM5RtNpRRuVViwfhx0WvEFx0utZ+lw3LBdf61bCBbBUSZl6bkdekZL82JK8H
hsTxMqMzkGqHnRb0mz/RPDRz21YP+zNr5RrPaNtaq4j13kOjuYnMtKrcCLbQ1l/YAxxAfZ34Mw/a
LH2Oz6dE4iZpIwQWb4iKbsXan2R0w2GtvbEehLvZ4r0CbeVMwDTN26KGTHcVCceLjbXnbcI3C0nA
hM4XhNfuVfT43BxjWgK4KteANM3BT4ZYJ6yZyXoBAv55ivIcGyHgr2c/pFofRTO6UD0kRFtL9o9s
gbSZQJBb6dYduOagXqiSWmpz0xm0I5/yAi1FC8Y8alQH3o8I61pIb2QX9UqxTEVQlljRy2mpk9V+
sABnwHvKWqx6nzZYgWOxvPrZz7J23N7h9q2w602ZZRRH2wQnfSrEVTWJSUZ1ajh5RcGqqzziic2e
kE2GXNbNt6EdHzlH9jLUKAJENTHlpIPYHynR4VF5lDCPQFIENDCwjVkLFOzIrko/mfBdNp6BA09b
PHOzdgCgYPeED3hTUychA6hdh1FeI6TFsO2NgIUd+zQIOAkxSTwCoNnYYgpN1D1r+poCR+YL8Zqv
NSSr1pCICviA3jGd48MY/InHvqxvcFIk8uipVoxxRrYW6n7z49lnpre0o8SCShq1g2bXO0Z/1p1K
WD9EsFe/iW6beqvhh2EUCGBsKCNtgnuVn/AyEWflpjvwHK7PhHSll6/GclFDMQTlRM8hK4NhvY6T
bYXXQSEsXFqp7WAjQT0XjRSMqWgTEaINOfW9CgBlCTm2xeABzmY7jKAIl4DNF5qJFAWU19yV5lN1
RRARXwsH+quYYI7K2GzL6J6TjJVFtFFeFzFTz0NRwfC4DGopu4Q2JdcN5afDfrsYG/Xq8yfNp0Kz
EWNGRpEPNXkyRDtgpIXGYJmga4SiA3wJNHuZPrv3YKi1nVBy08eYWoXNsqGeRBVOzdeZUvfz8tPi
srZt4VEhzAMqfrxpwQrLE67zD6Hx9ICcLM547aqJsfZ2GIS9XXOV2XoyPnH2lLsYlnYMELs3sSX9
JIF2S69o5rFcBGjHSYMlP2Rw/VGuZbQMqMINpI5JkKzHYCct3CoXzT6+5rxLPuGwMJdSzCQnP7Qt
IqihveYg+1xuHO5qnBiyq1nU+n/Hy06BqyDVXeD3zxv2f6cp+pOalHljt9XHS6ho95b2fNqrhMHe
GHrbbV5Rl3uhTyOWD0mS7kWM+RQj0KlJ9V7R3mMy9JYc+XQiId1yxiHCtbKLQ3TQh4D+vfc1+8xM
WWEt7bMes1ceJ/Syp0pJiZ/KpLPfxjW2msnM8mh2x9EaUm0wtSljJOjC8P/dA3sYmWmoIpmHNUrG
h33ayWkUW/mtaqD2C4IKz3uIY0etZ0o+te8vDOarLJyOfhLidEvHtYyzPAuT1uj1PtyP42tloiWK
jIVyINtuEelBtnvVryL/sL5831DJt2N3FcJm//CY2aPwqJds+cjM34xbQtWFkRveA3zI0YwZVO3c
MV6LBflkawnF4rmyBx9gdxloPipkvbL16u+wE0ASnz3m2dv1gJxhFmDcgEmoBz30Z4gnOv+1c4mp
YKizTQVJDlrUYxkCIzLdnC6PgZgfwR2o8m5GKSS0P9OtY7+paY2cXoTW131z7yj1JmllgTGm2vgs
Pvb0467gxfsbrCu8S1CS+nyFv0mrad+W9cjqXN1IRryubYUrebqaCPFqMB+nwfUw3sT+2HoWxIsQ
tmcv56WtKJE6/CPZKT5vW/NLhl6EpVcT3tOU5hwDREAhYCyPbQR6OztL2w28QKE1vzOD5GxxnnB7
DZLhfz79Qy8gg0WwiHskQbvKarQUvR+0EN7mBnqg7fYPqsLEjddLlKn/N7ii+6f18MrHisNclGvl
PVCRtD93xUvFqeaEsFxyMCCdwXbjh71XyPVtHCfzxzNzUdaJc+zBW5/D/5ePNqhwpcUgdU+k4DrI
fK7naeb+x8pec4YiubTfMzrSJ6S0VN2iAwEHYH7vOWhVfOARI7xRLvZ4IyB2EpK7x08fGohTl9pt
K6IDmQY5EfsEJZpbRQSBWnr8II8rUUHoJZCHtipDUIo4HZfb2jBzZAS3cFHt6RB3b3JKifJ4r1zO
XRS0V3spkP6ZEy8mF5yoYEla9LoSuy8PtzcWIboRFkVYKqN7Ye1+ws+K1NFWWIVcYrbFelTLmF1C
9wakcL/WH5XwLUyi5ImXCsyClE10gXqh4sqCAjYto+vEFkFhCTN6GVcVjdyVHpy0NvQaZuuRO3cS
mLmqlYOzz1kcWF7SPAX4LUX1ri1KmQ4kp7j2UtOElS2C5AgQQHIT1zdDTErylG4NAxz9GoHfLIuH
zxS0m7rkCItBx5uZ1bCZxo6jBEqjfHSYgpqrHO093nZorugv9vdUNgiTcyXhuqjBHvEfxN5mRRmO
r2QQLHZ/rP6q2A6/vvx7dwBfgbmq1HkDF5ZiXSaF3eZybMSH6m/uNXFcZpHz4ROyJe1nsqP4J4ez
TgcNkX7T2Q3UKllT/XRqFpMmQ5s7rShR1cKuac7PItdAgyC61kVOHgGFsFyOW1xXLbp9uCgz6cwe
+yOEyQe7BmUEJcppjF5z7Ou5nZzuxNTQKRoRhs2LHkgZGCUzanMtzWH6EB5FQwPr6Y7/LelN/Q/t
EE1w11DC6HfaYKL0TRh3PjBXMp7pArrthO1xozjqxL02bdRHGF1d5rWMaZjOemfR9diF7JJLwz/E
BycDb+UVoC2OVuOIjYWCJsg1AjfWu2WD9OkyBAMgnI7Zx1Zkiu/K7VBtj8aLHsExJgNol2xHJBcb
at8p0QBE3L9ddn4FUtkg6zixznXOa5cTwD4K8eVC2odg0HM/fkh/bUu+xoxEZ5933Wj4Nxgl/ry7
ESLjrnnJOnr8HnwtOjr9oTE0TX1lSbqtD6tuzmdDqdoJlO5yfKgkpKhZP6lSqVioDUL+U8Vfpg3k
HraQRhsgC/n50QoiKULrxyI2Ybk67IyX6o/REb/tmvniGdafo8aKQR6/CkFKirILFUYIR6i5vx0g
6K9Jv2HWNNp6rbK69PZi4oXAe9u65pFV4w7OzWQlAtHua7Zv796qcKPc8qsQXTvInjEHVQTP+fQl
wpRUmzoqRQjrahvJCknsObIgw/rhr606ga5sUblg2MgYgFlpnA6N0oh9s9DZQ4JE7xlL4T7zc8lS
f/nEKvxbRbUnchxhe3lT1XU3dk8nP2bonchEDozGCDajH76CQnTuYyGNQXuTagZvBPiHkRRFXUCs
0MnV7RUMaf32+oXhBRMT39YeP3W7j1HAVbBN5AxoVMiiS34tsgUSdiGunSWN2jp99shHbwYV/2U1
b6vNRRJiZGSqHw8irGWkIjm8GUBTx1ytwKmY0ghgsiXj3eifco781VJoJmFK0lk7hJaB2Kx896xc
cAfI805EGfxidc/gzhkT+EM3hvievzhUCvqmqCGywOU2aRltHq9Km3CVVhXG7fALDR55gPLxYfTP
Lo+Sda7rkwmcE/LG3Ws++MWhCMwPFYfGXRAUQbjNQRVfTwHkU2eRxPhve8KyPRBhC7JusedmEt6V
/9bD4TZt/9uHuDDezdz73p8EldsKkwsb3WeAFBFgjO0jXMGy+zsQBSMRV+pxPB2HLGbyCNOwFxqw
3j3oNpP8zkrFmbz4fFEZTDAxYH0dO9HsCwPeggg9kyAnTR9OtoJ3UM9687hT5XcVNUL3WJ+hoK32
15Ty6QxnuG3Z9mgIEQmVs7I8M8gra3QBF+0LWHRnHLbo/RZOP/oRPe9eTCes2jXRARL15qoGyASO
hxKGC/rIbInXg9SAh6i3FWixfmcKQhaogdi/tP9G6HBqjX/sSGrXsVLSEcZ+7B5miUpeOTPfaNPj
d7+H2jetB6Y0XysukuNRSSqVx8QpqJ60TNZAacrG6ak5s3vkD6bfdy3JWRFnbt1njWOd8dtiiACX
ZxWCqMM25wFXC4vN8npf3W0Zpaqvfhn5o6EqREX4LcggwsMHqYF+8Qut3Ay1wDNFzj87xXFlRvLD
JJt4cotIlfSqHOVyQVpAY+2dMJ5W2WjwY6gcDSJPvXLC+sQMCnKx6UsFgv3q3KnLJJJmMJwRZCuZ
XXnY1CIOtaF/M90KqOkeuMtHYBVTqZqpHTFzQUxlNbEB1RrZXQdk4WY2+qfZcedVFtpQTJW+u5J+
yMODnaGCxpLM6kMj0KJI6YXFo7s/xxAqCxfGqAOZ1tkKDQt1rwG2AbGQYhieFcqY98UcPNKWsjSX
GbvdBNQsQOACKKiE7Hae4Vin5xobCMTtbQyHO8wdjTQ6feji+4NQ+wlYLKQKiC1lhjhl2xFzBef1
SILItv56uPqjfPIoXqowkLCuBzsE2ggMCY2PDqIyGY9U4ZM1Tk9H5kpbQ7L4gGclSihM3ZVDbFMv
AX0cRTRTxY+D8od5AhiWa+XBdADuJcBh0dyc8ar5U3aMGO1Wc3RVRr2raoEXh0H7Ja06sbfiqeNn
ogWUmjb9gKG3OJOgwRGF0MPmlsVQgsvbNkDr2xHixgV/lAezSckmBcbc3q0I5s83AMtRCq99sTwF
HJiq3b41c5HpK0/mp4VIrY0Yg4mAh1pnSfuK84vYFqwph0cL0PTaLTyT5YR19DAphtQr10XXCBuh
RKgnncj17TJc7d4hcG9PEHXZf4+JiPVuz1Dy4rS9RLl3gnybxu/bF1ue3PWbLeZ07p4rIPWlMoFH
ONf36VnJzkvLX9VKuKUXDGIxqtfTzLYMGC/A+Bfp5dIYKeLAhW3F6cKN6B/CuUpidqisB+PDSyV+
T3HQIZIpyIo37hQOA5mSk+k+DoV10sO+18Vyj+ffje8xj2kD7r13Lds+YRgarU3l1AnF92/HIJKq
lBIjgNTa4EWTN0sdCVZWBFyk1qOcA8Dnt4WxoTnnTnqn+PCv9hcWCyGwtXWYp2dh1j7oo5cV6jYF
nlXr2YPlb4c1hbZx58Vx5guvGC60mXOt5Ez3g8a3NCT8P7Kh+E737V3FakMBt9Y4XXhBjmiKUeb/
fST8sTA27DmwZprAYbkP1yOeav2VP9fAaHO3FtLECihdmOTKLaJ+F0dkId81XKA2X5SzFlRFQPuC
eCMokt7AcSALlKdbkqLkOVYm5Gqha2bAIsLszhUT/CceNBmw5Jl9uOtKvWKUILMWa7rH/fzcTK41
ijvIxLTNP/EkZQDOcXNs0pX63cMQBYVvqm1Qccq+Ie/SiGmc0DGCk/48dfRUGJlgoif6JKJIvCjl
zLMJUEVI+Ga4dA9JqpM1gw4C6n/MqLbMHSe2NbKkEnIofQNAYFrCgmu3436rKjmkIkEIZCXozwWZ
XR48lfZAGvm6ibqh6meA+4IN1zC3scCRxUGhRb0ZFDytDZSaCNEbYLplLNfimy0cv5fWG+K64hnx
rxiAlmkA5KRhro+IvIabeulWbclRaZHKMRTc5VtaP3ifF+mf1guh3Kp2MXTCz57CLqN6RUwNDcPH
nAEpg3BGqaDNf7PVwIj4Z33ILv5AAw9ozocAtzF5oiDblFCPUonaGDni/7KkO9Shs/nA8jGhR4k4
TAZNF54xCzflr1e9bZaTknqca/hcil6edPmSAyvqH14U5ls/Xr2TDhC72JJDzyB96mbxOtfywqkW
i6X3+wIdfLP3woXSOvpG7m1Z/XwodJu+SJFAFGD/0w67OhcEMBfHZyY8RmOmst2OT/1UQQE7/4oS
WZvuZIVIvm72kVtgMW8vKw4ePD0CVBV5eIXcG+Dx8XunjNKQYJLAN2aMXTuTUTCHS9NDa9TGbo/0
/VVZE0iQN3xjf4xS39sT17DY9lpDUtUHZfz49dv+cHdlfYb6/fyypkLwRTx1lqKcnnQBb4MQNll+
c86jzMtX20Hwq/+T1t+5+Uj+LBRkDJ8UVDPBw+UuWo4atpxMeBnQddqBZT98aWlkBWOVi9/9dlF7
+19v4s2XXIOQ2ku9XARbJaPM1AHpl6CIK8SHw17lQA9GYs9RM93NEy/UBtEvK2yDZ6ZB+HyBnRew
WR8zg21/4JG/1yObJj/VZiqAwdbdLKkLU5wOA9RcfbgRTPh9eBx0Pb4qnaZiKwyKC9bOUXDokfuX
Vd5gw2+s0+gv0fZmJCBqa+VIurXVaQaMAcK563ESn+R8AFbLwhW7zyay8ZnjTs6nmYsxnfV3IVJ7
E7S4UbV/HFy3IXJRGYm9DeNIIViSzIlOc7moPwKgKs/VoZQCuMIrYKMy9AQXk1osgAoHc8Tj3YJL
kxBSKSiDptAuJ+8u9XH3ko1o4B29mWhoER7ZrjuZw1lWYG4VgEZ9cyfevpfMGgxGYeGtEkOUpVVh
ZP/pU7nsDrjBIYWUu3Cuug2Fxbcr+J9Y4dx1bb9k4nHpgBJTZ5NQtiSD8RS59ok4CXESbWrkdIOH
bfAaD7nq4xkluADQZg1kQDMpJ5OlWmOlY45b0YJFPHnqB2FTfd+KQ9DJYufDZChDFozBHi9vqHoE
sa/NrUI8CsTCUyoDoqBIX/AEJDCrHcwKFbWwzwbRogop0t9JRzA7FS7XeBxrvgycA6if1IDywUpN
054NJcTH5jU91t0HPmPN0WZ3FuwzUOMSDhJFV0lhOw0ikyJHHrmb1bdYOhshMQT3s/e7wm6XY+NL
s9DH9epQ9rnvgnmV2TOQI+vK6LDU0YRrYBqha9xjetpvO5K1OEkRUTCuSVNtoAE6HCRF1B2Oo/Gs
quiVOD1eL6s6OdZeMYc5WTkkii8b/0U3WX/W25091n3hdE9eIbDibmW4pSsCeUO3/jn/3IWFFf0s
LTP+NAzWSLW2r+B9nmJd4lC7jF9fEh9ca0rv3z4SYdGmO3TBItQ+OqO3Ca6FTlNV8JXPjglOUgSU
FdxGQrrIM9zSCskRwWXZ61tBLyo6JiHdWoT+ABVGAJ7uHSHmVMgYm4qRHZzpoZP1y1KBo4886S7P
fb/7/Ou8Jsm0hUnaXIgamhsDUZHPShCZzGPp5HwzUAP7SpXn5YKDeZQIsDRvfaUVwPb/khm+su/9
2lCcGsTQJXDXlHwUIFqJYozQIpcNz0rmjo5HnJSsWkRJpTHBS24pFxDs/ujKAcUor31EwuHz3zWt
aZDH7Mm6A8eZxdl8YHt50JsLdBtPZ5YSxJBv6WTubkbVIFY4kwcFl3KMptw8LO9qE1wNs31MK5ZF
LKVorBvVSQdfYmIH9UyDFas3TDjgPWJ6vEpxmlyvZei0VXyf0XSt6tFtswTXSP7yjLLjrkSuUpny
ip2z80ZyLh0ROj5Xf05Bee7kNxLcuCprxWKFOI31z1YJte/J2WTUZKO/caAh+hiDrnzLJPdeX6/k
f8D/o8jzrxfkEbdUYpus3YZEed5NQBFNDonLiAi1i+RxmyR/CTCnN1f+bW38wQDeqMaWp6fMQITd
bYkepFEt2luvXZ6hCI2Mk4gxt82yuGukKSQhOsMdZbCnnBixYnOj4zJNUWzhcSxEMM8wMGNrHJYX
9WgFMq8Jaq81SctzV5RkYqW1dGSzkwHVHpBKepAlYrcGjxE32a9kv9k/pFODwROBL6Ixu39etCfZ
xoFmfEXSzZDcFIgaBuxTRsiujgwTPyi4kCw27BzUendwN/PRf1wtupgiJFxGo09j6AvcLtF9peUB
5Qg1c/XIiFuPP/JMLbxtvdaoNfn11f5G92SB+SBiTLc5lJ4jfnyLzK3XJJsbxNGXmr2RtUJGv3SE
ZHLtXyOOBzpUWA/7BtLJBvDrb1OaSiMsCTR5AnWhplUfyHUEzQm8RBwgmgDNdD79UM3bCmyHgKaF
5O0M/Kp1UEm8LDwnds5W1pMis1NBigOOiXkm/OxRe0Vt0C9C6IIt8PmlYqgMbygyHuQ7t3FIycUx
kAlOcweLOPyFxPC84qAErH7rH0Pjd2nEBG3h/YY+0S6RksevfZolZXxKQ3K54AoQwWjrg8v/UrMT
wcD0oumooqcK2IIcZqHCSMJ9WGAETu8tx6Rk6z24EEekmH2YBz3ddO3nJj+jky88lMR2RHTQQlt/
n6tGFQjJB6fhYw3pAhOCvpJAjdxBqlp951Kcqdn5MxykpWWt/ZEURTQM7ZtfavukSlu4cdwPKEQx
CPXsKBrUvrmuNwzmCXg/YFjd6RxuYaVRwjmpU1q6ZQBeTH5Q9E0DrtYDlj/x4n5KLx9s6vVQNmv+
oMir8qwUz8pTJdYBrbfy7cl6RQnGqfJSu9hi+d47syPtuQKqRZM48K+LhiCL2i8Ln5iDxE4o3AiV
hJxlDPpEO1ad7vmBui8t298N34QuZE+G/nrDzqnkqcZMmphVNBpY6v01RJLJ7Ivn5SIcVreW/lV9
fTBPAY7Y+s6PRGRGi8GHaTzeUh8sb/mgm5Oz9ZXUhkakiG28ZrHePQPuBmsiDz4VLPIj+lETkNEp
26OOMWgO4+5fRd5MTavQDy9sJc5kTA8Rv1j0F1uy+Pqqoj+pylWPQ7eZRo+GleLTiQ1WcQ9Dl4F6
EW/DEb3m6BLsQVGA/qHe/Z07gW/8mptc6E/J9nviFnj7sr0x2ua1Mnx1Fp/VevdgXJv20R97kwMu
qmQS2FKjOcGt3MgImSHdjbFRN0KF+5hTWZvPc6h4CVbOsKjD/K9xsysybDw9ElsDwJy1xWlhVmmU
JelrFN/b72tga7v+3oyzu1cXdXKGgxoi7GOVzlB/7Y83eWRvDGRQ25HzNglTYnprHNsojaXXtUdK
jZCbpfx0YL59QxB8u5MugYCWunuuzz2yLh9Htf9cq+Df5bkeSXJ+0b8H9+EUzY6UKTe0hxCliYyk
H6ALmHFUEvkpVY3PnTOebsCaRO46A7bz/X2dbOsYo7DqrswOBeohTXrJqyszdIpIatkNKOt9J/t5
KR65jSKf3CscZ41UxHSd0ISXwUSTw4N180/lN90k+h3+SakuCx3xlPqWxlVvUX74kFn/rzmskWgY
Z8/hyeAMNEMpZxm43B3MeL0Hj4mzNYOxYT5yPfGngaHbmHC/TVkAZFUWESTOmYMky09xTdto7piw
g5/xuh5cESwdB1XM69ksKKdef9eJey6KjeWZK0GuV+l1hJquP45KonANbVrC1zO1PA1vl6krKTlk
eaSL9vralzo329xDdHA7cMBNEeN1tLCurTHfTzdgBD9mttAYqUZqWi38BwZoi2H20tswNXkLvyq9
JV3mXGYbp8bzUh0DqV9WZyDm45GXJquHcenfS61a8TIEf5kjC68PVonAFmXfgaCcHYIPbVlHQgJX
KpCU8IRdYQt926f9mjuRKPpoGhIHL9CIb1aahLLPCEgJuSAk8ZZbIUE4h2HSfbq8ADN8YP/YgyHW
AQIOK+VDXbC3tzDMm5mDK1r6tFKqYMtzn2I+LUBKu/mrDTGwUdJdLX+/adFda5ycCW8a1IkcYloc
25TP4R7xNxiqKUAUiVp08bmuPhK7kDHNDlNgSmgA+SASGjjIUmuqcoDiPFIHiT7LglW3IqqlVlfl
kGkDPqBnK9iL1IxpZWdXppjF+GPAivGezeYKbA1h5iX0/UhXCHucirX6vXq2olpwyPB6z7p+s5MU
OE/7Rq20DCXtiPIL8caTn7nrJaIUIiUR0lBuUjKlAMRFom0lSr9t3BBDgsYWMDsTfn3lvQIn7WnM
RZ1GAvc04id2eNGguh1ILqHbx51pQW6KbuSyorpi8Cp7wehjornlMoqJeCYgx4hChJwxRChN//dv
TGoYw8ayThlHqSXA3vYBAJbMocjjt4KOdXb39n5g9ikCfT1VR5aAXnC34u4x5URC7uONOJkjQVF+
EJtr7n1NhFDcOY01tJaYxUi97KkLKtAyA6X4SLG7QtxGEMLDrj09W2e35DcC/Q/l9aLsZgsQKV4F
kdOPL1/aV02YF8VIHbk0721/KdYUn3NXdrxURGmaCzEP/PFFPoE6Q5Lh32Y5TPONu8ThQcMjqfi6
4W3hm6MiZiB1T4ZsxfAwydiwBWCdinq/DMRVW9gxNgZyU5YY5gfgcs9vtrvm5CyfCIH786wnUyPC
rAw9nbPeePyHeUomqWnpyb77z84+NQrvNFKYGKVcP9TSI2PYxXk8x4GHBZeQrmRW21Hn2jJCGb8I
mqlhEt4Igxrj5Dvu4IpGVsANAiAxh6rg8aYZPHecqfbBVGl3VXpVHZCjxu9HY2k41sqZE/yyDh3r
IiMSt5pTq2IUkJVu6uIWkH2bTZkV2X/yvWLSiNQGUGS3HJyGHYcmnvjoftX5b/J3irH4aWmp3bax
hY5RvExaSdzo443WkB33mT+iXR4+K0juTNtqzKo5wkAIsqo/6EJyRe0gjDbQl9nu4B4kgYrZTrqS
0a0S/4zZncFFBeASpOyAYv2HGa+EyM2B/+8PFF28Z5aDQ+iy7s+RIg549RFpL08xI17CiO6umIXT
sTq3Qltt4RFsC+AY9B5fTEfJxOravwZSMdmiZQGWI0WWQ6Oy45WI4R1XhX5tk//Jhq0CBdhK9gld
wbeToX/Y1aKdWROF9K+/maNifBvo56SUZqK1mqBfui4lM37jfTWIEysJkb+mChKtSUDYmGCxiy7z
J12KVkWSRM7Ub9fa1hHGJZ/sM5kvKTJBg/klRY7McvvuZnO/NkYYKiqnaRUsJKvStjJQc93S23W7
ZnaUD0Kfj64SDskts3kvoBmb3rZ7NrGH0ZH9pa7+jZjFufz3vAm2crDRaaaVSiPvz6s/bAi3OIq3
4IgDWazBpHjIUO8ne16QvxQfAnd7Vq852sJw5iTZiq1hFWe0rvHqhQY0mdDv52kz353PNnv28b63
k2ByuHH3CNKoVRjGElheeXWBMb2uj8Cz8vaNdgusn5sorEmJfGtmIQUzZZQWXFUoXvcuTsA1v8/4
PlFwlnRvszURCxkq6zb5FOVdln1GwOAqNydiwjKootJfDzja/68LgI02wuN9VjSRdencCO+/YGag
ei/8r+JP6BzFT7uWJbPezBWf0mHe5vEBPp+ApOLfB6EPKfhjY3g1K6XxXunSqfW6VtKQIhY5ASoW
bKZaL1Bvq/ZC2JxoXi6+yxu+WMv8PMrdaKIzIvZNt1sqFSynKEtqy4k6/mT2kDKgUxgW9iPoIJXz
kegpt3XYJqmRCfe9w3n+JadcSuAQ19MTlXyHX/KjOgLqt9Gc6LmgsB1w5TwuXD1j5NrSA61yuAgT
pzYHHi+jfJr7/Uw67AEArashQy5ss2tv2B5wH+QZHiHZXaJmMH4lapyOxf6auov85zdHcbWXTsxX
FS6aVoXzsNZAjpWLYTN4JFT679z/nJ+XDQPoo5zvjMd7b/PdlGFev5cMz/JgEn6kMwOmzdXg204a
dxHs+L7/8eF9dNtTG8H0zlADxQxhYSYudAxqdnXbrtaFvRTRAAzhE4hKtvPf83DPlMpqFnQ8q+Cn
Fo97LYb6FnJZ2fBeI5JyfY1mvZ1Y1/I+b/VfoR58m9OvNwA2srLSMVd7Lovj6wIleqJbOpKRWGUF
x0DIHiS8SU05tolw9mJm5p+yq4oEz+CJv/AmNUuY+cbk/nXpSJmJ/lXfchQCNNKgnssU+R8isFsW
ebLs8abuHenkD0JnXlKo6ZVVWXH1pr54RzxbXfFYyqqt6MXjStXZuuP7U3soV2OxpGKhlPHgqMvG
UgbphCAZEX8eOHXROj304CV8eqIATHebx7/KzY1iyzQYfaP0LZ2qz4ixag+4DASRkr02htMbtf6H
RjblfDOGTlIprhCW/KbWM2wU+7E7nbICxVlhEO17V3V92dUZiXjN5YirZ8hOVGGvZWVRBfQ8P5z6
xUGR4Plf/afC2nHDmaJ4xTpELRr4LhaVkiKFL2xt1rWy+nNPGAtqIa8vC7KvvWcAJvM8wIn0HcVT
yAWpC5Mozku0SQG5YRp7HIpAm2YUaGoaaUlp3g40fzH7oZ3QmWqBKVpM9+BLTOnzGtl09I2gsyUj
k46P3Bg9z6aXLQRNuCbJGC3warloR9oXtH//usP7oEFWnMM3scVG8fWRViGgTAMTzeM8L8sz/qkU
AIngDv9VqwGb67SfyKcDxU0+U7FgfXGJmTpGFL4jiWhQAYJVGKzL5C/usG6oHoR7BvTBF8JjbqyC
wZchuXnTBupBh0hX05VQLicRDwGNeYF/azTcRjUEuET6d188MRlMbry0kJIobMPQf/UKvgR9hEST
jP0HhRcWvx85k2uJ2YSA8AbT8Tq66qVryrn16mzlUxdN9V7QHLxek+KUnFj1xqS9ky5RVbu1VRmP
jSdKvKU6q+gxwagKFOCLZFeiYdNyHIvx3yrBf4iGpBnIPDd9XKf4rIBfXNM4z/ChNV53qmZPldx6
DxTVru7yciljDvLQPIKtziCmWlvpFZORQXm/Hb9C1ck8NOs/f+z45uU3WwTFgN8NKTXcITUJ31Iy
AXOGLzD9Bba/jG5nkYiLXSIBvnaES3O0QSMQ6trqG20PRz7Sp5f5k8nO8TkEnPSJGHVIl2e6/z1d
Ema6hkzPYfnigFtuoLsMJsN1RIs+FjtyShN/DJVTP6lnh4+B0GPBuO17DZUVcNCLcrA3laAJMJvi
p/Bltj4kFeZkOHJ91oTlNCWPdBhFxC2gSG/H8ZPW4idEg1nwawDOqiDzu+HmSOys/VcT1ykOi40Q
dVplK0sO7KWCx7znSHjneTIOC11D1XfnGVpN04dom50XvmlfmOPU2+qyMIZZ1BVIpMGVuRyBm1+/
Rh/wdNV4MZZ1fR2LfQ07kpxndDPnoBopxxhhBbYF5DKNivmBesgAMfXd3icIdsG4fFiZ/pGPceac
TqVAcXdkqTSae2y8wJQC/Inj25OQI/UtL9OblnWVppw2E7IJpbwnxgjTzlUO2JvenewsoUBmh7ey
eP1HKe7RQsnRIzQnjvtiJmqjFas+RCiNh7mU+Hr27DM6XxATuRLprsbEHKfRch5pIK2hE6kIVIaC
dWFS4i2UU6v5BXQ6sV/CtByPgi5mJ627wg7MC5J+nDSRvho3JF2ykazCNn2OoPb7EHRqorSE61m/
4hknpSZYqoDL2e0g2k5WpJ6NOkUgXnCKjUg3c+oy9Z1oOyzUh6c7sh+gH++j5yHVPAj2vOupp7i7
JB22kwarcQFSKkjKtgFC2dWmYGF0+TbXppLlouKGAOc887xIytEYqvY0aULW2+9V/vtLafatarMU
I0RrLR2k6gOgMfD0W/YlMncRxhGD1lRU7A0Fj+3m8bw2iaxZ8XygkBF9teH0+G9r25iCatGOleIG
5x71k6pYVzI7crnYzagSIzA4mGWTVzRCiURtrr9bAH6IWrjiwCRKgmaCfzvovDQamIdidM8uduHo
PiBAO1TcXhlxPWsLczMWPYUvLq4XYznOLpc/hc5939OFZaZbVgqjLCFt/FfQD8zlri2/8vQrxfQS
I4G4KgfJY9KKRDma9U+lKd4idtHDLuKFu9AFhPzL66wJX6lNRUinT5iGDZM/blILM9WfyGv+uZGN
Oa6C6Vtp6sLV+nICG5qr/BTrZnXp/HYjd+flvXILdZ2T/ZIvAV/QKdUG6NOpOTk9cKokdqfKvzJW
+ig5xhjkdw+0BR9GXTyiMElankgQD2HjiwdmZ6cMROpxaGcicuaEOvWwQ9jyQUgA+ECixarftpNJ
aP4Cj3sMJXziytBv8I0SiSEiK7oV2bwkHCARy19HdXvhxzxrQOQjW89D9BPLuRNbmylboJufzpg8
A9GQc51U4odJ3fxjH6JRpXSiiPLAgm2Rj03/VxtImq7KivuQF8N/5T3FAayiry7wuqqBOHbbQyQN
MN3Rlhrlrah7SVE7pTpySImgOnMpLkVMrHUKB8KrAO/t1Z1NHMSmCZi/j1Un8wfddpT87LhgZLNf
gm0I6sr1hRCtUS2rUx29om9/lQLzgx1SgSAsKVtcGi4A9W4cFUm1Q48yqOBt6ZxnDtsAaJoDWUyA
nr+5vzc/BPd704UdgT+N/qIfhbrJ4RX89avyg2lDYETZZurPNCefGaH69BcU5ThENfjLoFPYv+jo
ZwMDIPuXEpFFp7xc7xwt4Gxyx1030hVnxxa9DCw28qfvG0XZbf5c/XEJIJp4efA4C6j8+gV4JP6z
2gNS4Wj5tsmYqOCg0b2ipXbGGzCryT+Y0r53yelt/NwPq0rG4M+1cwOalvNUpI1St805bMd3DJ8f
ozWN+HkLD1lMqp99AIT5KOuzn1LrTgXiyH9cCvI3TGkVc8kubkS3d3fYjrT//VDFBimw2CJuEs6j
axircDZNfNL8b1ufKu8r6dw1V2j6X3tH8pG50iHW3gpXbrDHV6HtulnwZNPPBeV7542dFVgGZT3D
8wqRrTCTXoJ0Hg411gCIxtuAxzCUqkVKbFH2bSXUMDpERoyl72aXjv6NI+pqxTvvW7GyQrSMlMf8
TUjTuyPUC97QAyoxodFMyA9dEgKj7QipODQGoKUUxaheJzh4LWlz++J6STuhCuQZdWqZegleWxDe
pyBONxG4MrZG5LDypafaTJXDnJFmJOp+Ps9vVr6rgSXOVGnyoPk9zYvKL+2iCIfRFftWFLMsICN/
O/VbumGMqSMZTKv02elIZBcRQQhnbChJelzAqF1fX+eFl3UnB33ECi0bMzs0CiTADEColeyTYMBu
3tFHuklVFQpXsx5EsHPNQx7gPArN2FIoExFELD4B8Z7rNQUl24Qy5jEWmG78ZACYX5v3gptjZifF
HdJ5woUWmRuQqg3vi81w18A8eFU2v+Luvd5esj1G3evCCYJZ9R3DaJvzVtB+jwN0pR8gtYtF9VgJ
Q/rQ+tviLLx0YjnPvUTfkBgqqcYu48TuZJOoWVu6TF5IbPwfcOaPVzXNuSZ9e68kDlREudLaOnrd
xacm/5wLMuYXw0B1mlQzSkDK4cwX6YaKREOo9I03wy35YGTeQShkvs8t+SCIJ082fitUa8fiiS/F
Z1EO1oSmX/cGhK5V39a5dkBZ/jRWjMN1H7LalI9xgQ7UBAtHIyyFAU2wMYykiPCv9rCeLmhFx/zb
58RqUIpyTg1O5ZL7nZcZkC3ce4ptkYrx5decKTmmmtMIM1jK65UrjTnZj5x6UCVBTOfJQEPR1ukS
EIaTg1k1KU/uJkaL8SHNbBdssOLNrF9dQ/iEwfvcoZl56/eetQi6ZzLFIs7yzaS4BhLBFbEIyFZv
iK6aGvL7bhCTPN4vK1PERIkEkIZ1kPPs9x6ZtEIzL2/O+5/xO374mCjaOenYhBF/bN3eGesWlhm9
+VG7ostBIdJG+82VEtQA23tkLoaOFugUF1o+phjYKYrsMIYtJHkFegT79CT2TMqmo+H+jW9JiFXN
mLjbs+fJfSbSKKNzIzs6SoX1Ca5p8Iu1LQ87A+aMZtMZy8W7sMxkfkZnwUu06iDJvSc3cPa1bZQT
TRxEjQkWnHHLvBOw45iZv2OxAXlzLlDpIkE6uwjlzznN76lAjr1baGlDuHTpWDxB9SKA8ZIpOoI/
gDFS/KvNuMWXFtm1va3bnyawlc0VZSlC2/Hb33Y6nKVzDF0hGs0jbr+TYKo9XknN1ZS+rgdM/P4A
29ttNBqEO3K+MX9opyPrIqJSHEInBXA7v7sMoGDadvhH0qPLtz63hs5f6NCOhNtSSqb5SKihxzkE
V6pJhrwpXNmCjxI1f5G+da14YP9tGV5HeBoEOJ5BT12IPJj8x5FqdELDNM3qcdDmzwBn/mS7dPwG
pCKVqM4pMw9cPS8gJ061tvsUUqd4Hw4IeSrhD2q6pKOa48fJ0UixwfjSua1GNIJF0DS4rZGSZHIb
kPCTAuxSSpjneuVHpdWMga/Eo5byqQGl7ZnTlPDwCDc9moM5AmPaknFyO//MsPAVRpDjv1daxqt4
hDS31yS0eDN/fXey0B2ZxPyqbcHpBxgSYzV3zoB7SvglKq7m+dORS+lQeG6eqF6wcngb+2K2VpfR
xBb/FkIXIydavMVXRw9foFRBX0bgtgNIJzszi743NSlwmMlkar1HyT93eP+IhC3KPYa8FUGwLUPE
fubVKesAkjDnjqVvU7wZSxp2WF9/h73D4TbzAohw1DupoWFs45ZRA3qFwjCk087EFfXjpPi1lYia
W6w1edcED7nzkCws+JQPZck8G4ohEyi91X+BN17X2gWKKtQSk7EZlYrJAUuxsVTRgLBT7MSjPfVD
B+Mc1hN3/9WdPRZjsDV/YFakc2PRzc81VpjyTfPnzObKouoTnrzdO+pLqEPMhMHvNUJew4r7k2KX
eb8eSm+0GtnsBzQUfBlVNzTRFhRgfr07DfTbCvBza0V//WAxaGzlfbv4VvXvgq4ibg/coz5AYv/W
four//rp68zWvu01DpCqSurKqKxLzUvXDwkj34xdzzk0qVbzh1fcBXNknZKCui/0zGueBr+rzLFo
XvZ5PoJtz1pKH//besXE0o7msQeG+NajAubYJHIDpE4D3AU8nM7c1rO5C8WPC0jY6dcMZLBeCbAZ
7Amw1nFom0tS/okuEVm/brhs+lSGdcP8oPH8AGG8wnIOqv3iH++pdl6MnG0q+XZ3ZFiv+QDHvRf1
4SbA1U+w9tfW/ZmTuYWIB8Yk+hbHWGjraOa5Xq0sVJ6oWoMZVzGX1v5mGirQK+qrbjXnkxq5LZM4
tq5L24cZ1AhsG5Kx6rkVJEe/2WKrKQE5LznHKBfjvbuvaKcc6vfwlA3yl0scBKM8UYJwnVXzJmzz
1NeG5VnXgACjaQ0hVlwZrGy8mjN40A603YX4m1wEdOGXLGYH0ajK9DI8wlMX680JXtCp+hF0Kqxy
wSX9+vyL/iRuWgFmYSBFaXCbwjiuxld56a4hUzuGQZNLWQW7qbiNBhsoDbIPBO8EIPYgbcqcmXe7
4hEnXJ0dCA/+JjQAKvdsKrqMl3UwWpCHh/vHgbcZlJnF90UdJGIgUepPQlgZyec2cFmCvJ5QqW7r
FV5BeRJjMgGjb3wWR+3y4nZackYOkPVM7W7iqAHAwBTyxCmxOEbNu6+1L+QnQ5Db/JzOQYGixaQK
QURf6kb6lmEM5kUrCqtvEXzj3zImLAL5D+rXdJbsp3IPtdh7aNxBZxqg4PxB+1MHY6PJOiswGWY9
WNWPkjz0GdED+PXIhvBdZSSsdgnjLwGOsyM0MWZiQ2vbQeuAdPzVl/DcoUKTFdr/DuqxjB8m0lzi
Oea/oKVvoJS994NswC9xzxlhRyhM72BBQHyCw4eXIoF1wgy4v4NZtvFhkQ7/UvXqlFvMIlhttIsG
FuH6sD5K0rEsyx8uTw9Lm8MZw3NnJB0oAv9pHUTNRxqdkWb6jvhx1S/PAV2aruyU2QaY4JQLRroI
w/d19J78EjN6kWln0YtoB//9+fJ8KnCoaaK/I8ckfJgT6ne+d2zpsdI83wsxOQF4ZuECqYtovpHJ
ri88xPSxmTrm1kh7LfyDbpacuQVq52QjB7KUBzddtWq282qF5O0WuH+xnp2caWh3a0OQO5nbL5BR
wnb0p3bhEuJsc1KDadRS5S3yazUcFPGxSH6ZzA7Hbave1MfNJDA489e0sRAhzthq/Wgd0MulLmNX
lPeC1v/sILLE2FSW51dk1thQvGlVx6xf2tzY9ZjdiPm+bVUpR1SmVkaH8N7950Z+YjFXk3U5uFb+
0Wms1CWi0Y++KTVaoGARIsQ+G/L2jljBEdNwy3YfL3QjPsglbBA/DsTj7o84krZNke/R5gWOeDPC
SHsIwPfTYCgpNrHq+UwmO8iXfDvCz9MWSPUfY4xsef4bMEuZyZ5H75RVp7hPD0CcrGBuYrWbNz6g
gsIXH2NlXIpW0GVa+yIH+VbE6zUP9kg3ktziC6Y6eZC3qpJNELFhF9edia0po4NiSS1zortnKo2c
bzu3p1BeJl7h3/5NttD0+HOnFZlEzb6SytKYA80bK482taLaPgkXOL53MZz+mi+uro/7fCjY2d+D
L7cksLjXqaV10p0j33+cgOxPMtFyzWBy3e9wuKxY17zlkfRovsMypVMvKOX7aLWF/NSgU3GMgVd4
ISgzDUR/EPV77pWyGkVGRHAXMR8wB7LPHMfdglq8Lr/Xy4yubkWq2oxeDZLymPrn5VZ9I9AYK8kh
XO/qH+Yepod4sUbm3KcL8PfOt04oO9aBaMRRRuGFPv2+wdssGtSoiBAUJZXwR4QbAyF17KQqiBw0
NdgJA4bKvbFw/2J+NvE2vUt9oeuExYtTsKAEkmARVhLzB3QqV1FBaeCW7+BqbiEKfDrCyRiO6FjC
jnwhpJSgdeWyolMQDuGqB168mw5dXIZbWyIu4vW/N7UnkmJvlLLMzbD/y7LkNHLpGcRGInAljP9x
85Do28J4E2xaott+679b2dGSfqtBCAlLDAnPg6uA+Ti2tOIte3tTjP2eIuh8MwAktrHrLHT6r0cO
Fp86I0N63I+pjd1bjwbQjfUV+b92b2kkIy5kDs1qeCcW4/VW2J7Ik3H5AaSKwDGmOOLY61wTv6ZB
HWhK4QxmxmpQcAmEZU+EZeI1nznj1aOiDmQMVKA/kCfTLLeCHJIFe1OUTgWCa3FtuZkxq9GywvNs
Y3tESZuJhecxPXkg4kpWO2EwOTD/nK1iOvfnof3jeLaYMUGpMK9Tsab95H/4noaWsaQngl57TB9a
MIORpPRaXDQApz1m17F7zQl0JvrRWniqGLXhCkKhoRej3bDrM/atOADt1q0jCQQ49pRRyI64IW57
h4VTltPPDuL5lYhMVIoSOU8899uUaqdQt+ms1dn3pNFk35leTXTkXZ+VTSB8jKFMGLjOypsJVW2D
KPw0DWUwPZOXcx1Rm48cauT9/HpOjNa/tFwnG0Hx6HjWol8WDR021/rEUcu2X3QEymEcpnsnwcu4
yAflICKLSpnVkbwrHmfp6t5NtiAYLN9LMjbyx/TkLaVqejgX1Fsc7OGjSxKajAa3VjP6/YoCrePk
B24NQgyet0ZpyFEqng2iK7/U5GMVnZPg/P0kS9S6AIOMYaqlmt50asq11g0w7bBw4PNEgZPh/GsF
TEVr4nrt1wq8CU/jNY2XCoAq08lbsrR77fICOQdiYVaS2kWzqoWKJnZmhhkqFr9V/quuftosN/xz
fGRX9IFBtqGj06XcWKvGOxaBC91ZQMbemJnsB82bIX0qC2/8g16rCuazQB670EU0SWsUSwueViWe
xYFmSqzUtqJm0OkfuD5+Lrf4+za78MDGT6DVekHBxIZ9kIuaLehSeR8FrFO3Cgz04nZeY8fakh+i
YFD/SHcJ0A+L5cmlWznTELoGdxIHDJOpdkPcKJc0jnwDueqkXjRZYiI3QwHr7MdTjupB65SR6IJ9
67hhcjoUdCsEUHZWPiXQzBHIaVRJf7Q4RVMZRDWCFdfydKbEJT8ToHtq76CkjE2pbPLC5tEc+hvJ
2+b2YOE6s+wuYfR47AX4u2ojXhlQdf7aAe/RM74M0k1QbEmfu7muF5vEUq8CE7zBNgIafSBBjaqw
fnGS4HnfvzqvzTYZEKdapbI6QWKaC7iwh1q2xT/v/Rc8QIja37F84cvFRs/fvBEoleCmWxyia0f+
YrIt/Vl0GwR+IC3uy2FaKvzHWIRHzJFhACBYxchBHma5/2ZMoXBkVutmKMXLwIS2MDcbLeywL88l
Xkmc4uwUBqnKUGKXLEWCd4rYOT6GVElTUo3J3Gv4/hinj6ALMUSh31Rv9EwDK00z1dSfFB1gVdfG
0p+2NuYFvpFCWMVK7BLjLmZrqjXgUBGsXnKHbEwqhN8BgRZGIUBulXyNjhYjls1HZPXXVDnPSn4o
69z4RhXVY67s6UySvwHUt1EpF9x7Ss98It1DrGpRYwnTUbvZ/UfRX0f2ZV5n9GvddhcWhKy6AHdm
TUzBXk1+FfNCFmJfa49fwc/Fcjr6lLwDJL72jKTopg4jMcD2kwenMx9slRl1wiFd+FvoOd9R4uS1
77E9l3lIxczpELe/l9RvN//yOiba5Bzw3ErDsDsc3qNb1NvkrF30vhZH8xYTWGuLMI2/40kNdSEw
+iZNVLGpOUfy9YdcnVLnpDmr0ysfHBMQ1zzqcjicSugPB9INFIVwtHunzsW2ExkJBFr/cpCHNqlY
HvOaIMR9Zy6swuCc4I5soEjTWBjnGJiIvkR0Gp5gpZ1i7uslIsZ1wLEs+5Rl0txfF2TSJxMGVh0k
Vph1pru2xTj+ECTnQDlz3thhqV5d3D4qn45Mq3A780pwUfoxc0TEU/6rIuJGYvIZcFm/HkXnQESe
7MYbpdBYiUhLaVxXNpIp7F1Eljv/qfS1FpXPu2AQtPyc9BD7ybHt7lAte2ONSw4g0yCh1d5iL/jK
HOtEoBctXbvfW9b8wwToXlJJBRfIRUTi9z7R/fuqCGy59KVEQVhFNw5pPVAQsNq3jw2qZkRkYNfL
3pSVAOcBz4gJxkr8ds1TdjeMawzI1gXduV6VPunK+Cy/cEhF2HwK5V/JfQXLmc7wvPDv4VaQ1cQJ
2n/5gRY4z/PBak2ZofaIyaHQLcfjzxSo2fxgWBQFnZJw46jEDmj/yo9Mcq8ZCWt0zJvNqHNTWQfE
bbGIa+Rd/kIiTrEPwntN0HO+2/tKkqZkIyeAsCTG+PWHhuCyaY7V/cjIv4vDtwIJazakdVMWeubg
ET+rSGS9ZpKjadBg+Wwp4pR90cerRNC7IaCf+f4//s8eYapuU2OosHogp9Y8iTZpWGRNxGRqu8Ie
HuWGJAJoaIjbe7eEwYNEr8kfTqxZIHeqEc0XukhP2FZt25JbRfRx2Oa2Cy2/mlYNQfGu1qRGxM4y
d0aJJg9OpENxL6EOVenOuQhYtABzfe6FytiDHmD2KBlt1TYZgZ+q40cVocrQXUC+hd1mRX+bc4aG
3GpllCYo9WZsSor8AQfTtUT6/A43xrXMnqzgy+69bYB6OUiEyFd8lT0b/yCE/r1EMJ/y4w4EcSkf
AERp5uLOGQ3GxnObxtqCzL8XeY+/AoYk7zA3VT/A39FspvmGArBT/0qlV4kQaXbWkaaRyJ5vVcgC
Dd0gV843R7SB09TiwQNsDMKiY3z+4qPyiCsMDxQ92EAX0oNNObRWw0qZpVyyHsohWQH9zvhjdc0r
8NLFVZ+/7iZ2nTu8/OUaL/LqkL7Y/VPS9Ot2ieluHH93W7jwAnyjjngU7f8vc6st6T44VW2bFJmI
LkU64bWS4sAlPzhbJ+GSQx2IJGWvsXAzgpBFXkAaa4aVfTzJ7P1Isf7HVr0phAsyAaASgsFnWCri
RWSHtODM9eqYwuClpuETwRDaooSDiO8gWKNu/GqBFPS2mNYGNGsRiA/gFpFmRTEJEOyPlhRbwcwb
WuHrchEqod/qfCcANmdqGrr19J7pT1zXTfPy0STUKJ2lLjqg5XTQq/y9Py3rCv4OYhRwUxcT/LIt
q0sWVfOVx0k2Pq3vxRSKxuEZ3O5HyvytIuk4cATQOgwfcVv5NsRMqA1N5t0CkP2sIvAI/zfmpNKT
g9QXUd9b98NoAEiK46jTh2U0SwxwV02Kjri6KMwKih6vONhEI1XDXL1ktYc27ZKlfF5YmRNZcRSo
kY17KuT5LWALir5gWUsQFvpbPIn8Npd2h/XmCaxB2BhXrYFQV/iSIWwWQYaBxPirtcSdIFTCy3xs
P2W1rYmzNUiVRCKSt8RpEsEcX9RFxVamxmf9ErOS4KUP0JxWqPxnVSR1U1vCI+TI38d9DNfpYec/
MJIfHY0tBX5NuXBw4q9PcZqfk+9e2Z/qNbfVpE2F/rWjy2zhxV/4Me/ScSXD/V6SB8TjpPcbu6Hz
D8gjS4bgKLPxufjtsZJSzd14dWC7y3Wbr14F46Onx7coS/32If3v6IrWkN2zxy8YSBRBPhuGEap1
uDQcIzY7gMlFMUASq2jMnm66SV7DoqUTOoBhq694LZCDJh5IDFR6YDhBZV6rzbSf8gzJT3EHhGu2
lGflVGiWI4e6LebaX7NUxpUXw4VeiFFkRuVXGeHPlLozhMAOjGAvngbLaFAfEdGSLyuYm6DsZL9M
0VJYls8MRRCDYtDjA7NAfXKgBoaYJ9oqeUK+IKfDNYGyaq0IlAiLc5dU/4GI1jvfr3mW+5nEE+jw
/toG2+opx/c44pgkDMQgYfOL8xqJMu4hhfXwNnQ6u0g66svtpNpD2NK/i+Dmf3nwvQaXysnTkR6B
I/LxOkD/Xsh0nBvSYw7iBKlFI4Z1aHiETXUo4GJfqcqpmcoW++owBrnkfBYXv2v2Jf2YtBaEcNAY
X9g7GalEcay0sfyNXi8IjnjjfXMueRv+CuXEfS3rvbHS1zsM3MfogwC1D//0nWqz2LQ3DnGZowmd
llwFJIoyjhyRSm0N3hQoiBzVND7yQd2OAxGXxLd+3XZVOQ6cDOikiLiw8GUPhlFlAFTUwA/QmBGB
DyYZv/pquP82bQinb/89wXxNYvqkRM0cFaivh0jJBISW3BwCgDcr3Y/JKoMwpjapwgUlyXSkUFNd
INtbLes9MBDNwvvdne2tbI8O2vvduedRq+qV2zczPmys5MTnGA9PdMHC67EoH5BpbIf8mJNb8VdP
bxxnRj/5w9HU1bZnpKdvQxoaRsyzZqvnv+0WjLxVG0Mv0lOtfqVgaNdkBqVwmXYLySdadl+zfv8U
/J91SePTBhdb1v6YpfUzf2Yy5PTsSXdpw0saR7LKgJp5zLanU++ts3wMQMwQZeVJWBlm4wvo43ec
l5COecjP9fJzlFXIqM19CTb07RAppLYPOkp14k21UWyp3q0idGerAL/zuxGBlun5Qt5wxEouDAnK
3dQPtYuvGfgbD4tbyZrjKE+I1UznwD1cD8xETumddua+a8SnEIjBMg4ovEOwUSpr2m6u152ZD7qL
V38WSn9U2AfHyuq0+hk/bI9U5Vy+PZCwR1Uj+o6X4tmnacJ+efPPYrH1NBEVjscGQ0HwJB54swf+
Nd+v/b1/DvqqN3GXNIf8JKc3277CVZJml5JvydlKt8XD3ptH5tSOObacIaWev2hzDeFstJvAsshi
GvbTbRGxBUBeUZW9g2VcKF5/pfNJ3ejKPUGUott+YVFzVh+4+8oo0zuErMmddlrr4QVA1xNpVQ6Q
yOkkhAaXZDaTWxqt+uudWpPACkbNcTlIqiV90NxkqRl1MHBwottc88t3cms6vNsMPRCHXqbNiEpD
KWYzM98qWfm4PA5tlBZn7pMCYfx94mUksQCLy7Wa6bq6vzOnHHZdYzvi/TYyBHdD4wnfBZuVCOJJ
5/VyqzTYSvfo9uuh5zKMyAbes9ui9P/68IpKeFrHcr8MMdhhgiVhMtJT0Bz54uN4ApjRC3P3DRGD
usxWLxX/HPZIAKTrCe2JBMZHpHpJyF9RawWiGDsCRrhtdweNx2VliPqvkBLma/YZXHdOwEy6QUWW
SHK48yPDBrwx/ftDnNUhmBaPN/r9gQFH8RVREDVqBsGbeWPlkYIVMTQc/aPvkxt102xTkcv8sBSA
tnC5fQVWm/dose01aYCJj1aTTQziEvkfsN3/aH0nsUAoyqzZje/Mh2RMM6LUkhO1Pf7KBOv3uGJB
SkcIW6nTb2hfJ/filnLdAu05RmV9qlZtiNS30iAF04Px2LsmGZw88ZBwI7tPoRfQEuZo/p6VR0Nx
8WUqjknyhPVjK9C9yyjDMV4a1Hik3hetWME4dt45WiPnjibGNwkzcPXGPfVhYI6hm2q7p15Q7vW+
IGOaUKlK02j/jKuhFIQoX29AQt60Z7+3kvDnS2R1nkRGn7mVuqFxSV1OxbJZmyW01RMGlRhrdg3b
BhqEGf94HDSonGuZLmGZ7uI3smDGMqIx5P37J+NzNsdIlECa5d5x5K/CoO74RXPdJvWwYO06sAqx
JyWgAM4CYDkdxCADgd12H+/EFfYe39JDEcpc33kWSJp1ikWOIaUkKONSmHe2Q6OXKM40Xx38QMtz
LS9z7QsZM+JUup3k5iPXPHsqLtvs8GRr0QluibOYVyf/QazGf2CN1KBtA4knYS0pXE1kyOKBaLms
v7Xeu0h4/UxvO7Qcift9RH/AGn9d6kNR2bn6hzcEwcCYo8YMnq0ZwZj6x6qeU22plAOemaBdzE7d
GxnGL8pjdrjwens4rIgpWZhvYe4kK66VZX0Q4WxRZPzH9tH0Z3glI4DEFs0zD8gFu0J9DVyF0rCd
TZfA0jecn5L4owfWw8nB9IZwV7c7G2Yg4EqKnCiPz5O6Ve58sjZIheOv3u7oqyMZa1HoFbGVrRVf
vLoQbUQIEaVnvZDYXo+SMQpY7uEKCHZjxbvY96OI/MEadw5xDp9RZukLUezuzxmGI7sZAQSFPwv8
1HSg9wJJ3VevPcFxfGhgvDRoRO8WhQacnatSBZ5CmRkxCrR+KnTiLMWISwwAf80/A36TXTTqSfzc
4tHj02ZJkbGTL/Dg3y3fZDa2JA+9IiSHoPELsIoOrRlpRzE5zE066Pf3Lt5tMkT6tX6fQRY6poLR
uyYBa9QEB9zIxs+5+L5ORiYKe58NZ2njAbUhwky7o6lAuxSUn6Z/4LkZ/lq6mInrPceMVfFXaVj6
rs97i6SUq4m4uDZE33JUUdTBvLvvjzRgztL41UVis9sBtUIR5qbA1ob7ClzkprGsU1GHNTjAnyk4
xNAEscA2w9BRa8k4ru0MjMGgnLW0oKI8/Mfy7b8u1edtd9nDZIvD64ikk2K+pgKa0tRBnrcTBrqo
k/gXBRbzubwDx/9qCd6xAHhPcf65CGs/qv43HkSx433RZoWo3kAOI9OsyXkvmlgTCzrMaNwwz9LN
I8h4PpHq7HExRylMPM3VIm24sTFxV4mbspnV1GKFEa+KMm9LL+uNNuY4W0tYrTpHPSWIVMh5n0zR
3rY7oyrNiRvhh3KD68OvGG3yHgAZj63E5E23fGVyU838Lry7rUlvJ+M7ORlOhv0A1A8ab2/KtNKR
yoMlA+ANZUzeX+9qyC7RPH/axH6mivLfsftWGNRWS/vS/oc5ghJy2Ri+Au5MwFLHaWp+UD7AyQSN
Lxaf/8FMH6yPHCL8BwHYeSq6z/YAGv85EON5qB0zdyPbgsSuB0Nhy4OCeSSSySk0JjaFlFbp/7H0
EQ20G+vj5dK5DUsXdXZBKBxirDFf4f4sns13A5MdSyKKoGGQL7Z/vG5V/6GaRn5+AhiueQu0iLGy
RxsIX6vIOFao0xBniYa8eOz0Onoyi9OT52ph5UYWyJEnWpXjpYHFhgha+UoHE+fscYrHwvVnrN5V
dCX5tfxcEuwoFichlaK96H2bEvWzH8EoaT46GZdM/H7Xg7TbmXLK7mZUcDSs1d4on5Viek949VZ7
JnnOUI4CzfEOZy3iOlS48KpP2aB134E8DHxAvQ5VX0cv3u6FcKr/gqgzJMGiEJuE3VPNlXbQICqs
lg0j3rndmxJ42DlZneRMa0ZEFBaNXau0rpyw4jDVaso0vkGRc2JSn1wKAq3rKW7oqzYle1QMyw3H
35ctHpWoOZf7rRs0L5eBOombGIZDrE54F3m9R2LdWOjENU8J6KLdR+ta3bUkzrOyKGn/MQVixvGH
2D0vkiAwnuRxaKAJEb/G6lvOQpSoAg00UznUiIxLMVL/+woybNmOBYqxC140m/jIUaJKQxyffxPW
ThaA/q4APorx3wQZqkjiVDXnuLNseKaZHMQ2pQsZhhrg7bZGULB3gTcAqm/Rf2Nh+VWWtppzDXWE
KtqNRkVzZEKQnRvCGnHCuH9eA0x8AtdJZF1ly80aICwu6z2rxuVU+5IKDM0+GaPK+d4JUufqv4/g
jYtL0BOplXpA8w1aI4nGfnmHA/6W5uJDH5JEGDD0PlYvw1pxq7Z4KYQeGj7Z1Ps4uJuMgAJ4mqIh
8xKSm1L26HK9g/Dw4qaoQ1HkVW6CPUcqEWTsqsIElHuo8bsvbbhlt+/cxfD0m6kc8jJzmxjG+qxd
IrarudPFzaN2HPWHv+/TkzdHxb0TQVeVPleLElFTpiujkMVezTmgc+XVqh6XAt616u9MIbdT3Y7S
ccbyLz+mE8JcmV+CCT2kqHvikMLriA2Bl0tQyc2FgKzBNEcBYN5ZsjwSaedkUapVQCYiDGaQ1Cph
3yR0faB3vzRvEdZqj9KjI8KIEgqWL5SFUqX08l8A8pwRiXIcLyPW3G1NcfQghvzfKJDTrO8U0BjY
GaPq84cWIy535vi0T6I9rVkoBClhRKtjTqKNbh+I5b81+s6/3eLfUMz1qbli/sKBFqYxVVtvNB5Z
jCnWHXMlrq1/dRYgZoUYr41RUTEte03xSDgzsIgyKZbp29Xyl9ukvTv8qQlXXIY2gqDeP0fmMr8r
E9SEnP14gUcET7SGIaBic7uGjABtAiA7tYSj+WZMZhz4O7ofk110wfFISbJEv2NhI9QgKzFjk7sH
0lzO+Mve4DW2gI4qAZlqiwwWuptvgtB5JU65YbGFFupNZJgYAaGMLWW8/jpgc1pEaMRbHKL/4Xfo
TNx6LH9xCHAV78JdUsq2BeL+rP5XMHNZdzTxiJvz0mQMrSKSRYE8a8bfHPKh/vPZzeMD9qLiMnBP
l2x+9muj/PJGLFrqgMfFYvj73SGCxWxCGnrbzdwYvjBN7BYVTWaEV9cZnfcj1/qZ7SYyS9LvrWTe
CWHx/M0nevoCQX/032Cf2CU34Xf81LQl7cnh1K6Z/6YIatwv7byjbcXaK+2Pmo9ohu3/jvkGO154
kS8ZHOXss06f1dTNAhMSBhDVluC6eVhBDVmrHUoyvUyscKkqlqwdc65c+a9F75Izu/DwxgPFBxZK
btwTrU+5y/FGL71lVORJWWzThNN9QbsI7RHwKXTwvJUubqciJqpEdmCCm3nJ5//sdTFpUZ835zJW
/jHjSG+9eqQ8QiZPEswEHx/7piG3dPheaSu0zvv6tVvIdMDBgEgJNlImBPQTz+Tx63IqbfpFu2fH
XB7o2oxpcjcsq+WOh1yp8j/uhS31EuDX3kIzMqDEfwTOEPOMAKpttodBZCW+zVsAJUX9VHFkaLB2
gJbypM/DJVeevJ6kVoS6IG0C21ED4YAOFIzEYVH5tCF2w+xHCL5DHHR+MWMuLIjjhfOmr/nokDbC
MqnJwMYtBEALPQ/hcCvFWTw58pAdwg0D2MpvmpbVT3VZRo8nGHxLxDLYima+rn5a+FA2qqVUyggK
pys2yfNZnFexORJ3TADicn/G5ThDeCdj5Tegco8FcCQQcWWqFjiMwWmD3IlHwlWd+eAKDEcKLLCL
QxLgj0GT94eeM7mLgM15pOT+0es1p1JemQS5NpSlA8FWI8AxyTLWco2Z5F35oAzDkQda/J5QvNH0
UrU2G5KBJ4Wz4SeN2TjeIF7KiTOIvJHyfv7TheZkjl/qn1QSa0LTnIFxi5udcNfQ/0mWs50T4tGT
Ux6x+J1+zKbn+Pp8aRY86ZzgXLH4GtfD/WR4w+h2gMgxaNQ75HhN9sMQCc1H9f0fvV8lscY7eMJh
CZh6QlSo+02Gqw6LzGaszH5KICkB/0K3r12JbBnJuzA74OS7niLf/8T691+Bj7ZRMI3vRfqYOIUx
J5VtXiqR4pmyI/I1DxxSKwAz2marJ+V0HmLmYs45+GtcOAMaaW+ti/C6FBHX3p+0KeJVKchxRxBr
2ci+xnn67x7q+rlMTetHZWr9bRbNAHrjSxRYJ0sWhWv8XedpUggmau3PUrnj5jbc5tHdqyLdkd5J
pPm6AtIdQlZ5mb711DzoVotuvOxJVW8cpp/ufIsmxVhZeHGGLUbU3Zu8oAqBh3u/dbxGDPcALw26
1OVxYnNDI+30Z2ig9AC4zffK+YIjnNahrm60jynG+XsefzxkdhD/nIF5Ax22l90MRR2iddelGn/U
pnt/i80YQ9IeSHokveW4rEg+8lvePI9rmAKTVvWfkAE4IQsQ4UrwGr3F8ZbUZexx60zbqLPVsiis
BfyekfcNvIL+rgR1CwzfFohNn+DsOY99WarKAtifFTr4gXdLk8ICJFySyR7utbBonylN59K1XbQf
s2jXxYzCbw+MN7TBEiClYxIugFmR0p5DvzPe5+1BOkDPXXrzmTn3d+UXT4S+BVZnI3tFhG1ZR57A
pV4zbMd+XrKVvTgaRrKrNTyRrS0mZOQN+emDj/GfxOpVbFFpH3T1UjCiLNcjq2McQibiHLQEPTRb
VjKg0G2d7pr6bwqYreMUUxdomXGZKTaZXIS9FdD33mpAwOguHvHNP9YFI7i8LyFtQfoEVs4C0pHP
EE9NQI6/TJPmTE99CTDRjBsOqzNaRe3tLbqBhn+Vdy/mhl9u6DoqnDZWuwRCLQ5+pJnmaCSLW1lF
mHTMRLmNXH+d0K73lznWi/S35RVCtdmLX2HP7RaLml/ayOmOMku4AdFJ6RDbzXkax0awLO/1pFgr
nAzdi4m1PQQB2rCucxufOROIR3SKOPLWlvt/85LnHW53U5Hm6A6Q2lookR/0G3E+BLwp4gTzj0Fr
DIku8acCoRms2jFLl8EykLrxAltulC2oFwEa8u9psbZXw1q6/28weCB5p+yc61OC2zZN4/rd81ee
Q5DRuPvK6Oo2mgO5GkfndDqF3/yDPcjI0AOQwcGI0ZzlCRJSOdpfH3T1YOihvwGfAuELUc0TJg50
vmsmwBftfyGd3eS1w4Pk02o5U8jW1YtWHEeZw27Lt2ZF0qzMYR4sUM/04ZzEdwK4nOUCV48Sqknj
DmKF1WKgXne5dw0cJa1GAw5KbKmtDZ/K992EaidKJ8QMr8XA/wLje9PE+DSk9/0BH2o/CWOAcyL2
JTyXg46m9acux8W5KDCFDopXdNRgNI13FcHARD1ucS4qV/iXfvqQFoi8g9jpQIvHbDSTNs7DN5ol
CBOgYaTOY4FiQgSjDC6938g4iCctQLA1HcFEZiLr3v1JyNF0CulWM+BbKUiZwaxsmr5g/3SnC2bE
bXOOwOZpYWgiNyAcsOulr0OmmmBhtYoyI9nIyl+WXP6gvM+5Ur2uOoJIHJ4h05TeF+qoiSNxW9gi
1POJz1MLdzOG+bzqmjRpIca/bFl1bmLZthUoo7hQJsBl/0EbCKdbt1c5NvSMxFlDA0AxZrNuz2hq
CCrMcZhGKBQJNn3B6Slv34rw+wTVXXFlIeOHq8vFbhxTxlDFxG+w6JBbpmBSefyOyJC51Uw1sEHS
OnZZq4pwxJ3EsoKJ9gk4vNdHXbFnlw0Y13yM0a9b8P2dCqTxY5WjUMtnzdKEKL9pT6OIpDtsLOPm
hGYN8Fo0f1zPie4WJOz8PSykHnj4V9fz0GHSzwOYUWR0xDYln0KsRoUAL1cewkYMAbiKJjLDNGDV
uxW4G3rTWmdyo9oVga0Bkqe1aP8wfrw/XYsJSccMUXTwqfv23TzM9jq358vPfixVkMPU0anSOyNR
6lx45rcJnoQknf6Ig5loljbLd8NJhVeS3zx0RThDiE7YrSLxoM2qhcAohdrOPMEAA3JOOobSlb7R
T9I07LvHBYFwMYr6Z526lfl7tsq3heyPhLmNwj5VVsOVHgWx8fd1PFrB04JYH078fQxutu3pUx6t
C9bbGHVFW4zATCfho22RvAekQ3z8TQFEDG2WpmeDv7Rollyjl5D7AmDWHNCkfUIey2d9iznT2pKE
OVknDko+zXlLmGHtIrY+HMTxdMCFOrsU2A6onUHeEVTE5SBLCFr3NcTgn3oHUYFubq7q3A8vjN8a
8tzZ3oNTLfFxPt8hmgRK7dur6po/g4T2Im93dllCuJecP9KWA47lyuTrB7jTTmVo++PLybHJrGYq
2VuYUQBsb8U+EAnh8Gehsmta/86NDiSnYkept2DSnss8GJJwVJT3v5imwT2LwonIoqlF1aiTlGRt
QJF/PyXFR8Xfn9NKrzxyIiJf4LbBg3p+YH6UGzseknkoxfybLj5A6WyoKv32+f4/Extg0GC1g1yk
JvrtTwCvm2zB0s8886Xd27g9LDqocB8QzvcOQnriHnDZsWkJGQfWWGXejXVhj9xw8dKehscCMMl7
ithYAEg1fL9/VBGXUrHDwfC8zoC2CRQYZSvYgcwEFTsX0bQGg+RsKqARJEwcRrZaFip0r/kW2HNg
V8TNBx6akSrBGuBwA4AXER6qzEspBfGyZbiuTm1MIuooYIs9OMSls3FlczXy0q/xheXWlqW/82Sh
pu9FRqcBzhxHdF33SHRCFIWgs3VwrFjp7vIp6F6PSDIKUn0d44Pk0BXmaOWVZjWpFY6tO5455pe+
CWj+mObhyma58Fb8Ows+CtuTfVXoIVS4d/BWerqU5gFVQ/Dp1hWeYJX8KVvvaIO6UeBwyw8xuVCL
4jkgTpPhLjLumxWpYCoMhNMnjbv9Ch3gJ9D5pRUiznnZGGZDc+9zbrj8WPOly7Ymev7CiL1iF5rQ
9UlkAih6Qne1njJucJzukjTMpUtnaRozv+4S9ujr74LjsR/4IUqnx8YmRLGjukmQjJytC0Gc6mVU
LNmal74+fWZXlvqPazr6LA6HEQ2/nFBnq2pD43Duw6GFO7uLEfUVukMBWJ5NPr5E6tfDN4cR8yvz
ZniBLNiL6nUAjVYXNyVPiEw6v/OrnK9nRfi0psl7sK31PJ59WJvOwSs5WLEqgCq7G5HAsQzAHrQ6
ZvsCABNh9OO+whDw/Q+BzRyRtnXK+NAthWer3al2Y+8iy4diPyPzjQ+9M1T5O/7tMB/0MkmlmKtN
ZE8Y2puF74Fd2U5+mY4isTrpVA6tIDwd9DJDUNYHZMLl+exFASv/D1FYKogSLmyye8qZTWyFMDLN
CgTC1B/D4kcp4YI1Pya2Nw9DfV2mR2EAJBx+eDL4dboI5Cdj9cBUEshCCQpAD7gbooOEOBuPYZV1
5EDTiEyAIr4ThcO2xCXYHJKimiXJIsL6UkXf6Ere3DMp4+twclAV9+7lOySn4c0+b1kCM9WPbZjG
eii/1MakO2EhvMJtKGMe63eCadbnL3y7wLSGkdwIlJqVmj0ubplpH5jaWf1fBP9DKtImRixmVev+
21pXMb0kasUr5/duAKmCdI9w6e8afHjDNaUtaQAn8U/bOnwwmSsBPJnbft3bh6sCzW7mszwMORG4
N/Y2BiUatybZGeyZH68dqCFd1CFMDSIund1EzsFM/AXn86UGlyyD21g+JnV1IY39aaHE90grZX0G
5cs5RNi92PMtrxTM7h65qoYMA7dVp2f31nxIOC74nFUTNmjqKkOKg+Qf+lcCysUkkreJsm6PbCu/
Ocm8ioR5H1eW2B0gENkduhMrwDGNljmF9qwSafKebZUHYEJZZDHPypt2s2GHJAdW4642363vwRAs
l5Mv4zx9qfBLjpEh69X6dmmp0UkvlfLy0KxzC69Ml+z7CEfVI2z+onESSVqC4yzojYVtHblypffl
nPlpmAu4O6KdYNh+W8RhjgbAblF9y4Tafe3jDM8qywOb56U5uJhhNqjHHh+iLeCGUMs9rFfcmxyX
m556BcKVenhQUvOgxnWWRNcM9vtEi1YJxGF15wvHj83wdKZ+ilOhjdHly6QutOVdatB+qY4bSnY5
uJAiuAdK5fui09mpq2FH2vgLqBHP5+rPRDsnBkSf3cCDhXuPOGz9VcreZyhz9FN/zBp/wu8xZVy0
2K8ZEiw5cCp2btNsGD3M5rb4DwEXucOMqa9zLHwC9bbjIGTrxyOELqQgRkCdOkfqeaz9JfI+AFUg
zZLrS4T5hACpOplrra4StHRAlKZNn9JD+3xDIGRa3/CVH6M2jfvwefbuH4VUL7r6qYzBS2/CwAgx
iMBAxg+L+1zNAePFilBUd2udBGL+QVaMwziq1yWLv3/NPMyocOzTcmc9toT4VfNPto2t2dJxN/cK
JgNjdH4Er+fUF2Caad/jvaSqMkDH9Dmdx3E95bOqWiTLps02usky/QnZyIO8mr5VIvEapbEElAgu
vqneqmHPmQXiTn5Hq7JQuKoxY1l6dJuF25NxRrgF6ybQEzBti8wEGjO7SLNkinE4EMxbrmIGV5zd
8p6th3d8+MAyst+H9n6/GRFqIRZxZ/NR2mi1JobIkNkjHvDRFZJnpelZWG8kQIFofYj5bUHRaUls
nxfLfKefLekYJFrQvUFOOHhyA/kFi55pNXe7PHTT1ZFrnNJpdYUq+OL2tSvsRBqs9s1q4GPzmTgE
QGMHC0hFwtXKZId51HBK+93XWMcwvXVegOv2LggUsNbEvLnuvlQl1U2yNXa/Ve8E0EA1zKxDQ8Sn
5/t1xWIt69HyF5Cxwer0J/iXSWYZPZ7hSb1Ab3bSqkWxpRxdUhfKfvI1095YuZVLIU3/2OzcynKS
lC93kKSRrrjNE8Y4x2bnJjMc+40xB0EytV2l8+k/JS+SwKamEnGDTSXwbRB/D3T0ZOf5B5HD1alA
VYAWfTY02OB8/yziWLRsD7J6T6lkU55/LsrgbxNiQjJlZtogyVHy/1VCw4fnAZfVlgFTfXUx18R5
TZg55Ql/YY1/+6lg3hNbZvhWKFLHduI3oO5KJIXr7ckv96GDrBogedK2Vxfpjj+anw/3A/LbMK1z
2EjIOPSWlQ/xNxwegfcphJ+dSLcNx0mrrcRcoHZZVytIpi0Ev2/2gv/P+v0CLB0Yak6F3WfUgCT3
h1TfkxJvm8Mka+5M0Y3qN/ynV5djoGPfe7TKw+rbnwo9a8U3WmDmpqZcBGB0qrtvGDT8fA+nJOzg
iWthLl/xHyAOrUSA/zwOYaK1k5Jn7x+ywtH2TK5AWkBZNQH55epCTirRw/Vio1yR+CAFHWA7JuGz
aJtHN3okHAjkN6qzIKNHD57YfTgng8fV4J5Tm1Np6gQNWuoV6zHzfMW8prW+rtnEZ1tg30EbTI+S
U2kbyM+8m1thQZyDfLEF/H9tkWf/ttSU1dd+zq3fPewrguaNB4pg2+oQIN5ogaaOE5wZpHQVIRXS
ymXWP+O64BFP1jBm9qaiBvqohCFKPdGm4VBglf8TfG7U+GENC6w7GfSzey3eHPXGl9QaKHH0U5hV
zfIHxU1Jw50+IG2/AZIYDaH3eV115LbebGnMtFWRKKsUIbweoLoy41bt9AhayVBI74dMtnu15e/E
f/997feWZ5TrEtesTC9N/uxSNsAGKKEHDwCLDxZFMsjek2bLNkaASYaPpEjKIL8NgResTm2dmyH3
2D4H1DkebiiBZubIO5rT8ktfCn25b9FlPbp+oOzFst6+7ip9vj/GDBqaHDL3jxVzxYXzLFU3OcQO
/ax7+HGBovlQxaU2DoKxbwjALOVZmlHiV8m+RA1Uy42hFspF0fhoBPcrkY/qU33zyjppGMtKepLf
SG4zYS0nICqvsorRK4w6cZ8DvDYiQy8auXnSzKUzLRMeIE10BDLqq77klxhAZxu6vo3z/2rYUTv9
J1rGoPq6tPHUSwwSzknEXEwA66UF0zBgVfvyBKFmIpOsuGSq0xbS58FIlEuyIQcc3HuS1ocGRngR
EH6R+Xj0bdPAZgslQMyWGxW/mGrtFj4+KUkHrWXn7GoPqgL6YOGwZOSJ6VS5ktaibBs5LZ1XS42w
a3+bYUHrkfsDOYrhgTBYri4gk4BXhS7ZmX8xMIMEsH+GIZVKkxYV/SOaW1ALcJOwi94FE9134Zb8
nYJfk+GNAEtCJ27Irock67zqC+f/0WMePDVl7FiaTFxh8Za1kUllGL6zII0Tk+1n4EuyRUTx6uQ/
syiq8w0Eiy4I5Ktw35Vorq7q47egy5W6Js1PKLa2jQFRTOWbQ/cqajGMJLyfB9/SfLLnEbdpdUtU
HbrbxDhNhVyTnDQjTP2F2RMks5et04SXeUy32bTb1Dp3oyvcDP52/psl0NnbA71W1wC885D+bjEC
IoVeLYT5jW5eNMHlm8o9ZdXbeu5JGk15/LGTQ8/ZXfT72/hOmXIj8jC9L2PDqt/ejuk4lL/zQ/Ph
4mQ4+xTbp0TIwkMIQtZrD2CQOl9gN2ECzCxkq169q95xWvuTi/nTMPNz+GfL6Muwug02eNkfwl/c
tluoOTZaWfHGnVL/Xks1s153YE1LSBzgL4NZMyS/O+0xGRuA4899CpdU67Pu8Xq+WRyuVjnmf4za
RlB41CkwH7P3Xp8AusM5y1vtzP9sb4+5+Y+c6tSiIjvbURYAHN3NSY0x5A0Let8Mhfc7+eTmVMSZ
pyzzZ7JuwRHGxweVY1YAepldNvz32G7KBpxGgiHbDD328DMDG0GUXI8YAgkDN/FitGB0yBFz0Ijg
0ECt9ZewvKM0cTRhZ6C6g5bcGcYC4xWSCXAAo2xCSc5U0dNF/fwP4RetABt/Gw5QiIEG5YFuhEbS
jSDWua9QZdu4imgVRrumW98Z+wO+kpweAbW75J4qQh2wfw0j+FEnDCceox1uNmDIFoEFhKLso376
093q2IuMR4BWnK6Gad0RTwscxUBh3nyl1AL4J+guy5rfHXiTNab9RC7FjrLZzCPC9O6Vssq7H1jg
lAs5xZTt3I0KNYPQnOq8dR7BdBjVslUZWWlhTkRQ9cVSzKlbXwH0dJ0aMU/Vl0J1M1XeiD82BTOY
gi3+TjyrW2Ov49Xfc/66EaCSbdd97M3n6GB2olJgVX9+5vzxfbjA9qKAJzjghV9qoVPAqponMxzo
OfADLf1CQypcjKM8zFJHPyECBGcqt0JvQGNnWJ0frtmMVOllDR1WWp6ERexYh+cxFq/dcYV3zkq+
v0cwlb/S2bV429J1lW+q9ksPERYncAOBDGlk/LpG42yymtbIrKm57fEpdmklYvZyurVoIUA0FVRW
g3hgYFO4P0X+MuNpL0Hww4qpztBdhVcJUvhtU6DXnyAuMtJh0VL2TMD1olKUTxEoDP4ewCF3fFLi
EkJCBaIyWbFCqirxq/B37qh5yZVOy/67LkSX4Htc1MwLjbdnh/SvLUQGok1g8DM+lUSCpjhfa2Yq
ItSNZqLkZgThPic6PPvXh24pG1rHjZzye3qCIRLSLXA1tVX/wALIwBFa5BlV/OFwbNGsxNR5MuVR
8e2jc1gkN1QGnM0GoGOxnpRvFvO4DpTUJega9HZJBUq2k+lrTQK+qSIajFVbWXw3nktEgyuGB81r
SEUZLF3HIrwj5TiiTS41N6OyNrJscmvE/u7rQoYFpWijo3A2xg0dEte80UzSGlEZyu4nVnELhm5C
Bgz2Om7p1UFH6JdgNt/H73W+zF9QRx3Oj3sBPNofQQiN0t5ALIID+LfXh0GvoE/zcEMCa1CyqtNm
Hx+nLJvntO9e/JkAjmJD/LTD/Zx8Z8fXf/XZ8eBTP0SpqhR3SchTqbfHlfVHsB3Lqie+GFF8PZQt
hgNe20w/7eW/Eb4FNEAm+PBUPQLnvUkGImuBMFrck9TI9pDEbCOIDnDHV+d/lyDZKf4N+UIcaRgS
/hDTHSj6zduGZCnznxKtewJSenrEqGwV989ey2W7VMI3sDQ00CN/edQgjU0/atthxFmGAsgXZDmF
ltLqftXkDMcr2fuN5gdWzJp9aF8VOIWw0D6655D16KjkBsjtl/zdCjPczfaME3KdaRUuNNWn7+O2
HtbDYeDSaYCpm/FpQhyPapLB+Hz1I4d7jUi1P6MHrSIw02alhcQjoA5hme1n3GZstdAl9AhG+CoM
cRGxoJ6UENTyh3gmlU8wlt+xKs1nN6PPye7ypfegcU2c2bEW4BipU4Yoo5yXQyW70E/vzAUF/0Oj
W/O8YmHcaGnY47ljMxnouF7C2coLKJ+X+q/difOfG8sA2vO6gYVy5fw2PFipAn6lhS9fnAzrL9Rr
CedGKLGsRCwyXECdIIXk553JI81lcoPPNXF4aOVnNfNG1e/dftqZn9HwX9+3K7PnZ10GwIV7h2ud
3wGW7Jc+y+JCFacPKxLk8ipZlnxH0olM2MQraOgA5R92tH4uFhoOo21TnsabXTVzcnUbIxs0ycO6
Y7qtnsqdXM9sOTtN0jA/lNr0f5cnEg5A53ivnl1rjYKo0NmJqi+By6ZPWDEW2gjjP/qgTn7K+KRi
P9eZuOVUmQLPAcTKKA0Hhn58m8gvWbCBniCnNog5wq2SWKN3SIDKchsm7bOc7Ysv0HO6C2NFxVJg
z03FdLhNJQFXKvGZTsJkaWTUEyFeU/MzKbV6I8eG+/WjzBpU1U6bXiwSoTeI0uDTGX8rlyc2hvCh
+4nvfcC0kGCBV4cjjqzBjsAe853lik11Ld8q5CHb8lFPCDjlXC3bqVsI84hEMb9HS/jXk2PutRpx
mx2+p9CiqCN6DAF0t7OoP25vq/oScozRWfMMIh01zVoa0PHpVme0nloTazfbRSaSKu2RGjycdrwc
Y5MBXpIhnNePeA+GMhxE0E7h+eqbBjMQ6SlcMwL+ttsczJIP7VF+9CtOItt6gnNQ0oP923aopLH6
1qG4cUPV/xZEmQTbJT8KAN3JqijLnAoLhGMo5Enf6sSbUhxW/rYIuTkZf7pJuiGDMPE3mmeD1fVa
/W9yDpC9Nd5JqlXw2Lnmskv8zf/itk5TQ93GH7m91yMx+2Zsz/u/94gAi+c2A22yecCHzWZrxTnl
MYsaxMApcbovVgk+UftcxrjHSzWqOnx446rvgnEDIqKxU5pxFGAi9ckXGRjtTLybFlNUkPV0mLSb
aAl4QjxnGO7GgPpR+y3YkuiDoyZ3d6GbOdlzU8IQEm4Jos/v/aqqTV+TMPIqxyBsaGmCelScOj78
zZX0JgHYBxkjloBZaN6Awoigjn4Vkg8oasQw9nYGWkzNAndZBhy8NBlvhwcxqN8v1HGPUVi7xmkk
LRIvYXJktQPwPeZ6gmDKSM/WrTiX0YxzmIOeTyeD9M/U4jscWUI6XmQz3yFVQZjAAAYigvzYWJTy
H39ABvvuo8s9H2wVGct0nPUf3eZZGYP+flGfeMH9YpDUkEAoy4oo7BjtHcoB1CEfdX0qwi3c1ec4
t8iwbgc/6kRg2paZb8XDD41O1TiLCMYwVT1ZaJ+sIqcDHb2uMk1BfR3+bvZqs0jjQPhTyEpxG/4f
UTgfPwrvsecapWeEHM/fLD5K0aTe8Ro9lSUT8NTdSAolCBiq7+fOEzwmBrKm1TAw2xUK55EqeuxG
+6Fqp2txyU2Du/MlpXxHdArQb0H3bugRUo6UdyiD3IK/si8bSLJuuomx/wAqDNf8xHjepMMiuaPv
Ew18eST2+ZptmZk4c5i4k+I323kKFu050WZ9pz8deBrzPRnQwjPTQPCl0qC1whCGpfg7lvBq179w
p0moAYPz90qwiNJpMXMrVpueEJdevkNuJk0KX+szp9t0cZAaOh1jTCJOwPbGqvETsnhHlZURuAV1
v6xLhHu2YwL2Z3yTloNDDsAACGzDQmQ4Q1FB+wbi95hRmGO0q5wqSU/dgl49hZB3vmCCVeu0/h8i
vbJdny9EuYQFpvBhXv+8+0VzeGQUAyAsGfF5igbKXFePUw/lEoguPFtKLdWhTQnh3HSw0i4e4Lj7
eeZTJJQ6TbqlQA8tKEVWrJhSyEZ9nn6qZeuAaWphMUsnOi0o/5v5F4KONZK9leYbINHtpwXQYzmS
RW67exOVDh+ym2EKjqzartH6AI1efPvTCFl+/atsQIw6Cp1l2/fclCYjmHzxb7NpXgzFMlHb5HJu
p67yMHYud4D0XTChgUelZttTWOejUB5C9fyBKPpNvoNOjH2j7JHPgfFsXZD7oj3bMiCuynsviSqq
VHBTXjpc2Hpor44q3bBl6J4KIzAbdskXccp5EXNQ/U7qjB7q3SY2HQvLt6050Y5ETxSuU9REelEj
8UUEXrhA7Wy8lOxQU6A4d2OLt+ATq2zal/1z/VnQ26jzLcgd0BnAmEJR7N6AAGMKVYNlFLy8F6ZQ
t+eBJrrnS7YhZ+V2uq0IItrsqAyt675qhWiEL2GN97YZALrI6NVivqDf6ysVCSAkat+7TNQ6XbhM
2CQ3jKQT9nw0yQX0fY1g2EQtP6GAUulJsR9xXQYDpsMLkymgtUSwyUIQPedh2PQTgsi5hILUGQS3
MhZbEbP71KxqHU9hRTGiooXrTIWcPCR9oQWO0TbyY/UFN78AMN9rioJwTsoPjfn672hoxVw5Gsrl
gX1pocAzCdetNhvRsE3krjmO3PWq07DUUVxN/pImEUBbhjZjwV1oGoHetz9C2Vb4Nn424p5n7ybe
84JToO4pv8y0i2SyX4kxxg2AF3dMl4PASUfbbOOdiFlf5sXr5f+jIVnwqqJfdjvZGvNtTi8L/8sJ
bUnz/UJWFoV2R5kr0B1GAw8+SJj4nYkYRx4v5iy9HT729w83a1S4KNyEiuvOsUOeyD7SOsonpKX7
HNdpKMjdbnCKle+LK2i5NkVmZtHY8GehxGDkPDlCj6ag4uetwrUzmwNVXhTQbtd91RTVtA2OmmMz
cy4p6T/ew3+VSMYXHY6x7V8tT2jxwgw/8KP4stmZCnDnT1oh/QJS6+34+v7WWtyf70JSxF9A24O3
tPx5RtYTJG11olGGPLZvZgoRm7UELy6dFzjkyboKpI5i1J6G4/y1qXGjfZnmBf/vU4Xs5f1TFBU7
EupDcpSHRXT0DI09oz7VoUvI5KjifOtiRYSpO2AnYX0RKbDi/RO8ncO+OdrbCtcD8p2hcsjtBO0C
3KnSC1UA/9mb2Mo9sjhUDkaVxU9ymPxd+eEnEksg35iLn2lbDZMEiwfReCxvPm2MerSyl+8lBVXw
AXofIIsBAAzcVpI3QYIGliP4te1NW1gl9zR1vZmmvqD4rHiIHR89VUNebi+4iwzXh0UfG6WjaI0t
ACjDAFhvz1fv81UKfUVIFRfmL7QXMvSsDAmB3e8ygBTJx4mZEzkseJBxhjYqLMj9S8iDj9o2vAhf
1TywlzBtybqhpJZUz5FatvfAK2vWuaQU+L5V7ZU4EoARGHuMTNO1exm/uOgiKwfxvoFlOLxc/jjV
O08xIetIeJd0IJfAA6Rin/9YqX5AsihJ0yIflDq/ZQqSAYqwr7T2GVtHUE9dXSGT8ZvqLHMbXN73
TniMmMvEuwEZ4V2AliS63kBX+aUvoVV/jmmYrys226/N23Ak912pgbTTj1MfJWHJblZDBuzmyYyi
MkX0etEm8qB5AoQDr4XJg2zlZ3oDJDg8zZPXRXOVFtUlT1Us1EFtVq5sZrlQzXGty7E51tplHZmr
HS/qoB50taaTQ6r+LXcPj3ZjvrDlKaXMEqMxBta6mwHG+o4Y18eHh/iyW5zhtsRM17HRtUbA+dTD
lwTv+LLmAoFNByxSO/lsmmO8hL2gyU2WuCBBDH4l/NkiROWxOBzXPNaAb1GdHQX/5YAeXA8sGOnp
GbpxpE8Fwah/fUsAuGJR8v7PZkKweQD+9+f0Jes1zuW9QZ4BjV59CN/Q/OEqK6Z2MaOpo4QK96Jw
bSkYcxs3X0L/hcSpHKpas7v6SuGLNOqde8VwI6m2nhzAdmnW5PqKYTeVYRvhM36Yvuo5H9IPgDdH
QHSKmOhk888AZNYdE/9sP47d8tZhFIGdCKOhUA2Scf46xALhKsRf5E617y1n7W3wp61zvdfgwBol
jlABy331MEfpbvEPyu2kggmfTsjULR2LI3xLIwt+a5Ea7c8x4MROLBwYRPYp61+QJQQyqNOCF90R
n9Qstqf87tNTdbziTw9S+x/Fahp+PqAgWbulTIcaHlT+6n8ihhAqi7dyKM3clSnoOGP27y51ClAX
A9JpMdEzKhS/65XTBW1P8KZ6Ko3JHuaBuqd+t5OQ1/VZfpNxKH/tDITtExN1C/5FcP4Iw0SZ3gu6
AnNFEsyGMelJNWlSL/MZ4ikcDG+ry5atnMg4vFGrry80d6LH06Olp1DTx64ia2s4PZLuly00djeR
Bmu5NQDrCZr1sXB4m17KwTWPfCP42Sr0H3H6PosJklx/hTMs+pnajXSODIUKSMrwBW4zP1yPnclt
oqzYXk+Hd80V1bp6k9M2yxnjbIHQFWqnnZaBCdZ/1hDWEhtIeWqZQNxH+8zRxaL6yWxhEv8RMn0d
2Ijusv8svSxNPo/7GMs5LeiYE570mrefPP08k7YCttKKkFjrxY784Y+KAYSUuXBJAzOWhNVhviPT
Bu8Mjp/bIWI1kFw0Hca2UodgEmnEMalTrQWsdmmrhMMM0gPhZJk1F43/RxJXJHZNdyaluOjNkoeZ
YcrWjiVQEF1kIWQkZVUVLvqLeS1pbAZtDtBG8PI3hCN4iaKppSdHoLSfWUPX2pqkYgqLcoCzaz+8
XtuBN1Iii44CCg/KmLaVXbBzMamN7pOzMOlO5BBqOK6pUd3gyJCtRCm/laekuRnZwmvY1gJDBMzB
AQ0E0fZSxEdDgAuGDiDjH2cR6bqZUjcmO9r1r4QQk3SjMTIab3gA0byfdd+gg3/wK87N/Iq7eDIe
qXc6SF8ALLL0thmjRBqR2jb9avJSHgBTjENveQtV5DlgDOlzXnvotBRAQTRXQmh6wX41kfNJIlYg
ar05HfvLEJwXzk3NqOg/S5IoMhZi3gGWmFFztXOMLyiXpWE2mPrGeYHfLChLgPt5g7rS07aqMmwg
PE5PdXTAyiF2VfVRHJ4wFLLjKsYgpAjy3rZ09kZGmDNGh4JAceeQ2yT53I3UQsyomy0ythlzKyvO
bESkmG6HNujV7KCEpNT+VuSktTrXkBGUGV8kg5/Sj6pyae/fyKDjsh88yT/FgTdLAgsX4aQ/ASHZ
nWl8aUDWKQ7Yvbt06MCZHZ8JNTGqEdO0M6kqGVXoXxt7qu6rc3m3u1BQu7pEVdAgifPjlrt4IX5J
IcrnJ+RYcC0d47TF6VaAhjwvFZwJBbJ1s5d5zmP8KQpcOQX6gITC+HLTjd5oX6sjIJV3R7bzJMEk
PgznbSsOwMIi+tDy4co536TZI7CyTNZvXsopUJYI//n6u83azsycA8nn3I8wKCKwU914AKiAIFTn
PfrnkR8CgH3oRBTjzdNwSGFzmT82wKiVuSxPfRoxoyAKENaYYXho0IoZhGpGFUFASJ0cGiHGj6g8
Clq68Yz9eTNJ75DjiTjXXt58xQ88bfuGliroVWSj2cllv91QmwbCn8FEYztNcVhiBgY4JyEG1biT
jow5JhSyZOiPlbxbB16fRrho+Z3U8TqjqckxHcYk5gslOjRIodAidvWF8dZ+QO7CFerHuPqJ3ZM8
D5B/CkAJKz3YWgZD9IRJNrsJXQX6Q0Aobtz4gGeCPO4lP9VWVY7j49Qp26csQz0+B2exb6Q7RaP4
V2+d9DTwqc4qM4BCEiGW8pq7CTyr0bCXd5nZGQMQOOKaU3qCUYKF9iGtrZgpTzMu2jgcsGv9+1yI
OX+o0vOInr6Mc4VC5/lnThBzuoNs1SvzABQfCMbrLhdphW7jD7W8lUZ7oIMOJHSAVf4XMl9sSGUg
vULSyVEzSU1u4K8OIrbBth4jgmdUcArPjK3Ja/esrdaxk7elYau/etMRhsi2S20Mj4gOa3pYmk+q
1+8i+gSfdmWrNQJ65fjQwSE1OBrLbpyeJSxmQkqf9OeNzXrQbEz7gnhnPWKgaY5jU6v+6sijMFTy
Y89rTKqJZvzVHq5NiINXj80QeH9CSv2JbNPWeP2ZO6EPFi4dRxE5w1OZXfEhv/Vr8aRRV5YJ8GJV
fSVXq+KBeeKL+T6dk027mLxQM+wiKBZwQA1dgv53TDON6uOUMYW3qrj6cTZEX5Alp08TclnqIO6x
wFBKe1D7khVFc8q5cvVD2zjbAi1rlrIty4+eel5k0ahbHXxuzDbi6gv/JLbq/1M+fsZSMij4vOBa
AsqAgLrJXqYyceICz/H6QJszj4DcV0NrJyC2iftB/OYLwRJ8g0F+NKCrP9l+8aUw6qWOIbs52Kr4
nYLESJsnHNxwvCMUlwJNeqxHppvVNyITvLrSpQAb02M7Pou2aoX/tBJOcRx2pBW5QRoP+VsrXciN
h5dAA7PQjaM7sAlZLifx+GbhV37hsi5CCcR4HQyqLQB/FCrNuPBH3wZfueJBCqKzLzLSvtKruwXX
4F1lyFsR1meI4N6/iInCb50ZQSx0hyIQxeWodt/yn7Co3Oge4w1+0w8ZHaHFawttnTmYDzWapzpR
J3mL0iIS8m2MeZFCcl2RJgL+5rBAPm0yEAQyNXTZlTgqoEAJt+W/CzmRGDbPf6RojP0vyFKkzbea
H01PNRIXRM1WdUNskL3cuDGtZCCtQv+yIOWbUtkDqYbcU9sXKUEe+mEWTt3LNCAna02x7mxgFWC1
0s/h+MDCVVn/YAoWoz4F1/Z1wkwwa7SjM4qo323381Ke8DO9nZVU6VBea2+ovP57yqY14yfARjat
KkBMnqznGF6S2qbwd19nZM3dlyDxiniOsKaBKXSr/vG9XdR/ciJUIpfygP5xeaPtMrBx1sHOI1hg
om+aRlVbW6TJ0YAHNeYX8XkgSJyN+RZKS7ztjS/qqujBsZuRqdq8YGaqUe7KFQHduxjLkDf7YCiN
WOQdnuXGB2FEFLDp6UzuWBkFuMv4LUZIEZ3gO1VKvLqOf6BnOJJsKQpW870QNsxE6ekLmpKeZ1Aq
ID2PxAy2iPlXtpAivWqni1pgXRVx21JRrsBQxlFgI5lLZ0BJlgXKNn8IpcumvxHUBep/ear3ls9g
Se5GIG8nqUmrO8yAcudhxylSL4CFln/9mnZaew61gFJpY/Fw3RBDaTg9/ibEVRY8IFbXDu7EDEX5
TEkjVFmYDawnImAhLZZyF9eYkIWKN5XU8No8Ka/1if2AbilHo7hIKh2doM3lBt4YfIjqEQWJFXAr
oqhDs+CIqTzJc60+e3Mu9VVLVhfGzjMXcV9J7IdPhLiqnqeFttV08Db0r0Mje9Ce8viAfgN8BTjM
hODSy8Ip8LTuyXzYtnZarPI2zGekfJVJlf4AiDwH2AtMyKZJHrDShw2233QJSGLOy6qn9xncT3ly
+PvClquusdY189OfCn5rQ9revlEmUfX4w1Wgb0L+ZOmt0HsLmnXTJEX08IvbJkYlvQ81qOdrL0Lq
v2CqXTsgCZ9nfuCJqRlvaQqo0oBSemKuNM2IGigy3qrdk7unZ7bXEmehljH6wVIb5G7HrYgrAeId
ED2uG6VVqiSbY/MLyo8pcvk3PVfWooo/9zqCOKsueFULcQRKP+5PBJ3mG3NzDfOslB3+WCfuNzM3
cPKJys5rgSxyp1Aa+Gu+Jpx34ZNwZNh1vZwyCH6ZIYz5kIpdQoCGIyQ1PlxcrjWmR5E789dFq65L
d9KbzE4sqTxprd79Ga4fXRxFv2G+lMCaPAGuJ8ZFON+ufoszCASiv/2I3DgT37dj4wCT4PwK6F2M
NcreSx3Mu4+Xofb9EnipvKGsFfTdXxM6EvwwgVCMjosf3MB+SBJ3d1FqsFwsn/0IhAq/iSu5u1jE
eIMyeEEbu6c4QPQJJdHXczcao6dFCmXqvvvElpKDyRXoytss/wR+gn/HXV7BgZ9LqPk+EbOo8aFp
aSGOYnl2UzvvUbCPoK1Ci6n2twKuNJjaf+zeRE7chLgNWxdO53Syad78/Jm7COa+xgoHOWr1QwXf
7GS/5C3D2EVQOFLTsfLyip5KutUBMYjCBuXwsy1qnVyb2ulejIyFfDwPJMFSafO5M7QrgpqPpb8v
61OPsiOFp1O4XkCx5KD5KIGT0lHuB4fA85Y/y/U3/MrBxVSpniwhwDwm4f3YQutg+BjM7QTXW3vR
sl1lodjshsvmkEFdqRc/PuZ33Hp51gcW4OyzJBvnyU0Ow5R/hpZ+ugs+6dR87QYg+ePCoPKVafLp
thzTsm229tDlw4ZQI8sIbxEZZWSgOsKzUVUomGpYejFxv0MeQN6V7nST+CXyNSuwUb5brr4ll026
feNZFFGaVyY6GEpgCWUYOnwETQKgIqpE5Q1tGhXjynIElDhVoeXtbZuQ3Rj8WDYzO6NFRrP874EZ
u7FINqv3USHeNIs3uBlz3J4zsAmzwl8jSn5ERkdjr9kvk/YY8c7DbVQEYm7fNg6zYbyYC3HvSE6X
7/GqRL5YAhge5V0eTaGfPFrBFZb/J69+aZ2ae9ArJiOVKU4xnLHUS503Mt76f5IC5IIMt8x1R1hg
51AaHTe/b359MaiWZKx7UA1V7EDQQfD5iIdi0yPNWmUgadbf1bUhaiadag+MBE8oQqRzrC2WKKsS
j1vMPOi6h7+DaVTAS+NMK204y9B14asevuciX81Mf4oLNz2DJSPqonK9Di1mH6f1QxRA5KG3uPZs
evcTIARnp9zjZnhpZGPMEBr/IrxHDzqYj2NVusgApNHZett8uLQlv4oHErpb8Ghk/jpqaOdLnpL1
nR3Pg6vvQ5EiWk7bHXtANKTASdchAAyDxcggRjFMnbS9LNbmB0jLvqnlysI/omfqgIB1AjXHqdbi
BLhHFf0Fq4pnghjzftjaTDaOESS2ltSVeEl67ThSmaNEApW4L4PY8kkjzD1JVyyS1p+yBNkzBNGK
exSeAhtj8COMFxsvlC+Mco7xoP5RLvKgtbvAd9gZTwnyTuZZ/RxayedvH0952nwDp2KED16mgAru
A4e+PSt0wTwqGWDZ/NkJboEtl3qctbhc/W74LxqRWEWzY6s7T5ZnA2pxdZWRUDYS5hOuR+07yKLT
/pxZ4GTFVFNoBjaF0px4OT8j01KmXudhw/DMtTS7eAROmY+HBGNHWmzo6fPrMdkC/HrujiF43MJz
hnkx69gKu7V08IMSBtV5Q8+8n/tXGbJ8dVUIo4m+KkVTRxsexh3k63bEwjrdbjgf+9KZpATFEwW3
XyrSezmcrnMbjpWvifPSQCe/9qqC2zWws2dQkrhFjA9wPT1qxDEsrqTgba+vVw/O7tZqEH2HH+Q0
PL2G3TG1oFBaOvMcn4DAchv04vdIJioSgjYOi8HfW0Mmlp/6NT8PnivcUMml82Zeu06iF3B4Bf3D
IAciXEQza0xdNuTGxYnxClMujSdTAQqAcibc+WPco9EKyIjm1NLNdbX4p6mcl846o3CVoe+09Aqj
ao9WcZKk8ZyOV0wGrXT4y6OE8T7TblLPB5I8wCM9pfwBOIsTtlD58569FHcGmDI9BtxVratbmn6D
fXh7yrj5xYhVPbFXfo4burRooqrd32hlqxRDqWiijT3lhyOg0Vy0C3IAQfB8kXEvgmj4R2mWPbsJ
ujUl7lGtg5UUY2qjpZrQ02fztYGoG0j88E+MTd6Uf9ceOfGX+CeZGj8n94GQ7kUqHerRxvr0l/qb
JSyaFzsN4ioHYUO98AUKRYGkLLgkkSrGL8oczdxDFlKg2BkfMUcBUG0yM92RqvsCKibghDa51F/O
b48GxQ7uNsP1ywVs509/ZJL6tC8elSslBtdacyD+ALtA+uZecyiCSNex/UWt0Gjsv7PHXRyysg4Q
C54yPLdPtAgWZZrv2baKZ59m6GY7Gp1g65kI7C+eroCK5WbgXVtihz0FkHuxEUAfs5q4G9ltB9fK
1d6C6KDC4ClclhIns/+5N9aWlWu4OGrlbpkclPlEfJNYjRL29iGY3clQQYc285WplsHvjUAl8sFr
aor6N/TWX8oSZcfaiApJarGklcpzEtCoa2CChEMEPLrBFXvjG5PPW5YRLM2nqfzLY1hz5T4WXHA6
uNCS+7B667meziQOHhCms7p4OgihRZe4rReVZzHJ5ZTPuQSgasfBnsvzNEMz/zTwq5sqQgmzCtNw
7qHYly7wuhspQoTQTQfLrCF0SUqljyxjDUK5hgtIC+6qgk9F/PD52b4DXF8FkzdUQOV/g3u77qJi
L/dLPAiFsXYKy1jAk3x8n/aah0ttoHDn8VDeb7HBGyfwEBbB2zNanoBWewNpfeb4J4lsS90bqsDW
+BomWOXyutGuCF76jNzIrqg8yl+XmuaJ7a6kKqeco7mZ5J8l+9qNEW+sqbaIIpDFZi2B0ZIVZutd
KcKzJcBCN3vPUcCfuaFqnAK414NY6E73vTEu6+jtfuKrvmFgG2MfXpIjOQhMPOP6pMAWVs7xVRLn
JgbcQhytKvrU/XXhLlVjgX48+ULxM0st7ZHUu2JSOMvvrtiktPVa4r1SF3Rf5sEz4mijuHVyVM6Y
x+wJIUhm19bMREDohPaPzvNp1hijW6QMMomtvCfcTto3tONsGSLG0JBFY/u3i6fDSlz9U9nkVwO0
dsGO7LdhkLDLzKyQLWToecIwoWHZCUsdqsquMRwCiUWvVuHWGZ1vLajXqUHXIB7XpNswqsLsKH7V
zPld+deyGORiBHpx0STKl2H4pmx70DZhGeH5P+8pv/i+AJ76v+DUN7kyRJ/boi1wvV3fIhxq+WL2
ixg9RRPpeFM+wWfhnwsCM7eQN9Ev7orIWLlp07QfP0cC6bnWMrBX8b3MoZgB8JlonFIAn81G/OUD
26dK+KAGma1uEUzyYW3wmQH2f5mgLAcsd6SQzf3ryo56ivdsje3kVuHqfmyKZo/pCNU+uYi4BsOp
iLmEfjt9A1inv7d262vg2AY5w3Ni38UINP4nx6v5nnvNEqe2YSCNIn/2wec25xlpoYLKte2Z34th
T+MVunemPJatrzlZLpNrljhklyWFvrXaLlTD5KsrJ3NiE76sfVhQD9M3has4DRVCqN6iMAl6dKQZ
PzkaA0KLFkvpFYTwvgr/WTtfd42Miu2D0piT7O7Xexl9VJ1FkgimUBGCd58tY/OJF6JlVi2uSJUx
Cauwg/YrWtINIx8SD0oZzjBX2f4MIUHj5KOPE95J9STIhgJwgo/JeJRZvJZ1FNTBnosMKxVH7v5S
7r9Ri2KbpeKhvE9ODcmivxzPIwTJ0O+Y8L6Kh/uiOY+zos7kqD9uIqBq3brHdHvcY3UhoausXQzU
2FPBikVT/HJYr85STAu5qXszz+vZ4pfyKSWDS5V/+yDk4RahdDCqQdT1zfAKc9QDIp3vRLa7dstG
DpIKOqjGUkZ99g1EbHzDeqC4s2NU4cX8LvDCBBA4yatBXFiIutrfFVarfD50lhh5et82ymHRMptm
ltAorIWJJwTjO+DdG7iT7bDRcNLkrMQ0rrcZEXKLIYas+X+Dg3YMmrTCFhJFiXenQNomVaGIjcXj
MfUhxM2f10uiT6WsHXIiXuCR8I/n50u7uvvoaRVd6ZHJ9ehlTSvq89KIEucE6bf8LsZ/Z9r88JrG
i8Q4UBwl3mXMaCkzRQERDu9Ol4M7XZRQAjOjPYjcanjQoJSgvNElhnY5RU8n59ITwahafMZ3cQ16
+/nnj/gLj7V885R7HJ0Xg55jUKmyy7HWb8gBRre4kp1R7QldkQ1w99tQZ3HrUAWlV6vgisoBBReg
1iskMkcQ3F7gZAUyRu2DBdFdO4JvoGoCeCTe7tjJL4UZXjI7sXhyI6UIjGDp61T8CMa1wRiT+4cV
gfUTgGEJdXV6L1QVd7iWvcU2oFvctQD9kHAI7SnONbu1Ay0RgCiOmdbvl0IXP/xxRJ4azZ3nrJck
1bDvCfEIwQW3FlB+Td6bjCrSMIoyiIwNoZ930nFMF5QhIw3yogOZsPs5ZTHfpQu6Tlpss/udiYQi
N5LlOEVS/BS1XWuGw9YA3D7Pkn7a7NSkGxLlOziSQyFQtas4uCxLZoCB3XE8Ph/3YeuqcI2SxNX/
ptuU8hde/nEx6XRbiOFxbtesnp6c0maHmkWum23Phw93yy1R2SSnRsNDSWs5Xh7f6/VeGsHpy/00
ReMvtE3pZc/cZ7KCszUxPzHP4M1tGsHzzPurYA/DbKpMO3myeHRREGPnl0v23pVr1newh1dOvFUI
LHzLVjCcqAOfCHqQXdsvFBrOhiIJvGx/QsOyHC5HgnRONYw7PURH8gksNLoHOBM7Acn7jXO2FI0k
Gp+Rw+WdWQAmXGdy7yAbgy3mxIS1Ck+MOxUX7Czdo5Z50Nvk4HHiwJ6efwpfw8F9mrGyuR8JCqtn
tePRMoKrGns5Vc3EKqHvMe5gGKdffEsECXcHwQ2nGi3KFdvSzU/bivFVd5lA8kQ/6xJyHSL+qS6M
sxhEzHV6vPeyvuNJwblDCYW2Ogh1Osu0bTGrMGUtl89rZKxzeUMjSTGuWNBWuc7oXAGOfU05ORYy
yN0HvGCZMAFvGltOdYdjyQ3b8pWFyRZsUqB6bX3dr2GJjR7z+WICwkA5ScHYNc/pCDaO3sCYksWb
xXUkPDJvdDgTFfnVaMGtYgvtoSRgX9Pjnvuqc0sJ/Yr2mNKVZ66g5n4b+IqIGcUXymsP7CU1Lc37
eGTb+GuznCsk6ZCvl+/gkmqhR6rk3BimzC34gGFt2hAREopULN+UudvBCQYU/FZ385gzZSOdJmry
pPuldUq7CN7ru6dnUoM3P+S0xCIPQfwad6Bmnv0+RdqeIN/yj1SRl0SiZfD6nYYrCA3f1XR+mCej
wPfsrj+owTo5P6UJbCG6sZg8ycdRUGL8mZRXcGauhpdaQbfgiPn1NUfME+aoLgRSbyh3UsxYcAvT
1t6VB92zGn5HSBgy0gUF1m/NjUIacfee5sO9mH1JrBrawoIEuNaIx1+Dy/gYO6dMOjgArfKwvqa7
0eIZxREb1ENzer/eVloGUYViysX68qIPqR3u7UHHpCuM5ifQgKtaEFAt0TpKUDI7IWecOL3oXQ7l
7nuR6CVxYcfDLQM1fUBn2Oda7hgJnbjdsLSW+/hs1wW7F+f6yqsNu9qmjbjOCg6TRXt3evPEwRKX
hoeJegePAvvQa4c6QBYA01auevaClxGhV7wVgcjZ2WGuO2MUsT7dXRpKnlbxfYRyUltw7tGqTTY0
5QLOp0OTkuHKWr9Bu6ZDloUUm8mMtvVFjwkJy8ov3mnkjoB06r0XOadRJPI1l1dBNkM2V63iFZzK
CtV8d0oNnxmH72ew0CO+Lblksdkrp7wn0B5B8uGCHdMZBQkmmw5jEA+lT7xlaRZP0c2uV0Udd8c3
D772ZyujlF5dD22XYE5mq8HQsmpNa1A7UeZfTEDvmo92ZuncT/G6YO2ngrHj3l/wfqtCGewzxwjC
SwynYbCTqOQRfWF4Hb/C5EEdJVKbVKLrabYyOog6im/Vl/Y3NeAhtMUn5VPDQdsAAfVue2DCGJcQ
7ssFCUpkDNpnDc+RWIugKOc/JJH0z4T7dKtQh/niE1pFb14eUMn6cgul1gHMwc+jcOydpN5uJEko
wwg+9g3khWY2SQSMPyPSGMIQ2ArKr9xkoERO0sOa1VNa47cSLTINn3fYzO62zind8VMX9wQMuifZ
2W4SbEPakcIwaxSoTOFDZ/0UCPvwbTi2ro4VlOBxQQoWo7EN6MKIcXIzkdwShfL4FosrWXKLGj7r
vYAhitww/q8hzEW4S8Pon1XHTv/08p0hvXXm4dUUa1ZuYUBAWrnqAVzy1WcCGXeoyr7UVVMVMtEs
7Gm8KOrsJ/2ynhFGxTa0rCGz6SmZav17XjfSPAE6/XK5o2mRQYSzA9SAAvsyOIOdq87GEvd8svnp
NXhWrqyTBzEeu516flE0Ak1OPoboX/JYsxkQVzR1m820xKexHuFEhrvogTdAKP9ypQNaEW9Lt7BJ
9f66AYDckSC7UKQpTm0jMd1Q+JS34e//ce/b9rOZvA3ALDRIuFNVLMXbdpc/ZG51FFUG7gx4E/Bo
LiHAlozCRo9QG9NwpJCnMmCh1Qm/nnqDs6v+3t+4S9bEqmNyzH/jFlEcj9YIZuiihSZ9v879kE8X
3xaB87EMTstOkyPLQzLR+c3Bzlk8q25thtZdsvPlRm7bLdTLwElD2Sx/4DHwAMyh/p1ili3xmrYf
AHkTaZcCEDFKqImv6z1d3vKRDyNdmS0h/MLzQU3IOD7B0XW0PjyHTEb1dc7XFqB3VggWSko5c3Fu
VUCCBR5LGx/Nn2ByqGeDqCLQ6EO+jBxfYDBxZ6Wl9GJPr7UPkaFN1SQNugLqhswYc/866NpnMtSg
zIjn+fyVoQhHxjxJ9bI5axbgZIRKVAllzArBBDChMqzILq0SKUwyJQN9fLlAnkWdapuYli9VSHdJ
GQBn7qt7mNhu2MFe+qnvgmbJLAZ1qXX7o8dWOCmbZtL3jmx5gYC2IXvxKN7xiL3cdjw7bc+PfKr7
ybZF1d8NzqfR6akiDf2PxZiXhWa0scVMW9iOBb/S+czZrbXQlV5VEx3aE71imir/R7K9sQXiWF4A
u3myaOJsKuj6z5yDTXCW6fUPaaooDmuvbqpR4WX5JyO3lhi26rtPOSufWRhZHCh33WKxigbarRiv
w/SV33PUqX5A2R2HSxcf0v2XFc+eNMc+RdCeTT7/9dphtT5T0y0sx2etmVUcEb3qvPqMM6ZBZsPn
HkuckF1a92520AzAHr5UQ0udsiFsvFVWMb4HF3/waIJaGey2agvmrZMlqGZmHtYm7J0+O8sVL0GZ
5RWzXklyGLyU/IioSuzEr2+amXEfl6vy4mQXYuVszFKsoVw4Tt1VIlFq8hagX7hzZTph1rlEwcjy
CjVkIR1ZDa4pxcIhl1AZrLXSQi8gjNik+e/F0vvmATfxACfGrSiVDAopMjw9Bc8aIQQcnf5x+waV
GCRJGSHv8YjymAFOz04q3Bo6/AMPKNi7fsF0kDOFnQgPvJA8/N5fK22xoRw0SHrN2vpw8HByeR2z
Jruz8yHIQNSnoq+iDPu0pkDmXJhyJNtwKscx3lwOgNDeuAMGJd6mm+h6sQI5+MFXXBdcC4rUDeab
ediGbYWVN27Le91PyJdLvKJuT8hkQzDK/0V5Zlg5H2XjR/EYJreWurcNefw4lwNNcIatKzJVSH1j
a8D9Gp8A3IQU/glsh26PuyBedVAiLed47z92mTq/zyPgiFEqE0JsNvS9EgeYTpE51q1ZafMsR4BY
kFC9B1eYm/M6PNnm3lRVjXBr6cHhmQGyt9F6QBnp7dYMlC51MVGE4mVU3mai4JxaSpFNNg/SDX4D
LYMp5I7G/q7K4b6YObsU/lY7UEQgOyNjgFwocXbzMPgXopTkKUz0bLMoeUyGteYPwCfQYI5pP3i8
xYbELVsHeZAjXdQaVyAFVqR1yJf9V4ygYExuFayRuZuH+Q9yCoL8iKbYwYm6M8xwj9IVxflFjLH+
sJpQqcXnmZ1kUDkjSpRFGL4HyJJ8IJjBaezUQAGvwgifd3Gv3IlwD1CazDHILrMMcW95V0cHTyn5
QcUdLMPGlqZ4lVeMhiVpotJ7tiiYiiEPOwv/Y9CB291gv8KmCaDhqr6opgiPo7iKmo8PmzBNk7Q+
+IlI7VI0yYc1DXnNDG7d9ZH/5Zr/OmxGsjWMD/yiwkuqR5paovvXDcQQz+KKyIq7NjSlmEoTvvO+
op7SIrbLeFCbhhINW/dl+6jXmyikSygMObgS4YkHhJQqmcFLvBX7kwyrhQDqGeTD4QNwNq7e5QmE
19czD/X+VrEIoLbylN4O7oyIR/G5vrkPYf2MEDqxvKhW/l+QE/Drh7D0VTjpGlzo4jKPTskzYWno
8pYvXVB4Sq35SJaSgpB8+ZLFYKbLIlgIBG6V+T0BGTo6M1ONpwdpJy8blhm5cXp/UMlvucOPm5uO
BXHX42df2tWIke1DRm1m5aU9fNp6FRIYcRTJK5SZd5xrcAaHBBDnUKBr69HHSyQlb1iUaLjGrryj
LkelwdLdPtV+LV5XM2u3RyUbDcdNm4QqIo6HpLREskUsBnxxChFmw94OivEbN7wIutO53Q1Xql2t
0sO4ky0JbCe30neOpYswI2vSE15WoNxJzL9ILmL5fKcNKXtCHIkLTkeTCpcGW16xa+Sdeq6gSPJc
lY/zuq0r5LNPLktuHXNE0hDrlb3rez7y/FNCTY7k/sp8QzIM74lykUawX4NWLARAlV+qZS0VLDg9
AmKI8ZUum23jUrQ+igUfWX5RJ2R5p0YLHX3g6dMpFtu5r5E32LXFZTjppX0OutHrx60BzebOooW/
yxh3jyyfGALTsWlfoTHJrN/hd/KaDNAPLR9rGVPkckFGzsipog+u8BEo4gh0O1B6oPme+rILFbrL
tgiC5BXzaiJ5xTBV7UgpfdrrQD6CyYSkrSGN0m4ahdPdFmrNT/QqPcPxEquSs4dMsG0JXlfqfwBw
vi82wXyrnGZFxaVLFX5Esn7F5dSjAr8dxwTVPS3xjWRBwpB/gNsTW2m/wTNKJNCQnCbyDKMKm7U0
kSwIHAVYLXZaBhQp5li6OBxj5cCkn9Zf7Y2Lg9gqM8inqVb9VeEKzAwLK/HarsIfl6gP0VMmJuPl
acXTSx7+WwNSXcf8Yuh4vZ73r2XaowMkCkOzE4J7/V35nEhHC2rJjXfhhxiqekucwk+dG78G+h6U
2jMaHfUwG/f5GNQ+X0FZb90bkaVSWV5u/sEeURe2llOR+KSop3gNyO2dkm5tevxI+xRzfR7j64DE
uWDVR9xhW/nFBQQmZvQXtZIagKRtqjRrgl+D7bixNnzenuN13Ygi4wALVpdq5C51U0KZd/CA/7J+
uPXyUxZUY6aQKyR3a5DW/2xupzY4IKDcVpBiKDXfSbX9MLntZZ8M5p2u+fXanYoR94t6dJwUaXC5
xnpIZ2CSFfgnZyXguYPAMQhYCdvr+1i0EraUZgHfmBLxjNPeiCyRmMM8O7pETCbdXR4sSqmFC1E0
g4A7YHbBZuhB5ciYtyxgJM/i+PiIxHahlO12d68mt1HsNV96u/khqhnayHSi20v91W2BxhcdkuNT
Jd+i/mtfkBwb8U8Zma9fulKBqwKwAk0K158dvkiXGRe4umh9HsUWTIJkqHU4P/BvsIS9itqhDxh2
d+iYjNtxobFZC069/YNtPG2CghnM2BSJFmGYDSOPiiMZrAtY7eGfkCdwAapQ2ODHj2vR3TkpEyVG
m6QtCUw46/1VKqx+h4bpRDZK06Q2n72yXskHy/dFtKBzAvoCwbQfinrc3P9Dzh20eDLrEWKVPMJ6
TeMUOBbQM8utUVXPr5O/I4Fn7WTGG2Xyj3B0yM3+aGs2JLGXvJ3LHstS+BLmSQdGcrmmuY5Xkz6l
rdLC44nLzp742qxZiGlEeaN4fPgmb0t92mrrgnZ0VzPo8SkaujYBq3DpHdUoafvWFJmpzyFcFx6o
QKNLv3WvAEhrZZ4uxiqU6DUvrffTYSkdofVPHIyGu/2APiQbysaMQLkP/uqWAc8fy8toAg04ZKa3
+7Ry4zV8K1n9nRXA/21auRMGAgyff0qpp46DwODjOlHX7WC6EzqiBHnCAp+NVM/JuHwCBnWZXYOK
xiVqe7tiflVC8V6izS7Ny21wz2oZTtKT0lBRX2wKESMR1mY7vZHIUb9tB062LvAQWDno8Nf/D7V9
mViC0bXkXKpKaTKaLptlab5XIg6kAnVVbWTW0KBGppkDJeosNNSj6tD3K0gUD/eA3wCbP1VznMO2
mmPNlLV2sol3HPIiUfd6WyW/25jvZQINRIGKplT6xoUbCbbeJ39tMAXyqPAqS8v6JpLnva1ykRhj
p+gmuutMeajatmCbgwp1CGNy5gYy/mj2t1zERhKWeHdtozi0OvvB76NSTiakkczQCebFMj42dBaC
4y/tMi5rwKrE7zxDcYKsBya/KOyuprX9HmxbahW7lJg+xEHBH4mqRwbd3qj9DkiNShfFzP2XJtNF
jznHD9Np8C36RzdjGT9jHahP8YkivJRTqNvDMyqxQiUPuLDg7m0znY9hXuxxagNs4K0rrPg/KapB
TQUdLB9hhgwAI7E5tluMO2ECusoi+zK21SAXqCRjZ3IChbFc562XQ9KPtgGtxW/e0nEdfolkbEbC
GJugw4KbcuN0jpKDrMykwvPRuRpG3kQySCIdGfRNG1Ahg6WWylTADWGYqc77b7Ws3HWs1sd/t3zw
6v44iB87+5FowAcvac/f7TRXcHNtSxsch3dwPxN7YEuTdroEnMb/YiEmdNwEdx21ZpF6u7/iQdtQ
etYw/2pR+QJsrs2CZdHzNcrMmOsUaOVdeZK7GFOjXyTX8K77iQY+R4LX2pMWMt7J8fyG+DLnCf7s
5PxwF90dpi0nQo84DX4O6hwFbgeKhIrz3boSedvtpBdTwcHlimxIf+SCFvLtmUgIsYbY+ls5Dd9S
8lX7H1jzm5ZI6MGPv/5fqFTNnddRLTalRNBRYOAziCh+dFLWraFfz0qzj8+N8AIh51z95N0PJukU
NWHykgzp+je1is9kQzwvzid8KZ38/uyMQEAxDo6lN2CRTJooMx4CJaZkk+6DL0Wm/wcf+aIu38sn
YowiFV44vvTc0TTCDO6XjjsI8KcIS8LcvPCu4/W3YLesSWcVPBolqtk5NosBFn0xcCwhq8KLcRMG
cIuZm/7e8ObrJ9GjyfVJ0PyiN7i5kY66xEjHz64gpSNu2rOChSBu/EvdGLm/aJergX/1HrfNeHaj
698Pd+fYgQf6Xu/jP12da6iSl0u8eFvlNcfFB25/2ducAXVmKE5lJOlXfhKJ1t3vqkBv2GAxYGpC
HF01gD3/obvp/o+NZY2KNTbbOwrP4dH9mAgGZ7Fsizla5uD2hsj2g9IetbvQY25J00EqPKTzRefc
O0YW/1qTh1b9vVdxGC2lXU+CkLzv7X7gDvwDZej6SiNxCDS8UCsEZhsTQlZ8pScwJa0oWM/0L2e0
hY5zpsW5JhAYwjg7ZY9D/jI0Ri2IAyWY3JWwEvDv+K1Moe5A5EJ0cm5y9BCBgSIRG9MuTywFFyGE
s0IT+JwyGyi12eeCCnuoAanIFv/sKCUpZ7PvctIxtR6ZqldW746Ssdv11w9vGlnGF0yOnsJZqF/M
sAzg8+ZhN/g3RR7taHvwm0O4kWJlBVojiuR791uugjaGJphgLyb0XNxGZEa+gRS1V9Eg7tsjgKBi
foaT8fCOMmVmVhDgCTFBixgnkVFho4F9EZ9QBOVkCUkSm/+OMxfCb24AyCTLyw0iFSsGreUAqUVZ
D2rqdzgdm+fF9hcXOk0mdySdP7rJFWRpIAKifFNK73sfOluWIG0mcZtIqKIa298raOnjc0B1VCoq
JRiq/4UhTEAo9eq86RcKnoKaSMQKhfOQ/DFoIPKnhYLxaC0mm9/VWscCRuj09qniVOs9BaTux39O
KjalQ6Ttyygcb6eixAnE1E7cXjBI7M+YpNSeL5Wx8U+YP4ewRgLTJzLXPcFXZwVEiWgBgjIv+0/n
z1RbZGvI6IjqH1UPorOx2OUNivt9A+iTC0gMDwpcW5zbv4/JOSWyGdRyK5Ef5H0rl2WN0o4/1BWu
v7WFI4ZNH34YNOoY6S71n3BeRHNTgY4JS1hvyPJ2prLCqWUUuQXLEsqY7Byn37VVP5cP0Q8MrRgy
2TQ8Lf4jUW9TqKQWiGMY53voiDJwUJKkjYxjQ8AePIQYnNYIsqwXIFoRfO3cSF5sigN8PfxZ98SQ
j+0/VnI8K/x2hEhClX5gLmSklIDUbj9voGNEg93CkpWP0KHYx0BdMKj8EaucCsuUGvb9Aj8RHvCH
2bxtPV5aFFigIdWgiZKVJ3KSwCbYDh/1lIbhJHVpicwm6ZlX226GAHmHoZDYt5LxLqpnasxOSm8m
8aT1OUsh1aY588Bc1px8aRCzuEYPRmAB2EzakPk3Ufv5oZGAc+rDhPbqZQPoSQEnjNCaWVvPNo7b
JECbhiXBtGOQOSLoiCwerjPBLolcTbB9QYI55fPslYRVQIYBCN75lcX/UnqFX7DsgHNWtQKedC4S
p/6Pdw610NHF6scp821rjBzsaKs4w0aQI8ojOP46G9zLD8M6n6ZvOXSqOp36yKSfz0Dqctt3c3vF
DKu6ZDkUqeJbJ4/58FAWAR7RW7LwRE4vRlNwM9mPw8TDt93HAnPbuyplO3WousJCvbygUvUr5McO
oVz6SlTolAJiddrfhE6xw3pxZcPS/DFj8e0JwBJuQinVgjk6H/H2WL2i0Ecl/BXvo67UvqHDQGxm
EKIiM+S1UEKKGnjMOAWGeyq+aw6Qm4qPIJi+2Nll9gGx8GEc9kAljeaeV7Le/UYMXMAsWhtINRPh
Yb0IE/LsyvN60LfFRAlbCcCmG5j91OV01w4WQyJxjh4LTRhXeLDjniZ130HFJdEJpQYZ1Qjw9QEV
2EJpCP4vpOC5LjL1GLGL9E/PiTOuRiME8ArvqECandGjgmmwD9YSqAURu352mhX431bVKOD8adLO
QrXOEOQe6CxRYPd3O8EobZIxPn0M2b8sutOII4AJACxqYrra2PUUk0pD/zciseyaiXcVf6M+uFe8
Ppb6i9lirdUijvkhRbYNY0ECgfRo/lZUfHtWA0u1rW99nEqrveqTpQJHgj/VKhlfng1RcCwoyrBR
Y3iSwcd5gTjuJunsdEYt5d6q2RL09cmxM78wfcF1SPFXfGKG192sJlfV/pZvKEzQNSRcBzke0MiU
9UpKWgXx7GQcjtGX5HAUemMChr8Z8hu1JitO/Zh6OUD8f4iJQj5aWV92LLXKdi9eSZRB3yeQAHZZ
ij8+EeyfV70+rnXENqO3FgB1MeDZ+tCFDrrvO+R7lBMdzsJRlBdt1arISOtlOpwobAy3LphU5jSy
Nvv2oSobOCZWCwzZx6Dkdrc+XPdVSpfC0w7GHt+ZSAZR50vOxzmigBXzWmz848wcYCTCJLoGIYkz
vDONaU/sFnWG/yA8ZTcmEdwFzHryD/O8AZzix7/o4Ob2rXYWs7cIN9wYmWOH2umDPOx/1LQCFmjS
ebZ8Tengkbqv+86A6+Oh5M4FLU8Tav9kCaTfTJDOca8fXLHrCzp5fRsXl7pjquoitbsUmYlLJVi2
PkMeKgXmoj/fg21vKtvs+VLeZw/rzld/yIPZ4dCLd0/sR15cLgWtn1PZNVSWkewIBxPLGKaBmLyq
U6ekyXaT7U3ydUPfZNf0IVsCvK4C0tblxLaXcgr/4mihMj6Jk0tae3+/TBR+VSqdxh7jlc02Lwky
m2TUaABTyT25+Xh93o4TJHJ+GcnwYlOYNo/XQkw6EXG+w+O7nCU83J2pom0KQxZNCEv0a/brRHKM
nvuazZ6ONeAGVsxf7qMU0cf46i+PzOriLk9AJLq5yUrFb7sXS3dazoOHFP+/sBZKuKUExkhRXGrv
HLCu8ewhwi0bJB1zVYK69H4ZOWat4HxNz03qMwJYbJ4T5qR3I+uvgUH0C+q/O3t9uHBjrM7Lnvyc
ZF0jUn6u3KVcTqrTDxQMmvYzSNDgYBL7VIPYrclAFrOJi2VeE36wtKkRFES5kw8CtyHHmy9qhTJw
0KVKzn5ZgkKHjJ3e1mOuY+6xGUkXz1FlQCUmQcXWUUf5dVoxBKlsCCwUPGz6YzbSCf6kUlI6suZ3
e73WS/CtXYaWlITmb6J69TzkYZUZl3WbybpvazC5t+qkQrOimwGMuRHBW9/eglRFNrnXUSetNZ64
a7wlHrGM71ND9Lr3Nc+BjaT2LMNd6YxvllNaV8es1WtzbmYBmpGlWMUPqKirQ859re1wV6LqLpAU
wgyKwAOKzVZVINs6G0ObMtKPBXlkKWsCD023TM7lRVK4dVCXm2fyhEDa8+StN5Gx4Q8LZGS8VTTq
cGgsyESVv96dPPe9fJ7Kb0OH0+l/cPgQliS4y72j7p0psUzL+aT3+XrmNibZvCI0PM+iHuZNt7l6
3GPWQxrLxaqooVDkAAtqh6ab9bCBJyrfwN4EWJ3tLtQd4ccJfs6T6rq5CZ0lXjv2n8WxX6Q+XRud
hGA2lf5tyCDMIKuGxqGHcBY6xOkXRFpEqHQj70+1QiXLnmKwffAhhV8+GZGvBLMYYx8Eh7O28Oni
zB5fxJoxQLnoDXDfYBOif3ClaKsnwDWC3Up24lF/AV0qYRHE+Xt1slQtaVGfKs1GOZVj+/RjARrz
43eHOJGW3Fq84/++8Ng8saetaJrHGmflY4BagRDIgAqkOPIj4+Bvf2217SLHygxXrTKjVL0FiGzO
rMKVhZFWkLBMEI8dxyZGx8QB7d+QCChkxLJvnC8T6mjJL7dWtO2B/DzTgVxiOIHZY5iX+qtYeC4l
B22qBD0UkIpKOgDXXa0/W0VZ79ZN5NosXDNm0QNN3UQouBuldFHYtPJLdxNQ0kWh3JbTFi3Exd9H
+MBwRwyCQzfkMV5kDjneBd3bAHtkvrmtG1EhQVD+rXc4h8Gbf1JnI8qVIaK/6EaUcpqFVBrXPDAv
hOxKfYuvFPDtOOhpmSl5SCYWUEk9OGTAH4ADScwaOSfzR0OV1pp594yoODwc1TOAamtqeFjxghvK
o7a1Ci7EAkCiYiD4s7oul8H/1k4vQiTQXGizFwqBWVHph4Tt0EB0DTWwLwodN5ZRmenuDInd3P9+
3Egqcg4NnIkjtAPF4exDHyIEmFvjancuNCb7RsoRHbAi54JAnGOmCacm5mAR8kvbczQdEbtjovgW
i17CT3pWGXSZ9AJzNUdfHBYmZIpBjTP2WjcGeOirO2ylyNLlzQkuhmWnTJt/6MNhIYUsGjPkhU8V
ldoDzosLLHq4cFdsezqTLTUe7EC6mFhRB2iJd5mPa47tDpZEIxuNFZp9WdHfSlf0zBK7bHs1Ahs8
gCnDnqpPzzVe6bhFJT0XCypkpix8+JKlNuXZcjm1Ias/MsrWzZ2FJHRrqUCbqrs/tWBfKcTS7TAQ
Kn3UcRx0ML7MX7eG4a53EOjoT3aj2i57erLlgARPR0ofzOAYE6IJ5NcxUNNQ/p4ETAzr9OYbT2Fo
6y1RFx/+w0FwRwjsIwS0nnng5ooVbANUVpPSgQbmyuTteEJ51x3JhTC+cdEG1csubYLMhyVMd+dy
oyA5wHFELL6RAIfI5Oja0mHIbTvE7vgcxVM2tHlGx1QNPAqFl51BVeXG5kRGFFQDOCtEUVspeOOH
2eGTzKw9SllMzvj4wxsW5VHhwPYTTCfWieNUEYD0UhwFmjkx0ljcSdOmzENuAVP7uZwFVu/Ffplv
9yWVVHeDYFffoGRuyE2icG4UWeb7zSGfgOJYxRiWec+sy/dqssb18B6z1o3dDR8B5rRMxrhXxKkz
OIYSSDuLrbQ0EdXxFqtX8qaYbuPslhaTIKx8bZfZ+ZFhOgwX8pV60Ezkvk0869XnQ/v7aip41I65
LU+uxzCs3T2WdzWfCbqoU2UkdV7vCB9IcUZ5M28ioydy2ayQDgyyjNqBeMk7l95IuiXvDPPGIBj/
PM0TG3wfZ4g8HKUyLLv5+GBxRpYCHndexAi4lolU+IA7bWEIjPwgTASBNZEXcmFfpGHnLGqj7vzM
Yw5dCE6V6fQOFYSbC+Az2VVZ4NJS50UlutGbKbtUfUn+iEYq7u7bXKAalUEX07YaAsX8AbWYwQqR
mbV65KwZGpDLr8WdIogBcoHYYmvdEpDQmAaD3bDMboOH6dWXR7bpySjh6HLVayYuTCIMJFbqYkGI
d2SUp82xeg3QhUlZ+2ukd0W8CqgMI//qdnivSQGoylmHSPjCeIhLJKXwT95nlqdeap9rcmauRex4
Gx7Hn7NBtwAz+Yq/DYxVpVnhDT9ysauwUPp4n4w2NG6Imc4dv79GZsUxIptRPCfxmGw4gwQV/Bbb
7z8Mhj8ABFi7GDqr1SQGlSU3VD+XzLm5nIeHdj9JsBiLmOKZuIx0AJqPsi4erNozQAbkNAX64hpx
JB8OXnV6slMiS6NacqWjRX+CmZGM3ZC60POPj6tItXXFEou9QW3zsiAeaclchbKViy7cdnk3ROYI
J+LKF/XTEzYqpvxqNYOcXSpkPzp/Igx/5mQBw0B+i5Mekul8hnsBRAo4kC1k2lSaaatPsrFxMG0W
zf9t7h1GPxvrjdbMGB2qYvF6OsJD7kjmsTx8s0iQ0sDsn/Ya4yJk/HgFd1fi143TtLS8EpwIWzQu
AbuhNiTy2JFhoCqhK/8PxZuPDh8PqJcowhNGYwlpcjT6bOjyovrzUWeXey5fmONgY0RPSXPfBs+W
UjQVxcmP8o1xRnnJDO+rA/FXhFMtGwQHMcbKtSG6/zTZRLS5ZnXWdi78JLJYQhOTcYTZaTwkBuhG
sTJLDyjl0pzWZ7o7jTHsfkAuITFxe/csD/JtswjvOPAgEJ8nEb5ZPoEBahEEV7h/jOslv9ox42hc
TU+i4+axMHaVJSw55N5tDfia9TyIc0h6lEfAebKr91N8afNoQ/8duBxpDBHOcyOCh3JxGYBRGcYZ
BoMdzxTo2DbMwQVDvMBnNLhHic4jS3dUACkZA31LMKdpVmfhjxK1Hy0eh4nteUZsqykWSUHpG73T
yxLoa3WCsPYRZQKuN6MmZR8jBQdcvDktk+H8uCmmjfCtrDvPHVGwOx7Qn3Ay2ecVt8l45pZm+QX5
NOHGVsNgtjX8IbikcwMsojrbKOQEzg+E7uE8MOF2cLMkwx3MegUK0+i7bMGmOjRjbkAhoCq1AVv4
sMclRVKJALHSKaNDphIqeuq9qrVbn4MG09wq3kp2uhO/5xLPJKWhpf6d/JPCiEA584kzXBlJDsV5
zRGklBtg6aVnzInAi5+odyMgOVSTv6UB5yE+YPkg7HWeRPLvs+VxcHYChzRqsnyweEAaADKDsIkf
JnbDgNQslv2TGi2R7WGdDFUanRooMrluPLSBL6B3S/K6zmwMbgLU0hbXGKJ6o/iTMoFbe69IVpBt
u1pByRWLDUgAhluCMqDdeyVBFKL2UUFKnKHdxQpLN9kWC81AdBTey8sSiAdwimCnCY0EZd+y/iAs
HRa/j9hog/UcBdawGQSwfu6yZKkTg0Vv6SADbpBnbp3UMZRROQcMlDcJZv0gTBQRuHKqjhv5RJX/
N/FA22wmGyztihdnWb1JXEbU93t1RrpTEOTy8ayHaa76kuwZ4w5PqaoTpTZZfMVYDPg6n1Wf8WvX
d1/SvUvizpKOR3Pb9va9J9o1rLmHig5xZCuxgMXj6f8TfkOTci7jHIhENCxSqaGSugFPNJKgv8Nu
k3QXAZybcQuQ7n7qvqAPRUQk+AUQoz4lIC4vIpqM2UbjeuxvTTc+ai9WtFV2JO/vnv9TtkszIJjq
02QsPBQD4Y2VXk0jE/PWK+XCxv6dJszbdWK2AM5EnuzCvbU1bSPOlfXRIY3DWReM1hrZUyH1QAhW
pYci/04OIBLfIkrTrwCeZ30gNkpUmE7bUBefFJ+3ynqSKFtUNqOZp5TH1K4N13MAVVCoaSuPG34z
T6nlPNyh5AJ9CC45nyVQyAMHrdFdacLFxkLr+MbSZEjKvGPPStAQ7A/L8qNZ5iHCeawdaqq8wtEN
X4qgmrjZDyCJzgOZqONhDwx2lz7VPU3c+z1rMzKRQh0oimI9qi3ZuKhTjlTLpgw7IuyHxLTsjGOE
KA2ZH7IkR201m7xfQ2VwqWdM4I9xkNwTF7HfUj3ShbCGcI2jKQ5ZuMRuO3alAreid6Z1kcg45N5i
BpuO9q0Y4cNMZkqkaBgU2pYC2N2btxSk5/W7qnNyI+9tlJQ6gd95GsWH5pbz+y0/e/DZiZZQaJlp
FTfcPM1lsFLU4HirJKZuipTf+Cz6FW82Hn3p7OBabeS9AKG0Xgzu4RxuxT9Fz1j8gNJcrZcBKBnJ
aV2VLkJA1MDRoFBqd58IaQRcdRtJ7DtXxZLgw6P6HjxmYDQTIbUUgE1LjRpF2tK4dvRNj9KbYUKQ
M1P3FdjzYvIn+REQs9FNLWUKE5l/0XJwljnm4pnCc80KUYiNssBhAtedj4v5bR5CYGZw4si8/7cC
Pu4bs0NwUC2+yfOXNP5cCelDmWD+AvCocrGkuyEa9j1/QtAK9RScZY5a05lPwu+7yJhBpvHkmamD
dimEHdg06HmPdB77KLdikzenknA8ihDsIAr+EJRaAWlY5aIqYd+/4Q3GFjYoUTCEg+IqJ2DOOWP2
alX8bAxjDkkPTr+MJrcyF8KKN6V3ckIf1xwzogl627gnEa+M+r6YTfsenVE8dlYk8cxuBN2biUY+
SKDJJQSCEhP+HDHpgPCK5FzpXge21dFHZnR7Ao+6HcBmylodDca1N2OWXmyw8JIhuH9vDUXV4VoP
KFI2YHjEvA3+AU3rsZx3W70FiMQdhVGI+SOhyoag508Tm7u5ZTwPNmfQhVxxcVpr7v5jwlQ+8CfP
x7AklLPaXP8fgSFxmTqLlbLlvCIE0+J4SLHSk5vsXX0nzo/qHkEWjfdZQPgfvb2YNWF0UeuuhlUa
BnHA4vWAVwN/A4utK1COhBvhNzNoaAm0QMfLPvlqafoZ4wvslQCmxzHeXkY030tWV4VJGV2Hd4at
ZRLHCnJHoPVNdpVOLZO7RjLCVa8k9E1fBaB9/IEvAW2VPRYlcp0YJylO4Qy3xE/0ldHvMJvP5PCP
RX9XXsLWpAsJRgKT3mMRK3tHS6od4MPvKU7S+ZmHwfduh/FBoqBUpGcZtgg31KyY1xMCJumiZr9v
ZVDxtv2a2jAts0O0kVspqgaTYfBgBJCqWzsBXrqrBXuuJdPb2XlTELz4HtYlOv6qBgHqyBsFYBDM
oDQtxnazKUTJ3A16zuO5SLsM99Rv5erx/pQHq0Lb0rNclnQMJuJJRaS3+KphcxGRAuJni7g1d3QL
57ZYhZhY1eg2coiMChCaVf5Dr3i3C9FeW3lisq5LpcYs5Mwn3ZykNvza0SjBqGCtTQSe3cc0h1ck
I9amhOh64RAhfvyfDH9E/I8S2SGUhfWx7B58H+JItbvbwNBrCReZ8/+FtLi5KgwbdpWqQ7bfyS7T
2Nlhm1s+mPMCtQNrEq+Xopm0/ucZUSizuNzlSMZb1VWSa0aiRFUX5YUP0h8HEuVeMq01bfZyE8C1
QnNXh4Ri9VwfL3P7pUTAheuBzPoo/DYh5R+B9Bqn5qCkHWeMe6voD/m/uyvEUpsxXb4cFLRuW5SD
NYH1XkSg7SdlM7dqN2C8InLxWMl70XUOiKE4j1CQDH+TZDOlklWYMpbJLoMg/dx5CvzZYnaeL/JE
jKr16qz84hvelF4P0qcgxtLj8GmIGxN/ksS7uxw3BeBka/pwyOYUSeqcrTFcTWqDZhGLwQWJNghM
czJjrFEzCS+jblpleL6BQmM0OJQJapq/WKRifCBOiNJ5Y/gqgp1nfEi+/CpBt0diykTB4t4NUZEX
TkoYb499hvSK8LvOG6DhIcpb3WqIN3QNoO/MQdIXdhV8ijQdxDSVp9x0gdx3kxF5ZHaeLZvaOOXw
PctQdtcl0QaDK1jcOFAnb4G4t0Hh+n0JwuHirvovFzk5y2Pb2ms+QDl8XZBgz3iQkgra5HbZ6HKA
5k2lutmQeMWbqRXi3NEqegvVuXtP0PhlnvrJwPxil7LBJGnAtaB56eHeGLkqt9UZfyQT6PTn+UWY
qyZ1wp1yUoFDLlPmaZj/Z/VmGvCfgBrJoUpYJSXJOk9OS35ezbW653WcmJu/1q+CpcFmGNjH1Hyt
Hg5mHnMxzWL6rHrhZWKkgN3ZCuLSjftk7cXYy7fLWuHLnZfOmU7K9D3YSikwhIkeyeIKqlSMEPSH
b23SemSrxk6Na/dgKujIMGZeKtx7e5zGDdEAUPFPn9eXE9smeyEO02H5sHwaxtUP841+2SSExJ5Q
dj9dCaUjWuvKRMz2yWy6wmUG6uJlrrNea1V36uGdlt5e1TCBxreZyZy3WwvQhtnMRhaVIEkyx/IW
wVghOYrjxiWe5064fyMLdhcfeBk1RYsyweLbE4FyDRKwMUkY0dl3dAsYpK9rdfAZIRIOmu6bNkKn
WbQq7+Z7HUbVt+b5CFc/Z21ywfIg+0nEBN5cDcSMKqznPW5pRJd5NVXjCIMqvcKs5ROaZVQKOZFz
c40QPMuQf7DBDc0e+NYSyIMcrzaw5B03M9Rj+QK5unSZ5auBsOHeq9tbLhZbqS5AvNBR/YeOSK10
MVxsu+0KCueWV2JNdQr8JjiNn2Tyak7tXH8DqBwtP7FQwYqgTZmQ/YMLtkzuvx8z19GzdBLt4FMj
CUj7BMrKOFaGfq7GKrkt2R8/CxzGUzjZE1XTfDZcl/UZ/QKnks0fi8sZNwyQDzVWpBALjGbP/5iO
YwUd5/SHdqArvx3zm9LrSoicgwEN6vIiR0jM8W7ZM6Kbk1FMHh4lWPPl8TFnxXadkPnCIP15Xf8w
y00ahvY5nk+kpm9WXfu/FuDXuao+O2VwCnxBd3q06X3u56UYCqmHUFvDljuxmsJ65O5pL8ytVo+c
r9fBm/16OIfcP9Kzm+6fMNycj4/l5+nIAoWVIMJJ9wj34IOxxaxLUnhVzLZuEpWfHdiwL6jcLOdY
OBOoTrc80J4Dw8yPI5wQyUh6kR5xHjfUFf28HGj9ngzOcfZl4XeV8OPODIy5XtqgNSRJ07F6bV/8
61PkZlv2TRLO9rCFlkbsmoTRgASMtwMMVIMpCS3vqytrfei+w7uahRbgPs7Csz+FVTMtE61M6nep
uO9v9641MTJ2SjLfy+H4ABU8UWo240iPl3sbP5xHMlu+MCA6/lfaZMcIr7zztDWxGjXRL5CIgVbC
CRDKYdl3u7XgZjH2a2yrim7O7EnQBveap+Uu3hG7nO25x02s/V2mc4OaKr8NOgIiT2xPHkPra8Ct
xws8c3t8yfRGEvmCsQ/jiygLUWlzaPrGCCj8hvDPusIzEDXkFXkACWU3WtiBuUvT/rs+v56y8Kpx
twxyRiJvMkwDe71i0RftZkoJ4ZtZQlBZe7iFT09QXlcuQXbz9iCKp/a+qpSqWuzy3jMXcZiGI1Fq
W4gMdED1fXRYreiEsNsWvM5Lqr8Nrrmvcufi63XYCAwWFntyEXstdiYlKbb8E3IQiVjSQiFVzQ6A
B+8T1H8n3X8XWZKi0wTAsS5nx3GUhqIp0/A/UKQ22b84hjCTljmuMTSvHyRla3AgXFvgqbmsgnQk
Kk/Lm6zBgntyO+hdh+paNju/t9WhmZ9gTR5ATRgDbJKMP/ROyOs+XmCu0PZ/grSN1sQK+Hvr7nyx
x5Z60OojbtoOSQF8oKDC7nLrOajhzl5MHeRk+idRXPML0yOPPevRRVgu/BvBHET/58mG0LJrDsuP
S/APPlq3Wh9xaRNVgF2vKxbkl2ZdkkQ+r7IwHKzORF1RLHywG9pNdlXw8frUtO+0erISis2QSvFD
bx8w2rkALFg+eAVKU0vvzwutwsyPCmmV3XA9NmidksIhzZmsWAJEV1avpBKl1AdbOh8AuwxNW+ES
2Bx51bic8+8dMvq2mIpnlSGVktBW3Ckcl0aw1l7C099BNwbbOOugxuD4Kf9yK/A96W5YJ9Ie8i6a
DpdRT3uYADYwZX2FbWSh0c1UlDpEaCd1+yuckhjleJrCeq8V/BjnZo8MP3w6D8XODsRlxLuGbchr
piXDpwIWlWT0mdx294IAlKmVnXjxkK0xgkjXEhtuznoqNKxaKEIBW040pg3Jo+JSI6NGMIrMQ3S9
N1iS9O1SB6Bpjemwjj9UxpCmPVmcW36T9u7JCCU60jpycwbcfzWYfh/sXSZO6ow8ZhWN3Xkf+QXU
8QdtdJcPf21rBAvahanw6rZRStWeujIC7F9Mk6KZMECPsMLSGWsLBomm8UM6dcNoP3Eft6CJwebo
NC2r9n0c31UD5eCPh0vGcpLVng7vYsusoWTZtq1nlJy99RLdK2JpG4PtChdh8/6gFVABPfZxgBgy
M5mnUacRKdOGQcHdQ0oTUra2IkzGd/6GAikmqSP2VhNP6+DMryKpLJaS6T4nWUOjSP8IEiekAews
TC7pniTaGQV+hQvwRKGFbZfilNW4FFV52p5ryTzMj7VTtGNhZldfPbs76pITk9XHWP5pmjm7O4nc
xtVF5zep8KZtlxYoD4JAhNbduFLhYFCmUM6cwzSh3Wkp3XkwQHv1PpvxttRf+SGDZrq5x0qJXeHd
0P39TnQZ5ONN90rQ+aIr0hSoen9d/lL4YnlP4nkefDOzQ4CpLdbLfcvia+Fk//BYVkDIKENbxg5p
NeuaKi5a7Wy2brinuSa/6sfKqKQFtoXKuN+QYIu55gfTGD4l1fd+HWb+A6zQXIwz3SQIQ603XehY
jc7J1Bm3kzlmmc8tRVaWG8A+qkr7obHCwQ0dQ4sFjnUqMtvHWrN9g8+ThaX04XjhUX8EhfGTesPZ
4Xn7ptLrbCcYoWMlZGiRw0cwQasF+lspby4/m+bZgWM4X+l08r6v2vxJ+pCaEvQ/bdhLPFghll1G
71ff8xx+i1wlkfe2uO2xIFK9EmoKC4GnSVktVQzcpWPoIl+nDM6MGm20T6sSJ6AKlbdVWTYA3bai
A7AZEyYSmQiVfxP73bzN/PgmstOb3NYBymNTAk5ZpPGX8OYx/nFkNOiAWAI5tQeJClOfoEhLqEW+
Krc/BOnP/dl/6Dju9BGFhr7qR44FNg3JnGMQztrgw/Bog84eG8jghKJ/ZObXH0LsQfOMZw47ISgT
DXT0rQxhFc98NZfYhNs7zx9HFbTQZuksrsQAq8DzJ8H+AhgfpBL8C697bWzAltjm7X343VakDXAL
rCIK71KFzgHlzcjl2dMyfq16HWqkHpYZ+8NEGCqLSrbVOaNAZY08OZ1gHfrB3M+Yzmi6uACCvzLq
vAKNeN1MJGqD4/1XKgg3KvCpqpwdhdhOtsuBbHiVsqhzM4gR0kqESxCyekBIjHCQEYqT/qyqk3gz
4G2Aq+0t1SeslZdEIIkXDsho0d2KQI+lkecWic5GRzbyw7M5oRJ18unYK8/tBDEjq3oxnkkdkDUT
8ypVfzNOxiHNNXbTkCxKLcweytQeNj+O0U3lvdRy+t30NXh7qawfOhkpt0EGZGiKYmNTzqVkSC5J
BPn9HDbLd8aoUSia02Qku8zcHbKXcHcCQwVD9QvNbEYFMJee4r3dez0ws+j4MYcewk3Pl27okA6B
i9amz0u0K25Jng/wQABA5hPldxleTBcGsgAqST8IjqpMkl+osZlAopMIfD943o/BedNec1uE1njK
66FXtI/hHTySURNmL9yTCj/0yhCR3VrREYwHfMvJqEXaLDupk9I0ccRL3gRJYzS2asEeflRtheF+
NVLaqnUK3wti0P/1jt6GqLTcxG235kq7/t7HNvGCm5t2NF+aGPLJTlod690BPMQHnKsv6eCKsGh5
L/V1LcXmZ065ffrypg4ibaaCeN8MCkRmwv7h0VeQXFNWMIy/pdnh8rzNAtpTrYnfid7EkSuP70na
JIREyz0uCzunKzTCbV8TD1QLs64ABA41Dq1p59lk2vtRZA6VCInL7pL4ptvmL7UCC++wfyTNb5BQ
PLyr0OqK8OUQvHi9D9sMYd5dGAjLxOMlrIWyNlY/bJBqiDAlUFvxCxe30M5pNVkWaYGCeJp4lHxa
S/srFdETZeQAvXzPh8OxUshLkTFQgf+riK0giV6hUHwkRW3jX1jFWgX664zJTYxQjmzhpaaNOhPx
o5464LK33pB7cV7nY3BXpnKivE6kGn420bykJk2mJclra+iMKoBmWCEumszXsxFjAyVmfD5VYot0
k4iXBnb3q/HSy8qgdbvNm7v0AoofAO1IQ0A9UdfO/4sHT7K7mFZDd2FvDZQvhBeJtlRqV75kO9DO
Mb/pG8S1G0NgdoyAdUa9p7477cyS1SjaywT+HQM/uLJfgLs7mDq542GNow/8wUMQYwOXiXVm+D51
f7l2RN1ZM16QfaQ9AsUbg7aF05m1jh32O8tCemmgLFSx/7wmTlU2LMhfgsWGNzJyoy+S0ogbH71c
hvif3zqPFkmtPPcyg6qa7amNtSaLsPfi4FcLNmGvZBdXKwX8ek3AbPd+BlxY3D1cBQJZBso0blSR
p6VIYoBYLRstRUvnoIo3ZQzoWpRuYtJkZjqwxaPQ1Oi58oodqK6/GsrRVGXghkUvtZQo0L+XH1mk
21SiFjSeanVlttyvhwA6uFRBnQe14JKwa2zDgKyu41nQeOO/Gwd2V+qPhg1amKG/FD+o/0oEqxKW
RWs/xyK15Vw0Hux5E8k55iXaaHb46/2vlZKlr7oMsDCBv9ycwqgt9XYm3qh5RyQ4J+zIP+zhZCHD
cf2RgHuM1hbm6JUtBPV2LoCiwn7vzraWBGsgdqb71ueHTaM7n//BiNsjTuk+jgq35tsjTOsLkotM
2KyUN242M/VJHzEX68X3bo3w7a/D1en4CwowTpOZ2FesDJPEyjR7UKWWx/7PJG9tzOg8JNuZ1TT/
4T0BkdIvQGgDExPSQTSP8rfJMREJqAGBXR1EWjAg1cM1tZtUIQEkV5ZMr35cpHx7BpP/QuRZAsNB
1xx0GL8fJ8TqL6hO1xrWnNg5fGrdUslr8cs2gornUNiLLXfaRSLScTMH5vJ7kg0Rg7/N9HPrxMHi
87oAJlftcn2s+599sKOZKOaqGBgIpptxCz8+Y2/B94zDZUEJlquYGB3ezd21Q9PoOuKlBKf+zDDx
gaSDEu3T/90HcSLH8Qfh/ir3egSg0a4s04sRDW4UKG0ym3BLxfkI4FMnIwourjyn+TsDONm5Z5fE
8Xv7cBCIfHiJUib/mOXjwWAgKWn2RdROA9Op+7oQEq7s80jT65Q3B7/JUHfgsftDtkRUqMUZNarj
3KQS8sl/CC+2L/EcadoMxp2214oqUWn7jgYlwBnXnj23Di69qW7batu1y3fVP8ms01FxlEqvn1Ls
L+/SnmWxyNWZlxkiLDZi3DWTTFe5Oo8XKgDThllaWNSpJAP2p6ThE+aaQDWnzWLoeRo5UGj7Np9d
axyvsp7fjsl9ShmUm95e2/cO3e6mSbicpGRZI0RK4NcroSR3j9DQ9SFcMqjPuHK/pdUSHpeUyiul
wGQ6ocZpemWdCayWGRk8UsrcCnpB+7LLOziqVDDSnljCB6ywEtXRzZmcMz3065rww+frM+jFiP+E
Lm+pveFLVfZFWSx4kQQuSpVYoAPACRt73KHD+bfZIbbfmxhboMpKcS2zVQOXKrq5JAeGtO6UBSYH
8G0ZClP+IC8RBTbd7zLFmwgFLrAGMTL+EiirwHa5BtQkzJnQ52nw55CvLd1R3H69FCv8lvLS2YKx
aIgk9WeWSgdzLZ/Ez6or9TZTChlY252bFvijCXkiv2y2c6YSRLSFJ+rdkicmSe5FNdKxa1jZYnia
qgBBvHBACxDrqy5zTgflpRDidWRmF7R0rrWnhig3aWfh16ZXDbjx8TTFStkWBk7uDKcJ7cwG3Xtv
LtKAYN8tfTD8OnaANpqXrH65gCmSLC9BeS9/vTd/+3pVczVAY6+AvKIhFRfweRamB6ptvjJkRQgT
YegCVazl8p21x7BpK4j6OZTkDSrs0MV9VQrZB+YLkm1DGg4tz1B+dPuXbJ2Xnq2fJMTFzhl639YO
1sNTtLYUggVzg2vnuozuqTsvx0yPtyqTzTocxP8tvkhACfEYENZ6BFx3smmtUPYj2wo7WKZ0FxXs
pgZlNwKJIgix9+/+/IYFghkqBSSf0mAfE6sCBR8rfjAOGP/kb0t83bV7kovIhYo+eDKYfVP8XznK
PM7uTpwbqlXJrMdfl3hAXP+otCSWesXNJR0ZOCyN5LD9k5KWRNB5TJouPAoBjKCPwUHeTgGWED97
FJAFJisvyZARecFs6O982hoRvt0zmMQatrU1Hod3ePfeZwyWFX6+0N6kkFZOk87H1vTsdjeDjUZb
j9Jh4QSMCvArKu0RPA5JwINIC9R6cuqmjeyx46ome6RMZQYZ+hlBIucMqph6WY5KBDQnbyAQhdv3
LynsKa+nnlqMZfMiVEvgHMLxcjqiBTv2BcNGo5SkB+y5Wp91aGVtrf2ylG1X/0/359xXxJTIjqVX
GXH6pyiZMXgSScnDr5VhUZPJizEtwWEIhmdmO1WwdrXBH7zGiVWdJe7DOggCfCbOS7uzwl29zeAc
la3GSKXRvWm9vZOiwdzYaW9w+BxtUZlt86EHdUl/cF+SIZBOyec1kFJ3RUyJyTCvQ3yXCndZRcu8
EB1sAk8q4J+UUjvOf9Gllo6IOSaM/J6zONVmBKtnZNL6Few/X+cJwyV1V1V3Lc5Bk5eV5jsczGOk
w+tAdcEIxxsjsIIuYXtLqf6fqxbyn/UJwtBX8gO3V3vWpitLmLEGfb5CxZHXsW3IgxSxMP1r5TOu
wu+Bv39UXWx7rPz1ndrKhCWsp04DMa1rGPzg2IisEtMaTEkLjFaU+sHnemXxqN/XrFTvc4TqAyEb
kNEAmeQpXZVHLzzPzpXaXBs0wcLFdZlWIHqM/BWkYWS4Ewt/7WqKjhm0IT+otd86F8laA2L7XLb9
KduLR/d9A4mlpIOk8zF4RT7aKELuCFhn+5vtK42UaF98QbP1StDjdNyr9VjQbfaIJPpDwwu8xZxL
tKRgwlIVX0f0IJL5XXwHBNPLNQks2aQn6a2S2M1DuHKgaUP3fiXKfq0g6mHPMGh5tV061ZhCp3Z0
bRpCOKtp4fKTsiPDk8RHioy5KTAjxeHHs/2obLk2xqnrvEfIw7kOkDwoF0fVhIqrwdsQ8eCiPYBV
d96OXMQsUdn+um41L2pd5AxHFgKNe1L8nzSpMpmIT34BmNNEOfpj8jSeZ1lFY0QmyjQHHGTmpHMV
EtFL/oBDKK2TLuKVTJ3WNYuVJj9WS65OtKppP1ZjzNVQ1LtFishG41hNiW5MwzWZ3p4tvSQ+7c3e
5zOSNHXJi05YIPAiBlTEax9juSo/1tuoWoEMYHre237TXB1um7OtNUmgqsYjmPh4GHkExrEg4iA6
Wz/lrH8UefX5k1EjDerqoSqbvh3n8tEUHuxGLUsCaaqeji3hhAl9ZDp4HG/HS1pGMhWZj96eKtro
2BSrjLUeB6kOe4tFNTBEN/yZHea4Hj9ZQxO5PMvKn69AQTdtf1+3nyTwFS4av1vVjlcCH5F/xQuL
QcmDjNZu5KGtqM2jNHiCev9GWjegzbTfnnhUR9QM+UaNftkkwaZC+aHxD/Lln2/6BIwTvCb7AN1y
yXIQe5frTJNAG6qCLuv845U9jHBPQAhhHFhxNEZ5mDq72DxzEiox7St24na0RS6eaqjnDdAtUzKN
FnMClWH2xQP+Lr980ww3RAcDfrJ6bn969wO6FMhlFmX7fHrJu7SihiRj5CoxmV4rPYwCqM4CvM1f
t8eqnWXtC1QxTOnKlAj2u6lvIHseyalqFYCOlg/NWyiUs4xEAehY3/MQhGcnYN6dpWx1oWuEg47r
bJ2DKlAhmCDlyGmMQmH2AnOpqTYLp6jP7LSwuqkEkOwmeKQhwhxSxPQr+qlO7k0mqSfG8hy4YEHU
77SzKRIKIV8FVrPw9hqzEXPyTR6Cb3evzagcsfgjnU2aXF7y6W6oXt0FB6pIKa63uimelbDvY40C
cR4rItTLq7XEuIRExQ6wsGRwxUKn1wxbYgkOg0m45tNLmMOvFkI8BElTPIZThd9blioaR0hn+6bu
LkUQhkS12VpciJzYWCKcB2bJns/Do1BA/8y/5xgDbTSy5ZP5K1rfVyVocxvonFbxT2Fgje/t/q75
V4EEO6V2dwDikDPtK9J3CDgBjsFE0KlCIQ1Q08kJZgQInloc0dFTHNY5bYJIi1x0banbVXb5M38S
1RBRRFZPesZOS+5YQ6k/NAKUEx3stPEYjmOIPHQ4aXOGTQ14VkE6M1xtrCzjNlkNU1iqlrS34Zmi
ggmtoBino/bJ+2FWlGfmKVRC3J+p91Tg5/M5KtHOO+1d9uuC6jZe3YWVIUSPworP4JUKp8yfbScJ
ashleSQy/rn1CVvzmRfZhLraWNw5K6l7EsWvNOUHzKu5iQvmAJweKas2p8Sajmf3hVIGNobBg3ne
ISLRJJHFZAgvGUrU0hR0fU7LF7l/jWUasq0FuuVLUmoDPrPXEuGWPz85NBGEuiVdjPy+rBQ8aCKF
ZubwvAHCaymE74RgAZPLVZx6NUV9pvGR6+qQkPo+R12aaWo5wrb8h/SuRD3M3rt3ITcBdCcN76zR
m7bzAVg3YAJJ/++BuBdCZTuKsTdgyZpzPcyuZfo5KYEOELoGO3O08zHMcLgKhdJgD6iObupdPysb
29d2rkpd/aWBRz/bFbD3h2WXyfEUGTTrGPeNOEItufw1HQ1AWaHs9F6p1UzJ9rlIJQpLZ2AivF+7
KKgWOL+TPVLFFZsCHQWNIo3pIT1z+H5LVjq155D/XPHn5nx7cNWLKIuDORxqGuxshk16KMAAPG1Q
lT8Ryy4wbgizQ/sDVCOxmVhjw56pCtRmDliNZ7Ez4ecdLbMh6RRCxWRuC4sCTJXkElZGSFz7WZvc
LRRUf9ciV0DW1rOeqFwCpGVJsAy/gUlizKjR3gGF5J0ROnJr5YGNwq8GiYgAbTFO2C6xWWVKbRij
4mCs8edJnr5tcMXx7JKWPUYsh1KMqlhfToVVaTm1GnlwbsGu9O56PaLTFN/azp2fLUBM9EWmHTLK
oNY+ZAzkcAAB1mOC6Ez8OeuOtSZb3GRzEsV3Xh7ZJLNHLSPADmpoRimiJefR3dNl/UbMY9mq3J4b
UYrD7PNoflWpZ0M46jCv1D28OJ1rG0F1BmBPVuuPozbgeNElEnC6MSKKibFgKza7Wfml446ddqyF
Ht8X9pe95AcqbnjVfKy7IkbbEQVVm7huLlu81c4yRwYYs/aBfxbCq7Jy7yvK7Lt44Z/6m7T4w5HB
ZkmfK8wUWcVWzLWE1WHknzWr/4EZ1QZQADZQ6HOPZkbsfJPJKNZAreLB3KXOwJ6x51sIX1oU1Whg
8d2Q+VPoag1b7oOxlMQX50FqiX2eKtYGsAkYbaese3PGT3OPl5JZTKYo8E2wQyQDRSqvKOaKLOat
S/X2yz/vcKoXuadE8931XFi2AmiaZVOa+PRAW1RdWMW+WYnnEtkFnfBUur0u9rkfI5B9rFXyWYXY
HcL9cdj7WBKWgL8gB3wDy5GmhCezFDFoSNOuwMTZLwPujipl7sTQrLMivbTi+QQjxdM0l/Clms+l
Xdxrtf5YYeZxLwayHomS3iCI5EFyIopr1NDjSkdfsBwihx0CBDvuSP+ZHDbRWs8gzDytgdIt0oAC
fxfA6kHLTbxbJhFQnm9m116D18/2Jr9idF6L8JvRECinQorFLKhHO2A3TAHNmLEBU7gKVpWDTTZt
/A3vIgXM0v7yEJiN5QStmIBtzRm1OhYtYCIHg+9bnVfVUoyk4xuVx0X30WWltn3D6nfWXQbPFZ6U
la/ltQWyJTjca7/iW5lsC2fnvOYgOzcORnbOEeL3YiqP/9pMJDF2552GVTbjwOeUpUeiDOxXP0xk
JlCYw4Ip/eyMXMo33K6stTpR+G36FP7+ju2XeLaydLvzHVr5K/R9ajMYVAb8kOx30QUJgz1y3ZdG
DUm/uE4TdW/fkZHiiYThLc10Zp79WxhncOq+vvWqaonyXdokOZdgkZZBkf6gsTvWrDPVIIujrrb/
Aa6mlc9TcJKAYlUbxH+sj0LyomhrbJ8DXDleur8vceDWH+ZirmGBVbl86t4giefdvvW9bXKOg8Mh
Rwy5l3NbFL6gfKMqxKE3+NM5tdZzKV0wbrEsQj3lgBT5nQTiQIafe/75yMCGavsvB1L+Chva9won
uc0pfUOfxLM//vxvCKegL99TR323gnGbr/ZambCx5KdmN0rX/MxOXObk0L3vkR68kUJ7rQ74kINN
gWd90YevFI1CIkfGIT6xmY1iD8JkS1SQlhXnFRZ6acliJ36jvO6yHx0kkt3J3RTeXAi80Xphwzvc
xqsXIBBJRazuvc69PKQccngomoUbYkCWiFGV3tAYxG7X5SzaXUW1uNk6wElD2CkY1l7T0vzq4a5b
FSqzx1/W7uV9nxhuQBX6u7okKPsrwgnao5fGpO2BNtnP3+4m+s6HQaHacVnLnq368ATnkDpgyMWi
eJg5SLp7tN9rR02PHhoIQitBjpOsPXwodQSzyitOkifG8JmYCCyjzUrmokg1KLFmrn6f2aJIpCdG
lE7PwQa/mPyLHi7EuthJXnTSu6KNDwQoraIyQ5vkeu9TI7ZYvwngirwJXmVjp3hr4hIzf9JX1oXt
MTc27ce+Lp1fcyNxfV4k5gZMaHpT65L9Q/StzTUqabEuDQ2a/x83Zn3+R6S7QLJBAlRkGh0fefOP
IDEr+CJTztFqNUwGSFcr6OaK3U8tNVwWCU/NrYkMCtc6VrQi5bDCz1/7obQtvjq+FdjD8772JCIq
+tP5ZAfmnmTDiG0TEKFNQ+06sPnD4kuBvd7Y5u3/2ek5Wlm20fYgtog97fIEIM7MKfa5lAlL7kMA
mzgyeaX/VnVVmAusnlur9l7Fdulo0AI9EUmrYIwTD5l/x2fFIoANj/Cjzhxniyx+/6m1fpH9tWuD
q/ti2C1U0AZKmQioIZGMdZoqlQQAwpW0D/VRfn3cQ0SDrawLi122LRwrQmBk+z3lPYYazyBV82NZ
K2RF2HQOd004Hlk0rqP+iRa2y/aqyzZistJyltcgy1qmvLHbdaf8cvK3sfE6cGsJrBwTS/4xq5se
gG1Y5OdyWzE5J2aj0XxuKdtnIEUeQOeRDx17ISh58ZMmkGBTTKnFl0/qib6MrCXfbQJK9lNU11W3
6NJjxNX4VEuLBjQCNfUtjfYM3kvSKZMCrjpr/fQPyulCwKsnf0FJ5Bzx0n8hVDUBqzYSY0h88ckI
Yrf40CQti2NhqV81oGMB1/r0Hw2M3DbZkgYPPgi2aHrWNNJVqwACny6GYIHbeaq8mhjPtx5zituy
b8U1LT8KQx0Fqu9F/Jgg9TOBMU3ygWB6OGU7qkc13/owmHxluKUt3unLo2ei7FvhpQWv5TcgdqbA
8XTU3hvfD4262RlL8GGC2Ufj+zag1WmSQaD5CsILZCAU/h2tvli18pld5gYabOn1sYIb5mjPlJfK
Eep3+I9pdSEKtZbczxAHCxqTb6LLHZukbsaFGISHgDHHkCSyVLBafaU0c+3fLljRywoIGHVm4i34
cxCabRvSMn4FLgjs8s40s0xYJIRqOdeTm1ljQjVPQ8auuZ2+G/9v/t3lV/Nj+VhrgENGeLkthhOW
TCb+QRHXJzx4v4fKZvudMWL4dTvYwleQHkIuNSvn4jZkj01E4Bt960Suf0v+HK0mpPYJZJpHUI59
nIG4mWQWh4gSxsU1lPFIe1pav2DYatPoKErZHN4GkM9ptJHKSgZnuedgCnvm3Z/fz5qxZM28gx6q
PBt5G7ZUKjRKabMVHO/H7U2AIoelZzjR8rHir63+eBUVLCdQpD8iQ7SAsR/xn/eGQ73FASs6wYk/
liPgtogZncgQvlS9lkYjS9wZ4h0zp1VzXlix5KyBfSek4gpCkW4nI8nqiVBJvjajF7R76BfyKthO
dIgtGRgW45jMuO7IiSKf9Y3JVgfviBRGaskeAfmEE4coMi5hTZT7d4HcI67O4BhRwP1atUtd6cmu
iW9gaSsfZL4dWAunZSoQuXx2agwobjumtuOT/w/jlnyvOEHZHe/P61XCcT5hUcNB51uFnXd7mfes
gyJgTxOHEybm6WdG21xzPcTKUAO5lhZgRYzOVIkq3xrunzmPkRQemDtav9QaA8W3UMjC0OTraTTZ
uJnq/8/khROxIEkIgZfkajXZGFt7nIRY8TzxGRpulH0JkaeASCOS03nGsO5w5KoIuoZ2RRr+Gqsk
qT8Sml8lLQ5PQtn+yERWw+CRT2ibhp8razuC+/oDWOMcWPLra558nyfJZieUWC8nWRsF/K3HHZYR
CQrn4PWV+6rtA1kDCSk8vU2sJD4Jwybm2zGtQWSKJ2QQVMSsgErWQ+Psy998hUWewvg5XRYoNoU6
kQQwR0brvVTk8a9p17Lbl30/2/6rAlS8Jdebocb5SUBUIOu50u21oVjMzIR4dDUuUlIRKepgmosv
V48mlsH2w30bsM6zmsMw456xCBvTmAwew8o2EFBgsJ1T9X+5uistXmnoPD84lyWH268mD80Ztrnv
miaRAG2rnnyFbmxTHRBJgfZ4tYK8krfLOuRLlI1Tyycjqm9I0bN4jYsi3gmkUNZaZdlz0ozyMC6O
pmEURTIsp2DFSWbSh5V1AWEozu8D5w2e2RWd/EZIHH8JJkZ2fdAmHZVvq5ODCwG68w3/yLmiQO7T
WDGzcKIlOjXUgRHQ0s04/xfNZp1VMkU54RhWhRYHPCFgWfAvt6aI1IWSu0zVZvwM82TTNXrNxDeN
hIgnV5QMdVd/4GN4ySKFSMOpB/y+lsd29cgUmxjwySfTAFf6CwcV2x7GClrK6V/zLA9zcnZg4eoh
sYYQ/UL1klPfG95lT8W09kE/RAAejBeaK8sj4ycslSOJ9JOHhR5TEVnNuyvzqgxtx7pgsTMmVWiW
z2bAXqf6fmQv79+uzhuYW3U7BqfiLIgGEg0wQebgeOaDZTnTY9lXzfM2HJf7kVRe/scBoBwGQZbs
RnSpodbQ3FZU/pamr54ck6lXDY2n7QBzzISe2oGbN7MGQjkOKeTl8UVNraHgz4BX3YoX7gBTS/MX
MEaMqoMOrahzQYurIcMO19aQuEEPRZ2VlUeYrZ6wdDau+OKHh7FHOPatI++QOeDLrcq3TOEbIBn8
n6G+RIyhHqHRbrhBT5iQuIbpy2VAFpxAJGu33UXu2v/8iZ/UH1b5OWNkKId5ejFi4aTJl6SjvbbS
Xsxa0iMlR34KDePBtTBXt4+ElbyzlMZIDQpP/ih0FwE8apk19EiPCj2GpIjSQ9FFI0i/hkxqk3Ez
6CHWnD1fxp3K5IndrvMczCt6CzicfRsHZX0h2+FotO9gfjNTfQI/2t44xVZTU+O5+pN15d0EKpnv
goMUe6QqQVaKMh7XCNn8OTkLn+OIgNBOHU7f+BEYpGYJwBWl1GoK0HPHHKVeM5wZMErTamWc7AtN
Eay8u/dYD6W1aZfLzNQXWFCFD6JOlRy21r1Q7llrFjQeHPnEj7klCag8Te5/kJSXaErI8qPd5e+b
K8Vh7zY0OzAiQtn5QbY/xXYQC3g3AsIxtdY4uBBQ3UFubEcOsW0a0QsonhjSzEpjra42KtKGg8we
N0ve2QRqSTKwVPZ8t8Gk7Nd3x8+nPE8wP3zCHAhphI9LZvIPaGbEfN680uAS5NpSby6GMzP3nCxr
uaFgX9VKNGdlMUPaiN8uilRlsMdBr6i2cXTmNxgFtg2Z2RXcLzv569ya7xqIy3r1ZKIvTamSmVkO
o784Nowm97BycGGM8M95g/mPvlD5ZrXeW/Vo03qZ1LBixi2zLUb0Xbi89mBq9zgj4lrCyT+MSeC5
+3j/P7vS3CiHwlAe0sBjyyz5cBRqPLC2VcSByZw8aY+GwOjb/7GR2FLEs0I/Eda3MtQa2y/Meqsy
HMwDpi4Cj4wVocVXKsSpoZyavxYIRjF05fcN1fP4xUasbtJ0Hzh4kpzO1nG3Jshz+thWUad/IjIk
fINr6tTahA8z0Db2lT3eX0lHxQDFvn75ysWdZxw7Z5y4pruHjLi69ga+jSkiilGohGEqMgAdgDPW
cUMwANYVLuds0tg8NqYN6CmQ35o1IsFOlVasV6AcwPOCAgf2iGQGPje4oW++2l6Yflc1iKtK8gmv
uzeRF2zfpJTm5Skcgh+7Xz1THaf+DldDtIuCmvyz4Wga4NEXFKAqodfuaagPe5U4TiIq3fzT1z/p
WXpr8snpRaiztekzBzFLEJFHpon/C+AQBY37DU0vHK3ajDlQqdE+q/JTY7XJC0DQ27tpLdvAcf9l
zKFxg1d4dPHqCfmbPK8kLQm3jaIGjt937iJvoFMQQfw6UrSfG5Pvt3nZHYPL6FAEoXhS2VzoHuAh
9gRVa+K5Cau3590DdNdcB1aGWA6ib2KRJhhEs6otVMYlO/7F1cC3LzjVdLKlzzsPdK7SU/n1uHV2
siZ+CMOSJCUP5jP2FlZ4jNPi+xXBOQxhgZjiQjQVuxGRtAz8+MCeR2ufWOrrU5pl5YrqtJxAEipg
09d1PtDukhdh/lAJ4hT+/3U+a+Jn2q8C2bADhxlu/aVB5IaSDPU3dD5ugFwn+Wf12DgaFWToNWY+
chpej+4QC+wWxZ/Pte01lkfKuEDBBdU8DHEk5dPFEKG49kyQ0SudAjeQ8GCEchKJ1MnMQ9RYiln0
M42nrfASapImtA9QoIr4aiXcgd/OmXw4DU5OmC7QY+2KipjaBM3YJDtozxLQoXVH/9ht52oE7XFJ
XEtl5qDsFwaQK87vV0SoPSCJ2trqjYA7KEIM94u3BiZUmzdQCr6HLo7bjpXeZws01uxg0cwO35ci
vV0jMxatOAJHYXxdFCMbNcpLTwaBwnc2WgyKBGHBjkZBFlSe0Li3GTcpOAKBlvaqJJEl1JOCUQAx
3y0tK2xyzKzHf5D68Q5riwldUto7aa5g1uMKxjgYziORtSncFXsz15FaJ3DCTUuuIdxRuGPYm+aO
yUHlK8Tsa/qr8vQ52/h1DXV6g+PxqojrJhgkHnbAO2OyyMemtTXHyfLxB+to6UkWAVFc6QaYO4ti
7/WTT/9b1MqL6Rl8Who/2i3RuHHXuf/lHPIhAtnLdYssTLSCdzZSiYOJMJ6bdrnhU4pcFc+lFEuE
A4aU8vVK3afIAUqbyQHNexolyUlkUANn9BuQAvSq+QoeOFgkbOeiZ3Jl+VNe1uDcJjQTsRLyLI0i
2zPNdUwtCPE9HBsBS/65N60J+cwYlIJu86U5ltAaNF0abeHwuh2b8LWPz75UwarkpDO8ETx08BQj
CdqwMbN4BztwsL877H4jvNgNdG+IzE1Tj4jUQq8aKEx2cIHbu8NWStHYZ1bJ9oWglZI/m4IhZ9dh
Nnv1gwIDo3Fw1Dqx7OLI4/4haiwqglKArSkXyz6Bxpi0/zuyF7hjjtGNMR8i25zw60veq45wgNHr
r2bcURYO78JaNC4KDhIhDk32t7VS8rDmRznqLHV2+RKDzLxk2/li2bRSeZiW3/VAHm0BQVZCwH5g
xor/hzObxTyBwfMB1bsqToCbvlrnzW46Dp4dGMBhtrVEKT/NpMAwoqISNtAJtXJonU/gJ4CDwfex
zB03Ka2UmsVnWa/XodSWjl8JvH7ARy9a0mqZdTnIXlRDl9x1//TnaQxcgEN6IBIcZcZdT9FxXFfk
8yqJ6NEJd64sTg0Wp3bB28D3AVAzqwVlCNjrJkc04bmbJE2e4mEYvgmMy111kxnbcaicsHnaDtyv
5OW+zNogLNUcSVs6oy4zGpHZSmnFtNx7/e7wya4fb7kHEptH6uHYwLAekAZU7osEWnFKggSXasLw
AGjEZTA7S9hZ6JMMVQR/Jzyg94siKy7kHpiGtGp0XbIE5xuXp/WTa+8t0q9xFpyOnL0LHRpsXcbR
Nm6+pss8lDnsnBu1XAtAr7EzMAxbzkJ7EBsnpJ4DRaOgnn4PF2/qeCVjFSPBEKsv+lgLDqvU6LDN
HAxzJ05XluCFgPq9FYb2WfFaUchjALZHgRnIFX1t63ukc6en7D5hxP4ICel9WJxPrpTH+2QVpeQh
AKoUiRHChXKlK7TMv7bkKgEfeDQ6Iq+BujlgKf/1ZucORfMbo1dVEYv0ey3prpCNKeWyR9J/i4Ej
CV6eKDMKqlffUId64IejFVhzCvhQTdsjhApyqSmiR6ciC9DD+D2Lz/8IGSPCnLFQ9vwMp5u4aL11
yqIKwlvMilyup2geg5h+zwpxohgHblyBDILvcTyrh7S3BNotZdErx6WaJ2wSNDp3twogVfcUHRgX
pKrmmau/p9LcoDH/HJCxESAeIHc4S7rXP6mrF6twpLtinn8ApFuk/tJNig3tENU+ezKOWOw0O7Oi
VvI0tRv+hASFxmH5HYa+iHMZAHy9ihUG1mpvosxOB4V3IfwjMkGX4HDGhWr7/DTGpLGy86jJlEyW
FsBcvhwLlgTbUPiSfkcpKwGiLIHJzVB2HGmc0FGfVuXaMq4jG1w64LZqRHvahltMWFVlPqQJ3H93
HufgN8CTDqZmrhXLROYLk0ylheDxmuC5Z+vHxt6IAUlkHuysd3PX1TaUeWsn3oucTt7Fxp+yluCZ
RKckJoOuzZYeISLCu2CxbGO6aNVZ8BnWpG5HAGc68ngJqh2S8c7XwubfX9onB21HW7vnDy7Md+gc
CmTT8+iw9YqVWT0fTruQ7qW9DhNWWmJ0yGEFPOq9o1adht6Lvt+IghCGC+x58S779KQCyFP/m5fU
zBGYhQcT2dIcHZW+VllivGtdF75C5+kGTqDsswYxK8Alh0eY0uiU1AYxwuac8rTMaOFapLnvVw/S
JAJ/j3kKpxC3Syq9YDE1L55kjA20HBIPfxF+CMzc4LY7nJ1IjG55m5bo+NCTcTFTU3dRk5xFO6sM
lGDkZP7PeNAkTkwSvaquD7UGm9DqC9ObKtyynEzSgB0AC1q6toY+A6U/1QE0P+a4HXJmH9znZRVP
gc3u92CnEAXgTrB26Z3GDOEZWbtvh1NW9c0oSJXH/U0fU+zqNu2gxKU8xjvrKpEITDjZmwC7Yiss
4Xa4JWSTqWskpBqoXTvNwDHASwgk0LRdasOoNjDwGBqvtsWqLalzFwR5d2FggkGETJzl6xc5dJqW
Vn9ha9EnvGT/GPQxLpdoZhazYYImA4ft4UsoB6sNSD9a+GNOX2N9Bl75TtI4EVfH+agAyG/dlcaF
W4guvrhCwmvKXQdGrhwLIaOgq0OrT0xVraFuGSC14dPeYXqXpMISSnVS6Rb7j/k66YDSwbIG9bY4
ZzUwPn4lyKJMHAZwnCLAwz3LmIfV6Lf/Evkg9sLhaOV37SiVTZwnPvqG/V7OP7CIHhwq/YgLekYt
zl2hAkK+uysQB+g7+uhgvuOtuOhnw3MowwCjWLfkDO9wpnBJyNAHiqFwYcNXcq6S4OplpIEyJNdg
DgzdY46VvLThxz5KAjak/IxdKp8yYBnQEtKtTg6tYzfWS00jGlSymxxU6sRsCtMrknCcJ7qkupcM
UMdjjzkFzq1tjvqx59jj9mXaOqrHN1DAfNObptFUpFOMSggt4VaTu1CEreeYpR9Bcrj+bBb99RhK
1hM4Vn4GeYl9FwJenIkXv8AGywO/WzBEuwCIJSdQARNCjkM83FVmtzG8GmqLLq/X62LFRI1P9Ob6
nDwTmsniBRI6DbygAf0a7xsTTCgVWkWtQoFZbo2yI10uAUYPrS3VnElKoA19VJ82A0d2cqxBJaOr
5cwRNmBJJ3TWne4rhFLlTf97DqzQAoELxz3XjPf0m4wBkkgnby/N68yR+VRNq/b+WzR/3bw44ED7
/Kj4CEDFRpoMzv7LKGjtnCguHnVw6LCS8lFubJUjdU0rBfNxeHX37neOzIpXi4sUC+9ap2BqT5mU
kNlgYz/AesuhXBy50Acg9Qw6rH/lY5HgD6GrEck+3r+SK+2CoIv254FXBoMG0dHZFZNraXrtysZI
eYvGS1zozxWYkfScPEHOZ+jcJhUZl06mPw+Axco6vaO5geuvtVn6Pkfl44HUrKT9hgzqgrRj/t3Y
YRFWTyUspR7SV9Zetbcm8CNhhxtRaJMSfSN1CHaqh8qfFSXj2ngqcG6bKSwJ/S7K91drRUXNQUnQ
+cpIB1CpT9MgdZ82VAyVRjjJvx0EjdP+RJtRe4Qg2qoYrMeShWnGZCMJiF63Bv5wpmcAIZ/4voz7
7ZgCsao9woEoR8h5GeJsvRFnIv9AbAJr/8fnq51fZUNLgGsrAFsoNPyJtD+aiKiWqBD3OVWsp/G8
yUal1T8REZijBdez8o/W3tFAM+B/Xhe7PUPZABGaEz1WgcapITGaa7P7yJMvNzcZv+a7heVJG/Sz
rvJiVJOCKvP42pmgY1OuOXZA+DxaDoo9YxutXCQ3JyyCy5muF/jn3yIPGicDvz1yiR5pqLT6up0Y
7O86fCrNwGJzhifmuVz7EKyPWSyNVUguzRpDAxNleAM1hyJJ28dl3kSI4faDkqOEWH9xUF67+B9d
ze73LuM2z/dkV6zz8WqJOzRwMCiPkSrv6YHEqjDvJKUj67aQ2XS0q092rFeo3//W3F3qSIKpxYRg
wcmkht7HvVYg0RJp6HCWzEt0jXgpU/aYa9XUQ3t/Q15Ue7GosJBeYohI0BuGyri8ZsGSSlPukqfJ
ATZ45nzb9zQO4UFCCxp1rqoT8RatjBy1vNB0HaBDmFEzj/eTgTTvMTgK2W/73SuLPmWGzXdEF+Nt
mlPKCE1LtOl7NCpCOV+CHXjHMXqR9Iqq8/iYuMtwKT1Sydhr3Myej+ySf8CUlSeJPt4w8mF0j+iN
RQtRTukxuxKDiXsFmLFXzwKbwOwF47UxRGz6xsm/guna+FYkPX4lt441Bm3Cd8X9L99Lce6N7a1n
4/xDm/mhsjIXAq7r9BvSzpaWQEQAM6Pvj1cX1CgSjumVZt2CA0rYTEZ/GvA5YHCj6rneeC5+Hbvc
nK9wXS0dUIOYP+hx2R3/6/H/mChtncuBqCRPK+iLx4qvAhFXeeBZKUVQDepoDNkWZ/h0uyV/OrbX
ootWowSxC2a2OEsbIkL4ydToD45cTnmc4lfusFVPLg3ZQvLmFJUXOZtqFhpml0q3Fdy8z0w2aJaQ
BJqftagCc6zfe53zkrXOp7VgakibRjBL5UNBpgf69Oza+HcD+aVaaPToZIswwSgVYpZNSH7JTJrC
6SOOjDOsdG6/UDkk9FAP6lJSjpwALjPIOAcsO0tB3A8ht1DlPYcnvr/fc+miE/OOW4PbBl5s0pbE
UaD8YUT7bIx+EOu9ZxX4IYBf7n1JBnl2C/l3KBu4Qa55jq49YRtdC81HbMQVzMD09Wl2EzTMWcnF
SbszJQBjuCkn3rHXnLOys9lGEuyBUeW/TlSi+5XrMds6m+/VZ/3LZ21GQ7fvk9x1BjLn0ipbD0WT
2evdXf/FE/FuPDzCv8ZAY5qxJHkRckDmZwzxEpTAHbRkQ7cKpk9xgVhJPaWjO7AcCLzMyXfSjC3g
AB/HM0yfFkHcGQ1EHqWHqqHTbHHxOURPoIEugCeOW0wtfDV+2piTalqbCegjes5xNmIcGvI3yvjZ
5WaEMxhtbgrORxnEOHYsFMdVRB7iFt7cfgvrQJ32Vi9WvCCiAL+ykH4a7WHNMpMHPFk7iq6aaDla
NN7dfsva7yEYzoaJfyc406XVfts9iNlERLLHI5p2T+HnO777PnisTVBMKlun95w8zog+1d/o8mGe
wJVzqyPjGVF5uXai6cr3hHZJ7jRWvnD05VY1ebZf/sR4PPk1CXk1lQFiJpO0tf7Lj/ZK5g//qXiN
ZtB5tQ03L4axJOZIxcVsLeNIGJTcWrseJugN5HOosZ/0AXAne5CiWfny418pEVVMSD1g4HR5vOBa
1unrmmYH7+8B7FchadDK6proGWuu/aU1jSW5rm931zsogR3eHMU+Y/P86PZ3YIe0uOq7vmIoKWgq
wOolyzMkhHpn8g7kcFyXfO/t2Q5AK8KzAMcu6IM8X0qooItK9ZEyR67rxMyG+hbK9X8Lg9YVS2Xr
IEKzFDrDUT5r3vPZPVozWXFYfDM4ElyYvIpMsTcsaW9vcdkgaqPWUCFMv6sgL8mHHJn2769KK/Yy
VPGANXv2PcYn5ZX8JuPm9IXWqA5RuoKJTOBE/5i//7pFR3/S3Z5g2zEI3LEFc0eHZnZeMXwoGzmO
tEyGGq8zwM1es9ktkMCVCx8k64rwT92HJE6cjHj1lbOmDenAIOgNudyc+SoNLKxuTtiuh6VXL4No
D+C6NUiSvdqk4QSnURuwK009CXM7SZmh25HKwaR5OclVEYgDh14TTCgGrlWaSawW5zT4wwpFqnlA
fmBb95Ht2yYevfgsnZAxXciUNAd9tT4h5F7WLoYQp8oSjiPSD/585ta4FtOTB/zsmQlhfvY4mXBZ
9mCj4tO7l05mmQ0g/T2goF1foFOju+LvDnu2QYfQsR4X8nSaNO6OR3+Ndq8h1antQUZN+3kTXvOJ
8dHuzkHQBi9EirEAkeXmSCsBOqVsT4DpJOhIDGargw4aTKH8AVaPhvRSBKm1Y5YNLesXj73HE4rg
qBpO9rD/wA30vu9mBSCTIC+bqHWtBuX6deNLINtEhIXnunr1C6MuS1IYBPkRmArx8T1Cg8FGgyXY
0z59BJmDj9SIUZCCxFm0FmA/1+kCKlF8qnc+wHyr0O7cgvC4dHZzuIa76DSQ2k4hHR4KHtqs7STy
bVPfmxpMHh3FlfSHjKAO6pI3lZjWj+P5iKNj+v8jw2WamfpYqWaqUdQBhEr67gXZxihNpeeXZ96p
5TleISka/xeNpERAkrk7gS5bbVlYtjWroD69w/qF0gai4L+t9v5wH1xc5TPjppqFPGWPZc6penbd
qRGYt/SngCEJ+Ls0cULS8N1VDybMXEvjBRIAotQlBd89lMycaXunspYfx/aPEcKvjIEG9yy1yf63
4cFMn4mbV+bRzo3jRGNzzQ9juU47R5RPKlgQ0/ZC00CJzHr4szIJnWbZsWxK2ifEg30znfnq+WPp
WMuymBBl5kbOCMtuhiv3FPMYKkIcl4HuOD+/5U87SBW53VVcn1if8IAD3uWUWLsuCD4FRzZaYWn5
DMNt4Q2Onk2avPr1Ln2IzvqROD6GrhJ1yMPLGdl9K9JZ7nCJBblMKPCUrzHpsK4Ix7ic1DK/ifqL
5nvDjcD6+vKUOSgcVUK1b79gMAcT//6imO3OSL+thmw/5WOTZTuHO00yre/mYhu2dodh5xFmuRsI
BoiMwTV5JKSTHtYPbBhHKl0toXEYKOKyI54+zCmGbwqST+d3S7JibLMnpnCPA2i2DdVT4y0nxh8V
amVJtZU64Ld8dvRPrqhea0Np65yz+NecfOtF70A75sHCt9E/LOtp3Mr2f1RxPLumgB3EG7C8bfA/
cvVOH4FWs7Mu9HvYibvBAHczgV0T4I4lS6XphXtuUhrCzJyybiHy2CCBW0maIpXAfpB118Az73oV
uigq0FiMasiM7ml+9FpqX9S35Um5qqe7Lo5nMXr74W+0GshMy/0luP8T4gLYP8geZGkHkD/Q1xZk
bhO1xzVFzm0RPiCOc5rgatA+eBAKu13FaTFWez7xaKrx9EMxNmQ8bAvKF/cbHZGwkneVqjt/aKHu
k8ZzJ+b6IHuo/7tfl3Q7WtGL5ejvOts0x/7zZYlQD+toeui6FTGFMMe1x4BPDj/A/UTTDFGXjLrS
203jeNkw0TTOe1W6gsJD+iuVz9uQIOK3uVlJumQ+l7X1Bu0Tf+4Cm8p7reVlOLsoad3FZf9kkv1x
3MmE0M2Hd43i5VJWmeXa4RBGWLZxVEzC6DkhdmRqrLWm/ghgIQmpSwRPoKYRRIXVn8Zs1R4tPQKW
ec17WnrbzhIOVKoinhvjcoEkWooSRmBclIFSMJ5yP+yaohL8c5e2bEfQDwDHp4vKLd04SWFxQqbl
q03+/xRejbWlmKBNVotpCZJ2oL3yDhRg0vJAMJhh45t2xV8mjl8e1ebdfyGaxgndwMQ1rlv7WVLv
IJBk9UbrNN6aPLFgadY1c6qlrnT0K1uLNBiQwaYzCOsfT0ZG6aAiPtBj8SY7wNcoom+g5ZorROhW
62dDrA3IgrTNPUVo9IV9Qb7sAbQHJUuv03Tae2yThz1it/uAoFr73cYtmeFnXpZizW1dsOg41YBN
hBtXOupP8B0gNdtiD3uvLc+wq8+loegNjhQQoGq2ZUyCtO+yIqmpOrhBOKQslEzzuhADaPRmG1ua
50kxpgI1UJre+yq2spiLbmhvAZ71KIpyrPBLt6zuzBsgJ4eH+a+uSZypAiLD2dHnqwNSg0BZI6zJ
SY/3qRaxQTDqziWr1fL/qNkBxNjb7FNa+rniEnaRNyN0Cmj4E4hQThEOYahLB93oYVn27sn/i7zA
FbGZ0NwBzIg9MFQgZZGMoC6Ym2MUfN40eWiSb7Rj9/2uG9dBxBYnz8xqanUB4RqRePx8cdDIU1mm
6eRFtS5WS+bs/Gk1qFHIMIncRx+AjZWB+b10RlA6t9s8x3APKmtY6fkW3D71SEvh2CrQxbovhrbv
Gc5uOpDEZtENxh07Fby2wzzmlt03thzwpmvHj1woTGU8bJbVmjqRzy95tVh256TyD8n9RTd5OWso
KYzvO/h2K3FJtPaMTpDdsth1/+uCJ/mHnFrlOa1xcBWyJclOIxcOCG4sRPG31KbLgeDG6Sn6iOZJ
x4Zu0so69+aFLeCw6lFzXwKJjG46NoEs7Xu0AB3yzS8KB8hwIqW/ZqaCCg7K4J8lGDqmdsi70T6j
z0wINFvjv+GGmD7MJb3Rb19HoJB63ShvORKaOOue0rZZ/tm/FOOLsJn4CMOWbQa4ZPLoUTqUSUvu
KLJBZM1zhNdAcnkuZKQWQCqahlZcaFWdtv1pDVGZxmiNYpmXczNJiy6eLE6Y5OpYzxeVtlH0ZrhR
OZMbroyPRR+VXmDO9MN0PYZqZ2BNFJekioG9xAgXg94h2P4yonDMv+S6ru24tz6uEx0olbCtCg90
/qvNYAj4IOKOsiD9mZdxn+/0tBO9ZJeg/YkIIVMSneVQHYLmZSxzffH9TLYxLCB7U6VtzK/Yy5VM
VzIssHD3nH6MEcvJTgr2U2nXfHRQlNzGvS7Zsscno3TNcWtsmhlnh64JrZm3S0dNOsq3nieE9f6W
1ECxmoNWA4vTdvWkhdUnLlqrCBOXVXjp0sodtHfN+yHv/RlrQB/Acq1V7KcqKBXFEYbkVKs6W638
Vix0eRMFtKki99nIZJahGdBZrRleekrLFStuSQ7oC/w/tKeTRpdYpc5CYZnTNNR10FINmHIw1u9U
KWff4fxiQlfb64uxOuB+9N0vN/pGuT8INlBu59fuIOWnK8xOZg0GX0vaHK4h8FlOIEOVZM4TiQ03
PGIuq7Pu85AIrVCU1jQXmV1+UK3X+Hkx0O7CGQ5tX4TyleOiUjWL87y/KEkt1NzPQ5CRFnxs/QcC
C3PxVwAQAfn4EJQ9smoVdPmVWJ2qk3bTeEUwCSh4R/xt/MP0wtlL9AW2SbbwiI0TJdtGKD3KXN4y
NPGTwGSIU1/+1M4ai4phtczIbRAwrx7HahRw2FgKbZpZqrzGH9sIMvx00ztESZm25r9TGm1M56Rq
IAdK+mBd5wxdkQWUgc4Ide3inU5l5H5jUhiS7UDMUoVEaMUwzqExCsA4idM7K6uIR9oB4sySe7/A
Mr0DEmsonOdbYI0DoeMVpo5/ODZI/CXpv8dYu/5zNQxwsMtmJbWEsg/huJEQB6C7YBVlkfsoQY/V
y9kYKampjRpl3AZ+05V48tgebQtWj05Zhxed98OEm6m6LyQ/jEfk6MM93DiJ83zTeQPW5NqySaQr
weVDU6bNNSh2rH4ItHkdworBEwNUlJu7bc9zLq1Ip4qy7lTQV2myEa2eLu5kKU8RqfW27KAbSVdb
kI2Wrg8vEIU3SPbThvMEFRifw6L+okjzrlN4buO7XWd5SvUuFlyAwfnMjbc3kBNn8o8n4ivALZoK
sbyvBS+BJkN8DnKU+EOjDmFnIQp7hMw8Ggl1wNII6GgHVNn9Ls9kRSJRcBlE9pX42wPWWYF/yKut
4MOGBT7Mp3RiFeMwkhiMWiU1v53hI+rdwKNICGabK2o16ens9FMSi/G08XS0CI+ViO2UakqkKxh7
NjvUwRe3qP/+0FlcrGurpMvGMFWtmLjQJFWIqoElLXakT9aiDuLd5wZ5JemK0A6JW9XZD2Ha5dUz
6lmRlZREdLf+JNLvqQZK/2MIZbjFoiwcvv2BVVOzr3AIpvpXM1i6jlD9ansK4s91g6Bt2E9nkdh5
ykaefojUgm8p58K27doaeX24AialjBZ7G3lkHOtaYDiG3leMX9uTcIwp+vY1uhbihqegapDp5YuP
haeliAQ2UXPZ2NmEW0rLSVh+wUZCDDxg2Jr4XI922MgMkuBwnYIfRjq09lbfjAZpXn+j7TapOPmN
P1slrDINTGEzyye+a13HlQmUZ02dqRwOvqyVDY00LCbCm6ZZrYAfYZLz7aL9M6kua7IORRGkvru0
z9yF1FgylkDNHILVWdIx2T3SF54FizxbZOiCElwgrwReSadRb1o+dMDTllDm+SXfVBC4rPuK1TJn
eMDqBRm1iR9v9A/9kRGYRc7zzKu/jLaSbGMEE8T4SSUKnDBX/8BRozzWOdSNAPvfnNO9yzsZk6a1
phyJO5oTM0O1JBMXLWp8U6Mvx3hcymPYj408SU2j1OsQzQU3mcLJ/a3+NTXMfFyYrVRQdUzZ54Hm
rb2D8Lsff33Dk3/4DfT6bcLEplCG9Jra55a+efC5PwCDqPCMfqacCnektGIAMDvKW4bWr8u080OB
aCU01MTaKMgFiqsTKYaHFYuCuiJNwuQmCH82vnt0u55LstPVCo8HvoE3pjz3nSd+chJyQpOfwVhA
bKPYQhwbmdpbyEbUNhmTdsxsC4dNKG8JqvVJ+z6NmZ1ZgOGEQbZB/Vnck3SrnYNT8+OFNJ/hYtjT
hnr3xoUPth6D79Zcg3wo0DvVWeRn5h3hjpeh90mkLjF9YgA+zAgDjs8NSmv42w3GnQ3Q6jpc1J+k
z1zdsbMhu5B23Ukp9jhK1R9XXZC/rs44vwks/kfAQI4WXwP9hlEig5te9wPrPbb96DNYxrlWQkpR
sAbAj87h8zFpHbyI+FyFPeiI0wB+mJCrysZx1+g2G4gGMFUTtmDHlrTeJHYm6/Z9K4Cqd1/U7bmQ
zyqaH4P8rYN6oHofgSqpOvwzzSRWZSPOnsFEI16a/0PoqNs/y+Y9aGxqMWk7qaNjVgUEqTu0Bvok
rsdSU2r0/9KEYrZr0nENdy05yvjHk6NNgdFyDS0ZwOHZ9o+ZYNb7inJnwmKE98MwYr6qeFxJ1m5l
MDu0KGpo8a7IAKHIN0Cku5ZZfDRWiRABQ7+yg8zIg1+rD3ZxD0tB7r0nAuxpjeT0jedV3A+4QZi7
9DTzKLQkKyn+DQwyhinobxqx0/mLQhu+Mn2LVkirjJ4IjUAegSa4FW3x92c8gxA72gLXG5nyAoG9
+AATmJhfDHS8XlaAnz4tXsDF1ZUQvoLA/tuV/Dp4KJb3v33/KtbCrouXo6SUbpb3JdIAQelXecPD
MDIGGu7OiK7jZ/0N4RW/q4t+YgPLILZi2IMhHM9tniGFaJTHUAqjeQ7r2/j7rJQqjdLAexWXjhAI
fLAPa5D/Bvnl5Phvz9Kp0yHPgsEYQNxOAG1NkDqhDjvJuesg3PLeix+gqJ6K13CaC75gYbnBfIMD
NEwi/5bpQ9tbMfmZ3eJ0zRpSEJHSxCutNhB70fcMgfwxuZGFlqtlty2GHM1b/LcGVuZai7CCQQut
rZ4zgQFbiIhy0iUmJ4qiebleLxGuzKAO7gm2TKEDf4OmqIPKutaEoVRWS/HvJSSQNq7BARb4bBS3
+8Ah5irHVTXbp6Yy2g/oSd7ybJMGIEvLDQKiTADyr/015extdxBd8oVUk+JQDQAXqgrFl4/TgZXt
GkaHXEWMljphtaUoG1xY/M2Rs6m2eaKzq1yxwYoam7/+kKaQ/3bfsCNjU7gGV8CYxEnsTqSPagHA
pTEw2zRS6ll2i/BJwpvktCIkYIM1OZOK1FX/VODsRIwDJKpZsjVMn93c01jaKsWIUxEUcEv/zhfX
lFmzSPepxJUTBRq1TPJJJvNd9xiRZhBfRYvtUz++iC72urcbRlTPlwwJaXHOgv2VpPzD3yDnLvGp
m+9p5uvQ0T/MiQeXeKpNmohKQLBQesd25wsbO2zYUIBBBEiIlfcoWcE6YqhtBmc/Km7dScOlVy28
QxK9xQiduRvEbmi4GXSYZKY3B5+LzojxdRLuCEZFltxb4adc6qnW0liCUeKqkmjXsedVBL4CYvwF
M22V3MzCyr3OCceKspGzI3qmK3jsKggXm6AqIgDfnWlQUoCifCeebavm9HCmHGp0CUszOYa4uqub
f1kPAHfE9XkWaVvrfrpfRQ8mqPZDeR/ixhN2jA2JnMyZ2TDCe4KEOypUIPaVQydAiHVuaY117NtN
1Z1mKAgP+9t8xL72BwIDVN0DTdZySgrbyjmKrHl8lxcCjwkdE7yS+NHj4TK3VXKWFUUZkgJfI80X
0w39oHSXmiifRIZ5kI2YyvYGDYJUMh+GlGc09Ty9KvYwSTVUkTCs3m7zufggAvD9qIOk6eWjBhtP
+mY0/X0Cu4fcTZAgnpA284H3hJOCPgWeKXCUsGkW8te10k941x9zQzexMuhtz81zWmXvClkJivYg
7sy9KobGhW1FcLc+XL0BRq8K9KIQPcaE3c8zBGROScrQtAwAVRXZHZxBPnj76Sj/+CuDmZwRPFyk
q7ATnDyP9guvIKZENlywDJ2Pz4rbezG/TDo1XUfYZP6KEQ1ZKB6cbo/RoijxiiShH4NJHrhiyJos
JOn5hRrQ0Zcw7FKt8gOag1aLQnzwlOaTNJ6k+TkNTns/nm0xoTIe6mS1EKMvx57GmvanXaEJz8fE
QeqokG2rSfu9UzTIFtVt50F+uVIN8YK78eEjRUFKxLMB9xjnm7lweYvOCjzcV7tWPBZP4GqRHTZV
9dZz0QbrE1mjjjNHcxipTe0bD+TSG5q3RFadrotTQbDISK0RYqsNqgE+XXI3TngJVsMpoOMJqWxj
vxQp+abRqJ1c3P9FeTkyA6w5HX589LA0UD9lQSvmdF7prCuwU8q6fjAjBXUbRCKH/NRdLxiqY6Qj
A7LgrzGr6or9WfJEUDwaof2X3SYuZIGrfH5uKTywa45e4nN/dJMrCgnzozKVXcSN/FA8zhWWO1P8
F9VkGyFFU/iSoJ0x5g4E/ITDkg0Z9//Tsi0pd511KV0C+U6MnQh4c9HA63rs9su5PDBesYR/kdSO
WkATgaUQZthWRKNxisZw+iu5VNSZWk1cWgiiIdgPRRyLuOv4mrKjwitRCJRL/5UuP/eY0+PiJyaQ
RfE9B3CpLH40qF2qNmNb9eqpJbPARNg2RrFvw8Ri1G1JxEP5DCzLMjXcTz7HMW+LjyFoURkw0pNs
PxMUyLKqg24mjebfTeNwndME+KwwgbTe3ZctpxR9K0rWpXKsJpea7wLZZxITq2ED8pMGNuG7nP2g
DvJ9pbkabEZVUeOMspkaz5V8BQH1pFJf/+MPeIvAZbnAGqhQ5mWsdPI803ywfcQGENEAApKXwB4/
tb7EwkM3NVrZbbNUJA75A8wD6Xgn70InP3id99vgPN6RORLVjUHV7abVrxDDotIET5yvNqygmcdE
HCUQ1n6Ab8OBJ/q1qRup2YhH+5jKP3CjVPNuRNosQaX9kw0l430HiansAD9XA6/TF0CeNvuxVq2o
LXtx94naM2Q03atxr4VdKY6JsdsrfErNdeTBuYKZASpa9ISveML+5ZjYYYqJUQdnG3LUMpi+S/RF
0GYzHXBRzXmifWG9N3OZp+84dWceTkRXN63POMWx0v1TYf6/JDxCnlMNjel/oJ/Keaa4WcAD7fXA
bD5zUo/4BLOJJH3nTh1RsuIBVKAIMkXyn37NVPRZxRvkbT+uBwT7EXxmdGlm5tB/PrZuaZF2Fcdx
QntQC0esMAuknCxCYhkX8/DkOzQAzV3wscVDxIAfMctDfx1g7cwJ1u0k8JPkJy3Vr0snjf6vDviq
I3m991Yh475dZ/nTBgTOMwCsetsDzfkpPLaOJjlxYqG5C1jeHzRe5WX3w4KYDZGHcCo9F5TuhBlA
WrQhBSQ8jssVUWPzXgxQZTH6Qlnu0AHpTUbf8sJhPteNofcHIr8zLdYrh/zhSx2EMH1OdRLa1+Ma
dXl0kZqDTuEq6svtNYw6/emdLgDxgzaUa0aS1gs87PdWskHEdE+rnQH+Tg/7cOIAAxSd0gsNG3GG
nILY2HYAIVbr1K/fABvb/iBfJ0cPd0rVWh81N8MCgPe/phy1B/xoC8Hb7v9zsTcadxLvhwzqQfDT
npFt9TPDozXO/G2Xr+o2cfCSBAbj3Ks9f13oQ+TyRixRNlQQ1ke7CwDwOH80G7El7IF3NXOBPZ8T
thMNj0rvd8sMLVrH6cHTHNDh5Ct6i2UNcRu8yymklz80uN72YpTV4mRxboVRMBKLCzVKgQc9eKAR
Qxw8gMuGMgddmZ3zfBvIEOi340177rfFgLpCX1V3eG9l8Nf9RvdCQ9+n5LM/B3vhxE9aYiYKe8jJ
aelOCraGDTgcRig/4XFl1jyng8KWHxZwSPFbPR+/1uVHoRurEKfZQIhAUSR3ujCg3WXPd2aiaAJc
dwbId4ARrURnQZtZtvbFoj8MpzL7I5OkJN45dvvGOE2V3q0nmb3zrNNRY7ncQTmF1CEdgzomoK8n
KQLOiGEvUZqvrL/Z41hpxfAeujTudgRHdZQO0u4W76nh7DaBQdQZsZOpU75faZ+hphfzSGU5Harm
KJJFEL9xusH0+p4nnv8CYAlgFlbAs2nEEFBpVqp50cif70Y1u4qa4zMvwOoGD7zg+p54Zc3pQa2H
K1lRLF5RpnWsEdtUQwQKABL41jgiK58vDSFaqzkXW7oKyZiemIEp99xxb7Hx56hN+MWRVl90YUKr
PFw0Kz4Cmicgcb05EiLamuzrhVRvQx+9ADNxcVQuuDydHSx1UTFGjLuvz6VDea7fKqlAkuYgbfPK
DU915UkVfCjoWfNWH4nyODnb9CtUJUxuFc5PPZy334SNZCBg1YrT5D2iFSU89B757AO/NCFsXUfg
eCqPWvsUDJNb0RBnIODppOBfbDEJBTIUheTcBJlZq49/6CgVjRdAT4w5Eh9NUOHRBX7WVch15e3N
l9gcnbKCZeMg3o4RRrmYLpwaO7/Osvno920+hD9tCw16uyJkfVerLu6C3l7/vOYPVXoBLh2bjN6T
NIeaUR7jUHrUfgBXo7lSfnD/FcJGzbCYXKHz8jigp+EhD3+iqKvO1bwSTre5YvZq699AdB448gRr
RSmcVeakLsVZm4ju0zGH+8o1czM3Bhg4I9pAD6DhnrZBXmIyBC64WlPp09N9lhSlyDaA8AGEIlqd
Sq9GGMjqZzfaY+9/JLP3IoXl3WOVMexkAM6qMbl+L3SU6fF+aMAbB42HqQPTJs9BVCgoUgyq6aIt
hClyKN4fEdrB4hdWUHancKvCrMHaOto5V7KyA35moS0bMxEVlKETwPLUs/TGx0Ybl90+OSWDF7nz
p0gu3JT27YuRwgtUPYIcAC0+OmjJ2ugApkbo9sQ66BxKtcl9qWEUewf7b0ki66tiPBxwcTaIzKOG
Sbcxx2/ohTtdG1FCh4PdR32LY9wAW1yl+A8p/XIAH+MxQWMNZxdjzbOXyE3DFE5PrhleYeg1LoT3
XFcadTK0bgUEHNH63pJYr5U8RuvEk/qPUfW1+hfTl6mcuaglKUcVN8VU/BeXpTOK/f02CiUx2hhy
I2vnuYoHiwk8BPJzHqRzC7Yj0QUXkQt+a777Ra2gAtMabZs88MBjPlatgNia3Gk4Xo1MEjozO6XN
5YIwgzkrurj2op7x0cMv3A5ACwZSg98KWvGiboNRN+73L4cjPVVAXawPUkHyS0vy2j7UioBDm0G+
uiZo1p1fma3XIgFu1iRMPVZcWse82mpF4+xRLZ87/y2j7N3smC8v1HvCh6n4I3g7bxlKEo0QoqgX
9MMhQdueXzuSESlv0zysUmn1Aq4CWIfqa4DNRZXHOosAWhYm3Oo85WJo81w7ykmd0NulWHNsHT/G
4e5dwkT93UBjC4j3CdJSnGNaHlHZCm4ViceKlJGI5RqqsitG4bKnr/8V4cWTBwMViAk4ZgABNmRz
BB67HRATjBXnDlSwIFO9ssRUer3NFaoL/XwTzL2pNhHf0efHmhKBiIIbn2od/EWMVjpVIE6Jma1V
O5xfTRYru7dMrPxFtqPF3jQXZ+qUWycsXQJLfTe/qy+tJujhhVS7eB8Ggz0ST86dcoUq9Dhbd0WR
B6LQhoH9B58KkaDt8D45VEY7lXR038JUk9n2KSZdzVlEXgH7UKF5YRzBDKQn6pQr0S1DN6loKPl7
GoG0rdxJ0xVjckaOuD+TC57pGCSJocqKsdCtD4eGaSNHHvU3ifhnQfi29jmujvEmfsKJMOz09kEK
XqB4id/CfCu+TG7wPjRPjVfqdu75FtW+VtMqS9MEC4t4vzwVrUT4HFmCuE4jRhLf76RJBOGE+t2g
EPqb+8w7n+4JQPkt35G5GlAZcmnpQOl2MqgMkOLZ1yueQ//MJzdOZsCaQgEcOTtLlsGeP8VODfKu
fxlL79DO/OvrDQHH4YPFyJ060OXhKTKV/XmiHVYiMzyyqLY6BTCzhvrN9gQAPNuvETTHNa1Oi39h
tLRqumKmdHfAWLVo2Qsfa57MMkjr5g1uscdoxik3Lwi6ZnDqsRakosTOzQTeHK+qWqktcD0LZexI
S+mF85b1jD8Gsxiy4G04HaIfUQ0KIWCIhPE2ZysEXULE5HutvVUtmRoYCS2uGjDm2HuV4jNb1hQk
AV1IzG4/hRNsmOwqh/VbOR+rxInpcRA7rSovH2rEQzgob+AE6wpzTsJYoXpmEgY9LOS5tEhfcgZV
1A5l1dnXBjCQlA9WYyjaavdrZWxkKHOIhpDcoMB7FpmAHCqoSzhwLWu/vZWy3mUcKLL2cn2yszeE
lf+kq/WqYMWOLntcJt6LWDQ4neQ1+Y1qQR8OuDQ7091IYT1S+QYRIJ6bI3xIW9B2eD+oxLEtiayz
hOmIf1ctDUP//LHB4MW0oMazX4qFTxaBX8t0zbHeu5K9W+iTfUM8zT030raAUw+mwxGmp3bQ4mnY
bfNcHBbI4gUuk5BzsOJZ/yVBrVwr4UgQKbonwY2qL89xNUD6pyCSFzwJKYm0TOuWUvBokZ/1U1/b
tIbMcguNp8f/f2nrWbyHUKJVe6kc5uC91lNz2wXOERZAbm+EjPVQE05ZzdGteOpfDjN4ofVdax6c
lo2fqXFU+F5YJqvyJ55d/l43BU3sV4oHadWtU8HOiuhChiEux1AVasRrse0RxKm9nSpZuMCJ7vqh
/T7pJ0Cic889Ld+Yua9gif9jOUE0w5FjTqqalmho9N1gbyu29ZKpSO1NQ/G2gg+UJX0JW9wlrM4N
ceSaolpbbC1r2jucLYY6fQ3Vk0sK5ICrS7ir2NBBRsEazi1IyFL4e5reHHTANo6l8k2X3Vzbr4+4
EAnD8Iavyd4KGMuU89uwPazecuGXv2hzpiW0AX+NZFUaKoz55q9q5gwllItHUAGt/7xy9D/DLcLi
yOp7/INAeS0xzkEqgLns4SHFqg9MlpKeCGoRdKkUw+EdVIK8JpasAaTFbJt07pbEuW0RwiUqDNlL
aDKPP1xNTlt4e7/M7KxS9s/TxySgWhCzz5bFDiHT1izM0r5Rj0Gn4rBGL3oREoNUoRMGHbL87Ba4
tL5e7ycyDMXm1LUgmAESSOmZf499UJmgI2F2aN7UTicRCOjZkR/VHI+mKKRl99GkZVnYIZ4Bw/AR
ayakY4KBL0jMTWDeR2RF3oOwfIpn3Hxq09k8xZqc6LCCANbuJn7a3ZLYjYQvOuo7uuj4OkvdPTJP
aMUCLKLVwL+RWypjut033CcoXr74ROOBl2IHN4jz77aedTrVqx75uXzW6I42MJdvjv17h5KOujum
56AV9eevGios4y9xq0f2rG5KEeInePbdraCB9itqyYdUQflppp/JzTbKOGEcrAWfHO2cvqwJH6yT
is/H/N+Ztx1xLZ6MhlZRI2f9FGQe8TNnxGmGOT+Eg9Er3KyjmcztCTt+KwmUhD6w1Bhu/qXHV6DM
zNY/k1IBh5MRQg64R4B2bqj81EJSxTHiSjKo4FVKKOC0lExjV4oz/+No9YXZtn/KkT8g0y8LfXwV
n0XGPdZ3Nx+6sSTRj+y9Y21QDgG/QRx+0QILHUCcquiDAlgBDMrGjw/3lB7qhR6Ac33hBMDg5jAx
yFXqJ/FAYJ+RPUAbsW5g2uH4xq9i1ZeT5lJHAelJs07phjSatwPe8VlHauKRRS6bW3E4KPqiJCqz
NlkTyyJ0MjjBZz8KGvQW1RGYyIcwD5AQ86tOxSj/ZB1vqm+VldbwAseT7JS7Kz/GVPrmEfynjuCg
aUUMMi9XwyKHm+VBG6xp2uvOBYCY4IsCRIpps14Kmjpy+YkYw7LpGMU6h//nGdiFRj9SlhpEHP0K
NulcoF6uhXsN00y5Yw9gvjO4DzaIg7UTApjoliS9eDROpVxzh9gl064zsw4QVZ/20QJGxZZESqQr
lynTf/8rFUg/B4gw0iDoYwR6a3HR3jLSkNCdPu93wjYhQlYZ2fOI9zSMU5WqukJ+9yA9tTa717Jh
GR07QG9r9e/OwzQCnju91SqNiwViEYY5XCcyWnIxXWlzfYWx73ebb7V73d3bltRWcT3zfmisjDCQ
Z+dBLTSzN2uRuYdCsvxK4G4Uf9ltAhQJzH5rRzq51PyX0xTAm5F83b9LlrY/N/Jf+BOkdXns0YCz
tjNTCv9YNAAWbGnU8XmkJRVHOszVI49ylb1wYRABH0sdOSvJ6twg4ixj3cCHk5W2tYybQIhHb09j
uXkQaBpqfnrpw1EH1V9GNc/Jp/LAI1/RVz4etVtRTQxGKNPSOO0oVZbFaQMYMyTF1tN7DYqC8jld
4LwrXJUa0jF7NwggRn/nWQgUpzecXySmff0bZwPwXLIyvWdjpCc4ZSy++Zc+1XPU0EtVqK1dO2Fo
GPcjj4brqqc1kfcwxIr9G4sUyoZjByjiJmESNKRFQsEQnUg09mb3UkIwfmK6J9oWuVqwUrHIBPaf
W9GDrJiLLbmFiZuvullDqIst+ybpJPzwGeVmmeFKkmcvCV4TFo/yeHVUp0XtU+GAcIFz/82zpC7z
z4Il/XQcluikB+LdLqLm1Tdc2QRPcsCPSXJxt/Ql7omknKi7IfdbAg9F+C8QqvT/w7NpwnfuOTmE
LG8FNJ5nRX9b6JMaFlBEFj3s9LiwQwr/Bix9WPFIwtmzmcsmjn3FuXq3oRq0kze7PPpuqCp/7VWZ
mr+OuzrINAVQumQirjS8FF09dJgNvex5+WVsQ8diVtonISHa+7a3tM/U4V2foELF4CujUh9fkOhC
0X0k9/7l7SdE8Q2yf4MWPP7EpqP1i7HSDifu6zYIukoBpylbFZ5F+T9CmEWZcpYeRMcT0lcvWZDu
So7UcfENZST/VBIaL63jefslwz+U6/2c5338qKgj2FDX2YF1nnbaFhBYXtNaeLisMo4SmHcDBWnB
83LRLVtZWEW8AKjOXuEZbdri7jznWRfO1jektx1zvVlYyMYX2A3bnWwTQBzSHrFgukkmPJl2jOc0
WmwW6VsctqT2em3fuHau92S/Euwi3PdtIxk9S2OAQA16fsOP5tJ3kLRwdNK/IVPJ9Oa1da+HUs/1
9YXzaK+3jAPO0GFKf14CzohyaHKBsruhXXjiMTTWonQcqnOPwG/4ZcObpT5jifuPCPtMImNXz0qR
F+1AlYAIz7vInFkHrW/L92a8xSCEx0RBKC4tT0d9uamTvt8STX1wZgQ+hWqUb8QCQ42TQggXcsPs
tZJjfRmwqDIXSCorwCFKTSYlySJOPYPndPifIzKmUIO4yrQB25Id75a2IlCYSztkW9RaojZxRDkg
iZiyqhODcZ7z84owOtti0/KP1IFV9n0DihHHBQoaA14DH7TpoU0LvI9i2f8coT7vEQUrZnWAxvKW
VSAfMWTRLCJIOV5M8QJuM4+8k34JnnsJdyZCVkwe3XpmDGlyjBaZXTc028qZysTny4QBJKF7M1cv
3YaX4R8LObNAdaNOZOCqif//IgqHqHMVPoqz2sC/WxmHLc0EjNcHi9Mn7BKWrOPRBmibZOuMEVXa
cYIWGbA2d9fFdm3FPSaxnFE+bXw54z0UNgQoPIq1BOlvfkZGpNQNbbpdTOY+vbg+WZuToEIX0Zsg
JGWuDeI5oaCQmuHfAHirMvfK99+EdEGg6pdKv3QTQJdlz4nQK32fOFQhCHv9JRWJEPLQHsLP90/Q
xV8RymBJNKy5clRwOt4umeXWRQEn0iElULxH/4ItBcbsc4ZBSqlWjUY1wtIpzG8cImN3dQyHOqQ/
uWCXGoTn4OAE4Ml44qCCbWq49/86XDMjgv13mnUs9AIJK9DJCRSbEukB0ulTnO/b/6oQOV2TTxVV
v961VmYOTqD3YrUiJ6lOINs4Jb++7hNpY31b6u1fcuc9omRPDumj4UIFPMmsTxn7HMWQ33yvVGw/
rQGzmPnyAnz3aqRS5Je8iZtApf/kdEnO69/mRLCrNhHd+9AgMhR3bkVcJatN/IV7coteH1TF3EKk
cR9okkehcpCU7ELx20k6ICFa7CbEZlf+9y3N6DHgT2NJd8gCO8oaXYK25Gam2XuT202N7hB5pqhS
+jiuXDt0Q+PGvqiNNt+adVhgUQB5FHeM93DaiYtTSYuWthAplCasi02ToMr7fdtZTg99RAxh+wWf
qT8XNDh+G9oN54cPr9NGOtlmy8ZUIDoWkVTFrpaREKM9HEVabw11TDHPv+ZQh0E2l7/QNfOj5UwZ
0ZYsbXiYkfOuGsH36cFqQqhR+p+k144bonkLbAZ7oEGWDh7OyZMNQZUmEZmtejcBO6NNDYFpOK/B
Fow7QmYt5UcfE+XaJMpjYDG6xigxPl99fI72TJN+4+M1CIjejDQe62UnQwLIGjXsYijw7KTy3Ngz
HMkuYVItu/oa5nx9pvKbCiK9L4CRprPHFh/YBkpiFZEp+LnYbav1fuOHpO2QDSwHYdsRSfp2l6pX
iUZG5d4MLTf4tIKQem37m0Iz827bZ+P67UU0xYEKdRz2CXdh6KhavmuSDBFew9w+zBuvf2toIw0j
J4WSmYFqIky5ZWsCZGnUaDIQ6MBZ7K5A+7DjE1hUL6UMspe60rIrQlTXyDngVY/2HrNreVXHw1rK
I4UbKXBgx1UZB9Fzq6WKtKdd6RvN7xER0Mn4XgURzXuvfNMXqErU56CiF6KP//mLW4lCx5JZW9AE
2922BcRu5uhfwK3yzhTPncKzQVH15QraeXOpatEfZVnMlWzoJOqZbOiLKLuWlM5XR/lScxzWiN7n
tIT0vSMKLlrNcqq9PtqDUlBC3ydFT+Br3EnGd3SzgrS4mV8ZuN16kU/lLAxAR93YVHwpnBZG216M
57xSo72KB6Xy6DpOq8j8/107ElXMIqjcgEyC2GleHhrq4BYa8XhKnLR+dKDmrVZTFYbcFSL5vXxE
fBDg+zK7O7mv4RQefipSE1G03f2iI1/WaIHI+sZdYJxQ9MEqSjO6t/PqrV0LUqjIhLkF4+hpfQIg
kam6/h3UZA7l7WdOOmiqLsfhme664tlKso0Ho7tOCEudWpqzl7bV/t+bQMMUINMMdICKOyspcMvj
YayM7cPjYbFYXejYSDSq77jNv4o7dfbYhRE1+6gcjFsscZhmEjhyuXgZIrqLktotaFiy6/R9i792
oU/hiSe/TIqIf/PhHlZglNwYMJFmwPGaZIu6GgmaoZ5mfdZO4oYG/fxnd45q4c4m5Y7ytoPeqT+v
c0v3cCVX1DEqk/1b4ZdErl1EF/okr2v24DFSHLSBSPV/4NXOOPgSg+qj3woJSbRCIOzRzt3ZZnA3
1NKzXJtDSyXwDRdxzyN50/0RcDGUClJbxAZ/7w6EzE0hHj7Z1E5W/xzjLl9e1jKqPrR7bmqjzG7/
YsKpTj54qvAIwcNAP+1zh8qn7AvYWV2ZSnomKS7MvencVVveFC+meiBlW5a42exRJBi1YHl0I1Sv
7tHv/A8DglR/39qHzo/r3XvRcT2FkNvHMbMbcJrPEGhyDO1kHyY3ZnmMqiJxDRRzw89/+YpV8FeQ
IoFsWf8M45b48GQVVhQeJkYzKuYFSSao9pcQByMi9StbJhxELD3zAVjFbxsyENvu32R+2gIrUVSZ
f/U9IQZ34T1UuPHxAI33FSQdL/Lyf3ylbE58u6a8+hDfiqSgT/4hnEBdqPzB51AZNmiullaKu7Wk
jF3fvD/kWMX/H9eSuCfttpCTb1isSlWTaRqZSx/MiLIgY3CoeC9kp36UTfv1wpiCQo2pw2OkxGuB
v3TcoHbvk0sZBzS4zykJMUbtP31cOzXsJOzirzpL51DKkLXXRz1wNODarjIxnfyobex+6AvDezL2
CZVbpp0W+ltaN0ZR0ORKePeMG0ZAPSbneMCcR34reLeowUjHrbJGlhrmU67OWfqOyU7tFPNJz2fY
skHWtkx2ArDGZVv40EkpeL1cVV60Nee85kC04XJ1Ts/OD7icAL/0S7VFcSNYZ3+JOWPO9Wu2Shta
Lgx6tirEXD3mPLhZMHgQmxc2OSsy7mUDYrSX+fGre8QoU3jc03B+8DCP1eHBjVZpgaOg5obZYG9H
1VfCLggGKN+PpK5mJPaud/tEVEblSCrhm20W2TIrKQZxKY5gi0v4KxNm0BWrTgvK2ZLDgWq/EOz8
22Baf2aY1ryPAJjRXPjIBFMTqekonwQxO0UD3Cd/7rJWfUy1Quy6pz3r+3MPiZ823nGi0wZH9C7i
AUtVGMZ95DERw6J8rTXHm48bUUphNhlm0tbrhzz8dpmwGQBrYj8vkf8IZBpneKWr/JvMZ2QmzCWW
AUsUahqh3rMnTSQ9oZ4lHvdtFJ0KEwgJc+RC23AK9cB4ZeYdOC32fZLE1r3vT0PdwpS1PSBIvBjX
RuE7TImlSWgBGakMOuCy5J/7s0OxJvUf3B6cqUFKwPtXB9CUvL3DsA1cuYjDQg7uItYJssnlhFgP
UonTRE1l0DV23ISdIeC6hnpnNvBg1eU0+zEZ4DXHmfLH2WlfSMGJCjHHoCId+RgflrsN6yC3skas
+ugePOcGwfbELbiuDL9I+KDNEh4E39FMajjVOgD89Krx3QKStCzdLB+Ia7HimFuhE04z2tHySrLu
2YsMYDk6W2/QWmG5dVLPW8/IKhpgYk752CDsvQsaMTuJ0qSS0T7iKptIh0/DqaSKA0tmRrS4AEWu
UWli0w6euamZzuQv+zPj8CCMEjGCUoPM+RMOCCc+PID1vTyLUExu1Cr/P+X1ehrU0dB5mx0tKCWb
GeJmlRkWzAlWGoNg0OgrmFDN+tpP2WFJnK4vGgWU3c1+iEoHkko0XaCOBOAc5zvMV9IheJTwGAmN
HzoVwTtfjBtc6/IBLiwudOt1C1KXSYyZqjmVtYfcI1fxpTSjqYwOgE39rFofRpu/KybmVuB6C0gL
kMbQCQVGVR9T3pjEB1lhuFSTmaVuLHC8cCXhtwxda4Mr04g5WsPP/OZsRyzCRTanMeh9iexjcwA9
RFxHp8OYucA1EfD2zg2Ni25fwpqrizpIDxJqaab4uuUNbQlo3vAr3w9+BmiynwiAhFFjmhwtvHbf
zE2GpzNPdinXv3SrUc2+NMHtpAnA3L8HDOdGFNK25a9llTA/e40fLYXXIXNvijHaZQNVSBo7Y2+g
IxBDTRqzjX/K2AVKvIkSK6z0mUvH6DuNwpK3vCsO0K2BVWr4ECP6Dzb5zvfmkDgAM/bwROs7nEos
q3ueYDIRqHsEP9Lafu/TC+mzEahB+erkiRCTzORAd5kSWAnTgxxhZzwR9boasbu7Gvsw1m+ypBTr
1dmV9BijjV5EK76dFxlz9MbtE7iTsDlbDG8YGKWHF8E/+RUxs6e5b1kBAGkIef5J0Q/dTWlOtvQZ
BYy4ZV7uH3AGI5bgJVxl8HycNvjNqhMf87Dz1oqyDAeatsDluAQjoUuWB7UiXxSeOFKDoIfgzXUC
kivxxC4Bot7Dqr5XMxSXtu20IfAMdREgfZ+pKbY8E9KO/rQl4fD8Y+HnE/K5KibiU/Bsz7aRkBa3
Yf620CpLyk4Dh3W/5DZ0RvU0bcvdJpKLsPT2rtLsukm9vGwzO+ptwtoMb3MVNbRStY9/fUIsMC8C
6MdpDTS1FjueKoNKVXrMShftxRm0YLH/RoaGApV2qGshY9K2hXFS1sQKohGBtiMrQrOTOVV+/Y4E
DVGQenS33FzfdKuJDLVYW18wSvhM/TvFKJbHgt6JMwQMC5wIlic9x7Bzjhmh+ewh93NrSwTgEPIr
d4KlBwQG+ihaYgWpyq+ypnYmDcEDKwHrqBPCsmmYiyiYWvgXHRU23rN/PnV9mggTwsBvtWvqyHtC
/WogXRD1aGbkzIpy22y2wPiFVo0JENuo+4M4l41cc0D/8pERHKR8I0BJXuahFFIFNgD0+4gYsSB+
/1wcK6M0EKME+fGxRGZ29utYOYEe1jSt6tYbu5jHZTR6hIeFzgi3MSGEvQfanjAoZsv3Tm1NBkPj
t+h9ioJrZ6J3l+WoqY2/9ckrYAHgNPdw+HsEhu7QaFzqa6fKrPi3GnVpzWqugD8Y0IbFsjAccPId
Alnq2h9rTAiropvmWfAVL7mYg3dZ99l6cy184wNIf7U/aPaxOrQP90Mq2W1prQ+fFwDIttqXB0lg
nV6bDJL8dw6QsyMKY+x8B6n5/kqtrFGmhUt9WSwodNtxl9xcFbIgZGafXQ9Grj4TpsRZjR9QMmGF
SBhJTqXS9tK15YLz5sCzxY8kmB2VyRmwGt1UkP1oQ0DzB+KG6a4oTq4//I0ej2qSMl44maaP8uc1
e5xe3VN6YEGKDqREVEuGLjZnrKMZ/m1X53MBW6HEo5lNSx8ksy8Yq4iq+t632YWhQuIQTvnnKP8Z
J6CzJpUEzkmyC3ukA9cGgfadH0Pl5SN8YkBJumLAYv0h49YumUqbfCfTk+uAEJte8HeKr1vG3xGu
dAczg/r1U/PtBR0CGpRU88zCzx5wrYljkYGHm6f4JCHCvHT03dTLHEURF9FiLxc0m/x87QISA9JA
9zaiOqD34MJ2kKlmzVIQKgmFnJA6fQzJyNCuJZR0nRSYL9x/b07mFEsECF4qS0FO8AF0Mrf5cxlq
Qq7R3U2s+geXew7FzF4ElUdBZVh8IuIPLOCJPBRJRDQ6m3K+wwJXmhoYmcX5sLiDvB8pEKSzC65d
NRfBYO6rr3hInoQt/jox/Tz28VnUAFAnnFL15v1uR0kY+SsaQn6wWRN5N0epJON1Vh3MZx85zXSo
Gz3kB0IaA6gh8BYLgapWSKFRtYiSKFx0f8XpBrQ3aAPgrSD4e+i7H/gs/grtu+SYY0ldEvradx81
thJSzJx6nTB9E+rZpoCNJw9f+0H//+IuPtpTeTaKIbMD/I64kFHAO+QYbQ75JOuN0gzD2gEg35sT
2xT42W5zwq7DE5neQ7gF61zKURooLivEtTMZqDXntQzzSGaO49Yt6FfOjcnaBgb8h4xAChHx3F5Z
xbspoNI2VX2NhrNxgJrs4n+Orha9PhvVNpORfzGqTd4w82VOt0UjgRBhUfPjErxwrzc4Qtf17gla
y+t1wLqmtu4Muz4U19Ih4pYXH66XNgZDPyqRkC3bCZJQt9OkHyvbd4DcpnwO63s6YpkBuA3IrUYd
a6dVZLgCbdHW2N38mgNCNhdWrSe3wkvg1210QH7Wi7hR53tp20zGeB3zjKtBPyOt94dRY57y8L0z
Gb2whh1Gexml2ylQ4pPP+rG+IhfKOCt9aVxcC/L2+aDM+08QbaRHfT+iyITNeBGg2u2VShEa9RhE
jKooKkglP3vADzbVvfhS/6TsZ6W6qzra358YhimzFj77g9Jf80mlC2Of8RG+dZR2aWiPR0qxdJru
1SJDwTByPbKRhL8wEOjyHwnQ873z5V/hof9dgzbkt9Zs+ds9IIrwuxc9Yt1lLhWHtYJISJoBTSj9
lkiDla9z70P2sj2+hg5NJ/o+IAMbT32QYAn1vgFSxMn6FA/ai0JWPJIpwlcdfsB8eZiGJ4MoGpXg
DBkINSQ8WJhHCk7GmMuo4kN4s54Zdozq08sih2Iy2hL8qpSCgkOMX7hj1Vw77WEKM1D2cqSoPJQ9
pzOy2FHA9EXjcri6jnkX4lRt21wYNeoUw68obCgTVwpii46Lp/9V1SFEm4rPmlFVLIe67KdcM6OZ
G5fK0u7xE+84vnA2kdKdiJ3kTsIN0ym2WVR2cEgc62OYkXg2G9sMsUX63cudzV/FJFrzM01XtCrE
f8WW/uB9B5qxLNPTelGIVG7CJvirECNXc0SIOmUS3QQsdQ2C5Zv/JZymzTYSVQM81Ko75tHjilVs
2GFhF1FDuICshlg7AViYKVJJxbrnWChfOyL4uXRn09XLM3+7YvRmXwdPkbgMKbj1QULCKcyg/ZlL
2cFHpNqJPm5MYnlrIE51/ESEOMJML5ZMil+cMv/4a0KXFPdy/+TUBTcYiq0j3gFaJa0Gqu2UIb7g
INIxGyj69rteMkBQNzK5Tk8QnqmjiUOk/aQdc1Vl4chmWUIQIUKAhTpkqQPXQ0ZO7s/a1SbmyErm
Tdnz8mVYK/fZtD4rFvUOv/2mKRylvITblwtdygHoeBg8A4GOhjELw/PDREH2bjPQ6+PrWFi9GCae
xpfJNELY+C5nYnYmAqOHwiQRrHLMw1WY75x2yzo7GpvZ4tqj35IuVH6K4WPQF8Ie/So4za4DLhl/
SV/435xE9RqQQOxF2896gSCld8f/uqXuf/SzGWO9uuhibDyZ0LX2yF3QZ0Va6QsduEA+4LCE++B2
de2U6JNHwVpvbr9TYu3GWc+3AM48V7OXZWSFSCkC7uNWu0OaSvFnjBwzBtUZg2hclfbn1ljMXiW8
aduFBlxKm+wOH+yxunsTbx1Lc1akj+bnv6h2iOrpN2hJppCWtfUIUx9OSlcdQcAGTA+XaR9PYY8a
SqvDf0Vh+7Z3I5ikTW8BSMS1569tYp7nhq6vwQSxXOSynG2GIslTO2vRbTM/AUm0FPjYAB9nUGhS
wF7aVG6Ukd0omppeuKHy7k5aF+KN25iv7JvEs36BRhOjxIsuA7BE2q6+AB7bdH1EiK58DByOAf5W
WkfUNnSlgvhFpbY0q8Z0SQPsesYl3F6u1QckiLlH0HV2PUDFtr1zwvyWjDbQLW5l96FcMmozS1Gz
86noRYX38IIIzn794CjuatWhkavqHT91uBCKTc3Dm6JzV28id3aiIn5EHgaWvZvMTg2Brf0xe4OB
Y13j1qrHYV+pwp7MkO5sEBe5djl1ghri5zeWRmTwXMatGmHrzFgbrQz6BfsQ+JFh9CjWxyQzFsFT
Uu7jXo3sGQrTDu/lw8YZNINVqWxJFmbpTFp9h726Fg0uqJQSY+bKCLyqy+c2tQj3tm/llYD1flk7
D469J4qtbyij/ULXDb6lrzfEhsk5ey5xjwlQcgkzScGVF+O7D0rqooF3dgq+Nz884PWZiPpZV9Ji
crMO51QcuDjd45gYV1jjb0hgXwBYHnBRqhH9IF63laTgtBMbqfbWVmxpWxZabQL+4UqC2ZG0/di5
XBCeHbQpvGYNPlB8zihXzuibaU0LvAx5npIU48tfM5il/TtT1HID+zKpHJ6SRy+q9vZdTciHSbhE
PoG7o9QrRJSdMhmPz2lgrpW2K9yh+JBGcFInuI/SdBJeLiL3MpDjmdjRc1GDZeIEPXBtk8S+tATz
GVxIz+tYm+wZVSquR4SdGbZO2Sr9BaakCtrvcPMjdTj9wW/n939qwPUoggZRA1KHHF4dE1mJLBZV
5HpEh5gd95/j5Rxdr/PlY3dEpjBJu3um3d/mcn7yGOp2dKbm+EzN6cWnGHxfQDfmWkEcskgZ0NvZ
M7UScGVMmzyuEwR/RmClhfDlweV46FGYCO3LStpgsT55kPQoym5lSLibtwoxqd/fETuZAB0GDvp6
I8ko2NKwJIowOOtyvSvatsCOtHX7xRJVjZ7ZjKCFpL7Ji6VkSa6Lou0QmEVwvTXqqouLBuKd+znn
56IbJFY9IjsAkSC9zVT2jU6D8NlEq2EZSt6T3BoFtKjWcg9mY6yLi9bKJWsQm8aFyC2XulFEcTTI
9G6OUgH7fjt/F9iVvVSmH7hFSPR6GINd+ffCDhwT3/ahPQbeU3LwBBo20k1YdpG6o/R6l1K3KuAv
0Q3yse1ZyufjP4xxmgm8KB5/ziAqnu09tqfn8aHfcz6dE4t2mOqP8mqH6HKwNG8ohUfTNNWroZ3o
OyQwm3afuZNOlzCxtb+cypZBTBEABg2ejF2Uu1Ea0DSAutGXUupGlJxe5kWrg/9IXSJ/8/ThbRMJ
CUD88JmRH1X5DscQaH3iOlfkAEo9Krx8r5FObwsuK5W1tRuObc+BeMMfvEO2ZIs4sRCa1/CIhHGC
v3zCXxK1W73kxKoGtAHpa8IKk51Xos5Fn7kAuoTrNDLX/E60oAShC5ZUqrK8TmmpOLRUPjtP75c0
MVtVSLPwyoVl9j56DdcoEvHKMj8Enl80Ac7vxogd78syRZ/mudFXeiX00TB4vQh16564xZXtmD4P
KtL8jVlREJUAx6E9DIogiJ1Y1J9TbxLisTypj4sckdkEo3CKxKybcBbRVQbJqPThFAmoCwYC0X+R
pFcs7rPHMd7hf4SuI4AH+oUKk+PzMrLPlMCAlaYgTsBfdVnZJ3y86ewPFY7BEdrm48Ko0dgZKUWq
aYK/pk9Alr2iI2+bI5KGFmzBQZ51FOurFbk/FW0OEIBHYSkz0cAiHVSYXU+nowNEXRydFDll4LvZ
u7a2I4u+iMs7hboVgUFgVqWn22wjvhoAqcYuA19Zh4goqSjBVaI2LrdToF0AEOEN4yLgf+JaDJuZ
OcT6T/Dy8a8PvQbsOlzvGQPF8hKU3sukeO6naxUiHV3mlk2TIuj/meZ0sb954lx2PPbC+6ZbqlQC
nGgDuza69fhDyeh4TiTPs5jn/9cDwaojgtx+paAuyRyWiBdWoHsJj3d5RAwvuszBSri0MLNbMZzj
vU625cfIqgQT5PMMP8c48+XLOYYmaiyvscYQHDKCtyl/m6jSGqt7sH6/hzh6tu2WwEicPsX3P4SU
ORgiaObx15K2CJbAYtG9Updko/3+Q6CTsBljyyI+Juax7Rvq0c62/VuhFwscP2qizGsEzTMWmSnC
6BelXp5XnbbdXTEd4h8plniz+91EYY6xRO+Jy/XUnPTGFz8ceahE+sKNHY+SptnodTAAI5Zwv55H
Hc/DfoCP3TwRcKs1eXB+rha+i/Paj6Bn7vDe588wBPYmljwoL5agZz1dG4Vn5N/SqZXSaOiK88jG
rCwU5fD/B4sAKBs9X/dEZJF6atAMN5u91qyyhXkIFccQhB7niXBibBBgvKtOcvggVC6FdrPMy0+0
Pv0S7gE3+hZ04q+5RDICiZpozV+9W7s8n38+OwGK59yU/hs+tXXHiu/gY+R4HyOvCHw3getFawoi
iF9cLW0LR75isQaGAb6tzIozefkGizM3vftt2af2wm2owJHXDgbopsoweSoxnLvfrguWN9/vSDcO
4p3rfASCw/OrsCLutvijIubhk66WtpsYR/YZY3ig3HKEz0ImB2GjL8JU6SOCHe4luGmM+xNLiRX7
/sCRWb0XMaPKy3hXWV3g+ox1kedt3bDscHlfJDOYq/clWNanXp81q/z95P1nVMH31kacijbKHCoJ
H7h53vkSGTuhUcnHD/Fzq012AIeq8Fes0CRAaW+WExl2eI5z0fIA3UYmgsTvsnyHm2Oli4MlFEmm
1uJfHXmyJmu/UvP+x4qEAawstUIlxAGoAag7Cg2mq3mhbFUB3B6eOm4AujM5E1Yrx8N4oWBbwStK
XYVmnuwMIVjZEr7j5e5+AdCGHnSYoh7N8AKqBxzOO7ttY8w8B8BVyaLePG0My2Cm/pM9xDIYzyLT
BusbSNbhBaQwMSIobAllVWG2z2HMH0ps0ch93Hsg8kzcbtWjzplQbc2Kq3U7l41z5EdoeQs65NT1
SCpgP3SMVvIUIgn+rtYrONNdOLbvHzkB9bP36puk+PYet8f1ji27aLgMnkCBwy6x53vM6MxsGPHS
99LrZy/9zHrw1Ldb6fhC/jPTUHJTDp44CB6+xBBRWREsvXY9A64Q4byf+SAuZa0Rb9R9nWa/xiXq
4vh5TcHBxecFkGRqByYugWaUnQzP5h83fkjIuujLfilrUwpe07MekPHYA4cpT/YG2kljdARVRsiw
3QtHQplUlMncUUdqmWh6oTQhSJKOTQ/oAP3NKgnyomYMqw1BZEAJefgSPtG/Fc+rh3qb5QxqGJbO
iXUvf+cAt2OTg0ZNmhZ1QzsVwzpojOv0hpYOtUr9ffeYRkOhwLH47FSiwbARGDtVsiGosR0asItx
OAVp8cZatv6032fBPN/XJK3WwkcBHPgeYvAmEDwDMXkKpecYOub+GRQDd69Qh+eMUc3Ur/LWyKTi
NksPJWEqhN9QkerqunduLH0FGkNcXnEYwfkV3hdcs1W/Yoh9DGISgOVJEhULjA8Fkgsq/gMXcRhG
vPQByIN3HV34skQhwqK7xxTynJPgT9w8J0L9TjtzSMneCFrLY2cKdfS9E9F8UnyEjvAdFokUZt4S
ILM9WD/YhKhOJGNRRZJp9A3IWWHDwKUMSbHR+aBp/xBRV6oCjMx+JJGZPjpy9SrsJtdCYYwWV4Fj
GsgXPGBINUTiClWMeYQVznQ6QDqskO6PAQKtBV862EhP5VfRFzkSz8UM++3gUkZLH1EHInDBgkyH
8sXFUEr4P/q4P+wL/PwoFY9uDRohqc5xg9ILoiDNvorvUymGHZxpHUo1+CO483CVKlldgle39gyX
GbTsHRzCXb22fEX8x6GYDNpCV3572guDZwhGIyBDV7XT5uQaT8VaT+9QxfcAJEpvu0uwKAkE0XTB
h0a0NSRV7wwdq9+ZFS3uK0Yci90W4LaamQAoUuznUoC5itK9tDWM6uz9GyoKKIhYSglt5igp0rcl
kXeiwJlaCMLB6xsN1O5SZqVPCcaxc/a+bP5uL7Dkr9r8TrFXmPMoQCJ3FYqyNaEPbOlDQ7g3xEed
dsq+eZ5JJJxezjwMLcaeMdfW5JfP30u02jaYeVRtMAaYlguOpTIZsmfwLWE7QoaXkEMnvcCYFTvx
w0ScNM+zBA50MkGFhoVa5w0ad+ZeCESDQe/eEWONQ0UZTXbqFCpf0iI7BhE08MdniAmTFrNHoH9m
Pd5jT3JFh5H6sAO8an2k2Vyo0VNJ7Th6TNXdYx1Lp88ryOk4NykvPjlypc3WevRePv9JmragUmFP
u75MV5Wi0lOiyma1NAl8BoEiXDQejsBKftmF0maQZUscfcbN+5MMtMKRMcdMv9d1eZ6KWENFZWEk
BxINYsms53bsT9qnwY6OnuOyyMZw56eSUfBGfzUY0NvO+6UNKEQfwvUsmRVyNFRW5J9lrzU/eZTe
td/HYyhyTT2k78LbaMgCp9VdDfXfjYXV/Bbk+R2T7xtgYFRUAYv2EfONpENQ3zSXlqO656uzsjoO
0zNbDv1vlWHb9j+BEwhlliePFS7OS2loTVVccEYYMq9airRngi6ofLglbdwfKYttABp5xZ8wsuMO
vRvZX+/4XvWRH882VpMTMWgp30FiEHaQyf5zoYvhCJ9LRLnRCFekaGUHKJ1IMhkmyCAb3/QPMFvc
Y4Dci6MzJaAPNwt7wGXC8jYjesPkTXbqvxgCLibpbI4ioq32rMgOn0e34fu+jhJSTPen4nnficee
0GshIFnpxfJZpeEAMzTUamgoHZZH/LmqGAe/M5AEmA/QTFJ+xgeAx/b8430v5JKRYXXUnZki5U3j
mPFjUbMQS1UNPxG3S4U6viDDoFakV+tHNr/Bpdd16XpJoc7JJaea30/6CsdMBmt2G3nONTGe8Aue
+EN/JDzoUUkKlwlwtSkWXtKGgCxujqSgXCYfBUbWqd292H+QSgGvwUWwws/PlbOK+TVrJlVXS106
Fec6pbF4XLYHgJx0m9PM13mHcPgTDRraChtypHi3CkxHoBxkiZlJs/hJl7HX+1w7eb7jf+7a29/h
vBdYIbz6TzSWbh0mOEOBkWHoSzc6DeczfgvxSLNr6QAQWRisjk7AmI2hgeoO62nRw5SXkhgub5m/
M+IE9yZg44ibeO/+W0OfQDLKAvmQ2k8dUl5C2+rwkDOog6HwTjtJ2YHX4uI5mXvkaWj5wZw0TY+R
YfPqVSMRPXKeXsN/SrD1qVC+XY0Zb7ejOd+zbVnaPxX0/SYD9Fz8r/qVEOAGQnYLV4oSToY6ahqe
TmLby+A/5l7xpRMLMnIDerukkp7ujKEmGTr/0Yaq6dnlWRsTOpUFSXj2DxBTjBTBo702NKsIe9QM
Wx1IElpgtM4czDKAa6vvUkMBv+lu63IDD8fQaTvUQE4TWGnwYxWFS2T5ptFORM9OGBnb7w4VS2T3
Nz3sJrcaURQQIgeq4caA8kTp5o84H3o2A73sQcSfQWWdUSjrpYtkYEgmdgHGgEEva29PtLD2NKAF
cuEtWXc3qVhsYVnManBJeLk6TH2oqJS5Xu5tEiIdgnEA7Gd1UpexMgNvsVdAy6n2BfZXT5n3FJ7J
l9Xg2BgnlUQYJd0KMiy1OhNJk4+bkBhDlXeqKcJmvZuQcmDcLCF12X/qlPkA/FLRIDuctnxRv54M
hDm6NNpK053W7k+u9Scb9Rlv4gbmSUB82IglKn7q0VMAjP0vKL/7EcPe8iigCsa2ZjHAyT/oHlNo
NpfQYCk5NIxOi7qmc/M2Ir/9+3pj2/2Q5PJFXdNwaZ6Xf38Dwz8vEU+jaHDSzMSlpu8HBb1HagM6
gUVYGRCnPA/ASIcHOqeu+kPOKCSoMPzPq4N0coD+pYMp2Q6iDUhSSFXQdvDYIrkI8mT0/rmQuxU4
b5goW5Xma1hvoEVKTJgrcuFD4Cgtqw4qEt+rgRbBU5i0/O73EfEFjk7V6HPlbM6ObqS94Pm+EVO5
ilCOeuxxmW7laF7pr7HvZ/oUK9rKK3ZdrSHIoQSIpMLGdp7qQ7M9qwi86QKEzScHSF/7I2JOR4iv
pNC/rWmFk9GspoPcBIMQJtnoIK9M33d2JruCklK2umwlYZ4bh14wV+zUdukAl4naKY4fkoiB3S0z
1mdG5/W07a2QJdNW3uA+c1A5pJ6mq7k/YCYz07Z5rLXwHCSze+XEJ1xFXVi3klrxK2CpOrBlLhN3
0Elyt7Rtvk/EPioucfyI/hImEKZHu/JBxcfHJyPwO7IcY35Gnu5c981MVu4Vx8G7uqikJfhwLmVe
iQdpxctUvfLtHKpTWjIreKZi7kRw/1xCvi3bfUPEbYtkMMkktgaOQvzKMjQf/QLz5d9p7jQGiicZ
f42sdPnODeazl3rETzfXpCRd8bimuKV6Qy4AjU3p20Ma7ovHee+4IFa793pkvfOIPEiH4cdZVapa
+oJEtTJpEDkmQ9bavhmScGyIM56bRGnLumZI1RSaOcmU62qAft33kVNrtr/RXCs89ie0ntdOSiI1
k/85nl3E8MFJ33g6X8ykxmleRaDOFjkuSnen9DgDIzgBc6mlqmTCUlIkeS/6xeJTU7CMp+eKmPCe
HTY5jNHoh1akogVzUEd2SbH3ddmfaO4OHjkQNkLWUuHskTqoXtxgeK36/eWgz2m8SMmxP83Anjky
7S5pRR72bD4ADiE8KdW4OGy56cWMS8Z4nA97cW5c686tldKHGokxS/KVSTsWgHI4vl0+bStFOns8
b2ZQjdBDlAQcjXl6hRfwBN4iDKuxphKFbJhgEui1fbXMhsxCmBeLNDDirqhgcUVT1pvsMaVmURhd
l0eCBEYRPwJr9PSuTCAqB1dikKpRadYcGk3zlRuW1EGN0QfHq7qA36eZS99LWe4cFjTR5Eq44tY1
m3NLOgaHUjK4hlCUg/Hccmsovhc0aDlvxNdXRW2pbdU/sbo8ivfbI4tamMTwtCV9Mkl23mYGtYWl
U8N+HMkwRJT8rrgm9Hdxm10WxA3hvl/ej1IUu+B+lquA4/v2Wtbkf+UKtXjpAGPOfMPfyZn2VXIr
/vQi7n5ezf5CqV+KvzGGHSb9vgYw7toDWaUrPl37pU/C8w79CLH0MNP5Nk7kDZ+Oa+7kdwTPY8H7
mZSSN3o+gdJ0CPgXWu+CLxnntNUgMTPsoN7qN7xh4n6TtD/tPyZXWN2l5n1os+9XJmXMtZc7YoME
+e6Qn97RFIKnfplnvRV54xykIRy5QEX3IP77iYrIHfCeX7xbXwssbFcquL/L4sdOAsJgNp9FfeM+
Ju2UeOhRqCq5PEhzh9eKKw/oDlpDbyegZ9/GHxRu0bt5iZc47y0B01VVm3ZgMnKuGaClnWNM63Nt
dyZa/oDGyVdFEr7WYdn6m00LpL+zaBMf+6Sq4GOn6ApI2PWS5Dq1vt3kVDRE+Y7JNRFMzUt1SZPG
JnyFDGTkgl8z18HvvMi198X8QyTzqIOAGhfoT1QGdpQiMDsusjp2YZZ7kIlrhLjRFxvzn1uKuTRB
fuqtP3RAiSTwTCHERBKjZLZ0S3okfmQ7nKGeiUe9Jv4QUFYVB7SreHaqopSLPGA+5pmdAsIkOMAq
z+Z/Pp4Y+oHFtHrFPZMdc4UZEhipmi3cV745hjdgYyoW6VnNshC5hx44GOyCf6RLaXsu4bHbcg52
EoBWNmwOlBA42IRGoXD057FPvFCUMMbY4kvw5SWUWTZQkEr7rkMip2vOpAQAR7wvUEWy7VDvnfqG
NEwPRHjy1E4C+f/4zVcZl3oUC6lONW4XTmBvAUxESFrlcyu2rSiZAzIpAZx+W6YnyMwgmrNvF3CN
YBDCiVqeE+e6qhfzNKHbnjogURWMdEosGXOMya/nam+eBwgucBnwvIblAY0/ttQt37tD9EYZweAX
vZ8/ymZI/Ke3tBp8knbrGTBVEf75NRaV/j5JR9IFe0McUS0+tmRB4gxmfRGBQnxRK0aUw2h1RBDD
Nt31duEzaLUizu0ClP6zOJfkJUYq0/raIgNf8vy8fxZRp57PujdYJ/CUkz9UOUpv3LqYjGa/dzEU
93tNFdCruN77EHkLgCScHBI/UkZLakHPCGp781zgnx8EHHFjtRUTReZaMOna4t/Lqp5vVVI+03/l
rKNQkT+7jMDDZ/Rpu7bf7rJRuIAPeO364OswvlxcldkTS6CR8mpWNc1C4SEozf1V+WXr7JxeSC1m
YsaIocuCGC6D+pv2AYfCRq7mdoMOxMWbbzJsy9e7xjsTajSb8Do8e6jRz+oxyG3QoeuXPhy2G1P3
osEHFSMKm4ejyn/lqELpwDRvrSEte0cDDsMD381O/ep/QvBq30Tl9Yx6MP9ciYe/O1xl1s01mNGa
KaPHLdaeFqreGCeAlowKvbgi2JnmF4Lq9DIE/B1QU9vnpHFECZivH4jzITdcQzr/dVet8r1ixLv4
+puksMBXSXbR5haWZRMypxvn7RVzBpWEFzZb+ekzqlTvG4YiE8P5/WxO9F0Hsw0yRJLNURYCViiI
iUu+T/YvES2jF/OxgJRsQMgmCvMYmGBjOMnmLEWS0rVwKG09wbppG24pQN8sy7NXeIak9VPFtOrJ
BwH5JU4X94wT9ByBj52x9rmENw3vMag/RZPUvvIXU5C+ZhFgrPxE+iPMRBt1c3SdFPw5DyrlOaP9
HAtouSkMolPWfTtqv69Rxn49ZGazj3ztsbZHu11RXkU1KO3sBm0R+j+zXFEzj6KqCNrdrny7DVKh
5YxrXY9u39dYnskCFqt9rgd5oZMaGIZ1QekzeECNxGxjlW4Zyp40uXjQLgYC1KGl7RSLGnY2bYES
KOtsjOsSRVOYTZ6CSDEI1sufOkLmz9U04Now5KmfPioNp2tIUqB9b+3lIvj1nRR7fC/hUVyeITg6
ZOoFr82k6YVkfFFFUhZsPZTjb6MPn/G6IUoIS7imbXWqFpmxKmNDzWPtTLRn8I1wQTFw52F+vYJX
yEfoybb/GB+8Kq/8451hnlGeWhudmVsAY3Q530jfTD9cu51t/9VTw0AP0KA+rvqQb/IdU/MMvcYU
kvTmhuJL2OBJk1EAmS7vYpve4LhxWGun5uBS+zPl1gCaxAZM2wTXUrs8SNfr4vZhcHTXC7+A0a2z
+qSebBWsHB+FcwT9JIUbB+iX+L6K+3vwMJV4Ola0f0WxSLxl4ayTCHT4gn4D8196NG0PGpG+0bqY
cOgAqpMIFoYpereCkjGxn1osjCl4l0WRtjclwC13zoKQHjBzAw8k28ikv8VtWD2OrZXCY15ot9bZ
Lg1E+rW0tHrkpV2ppfbhY3KC8KFEDByzBzdyeX3nqoZHVWnH6r/kqVsM+ypkN4/lomcptw+pwPl9
3uG/sUVX64LU+tdaVkUYHZM3WeXpcs0sgU7iqTdEtJGW1OtOCNJo/YSGkcY1mcTt2BbOacb6cNAj
9ayKIBTFkljiwx+oB9Ib3a6mDMcrLYwwfQ9HzzIavyVDblVdz4NRg8snCVGe95LPEMwHaRxsJO2Z
PGfsd9cyEzJKMvzl4bpGMA/7dAC6Wp9/EWOK0F4l1Z86m2DCmJkkGIX1m3NXVVz4/l7PoatWb2hn
u7Od2dhw5C4Dn8PBAWdCn9WRcN0xUXo78tv2khPmb4VLA/6DocBRND02juUkVmIEZ3WRuUMhJZW4
hMnHcc62Y+mL6e1T/4tCuIJbnjVje68K4oWKBnuSol7h7+6UbR2e9098BveQ22KJqmeeezqWzlWl
LWUV/Ji2B3mfGoIuRrjnlxhDSWTaAM+auRpu3JAtOsDVaqzBMZChyhEw9gDwZLMlvej6OO8TuFEB
PnnCuE8en5y1ak0sumoRNpnuTvXNSVSUblA/a/+H+EWiJPI9KcDPlylie+4zIFcSBCZn1n9q75F5
9aw6rDWSUG+IVX9a+f8mtlfb//lqPr/jJ9QqqfQ4haRcq+t3TpKH1ZvbXBw5lQriTJZWQPS0gW8a
EsqKsH4kxdgr26P8MFQy+3QPNrjgibSCvVOvg5Ik3O7jDypFVb+j+LRpH6gKd7z57F7aSSlnEz7C
bADNURzY59LkOm/+til7jH47HlHT3Lq1fd1aDXSQ495ChnT+Dkk7KTTxyfsGv7zp1lW+fQlMxvye
7Te8v8hjUsgKgfLNHH0hAruGlkH8g3tv/ANZJ+yY8ctFA2KgTE7n+gES0wbczPcWJ4cmOtjidCEn
G3arOnee+ALlctCQipqKthKIPpwKkcCHIes8bLpe6ezTE/qtiJue/yyJUSeucLtD6sYx+PhBayLH
cy5/6uc8xsbUTI1dN5Cs7CR63zrczHIWC2/M0doiGM7cKQdQR7AqVzndGIyES7s12/tuC3O4HzT8
Z7hTQBFT5YJvcAkVlsJEpEr8QIs+JuteeqfNeG1yleSlYmPY2zS708T5Pbr7VqFjQ4/ADrvw3+lo
Ptx8+jTfM2ZlIj5cK60K1xN0HO7qmG+O2Dn8bFFtPSRsyyGCpj22+Qqv701g7KDHvgggzMj0YHh2
/qCYW/3wZuqlJKN6eklLg8r6eAqH1zob2SAUMThuClKtPiVAJxbQP5swdA8xVKFtwf0UoBaBG8Em
pQIs1FyOZ2KCpj9Q+4J9sZHQwd0U54o62auyKa+yp/X5nhMhUZJJIwv/hotfn6W1j0pnzxJZjDrx
BP6iLIfmZ9Zg4FwRrRtmo74NUEe0YG34JGCuRJ6COGSYry65Y4lnvtuLxOGiU+d6+ELx8fCdQqlx
dF5N+g3E050/DSZBIu8nBX9Tzi+PRtSJ6T+6+UdPbSycV84CC6Yfy+iN4tvbeZeAx2tb8MfORP4t
ZLKVGOeN7/Y+cWn2LLMrh8KNusQ7w7+MdzhILmGuixtWWf/DN6T2/2cVfWsRAnvHWq26rv4zkIK0
dwn9iEkWbSppwd80O8NDJgp+O0wpiLpGoCR0M6CefVidJpANZg+CMv1Youz3uTG1ti5w9z7KYcdA
xZ+LCOwlFkgIpOQiqulPOcSeFLQPJgYVl/2QcW9ObSrdnf9sBSNMXUhN+QUnzu9Kj7F9ZG7BjqqO
Tr8soWuAtRgt+5Xf3mZfrkD8nmuF0KZHCm5C0FrB+plqjDSog4feOw+/Wrq2K6vQNZRssi+jikuh
39F4wJ3MZHx2MJQtYj3kTAdI3mPXODV5pVPYO2jadERH80I2B08E9FJCktv57qnwZbaFKL28GJqB
9tHQJjYo+NiKHrg7Zf7VtMyEuf7V7XjATNSatZf12a/TR/nMBXL2HJKG+O82WPqqy7+ck/cPjz9m
iaNiU/zfyY/xzE8TSIzQbr4yL6hDXVO6Zf0gTpB0V7PgNcSqCSu47+fVLS2+Nl5lHDDHER4Rcoyo
z/m5KmyfawfgAdgZtNl3F+qp0ItlFDtPF6/YpeTc67P7xwe2W44xxrKXRHv3IOreVU7trAXhmXDM
OJCOqZf+OySWa7FeqwyGmsUOsuDo7sC9itYnMYOq/2/NrEKviDupi03UQK4qA4ZzFT2OQPVQj6az
Ptnlpc7d8X7H+vrfSTxvEgBhmNMJuFHEN2hNWH6wdQNpeKk9m4FnNKogjjmilXQfMtrUGScFszxE
b38h/AD3GUoujZVQkD6Dvf0ptewKSngQuWp3ClcRwtvkXKVXbbNPDSfmnVkz+E3qMLSoDRjSPqev
scHzzYL8e56QeZYaRbEowjAru4awOAm2dex4qrLuK+ORf2gKzl5B5ThxSf1exdn0UnP9TPu87FJ9
aIuiF3k0dR7vjwqGMfSDF3O8I09U7HG0meA21XeH70R79HWXu/kvI/AB4QgIOYzHkvh3X5vI7HxK
H2wzh2qMy28KKs5nbBUjdgS3mbFCe1p82WtNPvCAOK6LtKeGp/CCdJHsY9Vxcdtbz3IEoNKvlsd/
oEse5B8VaUzQTy58MsHfogQY8i97sGmogKHM2VYuceJdQ/7O3/NqOr+vVZJoF7AXwPdCKsj1SADt
2ahJTm4Y9jkHO+GYqwloqrKY672hri/q/a6tKb5+xs3Otbq+LJsdvMnI0P60SHLyAR2vsmcyMjLZ
2xfjnVWgTnXFVlFDBbv2pnBL+UH89ijXpxAA4sVkm76Zp3B4n3BH162I/M+afUgblspCMN9X0Tfd
AhF5JWa9wuCYOK9k5cUs5jCjZG+14MUBlw406j0+k4nRJ9flVdtT1kyL0+BSDJuwkKJJ9JaDIgyy
Ydu14C1nXvWlXDu0rz/4QjSM7BUhjYkqUepMtAc62edbd8sLhgsmVefKyt8XjpU4PGq1xiALjwiH
lxA5qHQSwb376Z8cUc5T6VfumNV+0/8UGVHABH+6Pus4qFgzgX80cl2RcNuU4imMHtBWJg/6jdEL
nG7G8vWroGKMxubV7ISm1y2eoxDS3CNHeKfRtJXh0VtzuVhhxiAdyNrGX4yh7rGc5t8G8phMLO3C
MQ2d8woVKq3dIWxdRkob0LFuCg7bXD6d/IwOqVjH3RNl0Cp8GqjEwpQIfTcV9Fne4zTYX/PQyY46
DWPCT7wEqG5fls5L373CT+sK1xBQNKrPIlstaX2vLbGfCzWhX1bS8EhBQDQumLm6G9JA06GMOsCp
Aknlhedjfw0z2HjGuRru5npm8koDoc0gnsGdb/XTDhOJQZK6mjdMqFigHPoRNZwAqhFFYcbtupP0
EPCr1X9MwXeLFnke8AFgWM9VbIPAqgxxkey9iQ2Ba5RPkJH853+DDTs0Y13OAnKQOGs/V9UWdHGh
q03GLFiakdxlyeCYKJ76kVbTVkfchNDZmBm8hTaWxqIZbV0PvtDkO7BIcTRU7A42WJVRrpK3RoTI
fN2HCy8ofSYFijpH4P4UOZpfM39wVvvmrJyo17s39SV2sDUHYpQSI9Xgku2Be9Exrs3Ftt1qq5LJ
rXYik+ggz7VzbSwAoWvozall66KXVdM5AhYqMA7jBcrLTgJm9sTBvtyCcnxDlLwaGhNv503ziAop
gMBObX0zK0/61eHq+kRJQ6KAGAENhFYqcXG7WzKvfd79kDetyCIy3yWOG0ejjwtLC0b3QRPhZ9NH
ISUATqH2v5DmYoTZsf73yOKSHGu/4vrqkFq7lAYfGg40pB/4lh+zj5bKEBMF8hOT6NMnQDN3SNG5
swO7xzWyX7sQH7dX91BqRBpdBOTM1jkl3uZrXs3M69gS/jSCzLvVUzu7i1XV3YOLtxR9ck2866ni
vRhGRXMTuqOUCbuBD+2aU6KazAioiCOD3sMaXzzXusrw5I5PtHFARl4VenHw2sT1cpubwXDzcDhA
Y7lzjb7co/03DsX/XZUY1PA+CYyflfEAXPGNGKn120Msy+QCqKl0ZXJKcgnjXxWoXP6J+n9tfW2L
saRMOz8oZ220r5Hycap0VcX9b9KgdHJRcv8nE4sc5kYom4wk3hKNLVT4jfs/cj77T5HXwFoI06nZ
+6xEtui8+EHEaEXL09Jq6mAkumjRkpao6EIIPGjlBE567QopyP4Sm85LaBAO5POBIDYKny/5UAon
bznDO2auCPuoUcyy76u8RWFCstTaSUSFyHWOzvDg0SepANbiagZG9CTkZMmC1R5/ASiXyyNSxfS/
BRV41i7CTqvIxrnsucKnRAJw6mfTf4hiw0lyGVb4iuCTTlFEIMnGZvIG9QWPB7eRnqUdff9UY/4l
N9zjloh6TsGjAB/k/1iR5JgmqZ+W+erCu0VDk6FuvjPJTXpbsS4baQSlWycBJEHiPtbOHlw3C0KD
9XrdFxxtJnrW8xIdcK4RMlFDn2c8ocl+pnt9J5kYhUtMkuSqXw6IRUIZLRnCMBXt/xSv0eBmrhmu
Jzuxhq02bXBBcUvWU8rt2gz99Hv9NjhDHjipm6SpLOVF1EXR/khOuSKaf3VCeVM0Dll6bV9r/xq7
UGYfpbqdCUCrTiMotzTPSuPVmw24e1u2WQxncKvy9fdSyGI/22zNQu/Sx51f9bSe/R+FkQwbnDux
J6t7kBMUp8mlDhvJ4RFcFTmnde8sE6b6W8Z3nwzC5IuPEsODNkFKT7XRQUMXu0mAdWdoywQ6vLs1
Zoi9RvIkmI6AOab4cXCbdQDBeEQda55qAInWAVEllJ53biX4bB9TNj3613e3SYlQCl31SD9Rl+NC
gBvFbbce9UPMwNfCXASBf7z8SYL4/n4FnBB8EYe+YnOMGOHUdY/Go94J6PG6Tn6GeyTa2L5GER3u
Cm5HnTRRMlECR247ZneAUv/fPWn5s1lJPK8hfH4yS2+YnrQ6ZfExQHCnihUvfwGtgMyY1RhCZafJ
9bc0S0GYOHVe7V7EaODDrG6HBA6HmWns8aX57/0MVnp2IW7LU4DfNpMojveg46dIWWs7/PYJobM0
Vf5K1nep0HxMyClOCh69uKVJPIe+r4zrUGEh2JvtoMHDKPKFlAmlbT3mKx/llosq4CZb2bVQ2cCh
L2xr35XiWQ8bfMsGEs+DAXsQx06Hf2U0gd9hkhQnrfDkgaiiTsZtRS12Xg663i1WW2Yuvi6A1HSW
84qJR+Tco3ukyIY0dsLhoVNKJBwlPYPfAzWDmxXGIskropox2iavPLPIhoEpcUYk0VIyGej3DR2W
na00m0yH7GE3sUUk/Udf9mL4LcFhDmpdYwIyY5m3XXf8MEndcKCbj/Vh4fo6vAW6DjKN9xWTQU2+
e6fCODMWyJwTL6g9kjhbNemD8eBBTXfpyfLY1X30frH0/zLMVFOtTMiCHEj1Ib2xPJJnCS6qDSSj
O2lZfoncZegilEBI0wUksrgKZwP2m0pKb3sw5TISEtppTbVpXBHf2kaWBhfIF7VQ+lB0uTR0EEDc
zUmq/1wCkm/zAHWd6uDCjddQzM074ZHnZdl5LCWDBHClFjJkPGTdkHUbhK2zly5T8x8bX1s0VGKb
e9hj+MoNM9PK1poj/FItMXXJ3K5DZZOh/CL7uTECryb/Lfi6waRlriczVRLBaRZEBNdy4ULJNnSS
b/BvWa0tfeK/MqkTzjBQMIzK/H0C98ypaCFo304UQ+nNb2ADLEJCdS4S0mCzCuTKflf/NgjeeWSZ
XqfO7xS7UZVhFkENxWkSREt2wm/h1P8NHgWfUzuFMMKh/2zRaK/cx+JKflf70Egwn5CddvPpWk9x
5w9JQK0QLJNMWefxzrDin4cn25i6zj7zINcaKsIQaOimq5yd8Kj2grvDhLWPwZTLwsu0mX0OUSTz
afr5GQPR/m4CeAqfp2z7OSu1OUVmCgVwcDqw6EedwsQpMXYu6u8andiSk39q7ihN8RWwnFlyEWjX
xpqwROQ02uMhfnMamE2RHsoulEWnczWd0JKVUFBX96uHWcqBDg1QHRKurcDlFHFO2W8sSkHYi1IR
Tx5VHLDMaX6jvZ3Jg7k9pq57qFljrvij2xclbBkVLlT95sdoWOTmm7n7BKZT5Gfmwqo2P806jXxl
9I16H9B/6JamM761Nbrg1+4dZavh5741p9Mj0i7wL0tuvU9kFvbh+WOs+1yP6UcmZItEp0dq54np
Q5FyV/txRSnh/IHCklq+THsSxUe7+JSqBEEagIdJLJDsJe4gJkHkx3au+3j/vn5sleRPkH+Cxk90
F6ar9xgG1ytMFPYlpH5crB7Ooi4euKmGktgjLVEEsZMZwbsKD3sLgboVYa0JO19n5s6Ig9lRW5Gu
I7JY5sgerqot2BR6aO4VGQUAeNQBnmP49A9SGiM2hEMMC5yT4zukaYwRMdcbXlsL7VGW45IXvihE
e4bGbijdn74ljYGBeyNA051Fs4QKN0rd3aCMRUAZ0d43/a4IjN51KLE3TR33p9moQj/e7vtobfug
tkkaUTYsbS1PNNopPEfgGE/1FKcr/zhtVOtMUMu+QoN0y3aHlYe7w0b1Irf98WEvQSyDJU92yk17
aoweCtPIuDB59r56HQrEwj/Dwq08faqQqU2Xg5KPJQqgd2BPB/DLRbOSwvVPpMZ0zZgW5I2+kyGS
yB00vO/wBlHzOiqSlkFFDfwompZQa5HdeQxqw1uVLdS0g+7PZvM29vqoGyJDv0I5kdptXI78HLnF
fgLNk6y0ocbU1iBBhHkiSwT607HggOgefj01g7PNYPCF7OKszmmGgy7xx1IfmxHvBlZN3ZQ2kzsl
CqdZafaWQsL75teoiTyoZw07UBTAztHC2U5Rcspa7yCT3w4uZVyWPRr8Do2H6gmgm0nMjjtnwCN4
PDRWhlyarTFnEm9viRXHml4bs8DWWWXATZz3w1S8BvjgbCf3TSSQ6zRuGuVdErlGrnYoxHFYjH2D
2cLnsW+iYDeGqVJ+MwjRj0DTY9nKS7zhNTqI7Zvqbkma7eYRiUxb1FIBx0lEs5mUhHVMXQBQFdjX
hJWdXo+mEi1X6WvI6A0321YudwDIrSY7PMGSIBmI2uw4h1OGwbMCRDwtCFyb83Xm12XoYtwPrOr7
vmtqCkzxKpn+Bvt+WLiGTzIpma3+iaKXsdiUdi567HyqeLDyUTmJJYS6Fxm8DSX8fy+MkFrXmhgx
pKIVl3FpytWQQdH6YnvN7fMb6yog2Dxsa9qYPy0gOsRJM2RlN7EFGPyvYxbFbw0ggiT5tVyZV2FB
7l4KNVnEyKPESdKlVtxkHhmdFtUu8KJpKedrkl1s6488nuDfBPbMQvxseHUFjpcoeaeYQAdpgU99
2eKW+l0afUXhBTXzKphoEDJCaJJ0T9u7q6iKqi7j4OnxYzvCxbzBNrKxjYxaai4EMKsw6p0TXbEs
ZWbueBn+Wv17v//gB6WOTM1wRumrDnsNU7LcaZ4bhkNJ1pM020gQKMg9XXaq71ZIbXBSGrtNOTKk
Jal8l0Vhnkjs1vBJ1RRPTWWUh2KJTO1e/Pp3TH/XuJZMyhiEpXNb0QUObstljounl1RdOlVIchJu
Yk3KevvVt3u7y4ux0XHhK6Klyo9yqKvMmEf8fntdoLM+qTK+WmWP4wcCJD9PCT/VuW3zbzHpaC3L
S94b6n14+n4tPlMD5X3orFZIWg1vW2Ai3QHFbTK7PfDFPG1q5myW953Y8wPVaXOpPZfvA+bSS5C6
FInmTqc4tmKgnTPuDpiyY6PuYx5tMIdNAXboKCFZ8OohLVBP5wapkJRDjFArP64dJqzM6WLDO+Px
pzUfork384PXWyNm7d7I45bhPHFTjJ69bz9sPdNNbG+P6Nu03oU5Wg0FYyv70XQjgjEioa9sW8I4
fOSvR0WmWI7z3CWn+GbCsmhAYjkI9MQM+fWFzYTIpO+o3T5us/Nd33IiS/a2YQk9s4gxA632PgaQ
TFSDNGpkorqy2uGHT66h20ObTEXAgA2H4jy41JNPPugBp+IAnkgoFzi6MMHDRcr+FfsM2cbYYP10
5/nzEt5X60mB9oA5Y7caUrsvXgI5+YbOs3/35PaWbkDugJQly5UxkxSrZbS215/vcEUwTmdoSK/C
kYfyZUXPsTNhjHC7DurC4H8S+EYG5G+/9Ni9OqV8kBYrjEG8zLDVd6zI2jEaXZDVO0DohWwk19DQ
glMD/X4XTOcbE8sHmapV2dayrXkMAozKxST+7mT/Ia5Z2A4vmn0dPpInx/U2679Wea3PQEzLrafJ
6YzdwG3X9U/UrJpOHFIX+x9lmMn6Ucen8yl+zX3MWfijDcp07WpN/NEXKbsLVrpcBh28SDgxkVgf
e8e+1gYWxLhBCJ78DSLVIhy+p2BUltb1IckatsjRVJRA4Wag/LoBYMW59LXOZhMPMvjy9xi2EII+
d7iT0TravTv5I8mvuQTR3IqcWl6O/0jUW+2T/dsPAriG8PCpiFCEiqPEl0vx359CdwzjKQlCHdlz
XbIwniSlG8qK8ODXPBKczmEdaafvP26ovy5A+eHVErnGRl+izk+oIcPkxu8ZfFoxpYuiBjbl1bGw
mis8mk1sZ/cemeAWeEnjP3V3gl4KgpfFfo7JqYZAxUYAGqKf9GHLou+XZC0s7Jsk2B1Qwh2dgmDW
WlK1bAdGj9s8wnZRRI2Nq57ye2pr5kuyB4inR4iPe02vB2O85WQ2+QzBvmsPRuA6tPhSxe7COZJH
eTjBJ0e7o3XKQp0KF+zP6GKVvg6EHfOlEJuiSGSqYi1itrMszMKfVL4ZAniRC7s7qiGznPAXmOFd
xFuB/Oc5wO4tYYHPSFC7s1WBG8VKchLkDVXhjAKD1BudOgM7MSLqzjUiFJd2NgEjLhgB2eAujxNF
/CDQ6caSWI1YLNa/KTSlTpdOaLfbETCKzsdxmz4zFMUxGr8w7A/oMMxaiSZo457uxA5cL3+7sqW3
PWbU7vucobdkDtvUoShq5KULSoed0mPdDyyeu1xvJtB1DE8N5hFrQW0RRsHuBWbPBY8DrCJReS/Z
y+mLWRp3MuJ0Mn5DFfx24Eoeh5u0A66dT/M5Ef61naJT3f+iJzRL+jlCinKtqEyJ2/zmwCZUEj0L
iNdmBSkri9lZX0eBbn6dnxY06e7rlZtq4iLLz/yb9grp6XZ2xklKAayMaF6HNNx9pIyqjoKxhGrz
nX7O8l84+ZJfxAmbJicQvdecje6LGIT7HMmneMpjn0OVLkdakv+NswiB0pfdCm8ymtbyK7DbCtZa
usqA/nOK7BaEiRYBb+7VZRhYIuQCr4ckwk66TEQJEP7ZAqeyot2IIahZu0NBM2R4FwC0a7mppuKs
G0UxPIR2IolNwZR2z+ExAC9o5N55nQjZjfjeFbFU1/dzQU+IrwNe/+L+sA0YuCwKeKO5sWR1QmBJ
xs4zWvGgx7MIUDGm6lqC5ECgZhgNvrDY/Mf3i4+OquVMz/iI5yrApM3mD8rzS2TJ+MvHUAS9ERNI
lhwLtvHo/1ytRFMxn22tCB6CpPo4kyynkLg9Vqk0aVQ/avf9dTrcVMfXizKzWt1LDKWkrxeb7djU
/PV0i+P5rBTbs+yPu5PeG2+/65UlBUvD1yEWHA2f10XZwpS7xoz0Bgb/YwrmUu0ldKvOiZpik9DQ
8/0oLSvRo3q4hNgKWUscsWOW0K0kxdFuwLcCUXsJRUmnYl8ud9AcBrw3dr/SnVAskardM3N+opmi
fhnHbEI/GE+A7m7HTWXNW05fx/b3Rqert79p93qQ7nC64dFXs4oBuuLsiI/zrhjDxWTLjUI+zw7J
0axpn8khuUpU/cumfKk+BBodH5gQW4LJoPfnmPOAxQrx5lv5UDfOmTugxemScHHAg8dKVjDrfb4n
KSYdK31PlO4k1lgz0CTz2Jwd6s10TEysG5feogE0JiofTuL7RCsVNdalgXxjmiSocApmAqA8liCe
MNmjq25SuYW0/V0o4Z5yuLg5jhoUtYVY/c7BwDa4azq1jpECo50oM3BP+lTIlVUPM1HPz3qj90Iu
dqbxdMAaw06F6v/HmXrgqAWXWGIw5lsL7pKG83Qe6a61SWO6bWsoq2UKjW0So0eb7fMRJQWTsgIA
svAl/GEshOn0Ky8einBF6Qj9KaQlKXdU99p4yDnHkdtLSeDryVEsFUCNeP0TpBTumoRcIkE/wR8C
z4EOklIM7yugpG6ciyufsA2sRRldQUZTptxBVUuOvnjyTBP/zvY/ytc4V/fTNr/OAxyr6IQMkMik
8dYby0K/LIHqNlAFUzcGh9lwqcXV0L81HtG6C0ZASq1vk5iLQLOJ9EGuIamyxMsSnNLRDX+/VgvP
lwqWHdmIVxTicSSb413ooPJVpYJ7+sp9XDtjhzbPTBUhN6ZcHtRzwGjIDuvKoF+6tQAIRrqDQdL/
n6nsFdEYFXDk0F0rFDtwhhtAq5Ao7+Ea2X/y/PQWWahD7oiu660uYz/2tl/2Q4yhpxf6bTaRJCaQ
NR9fRr+fuEwbYV4MSl9GFv+5+WvmPc+kKriedERUprqfXvNUuWpK7WizGBiCQ3jGIz5SV8SknWxG
h6vrbdIWreVLHY8a3KkuLkUmCn31ntcRLvyNA5Hjnp4aKnl2D3sNWob+xjnIojCQyp6tiaTZAQ8g
pGgYlEjVqeCbUlJ8thKPGSDaFhCAoBjXkVzmV6TDxMqwGGz7ZD4wtN+mcaUfoYujgeC3ZdwgohGX
ojYTIcURVwe9RPPS6SJR9kCuKJYLEXal2xYWuiZlImshdQx/cajYhdENhnN3rTdUPeG9jsH2OVG7
JA1QpocnThXtUxcX4PEl0vJFh73DZoQ3U436LwsCBFFTXx5hJyejLRHpe9nErlVoJhy8ZUZhq5GA
WdYCHGjpW1tNmb1hGbriZvPGnZzexJItHZD5ALNSrBh7G46gA6Zvic4/p0sH6BLcvb+dmd8BYR/G
iLk3qsKs2gzGc2Y6DzYtfzfsPcTAc8eattT6B9+gKpCdruaDAdwx36P7/5jkkkXSFeYUGcq4Rj4Y
IgUR3QjMuiIB5nqYaR/pWbfpHj8pCCoJ8IxKVZwFOAyTL0qHjeZPYhY8HSaMZTcZrPAu6KFf8xkS
Bq9FRd5y0ZPYENk3AQSmZyD2Z0tLrzOLsvArQh5Y6J7CynsPRy2BZzxd1XI9MzIb+HBzs2onl+P5
z7VNl1gavzvHqrsZj2Xqxjpa/bQtH9K0jhEJKJHG9oIA60cOa/oU7G8P8PyRS+2iE8awIELlqYCs
BgYhhx0+61OsYLNAginj12Sz28mWMU7q2F1HRGEaBysBUIOgauWGGjZlY9dAKZWie0tvr/ntV3Jm
CtsPuGdUCQRKcuVFqrGadJvCDlThzZq2AO2aQETDXk4Qe1VmsPOcdK/SRKuKPQgevUb10s5chTv7
uVWqN2vCxNb0HAfVHda3ndb6mWAPR2bH5RaoME5urNgkdWqYSp3SGizTeEilf5mhcuWdxtaxKsr5
xmu40qhh7wlvnc+7MHN+htgB3lHzzk6iOS+AgM2rhTKGSvUn2YM9rrKZQwJ9xNWf56uEpb1LAJBs
RRo2UiTrfm6SqKz2BGFdroQ9cyPyOVuumNzTNBq6iDqqppegBgL03ChKimntSMNlTd8teO+kNbVy
BCfcLBgyV6lC0ev0aRAvBI4IZPwSW/83dfQVPF8kTYjj9jqz50ZCccj/2gdn8777RiLs85anbv3Q
fiZvHtgLK7mFZNzW3FJeyVf1twGZtwEQSDEOShTotFaVhguXnKwc1idrMrTzRMxI7+seAy5J7aH4
PBENJ5/Iuael72MgTIsbSYwvYXsYFWXy0XYFcO5Bijf+DfD6jDEEu2zMtBy8YROVduD0/NTylrlL
a75au3CtxaOkM004c68dADk/+bPikILxVoMt4hICxE8KEu7hmU6XTzINwG6fc+HSl2jjxFoxDOqB
1IdjFZBVAkLKAg/m4bpooHC45DvHf1j2Fi0mirdSECzxhu8slgLVwAVsPCLvKINM+E49vq3dOyBS
8ZMneFyvRA++8U4Gn5cMhlbskxgnhTcLZscxzHvRUpxF8yOGRvxWsApEVRTJ9j3hd5BtBKeG2gVO
q4amtP124Ti1oa85GLU3sdJwWLTvQ4oJ9v+FqyIQt9L4+HIj9tGFsP1TArVMw5vErb8PdwCuHum/
6PoKMaA2FT4MtUyzmpn3jLJMfGfaUPwKPknV3YtkqHo8an97H5Ue61hPfiYtudju52ISE0ZSTmVX
X4zGQAlKn2FagfB4+p/P3qGlfm4iGJ0ygDTClWtyHZLRnSn6owyK1/00ZQUxqpf/rVtMkK8TACxr
e9gb/dEWNZXmqEgK6UlzUBrmdxTAsw2hU0sqwjk+1oTbUvHiouvEoSozwuP98Z1qjStYOukdBoaz
yQX2JWmMD5hiAGHYqXKAgsIKczYpPsUkwKHRb1+G3lptSdIQ1cENQM702jSLBSFXhbY2qbDUMWgM
xoQQEux3c9KXbDArJ+YviNBikyJQyeo3+nuOW/fAdfq3aKuMoCH4hOmLiUDDDr9UAeZLCX8FfBxI
RjdMWmg+JDM7tJQ+0/O77Qy/XAcGwG+CRAs3ck2zUgWcH0GXgis4LtmQkziKRnWDJHEX51VNLsJj
mYG4YiOuUlyM4oVL865wVpwHxd9TkzMJ3WQbpYYlwN3u34ADXRDJZ20/YQSzcUyyK3cRF44bo+vy
pml4tqPikc2sCkgS4IeZJNd+zS1PXSAHCzyIS4muVBWub5dAWqsuNv0/OtynEnSx0tGfg9YfOIM7
bX37ry2aD6GitDXMqRjme3KUtNZKqF+5/RPqma52tvBnSnc9UOBW1BEcUqAWyZ1+EEY3l5juT/fA
92Of22hwrtNCkBYdBVAv4/6Y+91tTGMqLGohc3kC17ucOmUrkFa8rDX2I9g0VDDhDSZpP8PasnHF
/sMDfY0mc5viE2ydMq3xWQGPh+IW5BlVLfk1r0mHD8imuKMjaDsrlsYCYtPD1vc5xXDg6v/QNI0+
shTl7zVfTnb1feNtfkHOcF4UOOhRaJ20XIkaL/lPPZR5f03p2GyZBIIkEbgAAiqvmPTA1RBQWHt0
siccVUS/SB6vcLEabctlXZoU/zVPzNfBIPzs+s3qodEUQg8S6+xI91ABWKl78SxwBZSIusZfM5t0
CayqIvLDJpRGVI943H+/32v0CZ1rnWrbL9wqTSPaKzr9l0GlMGPWE70SggeNtXJtSCtYJYMHDBRF
HF91K8SlWbokwkehqNM014Nm+gvetMPz+kJtmbfLBE9Cn0qgcNAXOlpVDoQeN9Sd7V3x+WSwIU24
rJ4vQeCw60qHAdMxXij/fENzhMmpCLkCBv306sT/oGwyfeeuiT2ydCPrknX0UEjnlUkkaBFrymYA
TgrslEqevZQ/iFh8BFx+s8QbQ/SlnWCHBTb8yvZ4DmOulyOj8khC83tp9+lHqqlIGJ/APU04bVm/
WsD0Gz20EIAdQ8WCUa1H2wuk3TVF2+Oykoz2fttmrmr3XN1HapKwUta+iF8AceCAJUi+0kAhk8Jb
aeDVzrs6OgPdptKtiSVFHTsc2sovA6AaZfXFAWU96Zyg/s8Iz5JWEL2XVdsBGQn7P5oVMdeGD93s
dMq9V1AqIZUrt5jUxnfY+B8uG9csfkIeqAuMWChOZrXM35Lh0r85t+OFbOZFm0oVMC9lAVkJf/P6
9HEEahb1xbAfZl3Eg7rc1kLl2RQ1giLmG634fsMZ0ghqMvJhRxMnVqS/gg1aXWCf2/MWkTbISMWj
uYhSoGifrhKH6O/VcGWVZO+DnTiIxrshfJk0SU9hD73Q/8JbIQngvKlwvPVdoymyBtw58HSsce1e
0Tj3ehOnEohKcEvPDhldmsB7wHoIew8inyqu57Fh5836uZDozQf3/nc/w7A2trKH7VdvC0RsaNhV
+Omt2LxiFoTSjBAUQfMUN+mVEjFvAQr0Ddsgoi8iKyJRoqzusCUxXnRurWzA+IWBUAzArB6JoBnI
2MYz1i7MAeYIjwcCBZTbq+G/hfssBFcz7SF2G+ww9PQEzkYjs3I2hlMf7OCFINT17MxcqROX1Z9A
Vd5qisZvK7V+1+JX1h2x3AI2E167KkurhOad6+xW2pzv57BbLQB1Oo2XgIujMyuXNhwHQfUm5fRu
0A7UHQX5dKxpWSGc5B/z59cC2vXdEy3aKw/xR79N7FTdWOq4j5XuNSy6o2OTnQsFej6Ywuk8SY4y
I8QX4xIGWbJL4W5oUw58CyHaE+/ZmkQomdRsJtZWYk4yUlJLqd0YFAWFu2yLSrHnCSrlCgQReYgX
ZSC9vZcLS4Tbq4q+40Qg6Ko36DqUQkslaZjxgqI0K/+/7sCN3Lu6LkEDnNuaP7wb6QNV4BHy35y/
x/yxpD3vUANLVFxu3sk6yOe9y5+j6lkcyrVUu9Vx1NCgrH4oHQkQB8mF9HWzbDtZyM7dOJdTkjJl
7/1vOGRUDqrFps1/zozjty8YtoJZylZa2mUWRn3/U6kqPTh8nAmPp0esMQVwB9GxtXzAbxA9oRFS
4w1pUZ3q2BGa2/e84vSjsv++wJqm5PVJDUplTxZS1pR1N2yYcxiU9AG4F0e0WVUn43MfUY7roYbh
v8XSVpD6HLqm3rTT+1Nuk/H2U6O0EtEMVQ0T3WQDb9EfD9TYBTsAjjqJL0whXP+/2VziM6mxAH0m
1FCrdJ6TAi8U16p2JISMXH9odhU32zHd3Ud+x0GwPm+R9W+gOUWWeJkWZwREI0PMRnFZ2OyO8jtk
9osNxdTdPlHm9BnQq1xxFaKIGCp89CcQLEBIK3+6jN6QWtul/kwOE1Z+CiHahVaQmGtT66uFAf2G
3MyFzddRv4I1FNHmpfavWtN3Man/dhVtAX69WVAsUj+Feecg2xpZzJQJ2ytlG0MA0i82GoU3cMSu
7W0sAxb90LVO4sDpzwVK96A00msLFbiC5bsaSCv6mePPhenh0iANuNiCFNkZUHKTPwyWTHxtT9UK
XuS+bZXE1PkvCx5emRc9T/uzftdqHIE0ys8sFOZxqQrHiaguZw0hipYsrHEhn0Ete7xFkcF+2yaN
MlHqVGBOFP8fb4qpyeEretYVL167oiU/Kr+e/7+PYiMwKj/4q6/r1StJMTSZWNqkgXagJ+un5Crq
JBmQ94BcGfb2vKYM/FOzq47a90ephBDP9F4defq8CZ2+6ZaBzGupHIXND7YGS1ZN1PewNZHxoLhN
bIO7BFp4M1wfwkQ1/JbkZfMj9yTSp9y5Ep0/rgJ4WQTWabIEaLDzB0KPqR0XGsBT3VSGzkp/zLsh
Z68TyCOW/X7nZCE/Pwp1fAgdkKJfE2pZUOeMNevxM4t1uFKTw8Svv1lTO2HDkK6yXj6S1M7947Ro
seiTOLjonB+lN8DbcXs7dczllXAFd5NZNYaVCco5Wmcp8GBG5edNQb/nIKPOvS2Nty5qSwtazURY
otTBdjbTXWP/u5qaQWfO7iyP+rxpsIGd/xE5mQYCtYbJr5AAG3jqU7UBor2R4O38EssGcqPJ/D22
KEcphVrU4pOaMrU/7V5jByNMm71r4ZiTkAxvb0chsdwQfeoFHHLB3RjF60Ec6QHNhtUQ2GxlRXOy
8rh4r0HaZloOk548TLA27MqHqqEySEA9bBzTT88e+DmVD0so1k5R7Qh5lKIjHE1//S+saTLq/G8L
6F4M8zPUDme1ku8XQroaJsObxSe7cj7rQyy7XYuS09AmLP2hkz0v36AVmJR7RGi3UNwG5lNKrsus
lIDbauNTBbGvNUnO5w/n17V2uBx9ivJDcP0vSWM+t23XKJiLeHU7QPNNUwTeLF70XntXK5AUHuDA
E7ithDbizS01TTe4BJWlkEI9HDG1aJOm6FoE3JUuTQu03rhoXeG3h6EgVyDEUrHnvOkn9PpdJSuO
qisY6yK0KZXGpiSDc5w5iptkqHtQ7R4htcjTb1g4tU11ClZ+askacj0GOWXuWLK/SECDtMrXvFju
b6lMO0RqPrGd2z5cLlngx2BpawqBz135t8+8gtXKjaH5Z7O+b+TDyPWH3pdbehl1LHrAajh0eO5a
Z7dr6gY8i2bG9IVPfxvYcpUwBg44J+OLtH8VewT6PSLmpXFu7Ed31ryPNdlYsrL21AJZVdPEFxr3
IQWOA/YHyi7dzb9UAo+d9HOej7/H12mFTEb9wfXpYnxnnLSMvYjnH8YQlZrsYQoRVlf737gTNGhj
eLeiFpsYSCmW86CaJ+JgUVqmvQvWxyuFirDNq4OBqct9vGoQrgrWPFoCYM3/MJK8wuWOrBEIrQE6
uym6UNHlicNUhHkNVrCWFoDOMlwIj45Ox7tsSQbVV2S7syGZifiBREKWFfHzErpIJv+4CrbHzW7D
/NU4jBaQ6hrjnrbBLdThMSVuKBN6KoaUgrNgvveiaD4fu1nq/60vDcJ5s0S3Yt/0x04zu9b3o0mv
J6mkOyI3jyIIurcX/utDHYYv/661POKPDXVGjSpqlzlyRIGwKZ/TX8xtg85MupJ0Arwp6MthXUKC
rtBHlrUWpG574pXGeZcgMcD8HkdU0AvwottT7wrI/26WNqHzSFUi90oUWHiJw9H2sXujhECysXUr
tVZqs/ZPAb7uMkx4CuIxBrV/VtOZjyKLiQnk0UxG7VHHhiu7yZDyVg5HWy+oKz4lf3J/C/jnzHx/
s/Wmrd159v505+k3RFIqDA4xtdABYMq6h62kaF9WOl8rdngF/pLs4wFYqqKNgoTUjPujslyH6Mgt
87sQBPGyab0gpB2QXCoi65CFnqezQE7NxW9Zbn/ZT510/yEnoxeFcsTiU9MtuqtghscjES0d4dZZ
ZBqIP4u1Gr6LbHbqUBnuX0WS35UvUJn87xLbutUOVdLF4sTOU3uVkbhDKJkhfWgvryi0V6MNsUif
WQPl5B/LRU7+2+RciPgz8+qasTB2Z32PJPy727/58XWUt+ipm5iPkW/7lscCg9JNn01+dcswVZJ3
ESNyxZMm1c/dNZQ9EKWtM1Patg/9VZZpj9vxWtWrl7lTm7sPTFIjIxAzNceoXYNgNPpRZV0aB5pF
JP7kmWL3tgVVhqwPGqbcPxikUM8jnwV0l7zQsCYh6JQjgovvxIvBUajL9EOfXcfzZPnxIsKmeE0g
JskzV2sxTWMo4PjK/exE2RMeI0QtPBuREOklQww7MXM235aL9684Jn24EIek05o8FzwbUN01LpQ4
GCKkZ1ESRbjcC2aUA8OJpDafITOErihWlmPFU+uetWdgx3P33IdklLb0Atgu1bquZ+cO0Y65lMax
fZcjC793BZ9e/77GxA5nNhe1vgMmadzJldEJN2zNL5bDRx+lMfKbl6Em4/1zeVuqHvqvYAlRlAWH
jApNP2i3Peoc1+Duq5NmZsUGdxqO+seGqcjW9+Det6rJINVPWL7o1M5A7CXxJUOhnXI30Kc7oH4V
tVnspGlvd3uiPzX6YWMyhRpIvkGFE0jwnsGPrlKe83FtkYMEcpcgNjSLVLxPPkcqF50zaPNyNTmO
aCEB6Zm1h3Q9/3nE0Najbr+cFDP2IsWsWitd9uzLFQAke7MhWwifFnRsMg/IzRiwnQol9bsNJtWp
QFlkNMTrSVbRXhciAid0Nj2UOVhWz/LuvS46zwrY0LyZhZgKt57pq7Bng+RYchX2BrGc+nKA+qG+
BPJXFRIPy324sQQQduQrbwHXTAMbhuiXn4Gv8oSQ/YD9R50JBNEwHR0J998qoWQW5LCtfLspCjCN
zEcBPVLc29FYpE81sKW/2r0fVccFpyuAfuK8rVl+iKvSnl81uL8VCNpnFXbYX+cPOLHIRFtSIsxG
maLt5inQuSlrJPYk7sX/aJHJro/ghbBQ37OxCTOzFAV+HTOxlav6SEwCvDU8p6HfySSrCFTqufzS
wCrijJnbB6TyAVwwgirHBchhQ6mQZSVBvJkkL/IjwXoClHlw6DsKik4BB78Ty0e5kDOdFsrRyvlO
8SiXKSFY8cSAFm3alJ8CJLY/9oNi0LWRezwh0UKDitvHw6BYH/1YaLR9UNXf1NaYPSzpPNPw99AH
EdMDqoQG9uxYSwglGD5JzGqPeehfExZ3he5rPJIQzRRni3YWFlR8xzWkjHA3tYSwfJAQUQ2piHOd
Z6frex6VXEm/FUF0OTA8gz76wsHQP3NWmYWmhDMJ803CsAtj2gdRheTFwYuCiNlznDbOQq/P9EuO
Iy5HAC2QdkXATY3MoJeXwInZLy51AZi8KHoPYuTsD0D5UEodSTDQNM/DJsdzHsWYNzBv0LhLef/H
NLw3X+GECurXKASIwB5DdF/2pTrpZ0KanKlUX1Ben3opPY+GnIH+/kjrZ1nFhsd+b2n/aVtm2VpG
CsTgyNLt2xlijbtG0FXmseaX4BfLIgQoKokjzC3y7tPTrU3QO7mkHRy0S8hN+dDrO42EiI6xLvPl
GNSRZ432qOQHnPc+t+f2d2F39JEEHEap/LPWvcK6NAZ7rwKx9e0CIiil39/l8QfiaE+jIDo5TCms
3bbd5+fju3CAZw1pYaNgdOq6nswwwcTa4daZFEXYOZyKBdxdUeln7I1UfQodazZNTnAFz7g7UnbW
F0kBkmoLLtgbztaalMiL3Tp2fFwD3qQ/6fGq1U+dJZJlqMpzQ/M+vPrQvpfBf/422AF0peTh+xiR
//006Gk6YBSZpzEIoZjlT4uN00CmOshkvFwjewjSBPIqiPSSlItzuoVZIyqKNOoy1JRXfJEUg13a
WaRhOwEXg2+FwKtl4HsTbY5kgH/OK2SR/eyf/X/1ak70bJfXKED00/87wkHkTiAWCrwoOt/ujfKp
IgU6GDVD01QwbMwxuNBGuwwp0GwyDGGa+ZX9+Hc8Xln3kQ7VsQ332sEVJjVE7VC/8VksBtl+7UdA
3rcrj8FMms5NPkF00Mo8kHlrqTGHi+b4g4BxjbMMyzyrxO/dpwGWKeFf40m0EUuDx0jL3BYikUNb
v9TSNJxTiXZIGsR17N+klWM05qUhmN469HCFSZ7ILiH2DDlEZPZ66qJjrGIj3YayRN7xDBOJeV9h
i7ThuW5YEIzX50Ld4DOT3DBtng+RbPZBuvcYcINB440HDcW1iTwZaBrGE8SjA3mx8GgmLAe7zaaQ
LZl6lZgZuZHs39p656yiJixaP+blcPcRxLG3+91mOKiYQ1/9Vs4N6LFstRViI1A0ceON3dg95NNG
zQebDuS98DOJyiXWkZJFiFYf986O8x6T5ujbpvddXj2Ji+qut41P9tjQoWWl5LzRMxuMrEYY6v2b
lq4Xl5e7BgqD0ILm9oMPOxvhsWim1Gd0/ieFbCrIpnC4/tTBKafyFZDFgdSMlG+CH5phK1rmuuzK
wa8X/MjJwGVfNPQewK56pFWJ0crxEying9kaWrQdnpt4MuDTb4iaO+ABCo2p60COdZb+VSSOe2hk
NqCqzEDts3aiVCyZppk6JKHq58lIUM5R23uXCgJZ27mGJrGeCfV7jDQCR8tx3qr2rnkR2hBSviC7
oYPDwsx+eY/zSDO58t7a7+w/z0AIceiKl1tlsFgMcKcW+voQRwMP7qlUp9RhD25SxqkqQC2ep9iN
eC69geAaAQQjufXe3iJZeCvz9Q4aDV1vO3v+TvrBZzrNOTBzJsFUX6UfxPR/mbx0bMVggIhFWk4J
ev/LMwfSU7sTCkFTz1MBhDYwRLnisoXRIKjGNxQ/k84g3bYfnqL45prZebKZkOF8G9whwoTsgNMr
fZAAE4dyB1I6ArIjtYWVI07VMPd1l7ofcL3bHErmw657P7M6fc7lJqmoObcZOjsVC/It9tYJsGOz
gZzg4g+fdC2BWzCPuvWGG6RwbPDY5Pv807hlGh27KGe1FrzIediDFdqFEQgf+ONu1JSjD2v30jdw
zv11UmOglTo9nqmvaF35nIK6aslgPy7KzkbjbfUafBt/bN+z/85zA+/Nftkw0371fHCiiqH/4ZEa
rbnxRBnLYVkH6OFLKXB+V7g+CNKu0Pic+3ur/los6vI7c1iNoUSRY6yZCJyPamABYSjPMkjN2ZEy
P5qi9AzC54Lnui7fnRZfq5Oc3MHqT2UfcnJI76azo5GZrQ8R7JCakHvRwsjLvBdCGIi0uJg0dc/f
iFt8VVJhtD9fQlYcPSQLUUcaaSgqQ6Nj+fYHRxTzMpHJRxF2xQ7ghDLLXCewwog//nndZbHPwhnu
xhf7mw9Q0dRCUy3HL4kWxEVP+pwdvd0cVlnlp8bmcfEqts2QPLN2aebVEZTVl2Wndxtb03mEdQlo
YSbgkPwk3DEmgEZh3xyzcIH3kaHVn9IksRH2708dhi0NbnUHBC/dcy+f3/Qw95hafUMVrn7lKSX5
4w5Id/n++Ih4qwagKaQ2w3TGUnQDN9mj2fRvjYLomRU9NQOyMVmbXJyjGrjMqyagHvJBePbtjqmp
8ESgc6MV57f1Sp/1Q4AWKy0qg544IO8d4/sQ1WjWEpRFC8xamG9OvlemTTJTpwdnZVTiG3L5+TNk
0f4tULmpr/rthpduG6fN1g35OV2Tx6A9yQr46dvNA4ZGsd6TKU3NZw59tLCk9WnTBPYGMhSFyS+g
jAiDCNQU4R2GoCD1xcXammFn7xJH01TgvGyKBrJo5IM583KfA7NAy0uzSPCtXnEdoKU6txLOVlGr
x+PAmBHS2PFSImh0SHUfKZDtTTWM+Qw/fIl0UxeI9OmZ7USTrOFj3hNsHT1GPoxibiVFwOjC8XnV
q5EZSmX9CCD44SSe841o7CjxpScAGbxEh/hU1gAtzqidAUCHBOrgBIOFiakEGa6qT7gBHF3vg5iC
MaMtOtZ5+5VDnN6cRCsaJJAASkK+Y+NU0eTKJhVkfI9cs2KUUld7EurHUvbhws1pTemOUyAYn53A
CEmgnKIHUOQtwjVF2F0hGEmEPkdm41OyUHZV5QJAJ0ZhARx7D5drNul7//P5+cHZRPqMLz6+IdWd
IMYdD2/41Wg6rXRmqMGfcVvBuwpvqRIB+84KlRXMJgwtMnUnyfxv2Jls4zNcHOb7zdk6Xu3emibD
nf5BnkmFgZx66EI2tTRmWmdA8kGkuhgZrzcSz3VhIfwZ9/2fR6d5MZu+P8AdWJH2dJC65o9mt3xQ
O9FRLW6+yFjqpAtebXd1AO1XKDWMCPY0VTkRX0bH9zf0XSNMlkVJFLnxsqN6+rwELRxWEtnAuBcv
JTaCkDOYOR2dlbU8Cip6zU/KjUhR7O3Fw56mz+i3beDK+MoIyUXXFE5BetviStZtnBiKGwtOyIwq
7Mu+Z63vCVid0v79eS+6OWWgehXz53Xhd4beK8ZY1DIGhaJCzXjn+TNtgmQ7pFmE34PB2gWgBw2J
PNNCB5vvmYKWgNMb1a5F8Z2aRt3aAKNtxG7Y70H+yl25aY26cE7g3l7mw7zLMk2BIcvjwwxIhtDw
F7fO8Pz61vGmAR9AoZ+erPULaNIpmhf+gUFh2xs+YPYITuPrCeb67TEdvEi8nztw21nHltEt9bpd
gDwxt0dYNo/NOe7MeZ3penLhPvUE38WDdjuDUyd+PoJcG23a6sL0VSUvHToKy/PIwjAzX3kDGP1D
wy1q6f+qQ9cGNZy7JaJvTqDLRyEFLhYVNWAaAnzsje0DRPba/H6a+ybcrhumBfly/TDNH9/C8Grw
erSTc2OEza6+R+7FV9aNaURrmajkllSUNxJLY4N+R/2jsKQeU0ECJu8M0iGa/NbKZutzNkFqCwH+
SdzBw4MP23bH7gNMiHojcIfjZUkTybRM9mgOVjpfV1Y6dD1LhnI1Q434k566bgG84kkPCInQA/JA
GUtaZmvoT4cM/qLbSNd7grUzM42XB3VxJbJq2aQ87FUhBWlRGA8Ma5ByDXR4+wj4du1dnMJxA3RT
2w1d4CbHqaP8fXUaGoykuVvP3CwnNEioqd0t0Wj6hkt7ZorPhqfYoIlV1VsgO/5bwIk3HmuxD9yK
6TIAF7xObgDsCfilHL4HFi0LDEdlYx0GtT0vLDbFhQugYwqHx7lMi+4gU1amHOf2uka7O339kpRw
aIIWVeHTYEVq6d8h5PWZdcmP2JRue24o/aFcmDxi3ND2iYoJgblkJ4VvfK1KdAUgfCZKQU+wRxSN
9nDfdh7KR+JKdEvBhAr3vou8d23+iIfybjUJquMApZTuufGwijftnqNcJ63N3+1v3bRqtEoe2tNR
FZ3g1BTWncfhyQ+GTU0/4s0dVg2Av2Evxgf0Tam5gJnuGp7WAXMrB76ZuWyDIoIGHHfsfPLcLNLN
qU0ZCQJUo/k8Gf79pNj5OMhkw3D564Olm9lU4Rb0fk4W+SIHDWV+X8UUupWU+jTTDqBMh1nV25e7
otrBsQJiyEP1a4PU1YPAzZUaS+WZkuvaiHXkMnOq1N0xvJKGoKNCULMuMn/th6yXEOQ0fDJ1keTm
AbNDAvViEOvaHy73FWat/M68o0NEne1RaXCOHLdEcia3juCmUkkRsbKBx5JmebaWVKYnrT4Yk/sM
moenCkOjVB7/dWPuG/p5vqu/KKaW+fONp2J8iep6UD3NGdLG07xrrTRerDNQ87kfUjYDJnJhB3Y+
/ofLPCir+rSfIVVl6aVpiv93Sqiq4y8ajAnwDchgK5Iwg7WKG9zsODYk9r96lQ7whM1Cr7zpyMMp
f/oEmnH2E8KV9LzRYoe3Ne/uoqBc1sMP0LHX97GPYkdd2sJ1gACDM8HEvbZ4hSQ3OhFj33lNflvi
9bo5cq4wqUXy/p6KupIquvaos5FJsHsZz+03Mr6nsniBp9Bl85ljyzkgMxMjGXwIblrXIGjPQLVh
pb3H3UdCKPXtad846Mwpnb9TzAISHBtVRhjNwT13A/9TAPzu7PKy4BkcdX1O3bJGe3ovwSPH2awe
S+8dY0zaOs6tsu1gsmt/MG1xXnStn43qYbe+YFgUVCkUbDcGZQD/f0feWKp2ffOPwxq377ZhGCiH
CuCyqR8oVYjnzByppY/34e1/b9ETNHaK2Mn0zsj5XGGk+g060IWuVyJ+kL1o5RrFOQxJNeqmxx2R
aqR5kQdH8KFYJOD/R8anjPy+Qnh1hGIZAwn9lQpoR9YpfuTt84ohH2C+KbV2ocWcjXbc7WExn8c6
8wtgcBlwZfK3pg7EY+PaBsrTOxBH0vdJG9r+53ZnJKoyy2ESTvEOxG5KMH8s75299LvS0CkWgoie
30+705qMP3PoLpYHPPGQfASVPWiDeZj3J7t+FR7y0osOKjhUizC+TFw140r6iPYPLB34FSH6sS2v
xLwHA9zKW5sexm+yWxgBw7ZVHiUuZZjRTIZF6wJ8+zQn29LF0DZJHslNz+nMUlHt3HwCQGJUEVCn
dBOEL5jO94NFRpNnAbmWuHcfgw5dNicVDLtMg9nvfixUD8WalDbDU/28YyaI7XTBBwx4QPL0G4G5
ejkF3vp/6Eno/K/PMe4H8qoo1Ltveu1kaPHH0xJGTDG/sHnfv8GdTuYPKBs5OUEVBNRyRS902yy2
Z/ytjl5O6Y7aMTF4g+tCPeHHyKwSPGfE2dlDdZA2oFPGucVRbDbWz2V5ncbvhPLqL+8WiFoXAks4
SD6cx1yrsyV6qHpsoMWtYs30UV9joaYw26NMUEFibdj84xd4bMwECwO1CuNgQyK+9SSj2dOLs/w7
9YnVcWz8ElAqaPfHIrLSfW5WmIy71VrExIw5HE7toYFR80v8EreQg9Oe/gCHSJUDc7GDnKAf761l
ekOm++nRiUaJMw4/sXsd53EchnRqE1pjeOLXHlw0yiItEZRt8XBaOB+NSGv49iNGf7P03aa7wX/s
ApXb5VkieNy/Tx57Tn2lEi6wVOvovi90f3ENFik80gsHrAmnd5e3Gcxrty1KT4/OSDXuRgc93U3c
pN57jpTMprs3PoeCSrK4RkioPGlmD1vv3VzMuJ2a+Q0nZ3JV9xEMaFbYSxDKwtMDn/ZTyrC2WWxN
OUvBmHKsNPgxe3bpsuZHpVDEFbZ5ZkC09iCPmJTqRWF6c3nFfO62ear9zhSaJJyEcEsLhXKsDiCD
XHvM4oti5eDR8fPtLrncjAF154xNkh8P9ZIrfBEv3sgekO8BFn4Y7LvuU6MuT6yorUM+z2l89c3/
qaisiWkgv7VU825XBrw1pKg2Km9teu5qg36+vkGnd56hUBrj6pEHXzwSNfwgGmCv0gb785cDkOvc
75wtO/Nu/ie6oSc5GWCAjZD14aUlMs/8brHJIE9VaPT6sxTmZ5ob+qtANwR0hTe0hYmF34xtlz0d
tXWDEnSDQD/ZYnHFRgw317cNQICMn710ukkLRz4oJFNGoRYFk9eHZNfPaPxche95wWvaqRd9LlXI
P4eo2eWRg49NyF+IfVG9B4D6IiJo6vyVdBS1TDk7rHR4oQVMssuJrJy5gz7FRFQWSG1aZ71Ksd/L
hQhCd8CuNsA5myyPfDpeIuILjc+qO7OgLofdQ/+Zff4w9p/fvY5/CqUXvz78oEfFqiBcIKyLFQRz
ersU2Es5p/OH0lJnVR3bF77abJIuXgAj+o2++AgSgEJBhU8RhROKHa1gPDyHtFme94pQCSHEr71I
3c0iPm8Wm8ni8AVZeW6mEzNsQ2MKF02nbJhaYh0Bwol1PXkPhvj8k4EiznP4cGSqiyW5ydhbF7L4
TDid4fX8eG9w8w1HvFx0zHUpKY2N9uTzutEozBWOSZxC/r8+W0qlo7owoyHnjOZ9Q7EFDhhPAOY9
YCRfCP8I/RvhQsbYDUO4uAaoX1SF7HLxPt+CnA4f7VG4cM3zy03eHTwG9rzuUfSjae2Oex9bybty
HttM++5KWNm4CcaOtCHUnk6IuLq4hDXMBWhJTA2OebXUS6UbjOgm7XPTV8i6WEha4gwnBqOXXbGi
vtbNuaI+QSS+8m9fLHKFoy2mG8tzwmdS9xuXeZjNdhQS4hlp2RzSzLLuemD04ep0OsrbksRzI9YC
BnhuiNNtKBvSTYcswioBepaJM7UEBwbuDFlSkSjET7qN4YlKfhj7f5ZHjhi+1Kg8twCzxXUcFyE2
VPforXtKFdffzAo7a4YlwNyjGH4Qeth8QbMfH5MnmOXwD/jvb031rjq2RT5tK2Se5h3MeYsq/bIF
3jXnSmeBvgikZd0LTyKElx/PXYOwj4+OmMMMHjSxdBpqiIiHq7jRMDAIrP28t9yVFDrThGRAKw9Z
OFiRWATJnzOIy0LBCv6SEe9DEmUCH3YkcCHjsvKjyQACNduGzJb9yRXby8VHe7oejoXyXfwWotPi
AgqmPjOHMTJSF18Q0xojxR0hAyAefnpZBuYel+6RuT86xYOZaYK9hnrzq643yFUSW7GQv47Z+xWh
DxG2oCMZAIdr+8QG1RgylNfW5niVDSl+atHCVnILrFRfzLeETNn+bjKwlKDWVvIRKlKadh/FaalW
v3kYbYQdAaJcDx/yPzd4T/C3h0Z200nVMdaiZhaZXf9Mb00t56yf21HS3/MdoMXVtNaoEcKP3b/5
GCHZPfLPg+qFQQBjmAP0/YC/LsNX8D9HG1aPyb0wCrCDV1fWMZL0rHp457s5JGJ6tSf/uOQzVrD4
iJY4hRM2wqJOduJ06hmUaM57eb/iMtZKnoAbYzy7aRFkKVHlLAT7R4j1R/rftYIyHwBMh5HyFvN/
pwYzziAVZm/0lw3uF/HUtIAGvjfulGSithCzB0DmP/9TvqCGxeFad9x4Ykg/3iWJKw8ijrdaYOXl
+SjfTF0U7mTaVztufOllaYusxUQmCIW92A3ZLuuWbNwNTjTZZKXDEWQHFaMhLw479zghs72CGZxJ
Op67rtgAYV7/lDhmMraBnD82HvuTvq2WOocqoFpVhe7dGl8mNGi7/b5O6uECJmB3uDNBbpkzrzoU
kizkSTNYmjAksgAG+6aO1S01vxsfDCUP3fNKtP8MErxVSsDAymXLn7toZT7+OcFPLl1ZiOU2bMtx
ujCrmVHJ/NXg7XkX232DOxz4vpaKTJm4Vit3mCBlRJhj6Y9ILeOFWk2QNr5pJCGcGi9lK/HnfTmz
G3cO7nR9UXIyLEFRh/HTLEISVsubddvLJ7UMVvybX4MVTB+rPBpuonn1Py/64hrkcRcyqfbRxN2v
OuI//9ZISkC+wbRaObhTMJis2oN4+97OAyreg9w5TQQ63jxR/H7zyrFBi3mpvpLcWAQhizy2gW0u
PlsyKYWKr3I3JRxEFWIpEUz+NTE5mQ05KARqXI/F7E13C3woVAIw1JTFdq8CKAfhS5X0pH5DJ76t
UicMJ6j3jduAXGFZwxGDK+01y6XU/sNnEoWRTFdm/uiMzSAC1jYjUMJ3anYFqx+2OS6L3MaOclDk
h3levhnxFNOCNDQ6MqJZDXloll65NgaqLV7elPog+syPm9ISVHxVP5bOiy2Ay/WcT/8VR+jZWjgc
BBC9Vuw1EaZHGhsD8KAnYcJFRRdBfZldKMnEkdWRWJ22pONn9+tZxaYcC4PONiFlEHJNSycNQL66
Kw3CM5IfjizAQ7WJlcK6nFoZ5OhNx7YfTjGva+xV5JW8WvqMocMzYejNVDE5SH6EJSKnAptVnja2
7YYybsr29F2irF5dE3EvyygqJDVId0qFcNiEs3CN9xB2HYFGjxXW8HFaiT89z8QYP99lbsMe8U3G
4f02DMRnz8IERNQY3oBrS7qNPqtXhPQ2mqEHTq2n1nZ9juI//xFBS8SK324X6itgK8qEf/YANOcy
mJB+RFGGMpSaFjkPKK2WxsFLEQaxK1YLAlSbPQY//5GLt9J83uGGX9XIpv2yAswkx+fRwvBIKc7p
VMeYiv5b2+nEc7YJ8PTkB5WWjHGhiWx9UL38eCZXPMaDoenUAGqXGo+yx/NGI5j7ZGw7XmrsdgAo
lB3Qk8xBl6/q4dHFiqOxd9hI5Zi64MG7Ee20qr2jOXg0R/vP7pqX9mkfOKfQF3tdGK0DEOJZGE4c
x0jYZ4aH9lp8JQeKuSrfdol+tRFiPOnXqGQcsK7DL69i4+rtj/JtZWRTc01EmpqCzRA38l6yhpkY
G3rPamCOwkUveX5jlNo0ZHuVb1ASTdQkK9kwqNvISLLiKs6DB7QWIy+tC+Jdw6x449epGqunhr1N
sYf1kdtC6cw8bEy+xCk5vmA85UIqOC9CtSTvAxRwICQXWRGwqf+i3fQs1X19hjSffWPAp8fJ11ik
5Esx+Wcd0zIjEzDaXmw1Zj2VThiwZXFI2TxC93xaeSxRMR7/FFWxj/98lo8zqks+0PNgMM067Sq/
jzU6AiAzGN9wn7IXqkwhIaQ+jNmFNmMbfYo4Q3cHBqBMymKF49HteXGYQxfPlhbvruJZBlOEmamS
dRVkojQGhwyKGuptZAjBkfSx8vhwNKM7i/fVxW2J2dBVmW4ZM1doy8r3/LP3f/yw1Khha44rirTu
10D4aLXG0hdTyvb8Yf13sZNU6zu62a6O9u3bgcdkTpNgsIRjIlLY3u5Qs2iqGJHdsYArx4hHbGPL
z1JQlweoJYXC5Fynyoc3FwSKmtg6NQiWxdDVoJChgj9Zv3qfN3HtRUo3fFAfet54CFC2LgqwmCZM
qDoWXIo4eePjPMeIZtOHbI2v0/l+LM4pQFEOMUg1KCbHPFEV76Dz2CwWNUvaLQWX32DC/X7OZmu9
KTMWsy+SQnlOsEn6yzmmsg9W9yE3Td2EGXkCO6Op5A9gNgGV7VcSvKQG78PCM+uN4JiA8nlON1cZ
TsDk2Bw11YXyf1rzHO2qWeKZU+Wf4hxLg/LvIdj7YJbsLwwZWlbYNifu+qZ/McH8FaEB/5bj+L5L
jOEAsMjNGAeKqb50HHb3yGozNKcD9YvbJI7GMMnsSKXWlerXpmUBua5sFntE4EYQ5DOuYPIVd2r7
odM4HKNolouY3Hsoe+f8Tc5qHanB/drsFMwYpp6yVoCQuunTCH9OuOoQMTqTzxECPGTxOUFa5CeS
/XjV9pSCelGnwugfiJC/nl6a+Qj7IpytT+cbCCMJ94LTw6F861iop3rAfenSjxccZTX9qyP+zhlX
sXHj5G8MvZe/KZXEUs7RflHDW1fZkV+12/h5BLhCC+or9oPPoPcfes9FyfZhYFJK1l90n4V9jwIB
Uv7uJjtsNMWGQwl0bHfs2nrqW72DI9/T5TwKMIJ1XAWgRUjxl/d18hGjDJBDYLippAjThLHRhSXC
QOWyLT+BZiuPSx76jFxQ7wZYErUwhmpBIF5G713/MzH2rQM73j6hyrvIQslMIHtNaECwQEvEikTI
yWn3fuCATG9UgI7B4oko/EsfObgdhMBI3dlBoL6BKSaT2sSOoKX05s3XzPMSBlmKR6fu0CHsUwhw
AN32z6HHwvpH031JYNb/dwsWeYFI28cyidm9oy5ecIPEfQJxcRgnzQHMkxWP50+sjrPJy0m/9clM
KzEVOkyR3IPZYnwsVVs/JH3YbCarK3ibtSywX6sWVy1ThyH2CwD5wKvPWdQh0n6tbep/Nko5gD2F
2jOsbe+e8FX0zAMhC1l2LtVrqYoY/SuMBPsnsmkJ/i2lVMn4Zs0Lmgbcquvldb+0aBkAGSMjJGYB
P769sSgOf6inbnmCOisX+Ach03ZQYDaa2K3EHV9KjkXFaW/R+l+ruuaP5N6uhBl0EhhGFWZpRXAE
WEjqiLbdzdUlQBGRwQmFpt9AJoHFqe6ZVIR2nWeNKpSGYZEZDlFkYh2hOnpZJ2mkbEhlOVOZ1on2
Iuim+O9DuOpDbe1hMXWlD0BHkOUx9rZw3CYEYbCAgzTa4YTqOEDgqk8zqV9jJvOCJCkENZ4Sf02k
5OGwIpLpF+3eP+70B6kVBzDVk+bUah/hiQ8dp9u19WZcwctbTsytCrRxPQ+OIOQ810IhUH24oJZD
xQMA4AzX2jRb8ltiW6M0UWO12b7O2jv7q7l/hLWQwtRqwYEaTWNBwN4m1mjJeISJTaSa2mt2okpf
cmCVNTLXxKjYC+YT31R04Edkdf67AnQ2/W51hjTacvdn+BcDS6EhvCLw2WUAVqFI59Nz8s04VOEc
zOJdEDQeUDCJU9wI5WxFAQBli42vBTlisFIaoAOM9qx9OyXYVQMOc9LRQ5s8VoTZfjUzGQoV7pQ3
o9zn0HTSUu9K2d5gEfoigmX68hS7PfahhX7F9Kjzs+wn3SgpISR3WQfO578NpjqhLeXTK6Z3jnXO
bimbyFGY7KEzh7OQ3ifx2Yuy5C+2vWFwF13pSzjEIdwMR8A4FEe9F6DwpAS/+QHeD/AaEhJGQMpU
NdYBKv7HP1EEhDtZJtxYyM454kmu+JEbxu9Qxtj+gbh2GrihtRestdQAHugR+P4OZUcZNNTxB6BN
ubYsSh5m/lnTSjkKAhpmYgiqgzXHBy1fPJt2wyPbXGNjltXOhBSlKROorw56UxDY0mDFle6vxPkC
phhUObe1ONDC8eje+X0pmeLZPMhx8JROsFxCDeTyKk7kIgoMY5u486zgrhZUILs1lQMm+zpaLMOX
0Zg6pLzQuSr74PgcnpW77QdkvvvpR5X53Ape/JvhMyXO+9T5AtdhOQ74GCItkc3VeRUmkgo2P6BG
WR+t/laxjyuWzDECiY3vz+6nAIbx29dkWEB1ai4Mw7LlBBDxY9bYtqKn8sh1Zj4EjKVNbUS5yRKh
wGvF2rA68HWpkUyZ/y7bD5nJGoZhicqgJu5WQxkKE6ifoZxVhJFVEqpKGAbnFdq6DP9O8uYxO6O/
RVXYkQeRBoAKccRWyjXVoDcH9IMvZm64sAyZCmph7d+R5m9LKfae1QzGqvjLi++ZOVip+BdrL5iV
Y/FG7qa0a1YS8WhkDiQK91F3z2mvALrIcl31Ailsq3I1H/I3/VYZ+0z4NVz3L4Ii30pQEI1REa0j
e+m/Bfd69F9zYhXrJsFTo0+DQLiCh0MKjmVTAU1gA+XRgNYhR8Di0rbSaJRS1bPJl//SILHo7ziE
utLLDrm0Dw7OyoWEMH/gKZRWm6BqowNfeYN12rETMJTHunzamSJAytSdF4hbv5SYm4oGLd2AYYsN
Z035LSCHS/lA1ptxybrozQVAY5U0yKp+44xfjfXP4iyhqRcgCOGb9TN8n70THfGvZ18xLs4VQ3Xl
mejuJkCR1ooDvTCd3W/yFfBJtDLxVgcfPxkjoAsIZEB1QFd04O9sYbDo0wnuMOwpkmv5MfOPvuhi
ZVcZyqv1p/mwvBHFS6BkeMjwWcLjlGxv0ixy/aN+6HQe5pUHh3TO5hg1lxmEHvVdyqxFkFp9i6Ie
48VTzb7DfE0iwPve0dhj7gUqZgWyB9FR1GvW2bJXFGAvPbme0uELd/4e0EiEU5In8mJFeL1U0jMz
ja226gVhoJw9v97EVX8Wv/pH/27iuCUuTM3fFpg+7jJXYFngtDg8WvLr4AjqkmhKBB2VBb/WyLri
1iQa0kC5ThXl6irer99RJDvq2RMzlbMR7pC9cmJ6yJ/Zz9jYPsBikPr7jS+e/eZE5Xuk2lbN32B+
r9I43WqB4M2//xfzPowChk0JSAmGKkqjmqKwyWLa6wwugGA1JLIRn3REmJ8ReYiGdSPlO+d3wP7/
uh8bOcegbwzXyucHkxRr2IhWiTfDSYm6Q4RGw5zocsl2zUSoYLhxesbRUPob6jTqa2ZYZAMV/Azx
JA6hm5R5fXmbnwjpF5cQ2zl5mxkH8IsX1iT+NSJuDHqvPPV9grYYNx1hUsg+5WIRic97raw3YqKn
3yF0HS6lMJWzmLQL68JNznVPrDvEbBRF6wAvGFH0ESe4giuE8/n9QfzPxtmp1inJmXbo3c0xyHYY
vmSG6Bz8rSarXe8v/Tz7eIEb06a5sWqcCkIlT040TABRfZtpgfSMJ7lDfaTTYX/UnQsCyx1hB9sd
WwXl+cVY1T3qmEVcPb5FLPr2twT9xMnKQWtDj3jHxbmTuoBp3uYk67nJ2IzdlPUX2e/sYWrvZu2c
hv6mV66Lf6b/MS8AMnfP7MuR0nnaP/9kdclZ9OPy9ijACeIY1BNI+2oN6dWn01uwydKWGuFfaKdM
NlSp/SLXt0lawhBJvOqCrAfCtmUyFATaaxx+buvw/toxUBwdOaurl+fi/Tx8MG+JHAOrKXZ1C/lK
MrDttKCn1fm4g+ThKQiZllaPw+g6flM+gfMDZuv2qOzSB5Gre77l/PHOaRsATZ5M8plx+IB3+TY2
9DHYpfrrhiuVBzRqAR5FhQH3drSbtrClfkpCkx9pw2yYtlOEOLZ3wXSgVzp+EEUHAUQvHNaF5RGe
PP7l0e1oWYB02WiFi4pQTyH16CMkrImkd+pAWegitlyj5WaY4sY4dFLTfQfpirT7rKKNoC1YfO6H
RDqKwlXcvqZlA0x9L6NffB4q1mWaNhPt69/noic+SyiEnI/Uyg1z1WvBGlGOy0Kqb/MlDaLGieEZ
r4D08MMm3ojVTWCrMMW28pWFkCpNe3XphFlyeSUSGVGFEMdQA2VePkbW06epeyW4PQqPASRwNuek
6Npc5qSLWC9Ry34WAS0bhlCmu+zmWmj2y9Qb63ATZ5QBo/K6joIC90kjmB72G8ZpSbngHSOCxs/x
WKIPQON4Y0QRo8wiTR01BJa01yFNxza8nZ+OejcOlnelA5KYYtLKdDd+/t1gwywf5DQO0jE47osU
M21XxYZ+U2L4bQcytG7qOqJ4E0WVfsb8DjYl8vH68KqmEyTHqqbCJylQgAlam2HNQTw9ukQyzGg9
y6ahEi+NZuFcpykcLvZr3s5eSlIWRWhuGGodJBYmiBcDIu3OkT8JzZh6/jxt3FREEFHWwNWLpSlv
k1uIK8TKAmfAB9x8h33XBkOoEq05TndokRP1ls6P6epDvczJ4RpOpdZvBFDYGiY/HnWMIkwP4PP3
A3h2cpDIKPaoIK1jG6SNrDtrtbULihyTQtzCbX/rbBhVpALYzW5zdUitUhQWnYVEjYlB/zx12MoF
GntnH68kzwVL62tQdMk/UMQDIsGgcdCc6s9ok271niaVBauDN70mIg0ItzkSh9OIji9QbqrpBMNK
uT131PV1bEodZIP8stQjX4DaTWlpIHCGyZUnJKeHweRxNS1yGkMCwsZ+pioe/EOLiX3GD+8QVOHj
+DY6cN3Mj8UjfOC6JpVgZzrzlH00ApW4nULZ0kFUqgFomgSkRia5WXpuA2SxICJrYhnvByk5j6fL
gU1thGspjmMPEiIddGDjE4ixgTclJGcmRlI7+y0k5bzs17siRhuaPyFGiyf8fYbqNUMcg2TrpvbE
cfMOr5xBMSF2wOOVMtlRWIhhTFhc9xCdUfbz5q6LTKbRE4M+ZgB1wMXpfv0FHX1Gsyb2Zozls7hh
Oo2/CBWbZvxKfw+4YZpEMRTx/7KIOznG63yniuD1dVQVHZgY87Vl3qgS19c0cXuzcTsJIPf+bqHq
JYEZ/IWGoeZc4WjoisTfS0oY8F13F5Bk3PDtE4kykLIT1H5GVg4FErAHW18JBmRjHCQYoiXA6G/d
ZEpPnG3J0Nh/cpdJAZBnQk+0alq3MM/ZIApggNeu6ZtQgY3S1YDG7uq7hEusHdvF2cmKKAI3Q2Wj
8Y8ZHRXU/inFiTrfmDJ2a6+/i9y7cDLBQ02U689ICR+rVXFDYz4/uUQwVUdjHfXy+vH1xoA3sf0v
XO27nwY1jXiW5MyXAHQU3Hf9eDqENtDpN/Ayg7Pm+8M4kKejLCsToIXzcrBooTMaug7uVQ5qAwLF
M61qTCJy8QCqkCFcnhNtaPwTh6WZ77mYcRGimh8DuDDvhwR34l6umDMRhjBkkicfFebsss5OgHPY
ZBp4O7JKmFGSsSVfzL0ruvKu0nhkja4jrW7OXGnpOT2KOGUl9kPnFC5DUg36XbJ8MLCAif8irtlG
qG8rg/l+ZQg3DLthEYRCLlJoO1Ffizpi3iEmwZxkFaT8ic7kGYqI1YbFw/LbJ9wR6CVzIVap2yVk
7lGoSHfyY9hbMkWPVw7mlk/7jWt43eq+UrkHDwFXpl7HCAWb4JfQVvN3vBkIrei+2kR9wt/FOgRy
7p9dSwCoCN1ojsLpo3oHL888VAUhghfHteCzBiqLIvERActPJUrD8TPjqRwyEq5wa+D5AvxYNljq
UFr7ng1XVQomWuDGvLoD4XYEFOVZuzSt5XXhwz7BcYvWydFjzmnBPP0xvt3CS2kKkVvkYrNSndrr
oJYOoShOy8p8PCZoU8ESgBJYO4rfXp/BABfE5Jd1k3rSNO7PyYenRlAh1x5jiLxr5NFng2wevH9O
UqZZtunR0wzSJPXVAJPeleC+ZeTiPdxr/JdxjCZAi3bfhT3AvSeftP9db6HZBxkv2m8XhS1HCjPb
N3x8la09SijI5GDgFWhN/w7Gok6V4IuLYCEBneUjZYuqG0+0lkAdwKr76+OMaepN9eOYh+M5KkJ5
WZx8c0apkcZy+GtciEBwZK3173Ni2Hzxks0s0rOckiHd6QtIRoqXZYjF2KVnDOTWCj9s+VzuZ57E
dFQLibt9QMcUZYRPdO3qlAIXT2v7iNCOrZW1fMsrFUvcz7u9e61EJsc+LgBC8KS4Do0KmVS8kFXu
I38C11VECVWR/kD68spQfuJq+LPzv2wF7OLvhbOjpCVTxVy8eZ99N45D8NDdlNy8QNKAUkHEL+aF
zCM0GdlHVYmZ/6pHoxJqPXzpfWt0bANlrTHe6AqFozeV+kdq3/4PZIxsEFmwklLPCFvSuSrxjQNp
s/bHTaDqRVaRF9kSErLn/fb4vTUERujyQrguii2+NUlAQ8tFSJotyyXkt2IKLo9p3jg4k/f3D+Nr
snHbrCKF1xclj0hq0QR54Ysrm4KpJ6uIxSG51to3hYjt1EO7dljydOJDpnljb6QryOZbOF3A4eRO
ObyeF+mRL4EpdXLx4QxJ66qnnhOA6wq2+4n8vYhoJi966ZBwOyf3wC86ibhihLBsVM5XnTC/8zAR
SHqP1wB2D4da0JmVT9IVjp5LaH0X2VpyD+cVkQgBucB2udnaIZ5iwz7z9lpoEOIem2Vd+/QGHsTi
ROpOf87Ts+4X3c1FcCMBIfoIuQd1CDS/yR/Q4gfMVPVuIr1BZNmlu6vAhzEIoY/K+thFNVL96de1
XmrgYjfUiQM//bTdcHdvl4DwNA/1FIchK9Ez7j+11Yhh0wPl/pPVKhu4k/Tz4iRrtdK7MmN2OuMQ
ZHMJLOVay8BWnptFBkVau5Lw4GxUG/onBJ8tptnoJypsokVx5z4WZyS53IhHPoO8GX6dATE0luwC
lZpD9QQdZ3WiAyRPcp30Nwv9/GfVmSdp/PNQMkgpaAKrYqe+yQOiyGrO4ryQHkwZfO/kLsG94Dqf
eL95G35niELtKHnP1cziH6fddUcqorAW0sPKCktrlUIfnq8zfV+uhbuewGAurXAUFzgei58Ire3+
jfBXoYwBeeeG0v0OfNBjgocgmldZUOsDvK+JDKcOnb92elQQdiXWrvr9jZTHP3Ducmu6hBSJPR1P
o560sYd92s1AOUwqWNMo8DT+AjkOmDgGwe4fwp+qZCWPi2oWXQP+IEzQ1s8s3pySE8FqT2nEPL+x
+5Cy475KkSUdbn3wsWoxSxP5vPOOTD+Nb/jCl1xJGGmsrNVfg2hxrjPsVIF4u3GFmYdoHOqHubRP
u7Qj9h+Ay8KBybJJDtrcuucRu46XbRrR4oa4cOY8AMVdQAI+XDc91x8mg36O4llNDahhROliv1LJ
2UB64p2tmBQV/Yi5q3yemy97ky2w40VK9uhpxyohbuNZ8sRdVz9tGZzl5o4sPFhTWqDNasTdGa8k
9SMXvG4STelE4WDQNLtj5on/u4Pq4+sfXwY/baci6FOL/8cGJvgMfpaCT1IIONMjJ1oK8iujua+P
dS9n4GoV1qyJibZUq4q7CEoB/1ZwOdh5PhG90cWv2CDaIFJrTB2XjXs+1pHpjF7HcCDw1PWmiwLQ
hGcCCzaSCmZb4h/vMgMik+bgqjdXuctJZrxAXAx0JWfQa9Z+lWuPivUiSmx8EKHZwJaQ5+aN+T7e
nBv3A1nAKS+C5+IV4TrinDvzL8NFspLysaBWZeSQPnoWVDMiIAoGDUfRkzqsUEOCPIM8L3gAZyqi
PXWSYh+B52IRM6xxmPIlLjTYjdeURbwp6KaJGoPbGbQNrervKQDP5IoCrdKLqZyh26hw+b1uTyJq
Ii7zX4PNvtSyc+9KmT1tYKQH4/452jccYnkOiwV6SAVr121D2dmuxNUJ5LwRTqJe+OMGooUnHOWr
Rp0R7R9N1YiQP+DqRxR7VSCdDwuvuJcrHv2gkXzCOAaRMIrPR5cC0OozmuficjenRmwaiMlMuPKa
yZgbbjph+GIfYHwzvoaZInQ9SdYhce/K1taddUoP4z0ZHjpRtw5A/VZhLzyyVnmcE8UsRRwfK/mw
FyEM1SlahuBz+/vckAYgBVo5IpQqlHUEqt+oD+apr+1NnzK5lKo7PEUHJOx11EOvJOfBKqr0btFN
QysvnqPTcJvehzaqrQrBYdy4oVd1Ba2eMjRBIDx6ZBYtp0/dGL45ZuT3KyZ8IBGDFdK+aBjr+QMR
1nTXp99XM6HzjWGkZAuXch+xzoa6GLDyP+jfxmuay5nIE1SroxoSw13bxrbASWCYHqjxAJ7A/byO
KhEFh+GSCOzp5M23YPrpOnGJ4P4qIql3JqIcgr31GVUwdYsZn4ERWTMDe/Au6Lz/HB6Gw1U/6lGw
vHBGVvcJxnqnpdH9yr0bNw3mBD3kJno7+x1k83ErcuL1MN5BiVotHkPotPNvzkquMtq2zaMh7Tiv
OjSBZl4ojhWWbOEVugXpykI6s4OxQuAZjpJMB0qt4h/0CXDen87GNwupcJF3I5wvLBoTThXlg8uT
PThM7CGcOWHUNwNCmkqD+SvsP7O9lO+Oq2J2O7/cFslgEXkHSmz6GDkmXPf0dmELvoEq9GPspvy2
LqptzqR1CUVVUl1XxjKGMvXo36zg+ET0q2vmhN4q3NoxPKy/GKg1LqXbuLS4NUqbS9rMIsAdsucs
hMURD7v25r+f0ZZR0FB4CA1K7vM4Q+OimLQC+N5MkbROxHoHpFpA0/6B8bdqUZSzXkOyPdawDLkI
Xk41f5ZwMNH6oFVKcnML921u4xvm6zU7CxUORnJLAoXjICTodJ0Ca55DB4HU5M2CRUh7ZzzOhaIF
AmH5m2LwCQwG31yttne3Zu6n1FNBQINJ+bgpwlDglWXbtC3dXaEhX/HqsLiOqHjgj2ViNtGuxMnE
MtE4d4zAKIqifeBD9QOVuFziV/h+mfsi8kuX3OXHC5YaOOu0/0YIeSf8N6cg81AF6W59GfdPwG97
V6J4pgHTJJiROZd06tzua51ekNaiLAzXifU0zs9aQ5plKNYAarbxXk0seNfsy4Rf1IDg3afSz122
MdyItb2+7yKeudUD726m+FOTC1fmQJBYp5TUlinyuX9j/ETGANMGQGQLUuVhCTu++qNP/WLoHKT4
65Jlc4oFWF5DzdswOXaEb5q1rNpSsuK0VqTYb/KnR1KdDSTluSlEzomaSRrU2YtIAwg4pCY3EmnR
yQ6XUcsMEi7oHeSgApMMNx1aj11IBuuj3ZML5giboyc2hXhoOZY2GuYzv8A0g1CPbhDYMQwBcNaR
trsfHGGGRtGEPeup0veQDPk5bHoiQtO50ygGnyFf8P3YjBPNa/+3+Od6gOyNE3/dgjA6ZxRLLKJE
wytfopHHHTtyCtFPotJUkOG40G5j3xzS6wu5ktdyhBL5p6gj7nNIbkTk+V2GiG6+WAGioHgBQ4eL
dvo9hvQVl596PzMOx/V0yVfKvaSxhnEHsNhN74KzgghfxS9En2n8yfQ454Xp3j2+GiQ1QGpON52l
jBxSUD5kiHwZvDFQjdr0PH9S8UacId7e2vWyY1e3WG73dqphQ5cb1fZ0sOKchUDXWkl7O8JRvwg3
fJDueB05jwwLS4ktrkFuCgBn1lDSaOFV4L16B5zI0wvynNk9Hp+m6xpbYlQHPuPtJjXPDZ8ejNJB
X7Me089nneF6hzAHfUMIIPZ+EKo5yBHSyzSuOE2/jmN23YJwmfrlTBh15mB/jZq8qCZdOGkshTIe
/wMu+KQ3d1piCgSlil0oztrZhRP+PcjWvhG1hMEkvYEtPhqIzwrFrmkKqnfDy4bWjO0Ygzoz/o6D
OH9e13+ui0CMaCltsTElAeVNAr+VZPfSrk6YdWIJz4JHW6QKHzKdg8t6+2GUmbvD6xLbSieEQWyS
ZET3mmGJTsoc3VUkkayGrkeRWqiZgE3VGRVzRlG1SlAS7Hw0t7jGe+n6Mrh89GuPGEa0otls03Hz
JXH5FlXAzOkcPs+BaAMQnikwTwuaTsg7jGff64YNWDdOzzb1QafEmbVvl7MmB3MAw0x8DjDE6k4/
e6ciL7YfR3VeUsn+OG8JZ0ZV0IjswczzVqtx3eAI9tpQt0yFf/D+LC7lJM3LDNtgonD8jSatLKOg
HNtLCCBUXhkR9+/3k0Ghu1FUhEka/AhIcjZS9Ivn6WL3I8qxknrokkFDdljSluGDVmbZaAu6rWzB
hSFn41z8n24s8e8ZAG1oMiO6/CCUaxBpZzgPduHmbBh8Kd4uGJG2FNmJOQ0Gt0chZkkuObWGBu9C
Gj8wE2fPkvMQ5K0gLZ1HAxY5QCVEN5BLU+pnWaCotnKm5a98lZhGRpOqYrN9v0qRWF4vUJwMWZ6H
gshlb9zKaQoWkictikKqo4+dJAi7nQzVxEf0BZkpz+rMcqFiD4GvDYsDly/eE25GoW1RBdwV6Om8
uM/3CzUtoXhPTH7CFLYmFwXzBkR2ImYxmqrZNWbNp94uu+zqDw27gKciBMgGfmVPivEmLDM0ksL7
Niz3U0H1zxvm2Eqf+aRHi02i704AErU3yjGvqZr8NNj0TL7RRPqFM52iSX8Y49YzTfrnvMNkvSOy
e87GK3kf8EAFaO9HT+xzkCk2s8WQsHTIWM+LW20ngSAZHcjdlOSrtO4RItzpiMPL98F0ZO8d9wGW
zQeM1jGx5mHAi5YOAgDAehJ+1IfSIdwssTMftKZH4j0Din4e2PTm2fueqiHKWP1A9bLyi/5anDS3
rX+eyRFxZGqq/QZqNeFWK7mGNII5IqBPZ48dig5wPMVvrxfl4Lm+Ow0+kP7PW87u6C11ln7mP/Og
mPhrErrk0OERjCqctujVRzOaVAW3KqpvMbBgc21+IOi8qEf3wMoC4u+tJt8BDi3cA75B2vxRUnJH
2gc+QO0lrjs2wnL8fwPUZQooHObi/bXt22cwFCHMHtd8O5dnBNvmMI9vCO128zIFjyxj1ZKrShwZ
iW2hFGcNjcwTtkxtodbgRzc7sGyKVxHMhKjVL0td+vA/J2Iw9Wi9DW6s3SIlVtUL3bg1he2EXBQQ
d0hI5fxBWdOGCIjR1KAHAqtY7m3zX2IkT/difaA0duY4mBifv93CAUT5j2MDVNQrmDAjsQm9nrKS
E5X1K7YkHM8W3SmgR/2+ilQUFbylpgkzL4uxC6R5Mbl6IW9yx3zKw/iCaSp4RDnYiRVyB/CvorlG
Pk6ZeWN8xf4T7LW14x/Oaiv79n2Xdn0s3kyZipf1MFaDIOxTWZJGRaN192LgxGsA4bOM2b8ycqqe
cXVkYCdBg7XgVnBNmbO//WKOW+RGV2Jpz4Nl1HBmnQ+C3NbP3p7KFfrh0Z7DW8NNLCSwzcvZEyhj
nFMA6+RDKhfKbcKVv3AUOuEZXASJqtj2gp6a+F+oJbdoL89Fr3JH0DyjJ2fySGOy7qo6IAr4luyr
3gqeyaiH2iZIjrSlQ/3cF/jQWo6Dlcw9cn7FrMpWDWXFj6WZyqlRi7BS+OobZ8wB4RGnvZfdW+rp
0tTpVCspIF/8s+inDEGKEaGgGpZ3cRUIHjN1hK+MZThmhnZPpnlF7Zwqhul8PxSuzXVwUlDgOEhr
KEkFR5bLnP4YFGDxbcKMgvs4umcPnl3gLiMWQLvPFwAzQwiGL6x8/CuBTQHXGqahBcggRErzAhK9
Zv19etcmdiH5IXwLEAD7gpILxIF5xWiT68Kd660UejhcNyaMzo6rjzhS2dh0hCz2utViKoS8846V
ke9z8O9wlEQCWvLuTMulGKRzWcq2XQU9iIwqIypy6sgqx1luq+3Ay19BKqO4SgotBiz9kJ2tMBa5
t0OHBV8BgY/uUm7ghkg7wVT0Wvg1olYZQrcjJRz3pEweLV7fKdN9DQIDbsfEsjwB4Q+u1nIa+YJF
uKhFMFAERRnuP+oGC/2KG90TBhKr9asiBfkZCU6Bv7pwBifLTYdLuodECyUihRpKHwK1x6xamBGB
oZ26xg4EUEsO+T8tJ7+sOKsq06cf6amMopmTdhxCT13YCYSseJCFlC6hzrpil0BzfkAwJKGm+/Oz
nUdxipMs5OcQrA7tCrhkxSkv+zfjBULCRU3AF07FX2QmUeUdBneoPIWNc/NTtrjPr8nayN84vRTR
G+LOBTy2fXCx4GFrt8hXUA9okzS7Qn6/z4+HFPf5PVhB1cXt4bkJGb/UsxkkQ3C0Y2Y1a/o3l6Zh
MwTYBR95qSSxgBau3uPEw07096wW1FH5v1dDkrERemUFasymZXVLDrhfc/ox2Jth+GRn0YxoDsKx
GMfkqVuQ+YqbwTqNbheixc+tVY6R9UjTevPdw5vLSTqr0BFl7QbFplBCsm67VJtc12Y0mycsH+F/
asKCTfYp+WGT2FmcV8+UNCiAsBjyuqMo0szlFL4IxrwzBo9OjV70eRp61HWkAw5y8a0pshZnSlr3
HbfItD3qyP7vMol4b3jdHptZVA9OZ/ZXSD+Ho2RZx1eN+4je9TcTtbSQBBJKFRqwovsMeZleys8Q
ej+vSiaMaKLfzof+9OsIZkF5acqejuSpZU3q8etK9y0YfB36SZbuLMDKTrIBN20aszRwZk4ddnHL
7rmkwo52PCijcsg/ZWfLZ0fj4PZCrmSfwlJIjkKykthcQf2PPcZFFHQVg1xSwVgBnE2c/0l0tDnj
/glTGafrX6DGN2EDju0AQSRytI9N2Q713rI78wwJjNro+f0JgPCcSUpHIaPq2Otn7pgtWnZXYlvS
Rrs8yzz8try4ER6QgBaFkD9uS5UXchQgC+WjaeXib/tAuv2xNWOnmDfi1i2K49q7/djATMMfoJUq
LvzYt0RT3nd6mGyBbv6AVtEoe/I8YpT8G8cdjMJG7Ha+TM5hgNjMXc6i8XJF6vDUIjqHEp0R7gV6
9qKpHpo67KkwSu7F2DxQAqtfqRk4Op8fdigM2Y1zuQTfBml55n/52o8fBdjTkGj6lxhuaCPeAQmu
9a8dEaCMAURxXxIhszY0n1f1YKOdlIUAuN85Py/nevuz/o9yWin/J8KPfV0vdD8sbdPpLpyHDYjp
GQkEsM31JBwojuS3CVqbobYbWUKbXxd4tta/5u+v5C+YZdp2fSUVZ73IolAg8mGeJulUNNaxf2sU
SEnIA4g1nSbQX5shR8Ytq08csaZW3tG3sdHGoo1A9uRCOOSZXCBUCcJ+qG4UuIMaveQvl9hA5qbP
H1bsPRP7M/MGJVC2eEJ5gvScIdMnfwqaePR9+PuP4XeHmdpfoeXfCB4MNXBrgTPA8DTifL7z3Pdx
CtZawT4YPztK52bgWkZcWngiIv4IHSTDFC6NQslvWB+oG1Hb0l6KBF3CZB1QcX+eyB3fX5rnewK3
m1h6SyPPySkP2ZxHWj/L1r0irrbbOi78VM5yEGRwn7MTGzxsU7xEwisb67eBmYVkuiReEEO1Uy02
BSQN8iw60Fn57tmkKpbExPM5g4vB71ya5J7+bdGzxXJGEw0FWzwj7NnImeu48lxGWAhUED5hMjS2
xYZnQmrP5GfWdblLIJzAv7HEqTWSro/dSTMRM73X0jzrTV+nENBamA6msFy4H+Hk0J2j0/oIKk/U
m44EiS/SyWP0fpVLPKeZXYZOJYkCHcMfDMpKwLcUzDtHSUuAi5MSeKYjnlQZEtw0/fTc4CqH740r
0DBpso4UEbuciBEvmjeph0NpqXHP13T/YO/Tx5QOe4Xl8Fzpr7p1Eu1loUs1jrog+3uWgdBOUOK3
l8b4L5ZjWzvQapfMpEMs5UnsIRZjfPprzxCBoyeWRnGCbfvU339JumeLBebEGJEBAUDV4i/XYtjA
paRWCkuaLl1VBMEgZaPBf5/CqHvGyh0cs7NKM85Eh+95JPG+aOUrnVWrNSfI2ZzMa+mXkHFLONwL
j1Iq+SDjATwySC0kji1XtV2thDf5kMGU2kHFpPXlr+tiYcStVLlqd/H5n/GS+tHv8dRJ+lm9f6sm
UV+FahZO7VXQ9GnGaf1iQKNQ73k0fjGnU1EdRx+P6wTXXC5Hr85bN3lD9qFhiSKRgFrKWoLx1DCg
dTJQm0WJh1P92Sfpy7DTq5XemMu7F2wsXy+MkyVaN3kc4hIsDt6megwKuzDl4HAosaz5SpEqh8wA
JeklbMEWqwRMO9Fax4x4yeEBbK1HPMKJJ8avmNk7/EFzNR0csAw8MzVwdiMQ0kRErkebHTIsAfqO
pQ6dnyUY2n/eFCLEYE24/aAreknswoHV6QgbZ84wkL8IMmGSjBpytvUT0AL7FqofRIEA08YsSJgv
z+dikGp/BAmYpQgG7RFsQbmChFWNL4/+1zMl9vm6QLzSvEJr45VDp+AERGO2hOeXN2NTdUbfurcT
8aZ6ZFiV7/zcXQCdSRDOmFYAfBqWPk5EVj+TUUSEduo3h275a2g1Wf+dRlIb2OxE3+4Cx8DBysWC
3wTz0S3Zl9IkqlXuP7SnYy9VXuM58XdVy4FCnVEOiXz3hDouPLikLgHjZUnc4ftva4Td1rAk2I0d
+OfkbnlhiEuZEUPRgoPwbb/vwvO3fCxz+tyy0hmQ/meLfVVaPexQ3ANTdoDFkeR2b/LpnlDhKQea
rtlQYadjIPIRFTPAer9+qvKjZ8U/lYVYu+cL3OkJVOpDCNQooNXsQSQr3gxqW8myFyg2pfGfCrg0
3bfF7D4k6LTkWZGeQEqSZbxItbvQs3ba4EJLIMEvxbjmo0V/7Rn4rGk2fb3xjcqvnzMn2bGeYf65
dvKCfDjY+JdYvGbWsnEw/HiSKNZZ6SQ3vaTcRvjxWdIsE7GoxAWxyikaDo4dncy8ERgIqiJ0tQoS
RHFlfumHu0S+9zsQplT8/2OqUvEmwZBgEYbV6w0iwbNEcwSnMV3xpaEDik66t59mDUwIGnW4y+yr
wuCTe6jIvteGUCB8S1oOv3IOHZhq1zu1YD8/z/qvAlzer2a4wS40qeYtSwZ+37or7E16rogpPdGT
7lzg6kkyIwhNJA6qBo0GoR11aA6H2dKtLWKOtxfq2gMtVdrL75McnVG98xaSSfwCCYgc3yli2t5q
ba0Z8tSMt2FDG6oCw/bzkbC1QWHgFWFQvAu8bggDbQE7xaOJsPu6BqO1Cbe+BECobnu2kzEaEOli
uToaRwc/FyOJcCqFJ9+ao5viUAFGymLTfhycx0oHHQ91ght5NWWwEIVWtY8c8rodP54TIiKjl9ZT
a8c57DuBIEgALIdVQ7/Rh5ygbYOrkLOkFCZi5EWBUhI8WZRkgx1zR90E21T45ISiGGfD1KLTOGSJ
YobPVOuGA3/QHj3hxYq5BaZiUilWLpgHtjuhY+t7YaJBswGLgJrBKsOZ0dqlfc2ckEItsMr1GHXb
+H0qkoVJdXTx5RBKRcgnuqH4BNkNtLvT3AoUlXN4No5mTfHvVI795lc+/ecGtGED7ay3i44j0ZZQ
rwvrsWcRwem/83WDbjX95pzEAPLYuGM/pqWAte1ifd2yl8YTMR8fzMZehkQH+UvcXSO5NOdzUxFx
0D7X6+/DAUW09jab3sVhzLBwuf5Ej/FtAl+UgJcUWkijbfGETo1dlU4uWqsocdDOZOLPy0bUocyH
W49c2Eby2CycuKuP2kRl2e+PufslX/42jOp0y/F83BlN4lTTj7gGiGTrpKzIkXXWzYv3o61Tbahu
TiiLSULQ1AOoVFmi0nSdAvsqsjgJUOBu/XzXRI4PuUQ+JA3phn9arzBtybtCsG97t1IZpHDGhv0G
cAquVcRVVfFA/0sMgOnU30GRG7CWNxQmcSnyO2YWap9KilHAu+2mTUEoBNIUyYVafa9vzi0VWdyP
5pZIBvJKIS3PnGZgWIOXqywpdXSDZjXb8mZgAehDJ5abiZr5T8PLDC44SrTfoW0Wa32WETFd1yJp
tahAjaK83kvveNp+0ePO+CJsCvphrm09Rzqc0dK2HTegwGdL7r3qqqTnHMr7exC/dKsSZC+7bFYX
PxPT9v1fYEORMEImo/ymiV4dssv8aqmQz8fFuznXFEL+4C/fbWDgO9Qk0SE+fQLgJo09SI7LS50M
AG2kqQQIvdyhR8nlp6KauoaIKgeFAQEAF6pS/0Y15vJC7mvbOZQL0g5Hfa41xzN6InRMuAtgLic8
58iKi/SvR8mDsysLwj574Q/ecwUGb1wV1lufagtBhkgp1vtIX1hEJG8FKPCt6Q2kh5mA6qEeci9R
lCyTnbPxLS/JSeaRcm3DfZ1nI7xoA6eiySkeBGDHicK9uwPKuKqRNrQokFckqe6h0By9KL1RKR/2
Eq7gvTVcvHfdeYdYD6Fob9pRv66ifHGKVuYnZtT7a/W+wYBnvcoAJLlE5EregYdqPcBRXcehKXxD
iS1oDkjSgBZb4Mh2dIK5gk1Pg0i/d7xiqlSHqGPCbXoC2kJQR/jubu+tqdKoK6DLY+01ZM/xN+3D
tkn4KZzj+OYAKRC2U+uljDxc6SUhSH9v4fjjwJAAPkMGvsEyJwJRQVKtbC3TAQe4QE+foi2mLNGq
z8dsGQIxkdylesCEAKg1QnvNCh1aIUUoFAIwatAkhtyjhO5ngICM99pcaoZjxSYJEjhTS8y3wQhq
kUBA91QylqMxTLGDBXCMMtDEXwoX0Q5l6pUOjKam5ezFFo54RjtbYigxWg9HxQVWNA1m74AF7P9j
t/Ure8De2t0YWP/Kpxtgrvg7ldbU8YHbbzDVHxe2qpK+29iC4o8Wfsl2i7FyM3kSKSLS9cjEkNf2
BuQaSyvJ9O87wUFDKhckfGXOV0vvCT+hyu9BTzefhdrgDczDud88fZhcxPd7FFESkL9qrSHi+EvA
rPhohdTuD1P1TH8QF6R+4mgwZUBrpzaIi9xsXxXdaz/X2apLBMryw1Coe66ZLaW5WbQ7cROLcAXJ
ul5S1papSsskDynIJuSHbRIg98RY67nn2c7CnurbOE+bsgmFL1bjE8CAt3XxUA4Zo47/eUCkXtjA
58qmbJJxb3zLANrXCHzBZVWgrUR9WUooWStGusXK5CWDLonk8bEeyD4EhStDRhJBCTADcs9Otz8b
hbB7fwYsQdZuMyWPbWAGVOR78sfswSFiJEhRkzMxe16uh/U04jxIlCBAMdOXjzyazIu40+SBIwRo
qtAtFom0xAw1A4iW4aYsNdL2XVaULocuna54asgrF9mRVsQWTJJiFpF4Oe5GmXbo7Sa+Qdqvsbr2
MB7aM27zPFx7rzs7o8IBGOUjNt67YBJELS4+x1aLgRfaLgMI1KM9anlCHkkNKRJ4f3R75kf8dtmT
X1UElObaM6sXs4iH240ElIsj4WicSwYCGlHOPW4lyfwvtw4r3JSXZxl2CNQT+lHVN0IeASsQFhR3
wSuMcDqPwsnJ6ZDCEfczOKMOTmM8Lr9Q1n0Re+RyXMgrnK3OxSY46e6temXT5L4UPPnqwUT1YcSr
XpfzMoRkGLVvtIPgS5RjKUPlgU0xajjWc6k86mAsCHONsvcI0V7mbAXqLpmCcQFeaFP9wPs8rN1g
TlJEN+a1ZkFxhVEOAHINr8VkJc4Yr7d2PDvDuD1xHBjF5n8UxwQiE+VvLeMFy6cfbGOCMfLs5sHB
+pCjBNZbyzzHJzB3NGOx5EzCg23KTiByE48o3F6loF1FX2Hsg5e22fOvte3v8mTLavRmDJOSPhiY
tlxW2xGm0++VAqXVghVkVlQODYG+GDB69uw4+7Ykm7qmynOZgTnCSAV2ZeOqjbw8Qe59cYiBt/kF
lpj3cIanf/ywzf9Lswf3wq9mk2kqjOcO3xWCTZekogMPDky1gfP/rwDJbtgqiaptrR+cWf+7yzLK
4VaT78cq5xXI2dpyUAxiufj2GWKpZ0HntIDePOmjcV6J76iALuszMl2B8skbZjZu3AmrdeSD9gsj
oyrd6Y6JnL6nz9z1NesZhf+qaMlXsq1+BWPdlcoo6YfjROLZqMKxS8DTmLxqwPOblun5Omfh+Ooq
Q3XE1hU3/I1qP2eQcxZcXJ95WgtcfSj8D7yWzLMvvTiz7O7gm6R2r4XkzykLWt+OKOLq6CAO/8mu
QGJVQzNheYsiOQ2Qf1vOiQzUFRK4ZObMuSiEJxSCYVsFi4Aw3xe3952pYsNHIM6tuWX6wdiJBtRA
j920YdJWOv/qrDRXa+FYt3FB/isEP2ThK2+pxF6Yr1NkRKtxWYCJ3CyoN88DISugLimeWjUfXSoQ
Jj9F996QnvdnYP07tK0s0g5aDB2pEePmon0fdu/lraXcj6LuUh2eRN8i47v0DLGVH+5I24cByUe7
ZHFmq+qiK2+cA9ImOMXppiw5vozNpJGrzDpOjXhSOH48gEwRwNAB1erQG9oKCJP97OwT0tk5arZp
KGwmcv4ABWxyRWrruFswmsSPCHnbgBd6/ZW14Xe/D7AniQ6xbdsnuJBFzh+KCmGvgYWlh+4ak/8H
Doh/vjXNTEapT9wT9aqqlKccqHvl/6mnXIObFFbJcIGUkfYZteTfSC5dhB4dd3YK0xTTWsVdnuKj
OsezVlZq9XHSl/7CMJl6EYsNf1fuKx5/WCVybh0EBu1QI9hm8dGI/sEjonx4VaiDOvju88N7ap1m
fEGq7b4ffRVziKNcIOweNd/NhEvevTpD0Sz+v33DaOMh0vJtt6zd778+BYj0qFaJiCxLuVpuVTwT
n6LEAFagGMpfJdslbFDHRF91+6tkgPjjH53zPC1rIv5Lob3TDWw6bMwPqzp4B1UlRRazNvJj2O9m
3E2c3KXe2601t43/rKLHszNiyxitFlMRv5BL5t1V/7xNkuZQXTfpz3KU5WiMz7PC/l7AgWEBo5ZX
1Twpb5KcG83MrB2aXDKgZBjW2LNRlgPTNPgBuu+neqEKkRPyWlqs3k+hyLCQXSbP5Wi1hPUmcdFn
1dOXydDkvX15XfAvral97pyQ0de9aor7zhuumbE2Tc8xGv/gS9HwQGYKWREJyELwpXZIlYppQOae
SfxfakUnEcrk026Q1MAHGCqMk8vJTuM81k2N6V1JugHT52DmVdPrZyPDn7n5JF2JvwavTu1cWMro
UOeO51P6rXcpRAi0V9UmrLOz606wwgA/ZlTwjhOMzV6X7GuynQljS/IjTkL5X/PekuMIGhS5qCJf
Q9g6K8hB8C24LeZMFcsA9kY9J6XXoI9rIUxGT3WuTyPJcsWMyTBgx7N6WW+ANFJzHwPytZKnR+ky
a+K9EhXhF+TYr8/D0x7OWQzYMt3vqto5J/T9Hr6JE5l1U+F576YZmxsuMM/gtk9hAqZ1qJnqq+Ft
Y3X+4SOb8OlFpe6PhZ5mV+leT7ZU5HedcGgXU0KI2xmTdma1/RWVS2yxThQx6E4+SBaCB8qETygh
PLEZLQGg+DRuC1+Al0ckK7ytwWGxzQDok1k9p4tiiYhGfj3BxQPqr0uPnPTo+TqLZ8IQtvB/Ji1Q
qMAQw5TtB/ypeQ9XNMzREJ3BSrSbBpbJHd2nwighAOAvzTquIS6KHpjXlPBX13fUIgPeHWDspp8o
/Q2s5bhkvkQCU476+j+9Gqr28OVSkBuf/zwtLmA+y6lb4occ30DlMUEUd0ZC4XxdsQgni3V9lHb6
YVtObAwVZ52gdfqm929biIgmWtadbWqOH6JA81h0PTIBQPkO5Q9NMl+ejdBwz1aylSeUlL9M1C7p
OL6MwhdQrhcQZBsnyZHm3Cor8WfIJ4E3JFtgPzSNwAaVUG7ZtD2u4wI5L3+mFGx6nibmCjsc/FZ4
QdnedkfiknXsTEQ72nCxKk3Nm1AsbA09WS09rv/T4ORV+ZLvfvY4mNTdAwOqffPMOwwkSjRAzQoO
roMvvfjpttVIhB9hL7kwDCvUX+rrej6S3Svi49n5papnvbCB0Vv6QPOwGFK2oboKZUNajX/NxnTg
fK9nBedzHPzDEa3CyZic4+/YVp8TTX/UVhcRYAR/d5+RaJSGDAI12EAyxSd7tztNPrGiaaX1+Iho
BaJq9GsCnVu/BityIEvZ5xEOGKuxcXGjCWcLPZuCfe+CY5gtHjXLIg62SXc2qlKlPE7pYA9e/OUC
ogSXgW3aFAlmA8cxq441hcimD0xo5gqR/S336PFcvzlef/oCTham7M3P+d/sAcodCBXZOsSMEfvM
gXEmFcv/l3MOU8s/m66RfDCjTFWcyibNztgjtKUugO1c0yAvFDuzO8bNuoSL7jBbm7qZ5qebrbTG
ybntIeIs5QZoERQ/gyKM9W2bvkuvu6cUGnlnsoh7RIb0Ces1mSVbmx3pRF5h6YoyyHtG/TD+hciU
yNsZIbPEbU7EBeu/JgDfiTp2+huZCv8/5kiOf2QapnNREYjg8SwW/J981UR9HEMaSMg0So24xsiV
vANA7QIT8FwvIJD0P7Ds/Rs1qvyvWrbH0k02Cl6DRd2TqVN95GEAhp70F1+ioLWTtY4tnlmDz8oM
Xobl4nyeYol2ziRGFxxRgI57j4kshR7QdG7xREk8rfcQmLd39VJGRUbT9p8yYNKluqJIkgFKF5LV
9kvBXkr3udVaOEWJx5ze/r/bo5tSnr64PiMF4Oyr1ETBXZAofxAT1OLESrNjJRKe/ZAIL23JYQcr
z2XKB0610d+ISn6ryffd9Q00HXrF+QzxQw5tDALbhfS0G9ccEQJyQ6k7y0xgP0MQsS+EWOruHm45
hqZZHq4fXVRI0BjUKfgHYEXzD/3TJrklvfRjn59TEordpjdkMKA6MhBcR3X4o0zwVL20HA3SnIIi
SlTNMzawr3+7WuD6Alno95uWeZoQqBeT3DmccUtmi89PnTs2e9uaUAIVtVVv0YZgsqwrxBNcSUGo
cumHVHwspWnI+WMK39s1j50K07AaZUuPDiC4fEk2NwSO/wx/0ATaTMTR8GnzN8yvSIz4SoRkwOEh
awVCvpsC8Uxdou9HR64nOn5QXkFsJr6Okge89f+rPiRSxpdr1MpizfQE8kvPewh7aooFyrrECUaE
JOBg2p9oVZStRGV9nhrhE+NpR1mAaoFgQWgtpOmyAnTi4efCmiHD1T/1SMT2K36Cq4YUEakkaTue
dA8azHDgMQGQd1LstUBK52crbxH5lRxNd9CbgTikGfKhKjCaflwZIdN6uqz/ytC9kAjsE5/mozVI
l2kh/Zr+14aHFA+QEW+ndwnFO0ZjoSV2ObNguydmIGHkIk+Hd0dBqs9KenseRWzov/myQHM/7YLI
+KAHDSfaWGuliE9EvmTWV/ZEfUVjoaog1wDlbl1GEpLuKUf+Tuzbo4SksZ5UG2zDQJR8iQcvs+sc
yNlMI0iLuzjnQUfKSqEtsOPFQa3ijlMovFacoSRLDPI3brpljRQrKXcR+uLagxZaeiJ373DqISKX
7JkLi+jZax7JKkolAlAaPn8sDZ6/kRaWWqTLuSNDk7xCLYAfCJgWG4SYV9NtesJtZ8rGcodjnwLp
Oms4wPokPjtEmSmBX3/HMI2iJMTtE362T4pH/FTN2Kh+3Thn1BSrBH+O/aGyHAN8pZTWHOwHdBjF
ySMTMhwWq2FzToTjooAbsU0CtJszOMvWPxEp3cc4rYOCwaa6S+JMffcMhNSFNF3Ej5AnQZPsuhFo
gdej4lQYnojNF3MiYHkbu+vRjcrsKvjwdJx9T2iBpdd0iyXq4Yguz9wSyY9x3sdlcQOce6M48cCP
Q935w3MXU8euQTj21SRiEOvIA88wf3KJKmZxzaG/WR48afW94Y7vjEkOmcNdxLwMeO0hQjtiVhRi
DqdgQmCJa40AgMx18TWDlsKsLFyQAURgY4nGHR5wmtw9+AmskmG0NXr1FoixBG4E7f7BDi0eSAQ/
zVfaTzzVz6YcRSZuZzZpByvVYcCyAUf9+jlGQUfjv1F9gXPGWhVRpP6GmUN/YQf5IAGbXPt2BXDo
dIAarf/NyT9X3N60irrn4AyVX4oPovMkQKSiMI2pVYtTa3f9VRLXvxgoBpnhdZzTrspgBhEJLriC
JFlG0mOWB67Y7ZZ09udMd4kt4s/xh92cJH/sUQ+9PX44qfX1d73IZvYggQB9KXpTHdN6TYlPUg3Y
WRSxwp7oUTHYYdH608fXnlSJZ+I6aFPR6fPSBxqE+pQrvqUdcnpuQBRtYng76tf+mJVYaw0FiLXW
Hgrou6wjUlupwqc4Z7eT5AMo9R6v8dF4IxBrZ+X44p0fS+aB6MXM5wKG4QhFCNxSHu51dTmtKQrM
HTOXF89i+clFhBno8duHmeSvzvfnjVHFWSfmrYSgRfDf3uWQkQSq04qF0YzSyMJ0HpeUm7o03I9E
rSFgjn61vPmIfcaZNmY3lsJYkZ2KivhNoy80IvdKgf6paP0PEfFV1i/hJ6IBx6N7LNlmYiPOWQk+
uZdKSDlRn0Pg3mgyZEYky46k9BVdBg6DeVRpksRN83p+AahpO3a+DS6MSObH0Fk2edZnMrqMdAmF
BGORokylHR9U1YkRme/v7uUaM6KdX/MedxkcjOI2n5jYb3FpqW0B2Zyx0e/sYxvnB4jI3ZzDWpGW
Z7x6TWA9SW0Cel9xLMgzjpBwrGtcD+SxXRzIOEOvGHGCt5Ez/QP0a82D5oxeCMOGgQ25YR2cDjEX
/6tL/G1X1wT2yVQu4yRTUKKB1WEfJhApbejugDerIwqGQZPQznwk+vj2D9hqMIyQf99HneO4yxwR
SSaHXx8wEPGAK4k6LVbraVJcDQWwU9ntKpNC5ulKULBJ3Ly1IJUy01lByStJ3mQPgajpgdq0Ssat
WB8J2yO01kaSu/ItOCWeOvRLComkYpFBIf7QW6NWGyE3XG0yrTrCaXQ+ACoZGeaJpkxYoFZrKA2K
jC3wDSceFgAu7Z/IktWFoSXoX6WfADgQsVVQp9y2VqxAdWB1gxC0GEvLZmm4cfYQLoGX3iKHzPnK
oSeGj7mUbTyO7e1wBfq7pmfs+38LjRdtqfQBoSI5Sr+pwYhPKJguSM78pmAQr4NUJ4vjG7Q2WN3K
/iAAUpnCvpjmYqw73HmUGCnNiv7mXqJKaUFvx9WExwO0uA4iGWSnAwR1TUXVKN7658alQLkNWR0/
zHQHkRjhv+j0tUYjeZRrxek9whz5VUCSb4KhfMJHy7ViY9Q/vM6PX2oLqkhCSjGK8APFqtbrVNrl
6xHoA9XMSlxJnZKP8pJ9/PUxkpjfhbavbnI3aOqdntB10g2jbbKnO1LVLq+AX7dI4loCmXLBdV3r
Hd7Brp5qy5jxYFxwxPDVfZ2i3CMGO22C5669mQ66QupdAlTFChRCjbfWI1rFnZ+XHtZLPaveASNl
w+KvXYnhZUNhG/etIh2BkDr9lx1MkGgdRkuC8UPin5qjTv7W5vdjaBXV4g5T62tuepEUtChN8+yb
Mc7/nKSLyf1MTZ8RgyxJWXFpNDFNJrmHopwRKkdkVi1bWv+VdEhlAm63ShEqaDMeEYEfSU9vPGG8
cp0lmB8soP0WRdjQXVgccBMhuN5/oFybZk+umUvD9vpXRgw7tETKeYvf69yxoUOW79XElQrLYT3n
5eEC4whboeQa1I5u3a9VCSVc9dPwBzWlyHtqN0/eMJ31a3NplRJ8+TdeJkhvY979nIs/afDu2gkL
zuHwD1nBuA08O9JdUXe9xOId6zgnuQYRa7vR5k3NGRb62ycr79vQwh+BPdw+S37506IELJX2tVV/
ve9DJ1JjZu5jDk7WAMLRKSxGNjLQVs9+lG61BI3qjWIe6gDPPB7eybZKa4eNbFymp/MvFiVIFI7/
ibrkJwKLTDinCLhULIe3NXgo/FDjnAQI9qTuWT9TKHthQhnjQ+nybADAy06x8G5JgRNBDtRm2PAf
GKPk8MtbVj4wpO0Vy9X2Ojh/6J0zKQzK+NElMQ3phEQA+J9v0g34SD0sdrZnPHpATBiUc8TLTY0u
uos5u8/tOzAs4PumVW8y+6MPFw0oEqsSRPcmMpj/QeXhUj+hyxRD3WKr/WVktjev0ZahFzcVba9W
+q3RCALw2x7enVTBQJ4/pmc9K5Bwm/oYNEIY8LWZ+sXFDzwkaKugjJKwwW4bEiTNqAbx8fpH/2rs
3v3A3B3ERAruVOJxM3D02ciVuv4nQJ/HYwHtCN6H/R5hdTSPWz9mqqjSmJS2TT1kMBywzXQ63OQ4
b7dWHmsafFmDBLU3Ft468mly8TYA3gkN5Md0sbwIo14MUvPcK0HHU1DRw4wWkIhIBtn2macs9+lK
h6jkeThE8GbAeeocVh2IDRISOOw3COprmtFQkUcHf2IqcaetR3MCx13pjeibHwFoQlKFUs8f0JRW
WVHt3wa34jnkwYFHOEUiHhfgflnkYrdEYdVOfpz/iA1SJBzI5eOiGxt1K652YazxL6lC4H9y7yGQ
bFsRKAhCgpsFVPyVVeWqKRowEhnyrarLk+6uZRbpZpSiQ/vAJlU9VfTX96MmMH3UfIdAIP/Lkvd/
DHwH+h5GQc1flCz0OSjj0REVbgEFbmmskDwPBdoqwIj4HB38v7KTDz9X+2cxLdV9Spp/Wihw11hr
HIll10YV9MBhXeAazPLz8XQvM7uyZXdoKBgIxJH5ge1oXmzeoAoClWSNEYEY71Uqfk5eu3J0Inf3
7Lvz5nj6dzgM+dpqumwD0Zs4jkVMGUXXy1xXbm0qj5hKSIlSTdJJ5ksgUIA8AS3bMRpBqCh4N3PU
cZduIz+bAwT1MMfw6Sle9C+gzkesav06hpQ8R3aeg+ZCwCj60CpGkd/mqCA+1qU46h5p18pPQW1p
tXdOYYbAVSfKMBZc5Amk0LjmZQ+aXXTI63fTsun8OmuVZtAYYnxtafUqakQgVwqFAOyO/MQ0HsJV
1qg6K3fPKKEU9s0RPXeIGCBZ65tGf2LdMKs8RV2fKsMb4ItfzQxDExQ4KYy6gbKc+sBoxkdE2aiM
jKHEPgxBaLUrvB9fOCOxhRJRnieptH0XPqDebc8ADIDlLnAshkvooSRwmWjKdSf5Yw+ZK2Y+5jNy
WV9XXVY3+PGpDsxwbK7uHowhny7ZwCiML1vsJizZmgPKvGlulu8SrgyOPZau1Rv7LHoTdZkfoNo6
rsJpBcCHJqZ9G5NvkpuO3sgkH3zjz/CJweGhNFeujn3FG845Q1vTaK8gOFmF5I7pdP4n4keqHO2A
SBqaitUTQw/BZTYSmZdvoTG/WeqxYK5Bo9m+iM66yFL1LPZ4Ul24TNRiOd29t1XY5zJlyuIaBrST
629OE0CAhxPXjh5lA7bLS8qxSHC9HQ/+4XZ8KAIRD8sFSM0n8Va4CLRAmaQn4h6fC+dm1AbnCUG6
9ihMFAniSfxaWyfA9eABibQit2v8RSuuKy1GGfEqHAJPPw5beax59QszLhAMPMUQ3kNwET6+UYSu
rM3OJsnGYuQbf8uO1I7O2RAP00xsJpkbS9Hw3d+f3NHdY5X5j5ADE5FhM8bOUFTvlsO88GnbmCx9
v3NhHDf+rLuKZxKthtpv1elMPxjmik3XiWWYNmhCQeDf05NRGbUCeK2Gzo2kAuKMiyMn47hRr1XR
kamy79fxeeUBZFK+kSEjquvtq5JBm2/cBdaOCghTS4Euzrk4F8b2tYvYysvAf8smctB52juptHs4
Dx6ygC5RycjO2ugleZfUN4dgHfRcFXFUCCNSjD0I5mDFDwkl1wsBHPW/S9M4lxSh0k433HMNwZWL
lp70fmifTlUmcW6oVbFlaa8Mnxx07Ee9nKQWALVXV/dt5hQ+bCuksnJgfFmKkS3hcRD0/RiiS60k
235tOChM6/ly6yPfBG2WqCFRFiddlnrzizo2hNnJZHsZSrG3UWX9gV+iSIMyVuirfoDWYkrh0nqC
1YwCpPyu5ookWuXC6goghYVajZJIPF5p/eEiHFW4Eg1ZFofvQPYU2kNh62nmhBh7WGQ1r0Wyk0I6
oDk5kvrOZKddt8UNjV97VV1Lcsmw6dBe0hNVr9ULOJbqHGUfCYLZotxD38GfsRDFfA2OPtP9Tol/
k1i2/YDA4dCIQK+7sVda6619U/nNi1ukSBI5XZ6BxYOOfSaRbbAaUs2Su1PolvjTPs8uY7mw2fZH
trnBKNzMHr4VERKAOSLXGm2T+qguA1b069Po0Op5BeUgGgS2c8GsAy3VhS95h3tM6J2u5S/vNiA2
5P89//qRKvFs7dKAJBwGMfIOuPfFjz3evKdojUvBPL/kannCRYffBd+rIKgbCPoZw1wAP6kpUf5t
sobRgf3rL8GyTPnNgVMgHkgGhdxGPl1N77Jm5SPsynHZFYCRjpOxXaPv0fGFZbTYRpnpZISIwJFF
ctGAC97aSUl3BR4yWEj02Kus0eSE9DkgHWW+v6cTIQsS8jskU29y70pHHTSeu0P+hsUM235cv/i/
KLBldJl3ZE2zgXpJHQn+/jecMacNAWP+LQ6j/MdzIex8nYu9VUejoOqTCoLr1F/ZIJB+fPXUUU7Q
LDjXhTnKznet7FO6B+XsgF3hdPOOh6UxJBpPz29bbjNBhTJE8pmrOzvsOl5a+KAKAzPeEXo7x0De
CxS3D3Y7DjkFFsBItrHLUgsQkdbbyxITaTiY/48eGsItSgSFrbhIVAD/oyQPRJ5nqS0ykmBIGx/k
R5owZqcqQfA3tTkezkcOpM6Nllq38vutXUiVkcm592kpo5VF7Xcv4WOehgLLi8RNXjjGqUTpy40g
QsyWkqD2kT8DGDXlr/hCIazLWxipvVBThd2KiJAMmk8YNzqx451SoZONUiswFzF1edeUMW37+NTz
ntN65P1Ev8ny3jzvF7DZ4/Sko9G3DLc7ATu8yLwSGx1+AHyXGUIle7jrD37t6HHRAbP+fwF46GA8
SB7JEbD0OSyTsIhv/9PtJN9PJcYsXXPzKQyJhKTo7QkQ0sbXA2DuySLzknYQvBmfRFlDEyGYetw1
reM9ADwgurKo9qnwOsvYS/NGVIBVbTFAEvz6YdKc+r/PBOW6rEzPCONjyqvrjjw7/J8ukd7C26jy
4zjmb7TSU5Re2mec2gqZL+qdKc4b2HKaKHdJyhG7QDeSiqWf63C4X7HzE4Hrw/P167qORYrfBda6
PaF8mhRJpHdILsFQMhugfQCm3D0vvlgl8kunxmfzZEJIU8njsDXdXCqZKJ1O5wQyXzxMPSIWfcYB
LF8RbdkWP0te57GQ2LLcI8HRvOShqbg9vQD4eqyWWx+17XdMsHg06nzKa2pcurHM2zYJcGCi7EHM
Q9UW7YsUALfgMnIm2IzPQsDXZdy/BXTcMBh0xpy4GBiUIvC1TdUTZ7RmrXL5NCNCRxkoe6TOnMGQ
esEgpA6CseET792oujMnH1mFFra75UhZa0xlwmCDECRBZE7bF1fn/M3Bla8N5NAIppvXzmamZEmX
Wx2sUD1QRMJFyZ6DgXZzcvlg0qZXyfboSXBa72qy9OHpfbsGfIXpZuJRtuALztm70opfB9rmv8QJ
FzXCZQp2SkGaL0Zs0RayTGgDP2SVZV7nZdXPckC0o7WfeLgeK11VDD0tGCwmVmO6cvddA9sFypf8
7GtZL+++G/4fYLMH//YPURu9aT37xgSF6pHV6cS7LGFdpLSC0eV+lHm+kZqlG8XM3VpWyehxl7Nu
+iO968j9TEyOId3OpxxDo21oYA5hr+VjJqMpAJKp+iADJ/WVHsYdoLGVU5eMrNsyEjEtHAy10QJJ
uLyZdQ2DIhYl6YgT3woQQO1OU/aMbDFiYCUgCIrrDDTSU8VNMTVxOnsZTxaAHfrbs1ULJFJ91yFN
UsjZLuFO48RhGX2QehOZV9hN+YPtm0j2JhlnooC/YDTIOUq0q5x+08ouRg26Tm+M3N4QyoNGYomU
+ZD8f7q7uRnXlwzf4A4WSMEMaLSaYDeF5p/NsrKjf9PrVR0TsUZhAdid/m6XlgjH9Pzs2bsE/1AT
jP0KwD8VPnvZ0fC8r4+5JGPCPdKF21OVrNBY3Talw2sxcSYeU/Fd7FtywM+l+N91Zd42O+qpG6JZ
n/gJj5uQbhdxCnuysdWidtoH5xFpsh9w+7MPGscQNhiOrX7oiZKALsBC6APppa5xFf3SD+ThpBM3
4FtjTuVHJ0yYxeUyfbQpSfw5IDjYPli0ULPSncEw9cBRGSdZN3AUQZDZBD5CDDAKfVyxba4Q+YS5
TC7UfbKbzj8psI+/U8zlnA7u4pn6sv88Y0jEVBnLtvXIb7algAGGRZP5VudHxWDT0KcYfsUPxR+W
nebFGzufkhlS3WiQJ4GYg3UBKVdMn0FJXreLK3O5nj9NqTXyIx9J2PG4vHjSxiOCFmHCIFy5H7Dh
AbE0gBUqmJ1V3V60bGLm985rHSxgdtnMVkxULiALqUIGlONsdWo/lwWAGwyBtn1M1nQqGmNKh6vT
dPXx3g0lv3hybOdqkUz14F08GzWRb/FSa30oclq0orPJwLecVevffqNzeIWQV9zRf6hbbfvf/E/y
2ZsXnWw6dc1ssrzYzg873d8OK6A2/k4MOphB3+dV1TAMnNCRhRflrePFDMsfYKV35P9FM3V3VYNm
jVc0Kf4y2414D2o3Rbc4IXiA9ChmuaW3MeXoyj3R/bqJkBjBzS/HItjpcycKBs/fxZ4DjAJY3Q4W
EKxB0AvJNvG+8JkZzR/j56HTfTXxIcUliEShb1YgumyPfIahy05z9mQcpK7BvCgBFuI1v/ZoOjXQ
B1VPUbGXIKDD2QpNwnCLAoyKhEl01JLsfPlLgW2dAM+l+cw89gQq6uSr2oSUWiSToVTvCPUe67W4
uS6VmqEJGmb+pyoyIFrIVvjfx7EELQgpRR9X+0zKMuTdKbAEauI7y8pJYn4UfoHR/z/kA046WQL/
0GeXC30eu8Y9xtFFrv7IwC5RthwRHiKKh0G/sV2P3150bIkMKXV5n1CvPYcQa4G6Wq2ZX6bXORT9
JwPrvN8JbQpdkHs+JWprJ78g86IBoPfcY+Y0TFOlAZnKZIBheiQImD9rHazrjYY9gUYjrMzlMKWP
Qgp5+e/31HoIjcEJcfL+OgULzEmYCsumr25EcKcMFMY41a9+nuONZp6kTjL6ftWoiZYONXPvguoc
sheLKGT6u42CXjVnKq1H1H5evXPYKgtGZxP3/zl4na4enRGL/ET5a7MxGILsZziLK0SzztVA83b6
gLSGl3XF3YsdZasbvBzni8hoW6bEs78ggwkxalQsDAkVEaEQMir9HrHSRN+d9VXi7v0HhpWsTXad
nDfncmbd/n/WuL/0X2ZBMNEcj/50OCR6VXWe9ZB0mgExK1yDB7r/zhRQ6xJDWLbLq06C6PCed5Iw
QzBaTY3r6X/K1Lws8E4jTclUPAwMep9KTonqrIh9mhUqiomrAqAJQtT5pnqBe9MtUSSngtOnbdeO
e+dg1p+z7rIVsPK7LSTHbMMl+b6FQVJSOa8Ncur0I5VrE8Enh4H4tizdS1vkK4vpGUNXDyQ6DmxO
xIL5gcHETjy6SAc+BeFGIK8D8BIpPIosUgpuuyM3ibH8O4LDbAfluPBF2sotIk5AAY0MuH2Te17Y
ZFGQNzSuTGH/pZ6uSzZOu8zvWRENhq6MWirIf/duItIXj7Kls/mHo0zjkRbV6lwzf59FGnY8WWW5
JxQWiR3sZl3jLL+WySGBXzR7MSK6lBWTsXpk8RIjm1/5tAqlt1ueqWkzQArH9RXbIkF711U/SIHP
4SKrgpJ2VGf11wFsGpa0sOTrtoB3kJbLhmr7X6qubSpyhMBPU8WY0wviFHLBwi6obJD7FKqwAxlP
WhllbPzHHqYG5Jau1+Kvhat9LD7FO686DAefnLB+aXz2zoRm+vY8BuTccAXpVd2wfMmqb5orS8TT
CcFtj925m6j9TaZ+SFBN2OKFConb0VVMm/jn2ydYz1lzHQP15O23z9vCGqdnSeIXA23gCyCdraf1
MRrKN4ZtTfrONPehFRzAn/BZ3vx07ZxEIa7RUsrUfAfyg75rGAbX+U1EAC8/AmRr+fXkdHnwzdc7
dXf8cqWFxxWXok042xwWsI0AIBtkEAN4GvIohthHZBdxXM86/SlhoFtUtb6COjxvGoAfu14wlbQ7
U8Kl8M3rXESFn0BN3ouNbewVmZo3ybjRlz0+iunwxAbkfK4r9KujYW31ZCPDoybjaK3HDX7wCOCZ
twf3QgY/Er2yzVuQ2yDBaF7ICIOk1Z1IZs6xz6Idj+GbBY6EyOIjP5iQyj7UqvHKixtyo1d3YJO5
VI3vaAlCjgM/gUSHy3MSiR9RoHVfx4jLTQuGySLka+0VVQDqyQqf59900iwoNDMwK0xY+BRsIAjB
PIEdZvGSlDhD6p4OYdyyko977euIh/eYgKq1ogmHmRMesUlr4LpohfyX82LOZ7w3uv2Idar4eK2H
aO1fl+2FFVPw7I2e+682yx4pJpGenY3Rfo9jEFO9hSEtTDzZMxgvoRs1GbdyKm8SokAG4oMA/ZKg
6bsvVlQghVZWxOtPK3uIdOgmiR1xXliJ2ZjZ1e3wtoPmMdlhA6c6YKhgocKaHVoiG/6KRrgDRVTj
81t43TkAnV2YgFlsCVOH4DnxjrqyDOcDrMUzSLbL6/MVDasN340Zc6wkW3s0a4tMYVD6BMFunTTC
vvb8OXexv6PZ6W9M6Ykk471ThAJd8bA0jaMgm0qCn4KQgd2EjVYFhxs3Z8/TLsAYndqxJckVD41G
4E8meY5XbWhETI+iG3GwGaMTrP655JeadHwYHdA9bLFlAuFfLW8s3MJC8Iftz9mz5Yr7Du8m+PAH
51Nc5ow+tPT9gLd4b2qL6DUZvOJbU530eeunvnttZHi//vqCM9KTyAQIbSccbcwHqyN30o3z/18G
z1fJiofleWCPECdSUplxMOrtwzaKYxqQ0lL7SwLG7s3jc1OK80xZZetCFXXGpN8lEpvjXKELRbhh
ngHXVIR06fXxErcPRfj//JzJuesaR1sN5Ky4x5C+2wYIl+AU1a3ALrOcMeqWxG9vugeTwS9g5fWv
j8w+JZJpupOzrzg4cfd6i7x/zwL2JrmRD5lsqg0zasNHNB99bcHmBMsvPvhBvrJVaZ1PTxTvGzUc
S3rgYEESmRbyuw5Vu/zHsR5j/aT6ir4NY1BIBPk/5ymCXQyJZqgCbWz1QVFRsuVvHz2ECFHghHEC
6Dpc/QFSLHQL8F+5Roo9k84YxihCik87ky2zr7aa8SdEJQKATnQ8HNVQhKZ0IZKuCJHmrno7rl09
dj8TVzwXP0E5quP7QX5RrhAxILOCrNBpUDBkQMS3icda8e1lNOQF7tTbGkQoeXcc50QW1ObLYMHq
EphNRDqb5iEepuCbeqgLWrTo6JtwUiJbyHBEnRSizixC2mYZu1Be4In3dR+N0S1/VH7AepOp4BbC
uxX7S2p3ucO2AQxqbv62jWtpkvgEnOGFQX64OiGXVgTPI+PQAxja3ipbE23jiMPWLA9IFqmaubeS
TxRAcVDg7/qKm3rByCzbrbowjGu2TWYYWvjqzU7JfZfxK0nT52ycZ7CURBnVwwrQ+cVbo192EHBe
ljjC73hF3bpMHXWRVl93iBVd4JsKlNZUo4QfHDnNkGDp1iv0SRa8EIzkChQ64iSq/GC6fjXiyLBS
lg9LzY5RoCXCWN7/B220jhwAv+MDbIDMBq2hBL8lQY1jD5aOKKxXzKCwhjNr7A3PAodecDMS4Wdq
bMRgwpgx9vQXuny96SvsZnHzAsl3b+E2bhtJqtkMdJeY8EoNQW5G4iV1KrOm6XSft/+2URRijbe1
RyasvLseGr/5nzqbx+ZhJBPz6vYAxw5HyJWKYJKJvTndqxVKv+xx719yd/Q04c/61j3+uh3qL3c5
oZeVwqwYmqk4pWWHCobMwuntsLMlYikYnFssU4OGeFQieY91x80sIU1X9g6VJ+fr/UNi/EqwzJ2E
ATEehIsvZVdpMAdi6CAABjXORdu7SN2pZ0by5BgH5VfxQJVqtC/UiuI+kCi+7NnDnEhp9c7NsUR8
ODa7lgBPzJpcetoTkPIwjeXICOgpSkAOw/Hik+Mg93dZHjD3a3Z3T7UVwEleLYV+G5QYjm+KVL5G
veyezjMyGGzeN/DNPBLD9J2NmK/J8O/5w+0I3Y1A10yzFq+aYOiVvyeu35002pTruD5JS6Sr+yFB
mAMfgBsTyb6Do40PKlVv+zKjJng7nvCWSxJSHyNgroFq9w5avzE0bTYndg8GGCznalKioJqzGIfS
SYiylQeeP15qIEhfzFhyBI4jVdWjcBpUJcTz8t+8qUPkqyoGqxOw/OJK00oxK9Tsk+XrPkcNmiQS
7THgDAHYPcOEnLjXA4th4J7+1bjKc/idj4dTViKmzjj35SCUMHJ983o+llTcnafW4GG/xqtabWch
cLYA+rAkjZJ8kgPw5mGoKuGU6AzEhE+OAaFpKf+sZu2jfRPoTbj1BJxG1cJZRLNHtEzvVBNp5zue
dNkOYjuVAhv627PrF8Ws207TlkTLg5hB1QcYPR+hSR0AT23doZnOCDG5DgPI6kxm3FXhiQD3eQif
mhj3lEpPkEFGzL5QYIU9/9+jP0DK5x/5e4UdxXHZ4OZMOPt0HeDVo+938CEb4LiwQZoC06lk6LuQ
kymTpFb5h48ZAMeqmDZTTdPolsc0SKTlzIpQvPJdqZqjzfj3KgEti5AOvYvHL1jWWy+0vfpxc2la
tX9lgIkIoG1iu0gEaMyTk/Yfhgq0IoTwLUVJiVgrQ01uLdv2Wm1twYeSF1WeVzJtelamfdx2jv1o
wepGjXHpyXIUD+FRlGamP+6W7TZ1VopdI4UzjuUvMPnSF+c1nTHDzDz0dmGebO6E8aC4WLpDqrf5
XYcXe9NK7saIl6JjXUW0RNScQnqFgBpxY2sa2gn4SyzuYvHB/VmJqrVW7HEd2XAzRYytLjz+AToy
+v2FoDE3oSm5IxXdXgzizc0RvezfeyPhAMr5xN4zvASMx8hVFmfJBepj+2gR0z8zCx72+gn2EnLs
SDVZ3QmvbvjsndD+HtT4BhoBkamx9RISXAQA9syiyKfVOlesEZoNhEtDaLl4LhANQu0KA+nSX/rq
fW1/2hSTv4nQ+Vs0ClwrssdBfoE6zHZQ6s6D5/rKWx30SZK2yXlhZUVujFBtuavWlabgznY6tMgG
SRGQlU6+dbJJwO8ttThuiTCUjr5MscnYoqXWJsejQvPduwH5js4AXD3xLWGIUS/cW1b730KBmOHj
HaMuMpzg2Q1CrnzceMNMhQZmDPudI0w8oYN5bEfyTtwuOjP7YCpcc08sPZqD87DA+Qhr6//xnUp/
uq/yi8HXE4ylJXM53gLxF23Zb8/ph0oR5etyspnryYqIITFlJ32pscLFu93AV1cIAobUoko3Tj9d
3bYswJfQPSZE4UbrDz5FPVGSql0uT92i2IDrp9j8oK8ELAuTEGAHg1kwZ5+y7c4iBbwAX/JKaYVL
UqnVO9zMhKZcPBBAQZwYkUCCnkwgfdTtof7Yr66altIUOTRUZcOJ2HdKxr5SAgWIsmHygQvojDW1
zazRZisbh7P6fVHbRulw7uiZW+h8qRbqAm/8lqNacs1exrMDStxXg6sI4oq1k2j44A5VjFUluBk5
BKeDTg+ua56Q5HlwSEHpDao/Bi8JJODWVMiPqpnoZrag4fzwaJmLT+n+Ua64TUpsTSICeIlJeYyD
kpW63s1Wu1fe7/SiauyILNAWF9rcrRydnlLLfD4myTmWs0Gt9SDS1rByWEh7t7q3hCZ4mv7JtrwT
VIoiGHFfMWt5J5JT6luMdMEI6IGGR6OdTpk3JdaTKP0ZN3mM4eu8dwG5Lzpd7oFGX5sFbKb5AzO8
Df0fJ1iejb3VPWxOUBhvjXbmsxzeekbzRol8cJPGPX7RJJu8ADvnE+U0Oepfl265IHzRvPoeRHoJ
TR5Upo27HpOy9YL2Kxe3U84mFX5ixMrfyrB8cLIbLYlfeVj7aWzWc2cdnR4oYkKPgSwAEmpjK2NS
sEbIu6/DXzGO/FCj6qHYfQqiGyVfwH0ipwBV2YeLMt/IBjReqSO6oPx+/dvNpAu9ENUIVqMtcwGY
Ejk8NymYoK9sHQJzNh2de8kSPUgD+V3iGRY5W4vbfIAEClg87LqoTffqWD4diQHLEo2jW1PEo8yc
QnAaXUwWiEKDf1YnHmNaHKIiUzqtX8Giv+Q/UEHmCuEfkmI8PbHWrLRVmYQusEZPGglc67vgaq8Y
aeZmlcnbrITF90/89wPHvl6LOJWzmFNF0MiDnoy/V7IY5ORZfiKyc3fCMFFy6jDC+rJqMJ/TeUeO
nKZroY3tKpfhUTzOUtgJVvZTgQW7J0aUlL0pJQtGZr9sQRjgo2eDbS3d3Otz2OxJ/lalq5B7mEOY
+4/wyRypfEgzpOQ1xC2OmJgcR/f3acDAOBUvnJg7b3V4yx5NwSwF+X+iCTq1pXnuSd7c9gigWZpc
rbhw3zoL0jU/Td58TeFNGNn2f3QDNIAP+jd+pEjT7bwVxhohTwKeiAiX5XpZJM9cRrFCk1JExOhz
RGB/pBqZiF1G/BSPCJYP7dbSSoQBOgxMkwBLkvgVliBwV0Ht8QOWlJHhdPCDtOphUaBhokWcrkpz
aGgBkTMsZRuuHyn74Wkxn9+oEzcmp6In800c+7v78rIQM3s9LtLfxFOtBGCqXK66fSfpmHkO4PcV
IGtYJxg6aL1vMa7Iegkb45bdoMB86X4B5V11jpqKlJ8+6jrncG5dGWdtUiKxN7RTn4HPiLgccv82
ZUzrt6VbGulW90xUK5DFEwqoKycmh6a6wmTh0SxEKaeuymuaNxQOAO8l1t4LZ9kMbZ343cOhR05C
VV+gsu67vksK0kuw2q3+jNsQUjF1Iv2Y3MD4VhXqea5DNSgv6sDgZhAlx1Pq7CYQAylupx6mQqMp
OjM17PfKxe2nkt59kqWYA7CeYo9s2z02YlCyF1+unM6kb3HOxswH5/DSJOtV89HB6qM+sdcKAQJT
XgrrpJLp2X/PLZw76wskFqrV4CYSbRhnClHsj8wxfYI0BATkJN4/I5KvbB6JnKOZ2XJapPmQmo17
jo6yneaP6e44TC13QIoGv12S68aDRnbXqXb53eFxBhmSbMkHv6gVS5GhEy6YEuOdbb0biz4eF0sX
9yil1n2KJWQIiOXpymQh4O1WVg867RTv+InMLKkExxn4cpxhmxEFJjmzhtEs7xTddBUwQmBSFBxG
3oRdhCPOhKshzRXBtl/QNoAq7fIK1pAWaP+NFlarUVmJEPfiwmU2MUcvqgL83h2uOwNabntLMvZi
nTyosOvHviWAeHXv8JY995OS5qD6KE6hEZ3gelgOGWT7XmjaKTGCHSVaNY7D1TILAGChuU2oJJc+
JxpR5QkOj4M9RBIUJoctMJ5sg4YGLpXybX0pxqhdq0czSyIvYVJQ7PqFriFswuBYDqb7OV+CFfpi
HKQwYm27M6sicOkILWxGpYXaBEvbVCZ0/XV9Nyq1rJSLj9vQEqdOs5FwAsNR/Y1O7BeQPXGqXoie
T31/FwOaOsJYaEKfXeJbYX3r2O9IL83C8kgtHnkd85ugg9Wr5bDCDkEj4N/ul7iuSbCIyd6sO1ka
SG4sXdqIobfCVk1MxA+xRne4hTBdtGEmKdy1dRVp+Bs+CnhgmVUOGVFaE3GnuJKEoLZILRizFpQW
oLBdJ/faRRs/YmyLu2a3fCKjgE4YCGbep38DNQKrPU/1H/jeTrOWm9BAYai3J6Pe4nHV+Z3HHwL4
GuHhAibPCMqZRYDX9Rm75/uDVQIdIMm9uCjSu0xOfht3j7ZgXOBTvjbnjsa3rSE1AXtLVmrjBtae
cNOClExHy3dq1PYit35GH/Pjo6Pxqmf3wmEqV6XKr8zh9M02G+6vptRDVCIVVQTbh3P6askqhUtz
E7jz4QYsC9i4UgX0WW4uqTn9UaMvwgdvnuqQj1ePKosUI+fOIhHtjb0ODhZ9GaxQQACLaHnGuSeN
ehbmUrSkZgstrMtoIpgeuZ7MTZNJVkqoNoLs61uATJsmokvDzDzcGG/r0CssU4QF6cqjoWebZng+
3L68T4GuvpMhhhoIEzZOwiQUPjBRNomyCYeUw5k+aaH4PHgEZgdoD0tU8OAInPAJgFLgqRm9szJi
5q7Q5EctO1P5jdcKRQZvYnEn9t4q4T7VglPo1QJMDllinPaOkicdyjgXgW6WBKHqsQkwxxChisfO
NjGrYLfsvTy2rd5IdpIVfewvdxXYnsBveUXQgo3RmArnMk4U/MwxOGk5yNBpj4/9dcRVgSEAnz3x
ff9qXuHaj9HkKVRmNiT7MvsUEZIRI3hcPloB+GeW6CgWRc/y6rgOiHLQuEHmDReuxOMTVW0PD0XP
KWusRI3sJm1lFRr+t6fwgiwKoJOJ1U5Q1EBaWSgfQgD92yN8njOD9zVYHAgQWrb67Jh0hf4rxrx3
ALA5pjGP/JkZ6YnOZndxdEqchTbiR0Z2lhHohJGPeRg0OjswDSXFJHhsIRM+4PTO1PEYt6ZBHfl+
aD7dM51z2R8DqoSmkfpWxYU5oOddVRW2E4QfQwL3uSI9IicnlxTsQgbW693ksVE280Xpno2+wXy/
Zfa+dqYV5y3bRavm/7gBOPfxuF7GEd/hB+1zTJbJtawTdCgFXewCU4I0jsrYOzhc9nJAQ12w4DLd
uovaZBG36CThtzXROZYAm7GiYRvp/9QcRiNVHuHp4C4WAsNIHrSFxONpf9R/UdOtpeMcRV03d8f7
ph3hxB+/FgZwRkxxkUQ9ES5xiLK1Npanr25Zz2dXAKCgqwFgtapB9U+LrjuBNFaNad2xgeVevgLZ
HJ/oaXwjJFdTp6JnJaNxN7n5JefW8mk2l3tXGTaUQPAvzttDpX27wBjx73yTW3G+tYhleStliqA5
PJRQ4MttC1/SBxzv+W4bd9Gyc6HcX40u7CF8xPKxgj+oB32Vqb0B6Pt9TjB15zrb+pGXZRJAbfGM
Jap1VHzUfhnuAKjYG9hXUV8s4UnF3R9CUUEwbMZIFA6mUgHk7gdszAenJCj630RMXmvw6FfCvvFI
fpqylkEc18RwNuBiBXTI+OW3EDKHFHRzyqLAS/W/gY+dFU8b0W4Xyn+TL2iKOByOw4irvlV7Z5rl
mxZA9I+P4AXhr1ywfPvhSODI67v587b5X2hIFOlY4bdbBIEYwGhJzijgaIUJARaAzc7oNC51lhtq
qtgxk8CWK2Fc4VFht2nAMMdrOan2ihUtYepz1ZwNf0aWMXecHjF1RdnLse/Ghzua96v6PBWDXKtV
swjioFXgIcWAOCwToTNow8w6gMU1mklJbHjsCxwsU/2OCMO+e1/53ukFwobpbiSKXbddQfvaKiVs
etRoVT9JsSXpZLthg8Y55G1iAKmf8/NrcOjVqa6KrMKcIEjzE5cCkwrj2dbJJ/z5lAGdvYKlSmtS
CDu0v56Yg759g0H7XcUL3IwFdc/aEVodV19uaPWg+j4PuJB5Ioxu8TjEFrJUg//xOaQLayZlxk5A
7vAuDYBf1gDzKB8e1045fJmPivfkdGfaxfJEnGDMfDRaZ55idTL8liQtb1L2cyUAsSQ/XQ+036uP
OciSyRTruWMMag4jNZgQ5qybHBDt0UQvxTeTatX30Hj2whT3GQ/BT9bg3A0PcoKsO0TChN+iPXbe
AUaMATiLGZJl++yTPwze+Wbv4axdJwO6QmGnBvn/qPB80PECwe51sHg2pdxvChbnxTD3XAQEYlGT
799E9gMx/BF9bXAt+vH79RtJzO+IGegMT3icNzLwT3UHbv9N1tq7na9y9qSQv061Joypqasgb7hk
IxdvTHvkA46U4MYZrzbLwL+KUOCVhPclWfSojhTS372oGA44WITfbfUO66Dy9Xq6wCPHgLu0Q9r6
9QbpKRZQhY+MmHnLlp+LiUNWF+GTuLLTo2GCrkPRhkDXHUCwA7Mm2bhaxYW4WNZy1H04jpzf0sI/
huvrsxyS0OXDGG8DUyyd2T6BDaeB26LZaiSgGInddxQpZ4sKQD6Dd23UZIV9pFWQh0vivqNPw9ag
LQefJGvlYSOvbZr1hTj7Jt92QBUTKUetN5+ij7l123NcKzsbP184jvxpuTmgH9crcG+LUiUMRzex
rX/bS/Gw/lafMo0vg5XDNSFOXI1R4x5cqn+CvzpR3+4ar8rggmy9uW46H7WkncQsH09eR8HjXaZI
Q9UjylcaieNciCG4dDSYgStlZo2tXQaoI6B5mhJ6JouDyusFFPodWXBsXkFoCs3LpXAeBfx0CKEU
Xjl7wTcAlOcUObeD25yqNpwvP/g5OcZ00cDBC/9YtyO9XTyb4ZxXe+QVou8d4NvzFTdcRX1JFSew
6KyVy0MbMX8tEof6CPArZ60KQyfvVV+nFdalEZwqK48G8vi2P8AiYpxSxiV8npbiHIrgGck5QahW
0wunpLVz0NSK/eL6jCUSXEMBOdotnPVs/zOPUMkgnPS+XFGU3A5XbiOZdl0p5CPYEFIB1jtGjiSX
Ju7vmf7urLf5pt4nJ3638G18NQaMd+4KbhimMfsL/Du+AxHbc9cnxCcF1+sNM4iYgA0A9CRyEFJI
CIxF8AjOhGibL7jBx/yJBXIbZINU3KncnIiS2GIfBnxQGe/fWp5ow4owww6k372Tw4yZLQZmr4Ub
HTfUSzvIRl4llsx12nQiSjcww9QjtYVGcdx1vVLsRrgx1Icm6DkJCOUCNzn8pZydJQh84i1yMFyj
zG0qXVlTVpXK51U8eg/5MyZFTj8q2Vuyr2LtvMLJyWWODciC4+2sp4dpikXqoC4KeJ6YxGwBdQm/
vpe5dFpDmV4l8q1lqE6doyDaegk9OAFQlFJ56BiB48up56+ew6DycR59fkGBY5mUUfsti+zcLaFY
EOVNQ61yfzHH5ZVEpSQ4Q4xL2veavJk5jniXNBmYaObMvWdk/QZu58dEjLQlurrZNAsZZbLJLik4
F9posvkACaLtI4rdkUQTBRcL0ImouYp93VSDhdF+t4zlI+v1rzic9EjKcCjnjm39Jbq/+qsbNZCD
8je4kZv/IJJzdMxj1HU+UJvk1MAh1TcHSvH0poK3Fogq4LGbgK+gi07mlhtXuTDf/D897xQeVQG4
A0h0c2TouV5F6RgkKnYdVD6sQ/ua94Ekm121S4BZjpfZ9WBryxRdxVuC+NSDmKgDozkNua1kzgE7
sAKAg5CUZF8GYJazWCVXn8svpvtwf87BJ2wZHMRUZW1DSoFS6QX1/wJMbZfjDXFR0P3M7vN6iEa1
n/4c1Wju5ySE7gW6Caq9lU8c9t9d6U4EEWqTK5xHxiZpttsbhPAeYBfo98bPRPUKVTZaDufXqjcb
ZtmyhWQN6EEehvQ/lUx6531iu0tuOyVQq+oNK0JotoWJ8OuTvxtsdwwd0Z8BQ6EnhWj54vlZRC5Y
4PlrBuFJtUT7Q5oJI27uJEXias/eOIg8Usd1wyX9SmUySv7+XkJ31noLz64KB+6Ln1ZnXmgpuJBe
obO3pjZHJGKqyGd75nAr1Ymkprln0HwulCfpu+kn3v4g5MQ58ETalmai252ai8Oo5yDU+GlBro42
cyWVXfj0RTtaFWmzU0JT6fS6opRd5Y90F9I+ZqLggNuyDrdkLOEZYwB3mjuZmqcHqSPbNn4VUqfq
Zf/t8fxuHNtp2pVjNt25K/MBjh8N/Acz6b+O4Ecb3J3+WgVvQmPsriYVIJV2yEScCzBwGE38Mqh0
V9/AETAIA5CN28ZBYFZQ+y0gfOJcAAQF0opigx6ssqtFdHw+Vvv4n4/hNa6UVBHEQqkbzKPmTpHI
BzwPiq9eNENbELJEZpqb91pQ0uXHnTNoD7M7sEnL8Tc0i5BwUd1iViNGjWJAX7b2xXRtJSROR3F4
vaFKsacx4K9GLMRaDd3dOJTrclnhhcOzjIYGXMuenrBO5BWPLZPjWBFX/AmBmKQjQDWphTpn+Czc
wZSpgcGoCKorQJ03zFMmm6x51LT1GvHUIuQR4NKkafjQ8SGElJbDC6M15N2BwjIvLnY2WquVvDtJ
/d3njlYlqFHFeMzNpiKLcLIw5zJAGwmWzb761DxGZeTYJa3SENmr2hIy54iuWf8gOwcTJa87c/N0
E+FguVSNEsq4v65N2436/EdvL5eXI73ghZfKHq2lgFdPdcKt27N/ubI2/RfrRd8AxshYwr5ptIeA
W0iH1L70ywxlE7vU++6pyF5eDqdVW98s2qxORYUW5fH3v2VGSCCJ3hTxjLU/PogYx2Agl5P+9Yhq
saAoeoqxh/XwCHFbfuh0Xpb5WB/qKSTuOb1fRk3v8mffpU45jRoO58m0fiLsX3TOSGIGVjD3/znx
ISmQMHKsvgVgQorcExB80e3151jKxYquHmbdamFxePVGPekX0XPPMAFyUjCIaiTNtrcA6OP3f2V0
8gVXRJlNjX8f3ppUqTqdoPoUQyR+pugWVhpdcckLJCbeDqY7CBvTX4anKiSCljtOkZ6fzEiGmK8j
azChua0oY/PME+fphSEAee79V1YgnFUjSOv2ifQS/WndSbl8VmZbfJ6Wn60SC6Jt+TaPZM/2IuTW
XkHhAa73Bvv++7AzNZ6RTQJocjXkWTafjLmESoMtVazMz3JEJnCJ0M6R6+/JbDZ7TDFJW6lyQ6cu
5jQdag7tXp0b8rDopMFGb8utgOt7EQ6qm8gcGGx0P0zpO/ibXK2UgPZD1tZcnI9YUR1CjOBz4KEz
yl9JD/HZQy0Zj98IPc8de15oTbn+EJkKAbSiDRsd9v1B4OexYCAn4EAvV2CvqXgGUPeYBNGujrt0
RarkdPZF/aqC5fC9KkxjyBLcG397ExL6lr4PrrGJjmDtN799EDYUaR/1YuXTm2sPWe5/N8s7kc7x
7IxLPy3K4luTc2P/5iDvnhcNsExPc5bKFB2TyWapixTaSZeJwc8vnrh+Kc5iXqQyxx6s2wPDfRPH
cIN2ksHrANWRiDooyZGog5Fc0EdCp4vr2TgqzLai1f7BoGumF79GS0eWX9Ed/UiJLnyygLUzzLhb
BeNQhG9iCc+aOBRMgH//VedZvP0KWn1fTWkjZ/e0AHg2U//Qs0pHLqv+t9dreKjVetSIPljbWfrG
deN31XsPiz4mfUwFhrokcMmWhzx7urOf4oIi9c39y3Mgz7Tx5fM4SzxFTXfBhWEgrv85zJn4uxsV
qajirunrKXdB8Hi4ANXzt2l2j1+In4FS9GQEzYrazplbVEODkLOQyRgLULQOSsSjPWrV4/hwMu1J
DeevYDFwd09Owkg6ShzhIz0cVVI3RYlD1+BVYQH9KwHwOIDghArcF7t99e++cn0QhT/NN1N3jcEI
Nr8q/ACrU9dY5xvsaSd0tcjo1sbs8TlAu0uQydYDtVuS/WkOlwmcBlArrwyseF8G/fA5xHSwNwr8
+Il5VVkGc8EvL4QSXdW0aS50tV7CFAIXMbuTVfFRC5ZIOJ/BH7GMIlirp8NSN/F5a/setOrTW02E
ky1NukTuUJM9okP128/DMidHn9kOCydbylCVaz++FsY/5wFTAYBYuEOqCMzuvBFGgKCosdwVwu/v
9h19W01OD9+GyzKLDhH1Sxt2jwccMcIJxkCmTjuozKn+B2742kumRDYEH5RoBPkydI6ZQRSkEAo4
wvymhw7QM8AjaVjNPbZDpsoZYItz1dFE0DOKJsaptno06cAQwQIlxGYf7rOlXcDByd3Uj9uRRNr7
pZ2H8NxyyVhxzE4yPai2QLDEJ5oxtk+T9atliKbal53mSmYgwMKhHgGbkzKm9qdqhMAHKhri6tBY
1VOIk+XOMRsE6vaxPnIr9AL/eBVxNXBBbtAtoq/og6Jak+fAOnBoMmuM0kyyUDuX2A/BsLG5QQWz
T6e6Zyfhr+SrvOQdbUYf1a6Fpco1QzZIpFaS0eP+Ng8Lmm8IqVL/HlyVZezSStMxtkW26I0Du6Qn
cwVnoRM8sT6KIjFxBuk1Fc9h3nNjxzS2WH2ndG7KIfEzSSeVtCIjFsHc28UGQiMU1aRn4Mbo2jq6
cCGHO/rLCDY8zHyENDSyAs4HmqmxbxSznTjOZQTkkzRahqDm2fyHn4qmRtHx1o384grq8mA5b0jG
ofkQFHwtx+C0gEWD7ux2+bkEW9TDOKS2hXZSyWIuYw/gtHZC3ZwkYUrdgJ6kFMHQaq2jvLalOvBD
k+wnF5JCcBFZSa3k4YXj/Mg/18P1PK+bjlcpdSWIzog0tvtNBgH1wKdGricBMbb7sx9e+OhuWV95
WQy10T+mfC6ETThOih+D035rytcHCNWr1io6i9mHTjtjlNY00iBcKP5cmZUL4PKd5qjY2mP7jOJx
vJVw1p9jRtKdx0WDJP41MW04JETFKphflvwR666zZ0uH05OrXVf0sG0xBUKgXD92aaWQlWNVIGyq
XekskJYLpOiyaFjqXHMBOang38dOcBhRKv4BFlTTFhU1JSO095jM4DgQYQljlai2xv2mkgkQnAdG
dnf6TLEzLNnQ7jdoqxnBww6s1DKVjf8PiFNnJSJc3jXIVbRztS0G5oZU+mkFdumbfSGajvAyIp5D
GL/WQCrZKRCnvuJeLC4rmLxvaKC+STye9EGsnbdRfmJDbZ7+GYH8zbYOtvIXtHjyy51XV/iejTR5
IUHwtLq85Loc9SYMDIsWJMpZS/2F141dtrPTo6D3tv7ZCIv9L1J7VnExoeteGyKxkCRFANTIHA+/
oYxGUrRu7H3ts5LxyLQqjvwM5cX/J/oj0L8iOQMnZbaQ2Iw9a5WJYm1d3rncOCj0KgeNHZlHOf1e
/ojzj5/q194pNwjaTJ/s0J2vbN/lopNv2W6vqOIdT7nuIWHfp7/783mpdxzJS783pwHr0HaejQR9
02d5O1/L6kNrinC0ItPdtle0qVy74ha8/u0FW88+wMORpc1RNqqtUK9Yi4Rrt3q7J6Cb4DiLcEwV
/x2Z/xdqTGTdChcF2Afs2V9/U9TRIE0oCxEov9IhlJw/rUoHpUZtwIyuPBpwGZ2MqP9WFSJeszeP
KN++Bn+dALnIh4Tl0BMQXaDSh4m/GVXbSFkmHKRufIfpIsyQlLHnSdkaHIK02Ov7ohOXCpuyaa1t
E5g7mqXDFJl1KQr72/T1PGiaWTHNXN2jNdAilbbcYMmnzBCTXRR39gZCCAvX0mWohzwG+jy7my+R
L7E13lAE1Ez4hvvdjfRgNWt6pfHBwCFv2Gn+8gxsx6vZMU//yN9KObwsYZnOpcPTsGznEua6YPBz
zrkddUpHuRGsUUEgHoiSRgHHOrGEwltD7bqbMiuUTEZzezXRvmlthCQ12I3cD11cUv4wd1y66udf
4zwlltt58GQvaIHGIGdoSLJxYvobUAk/pl95K/zriE903ngS1b6wopN5pSHF6qYOZIDmjckGpxFf
eJjVnH3ljThJfNcDUG+iheRFMZ8xI0PybJ4t88HBrFANhlrAYM1fBCcZfNFHQdHSsccSkbzaNDTk
zB+bX2Q3PaltyIDuRhjIYF4QL8FYb57YawOv84iAPS7F0+xSABXm1X3wAA+W4Buijn7ZK24Bdv32
ehR3LbotU1VdcEFQLJd+uDKF/AVDdXk6MZRFhyPr6q+YTosttsKlq37ZNC6UjvPp3oFGxaHgTzTG
6LGR4rKWg/OIGb3w4/isjUth9ROpfxNuxjE/g2/NnpWTcwkcYsVLFm08JpFfihYWLF5WSuAlLOrv
xWlFUlB3uBaum3KAyA9jS1EVas+hMU4/4cgvxIIdlyb5pw9OcNMl0SXpTO1x7UITqnDuJOY82gUK
OEUSA1i3jX2l8y5VE97zbhxQOAIZdkWn+Iddc9h42FrRKQNys6Ccc/DriEgUjQGCUs9CjE6NLAsN
2hIuXpDjl/Xw7BD82P1xaH2mp+4ENtz9xpXONjp4oIzUUfiYOP/wUXBS5w5YLSzWF8dY2ugAMhdE
yvKhszVPafh8iCgC4dMQIvPua7ytUca59pu7gQoMBhLGVFUu4w30FZUobq3LD9xNlBZt5/Ex5iAU
Y93G1eya2r7uklf6IrAbNIqEF2WRNEWxKdb3vBj9+4jJDHfbs67tVKi60SD2FbmvHBteSdbhStWU
au804Wzz8OkaZ86NkVQqm+YY4Ipze1O41RZkC2xWZv6rIPijnFEOmPFJuOH1DX0lrHEnb936dIDE
1PJs40NaDGBz84gfI/OiX3xUXPA5DaG/LIsvq4R3bG9K8IkB1dbWmaglvJLh6uSTPzmwjNsZAMAf
aCa9dYwmQWOaSVVPGHLTjvAYEptcbesqm5M5iIqHaSZyUtAgLj1slisb5vLFhmMyKLKYENk5I/pH
BOR8ZAhtkJrc9SNhNoKJBaIfzWghQQTEAl9uvMiDmp1xW1JiBad4MdKy+TSMDjXKIYgg1zTOP0Po
0Pi52owK3HvXxGsa+3wf5IxtHlK5GT2dos+hX1s4+365rtULTeaBhjVH4WGFyqSLNTw6wRMHlVHh
Uh28RX32/EAzkSh3c2uDfAMvaCJHRchergcZiXHDoLZvWC95fshzljE/xWdSs7J99lHl3tw9uTCJ
7qUBIKqvs/YJEOQJBjjIGTr/KLKWjQkwk5m2urBXQsYvuOYVQUK9SIJFV25chEnql913E+dAZbvB
M3EL69+fc3/BF64XVb7jtsQ5tGf8PIfQd+/5njTI0abpK58nWhaMxhwfBVSjMU99h8tPdQ5a4fhG
ICQk6Wsd9ddNA1HTDzcZ/9x9OoGGQTQIeOEeSu6h0GJbjBBVv8BDmN6UaUhZECm+zTBK7a6jlJgp
xfOUaS4rIPoW/IhFXEwPNO92zpM2O4pZSNodzZuXsMlasVJO68muk63wtUjie/eyrzEAVuoL6p7e
5bq01OckKY2WxpIc58EydyDhdZnENO1gtc4EvJCvWtbR6CRFyM5bRVyYYlT8hTjj6z/mJxq/6V0t
IR2FNzdKn05mti5m94ybUd0YZLc9sylUhZG8/2prsoiIvmLLQZoWSTymRwqEc9wtYiHNkQkYjjxg
v/XineV3PKIz1OGjyvR3V+A9ewu+FGxYrq2eiOP9H2jysVABengYjh3GHVUoinjw4HaDXfN9qKpQ
Cd0G2xj3GV86bS/zY0zSiCiy22wXgj8dIsZfs6Sp1FRnH+gSqGAs+E534Qlk2n0OSArjclGFAd+F
yRp8TqZ83KpS6p1S0SAZPIasgb1878HPp2Lr5Jt81lKRSEJ0ScUazL7dm+shsqlyPuaARdsB2tMX
GI9lfzVR0zQXzM2kCNbMOhqGnsT6KZZgYqoEpP80LcpI2FXh0ZYXpYQWXRihUFHZGu/7Gs2sGgD2
JxQO1jHF4QAnH4KEwpMAQtB8muX+jHrF2G4y92+tIwHIMvzMOxvO/YYkt6eAggvnUUdb5/23/miI
I7jfPAhv31Bo3hQT0gDnPn4KvQU+OmQc2ERR6kMl1IAnl2VYYcYDKTSMjYFIFTP8L1+uiUM2k3+t
KvWqXCkhHuxCsSb42VdEOS5peq/IsEym3Ulxee7sln357tF072py14Z47Lwec4t+w7d404pjamar
Jys01QMryZiETVE/5vC5eE6C50Sjq6ucAAQpcpoCnlhuA6sNTFqur4HLtdV9L8dA0bbWqBMH06Yw
P14SJmXvJP2RORiCKlAsEHcN14AWOgt/ysxjOMKwpwGVriWdL14R6Isnc0ixLbHmn4ecoiQnTNG8
m6LfzqNCoOAz/yh1Ab10RDVf0N0tleK5rD7BeCy/gy7goQZpotKWMVsO8lePh2kPltR8I2JwQhHD
kBtfzxRgk8i151S1fW83ObhA3m7YUvMqxDwDpGb0QSM9B+g54eiErD4IPxlqnMGQ7CjTyKcshsZw
jfY/OQbqGfZrKB/fHBcfgSw7OjR88Bo/xRC7NNmbA1bmDuqu5tGCwfrP4jjcwwsIRmw1vt3I26N5
J/H4aEebsUB1AdAdiXQRUKulZ1w00EXcNVEk/jTmK+rtOG/f0V//aZgtQke5HCXGR7VJOvCtLRv7
XHEjdcYG2LqHwyhhZWTWdrrhlzUHAbOoPwm0WpHKUcBlchmpaQubCP89p4S80EZRNKBvHLb5/hPh
IrJSVA0FP7WwWjClz0AyIyrpGSBGshkUQrUf3EJF1TbBR1eqJKOyZ1/7RnXpICRVCyhTB2Hy9DVR
MRJNoVvNbbV/aAVgi5kVEhb+A2nUq64FzoduGPIr9qtV9slD7OkZ0yWz9dYrKEggUepJgSvKZdV6
bqNxaNx3PvSexKkAduz++QK+tmkxci4z/5Bvq6P5Iz0XYuWjTM2L4wwYbzqKtFFomrQq2Nfp492T
BueUs1f4NYqiJDlmhGWHowY7nILDajiPnZyOJkHHyCJVcywI41q6f1/LGNWLniOVHTuY/K4d6Vbi
tcWlt9tlLnvUyNiblOb2gc8+S0nchHnlVxOc6Jj4+h5CQtGsKRafARIRvKcfLaP0xvVNr3Jt8A3r
kcfsPc6Zekw8OWAFfBmRdUlqPUZJBmza5MffBYaPevpBAGOUWy2fxn7E/zP5MX241OpnETe9fbnn
h33gwgCd6zIKl3Ak2RDFd5jpuGuttnk9TZcIxMaHLH9gb+4WvySwLN/P7Z78uz4JKPtVv8Vvbrab
e90I6CPaM2fi476kovDkl/jTcCpnxlCZJiJP/M+SKvcMRF6eyhaLBNmeChwcjP8mMMXo6/A9LULB
qdz9LH3EncwdFUYRIZQvome6npV1Jhz9okOBmLXCzUj371nNroZ8of+Q/636/rytML/gn1P8Tfdk
QUw1AH9ttvbZX6NKcBKe0H3M07MHfEDBemhGXQ7bRFoOu11bKKyelzRbH7n6rkErpvQnPhVDUKCK
yjaB/xDDGy7UuWf1T2Mm1gvOr7WasTcMonFmtpgJvn50n8JoWhROBiZwJNj2vJVPzSf/A+fj+iZe
H9GWPADmNN5OcWTSWn5mE5Q3Frn0iC8NillIeeSD6LY1gl0jqVdP9djQYpGNWKPhpvqJu23N7FHw
83TRNEINYJwkwkRZI5T/tDkpS5AKWY0+CIeItqO/n7wdFoU6F1c8xXwtL4xLuWUfT1H130ck8xl9
PQsa2f+paf3X2OmaLdJccl1TnzyBnPpsojozIBn77q2Sb/GDp4p9b79KPy3HZGOtdQK+IRkIA34U
LZB1+vV5OVbUT0xU++U+TkUpa0C40dQTdt2OEshy000ixBg+vyPG+JpwC88pngQz/1WFuCxl4oSn
IFMqcZZETgFWTxgBXhBTiZkn1+nl2c5JtUrd9TN0O+QZtMXImbPIZspnXSTHN5d1h8TpTsaOKuV7
prKBCL2X+4Yekk3a7Fj0CKZaqH+Rk13yAqE4Kf/vz/zykIR4hTaQVnp+Nkwu5n9bX99hfzxn0r9+
os/AivZn8rQ+bBCmqDOXTl1JuE8EoXr8Et4f9GOS9DwVBTrP8roZzbBmSleiw/sw6i8ASdwrsCPY
Hlmpw1EDhNpZnNyoSRTE6YrK539rbkC3U2wdt9eRftmVQbiz7PiIMnwlG9nD7TSTHTbAsNJZVMva
QjcnkY64oNarSZ18Itb5uCiRmmyszonJlx1cy/TihxLH2Qv6b0unT4nfSn39yul/1ZFm2kPKXELb
OIZZ48WHwOUIpGTcqcdxRK4e/QipF575o4k4lOItse5WyiTiyT6HdG2HHutjOPBffvvIBiNX9mQK
05D8VHuoA3tCl/G3Yg+LlQp3s45d17g4gkaEZTxTXTTBsxTsEsdZB4PzgwvFM6IH5mcSyAI7Ufog
PRXD+qmyoQMfNSaAq6pKbmoqhBdN1doOX4cq0R2QiNZnB8piMFLGJLc8zP6+/Cw5JPAjtpASsWeh
t0LQPRCMr0Qo09WAKQSQdKnbHL8X1bV6AXfji7Qz8ujgLmgMKgj8bsxqNWRgbHHFo0X/cVi7aAeX
sXkHKG+pzcyVS5lDj9tr8AgEG2x868PPuKvMXA15q6JHmwDqSuHJgChXry0TasL16RLDHhJ2pshd
08ogKctTUxZ4/0zbJlY39l8qhrJoM8ZsjpkSUjHaMjw6MpfB/oUo/bWI1rpH4RFUptlR2GF0XKdc
HscvBHMvD/ghxxeOPU+8Dz8EfSIUUysW3duUmW7jaqT0fPssIRP5tEaBJwRtkgsQ8iJHd6zwJHW1
wboVdZ9dBvf375Spkna+u8mSgedKbb+JdPJxI/ZhGe6S8r2dQt8KzZoXSyus5NdjOvesy9VpIdKc
8MRsdkOXKSNBVhgzTS+KCikzyNRHgoXjuQVIseewZWgUTtrQyeq0GVmbSNCL2Gwf6R023Yth5GFx
K6MpZaE6eQGXp3/QgFZ+ZX9RX9yFUS9y8CF/SOFaYNsc+bTT7JtvfOSw468Dj1K4yq/JEx73a/Yy
HlK/99fEyhDijASPG92kzxwh0v0R5A/MhvIyoPbOju7i7U/eXSBhz76E0FlBKXguzLP5JQrIRze6
jZCWTaOOWL8KcBXJvJ0L59OxYAe9A4uew2WCTK1XGDENRA2onZqGedNKjinyNCXNWfmLWg/w5OdF
/zwpKYiA83SLMfdWtV0iZsDr508ibxXvTlWCU+4IIIDjWZUH4oF7bk1ybHeRfYakLZdGzpUTTHWK
c9q44t64pTyy3xiYl4YSH2Ojo6tLYrywW+fO3zqdPFapNQM1SC8DHJ63gRVi544oWMxpDkQ2pmmG
u98B7l1FdCoHRFgpp6qxf6Fl4ryQ6g0dInmii9wS5W9Ol0LXZrWLesvEHAylJpdHwAG2AfYi7Aa5
EAOXZ39l0T2hVD5+5EH7jqHjFf4JF8NPKEeqMF8X3HyHUfCMiuhvJ4rps01bSJN7cbqqDE1oltJo
PqLCD6Vb0WRFwTStaB+xAlreujIfB4XlM5StmM9c8JN78wa6qudNV95ByjWTbGKKTjvuwwTUCQHJ
sCI1hQhd2FXa7w+s9VqEFjLgrHJSZQh//M2majKYqC8bApAFzr5eN/ydHSqf2tswOu2PJYnQ24bV
0G0UvUVRLX16ymsnEDHrQadfCfeg7Ws3k77KdZtye+X8UdKLl/a2euiQh9ja9F+hhEVprcOJxV3E
p+Vh8pObbYVX2DLFCF2QkV5enW2xPj3UuGk+Y2GO6UvCUCfDejm6cWceQkEuyqNif2tXRQTJ89/B
CwLd55SHy7w84gXXoH1VN+xM+fVO53oVeNK2tk1C0oawhABZ/sf20JXb9+ivs8eiWo5SWuY3YgRN
QnbjUHK6n4Dp73Qfas3NqkS02ge9GfXYRKmFFY6IFcCoHx5IFI/pzHOfQ6Csq+gUdP6OtI6ugMQm
eZc5RV9xKaj3yLzGv7+uwg2YWWkSjFEhJuoT+XqxP1PtlYjWPUhdh3qN7ZMzFev3cPLYZuR18vgf
wbV8QpZpEHDGaiuban6y6yeA+z7tm52R6EVJvbN6pM0vHrV867NjhCqFh5IK2xXnlAQxke64MwDa
ekBsRE7jZ/cnrAtCLl/1d/31ujPI1jn+tQLayb1+Qj5l7zGoDH4AEuIfa40FES24Wz0IA7VB5r/o
hfpVEHufu6HLdp2pP3WuNZKIs1hWLIpQYjhtW1D8k90hN6v+VFQk1lM45rchM8MK+HHftnrYgekF
NclziNib0yHlf7DoChRjmsH2JzYymPkeWDtiRxv6Dv3IGZSaB4WrWWYoOmV8fcSZNcMo5M7ViRah
+HfNNB4oRurx+C3qgJ5UGikdKShnlFUFnkpdJPy0wrYrvKBnFPVrDEuyqLEt34n8ibX0PhsMfyxW
9ONA/QjMlrG0JlaInwUXTbjOozUDPKgmOr/lJywxRQNpUxlMHWLItiiz5DCi5c30s/AzqfvHH3XV
LhQv0bDyUfewlbmbFEPk+nLokxU114K9s8ZFLtueMG/EFe2H8Tikts8INB6difn+bFzwTDT8ITFl
DssssuwNKR48y+wB+rDMrl04ShbyXbxvHIQW95DmCK52XOMZXwOECKbglHpUUPq7nNiZ6qLKlP5/
/OnoiJD0SD81pFfS9GokEFdaqpEk5rNpyQUQxeHyAHN/qcFiiOwkkpNFhSIU1SjnUnStPfhvPsjd
IQwAMy0e0ydyeyWBFgqWtpXPD+duQJBtAol5MBCZZ8Kiv3Pl0i00keIV4UcKTOy2VlCaaeI8LqjT
zcWrYbcFb00yk1f05ls9OyG65FTzzV8GWRhzt4Dxqr43zo4vjm4OWMjfd2GVtnRNN7an7kD7fZ6x
+S67o99d9Zj/+cxuLJtxwU6MXmqZ0owtuJbWXG91y58EKFdV4zPQ+gQBoHBqmavOxmGJqe6AKIJk
yXbIbnly+gjHUYJenpnoD7rTdWGw4jUt12Dm1pC+St31QtFg2L47KiTD+EPqtQwj/vo9ViR4QIW4
KBsL4VaCZYgjtFrTlHHpVCTdWQgZcWZoWfBgx0pNhIZBlmQF9FSU6nQgklWkcoX1JxlaYdmnZsEd
s51rE3neZF4U5xfYnPv54rzs4cl5+cUwKjVoPJVGujytXkip8sFs4GZGQeb2PPMnFAa/D+dOeBjZ
T+QfDahxlAcrO/Dj5xxfzFOFkQu0PSfwbKVCgDfYIE8KQo7duR6Oop6iEegkmtLIrE7vP1fT2bWy
7m4c30lkfUw2+5qWJuXUw/74WZH5o8wgcpAqCyQ9dUukCIiYlbOUBz2NtOAbBj91Y7eKNAtu5iyN
HLA5UPf+/HTfwhI4648CI+yGRz/mGmXBP1SHYxQHx8OODwSH6SPPYmIVX7uBiZInu1eLjY9FXVwO
z656qK/I+8L2YUOOmOPj/Svo/vaqD7rwlFo/AkpD2CFk9Dq3F9rOCQrZvmrrhqmnfMS8FjDqoLw7
R//Ow2OIzd3PFcUoCdy4hdCG3Bgl8IWAhrrQDrY8SXFEI2fts8xr+z7N8S508OemD2HJIMc/N8du
4CvxLBgECJkHosOmko1OWRb7C+5uUE73HVH4NAwOk4xcpCOiVjwVIxGyLJI0owrCe4OJjNii1zO9
6AgZVv1bhjzcWowDqG3c1csZsZHsY0f89+Kd6zTHlNzO13+IUspCjfM75HjjV9/cbPrQgpVRji8a
CVA6fbGzMev8boViv/P6juJgMtWeDhZFvf0Bmc0WTHyZsYnBD7xBbD6tpkuZgDurThzpT79JezEK
NMnS34F0obXdz/khNvA3sTyNVpP3PwSNkfg8bGzbO/kgmgdM8Z/sMb00b3d/qcrrTltNzW505Tyj
f+1V/y8TbJyFmCmGq2n4m7mfJF5ClYyFqJ45QJGvdO9W6lNZW9xF3oqsMNz/AzKelnKoqvTAyk+y
MwO6FJcYXb/+1nUMZQT/skeyPCdKPHAhiEBcCf0Atqdg4okjS3XZ8Uh17wFf7ZR1ygzNE5wGNdYf
pOfTy2wzq5/YyylLNZTMhjE1KChA6RKl1d4Cjb99z+b1ofrIxYK6qX4dsEIKUYQhMcRwljjEEfKj
ZIZ0/JhvPEVf6FeHLewxSX5AO+JszTL5m4LACGqjIcylTxG3No0gqYMcBiVBaLToTseM/qLHVzHG
sqNwJ/DOR6dDavF7IC/q2FbQS289QZSX113a6Yk3fEftOjYe3YiQkOpLzXJfcrz7kXQBfV6c8yO8
bFjHRaHkYpkvnm7FUHR0uQmK+iVqw3HrOs5StdFzrqC60Y5UhUN+/T6W+4Kjnm7dMNdcCMuc14r5
zkkZ1BReHL5bJu3gWAmxvngS8UHkXQUyNDPrDWM2bPyx/xIOR/CK1WcMW6ZMte+TV1QZR8S5cL1H
3lAoOkY+5ztdzGvE6Ng65jWnxapkFC990IzM7rHTRnkB4um3z/2VCbsvwbeN/WibBGg/oaAlCpAR
H0RxPBoad8l1PFMVVnKzjyJXdmoPtYp0g+bjcwZizyYxDy/C/sazHA2zAOgiID7A2/BkhDE1/X9P
LTLQpMi9J8gHNOdSLHk9haDyKi5H97R7ZYlV6RiWZniAtZKTnRRyqw0mA5yp+I4iRuCorY/nfwKm
ELIox0gEOdYUCzxLxkKEVLx37a7r41JHbMCLGMi4vXvQMqVc2vgK/JaOlfRAO0HGYIrBM4wDJd22
H1x1duqO+0C754a/noF8L5FRjS2WdQzsTZK6HmgtUIx+weRxjOTlbIvp9E5LrLq+H2rMhfusnlb7
36nLZ6wLZgRwYw4hSoglERQAyQvPI+xFojTKM5xpKjmFA/98OMkXnzQ3M0i0Jdk6DXu+EbCR4Hs9
LTjoKA/I8tltKp4ZjYaUXkg/wEQf7GxuL0QEcAXX7vCIHcHnOUUm62xLwn4FcCVtEylbrwrBMWUN
umac4dtXeyO27xoVEHPOXEhfNGaF/x4TUZj+s+oxAHrmIb/K4LMvpM/UAXA6uH3HSmpKwkFUNb37
9bUBjHtuL4D9jrTSDqiiNM7IpjUfs/MkcpXgZKzEQCsCmszE2F39bHn5jh+ekYUl5jfD3LkSF5Kq
AyJKamaY5lt84Hva45/pUkARp/eJE+rKZx9E63Mxp574kwnivr+2aguL30pwvvrQJUu5G8uC+mEr
cRqI6NVsCwVSLltFiI8GxETjVyXLdI0KrHBzMT41pXEZk3+JccyoQ7IUna1GytWeD2g2MjLEgpra
tAW30eON1wQzh/5gmHPqiH3JWaWtAD0JvQVvzu8higJA9JdwJVbtU0crtFK0f8q30zEyBVmyXZzr
k1ytwn6GYrMGrkT/DpdmnRfrONjlUvLNNRAi0Lq9vE0W4XK9oiNmlOhCGxSdeBJu4siZFvRjSURv
FEcCoDFt64o9HsoLWHtyQCecflZjK/UzxPXQkqLh8GsNiJDtW4OMtJiTSQrt6i8wmUnaR2CPdNZx
EipODxhdXsBWe/F4h/u4VC5hDEMyJyME/TstF/arJhrNgxWvGvoWnGgeJdTALpytLckEW87nUPt5
LroxAqvoOqoyunPVzyJiu35JuUn6VZFouPcfmy+c95eLYYhSly90r51QomPQTKAP9ho4I3krFinX
IIL8ztUmorgl0B+l1bWnkQdbkxBx/kmc2kyFzvH1TLgjCghkWOMp0znIOzm7ycMRpyHR/4gfbMkr
VzZlRCT58RfaT7EeCgUhf/r2DKHoxMh6QBW/vZtVECIOnKY4qKPk2t3OyuC4XB5w/7N5VdI8kZoB
F07wxjZzG3Thcf3aCqe5oPAayIQ+mUYjq2gCMiv2X3DBt95c8RbJ1So9v8z/j51OEF4uoaPLH1Y+
Ck9rtFhEPN6FUnE05mjhtksQsXxeFNS3JAaHvYqAihddXnWpbfHL6/8zy8DDbEKx5ZQHNPI4W70q
9YlAiQPimPC7eLfpJXCKH717MmwLH14zMWTLawiTU9cN+BmsIn2JU1Eoyw9GrfBzcQwo6Hz/pZrF
SKjHmd6lF3u7XChuIy7B370wL5V94JeVlz1H8BNCBBd0Bf4EHcUxtgB8eM+lA+0IplS9oFPxXnnr
cZ0OcAyFpeF67NtPcqtVYyvzUaFs7MWXzFrgKFWckuYVC9OZH4O0lSekiLNt5aIfFrvcYY2xRls3
EwWZNhKuvSSWsrcr9KxEv5BqfCpUtJ05Qvb2RPfmVwqwvayxp4ALYvJbESrmzRJf7W97e/CPvExA
CWYp08QiOSqBPhLmXAI7k1NEpDrDeSpuP75Us8gwq3TYeSwkxkVqOOvacDh8rNQVgq4gQX3lzbr9
fjg20gLA+t1G4pWjlIaX0nt+rOWmBCL05PG9BkYW0lArygkFg5o3ywZ8afbfp/sjvmJ2xIwkRBfq
O4NCyVWSLoF9Q4d0EjOL4UVreEk6LFMOI5wUn8xSfP7gcXdBhtPTeKuwyvRlSPdZhhtEO2eYT6FY
fY+XSZg8THBNUyoFjbym/07Z3Ete++TXe9O4USYGgA2GIDu8RFR1pRutNbRzQbCQPkh4nDhcOXCF
Nk5xwanCAMdSMvwLRAQKhgg3ETSd2q0fzx+Rw5LspHshB1Sw3745lozqaOXIQjEXwfgIN2+MERr+
Qu5MvhhtZkAdFpBS+mZyPxoERLsm9CKJ+s0Jr31RYfmfmrJWo9njWyZFMn+hINdO922FGhL9tzC5
AwovhOA3wEisOgPxUdd6E5o0KaUnaLx7LalaTGXlO+9piUlt1r7qH86evdmkA4Vr0uxu0lhUNbK1
kqeQBo0PJAJD7YCXlJSfC+neSlj5G0APoLIYzIzwsZCpzjjxQ2thIO2AEm7dH/+90BmA6/95KwJq
WdUxdnM7gP4S1CjubwZBFm7SZsvcDbuM7U1pvbkpmQKB/iCo0ffMlTrImpju1NmzLx6nZYrqX5v4
hQE16XSVmqdLvpdTIZMyfHnnI+ZqG6AdH8FBWZfHmwQf4aBXISovSCtSWLUV4ikNkYFsWhG3MeoD
8j1rY+9hckUHURW1C5/9d4jZjaiacmADQ0SYaPh0Vw/h9hCn9pkgpceUIQ9mdjPxO/XQDWWYjPro
LwWbJEPSJqF8rWd0KUeKLWQdu6NHNLED9lWkVOr69/73M9RI02l3TaKlf+gOmpY0/fFbql8gPQDA
xWAtHDSYLfNYOz2C6YWYhES+SoOLpeam1v4FRIWws4cfR3gmiK2tsl95WU7z4sCUUkdvAKQZRPFo
O1zMKLmpTlrxrjk9bjNmuf4tWfhxkPvHp3BLF8uFpNFaJDD4cJr3CALP62dJucqeIC+AwUQWOCRG
6gmeQz9loKB+NGPeSwca5F41DQooJHq2gp5sAG1ojwL/ekY71YPNbMwzFGYzhnV16wtx5GC5mV4w
0rpPakHj+KKaXere5lmmegQWbg1c4Uohn1bLcTtQvJaUMAH7yPYF2ST+h+YkK5lM6k2uoiUCCSTg
gpprOd+oyULeIcrzmOY+1J/vEbcm0fRB1l/jbWOmx8t4UyWfvI0pb2rHG0WHDVN8Pe7EfY8wFTCW
NKBtGV4tJSQEe+bWlAHq15UgiZLoQ6lkjoOYn4DAfxsUlsuBiZ8sm6GrayOHLmM2Jxkhid5/HuRp
QrQ0ahbWAqOuatt7rrVLkaRBb+fHW1PvrCnjajxxUjdDYphlzLyGdFZhyn9LB5U42dYx/RFSda2t
VHJYazJzLWXhVZ7qORDrxDxr04n17y1qTVksnaGT81ppyYzgxZ0EUsrY014OldPsUUefT0IVAQXy
8FizSXFBxPQLxAfO/1q/EJVdvJFY26wavmiISrTTDiXaJnUtzfeEDPEB5CLOHsdpdtBNTm2MFhoB
ggygucKg1B69g4SJv64A002Ebgr7EOCXqyxgyNJoNUCSeWmvixXMmkywIqU0Iop3xERqMaWm5anl
spuqCjGs4G2sC4KwQqL7++7mAPG22MRgWz22lzabjmM+KIl7kuXoLl2dLHaQ1uiDgYOSehNiQFlV
xB6AGRAkjCJvsb/zU62K7SeVn0f/X8v0eO9KQqw4jGddlPPC68ysLZHLa6yAX+Yr/x9X4rMs3FMb
yVS2WxhR0aCO8N3D+O/K5GMYsJtSjTHzwcCw1hd/Aj8FUrFcKsQtDMqp3whCaj2Hz3fExaTpl6xm
cvplLcfxoqM6F6LIUHkOHLH3O2QbKcPTn/2LaR4i1izAX+6uxcFT3E/sk8pefOt4+OJ2DfSVyCvn
zgVQvxP5cckFXBvkpH7XwSkIcr7UQka6k/e8w8+0GQyHr71ukhVsXrObC90mtNAu9eP/BQRGu59F
hbDnCzhtis8mXBKCDbHoG58kZYzh/KFa4DeUWSG4vK35bQXgHmayaKQ/WJQHzWLIAdytrpea03rR
kc64/rrkfPo9EtM8HCxZ55WuwwYjeFzOdvWdX3SQ0pHkRcypHmkW579jT+AP5+hsgbiHbaFzDjAj
hGvYm//2EHf5r7dtOLCOKGQE9POwdSFCbrX4z+r62n0GeykRFzZHnDZzOzM2EHCqbwNs3sqPJhUF
nF48cT8pBGa1IAYWrDFvyh/ZiCWPLKwisXtI+rSFflQ0F1sm5zjMwhGfjxiEmqUnNkVraSH6UIM8
jmgWnepzIcrk2g8rnSV7zP94FPdSu2H7SBd96Bsb/EDC4Zdj7FyvvO1dppB5VOfNLpmP9nmyqG1+
0cKuIgSaYmqHBCI2hpPSyJIcOFSsvDD9q13ZcaxW3sqze6wjhZ9biQtmEsifl5YuVbq5LuO9aTQo
vERxebEzBs2WJFgnf1BBplQvZEuNrveyfCMcqK0Yxr1eB/3Uv0c6SnMj0/5Vqx42MgxVDRK+J2gD
1YBDW+xF3zYI1GhxuzdAP9bwfh8rbts/yUtrRjwqUXwiT1s6rVjE/LhZN+M5Vkf48uEa8Mb1J2UB
iu3zC3QJMz69TkHPTBKvMAoPSXKWGFAo7/Rvqoy0LLDXO6hMV/7S5MI3U0BazuSyR51fndqmBnhF
kc9qczO7NckD/XkLW9MZ5LgJaJP6vagf1K8nCOt9PFsJpjjhmxvK4ZPuJC92+sqvu4fRGhRRHq29
1jXlJbbz03lwC/SSgYH3vUG4yuFpp2+dBW2w1Jh55DY5IQIrKm4KFPMxnlipas7KBozid0/LrwvR
eJceAe7sBr8vmF07n78l9MUbvXM8f5MZHgcD5IGNoaXMrEIQcKCZY5SzNZNiLHkdElgW0gh4CLZ6
KQxJW/wQwLIkagJricWwLS+diDoDxE3wOllVSq8RsBU6kOALq7FGu/5aJRTAZhfo3kFo8/9aPfGP
hyz4AgclJBrYDkgM/emfwpwjW+fiJutPLO4ZotaaaXCgZfLBLQhxyN/8ZDkDf7VWKntmeu3LbvE+
WnqLZ0w2aRpbQgzc2qt68hOYMHcDcNELIEX81VhKJTC+wZuxpMOhkUMfwjwvX2eoc9Dvj4PBWjD/
+NowwVRUZsS2s57ynu63Srhz6W/jJ/QXTipBzeDr8sVATT5LWWyN77A/BOBWKU+GfDd5Z1achkGz
NGJFwi8lnBoElWXEql0xVGWmMJTcSoqH4J2/q1rkq9/SA7ao43PGRVYix4ck77pzVrdxCLpnJvOu
4QhXwyWCqm9m6ponoZ6Lx6HfQ0vtYMEJsq6s2Tgqku+HZ57BJ9BRotJAYZvspCC0aZqoynwKLKei
SFI/feX39umvKWvr7kglLjYykUoLUd/lN1Pcx3AGG//qo/qA9r3LBw9xXc6n0JNKk7Xx2R2Z8X1h
ydq1lUFPPqWaj1h3R8/XlBpXJsl/TpG1G/K5/DTuhCmJuGDfiFxtR3WQmfI2jDsL5DzRSvJzNT3m
5iEoMf0nH8iVcxUglSQyMSWdepx5PYPpRLTeTeVxeHNKFNHrOkEqUE1993FV1hisYvm4uXRrujYH
RfZvYaAygpWrwnAjn+/oQHJrILPpPNwioZikuoBxTvXcR56IPmOasbIbblD7U3uT5U4VwpFKoiyT
IrskN5BfEqwQR/UP0qm0xP8LfHXntuNsS7KY3EsU510w/DAuCb0HTLKSE52WDY2Kaa4CJ/pQhMGv
dTYrqPwjOW45l6AmQLh4I4jdgZF6RKtbjSBiOydbBIfmayDjKS8PSxPgMKJ56Ptre20Swj/s4HIf
QFSQo7UFkXxl91AFf0+wpTboyD1ASlo2XEG8tG0Ed4spBn8kAuNIp//ghK1qhyNt0N/OoB1+iTLR
IIyeTxcYglZdai8F8tDbJNWm2IRzYojK02z5asdKcU1LlZOAIN4OL6w3X1avanGg4UVxT6e1S7az
/CF5OkXTQO66n3BnwKuUFThpM61lyNUzi9m8WVav2WtFJvh1cLYOlpmk1U9GvSQU9itHJ0r9zX3o
nR6M4LA8vNZvmEKDI08LdFe3WbAz42GWAfj+AvBWm7bZq6xQdJqpmLd7041fWSire8/OCuLF29GT
xR/lJZ+bjrbkfphDc2hifDMwHSgBjnk2bR8KkIMSx7kbB9FAzxvRRqclfmn96fTEPiF0/HDqvxn5
fNH0vBUhY0alzAYrcJvId/0nemmDi9PuPW9hJXWF1vOP+8SLnaZ0Qs1fmgf6Geu6IGnQelsD9rrD
TZSIP8BYGel4ZF7cah1ge1WC43qbQnaj8kFNal9ktCB3VdnqmRxd8vw69Q/xhDSp9qkAyNjkc/90
FePEN0EzicdI2T3O5WXTFqgiK7rRgVygkTG2d5phmGzLqHEjgqoNku9X6PPq4KzbC9o+/DaQfm+i
Pe1xHixrdTHS2RLDbz8F+7FGxYhh+c1H7nk2MgwR5B/FPdU/YJOI+MR2pz8hk6dZjB9iCuU6FM2G
1RfV8mLIoyySVGyY/DaR/fyg0haEUt+JOpZ5XEQxTph3kPDETL4CTd5cRxNKkD1r8wst4LDUlbIZ
2+q26mrPYMl6niVuGHdRgMFPAtWfiTqczneZUsh7ra7U+ZykMFGOslN7Xy7zWScZE63kg1W1piHk
cvzwHRHGIh9UWV1/OqBNQKFMht4QjXXaAXnVKNvHhU451yMOmkWYBr4Z6t6RDXblaGhTN/bQCvEh
Cite0cRwn0pdKxybzex+abQAHd+dEHazCVU5Uz86fMIyOcakVhIufOCpkxpKPNqpsr6FMpOjuiA0
/3mvmsTCrhZ24MRHjDtOlu1s1Qzij7nrwzDW0/WF0vkketuNKZZ8m31P3myN7VtFpAG0x90vfcnp
sLvCIscKWC1JNDhwfFia8oyltdpxC74JwZ8m8TRGXDycbo2X8KHcjMAohbxpTTFpkrdxB51BYCGZ
yt0TVwkqWzVuTsP0M1gvW709g42SqQiNEYzTG4PJCug3xchwXX3uWCS8CpJj8WwXYEzdtnuL4gpl
4G8/oGdrOeNuaF4FYXVTAT9hKv4emNEfOT5r0rnTC29J1uKFqFB/fgkW+2uQg7ZBxdGNaKv0yl9a
RKavIT5kNe+x3BnKe1sNxbgecRBk2eoqGxjSMWtKj2KYnJ/+HqFn4fDagG87uy5K3krcog0I80p5
oTrrDnBQQXYCLEyxfS9dFOFN7X1dXwHNPUAgxQ1sWQrUUPc6BHqO6lB4rjCLM+V3vhlrG6LecK8b
DlUWiLo+pz0icS55sbRfmJzwTJF0yIxzPHOafzX+Chp/lC7DqtLtPnnoHdbhZhZljUoKCv1ZCtel
YXI1ka5OeI3/WmCBP7KcNTTZPSxidC6Hin2XkEPE5bbfginY19s6SN9biDadCMQIGv69TXoHkkjm
U3uSxrVNjw0CYneJqLDriTCXsf7iEL2QoXANtR2Wi4KViV3JqLAcUGvdz7NkjtUOhUnKG/JmnDEF
pO2NGyYwTr77HoFDxYnHhSAA3hNefI4YhL0XK0ew1ekUVEUxtH6EQ4e9xJY2uGiSOFiBWB1tyWsU
z/RnleYBV1hvCpw94RFCAWaFuTvAZMsSqVlOuKTPZx8FuQGwb0pCd4DoStwVlbGIj0fbfrB4HLZ5
nS+w4mkIQvV01P3WggmkoNOwnk7Bb0yobeI2N7QjEh3944bAEvFWQUFA0iRaDkUuFN6TRUIj7Z/w
LyYYhuugVVW2MV3Q0Db6CbAc4VEQOED8N9N4MzYfOw8Z/nxWPTNfFi9CAn8Ins08DZmITzsiLxCn
WZp9npxIQNsKPrgbDCf0fBTqxfQoiqfaHV7kyJSG1sBMx4GmVnwrC03tnlHervH1o4zX4T01opRq
VtykLXdD3RYBO+9ijUrmUBa+/XMiXX3QN8YUwkdaiqb32/lq62hyZZ73hGNI8y6gsb5vuz7AFFsI
KiaDsK6TI4i+rSq8z09YtlJXRPaPSAon5DfdFhzpmqJFuaWr+WgYFHZzjF2EDeEOVTKTNyr5bBaG
/iWgQrKSe2MGUsCx1MLJsoyymsB8C0hORlLRB1FDzuzWE9WpZzaJLiS/eugy1v06KL/YRRUMW8o9
v47HYuBhcV01KGttaf/1ST3XOFmJ+gY81u/D3U9p+eT4irXjpKjywhzbKS/zSYmwHirDDdhxhddN
weDtVTs9oOXY51/GiLFLEWJZ/6yfQZXjnq1USi0xpS1S6ExzkvpCYTmBKdnNYP4Zx0vBOm9XGAm4
sHbWZ5MBXNhYsti+Nhqad4leOD0b0+gb9HZXntgPzBgyXvgQ+zo6vuw+JZpB3zsLn3voUjbicDx/
4OjxvjCL5EeJZTvvl8504kKUR6mNCiogtnSAMS22plxtCnsMUaxBAP5ASIMNZ9go8uSliBjndyP2
gaRCk8TxWqRo5cQ0UwV+cdNYhhdGMspRAN6wI8PfiPCjwwnx6ZgSkEtHvcSDYDhvD8NBEjpOMHL1
HZbSvAvDaNnS5h0/C81EQorhWizblTao4V8xl05UOXyh0gmAORKo4jTGd2ttWNml8Kj749z+KDg3
1CAQ082xjI/iXnL53YKKffd2vwrG4MiOBJaHJnYSPVZONeUiNbCab2AD+rI9xT8mJcPudlm1S3Xs
+a9n5kqrEH4bj9R6pM9CTFuxBewVfWTWWWZz+u3Esv0lYkzUCazsv+WjhKOXz+wSYM7gAOjaX6cc
yJ5h/9g7ezGnmPsiQmOtAjevtvJLeI5e3b2HFfeovyldbocSmA7wqiDV5J746r2jYtGFX4gcap5h
OmS9yiUrvabeuk/Xni4QpLQbXsLTYAgU7jHLE4BbJj2OTWVIa/1Z7M4O17WDUccrPQMbDYXq2zyd
9a3/wJldLzEaOk46BnIQRhu+aHefHj6c3IaCiJwOUmpZwdnstu8Bb1NyrWiyGD5xX3OlBEkFQ5jW
85OvUs3LAbODqyOLgBRGJG3m4SV7/ey3bJXut5CFvF0dvwIW8KX3yrs3ORnxbTM1doR7D4sklDKP
0MkiA53+eQLtNT57xPZhTSdgkbgPoPQ84xJ4E+rxSk/8GfAi1/pThfEts7l8+QKikD6QrH/REEd+
J2qVkAY0wLer9QTX+r8mL0l1uc1OCWNo8jMx/wDD/ybvqUuQTeP+HwF1HJGzg1Hbhn2avB0TMYZI
5DEe4G/8Dp5AXIDmWs/mXRJwK3wMtBUSf1cDfTKznBJi7GU1Lpvt5ssVmy/tYN7EgH8u+5usWv6z
wYNsDStin9/X60WzjWJ6DGrHKIC405m+EJ0Ojw5tdB3WY28C9qHQuIo9bBb+fSa/0whqtjscH8Rv
VBBFXv4hUcDilBcyOnq+uQO3OwuoOsdAS1+qbnaTmk9ikFqeFzf+Wse9WZk9CAryWD5RIGzoWusb
+GiqyfCK1LHFtIyfiFZAinu+DxTYAWWcJnH+wVukiLo3fj77q7YZDrBKtdzML7J+2gMqGvYtLKkl
XckO3IJfAj2ztJBsxgQYaKzixRwO2jTxHnUmMc+D4L38UKeCMRsCP01FPyrCfd5vWD+9tjOVkR1M
M/dQ3kJJkZJ2Sx5T16ttapjWK4PpcuHrvEkMP8L349aASj1bvHKKTvejtW8ii/JUj5Wmo0V12mw1
Q9+twlBePJjDCjattcEuYa27HNSvEtfv6yeNOUKexBsANbEoDm7B0jbGMXSs5cwiWBYRv22tbyc5
DrYa1Z1YPeh6D6F+ZFBeDIYSMg8agMhPSZNVEz2wjGkY4RffdWbLSaBRtGQyYd1LsnF8TejfiRZJ
UXzKBpsSeHExsr4pJ1PsfqC/fCjCg0X88OMoBVNhg+qk2zJFzu9MtMcuKmfLadvPNmxAgp6yco3D
VkIn5uPePkeZIl665GHa3BOFdYZl4ME6h/ZSX8NK2K8NnQwe4SV6eGCAi4gLIXiaZOl3i7R5Je9w
MB2bXbjAgGavjTcZ88xHDXdnkhLP1BVfpN6yRfOU/32ngcDM1Mx87VeETtDqN/ta2XD8OZuOviDE
T982NqQgqTtkZmINYCITVdRuyXqkA6D5hNTe+IJoB64laJOsg2bEWKG8WkYout75DUT3NVGZ/wp8
6rvm9iyFYmya4keTVpXIDP/GEtGQQRz8DuC41yfSw8hRZ58LVgH0aExiTXPfVqrf2Sp52Tey9JZS
4zgqGG/9lPc3x8ie13264Nj09Cfvlpd/A9qAlqT8qjzggR/J+8U45e268oYJO94ZTtlkEMW1kqLV
R5EGxOr8LXdLw+syAWmkO8A2I3jQWHpAGidp8pNoDHBXyIV+m8OsvNF4Tng/l1uqW7gvetqn7AgQ
va82/5xtY7VJw5fkIjRKQfAg5Db/Bbc8h7xyc6/Ylgv0zpVe/ESQ5YJwPLKlPZ11WDNhjciAK65Z
PlAPC0lA2Htfy2oaRE75plDDXyGU4KncQMzyMiVJpPaaHeaIKeZ9XkM6dAwmFFwb+kbQVH0KUSZQ
4SzJYSsj5VwILR76i9M7LvFcwcD/1pdPLKF/AYoj+uFhDOZpsXlFs0mAuqXe3ZL1gtJUw0RildHv
pVSBTlCdt3g/zY5XM0jSNS59iNYWW2Qyh73tOwGHP+++Ad2kgJjuN5eSqgYFyo0jRp294nuxU0bz
VO8oClW0hOW6LsP1k8OYpYudOf1RdQFoS5PcpsUQrKeFID39fIYFCHpxmrdtHJxK8ZMm13Dqc3uv
8BXZm8kMpJicMfVn0K83+edSq0+HNomPVGRgeDSwlZsgknNJcJw081YKJx0ymqiwU15q3e62PeZD
qGvsNT7lotU8xTjeVuBswm2LaFx1RpyX3VYQ9G08irBuazj0UTvRw7C08k8N5vN6n0x2JrCjaTOo
QItX9w7E5kQa+/1iqs2xRxCbmDTR1z4cR8q0G53cianc6Euk+l9Pz+5NMkHVpE5dqvIh8NGgT5g5
ImAQD7+mfJ+peDi6ec7DpbrENY4ZAGnFkVh5dlZeVTHd9+n3IjTNSOySIxNYlR4Bd/8lcmjbSh9x
tURTFeWAZ9y1ohhszttQDyPdb9ySMVGl6ii0+qYRfENm8jH8JctKTrETfqbZz71QKFN3U8wNqJHd
aq+5ofVUhBtmYDDtcjm6zp9SxbilTez/Qp58+eTsDPdEUv/Q9NKyLZ/2i55UHDUyGy4t7P4m2hee
Kw9SUqpM/JO3iBQU6nhjQaKn/0sZcIIWzxp3DARfbeb3VxzMtPHrmcxY7sDzsIDj6Z5xKVbkJkgo
8i4n72RaQJJ2cwBL+yA/y+vSCdJKkzgzkmxzsHIpuEyjx5S3b3uSjW8fDfFGs5BqazJarXF3exGv
7TKgWVerBlSvcQOxRXYnMemlwmDc2imDfJiUIZRBE0AiBdWZjuufBkLdSivT+7TJVxbE0Im1hHWt
AUVwCVGkVy6lhMCpooZg9kp2k9hP8YD/9+SmTiELyHj8Q7rB6ly1teO1Yfc6siiN2RisTQmNtSmb
xy1PMGXoFucImrAGDOYtZay8OFpXq4u3fRP2isz5xgxdTDaw0gdH8XhOt64fnD64bDEcDXa3D4Ls
IIM5i7rJjR4nr1XNR1edd1c+RXwmLw+Pr8fiVnUzdQ9khuznWyyR6yHK8lPecsTgbP8rBN17q5Qc
4VXhtlSbPjC+HKMzy7xkKxPQQO1PlwSzgYgpCIRkZUNmEY1veDLBtio945WsAxHQ7osGSXxttEQ6
KZk+mGaWJUbCsEKj3W/UI62PCBZRN6LGfrmpAT3A+Igsc2jcSiTCjW3lEM6eFYrsxLRYwAlpuCnc
T5A6VWLU82CkwgQ6qj40xWOZkyFdyWpeufZziS7ENXSvC96rV30+aAvRfgflW0EoiRecOXsa4M37
k/b6pAnib9iSgstYQKj4Vn7ypU1QjyBtAEujBs8F8kJc6ZE5DyIxp0JEMdnCGRaUeWR+HRnaZJEq
aELlLzjfkQkGXyczufRPHszha7zF+kjE9bdu8WOCZqaIloHHWbq5c3KDjXLLt8Dox/uA1jhkCiD4
OjMTeH2Z784K9I1vYNzpcyg7veJQe8eC0XhdxfQL7X7s2lGviZx7ahvXSijrXB4VY/cK4ClYQNwY
yGiYRlUC0qT/QJZht49v2v+obEYwo1zAtF4zldfhkX+fe635S+Ptmz88OGQ1aZ2D3m4TPuGcEsKW
xM4hLJQe+dTGTk23qC6ozYK6qNUT/H3ObXEXi7/C9jHCWZs00JExHzTyzZMiE8ITRv82Ndrh6YHf
bcYjDOoZJVddu/6bmsbDuavWQMHMrS4FaB53cTnYlbLEsFtoEK+PX3mNlCdB9pY19z45EBqT37LS
6VTJZaHDgw0bPOswma6pAyYH+rgcouRNwnrAC6f6JSHBslbr4XC4RzIL/M32ucdr0d914vlWpigS
3bECedj8/XDSHGtfArAyPOSQnA1jCJ4E4TWL/m8oIUOkpPdAggUQLxmQcq9+/FfRy3YZZajAWMrM
N2Mwg2vcUR/8s+AVo9eOvl8fLJOZH0exKP/lDggZMBa1RoeDe0M1Wp90bitdQ70GQdf9+Dyctnpf
wB9DKbj/upjI6kkJwAeH77bzqTeOrefNZ8BuwhVW+QaxeOrXO3ocqeGvwn5z4LuZ4wCW7N9EnuaF
a1n5D5C0hcgXGT4kxwhw3/vbFm2EOx5M5Qspb0NlIKiR0h3F2XTEbJ+K5mhhCwi4lDfp/USfDrm7
ddKhNC3vFmZhwyYtpe880wkUUOoIgwPePf44mydpfZIkeAHRgs3+87cy9xNWECWdgY7kgs4iR8Wh
iZIVCFmA9xWao2AHT+CHMzRP+4fU2KQ4YKv8lVsRHqWnKWRZo+F7mur4VOjVe2spAUsQSMC+wdh2
ZpeeUEHDd5vpP5PhN3/qR4D4ecyC/RAt6aAdrffQMLicFugkXdCbt6QkEOwBqyQT2L3msWyUqN1a
6F5sEfHIVt5l1I5VY5R3PNVj2o3UN7aePvcCZ72L40xo3K7B4Ksk+yv2LbR2TMBIfvfzsYoHeAeQ
7dReCoYvETRizXTffEk9saeqEWiSdwn48dJwZcIfop9k9qhnLDKcdj13QWkUN9yhk814snWi4buH
bwAElerPIImCZmYipbIOMNNVEgbLhfwvPJOQl3MHOkyNXi/sJRqQSgnQP0dU9Nt2Dd9H7yWsJUyR
N2W8jBD8q2TQCAOijVfxG2O/KLPYn23FujhpC1GKzjLkk4GyqC/jyy6RJiuQN2rfMSq5LoyRLDqi
1Ve6eo6SnqPlt57kAFWxhYVY0ayn0lH7fSQ1sxnn5PsNMUhAmVuAvjE83ry9yirynTbU/3RuWJs9
e1dKmyGwXwr/xrP7mFOU1BPkOKK3EteePPZ791YPODsqLp0ZwCGHH0vtQwPj9y4lgP3xNFate307
IYOP5/2eztCnloKv7STe7WOmcetpgzHYm0rTLCSQ3w5WPgur74ERMR/XAVQwaip5qKVgF8Uw8t5h
pGAkhGt7mT9AkTw/bSg06zX7iZCwz6hkQO/v5Fqaq6FinqOb94zzF/HWD6eUH1c3zvdlqrU3prCk
4fq/aBVoINRif72/me1HTdvDXDF8DjGbJyRspj2/FVOp2vCHkMlMK0zw6R+BThUw7E2eJHOnIGYn
GPonmqrnp7UtSafQV99+bmYPccTL4WXMmePtEY4YgVaIAl6KIFbbenpc8KnUzbq21C/YFqfDKl8p
mHVxVRwHmUpJtgEyIXqB6VkWXiHcI59BbESgk2j2JCFBx//cXj7jhzDbm/vZdmrPeeP3pfTSHECJ
xTp2pMRin7F/q52SJyJB2xqm0nuDK49km84e3z5sGp83vrqhURxdHybgYIXq+LeL8u7aeIS1WoB5
96uxI+ojI5IoYxu2fmXjWeWexj3d51F4inOfw9UFJZB9Up1uGhy8M/BudKR9LnKQnulHPd7CRxOZ
jlgTKelqw0uD8CeCCxMRCOqfi8RVTvbryjiIvOhYP2v0goeeawZMUnnoEgvWgco9gBqGvoWasx2W
UbOh6zBYUyMrdY+5CPH/wFTdJam5akCqGtkEA8EZdsnyYJ2MfM57R8llpplN6gLdIOxyL2PziAxB
1PA6GCMWVG0pKM7iIqrl/qC7PTpadrFjG8t/SyPRgEJ7UeZs9HaD2SO1xYchQJK/mtImPPtVyhpV
RI1PlCgrHuspUExl11s1yUKf2eNihZZCEDVKHprzliw/96MIG5635TWgazE2QqbokTXSDGFWodJL
LTW9T+2Qc3+99ukntyia75VIdWWN9v5bLbyuDTadpK8UgS4OA+4PZALWqDI/GMC1N69eBG+aeBBe
0KAr46OpsEIZwMtg0r14LjvhhLw3bjnFvv7LKB64/+NExmcGf10lP/myBMDbML6Qq2tRMnJJPzpO
aemWE9EWRApdcf9k0lVFIuOD9lVskgcmOFVSWyVy8+wnGBon5qWxT/5AJQe3YMUNR9/2WOEg9CY1
CVr4FPXWSrzlGm4TtgvRcvr6yVEeNgJZQFlPkxPPZbLHOWbQ/84hSCkDrlqnyf/sY/nM8TCxxDTd
omlVigoClUnAAucNMk4jCJwb8gZ/JiHN6LpybLbK7qugJl7auCaYhpzAHOOCC46zNMMOTe3tgb5Y
Q6Jz21pzwwWFGhK3iRzXY20ztuqS1kr0I0azuztp03IOHk330aviWoGSwF72jHeRMr/ex7VIe3TY
J94Y+ejhXIDW+v/JjmpsHhWaMDXw46a4zI7Q/yRFxOZFJHC0V9Kc1w7KJl/wY4xyg2N2rd1RU44h
Ck9o/6oYkNMZwQqmC5SRJeebOf0ld6DiZV8pi4NkzU9W89cmLOhmPAU3bfkWcC/GaulziMZP8LS1
T6ZsJQ0JulB/psKzEly6BFuPdVYHCOo2K+cBGFWcuvNzTIlQiK5TyU2UabDpkp39fTJKhU3FZyH5
y/6Y6Oy14xfxSD2h6IIFOOfNvch67idjOo8ClbvsBkLykNtmpNghgsxqLT7VqMSJnD+FVPQ/GdVJ
XmUzAkN8FDASB+i6SMukhSoOjn34ge/ElYchXCcWVGT9CK6ceHS4fGmwEVNYLR8/pAsZRycGcNkY
xochCCZbpGH9lzLRzJea6QxE2wuVR0hmHYSmK+L8BmuMferSK3xRC4bkgUuhmNN/EXg00mLU2OL3
jCTWdnBmDNjKfhUlyHEYCKfzcdF+2pKm6KtN+okAwhbpj/O69qkIe5MSY/rXVwaMeo1l+C1ylI8O
gszCVQ3Rt4iejYP+Wd0zhG+8A+tPhPHRUSjkxM238UADsrXxE/M/3VZJ+y7lVwElnlv/b+zU3+CJ
Q0J+Cm9FUdknlgadQbJehDoRSfM8ERTcpMIQFXq2nfvIfbXHswpZlQUjfYASiAW+xj7gNJKIoaih
QJ+ThjHjVMFXGLzKD9l0yrL0Q27vvkHS+JLQVt3U1ocyju3feg18+4owc7FaC6z6TC/TLxP+88bd
+u7NlHgR/BaWADI5iufn3r9yQYlsD3rGj6CoEFZzg7ef+6jwW89Zcs3DgcBQRrovNOzZAv7MVaaE
eOtXX2xQDdF9nlHU4l+e3rr4OjvVSpxYvFVO1qSHSmLPS1sQz80iq1XApRXg6pjbdKnbsMDmQckY
X9jPdQ1/8F7Xp1kcNgtZwLRmhkeHRXPm1GToOIcTYxih3j4yciNlcbDV7BrAqsAigQMru7Q8blYh
rSbMe8+1e5mxv6JYh7OatukG5S0V4JKAHVz85efjK5j2ukO4vI5xvXDfjE1Tgm/XzbqpVS1YUU3t
d3otNr+5ILmZ5xlgJt8hvNqHmOS7hemFCIp6KTOJ7AAFFtE/pzDnSvIbT3WrIzipc8Clb0seEJbA
Bg22KbfsC6c2ACEHYk01i59Tc1Yyx0Cb7mVqed55y0V/cF83WcbXTDv/gQQDDQrh/Y6DV3iTPmZL
zloL3XNP+noQOrp7z9nDXqdfaxMu/zMybM0Tiu+rivlV3p3exQk8VhjCOv/b/lz7NDWF/yVyebI4
ht8y78yHGe6ouTorL1mMS7WrF7WemVBzWP3rdW3+R7TX+gZgS0isgAEy/X06dY60Ld24slxi1DlR
BfJANk4Oo5Akf45nYngAOrrq2kWHoA1MurlLJGG+zVkdWOPeK4hGWNeelBbN0qKQxk8donHHPSD/
cpvbssdj+eKFkGrTlGDWhv7GXZHDwGHCIqPaufx4DOLgrqJnMNk7YfxmO4ZJZsie4hj+BIe4AyZc
fC4l5CIgqI32iZjabvf6MXnjdF4eq5EJF0LhN8t1KicVIYovzZxleVF1/h7AotohVfCJT5cL155h
4SKcOKTPSIyYmwc7xpy3Svhk3BybtiC0L6eV+XiG5bwL3a/hCHMdriULEIbU6jVtTD+AREBnzaKm
xotRU694ucHe3XJbAgijbNDGvNb+dDyAKOlJwzRyTKCxv/x+Fz8EyVQwoW3E47fgcqpHbQL3cxS1
iYwX1uXLOMSYPkq+FvKLzIHx7/nX5caTdY2s1nQHyaObtfZyyzNwuhaIrHD7oB9CZVweW/JmCiBB
Vn9OUCzYGAjrTG+tGwHPEbwLyfkdzBSiZ+CgAppgRfOk4NxHabVh/fiQqrudyBqFiiR6OnCZxavl
++GJEt2vP4dbfnXcLRO/Qxfe4KEbXoP7TBxoF1oZ4EnoXkuJtTUgHLBENJNnCRrG/vuZvtBMyqRd
0iMZfitHBzHCW8igkZpcx0HHdXvBY+Y/ufZd3flbj+HE6cPuY9gLG/ap3bqE1HELq7/JCZcSaIW+
tMqtCYEwHgO52JcqaRqo5vljOjrqlJ+FZOmfYr0JHXrQ6Cc3TEEwQOjcxYcmb07cOnr+whl8Q68e
n6CrQF4Tf4XDCda/vR7c0d3RVb1jOQQ/kw42FhrzsvmjHQ5u5nn04JQkc80Kt/54ZSRLu8MGjhSl
A0ZJEuV22/6IrKU2Utw2JJOIglCGN97P45NkQa0ePv2Nkv/xH7XgMuhIePq4yBBqh2INNUsCK9Vj
OzLWkweivCUmHAUzDFzvzN1cOqufABHlzj8XPF37tEcUER6bC0YtiqUB8ij7Sm3NkIvX6dQET0KJ
Tqae8rZ2JaPyzVdh+0kmG9Q79EWVHyTYaCF//VDLM3RIUNW/quPqxG6Za66bW3nZ+R2bh6+nYZ2z
+uZVPDhKvLt5MrVtXCOcInmKf3FwCILWPjX8RuQQZvJC4RcsXPRgnZuXLUNmdXotwmaTp1vImBc2
sZWifWW6RXzkZl13yYaGnVR0+E2mbI4wT+LsGoypnsdVAgkJTe6sgKchn8CN9ls0Npw4jaAfCEcl
J3HylDywNBGmaFG9aAm5slel9hGJiMZPUfZVi5/u5oPpGOPzbfGG4nzyEZTBuKU0wCHmpsGhegyU
3LFef0JTqYwcQRj0EjKFILUCyr90NVITQDy5J+cNdGjTwQ1upbHBbZ2PUncy+4ELYIwZ6/I3nr89
dKriXAlqq0z9XlFPbGOH9FU69d4/uq1W/n8bUewOCXEjzmkeT5cqlRk4Ms7eXR/ALbc5BQ4VoILg
xcLoF792c9RNcWoKFCWBm4mqe3AW9xzEH56AUmxLwae5dusGxNqace/6BRfNTTOqMHeO2VhIwrtK
25IMICtlJaVbj+FtV6oqMesE5WbUoWFcw50LCjBSmxfQGg6//eicOgPsSVy87BViaJ34J5xl7h1K
KIxwwgGg+/hAEMNDpH5oiih/MDWQoki9GBiAo/qgpklXLe7dfWeRGPyEziEQKWfrDkXu/+p4KBOx
Xg37QLPOvUm+rDI/9n0hUWnVlKtgxIFGDH9I8qDOQHuuLS8aMOo/U5BOtnS39F7raePdgMAazV+l
HD+ulYcsCpyikMGwv3sC5+nV3oWgAkBr7J2pT4pHBtQtGb+RSjnbLOIV7hhJ8+3lS3Jg2AUttbhv
aXN3JApppIli22+8dIY77Z0uYHfMGCwz4pC0CaDOEj7ot9Mb8TTH4HO4Dax2rF9hHjxdkMXxyInG
93m83RYaF4sB/6HKfhTw//mZ/8dWZQVh7M4n9DH/geQaoUJL/Z9c/HZ1+wxw8rqzAYtaTGV1aIAe
7BNbFqJdqOPXwpMW5dtiHI7QAdJ+ilJZv/4xD/BPNismzNMWxDAQcts15E/IlEmWUXubZ98Jf83I
4KEazQpLFCNq+F9tsMHtny4nPH1BM9z9MkomI3DqPMERWSPm6yVToBznC8rAX4p0i+a7SuB0b/cS
F2kFgAOIqXlyST/RKrfu4N0OIdCSQUEBfydDUE7OC0cQkxvbEAjVD4Gb+CekddtPd6JICh1zL341
s5/HHe+dGkeN++nuXVamzFC5lz4I6heyBG5QHiPwXcgfdSHy3jKq36rPVN5am9BmYveecVgCI1uZ
OiO76QN0uV5TDiAF/+BOzkSLXVv62gxlOU7LEuoTYRh3p5+WY+yS+/4wDqQc+Sga4+MRlW2ElpGN
4shmv8s8Q20UtbkL0JCDreCMBhyNOhbb7DQZdRPE/jpbaYfCTEgvfB5CqpnwfglJWUF++K4zd9a1
/+q6dJgUfz8wqIQn++7lm3TfP7SiVd54LSsl5oA4r2OMJ/OPCafzGaf+20J5lDctjIYk2pPuK7MD
mZ0L/jyl5zUIAhmK0iUe+mN5JWaa0H5lufTi248zekoWD5hcCeNNZruVi/2DGpJS2vN4awEPTs9G
vqvGVbwQdyrelqbymTlDQQLAjuZ/1nMybrjgnvA1vt5wAi2PvOFM+vLfEcQlx0K7XyLVL6hY0anr
LWQlboY5nO5ZQU2kTmlaI7FQj+R2wFc2j8FNfi729bTm8ixREObFOJc+ljgyfB83p5ErI7JcPWjZ
0HTXFgilKMpsvNW8pNbgOtA4jh/0vXMSg2cyOQBUVFbQN+Zpl6vG4df11Rjlu4onPOKkM0oUGqbg
k1xUun/7LVdCjOx6qf6rtuqF6zyUlcxUYl9ZX1ijzF2rpncyLF5q12cYKfo/RfUU1NuS9EY8x3Cq
wi0LjTgTLlH63fERR63yL2O+q9IT1ZARH/Hc1Q+oUyyJV1q/ehj6tzrwOaz0oalUmC5aiz2DRWD2
g79HcjS64kLnzvhpOVgZr01J1ZxHmZeTnScaqwVWe0tDHnlNobjyAPiaK1kOh7z4EENqsqgIoRkZ
W9HU/fImFnN5e6EF/EtuWTHevSJZBSS2nCde7kkEQ4+WKXyNW0Fh4MYOus4q0b4N1AkvZtzv07Rd
cCqTsc0bh2PpaS7qFstOrJxBcXPxhIUEnSMBvyN67ORCk4oMPVwePvK8tuhNxiHHQ1kCTm0ZObIJ
za2GGdq1Kl8vvPAVC6TEAbvX6V7JNGbka5ML+Y0aqsmBabvNAdFevnC/viqobm6Nk/jzwIx7fjgs
L6zNZeVzbmp2f9Hvq+Ks/d5lV6+K9GOcCxb/5I2rYfCnyh1LeR2HpEDkpRwHDqBDrxZ3rPGrmIXB
JBAYV+VUZ9hPPaZQyBVL+Rg6x5UD8rsOM3JRprsVV4B9NIrXY7uIE/7WovlPGEZTWb9xnZsnVa/N
uYhYgqjOj8/Kv44Q/G/EX1jpDcC8ptdK+XO9KvvpK7+xJEUklBb+AaEbDNVBPdmukn9J8hT2b2XY
LNlr9y1CdYfVX5SlzJKSQOITMhIY/4AY0TP+P04UmmOiPyC6uG6YNrArhP1BizaLOVvhwdjQ7k3x
/J3jkkXtIYqJyszauG7f/A2npyqMmkxf5SLEzX2+Ejxfx8lqca0fmQf/sCkZLwOFrVLsWhFXdM5u
TqgSksdRk3xRGtBiBjXqbLvdoL58447jPBE+dA7fWMw+uTf8ojdvJrRvFsiD5T2uZxl5Rjb3rqBc
cxtfBAbxMc6dh0IoqVgzNhmHAd/ACAGzuwluJZ2wG1syDLF6Xjh7Ba7d38U3JaVmpdmtyIdbYfR9
Jz3ezRqDUZcwX8g4/u/ipRpDKr+qdAR1HzYYhBHpVKT/Yc9A25vYj3p8GdDngmmDLPwLq3uq78SX
5Ap9VYEDGcbJRMmnC3Uk4l9WzyRvU9VIlixkTtWSsnAd9HEY3miLP9hBSQh7/pEUJwglgs2TbeNY
YuEV2YeU2zl5bHEPuedH+wHpviYYKmVMvfss+hVXhTKsgAa9j2ezeCMWhAejwzMcQZnKJS0I0ytO
TwQvMfjA8Ye18oXbwigLoO0aT7sC4NDNRVcTVGfgzJDeMT01u9eybMk5klLXaSwZbXVNzGfVu+jm
agIgPMysBIq4t8fuFRpjF6g2omtVt+TdtDjknre5e8bqcrkfQF0iLAKAiENZUyPQXO3WQbKqAJw2
9mEZ4vQXhBA6BamKcZNpbPEUcmFf/8KEZuiS3mID+K0CftCfIuYJ3DACqH9s1FFTbdF4f5knjBUP
l4I8YF8GXkhKJa+PSx0eqFRBdLAaCTqklV6Mqa2h90OSPefzcVxqmKGk9oseNkShpfaoASdjRdTD
jU7+WYmRGhi2rBepSJ/iolWw9hBPjnGr/Xe1XokCdN2trZ/LHxs5V4nMn8zflPTnX8XPb+VxZ3iD
RDqdWVUryOWmCN2d13RhUbawAbsB7v6s36U4HWicPdtbM2Fh+0D03aaDJuTCZDjn1HhJP0RHKP5n
yRn0nygTanaZvxGVzc6HBVAO92ahpT455ltVsjPtU7RDwCqmTp96UagKBQ9O6iJJ8IeLyc/dB6xA
7YHZEFqD7CAup1ET3desmVEleT6H2t87sO+tycOqgD6tWveYGSjnCWlt00nE2DjKqOjWmtDV2CD2
uIcMROqOXas+e88GAAi9ypviyFwKPWGLUT+YCaS2ApmTBWU7dH55rqBoJvIx1K0gqYmsdt6UCyDw
qiAV+Amc1z6UxUau9Sq7mLvg2lOjdUPCMBl3+s4m7Ey5FdbLMsjYoyD4HfbLzNMG+WyjgM2Rnkdf
sjo723GW3DyK56YCXF2keH3H6kdAYo0Lg6xWX+V6Wu+BWozd2VDarRgVG5jiFHyZP4Qs3Oflsean
ylzEWHSQ7Dp5HJkw0pJ4Pmg/njQw2+YD18CAdyGPtkmKyAxDVebpd9OuKz5IDx/Lb4PFcxS5+oFP
mG04bd0MZCRU0NDenO3uPL1wZ4ieaLkPzNKL10p660VOrIHNIcUVqDY4m+bez+EzuRhSA+g5BL2K
FjucChqyQNmvPRorM216NvzMFcQ4ehWpNxgTJnfWsuH2iPp4QpXyQY4xXDQwuEN2/FEA4n0Li5ph
3B61U/EQxrbuwLoRW85wUiloFDn7LIHm60UNBzh2LkL+t3oD7KZthIz0JcrfIL2s7k7uHLm0D/13
VjmHumBJlu7FQPHDLq6FLLCbK6TRbvdGyo/d8ofgw0PoKmmassBWjg+nFBNCCZaWc2no8Ji9dEA4
XgxlMXPcmiT0x7m9MSH6Sq/1tRSU2w8Ucl+wRN87n3zuvTpBV7+OufxbEYspCwxfjjvX3N30L+Gr
Pc/fpoPySGegFo/ww2fjnvzeaJM9OfV6iFBUVBmQ3BJrZ+QeGJkFUbuBEKdMsmTM6xwn9A0zt7Rw
4ERWYVnOIGHM5XT3C5m9fsxhar4qzrPKgcD3LwTI6WldsBc5oOx0ASGseHPln7AgM27DrKbbCG+w
i2I2kFtSgQxswGo0Fl8bTp/zVADpX3EIi22/bTDgNzjTTbF7ombaEU+TtzC3uMKhwwV9VmXWWCg0
lEbNVPRAJY5q9pH+HqqKd5IvInOYgkl3dt4DQWADrTe1wVZoX8LhXpo6YdQoDBfEzN+p6mrj6T/B
jY1K7iy92mAHjsLfo2H5QWPoRJbJyu31MhCS0WDzwSJnd0UPPNVkbkMib01cBUgktBewvyEzzrlI
191h5Aao+hhKtkKZ3l0rQ37LknTDjgytyFe/b+KkgQ00UncK9Nd9CHy2CvvT2AbelVil0bSvijA1
hymlMLqmKjMlDup77Uu/HKw8XEDN0wrJJjpPAXdfdKNOUYV7uSkwmBs2/NODVhnPCWmmPnfLfTG7
lFxEYUb0xWUz4PYKoehBZ3KoRMDGapcpqO+dNwXP4mli7pyzfjZm5St21VoXCIqSrUMXd5J4owor
iaEHLxjaze+EWwsj/Nz2wQA+bGhOh0IN4ZbHvZv0rxXvxMzyizHP46xBSHf6cx0hu3g6VMjmsP6a
nMnMK4unM5RdGnPKTUHPBhYdBRqni8h8QLdKxGqIceOZZacO9HHPecBHWXbF+fOliWT47J1OERVq
30gJEFZJIgHRgCBD/tGr/wi5VDa5mK+S5om2udZP4MTpQ+baoghc4Eok9wCXjpISOfQlcz+c7S3T
OKIVxMHlHNMAWBeqGV8xrlmqTWlIJad4dPyBuOAl8tVDdoZXsMJPycGYSsz+Tv7bQSfDUOewMWZl
+EplgImkaVOKXaUZcoZIyx0rz1T+ep2JeRm762dm+Pb+lgWCTR/rPWpr1pfkwdCN4fUiDNyyQWLs
JY/WMiDkZIfnoIbxUT8o6RJlsgZNmWxzGjgKS+DZPKWpF6VW5Zy7HC/CnLKjwWjrO/UwCbNcEDBG
rwQUk5LuOh1phk8qOjsIkaZTylXnleUc71U3dzlXae1ENIZlBelHUzTTZFeq7P40E5V9oTR0fKAK
Tmq7SsEg9VCkft4Xu9qPPtukV2topoF62uuSc8ogH0q86fgLHHuJ5uIpuxwdp7uMwZOF4/VkB82J
BvA1g80yl31R4A52CoRfIcA+FLQdq8H/wCRaQvv8gbYPmxwH3E8a8bK/K/UtZ1kBNA2MbqnDI7EI
wfVONg52UDwzV3T/euF882igCalX8+JWtrqXegvlEVg/dQo7b3fk/n+7fV08XmUaDUwE1DQfNgf3
fVUOv2AErG021lcStC1PEk2saLyBsz4lW1lwSpGKmxOsP3nx8ay79hKnMB4nomlEsUSZkIjw3HFt
+OwtVADBZNRjUjDRb9WW51Xla+BIS8B0vCwtusyT9u2ZGIVl2M/njcqKnW6Mm1v2B3E7zjggdjFv
L/bSPIEffE/sXnx9IyUsXZUOeX/khiwi/xt6zYIv4zk8hnWQ09HXfwEQ6rC7CjFG+zeGC0DZFGv5
LtT6NHY5Sb6vm7kXqlXjCQVrwuWgti+bo7VEJfYqTTh6DFMNEdGHkre/ULrkWN++vr8rKRp9lPQo
Ki/nsSna5KKuvYWcxDF7UqOq0lTGq2ug20LYvDu1ZwLlx1Jf7yuFl1XmrwcbiCpWvSmj8nzspd19
26b+tAzTwL+7BHPGwZJsdMUm0v5iUniLokbY4U6z9GAOnP9YVvoCMguec1d9Yem4kLTfrr2ws8k/
BAH7YXGToi0tN2Zz38/DahnXEETFisNppuK6kNurEYj3u5eRtikBNBRjXJSd1DA0gGuiD0V/sJPj
NIr6HA6ZMzwOE/kC2eZx2B0FJGy7Qtkkdg/AuxgS4AQvmEPCEPNwjpNmxvQGV9pSFrItT67fjXHk
qwM1jVflnzktolQ8+HNNXG8HZAwY/V3pa4bqDKxmpv/17r4BT8DX1/g4JZqMYBy3PEidOreS5U8S
0h/MbhAGKAgW4Kh9jtFwbkGbbMT5qdcXJxtI82JfZM8Hdx6ecm6YJN4J4hOaXwS77sYrWFAH2W0/
dZfxhj6427PbX4cdlyunK7Ir5CTvXLF8okdUnrfpdbxfE6JHMzIMkXIYPAK5feka0gvMad0c9HcF
2kAekk5+U9kGIwpKAJcIKwxOWtNADLfLXvbOtjDG727LE0ycoKUiwXo4ndCfAfjZrm03xmRBWfYS
zOkWzeH5zEUvBmCqVvqfGISxudmAEK1W+NqalvXTzZpDwNQbIv1NXPSgagbLpCS9PERTvPcAq95G
sZkPL2GUHr3s3me82JPXOvz7Edkq7pPVe/4OnLOMjoYmreZ8IR0ckQ7pYH+3F1LlMbOs0lq+lO71
2gkRkJIR9YWyYVgt4fb3T377qnBYja8K1Mq8tspk+Et9S8nxZ4Bz+c0/88wlW+f+vGmtnQsWmFAI
0wh0UmZx8jxPvXXR60yCsl3UWGTEHRZZ67fzsxBfrK7Lz6MTFZScJ8X/PQ7Dt2mFHCjVFcnS8og4
cd5gJ/AwjrbLRfYEj6VcrpibCPOWb4BqZrakDdALkypHm/s3mHHtI8Rs8e/fStbKsF+lQdglwemi
A5wtvYh7wiN8XH+8rX7WqPfZVkMyqIe/M9mtAtqOaeXAGN82FQeI9phWaZVzCDFv6t78+89YkZeU
fuX16BkBcfi/Iuvx+lCmSeGmcoawuZsIBVL3zXCqH8oLWkm1U0ZKA38JoXOYsuvPp9d1KdGx0dPw
QaOAFjGZjSkLUhoApjMh/rQYtqLyZwwwOFBBNkLIRun2+fn+JzZw/mzxhqMrcl5qlKXOnVRlE9zW
eRtNEE//KLLqcFNr8CmTzdJWjCmaQoMzhYIo/zgK6l+TfTK6hQErfjd9GR/q75Q/arStdDafTDC7
suFeBxu2LAnTDtMPt2S6lleKCW/o8vJOb44lNN+h+0av39oJviRHNM2Bj4vgaZzW1F2aCtAs0tqh
xFWQBir2T3SJ/6YQk0W9SAH8XO7gNUg1U1q8Xm7OeTG++vAM+3XWtarV+sDUZ7ykxrGyCoN5McnR
i+bIQFieHKSa2y/GqHBqob7kCyrd2T2ZphlSbTpAVi9U3goK/ukHbXYgDmQ+HpgmIbaCDdrQp5h9
ZPkQHEHsseu3Z3GO2ohvqfbkkAZQb1RpJBmw/kYej5iu/IAsV/C1zKikNCcJPkmn+IuSoMMxvGQ5
U55DnH+nP+mKm2PBObuJxF8hieZN0fpVkUeV7vjIkWqGHfv1YsqVOtQ96HCBsYcLfgYnd5482pNF
A/kx9XPumbLRQjFDLAk/ey1ENTZ39cOmfb2pjWiRBiaD7FQbDnLVr4jT9reUnj9cPspadAPDoij2
lswLoTXM2gI18VFCPnJxpnbWDK567OUe87rv15aPEHiVSxeA0SVRkCO6KdKmpEx0rZ3JeNdkXg0q
G9EULt9WYrLBE1Lxn+krrjxeGKDPVZ0H+iDup6ugzQ3T9rmUuFj1Tr2AXYTBGvf9qZj/aP83re2E
xk36ZBpD2yumqeOW+yVGy433CXdJJiJt0sYKqI5IND9CPUzpju36bOCelkelfPjmTjlPSGXQNUVE
zcpWNBHWE/qq0c2m9F4f6bw0GfHWQqiQD1KU+VR9/12gHUjx3Bg9VaT9UwjL4dH3yAKt4/eHvK6S
HUDfczotC+0N3Mrl4oF2YfF4YosxYKAlU2pOw9ti5sJZ01luBs/4cIzekY33EbLa1GejTq8sYcBU
QaPWatxYnuBFhYbPddPPVBJPs+ch36BCpa0+ZK2sEpukRQ5lh0+Bkn0nhBUb8ICSWT/K5yiuIVbK
iZy4T5uUqoK6/OH+vYQtjsf6S8CmLGSH2+cMUdeGi86ZdTvMLPwn+WaGW4XVozUl/bBv2lfMFPIG
FjnruN8WkZ2N9gIR8c8Iza1pkL7G6tPF7KbYtJYrAFjcP5lQPf9M9W/qn1jSoD7QoWAkWroDw4OL
VRPpJw7B3cLZ7zBMcX68l+uWW8GHd7eiEYD0OIkuN+rS1UO9JiHIegYLupx0UlBtY6Y9BLaUBZsh
If+6pnqkNlnx1fWJ+NTPUP7vlSBQxK3qlokk7DhgEEJPKH76r0hX3cIpzf8DvuFkQeZ9xbT4U10Q
n/su0Tz3XX/yxDTDaNoeMPHPYoWhMN4S8eYXBgMhXkK2WgMyeMxr300BYz2zXTk2c8bhslWuI0d2
nORDlIOfzoNvsIDBZr1awv639jeStItlBRkzoXQ/ryiOWSk05oRHgMd8Xy3kymaGhJK0v6WHgUbT
cd+oz0oUeWNdvHAvtpVaxFn75x7NeD0LOFpCr8dv0DfXJ9cY78/fiqdhAf686t2/+9VK0rJuoriz
Ous30rpU3nCnRerfUVyAF7pGVaG5qGYVPr7qgDmTlb8IANsiP4zg8PEKV4r1B+JQql7yhUfWvfEq
7/cYkWB6QaXxwgo34sMPGh3BoG2zRFf8NyaFMlLVFmVRmVG+XYmBmQZBwW6chRf2ry7hS32YspJB
fv1yXwaA+HOSVDQFrv904dXFATZSlk2cIuRKAkvD4UeE6AG9jbKc4Hm7PXQDCbmKNjy93c9qrrAR
PL7ampz+VCn3NV4UG8Y0ZTj1kGC/RzQ1pA6JuZhTbHFe1ZO6S4U+mmAhvjN57aeL8mVrKtrvl6iD
Ytf7ymTHjpo0rfBJantBEb+JRsqpfbuW8ng2p8VmRUyM4MofLD1cxf4pbo5LyjwCwvLyDpl9bP5Z
5rwwX7Ie6Pp3ZG8mmSwNBOkZC9Yhgrewt9AMJ7KK8avfBi+BCm84IsCN+wIZUNcljIVJzoEE+Gwx
3Vq4j/3pSER6zyi5MoDfauq4BwQYQdO79N1Kd19YPnMNw3vjUbLml7PFjbqJ9uHhqJanrtghbMlM
tQ9rUk/Vw7v2OlZ74O2pKWvLaABwmPgw7X37kOa7vunOc90gw05mZ/fcBq8N1wnPAWIvpULtAiFH
NERnDSNWa3bbLc7AQbzuGnk0L9KFBTO/CqcUA14gYZ5jIckgSH6X0SHZ7wIMSBxuZ+RwU47Ylozy
ECwrNIyiqJ4g5AEErj2OHLVjOw4fIzfnA46+AvXFYbpypc9S1aUv3rLkYtxJ/IVTWKnFQb+Xdc4g
5xfp6QWZdBldKJ+9qRhNnvpLYmytJMTgdriUK9Nf7/0x/kpUZHhYCiObLXQ2d9onuCrBmZGmoQOX
hUVGB8G7LLaProTzBrg9k3FrivW5a3S9BH+MMouXKx+oBDG/uRHX2deKs/3y4HhSwmhYM2X1Mn7/
g2YJwe9OHnI/bDyT/iwVm48C5qyXcOUxTZItmy7hYrb4vyITT+k3ZjLm/d+5HW31K+5nVrXim31X
Zo8vmjPd5ZaBskRuau24Gi8NH+LI2EArb++E9AxLcKT7kdx87QPhtm4h/NZoDOtLcxnb9yPC8we1
82LTcpntLBdIDKc7LHz0zzJpITmoIVg6x+LcnehCqEEqsCbcz+P9uAj3PnlmzLxAl/96VMWQPaQs
wTDy6Chw4EiQkHRBSZyO0wYn/7PUox3TvWYnuAaZ+wiLLgmdXQziWcN8LG5xbyLCsiwJ4fBvdW1E
dq3DXjK6w5JO5kjj8wElDTsqN3GwHjHse0Bcxoxnr5kSJRWDSg7YJNLyR+/TKWNhYfjZw1XBi8kX
4D0II4MKCUEWSwtmLsIJ8oOoqxEnwgdOPTfqBnAZivoK06lzsMqvtmJ/d3tcO++9pfUqYh2witFM
+ampYqWCvgwFNHr4Oq0QaD7DWXR+zH0fbzlRzxXeKC8o6CQqGqEod/CwzpT5dZREsjKONxYhNI6G
/B7oO8c8i02bW/N0pdJw28Fy3G31LSdcyIw5n0kI8c20nR9KrVn/kOZ9w//7f0YHqerFPy667r7j
7Zsw+la8B84w/ZfKDrp1blfrIMpmqQkq2Sib29jtCGJNkmHiB6l7l/vVj9/L7hEAp0PWQfCo0XQs
XFSTFoxoFld43w6UcFlit3f82oGv3iLhj9hp13QcahQiXzNBgCtnJq7zGoL+vWNQAvmtjhVHN2IC
mBOjKXiapzlP7wGr/o+ab1++rig798D6xtpbThB9Vmnh3gFgRRg4Q33227UbHVSkr/WxJy4Dj/uV
U01qY3yMLszyYL+amYldnRgxTjh45KEDoI/He+b5PCNxiQe4TwLavVpuNbHoT58scqo/Ftx4eovD
i6KA1TP7bruNUrYWC3VO9D5QyzV6uvQsv/yXMHY0ttYQXOEzAcAapyX4LoMOJt2eikOOB536PlPi
XT46EGv0jxHIii+6hYZQ/SKPU/3SJg1NmbXRqXlgiOdmgwYoMcOi1LK/EqYzpT7W0+WLKYh2bzgN
TqD2EbKv0XGuof9aYGNUze3ubqwzBqQr/xzHfA2FG4nFQU68HpSoHEJ9Npceiumv2dUjP6VMjmZw
eFtXcbwRjCaB0Pk5AB/tO5ta37/n0WdQqfCSfmwOyCzdehsxzIgWdwybmZfD5+MqrYRYenAV9fwf
vzSwIiaLXPvVvENrWHrTHjE12UsM8GLOf/uGACRnZFjyRVMSlnk+Wha9soS1Ht5Jg+0GtmIW+x23
h2NQQfW/mG/zkWlJDz70JadwF8EcEoipH3wosZTG9WWI0zvlMIBkhyhn9cTlKp32lWj3YMMInJz/
M2GYdwtKKjFRFC8VtBdvT+s05FflfswmgzOOuHdaQFpld5LWiblIy31iMHOLA83S7s0mEMd88mzr
aOmUTGed25rYkMDq9d4uzoWKN+Er9iy69IdgUsVWyDras19CtexK5Rvwk0RwkLIdibaARPallb+H
xyh/UBbG1AtkWyKqqwXhFTfH4/dv152kzqMHtm5hRe76yb7U/634tVxelqrLBTPZWUhE4teH6SXy
yjJ35jYRyTDD9v+9It47gAfQZGLn38gOXtxeB8MekYGzgcES6GSMi3j2ED1t/WlXUIjoPqI5cLVh
nhVVKX5zu81FjtUjerCFS7GNnANbPkerIpgllFq6I9mEFnhKLbSmwXtjPhXYuXwpPuTMIfMkKUm8
AXyVLIziVPayYJKWjuFYGEiaha/sbu8uIuByQLxr8vVpId++6uDyXvqKdUh4nNGFmTlxnWbHnb94
2bFnM+BHxuTJA51o7HH5hlXhvSBwpzo19MdAd4ebncqbQNkoIzKpk1zp3tab40zDT4crZ2ZrrsAe
K/+fNVcLJPXYJak0IKAJvYLic4pyTR775Sg1MmRTo2awFeESEmWaKevtkRU8h6SvVznorerzI2Qo
XRchbs1L/mFCK2sejuUGY2AJC0BRBiTvWSbOSdU7XZj6tKr6p2XY7mJXwfnoB/wKJFwqDEEaK9QO
4luFMHav8JOMcRJHh8nU80E6w0EJVfjKyEvuM+sUzIjHJsDEfJsmHHSgrOj2+ZcBYf+a4GAnXYGo
sLj6pEpAjg9m5VlX+IfYsZaa0melkwJRoyMsS4c0EwtmQwPYpvzkdqbOvddD+IcKIrfR6awz7e9m
NUceHi803G0INmgvpu6jS/ahIDm8vottX7JSLCtVvvk5Oukb3ZvAnsNAxgDDO8IPX60q/awfAO1I
rsSSPxCU+VILzTuAa8WpEV5LNFaID29KR5akrHvLmxlTFJWRbAm9vVNRB3mDeLBK9LLjTCNW3m69
Mu4oEHftbNXNRpjryi6wE+6xcTjDUeqSWNrrn0zFGn1IlMf0RvF1iJX/QeiyDAWPvoEx0i+bGbdQ
kcWip4Vn4jqBMOiFpi8tWPpLmpgtkojwyn0IxY92zTcs3LOL5dmmNFD92BMhzfzAXJW79MeAqOqH
EgGQaRfLjL/hzw8wx/vraf6xwo5gPcUrolXeTxam/X537WQgWigzqzi2ptXYU9BOY9ge8OXvKKA8
Sk6tKqnFz/F8E5K+jjJBgZjdPG+ES/ytwtf/g91DB8Yq21/qv6BpLoVxE8vxYknCV+DB9ouBl1ap
HUCsCE1ltxsYTpurBY1VIBMS8Q/9su/FG75D3E3J19KNjIwL88TyWRCK0U1OiT2yqcRYQ6XN5I+V
cvkVF5JmPmDUSONbpsm+2unb1lzHGGfLnaqcokTxOzlpKcUQ+KUXOfxvOJOd3fREm61tmANUCoXD
EqhymFo/d9bNUkOVudrMkk8fjiViMsEPORHPtxh3+bolwJPdt/j692VAcpv/BX/WtediQaffL2kr
kcKjdXtRKrzdZ7zJHTJV3Ex3n7+4Ad0sFBW7Bfv5gGofGEEYv78eBYcTlhat6g8YeFeV+cQUvzhW
8lGKr7qeQ3MT0iusLv61Qut7e6jLANhD0W7aHEoZTCl8zsqH94+kQvjKJdH5N1B+Myz4ryp/U1p2
HiXHHbAHK4ezr+n6TSbXAitSXxNL9jiaP5REr7RxEVKQ3bFb1v5xJ7Niyq0wgpPjojCI6LZ6Fyjj
KvX2zqwyhbfHQ77IHXwUVgFTAd0dWcZeYYyi9AICcmPzXaE5gNqtvkc5XfFOI6bEsnaM1CpIySC5
0ehhAjFYNNLO1gLx4ZusjkjLRYcFlvg+apdABElJ+3IkdsF9QY5zhbLOzGD1BAuxWOeirSEw1qy7
G2WgwoGPgkn0uJQje/+Q/E86NP+oqb11HIwJUj8tTlT2iCRfLtQEC8eLUw3++WexiXcJmALD5tVu
ntOqh3FI5tKdyVIbeHorjowlt+Ir48xzWodcvsMPOMg4kregSen1PmjDGaeTDiwC892bKeJQt3rp
5w4bDcHQ+lOoYyzovo//XPG4Vl3aDvovXqzPQugsan5A+TdCLnVxyN9XMnh8D8ovSMxLYg8dfl0U
uBWz8MFSNuNlKE95poqPsD2soTRXLU4ZFMP01jYMQG0pfIQrHH+0b5IIwptCMinOb4frfI7vyJBK
dOn8fT3V75DQQJGJzxRSEFkUFrWhkYQp8Jlg5FuGLGWHoq+Es9XB+UHKizmnAjF5AvevKWFxUnjH
R0ZSVxenufhljN941z6p7N3aFzACVGv3i+Z/pqhiSgjJRzvEySYxVnCxwSNx/l9qLHHnYXjAC8q0
PwV0P9EZYHM3K48LDNR3k7rmK+fBS5o3FNy4TFIpyZBKbnTDeZD5VKNCJ2WCXhMOK+5Zz5WtflYk
YR0CdOU9YRruNk6MRYaaQrKJ6q5y2VgkInZX4mmyOJRfvved5ah3ENEeVP7vuZ68QKs0wER2MMFi
sHYS4Mx74lUUvryO+HLE6L59XDfG/MuWafr5mTCUgiUxHSU4gFN3r27oiXV0xvuCOBNbZhmQTnIu
msF0hIPXfDAnjJqM5d9BuyGa2hRZBxTQLAvm7L3acK8RDflLUoz1cTRU2hACUObnzRpImwSulQQ7
nm8KoOp5t7YG2g5zNTyWFJotgF3QqA25I2Q27npvvhgsFiuH1gejPRnR251oiMvN6sYwqXjqO7MN
ceznn+qriZRLE1a3mfRRNsPmUpUrdAxZBXvXrst8hfxOHof5bh2QL3bUzu0/mQ6zLGan+F+qOvem
djlyu+EvFDQ/OZwrm77WT4qTeShWoX9qV9vgE63ud9qjkjPeIGaIIyrH1Id1iXb6167IIiIhYR1B
t206PXosVufwFyqsZCDeLmbwb9O0cDjJfPR5JCW/HII3EcxB1gY6v1Ois1Yglnu7YPG3K/lMIXcg
15JMesCMCYkBRJYDUH8bi3L4q2zkZg9Hr4NHPchv3fOH3VZC1HsoyT700XMt6jKwK1Wm38ADUqtQ
WMPTUULLQr/DE8Cu8OtwN379eoQ8nft8CsPt62uR6ZJG/cpoEPexhwK5JYucCXmFI1FR3/soYBlV
CSvv4hp4/dJW/G8FYA7U7WnQyWQnQUVK8SLdokypaTc1mbunf1g/LS0rW3JNSTuCcA4zbQn5T8Vq
d8otbiZ8mO8I+yUQDR+uKjdv8OuJ9kUSgnWJ/PQGz+QgG+7cq8/TqYLqjJzJykNpCBJnPbcXO4R/
+iI0PRzpcP+Z1ZI7/feCBnxfm/bLdfFCUbWI/9q5OxXLDEm4LyOpcd9+E4kuIBEfAjGmdWF5ruDn
ikyXj5WydY0F3joGzHpLx30J4To7hkZbVGZcglR5b4d+uSm5whTue3A9euiEx6HCzHhomwzFVPH/
C9cpMZ8NRo0Nee3v03VASxy0v7ARHH0ffQ572co0tHX818zedUSNd5IO2kW3EL1pZc4VHrqB/LA3
wSPNevcaB35xt4hRcrrJtkH3HySI9tcpwEPH+ciCJR7u2+R8xBnIB9XBShujpYpu+JuIagkfCvbx
PiXq7ZwQIWn8N0GcrE5c5q9Q1AvP3iJvZMX3wfYr93kiHSJ5aMi5iS6vjljyDuiRj5WNm7Xd6gs/
ty40g0KCiFmXFRTEpS1fdpy1wQuerFWtBJy7nwWMxxlNILmdEgk4XcerV9hrZZAJDV6exNmF9uzB
9hEbuh1ximjlkWr6Ls0DfrF20bxEzyPeAtfK/8vApbPO2vgsBy5zR0cFMktQUKrMRo7utlGImtSM
PiyzPHdE6qQYMpYk5PuV+l5l/HY2bW9Mi3xQjyg7DR/iUX6MENk0DvWo8HwbqidIzfVlq3Qfz8vQ
7dDzp5GVK2ZaSloVajx9nEwmvbKo9AAvY8J2bdQf8UV45ECLmNR34VCXtbnF7qkIW8qQtzUVw99W
cwbeSw31Sxuq2UMs7wuXdUKNm2HnKzCpEqMvqLdRgYV5MlMX/pinRm+u2yK4ewaj72bv9U8uChW1
+kjSKQ4i/0b39WGcU8BA3c0aNxlMGKw8Q8sikSqJJk/g0sjdFfl8KHIrPt4PwZjNUyCHortRaeLG
jZc/apkAu4Aa8vagSIeLNNUdgK4ixIj7AdWOUhzgeOKlWRXRx5xBQ7L33nrBgxnhedEJ/36pxnB3
AinjuYss0rWIIK7SzW9itLKF4YWWCVgyEBwiO8I5i9pl90aLy1atQrPNLewJLcx6FJz+KTjQ5r54
BFaS7AWtyxeAPan1cbrWMrW3qDRvOdHVwJSdwG1JgLfrMB0Rs92aXyfoTICrMO6Leh8LEfFAw/Iy
inmu+FQIDIzn07owT1qZ5UipB2Uoi5AidQ71tnvb6iAtNnKTf0/CQ9l+O83r9wTFrhtSUMg6tJ0J
3vT7ZrW2tnSq5ZRs0xmEqwVjUEZM/exvhWSChs53bv0w9ExWqNNjl/RJYRXMR8PZK+Wr9jXXFCCH
4Xv0IhSDK337lUts6U8bZXvufT+c1PSlS+Ec/aKtbgW1ErTPTNJSq76uZcCjAj+PLD0m8RGiY4gb
vjzSinyrjIMF1WVntcX5yeHYNntRFjDsO8Sqmd/hOJ+2FjPbQd5HoYhfbMF3rYn78zCwLWHEik58
8jAJzSN3Jvce69X0ORZc/wB0pISJb4pvPUqQbodaJkWlPGr1hcmpHTGqc1VJMSw1TVyXaxnUD1Gp
26aJKoZtESF9r63xiY9ymnULLMWM0EKXhjLwDpZl6TLf30YX5y1XCn0uHNqBKGtsY+jxNFBmjimR
nwh7Xi5baN72wmCp07aaXNSq77tAK4LQTP989cy4H7EahSPWjWKHfYjYuQ9K5Vf8jfAKFXtLDNWi
BmzqQJA0mTpVSvjbq0UIVrIpMf2VnVpBTCg94OhJOQkhbXbg5Dj6KBzH9lx0+w6Pd0arCCajgJsR
Dzeu9hJd/uddbLo/e1zOq/AAQrCmrn/NYAUkIqBgn2S/WDtkxLwlnnEEh6eOUxd5VrRJ79MCEAiR
RE9Li7qVlEu3aM3m/YabWVvYFLF8LE9CyxhawR+9+QFrU88vHQHoSYjZQu3ld6nSIGJDWRj65N5P
uNldMOcjYxTtEwUg1uayX/5vLqw2Ih3EVMLGTT5EAPalbRROA55Lm3fLfsH9yMDY+xXZeC6N7POQ
ea5ZmqhaJUg7b/YOrP7fnvn6RhfKA3q2fiyo6Vd6TMxO2NB1KXd9AwPnYFiKpB5kpbTy1Cgtm+Yi
36+4/RdbJnbH5jgCbS2mKbDEHx/IAa6b9qGjTaL6bo4cIDF/kb5AHNwtYxiMCX8Jbz4XQdsfejCb
VCzYkTjJthAtgkthdFpQAeSJPln3Zy8HJPFZQyFlj3iq4YpPxQ4CJOj3F4QSoYa0TwCgU85ZeAA0
5pb2VfuIaRps81JMiJTetYC5sjvzzhuMvALu0CJ6tr3/HrFu48D7BbpCVdQyVfyPP58veQs6/cBh
joMMvo6P+HlSiThiQoobnN4EoM/RNLbU6ssRdfBvtYIrYkHPGFNyXUexCai51lweq4osWnb/02K+
sv/Heo/qCQsEHD9eV/QUU+1Q/1x9nC/kzPeqvnHkpfpIy5MZBYnahskaF7CHfs/D9WtutQgeIAMH
z5zZXaEk+loGnPdmBm6nO67s8EPLaQrZwSQFZ0mcE5Bc8Pz+X4bKdu34rj8mY5ZDTv1KPPbjkxAm
R0lkwFYnDOxgbn3zhk4xmP9bBNE9QR2d3uCpSWZPcP/YHr4PHQlFsx+XUR4zNekpSiyf1L9QyWyj
Ou6OtxjDPhXf1JMwJNa35ox36fbDWu1YfaO3bBMzADSzeJ/vtYczAr2VKzihiGADscpJLIiR0Nzn
SvvM6AhCe4LmsP8r/oNaJl6ObbHJHMAhOT6x4ZFYdh1qKaLOb0nmr/gma9Pr4/HGKHdLaMXdBGTd
aKlDxj/V3PUd6GAIj83OIAxaP4u7FkE8ActztHyF1HTMIq7rmVB9WS62fNZIhS//yk/Ue85c9I1b
N3hj9ihuhO5U7L00k/gBur3basfF3Bd6pMzT1QoD93RnEThLOZFu5CmrEgMF+6y4DhlOptpwdzoX
Fpe2zBRwT/sqwbAsCrTJXZT2hj8xNuKSDzsFNOZOSMaTg672wvM+5y/TcuVN92JQ02PgkARrplQ6
XyT8chwErEtBjQMa6IL9C0WWd4DNixH9tocNwAiCyUZQVGM5dKCVIqbpGYLVm+Q9chOgiN9npq1g
9dSilV+uDcOF7hyAkcFAe5VZbzkigr7udvlFy6XiOEDAhOIG3ctNZ4flXYlcq6Kp8r6tJ66jPW8G
jb06FxssCitN4OZtvK5pDmTraM0uhwKNxTeUqKNEyd9DFc4787e3bJvJWf0q2s0Efh4YpX/Z1jN9
DQl/yJcUza9D9Sezp8mcxPyLYTBYJj6g2/yFnTZUAzcj0JNoyKIjunK97zHC+synGeZG2Xf1cGhS
HoOyFb3sC+j6nm8b3khFhLvpQhdG/ck5MnYOCPMEbzdwKtWYzSvOlO4pJ24NSThA/fopfHy7UWuc
1BqhLrXmY71nf2ncgprmK5n7RlxbfLJE356cmL+wVs8Jizi+2tjZ2Ly86qathOpo+F0sl8EM6Ljt
UALZmM5pvsOiWCflrICdnqxzbRY53ZEfTH5CL0j66Yo8PHTGkjxdo2d76JGujMcffS/KgoLjEy+q
reBa/zKz97FPwa28a2k1Qfee0TCd/O7TXT80V8vqgYjXyMTqLzKTRYlC/g47PN1AvO1T86doFHJx
oQWumrPPh6I9xXce0ckY6fr4y8ljTbh5JsRK1NOYpQ7JAmEM0uUmsNa9w5hnJ8SpE14L9xpr8rGU
6HwsdzFHpjXXzz+qFwt9yhnzMYOvtNXuMM142VPST9GpB1ySAiKgljpUEZKTDRCgI6JWfVXf6HJS
Gy0rnEIVWOYBwPcyAF22P/wxKkzSA/IdPMmUufu17n7QBC9HX4P6LkBgxMDpn9sKh4O6K12ViApc
NRDb2h8WipqarZAuIsQBeBUaestl2nO4NVV+ml5dGLvMUgwDUxRA8oy+V4mT4SbNhlUsOErrOGfc
K26ynboKdeD5ahkuBuf1tm/xpBC/BCH+06AUdLENnxTL2f9+iNCcBNoT7/Nqgqw5hnAf37rrMIUl
QslDelLZKWsVIESsC+EQk66CiiJIKi5xgcnGwwcwQSrlVxlSfMXvOW4Hdn4fHJsTVZ9Lr4AzTRg2
t70rFDSCAwsvZLtWevjGG6EF/JhXHOD8KBEsMigtBc2y1HGDVgX+EtHrLq8RU/CQmHNBckGOBLa2
2gQRwrkmbqGrZ9KW8lY0JctNK9jXWnetV20yhdFWzcn8kQu+SURPna13XtlzAfMhXzqccPGmoDeS
oV3T708XhE7kauT8w5R5GNwMwqzrQMkaOBhmRcxzD4vuuZpsouc1c9+JOWYl2JjCA4x5ZkFp/iNK
MxwornqZageiIWwnnUxhQrr7KUL+DE7wIK/yYugiw7Ey46CwJgwhORSn4qyY2bDYaWZ8Q+aZS/lh
71HKPMOgaIDMiCV77hwH5l4mJG70V1KBD0Th0D5osXlzR3/Oc05BgwMSRsLYuozVNgCb9zxo8dyR
G8O/qlrYUsS7KCl7Xy0jq5kv63yq8z72YaHTam4nXiWkWbog2IgfoSa9Birj992sxRcCO8+YW4+N
HQ0jPpK12SddM136UX6IsQKWK6OCxPAaVmoHAdeVW/pjQwCoGvtdNE54xNDwNOsHbBEKDdkOxK6r
s65/UQJlm+c0oqZX1oTVKhznKaAsqG9OQ0h8M++HMXIUcuJhucLlFY+nxQkjd/ANWb51ACDvb4EY
YopH1Hy1XJ+cRJL42sn5V5HPPKFpX7OXRvoTovIkVhN1LR7PHzCnhZNh8KBxEGHpHBKW2/Xzx4j9
hgrWHq+MycMHb9z2/jYCFQoBfrv+oJtnxTnNJppySxyWM5LLaF/zdPO4z5Igp3LtXsU5PWOTwep6
Pb2KwGoZlRY5NYLN03p1b/qvXLuUlABWc7L7tgPRgL5aWYWt+27sJxKnn+cjUR4jyqem0Kilqowq
HuxOa/4F8D9EpmvPI22MRbUUa6WwiMSvlco6DwA43e85KWrv3I8DZSr7dhVohiEA7NKg68mjeWMw
IXGwOP6OrOyh69Jq0k1SQBL8ZyG6FA/PXyl51zjx+3AezJlcGKSUOrNStvZBvaKFPlMchT5XXtpv
yNwOqsgG3KyymOdgbNvckP9zeY/3IvYhKqs9A4qHKDn25XvbRfh9t779AQ/4td02PsZNCM6ZMH+Y
wgvwontC62UBShfw4jxArTmXV/mG4vTHXbKUtru7k8UYfdwNx0s0u0IRfxIP5jxWsMwHpVFmcoIt
nwlKOZoiPsgDnHM331/mcB/9xZcNcizsK7F1U7R+i+SLARc4Y6vHZwFBLg/nClRQXrGQ5gURSIH6
QnrJ5dB1R4htxo2UGvCWbaHBejvSqLrmdMn4m+x9jYx/IveZ2wAJp/IBZZw9S8qBYgX2PXmGiCpA
JKwCDd+pjRBdfaKJhg7B0pmg1nQqFyPv1WCN8/Zghws/jOiDaY1liZaaiLzOadshojJkJnCkBhBn
IE1oCeeAG8Yz1KrcXx+QGYkc+W+0OccOwGIxh4c5tF9F5R570g2CF5yZK0jubyThT2Z2n5xn6lJF
B3805bjMupoZUfYAaMGAxtBYZQ/AaHC7n8C67q2506m5y0qfMDBw98lpyfYqlBCo6deV6oxj/njB
IAZWBdryt/QaAZBE6h5zjvIOUU3qDoyd3RuVJFH9DiYTtZgxzBXTE6dqtyVFjiESFxKo+I1DIP0N
xcmlu0B17NZtKX80BfFYsIbCv95dlSPtwQ+teMLOFEwZZK7X5vnmQ8khLbhx75mZ/uD3h8Z7iMiQ
0OSP1OjtaJX71bhdIijEE2Vqjh6CCoPCKztQg2nK6ZJOTVCEXQQFLPN9C5zN6B8ig33t6atu1Uvh
67Ac84dS2Dt8fpbk2Fkkm9LgsOeZCMov6+TfYEEenjWJkL5bPrXdeF5oT/MErYRrovIu139eFJRn
uyyVr3yJ9Mn0+TJ6+PmD6ZnnOWnfgb7D6tM+MiAfPwmOBgsTbMwBXCJ12N9l/WbAP0B1tla7BaPb
FCjSsKG6z84DyAe3pIfewW95S6Nn7m06evNacAWOAZsYLXMvCT5IMB30NZcKzLc2eNoWrWQVrRGv
rOVX+77qSrnjn197XhQl6BmrtIQPZ3l/sjhTx8+UZGE0MJatMzJgP0wE7Piz9zH8+fN0gW2GX+cx
vqfgcMAZcru9HB4MNn74HDfBbY6Q0R6Vybs0JmqxfWQkr3AG9TIxYgo5TVfTnggL4enfaTb8mrDR
zqD5+FYe8UFT7vyf0yPfVFdRgToa8J+Iyc1OM6u2Lf0T2fj58EcG5IYyM1D4BDZW/vzRX5ElQf70
m+ZUqnjWqoNcivzHEcqL6RtzCuZEEa9V1XsEhi4oK3wI2gVlJ7aIRoKep+eWVTbXrAP4L1e1UrSD
0LCLUhaTNFoJBcmcc3bXbLBpJjDwMCWIhlLd70O1H8AaUqHekyb3RPqP+LErlngolLnf99fbd6Om
pUzrGgJ7nvN9ZjlP23gmYNXYWKqpXcFBRgZ5DxibX6dCxu148diMWKPe0GqfS+rkugDZ9xdnlCk+
OmqCe9ciZG8xASEEtBHJVT786lxTW1udxCsQXdIYmaNtHw9bc2Cfd/IDldKz0+E8RO1XDwf0uQKR
tpAXys6LfVHcf1rn5xqR9nTum/p/S+rwzB8q8bLIunnJXEIYVQDXBqZ8ZxT/JwbAT2oSl3RVpC5f
n+OtxImnnvP53G7RUEsAFbATe10jcgV80pJVxt8TthebLA9JxJI4gsrPHTxurSB+9LF5xiIJdszr
sgHIoYuH2chSUllLpbkz/0xTDWCO3DhACHpJn0gz/MC07/9Q6C2ncPyfGItmDafJerVCScnivDvK
0DCdN81Jyrjce5jE+Z/CGKF499nAnlTo6wX+eVEMEpEt6V40txsFAqIjOixZ4VX2/i8qHwZn2OSK
nzsAUhd7VVVeVXsH85K//yGaC4lOicM/sOPCOeKQHH53OfiXcW0PZ8XH6MQrTn6RvWdYZBClPHvY
7YrjMI17rHHWnruXVeUwsSQbw5QF+nNjVjoUB8a8cnaGBibG66fJmJrxW73r3t0kfw7tp0DaiwSN
vGd1SAYL/rLFl9atRlaQShEq/IUKIS2DrTqrt8tHxhOa/KuL+al0jJy59cWB4JdL3KTP3jvev9yU
fjcxxu4WMfHEqeAoD/kSuu/34xCLg4zmSt3iTiO+bdl90Gb62E3ngt4Fz4X9Z+VEZTGXHl9VwjXR
LzbhDoqar+zx6XKGy7UEM3QOjDBEzDLrBCO6ptqNXkf/u8vRHA6e1nlOs2zeReyPD9DRPX/jRFlk
HsXhAN75NyYHS1is+mKgTEx55uEzc5s8qSUmzHhCzFS2tgMeIBvuzdBVLp81FNcBY/s0m/k4Dwmb
o6wkwa0KH5C7KEgWvntHkBGhLViINm4Q5IPyBE0ERNZJi9ujt1q+f5xOY0yLy53mMT4HXsblsmCy
zfZmK/NuFylbH0Z2/jyPUCplDW6MapzstaMYRGpAyrtFajT/myD3gU3MMFBIonf7hCP+k6A+s/re
DVMbboqgF3SwWSNZyMYNYW+u5w3GBzoapSjDyAhP17lxc7zVPu7ix5o2LkcG8uWCajpQqlPG8w0E
KIOAZ3dk95AvI3YWYBRZ3heZJf6azbKFuRtZxUzDJ3i3MeOSEyk/0051ES4VCiBK/VSPCYwdcTt8
a2gsdLNx1bpKvC2GF65CIzKLJ5OuNiDX782QKLVZMLI95Vv6ipUscdJpIc9K7+hY13lWAu9AS9L8
R8ktqrZzyp2ZxlDt0lb/yLtX1dV7J3kAmEPrG6yVK7ebdGcrE1aG8NyDWud49hlV0k7/4vwRmlpP
Thf/akbqfNlXehDQUX4mNkSd5HQsRneSnXUMHrS3pfW+64aiNr6CJf3bXxlXRJAvfYZhmGEkwKot
jC9Dmyvk6nGyFee8wz0gSqGuKRPpDSr0LN1pQivFKol8AQXEaHEbcLcT8dWBnghVDdhKifTJCveT
iDjzFRS2DWY4e64ebQn1AQalTC6vtGoKtDhvfDAZPS5VBp/qjbyhvi98d6hUlu7EHjs39y8oKzT2
XFZQX6bx49ZTruIvq6JmjXbs6jnehnGQez+TjvnnPU5Soy1401yO6MocJcLz5UI79RyE6F9LsDuS
bYrPy5qYzF0kLjg25+YlCa+4CDROfBh1SZN2pzjqGVZqlVxqdymfmdUY6H3CbJFn5QEdxNHherEu
0aH+KKpob6rqcx3ugBdNTzcX9UrLC05h+igpXvbPeKE2y9kJv5WELfb5cq28ymqC8DImNF7/U3X1
ETAK1ETGTlsM634AfBiHd75ej+Be/DhhQRToH3NP8LaimCaOG9FZsofK9Vth8LT8seGH/3xi3CjM
vWCng/aoTxYuWjYkMm/QlAmhQqHrn9HIHo0RQ9GS3rfuUANkUIPvDQx0Bq1QS6mTx6bYtXsdASb2
zQVPa7euxBZ8SluV+og3fuMVHWQafZ86cR2HrKBi72PCOlnh55DgBNwVMxK3HOrqvVHeotxUttTu
mjEiLbL6X3ZDvSvvHT9xwtRs1oDzKE9nkPOqmg32Ba30v6a+jBtDjviG4nsM22s+jEOjQQHaW4MV
yIRQwW7oHcXbR7bSP4ncJwAfpkMuOEZ4+lEj1a+VtFrrzcTPKNft5er3JnELL2JmU1xSziTs2kzx
VkXU7lmpnYdztAK9Q/AR6hunkIH14JWE5ndnNOEtoGsvDA2z/6jZKmSv5cH9cP+IYML/t8cLvB/8
uGJr7YTtx3j0WtaA/dWMSLk0jowjvaz7r/yF4t4AYjCRySnMTx8e6ayyP1U3tug+xQnF7l6Hxnx6
cPNPgeFNaTMcCMdAFymHWBbwb4rLulx/UZnH2qStFu6FI+EuZPk29CejkG+X6V1P06rgPA71ohBt
/oqTkdxrmWmzV89GospsQd4CDvaiob4/skxO8w60Q6jruxzCzZKCz509/U4p1G8f8lUjmBwMm0AR
prjFKsKtJua4o0+iYaWX/WFgAIHNDb4BcmXmxmGe1RcEMoaTZVkKYzJuWIMlwaNXQT00BYrGpPLE
Vc+tuFU5TbIjrDHXDhk78OvTUgbOhBq8AqaXv7X0PGBJ6eTZE703J/+sko6YU6T5OVRR21YziIZT
4JYWQysf0m4cmrTsBG2okFkRqE9erlODuNoxOKuOfe1OIfXoE9XdbZEiEfQkrvpBuBP2LrzPMSK/
8scBgtzuRWqqtTckWaozT/q8rxFuUmA2XGY3cLET4VgpVHKH9/X+hVzfuQpHJoaSpJ8vZ2IIKx9n
L7XxG+6/faFf9e8w3+wr6mgZnCmpbwDqP8TWwxI+tUEEk+RYdLzuLtOgE6DL9OAlkQJE9RNZEIqe
NUK4tweGvSa8oKXYDLi9FzhnmHp4eq3eCuEDdIeqvqR8gVoGtVJ9u847B4RysY4evSWkdtlRDA5F
5lG9hIPZER96PtjLciX1Ehi/dSF6k29I/EWVbGiBzSPZ8wkiQBFgEIgA2uKBTxHzvaO28wGoxVmv
vcgiVOQwUWm9IgbzSixKIbwRYfGn1KSca/2XZUU1/ImQ1X4v8d7RCXE/w+LvQxGvsbpT8HNsLJBr
p8WAc4iqaHSPOzqJGCg28cyVmrWiqKgRHDsRPQr3vc9Jau71wU7pj2Iq8Acf5LNkj1ziGFeDhZtO
F2Gq73xUsScQYUUn3uQpxjaqw1vJT1cPcSJWNxAdAjd0kCC/oZ7euYO01OnkKO+PAyr68Ff8iuvE
MsQUMWbV+oOeR9tk7DJqVijNrmE/OcOwxVD86iASGd31UNXRiNUVliopQP3JZ6JCD2ZpkNugzWp6
s2oTMrbLpt4YpjsjkZvIQ01vZsgm6Tp6SEGMscMepXNmhutd+77eOSCX4G4gUYvE4C7RKui97jux
f4LzULcsSH/cTIhDMOFH5git+hEvS+IHQ5HZ0A68SRuVg1agJXr3go7iwvpgjRuVRFgJEmDWexSd
IYgwtS0dBl7WyJfy4aY7fxjdz1xmLcPQfjZGLwkKKCwVtpyAry7DAthPPp/QXn0Dzp8Zfa18nvJ9
XgZKmhVGrK25LcK8GW6ZOjWyJYAP3zfIvDb9YqdqyE/pkPA/bA4921bwpks3GWkC73akP1/Pi9W+
elk1P9quIqxvPhoQNz5NNrKJfd2THsrhQSLXdYQpODufK9Bz/+fujD7AeRN0npTXiQRyXWZfZyTy
Ak/A6nHdi4k/Y1/HyClXCqENegYBrd/j4pBpGtpT9LnBLlrLT7Qhl0NG/oxt1TqIa9u2vbrakGSs
S7S448KLA+IgmR5ipVyZ8oR2l2fPWctfEkiMAhCdBnXW1iVmKrmfplybRxgMGEvYVxlV/449DZkG
5yMrsziELW4HnqcaohEumJySlTPgxLxV5SUj+M2iPoGodWi+PUsUBLF4thp8k7IDC/f85PsmkRsW
/xXvP1FNeTlO6a4FCCyGqQlAPCx8vvYYI8d9Ow1+uqtgT59H9vkSI6WWZQHL69ThL9g7BmuGmdWJ
wL4rwtEqNJqRsaQRp9WikWN8vXrwI7+y8sal+RmYeLa8MpSpg/JazcxkForOpl9rTmjeF0fhrk+Y
Opfp5VzHVX2m0KMsjSmb+x/tbqWzxKLxC0/hET4ZYG110wER9yaUIuI02yloIlWSJ8pzDj1kOAUW
I1T3SecOHLc2T+gzPHKy33rrxLr8AQF4WGJWKDHsom7fN0cQ12KsXM1UlRU2p3VvFGXjSyEtdvsp
fCFsoLUgC4OXIkmz+oL56wX3i5XE4Kq+6WirweeeHjtUaS4p2QToLgQXpmmiZ0eARQzv3Pan/Ggz
5k1B6SJLZqk8TTELnvRpCJbFD7f/89cFcZsaJI1HkbsWt7yJI4rEr9/liFpXFQy4HQdh85J9Rk4t
awMZxOP2Id5NvmkAg9dzAKwvG1zW1mp1mAjKP0GA+Hdv0ejt8heGyX6tbxJ5KOtEm5NDHvxChzor
Vea4lqBNJUkYslzpaZ8ucj9gy2dDmXCt46dtJ7Fg6ACtkB14ksLscKjgLIGL1Cp/AqWMqoHq9/iV
SscYOHIgk9N8EYFZlGTlMTcyBt3jJFmoT3lqNaZSH0WAxkkxQc5hl/my2tz7cP5jLTFCJhGf/9Vc
0xA/9IbTYf5SHrI754S3Sd2OO7DOSgF41OtIvdEcLbIXEiKr9Vdgi9m7DB7O8w51SaYy1YoZkNq6
KHKtZUgZ9fTRfRRxq9aFwh7LQw8F3kchHS51pWbAU7Y4GEzoi9w1JyE02j7/aLmAwQRWnDKHErIT
fneHS3YlS0wdVy5QqbgGTBPAux0p3SeV0L3SWpKOWC9TvIrSEj2yfUwShATY6CMas57jnJcZ51OL
r9QQQRfqg9E4xPkvbKYd0HI26WqXRSDDoWuga084vUSgfTZTnITMnCyjeROpHIFdXCEcawwxqTaL
aYjsPmyUsG45RH4dq/JGOD4jywGvV6zIYwJN2p8vBno/hD7WlxmKUPze5ZoAlTYCyPi4oTDla4Me
dDtDnJJ5HuDTTN1LcjxP9T2cNQ2kEZYPeNo4DHcRFKoYOtb51TBGo0eVBs3SNko7WDTQEk5QRksw
2LKjj6X3OFw1M97aAE43CW/lc3uimHxIFN2mKcJ4mo11Mggos+CFz7GsQWEMesiqDe8IFnebChT3
1SOB7wQ+bDB6swdb9LCvNd+rhZTLVmvq5RvjjOEIrabU0KEXAoUPxiW3MVnFR2mBQvMGz5ii6ni6
AwlUJJAJtDZTHEMaseGRMrXVw4bgUSJh8KxGMMbepDDWQxXRZ2xsPzVaX7QNCQWNREJDY0Ajf0dl
qqUECcf0nAS40xrvmluZcbzPbH+Q1fS9PCrmZ50ZRwrynpcPz1lqZnOSgZ+fVO+LJsM6yMuoC2Vl
9mBJ9fRZY4yAAqmsfDvHBEYGXIzJ7dP5aMBisRxCXQoSHsTAjpRzyT3y6ALYFd/5k8lqsqf97VD4
hj9SUTCPWT/qXPR8zRv4K2Tljm6g5l6pl1f/1qSIFRFu9FJuVgpsrCYQlb56epFZhemO6vDZZ2iS
qEgh185rLLnLUPisH+72EvdzsIqPB/NHo40b/soLWwrNcic5kNcJ/peQFy1qAGD/YRke9VV+L5im
N2SFKkI0aM8N0bmpJXs1Rx0Jx6xLGKH4CQRacZwuz5nRxl7W2mXHq0FkGJagVWDlkrtXOJ93l/RU
/8ArZwOld3iuc5OqloJVWBUXpXCv24fj7w5MVxSnp97OTbz7k5yY+t6rLu4foanG3o+pNzpPNWVf
cWH5cWkT54Qp1cAAZfhEo+8qKq5qoE+A3iCMSypJ1zkXmOD1BTOe9NBkjKjmiJ9RJOFJsVArzIvq
MrnV1OelIkxK22jhDXs6dU7VoxAw+Fzr010BgyR7DxSaLVBeKemlSFccAGABUIcDODGveMwvaHsh
gHeibWJzTmc4bBp5euaUzF3B12AD22wl2pmSffeI61wY34219AxUDdU7YX3nUg2xaSSrzNis39e4
udL5rMtviEENA2fUkADn5Uds2hn8gg2kcF1e+LVLiUlL42/2MpZI2R9xI0K0doHJsYtCUBL1d+FU
Bzk1dLvQ1q1wBlZ3cwpVj+qN4kU+Tl1HXl9Mot+jKKk/99WbQw6rjaJeDH3eXMHKwOac06Gh2NZu
/mD0VnWSo0Gu5scg91FaBYkywzvPIUGGZbdHMGrHdz7jYkm66e0l3VUSyImzBQb8o4Z3a8+z8Nli
ALGhASCmpApZmS1hACEb1Jug19lJhvY8PTvquUSn6DKGSYTwUyhnieDZcRkAcCCgx/4IFiq3b53A
Nq3lGKD/5Hwd7GWKPGcRKWQ3nMUoVI31JFQDgQMKvhm5tR9iUI5G8n3LKnSgku0btw15NpLIZ6CK
3vHMbIaXgB3VloKfF4lTJZk4+qMg2OPCvx60aKOkZT23t7EZ7Ks+6m/kQ70ydp/mq6hIdBaetAUH
KxS208HwJc1QY+PIqkKWH9AMthibvCgt3zVSxhPo0SfZMt+4FDAJPqFC0h85cQL2VQ9Ry106M60H
09xbKy2P2qLOKLnstY/nekXoPR6fZiZxwRwsWWl9d1BravJAANMi99tZdoLaiCoMx2CLl8VmNZq7
FrpAGP4bpB9v8fNfF3S3roBF/nwcCPRN2EeBWG/rW59MlnignzWVUx6dmxNh5q096bC7K7XG/OMy
25dSEarqf1JsaiAPSd+HLOantXv2jjl4h7RZgtWKsW/VTe0hrZLXvJZzo/OsooLEqnTPg9S/gSc9
tofElHsPpSAvzgr78FCpiKL+TAq8Bbz4J7UlMlH2TokfeLTsvHFt6pd0TVXCQnonZW24h7MhqnS+
jIHTRvTQ8EVqlY80nX48uI2baJY0sRp7GzkAh7mjWlC29W/ffcTyfJKV/wsKgWlADRR5PI/JCFtc
zPP9CqFSijLfCamsFDrrdbJDoL9fjTBCF2SGLUUKh4t7ajJTqdPuXme/vmRqZD9Gjl7rfsjEea2/
xmW+uHYx+L0GbgdGQGKegUZKncV2Ug9sq55/AWKEbtWpT0GPG5Sev325C9dH1XBm1CUeujnX+54w
S6Vae7ih84jClh+XbZRLnSD40e384YKM7fCdmE5qeksWmRrHo1GSilIl+ujz7AMJmOjNY1R2YaOt
FHt8R5gJb+XYG+Qrr3E3HR+zakRMuak9m6Uja9Rsw2mZ6unkPYJZ1lICGod8TygFUCuAv+jhicIF
iMGxdDa0ly3KyE+HgfC5qEH5svehrS6IEi2S/60cyNf0jByIiRoubLq+m68ibqVvBBOjUpbV/EVk
liYdDhjpD8aLEuhyZNChUN6ViowMiApFANP5DRjQTXVSp9HSRcguWrbAY1LMMyn0tGrBfNU2/gUA
I2hrE0O5Qi5Zr4T/s0x9+VbcJdRYR+WNhVuaUbQBC36UVSVaKMgYtaEgK/CpKCSQCI9ct0uRTwHs
S+MDfUUwFckQFdZiPtT15NT28Plmrrjhz30Phs6aV/roU2XNSLFHNOXIvjBdazE2fe0Nni65MQYY
MY2YWPnWPip01FoVhgyxzO5mvkuxmM/nmO96+32NYbjZdFxYH50oRqLiJPB3xyX5HQnKe4Jhc8ox
dCzoLcBB4hZ09xmS8HEzWM43Fw9otjdWpOsh0/ajba6G8SxvZSlwTzpMBeh1QLj7n+xqDfe5Gyj0
0aOap1s0dFdzPgmXMEWOKtlddSqUnWANr3kdRQ1nFGwNgfvAdd5U6OPMagqZ6++531IUo++uhLTq
GYXxKrWpalXOfaTCllgi+d2/yNraVBtBD5TXMVkekjG1IjpPBtmQt4K7Fds+zOK7RhDSYYJ417PR
cxMvJo9ahtXRh91tBM3jFZMKZss2lalNHOx26CbglqWNLhnzenAwXxQvwJaMRpPUB+Hz3iCX9aDx
WRWmOI+sHCimGJJY38iVazcNSN/MQPg0KBtwmxL0WGMw6XsvaFcVIc4E8A6zQTUKmzQ5Q6cl6VnB
iCB3GFM+66KtZ3ThRdFXX+37zd2+ZDyXIv4FdEnZjSKkabjBRG2SPzkyB83pWX5AF99IT2rPZUWe
a+goYqvC3JDHdpVEdKvIBpcjh1mX9B55BrkSE3sghv217H+BxGJcQV2bvGDHvcVbXwkg8HQmNVXS
NOnSWlVIaibMc7jVQ3zXalFihENis1FZrscn1lZZsLort+WCYAamvRqNS5xoTilx9ow/cVZVtxki
CniYM+Sqq+yRM8qk03Lfl4a3C8LZlUJjPQZY+v2GlJ+MzJ0OvEUSGSVaatZErcrE9YiuRPXashAK
pcI4VBB44hrW/hTvwYrFF3mogDCsJ7+ULo9VKq5k5muFi4/mSVwkclCmLqmC2JxAT9E0kHIIOcLj
Yy8mCZZjy9GjZKhEjmQ2FQDq0seyFvrFfvWU0JhE5dp+7U9vLWo3/DOehuwEbRZpK6iC6RW7+f3J
rYHgL94UYI2EQbADeHOjq0cSi+RyFgffbQeld2KiQA6B74aK6gIGNMybw2tT6sljLkhqfGBC0/Uy
ckmbdppZNxw2VvsqtMAV58Pj7eGMCKFV8wknNXW/nEBn6XAnbtejwz48dl5+FdcmEbqIma6V9XeI
YCQ79mqyWhV7N662IL+daM8qCh33He476gzywlffbM0KjSqM4ZUKB8P3fSzF5BEHE45kCrm10nQG
RUWX0TG1YhWmnxfUp7FY5rrpM6ggKuXAaMvSFk1FSf8h/5O8wWR8lBDIqb0ZBGlQoMNpQkuPh6tF
5emVNLx15EiWeRuX1oAe+B7zXt+XalDCGzv/IOqf9BEIMJH5y5V61wT2O4rXJokGp+T2mp9R0eeW
fCI1yIvfO2EPed6h+eLoSZpXYoaJTjrqx1C8uIQARuPFg25eMMpQ0M4WKhQYKa3Qad73FBJpOHjF
4PlOF+codN5ogZ86aRILZSzGhve98du07APki3mbrftKC9TVLYvSX1pp8eBFsodDoaHYW8Svtdt3
zd8PR5fotQRL1SRj9fmvUX8CnGXwOlGK/T1JQ5z9jW2cGsleTql1RI4+Kuw4LL4gBXG2/a3P06WD
2YGixCLdbENRKu9KrcX7hGIRPFhe0zedaL/ILkfhhDkXdU3bXRVYftE7+ZwhWFbq+K/FsSk7kpHl
WXlBukWXyG6KodfcKKfqIKjtIJ1n+JAJv0/Ctg8PiOFip4iha01yUXIB6Utug9cxydCFT0E9tUmQ
9UpikTCfK7VWfFReXHe5v6w17V9HQ6jbnprO7QBm+5M9GlDiEwBkk8+eTdNxUBPllDPvWtCW0Aqb
8syxDu4mwlipqmlWQvUHzVF0V7RgXrwmQUdD8vxPmhuG+mGe0GkdoqZpjWc/qidDsYYAZVqis/DI
bbF/KEutYMZIGUdFgyGkIU2ZuLMtd4mzKT3DD71nqYdeOzTsCMmyU4gQGio0+kwloP02r+muHcGp
8qwLUQc0g+UCtcwWuzlETR+TDEvAshjyZpARpbgaf++YFSAlBNvpkD76/KktO7xowz6O6XVsIKVR
xKQ55HCYxblqbNC7NfsmA3nXFCVAfbPryQoZCGXYrEdGj0mU4JuX/7RjDeTmakbmWphNBvvRDZMT
XEC+X9nCGU0XZKXV50H6g8Vz2nxwJ4MH06C0bNjmUrP62+TLiUOaoEc2cVIfThleHLIM43qcdHux
+oCvnLxunyGyZVo1JgPz1urZyshSQaTXqWZd6c/oenrwJNsNKtThKCUJWSw3tNKQEjXImQYZaEpO
fmYijE4T9UCsNvyHZedKtAumMYjZIs4snxfGJHIydzssz6ARd5BkKcCcj5DJ/byXtCCsbb5yTN5D
LyKERnBELshgsyz3IAUAcM5c9JOSWOX6AaLpV210fbOZZbk4nrnm/a5nRdFUwfW33p1jX+MJgkHa
55/wibpWEPoGyi2bXJGg0aE2ci7wxWm98jAxsK4f5XO4PnP6BxmnFSp/7IMoOC8uIHOTKqaYZeD4
LQe+jt0Mf/LW07lfFVPZdT0hbmvoZl/iims0kcKf3oPtl4niK3knoMVtyK9wPXAK4ZXneKsP5P8H
aXEWMMUBmsPU2LtRPuNiiUPDX/td29NQ9100o5Otl3AdLGSFCvfE4eqTBjBrG/in+TMfa/6lql5E
Zp+NxZXzs6J/lBFGqSvqSa4jCUZGT7YFgJE43HM4Z+5PnTA5S5pysytA5JbbMoxOPdV1IfWFmKXh
uFBMdmmSlhRCFIAL/nRjBqVdQtDyBnucPJkJ17VgrTtHMlLtMUHA7W4ZUx3q9dHbV4jWoG/ZfRz0
luMSMyXOO+A4TgddF24T5EkunC1PedGJbCejOtZQ6VbMcWHLuy7UBpJ0aKad+bNBmQsQ6/5TIj/a
Tbf4UU0PK+ZPokYIP0OPktN98g9pwsEbtOJt9VzaP3gtnLt8lpf3TlkV5O/ulFgwpHDxEgE9S1PR
p6SHGI3Aw+HW5ph/aLxGbCZwAJHShbGSQS185iMPBydIyCtDRt6vtg6ZISpkIpY/qU0r03Q0vhnA
2OuTLo9uzWO822rKY5OJNDFaFOrvPKr178S326xASdLvFNzYXhF5HmuhOdt9BC7KLL58GizVAiEB
rSORd5vksoAjxhmNqMkuj7WsgPs4yWLiinbL12GfrY4jOnDlxf7d//9MG4USKnlJ9uqJDWcckUB9
Ackwn0scx9UfEl4hlnClAOcIa/Jni3W+e7C0eUmI4e0eLYDTVDaACBhkuN4Af/jdPdfbQM0lzut3
EYhiuhqSv6hlIGcQI+iMR2p9e7zs0cQYnyQBvOMmIq3DINKcs1sNXwKIbBLF8ZQEfGblY8ume/Hi
fdRMnTu2LsYucUccE73g0Bavt2sjqGAcTynDtcis/w6b/OnV6c9ngxftciTpOU9hr1z1wpHxa3zS
TziHhSV4Al6Fc/ifAOy2LKobFByH4hRg+JawY8gbz+wKlMrT8EdgsYiBRrcLG7QgM5xFTtn7Z8Zo
4GH4yscJJAVrtAOwDDntXrwmFiS6THOq9LtnWHnY1J7ashUtbksF/1B315ElwB8c1BVluXyvS9Mx
3OxbRBNCvu2DwKMv7vC6WQjf8fkWtA2u/xnIzsY7mWQB0DsmyD76D26s1SRURhM2ssxG9Y69smxJ
xlRUUYcuOZVOV0n2ZEq1728Jj3Pbgvfdod9TVP0Usb5XbneHs0BVM5n8DEZAkFgRNthFnidew5Av
FXWv3DcmIyjJcGgdE+3tb9H+Mpkrh0Y5Ra/vptwO+03UaTv2Mipfy7vMGetvtx06N7gqJJkEklXG
RjEsBJkHI6Q5UecOSIzxVIV1WflCIRPXopw4c34YS9CLTavZLrnpUasQ90GLsFxT2+LP8fDw1cck
HTQ1TPie0Z2XDi2s0mvbCnJH0DC6zR6gn2ZJvOPEAVp97LiRkv+ga8vqX7UZCO3xH+xYMOE26Q9v
lEYR1IiPDA/B0yBb02ujVOJiL2NcaHr6nHkWplGgPMHBGuqzgAtDu14aJxq6WtivapFIFjVmLn69
Ell7yDl9N0eDrbji7UyaQdn+kxNFc7gcaXjivmruZwa8aYT952pco2Yh9tVKfS/n8GO3z33/oEQr
3xJM2jZRTj4QsC61R8txXm28/aHhfmp635JxlB1eqWjRA5zq9/zstBXyv5GJjHwRzSg4wPwEULnz
zdDODNRX5WjwRODdieHs0EBJIuCLyfLXCohD9hqAlIvjhqyvKIDbAr8Tcucp3oZvWnDSQuFoc4I9
9rH3agQfa9xNt16RcBsje/viFRmB0Cap6OXlmemEDToqCGjDQoTi14HGT6Y210+QQDex7d6sFa4x
t0p+bDik+6S/37w8hJtlaitBeWb/q3/nitfXkaXEiJ9w0LmEdggOgsq9cyUfLToHmM9h+itKqyjJ
NHf8oPbaNlZ9filgfFa6+J3MjVTV8SHgdWwKnj85LBOlTvKuCnyRBq5wEINanDqP+Ti481YShCgb
o8kNUMX/C3Wqi0mrMdMNiONfgjQw3bmYmN9Ca0k1VVYNMLOrsXCAX8vBpmrrPul1uJ3kKvVp1GyC
ABbuadNcOupcI+BDETuqgBhiHXiu9whm45Cil+D0yrknylOdvsefa52SCvJf52xUXeZvt6cxQwJ/
rdXDAbrb98vLzItcgzuPVBp8NrU+Xex0fhmE28jVG8J/872PERZHSnf3k/xFcZfvZbggRdozZSPk
AKFcl7TWwmXDNIxbfGfd7+YSo13rh5Kd7Gt8Muc9BmKp7a3/2SYnt/fwweHxl5HmYnwtWkEOfb8Q
orZRcJ5QIE3VvgHaHFt/3t23XDu2OfeARJOYKGUlRt7/00/b65TSBT/lef497ZVKF6tX8yNrO14C
Ix1YWGq96tbKauVlNBTysidsUeQV7fPFVhbPcnEoK+xzq4y8f+2J5alv0YcvTEnZW8V2C6K4CJMI
CABKDsVrwWWo3ezlrarFjmN5kdoThTLdgdtHlZ0OsSM4HgdxrKoPfkRFGIDjcBXQabiHNbbGuYbR
JMvIaLFyl1068LRr7/kyu69/X4e4p1uSV+9Opx8t68HPBI7n+45HZj2MfwYPy7MnoS4S9Ent4l46
6623tNFZ1JsA34P91z7wQ/h/U3oPKTHX5MjzeLDfXyJjLzzIzD85kniJfJGqfYKHK91Gfcx+M5c+
SP9wiEeBWJ3/hZ8H+bVvA9reFjBhM71YvySaIo1THW19dDh1xpdENJaJlbxs/xgzVi1nycETHihw
Y3KiCTO+VvLk+gFglzhZII52HNcJcIEPwlOsVyWMNrgfTrZrDi5EbWeWb+uOqHSx1A0F1YH0dZmO
WzDr8HKEbF5gjThfJa9V0OwAn+eag8E6gMb0PEv7JqxL1EMw3bF+m00c/W7NXT81DkSIfwRcdITJ
NJ5jolYjZMr2urK+FhZhoEmUwThSlji4a7Hca7CpDWj0Gu+acGmq0XRISbnK/viHOeYNs0zf3veM
aQ+MvONKS7mitRY3kvV1HydBUdo2ls3QVI2+ilE+GITnX8St3qSNShutgsYgCcNA4hy6aAPUK+ot
crb4A/DRXOlmcphUOMmSeSmPLdL/x09ekQmiC4Rx2eiXCfKuKtRK4xJlDT3ALItD4YvEZ0JifCUg
+xaLLJE3ZSs/Wgdv387PAKcJi8vEeALADSw1ypjcDLND3G1FvicDC4VoIiX5Aebq3zronRbTxRxt
HoDOAOF5ekC6bmGAII4UwWvTGpkuLo8tYQsVmvrl+7Ec8L9slpJ1QlBkJFoGWvVk1Axg3ie/1Ib9
kZN38kErLjakeKB+HzW4PFheIgeO/PZPPz49r3cdFF0VXmbo+P2NQpZNQVIixPL0zw5lBQJpd62E
a69/PAp/ZbZ4BFmH08zzo3eHe0SZD7ZVsIJmg01PN2ekn3KjCXQaJB5ofphPmWX+YoqJD5iOk4VX
UM08M45T36aLv+dHC8Y7bT1rVYWX/9N5zLZRx2cEtdCJxdQ+VFNu5cympDH3F5JYOzcI7TMCQW/i
7D8L1o6+qknxs0S6vJJbjAs4hQ5WtcmlcOc1t17AaZfh6KGqtNBPBmQMOhUMFlxAZSCe9so115U3
WVHGqbUO41lwI9hSI3LD298fTJGBpl7dL5uTsyVU9JR9sY//4dW9DR3p4JnICcJBw7i3YdYW+cEi
S55Z4lLMPnfQh7zuNopLD0dlSCFREt1Dzq6pMMg+OtPBpBwpUXI67y6XW7yjdIHUvNyBBAiFl+RH
z4k5nUUmUystxre33efiP0/lLYtQMoFw/NX6+09YpP2HtCCx+BpmX069ASOdosetdGkHdG5dddCE
308E4NbXPrYiQ6oTy9gnaI/pYZQdt3ASmkTBqR+UVoWJp8gcCwcsSssUiYTtTGli8q9H7jpVWtRp
OBgdthZOmMUVpToQk4qZ8x8BdIQv88hRWOECdQvSDsm2ucbkdHm9YAVOdlHd23VnR0rkhnPV1EyY
AhbrS/iTzFzoXCbV79YaGtH83gidMtiWZZfE8x4UBFEpf3VTZBJPz8dg7hQmCVzIJNwpu41x/FUd
pyqTz76sHsIWWD0ghI09zg08nTADerlY1yzvzh/W+9Pi6UrIZJxxYfcjH++acpx9DdsNrOL63k45
QhBDCmVPYDGKJecL3vM+4bi1j2n/xImlfIKdMxw3DKjaDB/TVqQj0MyxuOBmoli/6bnIpXggX557
WIeEAbvWJlcjeS7WCoG1tOaT6FqJUQ4ez4KrVpLG0CLdpl+JoRkljQ7b7Xbx5tA8hbbFQcOr842E
/6AvbdUkFS04ENlbFO5UzATMagNG2kL8mTxjIAVp/pCx0sDaM1b/BUA3MszTZrQdRVr4N4bXccv9
eWqiWD58cNyQ8Gtgcs0fFpJJ9ad3Vyl4niUGtYtj0Eybll+FXiSuhd7hqjcJCmASDUGYjSyz8tnK
11wFSZFHkTZ//paV6JZveBM0v8Sqr2iPf6XASXiBw+wa/i8SwNaiTina6dUyoF9FEs+VfexkmyH8
WDQfX7sBQukmCEa+ArMo0/bKppzZN4yhdw8uWbeBb9cdgZKe4qa8stBqq73w4v/Esgi3xnGcEWsK
a1plJjx4nuFZ0QSvOlJECuEpVcxbwwgkAGmHh1q70C9BSmICKl+dvj8AdtRovqvHuj7wPKvOE/7/
/qJEemKHoqueGYOEJz85S0izJgQPTno4adBQNamubmXmcA8HgzjuPBLrbYHpKp0WcayRG8UUQhxf
1HoIq2kve4/Cow7hH5xEcNSsBccHSG88a81oWzZKyRZ268kRIpmLE26wkmgegeougAbsHrcDSyzS
R+CITjqdYp6zffFXbnr4i/RSyDnhRKTe2lSadMT0gcJ8xj3OqlGIm2XLPflJQAd3Fd0NijtRRI0U
lMHIR6Wiu2SVIkMUUTUJ/HVH71SCGYEHGDJ42/whdIygGuAAThsk2GXoK9mQJQF3fuu9NsSmMXIg
snw+g+ofuzrOrLTLyTgkvVk0W5DUDicRsb92TKolX/xOXLsbmUS7RjmtFzQUe0ZIx7UOPdMBwBEA
91Okwk314jKvgbWzhLMhhKMeQ7qpa68c+3Omqyo0JL7A7QZhcOTxinXte28Ug6kCqUEXxZ92ag5D
AIGqZakbmSX9zVHKZGi1GKiry70yb8ctxPdlEwiPVtaEEGZaoSSriS/7/4gRXylx5p499txBcgtu
50sIbhTtyhjAQTUww1nsX7EIth+oTVdDKziSNSbDLebSaEqw0dJukh45IBWAMZ4IPL1+rnqOXeh5
jn38FZp6lIzCWcHNScf+97GvOt6E5seFL0lto1iaKEoNoc4Z0GG6B8d3CdDTEZjVASS7uQ8F33wB
Noph3bCILczpZgEehOH8/Qf6sVroKNNxq3RBugmQ66nDXlJZHphZg3Q066A+FHqjFGm3pfMR28Mi
4E+W9Uk2Lhrz0hWuBWBWHAybxc44TvwXMu6YGwNr50ZwnEFs83GlIZPoZstLVAIHykQXoGIp7tkU
AI9oeOBpUCTR7nNTzoRzyssL+AJMrAoMkBQq6JAkx8mGAoMZUCfdOpzmRk1tpENAcnkOGT10SrFV
bs9uaZHvGVOz+0mATKuTxjUFHBb5fRd/lIMFxhdJRNA94XR2KjwfAljWaBnWRmvx2cCpg/x41+Dg
nrjhXLEZ34zCy32Rtib7SrkL1zScIWII2rIpYWDz0PWoqG/vxIkQD1nTNkP3BBAycip0T4/lD+ql
fK7WaNPv0eikAQ5gMNJFphcIIb9iB118Ec6NAYQBR6rxXnvDKaeidsxNPhiZ7BXFEHkZkY1B2glL
kckE2LoFV+jXIlU5ZIpiW29W46cx0K8jOMH9QoHnoql5voHP0TTlHR6Fjmjmd2pRW8OLlTG/5rMQ
pCTxgzj5ETWrrDEI4+AClgp0mY4V6u/nFsJcE7/L+EdZJpJgzLUwro3YGJM6pqS701Fh+OJrbcKf
Vez3kLLHEg3ujDhvgNQuqPUyTPgOm+O6sw8VbdlST7n11z/Qxf4HIgPQeWggO+2DK0ot757PvGCj
nABtJix7XIu6z9+JXZVH2Ele1+LmehkOYaOSRfaLnAA4gYmj5xQKSqEGHW1luHupBrk7ahCRS7L6
At2X2rQZ8H3LRs2SMxrDPun/aAiBlFLdykc63DxXM7sl4y7rWtxtc4pI04fyNKOKXsqfJdlPIMH8
HCzk5/xJacLaKmqh7Rs5c0XiGqiZQ5mvKsl1hLwicfuhq2cyDqUD9c3oUcB1kZAsqfy6/bR1P6ln
QYBLcArECev2cwDymAyQ2WylyO0SsrwHGbXQvBhVBiKKTy9duPpe/BtXSUYNNr9rX3023M5/+s2A
yyCCT4p5fmQYQV5RLXvkYDJXriH+aTAXYjPUCx2YYM9q6ZazkrwBAYlisHm1XnCB7a3R855YqDNJ
u4bzPFnLRCpWTIYjhYJLp3RQr9ybDzf9z28Drxl0BDDmwbKvH8C7sdcI3Y24oL12H2Z/ChaGL34N
Grkh83KLal4fMeLyulpa49fXr1kxGVXtt73IxCyKerzlcwdl9zCFyaz3Ybrbz7qkvd+PQ+5aoz3r
OOtBc6Ig06qFH9scCEU0FvenAgsmjEGbg+1s748sObHhIztU87RpoWWiJMHcxg/onVXYho3s6AcC
VToRX4KnB3oyO8tBmkxBCn8vw4H1etB5cNzhDMKQLyHZEuj7xS9OuNgZzT5cqn9Wq+6AIiO79SmC
VOegkP5oL4aapPQNzLE5S2iUBuv0YW5aCXv9bk0HsZVqt90YxYzVO/YTy/eRfNpILGyfIH6d/jGy
5e6N+fz5M1bUAl/xxSnmib7TTFFnY84tcYzkBwiZqrDxctpq8fSNmca3/OTxsXyplFXhApMn9JEA
LSD/8Aw/+T4/MADE2se3PgJ7j2XUUs0rvwa1unNt/cqC8cR2XEGg2hRrT81TJWEB0Wvh0q2hcf2T
QU2rXWqRxbE5ainakLrgRozD4R5kmg2hzsdpKWVSVO2EoKUVL1SkaEs2j52NqOg1CRXhbP2k3dtg
NsrFbYpAl4mUUReTyVWnb7d1qJOBAc3ehAU9/NsA3BaOQHVXoussZZ2Gsvki5j8u8e2uCaLkJ8jE
g2y80VqJKoRaAxki6+8+2lK3OPvWISJJ2MI97BQi5bW3FT8GTdGXDwiJlvEX+VxHk2N2dzL+OkXE
/rt2aKCr1QCkubTCc/az81AT1cQXrPNlfb/J/Fed3IAC5ks5C/FUhzAKwMV++/v9kohgTaFLCd2w
78DhZWgx1lARYyk0YlpVNyqV874FuiwtjtAKld6SI7T8U7k54drKY2TX/Y5MbVsNH2FDKGn50cx8
Db6fCvNvypNGJ4SFaCZGOhICjAAkFaWBC0MstL/Y/raA4Nb+0gzQ/UXu08GpdMPaoOHYs19WHiFJ
T7gl+xRGQTiav2IHatUzW/IC2ixLjKDl4HKG4QyKck8GEiof+PoA6cyc56XyHf+8LNWQNG7eVjsM
Rpsx9y8cJ2at/9rSFSL2l8S/Jnei7Me1KA88uLur6h9UET1H7S9+Z1GK78RpnUFNb8ZU2tubpbcV
/XVS8Sjvrx1hNPj4OQg523khm5LlPzcGuPR4KpVpY8/eGYrRRG/aSfJZrtChlm2Hkea4mQMkOnMm
yRnYYQxH9U16dBEnDjoTMwtm7lA3tdMLiPSy8ZTos35/K4CqHvMK+3CTFvl/R30ilLr+OU1HfOIB
r0V1p30ff8HBjOEtttQsB7qPc8acWIllN6qTkzUcwuHm+r1Um8vizsxoeMuxJjjd7rME/CBx8oGZ
/NF/odE++3O29LYeUAWbO8ZkBx5GgH3fXoOHy5jn6KzSE5uKhoTfBRBt0bF7XMmlAkjQNskxomgo
o1N/gErM90qFkYIhX7Sx2bvnKhs0BNXPgiSFTzGRaAlCcY1BFZcFVenPJG3aIKdUIwQvdE9Br+Ve
/LkZ1+aOP6HO7cx93TuEGNaXjNKsH8q8N3kPACCCqNiQKbs7RdHMVNegQtyJCKSur20RTVFZl69j
YKH69x/APhNIH3pyALNj6YWmpt5G1xQoVT5ZIMR9AEvv8udM6HAdrH52k/XM0nrJlFam6SBhOJ2D
GUar6WIMlOgI0WEPbxEPC16EeFdolryUPZhFNHzQ55v92HxLJUFUVSKPJkFuDDDL7e+kkAniB2fw
fcdtisr9+ADiWYFxEaQtV8l21KKCdUmJ/Sg10nm61hh1eukU93fUP2l45NXPpEB4P+gtDWQMv5vE
b5bih8kQARNRmhDoDId9h+f3tKi7pegQe4vePyvspjwMCMcUlEy4g8gNiCS7NwT9ywdC3EgI8em7
dg5ZqtjqiothyP5p4iCe2zbJf0VLWXsHRlYTsD6gA60IR/RcRj4xJ3MoyNf3bzXq8Gnw4k/Jka1z
ymkqw1stzyTNx1MjOS0UCEpC9H0XqTJzRsvRUzAMpFuFBsh0m2hCJy5qvmsS0nlTL1lClP4YcEoI
MNRk98qtnJ9cwoy0OgOvOUdVPN1ckqM+X6wv8WzqfwEXHmC8nUx+XcLDG8TLpDmD8azKXeHZIIZt
o552e4B6PA6S6Wc71Hi6l71b8ncdbg68GLJD5kEngWJeafSFYoWtEcfNE+wNrQ16WXlGIm1ygyHX
TJ03CcsoPgz7JV30PZkUvNZt/YEVgAzrQChRoLmxXyfcrElsvpV23RC0vctnCf5Q2ShjFNRuxoaS
hI96trB9OmIDffJTlpwNa36HZNI4pbxx9FoJPOmmhUaResorAFiOq/LLEF6A2OlJOEMv69M4FRfG
8xjRQlHeWvzY4c9/ncngy9+fdvJsUnloobVaaqwrIkUrwz4jYkk0qZg0DicTkzESjUF6DjpQpjUh
Bb7ql3tVqxe1wv68P6/eo1B4fi8bF3uuAll2rgLNgM5uTe9PbmOzUiOh4CK7i/5vLwfU/SWN19Js
AHZfW0DibQF6CP62TbxO03BMRdm6wi9Penc6FQu+LyjSrR7ulG53j5ePJMt0agDmTBFRKkDGvjif
4P6tsHDEV/eQ9FqBSoS/ECX61t+gX0EZqk+msu1eB1wMPARFiJjOEDfuycntiSrgtnEavl+YPnC8
VehYrYWr/gO0YBru5Jz6YOMTpC/TNFZ9npaXxivhFYOLNmoLbdCG1FDmTUnkrou5jga8kzxEh8Qj
GSsD8+lFKgoScBrAqihdenUH8EBEtMrW//HwI72Jf2+3pfidoXDEESaJPQuJUYFVydY9evxCqGqk
x8nODxEFB5M3vSuRw6ldp3RjwXG3MyywBYl5XCPcjfza/Kmg8HwU9xGOnrEfZJmCgnBLkcrBx0aj
Ye4JzkZp4hbotoHK5zGm3UIVrZ2kzZ8YnMC9+aamiXGQHg/oO3Hf5beld3KjS3VJwfQREUNnu5J5
fSIgpXvuTSN0majDj3VoE6VVQPGtOqkyRFxXHMFZ2C7BBhnPUWOs6/+uBI9aHzgtYfu6LyCK4o9v
DtQ0l7WOJ9Cg0p0MUGFlePIWfsj1TLZTY1dBRokcRuERkpS9Z2qAeq8NTXeXRBTxTHMT6mq+2VTA
aN/xLO9wpfSeIyTBVIC77fDWpRGLqX69OluE0+20K5MJdYZjtZ/+DHVhnbt3kkVN12Wq5MquFRIO
cvQI1KOI2cl1z0PAeGA3coLUUbtKCYx5XBv1ynHe6jH44QmlCRDFlKxvNIv45lfU20p4+AWPysy7
YQT0QggJyiL0z6W9bHoRl7oyJ+w3XG3jE5P00RhO6MFXg1iKJwPXvrm4YK16QF25fRXYpkrUrdZZ
4FKpjkLUjhI7DrNxOCfy1A3p+3zS8iEvtYB8hoc0Q0/0nSGJ1zi8cQ/sUgLUN2xsghIXt01bpZgw
+MpWE1kx0ekv6ueFvN3FLA3L60qOiPrSh8YFXkUD9Dfp0Yf1xoNNvAotRlDb8lNtQImmlGGOlhBP
Bca8EA4nsxfKs/yq/WvItbMWdINi4WEXOji7fkMvwjX1zES37YEjDr9G6TBwY67wgiUArKOBSrgQ
tdx4BQExUlQc4Qt0cSrJ5IYEDeDINlNCbdAVzaD2BQUtVa9WJr4tR6+Sae2R70334uZqf81kY0MG
KXLmLL2OoEDahZ0URF30JQm4+A7XT1MswYE2Wrcf0WZm4dNJH/J5CA8Q03H7BnToIn2RtReTYDD7
0ViM/yOz3pb4oHG6FXfmp7xc9ZQ9zw81H+yCpF/TjABSe7Ig3e9HGnHgNztzj2LVL3cMtx6WOnok
TdAIoigFGTmw6XRLb5Q1Um62EJiESyT3AzSHw8s3kV1q50zcR03m0hpzmPFU7+LG3mBH/4IjZLYS
XNHcv8cCU9f2gCFfv4+CcIclCwFn9Rf3Ix70o2i0BGPlpTtRVIjzhSnXxJSklb+cj8xzozo+qrX7
qPmxENFyOsnm0EGisYHOUeqCZVHGgN08Cz0eqwDHN8H1L/g8HEbJJvKcE5Ul6gpJOhW3PPp5DxZR
zMJVD0t6rKAkPdwNk4VeXE++bQHZqOr4WDMy3ibRNY0V1yicmCjXCyJXCH7prY/+F3zkemVjt1iv
Rr+voWk/uuF0pedXrIPJXDX6arafyVILhYaD/3rg6rrU5C9HpnpqJBRPsGXOmJand5TdwNvc7Nb9
4n3GHVYBK/f/o+uA49YElGGbajgv2tBvYC9PcYsfMVb7gOjNukLeFO0cXuufj583Vl/LUmVshNtv
/X7Mq1kFJnadxxtQZfCAYV5kLSrHmMvlJNGXKy1ppH8/WenEti1w/cuIHx6jkNjKbtSzv41F1tOd
nYdPOIrJ75PeuNVkqV6DdriyHEYKxIH2toEVMmiBhjJaKFXtO58bivrRSKIfWALb4Gjz9d+wvOY2
LUUbrKz4IpnAVYW4jHv4WX2Pcf05vKvgkIlTsysgmfQrQ6F2XOpnghmQYL6GlYfiENOhZ2JMdAXP
88fIODf4CIcOm0mbY116XfLOZWkr6CoJgr8grUE/2dZ4LqBzpO7XyFdj7xn19caGfn0fuNvmLoWr
Eo+2E9s83zBwu+9vFor2dVySPUGzOXWnBq+XGxSwL38RInbeXi4QadSKtwiNN0R2OuqMI/CNL+zY
DQ0WGF3dmO7VTZtMMlb9XtDVVqQDbL6UDyYsXhC6Bg7cZiAZwK3XaFWZ6jda8wXcWpZCeK3QDfV6
61/00rsXeNf5yJRbkbyyOXPb6M7FAXYQ4L2fULE7AQfiuFyKi2z56rIoWDQTXNVJ9eYIR77arzLo
JA/y7eZDfjvVFC838xRijxRCHzNI4q5PBhQBXGD5GTJ+LosE1UJuCG6GaYLnnrZAFJFR6Ix7wS4M
pH7y5NgpFi/tpEMimtzeJTkfcf1m13L2USu6AEvouMJ+Q2D1X7UC5Ro4AM+ddSGtJHDpTum/SyEQ
WTH+hVb0tRZJrsni3r1XrGZw9LMCYSuLZAd/zEFKRrbUs7ADBsS4pm0CYsQz2Wx/yN0NjkFbN4Jv
mf8Ordpw5WdVtuHsn2oLafl2Tmiz/yGgsooH2V2hqgNaclGEconcy3PdYv+qbJmfT+pJQJFynTxo
WVfXXyef4DuWtaB10pke0ll0xd4mLmE/dFGe6kQEA5wHzvB7xjXgjnxtuyFKYnd2/ooR/EObDxhp
uFtiUTJfQvBW1RNtpAtk77QOYTJ+pUrmAKBleAFgjKI43dpsVG6jXEwxTXetRjLu1RDsg85HKdFu
FDBepLN84R48cR9tL5X5HUPT9DSqlNQnFzf8JhFtsDqumRqCrzfDotpLXtdab5Lc06pPfA8SSgOG
dzdHBZCDpIRV5IpocINRGPDeRdm7sBCA/WRrEtoenquLbKHjtw3uiq8lUjdeRoLzsmyPiaY53Wx3
zPH+N8JNg/m0BPrejRHnsG6sE08Fj4WcKglvrmh8ArRJCU2Rz7OzQEg1+aQRGYcGfgIutYuMPERH
0XKZkCCaZHHBJdYKJNHukKMNcCx4TP+IEjxlQf140da0bwWOuMF0ppuix71Ey0ixAQ68VIQwSM1N
IyMUwsmYzRhPFB9vMsqyUbgpaJzaR7ZusrlwxCjKrTgCfVwL+24bbjndT0OzOyPGrDPDcius20r/
NKHZ+8KKT2MXumYHLCGAvzu7JVzVnhnlCgrA9t9aCxD+H1jaxTC49MIEv9/SzAJac3+HCFDhNH9K
HA3J65eg2wEoxcXLS7abg5vdm65IffnC5euXKHxjOrOpy73FfRmZz4UcDagmJGAwVQFEqzBZzieH
kJZZDtZVw1EcpSFblbFSmUo9Iluw5gOZusb7eGgO0j2FXSjT11K1vkf24S9UVd7gUROYf75SACrC
krOjuzoqIbt5SOys0n1M/1NaWeI5Y6JxcUP6j4y/3UnY4QulVI3Y+0sv5kQ8lvqvBHXA4q177YXi
68d4lnEwQylhUO5ZIgJzgJirAEmXQDlYqxtiG8iITOzNBluEaOj/2/6KdIIzk+o/4ta6fuQZHh/1
yX43MkQiGPOCVublaMY7B03xiNroSqH0N92XclM15KmG3cezEbFoWo+jKFdI9CzJzcVdot04ICSh
psyK1BOLQ7QAiqn++HwtbXFN5gxCqQi5NkQVxy+Npm2dN+e4TBHZtYtKyfZXrcD+aCl8Jz6x6t6f
UT4iO0kutzFRi8KXoboQuDN5GX4ZHni6rvC2YX5BJPFb2pYtoAu/h1l0h62om1hQIUwFxFXCp+S6
JBmRTPNcf+4pExCP0QQcbtSF0f7gZOm6Z5q32+7FPVw39ovKtQHfgbMePdVIO5FE9c/9UQN5vQ/B
hcnJz5yLlsGSZxe+eeufqnPR0+GdUjgmzWOSWoX2NvSKobwtGE6FZ7AG2UI2lwDrT+8S//qdK/xw
Pzs/ZvpovVfrepGoZvSD6H6N/7MWRb+kWgSGWs/rKGzxzFFCxx19jf8zF/l24jxJ9OaizlDqhShe
s0MQm6/FUQPFH1fNT1/oEOtyOY2eQhk/eWs9xzeI0vB4OKTFFiyrNscozgqx5X7DaPQs/+cihJ/6
H4E3z6NHsG4iga2mjMOyhYMReUhwsGGmx6RCjBmP9jI84s4IGMObvYanwCtOABRG0I+K6sx4fsKZ
y/15gH3o5N+CgZ/FkXtjSX8nSS769+5wv52yxCog/sS65rKCSUoa6lcKc1nrpMHnVNzO2ePxfsSX
jsfV0JgvHaRZpZJ0pR8Gm/J78t6mDBdHeSzPoYmJZR4K7EZAdTyMuBqKl3INy0g0Qg3r3CsJEpRn
8ihWFMtZsldISddr+HoKqpz4CZeTtcXGq0ZUsKxluTtRLeToK3UI75cAimAmLbjvR92ddRkaoVtp
MjawF33raiF6wJhvVLdDJDs2WEVRgj//G75y7dZ3R39ixmZDL+k0yXYUoIeC1FZZrHMG+nr6vh3C
M9oqTg8MsWp0/4tjAzoCI4I0P/fV2ooPgKqD59jJkZCrCaX0yqXp9iJhYn0C3CN+g8V7eOE8IaEz
o0IZUG1GOKoGBT/WV+ILXkKl2xDoHYHYpu/TKaxTu2OcZf3VPRunR+PxQjl580gt/y2k3lpVrbb1
qRvjCtSdpl2v74hdWCw+B++K0JtwJtUSMkNd6uZw4wFEimhw3j2AKopdNb7NAUj93d/NsIEnuqcU
GB0NPufbrAo8r80+orK9phX+BK9iOHgR7gc7RGlQCeDMdfiLE1UxzD1wDYRijcGvrCQnGF7WIuOt
B0fvD5vOExQ175zF/TwF6QXikG9r7yIiwrS+hZFxM/EZn7t4UEEJ6vi5mJA4oxe6/hMCA3jfPV/I
uGMxUkBcExmsofYnkWYutXTwFgBRi6bgHikPvCuxfA/h7PGBolpcCF4Gm06U0E4CStzfe7Qfamhd
YY3lyXbDMQfHCk1V3K00eH7EREoqfK8D0cT/dZFsavAjBZnjlC5PO7sg8NQSJNJLDPsVCa4OXjI0
49b+eVBSZxSqmge5oczN8w+dWaM4QkJ4klht6SQzcBIGMeTH0etyb0qGR0vHVjua1ZEXjGv+fIf3
jtaaIEcc+WU1EjrMc7U6Oyr9kkdwtd3RtG08/Ci20eBOkTFk/CZMRDU4duIokYiK7A+aBJFhYOBu
aiaEpSVk/Yt47sF3uhUoBG8XjY+z7pROlw90ihK9icUJg0N+Zb6LdYE9Na2CvYY31xeox0ecd1HH
14GuUpbYlMdmwQ11SO4S49+lrFoyIcZkKcr6xACFFYiPzAafKfB6X0n+Crqb1CQWvSISCAzmDoBw
qKsxg2sdYYGGk9Fs+aedxpsYXLgQDsffEf3mT9uoac0AJe/QK+0Rsg7g503TGLeyGzKEfRl8zmes
26ROyBAzzLU4CuEWZ/lrM+sfjiCd1D8zq7auxYrNYWyWgs3rFIBn6ziMmhDL6LhZelijZ/iz/8x3
7d+RBpku04nh+Lgt5S3xVHCHnWuODkYVsIGOP6F1TndCdyyAncZxGwhSsz52XEVXKRX8Hhds76jN
Z+ZfoLvfhtr0Zo7j+su/2oJ/vrqy3pkHMphBVJpOs+3o+JWLp1n9gASmtzk2NSuwu5xpJfy4L0jD
ZSafJuzi1NIaoYS4YmJJS11T1njtv+F+u+SpA6CduKY3DmXAziRsRQt9VYESxFtiHvlDSaOEEg2u
GpGAfTMkWuocRJoMhCtsh5IYQnr+gdKePYqOppbKGOmhDF0k0A7CxWajhtajsuLMLOm5Fx/GqHhM
yPe5yzmtk2u2TrcjF6dbJIccO5tjYPjsS6eyJfd38MfprMclHz7xFTuU4TA4gktAtAatA78Paic0
5Y3LV1oQjnS8kodg2NVqHfwDg5n+lt7vkyoC/fZbDDvI1K9K82M5mHKV2Z7oyo/X6xEcFmNUQFnm
LEGCCi4ihvyVoH54wX97jg2wW1WpTQbZK49xFdshCMrB3jtvykQGXLEwDExdYh6kNOrT/zpL8pQq
Umsi1COYN3fgx3knSf013eqm/Ky/et6rmX45yCe8MAfoFBLIdeNJrhIjjgmh56rBLiA5CXNeo7lw
Z+NxY42N8AxtzwvhMpzQPWhgQwndufSDE1y/RBIEhAfCYws6uLmAV6A8VZ9TBnfDp8rt59aZxLFh
X8t9nP6w4svIwyskBYgOTvwQSZixfiBu64ZCQT/8bXciq1Fx87x/qXDcpveZ2CW8PoOZRs+bp9nm
k/Fo+8RBt8nRwDxRo1ZyoeyJpN6hSz3apesqSIIUm5qwIpyU99JPyHBZU1U7WZmuEt0hwmacHUZM
KF4PRnuD1EA66DsYyvK9aPjOp5jKDPsgHP1NnlYfBQ+alcR1rsroDM7GNu5qtqRjHJQYDSWnoVb3
UjjCBHkMoXP8+7WJlAZkjlSZL2GdgJprxPaqbbuOwJH+f1i5Y2g5hC7FC39CS2hcVS0wUBHqvSMd
vSFxFVcNgwdJZtZYsL0WifF08XPF+1U30XgI2pp4UHkAuJNpyfw2ZF5ncIvbwiarPfdVTLfAy5qy
1hsWgSn/YCt5YjXvgztuYP35blM9C1JYjTwj67NnMDqxmEIgb1ycnukkIpjG3I08sRBarvyKMLoz
csYgWlH8tRA4B7LqpGpXjlGCkSsx0AzfRORRcAOU43qYdQhd8jH8hbsERlcx/zuTnWv8HsHHFoKL
FIkTaCNCyXonpNQZuPren6RoSLbZFecomPZiheOPQTdgpxM21hQ5dMk9VoBUVcXPrxWj62yuXrE5
YUWMs+GdYME3zorZ0GYGalRKwpVklhJyeSAsCBGrrKnHDErtaEqYErsTFyXHQ/3ir6FYa1ogCYyS
iYVSYs8jTeOrwJ1c9Oi7/kkqd7Ga1JWcxT9nyCQD3L6pF5XvcCtbn7kN9HnqJxn1WmmXvia8JZ3C
EIETOHaLJ5Z+gyTIbswKk0/rQQ7I2eO4tRAVWuYhTV+5oPyeuFhYKd0Ic60mOSKHf1FZbULRVqZt
MbcxrpF9bGWl63u0XZOUTk4p96P68GPvDaZMLQjj81fwqJK30qY1FbI/JOA+2gkFJY9iQYS3TU52
vPIlwsL2HCJNsBm68D11cqqiSLgbVYCXf+IbNoJNEjCtg92VV7p/ZRVB5EJuNrkAhcsM4kp/dUhd
P3hMCNpV35/PkKqLBu+L36usvKJ4Mmnip3/SBX9QhmU4TdQYUOwuAf6ik8riKVoT4NGNTvdidroz
+4EN9ZHwHFlFRj0sc9xTTmQa8P/iQeN902EMHW5k7NmGj3ti+Q7JcFP3Ek/N19oJVkL7VG1GWau/
PEwcAAYqobR3S9xHIMnjGR54NzUI8nVK6kIwrg6dcFDg5xJQC5tdc70yFVYrV+xMuucP8W4xRyH6
0YvDrjDqoh22h8sqPvFu8ZbcXhnCC+IjYz+DMzwIY5w2TkAd4D5JoaTdlNZP+GiO1gAJVL6gBSAQ
k+Qxee3GvzwBVhdczNC0pHvNQZd8X/kFVR0rwWn4mg84bBezhso1aNP4PbSncCDZqLeVyfJmBuuv
h3WCg75cpDoC+QuA1ncg2sy1jgi0LMwYASYWzroLLMcCIFrpU1pEqItCC5ajqzGcnyXgpSgPn1eR
xUOuWnLBgNcLAYs24tjWDffZR4tV6A9T6A3oodZJ/4gMo1GgpcKPwEiuzX3fvbytVAON+mRQhsbR
fGsCEMVURj076uxRSfPwPQFOv1Oe1CTpBGt5xIF8Zdomie6fSVqEvdnZIk+Io5D/mH4KuZAMZ8uK
gGaeNDYq9Fg2vez2IVDz7a1AxLkBpeiQYEu/hijlbV8OsBpMfTac11atf7A5gun16qW22nE2hvgJ
de9aPTUHdQkP6d8DoTadQlXJgHI6+K9I2sdOnCLNydv12lbwZef8DiOHmsNEYUYxYa4GZJ+sDu9V
hzSGB7JIjHaOFjPa1x1cgNtw+z1QLksaG6meQ2Uvypz6LZp/zOcEQE3XsPCn89FqNBFaLPaiPaIX
27DFG7Dp1TYxLS0uX8rTU8uY63yYQ6ffBw8MyajF6sD7q468jz9ShkvU5JnadKrNZTyGMsXrHMC/
dfAiwjCJtZU4h0gkL4lWKe9kKjIiMmTcJ5694S1CBnTlwl81IlCHgDvmAZmP49Hufs7GmlFqYCZe
D+Qiq3nNlR/ZbbvdOW7RIOj28q5QjRlzzMOv1ZKNlGRD0SXOnRj86I7Yz1uQjZJirWYmcHLghiCs
VlQKiGE+oZFLz7qAubaHR9/fmW7T4wTuasDEOvxDf4LaAcaTt4AMABWLE6kY2pxjevz0zxashQhy
qwid612QuEiMNn06YkS3AZHZAYQHm60p7H+DCZzjnncBJYZc+BjwycBFTVJAS6jpI5oXTz/HhMAX
OlMh4/ynF4tSD6kTjDt8rSiOKKK7+laKhxtDMD0Axco9M+PTLh285DRj8YRj3+ny001plhDyAtTY
sDopDddwdt44qEC3f2Pq/Avu7Z90YACBFb4aICRHOitj2SXU92AxlTMJAFu6DFPraQypixycd8Da
tDAaglsNZJYSBw2f1XsWaMspDrfSIeK0GHYAPiB1fGtrjzRYG5yh+HJezwGUJy4PRCBEFQcLP06u
iSwVDqsY5Zb5Y1w5vlD/wXCxRnr64ak4N374sfqtoFKRi3OTSzaolcHNE/4XuLXvTaS7YMCeJFqG
fZYqZi5ldXHnvw28CoZDJGJkKiyjNSkCiMurBRc3jHb+oDHHDGEm9sTawq/wknb+ig5Lx7kGjKwn
gQ76j2Ozy/ft7hmPWee3iIHjz5idp9yIK0ZLBP97azeOfV2olvaYLeoYMXQK2dTYY7tfUiifHU3A
U1Hvv/moS/XQyh+rCXGibgxbfC0uCvVbqbjGNZPf88FuBMspL9pAxPb4MdrTTWoGXq9BiYcnhB5b
Wd8AgnOCZJuPAbyjuUFYnPm76V8RL177gSaz3sNwFbqYMFZLcjIPZeLMLyuH+qQI93hU8XjKy2fB
R/pPBx5LZ/65tr8PpcaDCnm/V6zyhk1bz195UVejdArzC8OSXFtHJaC+WHe5ZuAN+PrSsipQaNsD
tPF/txn4WU5Od7NIbTWQemOvXQ+ABQaVFc8J0fHLLO4gtNwLsZ+/ACvH6qyOsYkoTGfcb5Mbzwyc
rIpLNZuU6dWhStgy1sY432BRhZqCBInqEsU7sVgnhscB8yA4Jpb/B5nuEHt9QxgPwMCwNTHU8PFW
zZAOhltdbz4K3iaKEriXI5WkK6hF6SKOngYlTpctUEYmDgEOlKGm7JzFPWuELxjw+99u2atkvoIA
SONMchGtRqXyA+B3Asjhp0d3BfyWMtRgB4vewec8aRYKJlQLFHxs4e1CVHFxKiFJjSa1gDATsvRe
widxCTzqLRTt0JE8aB78d+9G4iFi1fzAnya5pxp8Oes2BTa8dVd/B6mzy5tItjIZ9/zCOQ3Zybkb
+F4tkzddjBOzwmp09SNnczpnc0re+Y+xY7Epw989lm32myBbzCbabyoOoZBCjb1U14PzMDt6Q8Xc
icdWqRF1s5fPnYScwbDRyWZSSumcM5jTmCzYS0uniFTIWeJQH7ajNw3vOjudv0HIcgAFVAQCJ39B
qcFYXnNDVNc0pL/JzDkElssqgrT8UeVMRkRFb13/HNaDErEUPcadOSP3JMiBqlaJ1wfZlJBEijWc
D2cse3+aLIn9Puw04+0jYMs3lLomGGdwG7nrCNjbqQ5vH5LQ2IHS22pj8rFFEJlSIMIX4Wetz6DB
2BLn2gcfhtCSbjjnC+WzgT7z8TGa6hYcRTcX6gKpq1dMyvM+or8js5rSlkhaSPC6n4TgshbDmYBy
R6/MvtLQo2LfZp87M3b9jdijsPcDI/W2/O458a4xJA5BgdQJ6iC+k+V6+bywkppt0ybzG4iQaiRO
wpUUo9TG619/t6RYfwRG7pW3c03OLeqoX0ZWs9RELamhcJCAAqcN9ByUOPiWzBpr8uZQrle8LnIK
hyuxkyKJdvx9kpnGSCU9NyAcgsRTwjrbIn+zgJ+/a7LK21/r4jxsmy+R52/F/4reqfOLw8g5e+Fp
U+vYVaIFMt3S1GMN2ByjHsvM3AVM7S/A0SzEHp76MX2+pM84r1Knzbz/HN6rzzgACWq+QUODHYoD
cVwgk9k6l5wfF8Cix75OWQNiQb19Hq6NpyJSJhWO9poOJrKVw0cYoGrynFD7BrfNNvKoTqo15cXT
jlo0PMgN9NrTsAcwcTI8emgoTsCVVK6yZVlS95r5j8UcjCgLrLFCeZajvgx1ZXfF9IGzHO0Ebre3
4snbjtVntGrpnNXfaRmab4bBmrvo3adNlGCa7P23vS7/b8tjYBgXkizSYnww71hLloaPVzfVKWhu
IcaGPdkcZKFWmf8ll66AUDRg52CU3Bbf1joQ6cYhsHTRQhDKLixZadbR/+s5KroCvd54cx95OXSj
fXAkX/PwHT01dBTXLdKAn0OCf7r2m6RnA+wKWtDOuNRnHB4cwvvVPs+mp/5HbFMB4ybLFO6l/bXl
i0kYhUrHnA244D/GAq2zOGEFo4Gzflsi9q0Xj785RlzKZHLrPu1ILBODcHaEUBWeAO6ELIZhUZ3r
5KzyDE3x/hV+I4N6FxI2R5KBwYbJ5RhdlwAe1BglhCVGYZCG4d55RW6yEnvk5tUa1zdqAN/s5jMq
TyzQuEXBJXvl16FTSC9dFRkKgelgJU+7k6vC2cxfrsXTVz3hHPcfTC1A2N94AzdBSbo3Gt11cwt/
/+FVUo+F91MjhSuS69AXwIWzjmEOxtqpVXsf/T9XVFFg7ZNsMNiZGPwvNvxX+QZZgVRTtqh6gjYm
rYKtV5DtyBd2GKQ/u0Gv6ZTR/lSVB4b1gDR10SI4+VvHpZ+qsIgOmgrBdtjuNNi9cki1T6WoI6ZM
weSG2ry4lRvyFH9bYJYvE4toWF5KxyDIMWhXRWKW9os1N0h+op7YA8SJChe0XdDi1CnuCsAdFYvF
7+viyWvROOoNkbbVYX1hbDVvsQCYNzP2qdsQXcKTfYpXh/DJ+ymLRFheWLkbCfHU+htMTL9A3Ebq
Z8w3/3eSyDTm7f1Tdob7nsuoG4PzVrBcOINimC7lq8Q5uQYnlXuD+VlZZ/r362H8Amo78TRrEiIw
nzthsiInyyYkm8i98LTxpAnrzwm9xsfxTLvAVcxJKCzxHbTh59z0PfnI0YXd/aH2fN7/rkpwlOp8
t82u/c5U3yYeywLyJzkTzrWXOP//Hwl9ebPgXRKISNkJaraojZqF+v8O6fVj3TCSzL+LR+tNK+cf
26Rjwi7mBBmrcWgq04uxoNqdcGXO9usduAYYThdNgJK+mlieVLAUpJud28zthbwhSlosItm/Rvv9
MQO3hUTe9YYGaKfEcf1oKpn+QwabeiGEy2rt59wbKpLrfF9ERbpIvWhoD7t4e+LzxAZTB2Ir06Cp
LwsOfLsa77QhFQuJw5YTxPpABDTe5YROB99q0GJTmg18wh/YvXiZsIPdW0JORt7cw4LC6cabJwM3
AfcooEjGQpXM4PDcutxUQMWqsrqgOuHnyTWp7r48XLLJqq20Q73XJM9U+TX5DzGYeMa7Jq/idByu
+o4+ERJB3ywOpGEhP5Kh2bw3BKbeb3KAl1x6DzQ5Lj/sIWOrTF6t1a0OB21LB0pPPzD9fIH8zPE/
ItorM8fc2y71yOsmt1PTN3L8WEO/ko/IeTiIfys+o1VJDdpP61qwoVKIA4T8rflA0ECZOQSJijD/
GAkJ8RH0NOxZiCGQC1ufnLQ0DixsAF6DTTRZDHopk/ETw79wsIkD9GcDa7P17Usr4ChPUw04J0+j
o+LsJ6zCcGp0sY0sizpd0oBuB2vEtZsJEDSJmO0qP5u9EsU7DrmDkTis4EV70MZDlon8ooAXxe/J
tJ1Pn6HXmgt2SjfGzRe7NjLHVzx4XoS4+3izXczf/cJKckRmxrN0AxtXykhFAcqd7ZWAlQmRwF24
IZ9MYmuwKQcjEZZnXVkaYUi/4Fip2HU8kNOLbXRC9EMMF1q+z9JRPDcUrPs3l04kmt/hn9cF/g48
b7aeu6i8aVsILfllfosTVhnqnB89jB/kMe0AspCuXr10qYao4PFWMY3HpdNNDDxkB251oWoygbin
2HQ/OPEeyB5mifaTx5y3Ti4e/B0SfDe+yqbJiV4b7GWIxJu0g81rBQfiVORsd3EBscnyIsqJS/Cy
NDbaWk9I2XVEWfPAkngER4B7v8wAk+0QEi7arE8m1VjnIqaItpLyCe/H4u8Kmj3P1v2yoh3na72O
ys5555uKlmvZ5Cqyr6lKDCDtB/8B9tv7TtnZ8UP77nQZsCRJL8iGnyR615nfK2G6X6YKVFnjVKpG
GqlwPO+Z3b66rIaL0P+aKyhRTC7/Y68KAqY4VIbhfpb3RUi3WA5p0pMruBgtsqsAHApE10iQZqbJ
aOKb3zgZgebyIDQwjCKOe4N/+8d6iEh1PydmLqhDTTL7sSfNx3hwutVgOJgpVyypYcicqEErkb0U
6F6OB0jNrGOJy+XJLF5b4rmIhsMqVDmgYLums3MitMVy7k0aRKWzuX0ojaublHFTbEckyBQdTTC7
HseF/1QJiaIzIrHNsaJ18S0pxVcHKfrRnZnIn9AzWkCSHnyFfVmL96QYFgodKGNCY4We/FqfR9IO
PiCHxvROJDSNtq7c5aIRewTF/S60t5Ho9CNLqsFYdPhnSvhG/nBCXrobD2+zvk4ql5v5Mp4QlN2d
Rwd4wAxrvMiHoElYW5AiWFzs4n88tgZm9J2zx+qmp7T6+nLX4S0bU3ALbElmdQdbem7yYc4zfXY8
bpBZ8Buoohi0zwgiefdBE47wezOszoSBRUv+S6u+KT/peldURcXs2qs7cNr3mNHH2UD500pRSq05
qmtz8OpFFnRKSvZa44jp2e8hp2FHutgUBZeO3woePmbibPdNvrfEFctOY1hdVUzScfl9KrjfSfGS
8M78gQk2ZTOHTTeXscs+gNGpEXv9eVMLpKA4UokJQTMNd8njJKk6EMd7OtUtLZR0quycujzWB6n0
ayDfz/enQnbSyHzdHyD9GSdabuIjfa3Ce3i72fwXNj3y4VWmAucziMgLcqJZ7vvHj+Smy/vao8jC
d3bH1SpChzkQQLbFHipUa03Piwf5LOz4UqgUZSU/ujuB5EP89Q8SIHcdyIPLZmeyy2fS8oobK22X
A/c4FZyYjfXz6RrlSZlOqzeJur5at3ku55XOE4GKmeFkx8ug2/wg1jcaSAOlpwPyIOEbkEXH/uU9
RQ1ad2ZJbhE+n3NbonGo/Via9Tys46jF3yHjAwpYk4uaXqY5UohNHQnymoOhR9oTyYKxmYbwx6MC
a5sDuJoXA9CKt5c0v9SUm7i3qIphNt1p4Op0v20ALp7Ei7/iWJp4hAJ3C6aUsO3MdDZr3iVAMDwc
wW6T4eGz0AyLHWGHuDzo52eiaXBNTaQx0ydoAyKQ2zgXBQfLRVLY3/ut8pIQS2H61XsBYKBIG5C7
Do3coXjururgdaAB8O4oo7PAH4t8pECtAP/rxLGhLKzkewEyPEVyKOhUB4g+Ww4rWMT1o9vNJ4vJ
lgU7htzG12FJbdheuClzckc2UXp/3ibY5iG4BYy88LgliJI6TlvWTZtmWNMYMVSI5jE46K94OsJZ
y6fdcpYQcvPB2CtYt97FdVrO6imMZtcfB+dqhAXOM+I2NmNZBtSg/Q4+Pe8paQfJX2iyk5s70p9a
7k+ZmkN66kTYz18lZ4/EC45RfUsy+nKRE8kr+s5hthkWP49gf0EUM4nLDhPOn1Tqj6kIha5jBerP
Lu2zJvgRoSbHj6UGf1eazTcPembJmP0wHI07y5f4gMUHoREMW0Vr4q4sjM2wRKvuiN37SmijXFFJ
TsQ48iAKlgwfHIhJCa4xdg6hsZtrHgfrrmXNjZRJ5YlhkTiTfed1kTd0Fxsy5sh/BwaNDpsdKpj7
2dH0etQ3RRe1H4J8u6ceCyL5UJtrns48eKTTQ0WNymhO3/eiNiDl5XMehd9+xfrSwvwZgL5x1jaV
pNVKVkb+56+MuDP1stvukwKG25nIxtC7dQH2+ngOLakTSrijm58leWwZHmbcLXSuBNwmL4Nv5XCW
zMilFLVL8jO8C/TBrv8gyfwh+BgtLMQ33zIHPgbsBOGEyny3/q90uGNjoOVK0jDUEeSDlfg3cjDl
cN/O3vAILrDeBAFZd6X8Cw5RMQ0NS1LBgX8S9f3I/Li2E8/JdYgLOL/3mNPivkvuCDkbW7xcsF/i
cKbSBvepkZqYZaSXoPjt5ugXjktmaQrL6A1AIVhXhx64f7FBq9cEBKF+Vk2IYTYPPZqg/EaqI9mG
uYrdqQn7FDzlh54i/RHlfzxtAtirMWRA2SVxk5jKKL2V+Mg9p9GhizZyA4HeIQ7uxfwXWehpLCB+
Qa55YeDk3eFQ8zv2lRDFhhSaFFJ+77EWPaHotpoI/QT+0Nr9UGWMOq+b/LruVSFqGhJh1vwGSrLL
jDA6kQ3Irl4TERJz+yHfZnZxBlV/iFDiYuMh7wyv5iK8Gb+h7X8ZDLwOxEU9JS4sDdmnNQEjv2cK
DrNS8y//8PNCsptFDED3Rkp3RCKlEzRJLJttuTTy8K2s0gxsGVGV+OaL6N2mw6hd4LfGHx/430+/
mhZenI536UzmOEXnhoXroS+vNUCUNjr4GX926iPqMnnZWyxMCk4eaQJK+nkdWzRRpW8yT+/LEQJ8
u3AIBhcRl5V9eCBBr7B5Mhuk97h1EJMuOUIjgde831z4wYfxLT1WEbjU9xSnetrtbwYlNKu96KJ/
ujRZki8n42a0tC6n8sOtEX739074gbhqvnNFqmQMCF+JSQFvEzMrx7DLh1H4KdKt5qoN2y9nFd6z
4NNE2Mz0jizQf0bx8KQvhFudPitYSzytlCW9dWWh1jjDJlTJAH6xqgyk2+RaHH6deHxEfzpGNgAF
NGzAa80GoVgb7EFEGTkp4/U5SMqC/h+qz1uknzKeIJ4II9Hkez9qDYJlXTP7PJa+lZ2vae9QKJyo
V4Hx2lsNO+bDmNpXWmrLtjdgheDTCm7fof6HBGCbjRmKv96QQda7IQp1uTHq/V75EBQCI2E7qnfU
eWBmUiPzGtTm92HM/faObzy27wHtKXttgrnjjIm6LT8MjnWgEEp8UZ30WYVzHZvaEHhGTOvrxNhC
6bw23KAXvxeHTNwzhS0yXS3aDe4yNdUuTv5KDpb5w2OIXWpTXRfrYjDfa3Bbl902spbTweTqSshr
E2xw34Jo1n77ap01Nxn6pst9u8Uf0mZtXS2hWJxmgJMtKXgzs+dVY1zJS9sEiqB4npJnSqO5T90s
bSK6DihyYjHFmK4LTREwGa/1ZkvoW3TrBVGzEMiq0jGEzTPL/B9mdP9pyH2aLKXq+ua7UaAJfq9I
gainJZZvisDvP3ZVV5escInNKxVSjSs42NH3bum61qA1FFmecWFN2rV8yZfG/gwGDZODDPU9QusG
7Cqa75GybUmPXkVs52u3GWJN6++/TECdNfwVT3YrSdNqUSUZOLYs6TFE3vSpA8eugTaa2ZuDrBaX
l3gPiEk3D4y31st9YU3jO8Ip1oC84NAQW+vysCA0TiRdhDBEsI82uwu2jWs+I3lEYK8IE7K/+u2P
fugbO4pOfr3HGVih9v5HdQ0dT2TWWHKRwjK1ZmjP98cUTvcVEAWTYxop9N7jKKSklO9wEOjYsIPj
HpZ5pO8J3xqN28PEAYGToMdYs4GkNOpinAdTqsSNWCb2TVRFWDE73x+EyF+vyA17ZytATrxKG10h
3vdd0yYJykbpQBUwJ4CrLbajIOe/q98zcI7y+ODUf4/u+jfUE73MFHugnJ5FthFt7wkeX7S6zhGt
l5sBMSyPrPgoiUiydIq3XB/eJ6IckxiGWEl6OwLpumrBCJ2lb7Q8Zw5rOzVEFffahPat4gT8t8t4
LaBW56gzfbbEyl3RvwR/badKEGSBbEusp2eEGbXcv9DcnsQp46y5ICet8Nw5lEK9cjnBetbj8c05
0krqF4gMM+3e5fR3B71Zb4HTrx2IKgsW0fhTIbwabkIqZIYbA7lyVBX3qh7tN5gqQReH+q4QsueB
8tiaz5jFKmILV5I+cl7B9gIh0wTydJa3tUKHiER/B+G4NMP7el7+9vSVIjK5EtwkJcn4PvgqlcxP
3YJEqV+uqRsEWFdNVgmdOeBLTK6cQWjJYvIdpddZz/N8155GVF9l9lmRvk1nmc10JOVEig36tjs9
O7dLijxza4lKEFQ1PXhhuEMnAYtxCUMbIExOLd4YiCUlB1l8fCAXw7pyQKo6C0pf0Th+hDorqwyg
xdLF/oovunctMcY29slQCfjGIWjm4v+wDL60iqRcoZqJAQiQfQdTVeS9BBTU4LOng5xQnHvz+Se2
PgYLQ+SqPEE17dllGxNNHUD0hQshJ6AV+HrHWpFKPW1S+8hhXNo/Y+MfE8RlEAT+3vJjWulhx7RR
68eGKpdYOLXs2Vor7eONN+aijoKLOFFrTu6CPMgjzhtFgRZ4fGM9k9HmxKaB/TshS0jhmS0BmdPn
O5aq7Mlfpu2NN6k5Q5RpGB/p/zzS8O0lTjf9dAiV3vH+0MNhA7NKk1NgJNgIxPcVaZiRw4eDhjfH
5s6OZsnWejxHt2wOvgUxie+iGKvlffyKpcKkWovxHZwol1DOaYFUpU+K88PMik9v/OWvIEK2cRv1
iV1lJ9UffJ9gIPAVbCBA2ls3Hmd+QEYmNwqJ3TDJ4uq//EEFv4wCd2wPw4TN1jzQVXnVrguB4OMY
pZtoK4v1SNPQo4zPgKKWlkpCoZWfMD/wpGcxwgJ2NoIekMrvqnTqLcM1Q0KIuOmEJ4ZOD24uC68P
60mC7ufa9rgZ010AEDVok9HqQsff8XVlFVj/wFUqt2tzf8nVYFYDXFgaRM5j65pX1Xi9EhCZ3GyF
HUqL9BitL2+1fUmCpVEonuJonJlmaMurpaWcYoYrGwlniWAdFREx5qlYZbYAKo1Ld2mz2hgvuDVP
gYGsOdifXTTFnKKOxXBk9uiWJkxbzz3X2Ec7PGQMqelhNeBWbz4QcMxY00V3OrvqL9vK9qdHmXn6
PF+kah8h/nyHH78dLeIdCAlagaMMKwZURFwyrLC3PdBpe5pcQo8gjtQjRoAp7yCuvQmVb1d9Yj/m
nEMncQUt3ohomiJHIx8WCmKHfAGqeSMioHczWiNgaXVPR3yNJ+bJx/2fBLY0HkxO4/sooX2Ll43Z
24EfvDVbHh4/nxd+XubQ5Lw7WawxSf2Mkg2zXCJhCSCUcH7li55n5DuvTdVonOPmCBw/vC1jc5ZR
hQgxcvVDj7ALteHM3sC+XHQyMGwlVEZn/cj/OXCJBa6sT30OqKEGaN+FyrHU6Kxv8r+UAUHHsDoU
KvJFBoAbNuMTySkQNhUuvmiQ4x/aAi3/r7xQ+DQJjx06BCxLgjNmgUtb1F2gmcOzeqq9Y+iiKuX8
yhvF+HpG/cqJE2/OlUaKpf+U1/NNKnJuhUUiQ0PLpyk3DuHKc6f2JHSNFqkbuKPHug2GGl4z/Th9
tjC4xKJKdA/wVQa4GCU2Pb1la0XJBARwNbUCn2WCA024N1DCc9frIC/sWLhs1yC41sCj7IC/neMU
aDNPRUIsLQVaEpj1qqBzRx4IdT3uK1NierDfJimAeSZHSklnWlnLSCvAEyFJq62hRyw+O03uTwSO
/KWmsBLldWiBhNrozPQl6QAgZIxjDuB/W2ccVhmGcnbgaFIkmUKUAKqTWUz9ibVqwalz8VXL1rMU
g4U2rXn7zDhMkOWGOJRbu0GiJj4Wm2NJ7XulE8aQufcZVEBEQG34E/xpQapngRqVO2et4mu5Oyo6
1gGm/d0tEF7LZnLkE2Zu2KdiSzfPRlHhCnkvcyfjCDZjaELMK6pK/675TVF2qTJEG4pwfrKGrjsR
E+qjWULGJq8CjNRd8l60vUtaW9Z5IZxSh5DSS/6ZqDXs5dfmpu+cYQDRBzySyuvE9KgGZ50S42A6
3awEmRiL6bY9Ner7aGh21d3M2AYhSpj9sd1GF7/JuYvLhZfDH7YZaNbxUrPWuS7+tcu5GAnML8r9
FSTsrfhdLF/dqygabs5L9pDvSUFnxpX0Uf4E2zOUcA++wZv6Yr8OC/KDt6fR8gTIaL4sG6shVN+Z
SbO++yJ7UbR2LJ+ySWzHZiwilUJM+qkU/FnwPfVVZAiucdyZGSXnwW3LFjn5F275wGl0TnRws8IL
RLp51dBmjW0OjrHA0Dh3IfkQoteEFf+VNauIlyrJ8ucXHeBlW9YcJ6B05B3EyOLJ09n5kiIAW7Dk
O86w1CdBbboVQFfYfzMr3w8nTesSYLzJ9WK5kbNUyfCG8tVKKDtJcIKgKeznrLY9Gf8Ao1VnLBFa
t7VB0rQF3E7SnBsSOWA81kFW6Afo6L3XaK/i7rFghebBbud25IowCFGBVlN8OlB0TMhaJi+GZlfF
SzfK6SfZA6Jr7QW3xcJfBi4s1RaISSaVSHI5qMOiwVBCcYHiZ3DheFGyc93dRdlLaGtYfrMx7W45
fULSzfRgshp9S4i0hnvOjBIMknnzxjkp8zen501XPgVrX1adYTbT7Fi4D1WCn52CPwAXoCyt1O36
FcW87U4JERmKgtLo+lGr+poVTVWietTn6/m5zinV8DjZvYfbXj1zlN0F53xQpL3jsXY26PWhTveu
U3pfTxaAf/Qt9EEKbUWFr3c0GyXjD23AbznmQcI6OJiw9IVFFnx+v0DPkheXTdHxzhgIJhnU5WBb
zfK6Jckdr1uXzfhgirQ9JtbuMR5Jhng8hdCbkJWwasRD2Up0UrxBIjqFkRC1QuS90zOjygGxumVv
/+3UVNR7om2wBUc+SY94paadNlvn6J3r3MrCB4WHIXXrwaRXCWT8D9UX4rps0X6D/oXBySY6Xy/8
IFT94+sKoPq5Ju8a7Jih3JBWYrxl2qQurXVSEbT/JBV45Lr0Y0H2epw9U/7FSddSLPIIdEmK50a1
GCk54c8c6YNyeoJ0LXJvQmF9t+A8Vic9oZbuIi3r93psaFAzmcBJd2HaGtkoW/Qz+eVDdujab7xI
b6aN8SNNhjY7Sf6me3SuMCBW9UppM2TqEBWuZfAYvyd/Q4oLTsiGj0yUBEIXB/GXRFTI5Qn+UcN2
vqLUR4W5skdXpdUcnwt0BGRSBvgyUcIbZAoCpGgCPb4U0ei3MK9IBJZJInL2Lb5p1MYLpQUSAy6b
ST94xJTCvxjK2FKAZ2fa7RktOZLihrn+xhnJs0SRlKSy5WEpaLWYHRrTcEo/V07gcKoxVqsr/HBH
/Mv7I3+G22+IZ3wDr19RUdUkx0JLZSLoL0rI9r5X08h1v8sCOpTNl2hK4erONudQ+TsBPqqRgr4W
f5FPUjDTtaed41DSdXBHk1Lmr+Rss132gTC3LD943I7Y/nbxpwvo1O2VuzDyqJ5zADhVxAjHCZIt
PgEXRfM4cpo6WIOz3suY1bnlh/C0iHF6OTTaz29zet8q3eWBvM37G1N8hE1XwhVC0UoySz9n0gd8
7/IePUDlhpGkxtc50zmhj6nkY206+iEYd69G8xA4bvf3RIfQQM59LM3b6PhIROQ+s0K4q+IzQoII
d6uerkKxN3SsLa6HYL2lF2db0GCIc2ZrKutfR012AdkKg3oeCEc0V0IKA5GgbeUzmP/s6JqKXGJi
Vglsq31YNSOL6+2kWdwXUY1o3pFWpRGcGw8Wqrzcv8rO3nm6UaPm8b+XtSXH4FZzyME+fnBsO9AT
/o2wCZnP7MFN8d3Yo/DH3RoI+bgdgdmIg0SbM3n5cA4oLsf5Ln84E9SRZ+DaV2D4cMi7eFNgGPlB
w0t/4rEVdUehItRxmP917vKHdE5PwlOLHcnx2o+RDebebhg+RokZBrpqLszFnjVk2U3F0E9dPYb/
GcBWcGd3dQYjta/ch+BHbfFoDG3HZS/R3f++4j/i3m0fWlDFZcnBNZOkMdOLSkiNQCFXxvr9H0/O
tpGU3qb0PhfCLcDLBCzK6DfwGc9U9e3DunOpnIvmF/P3Clfg5LGhY2OBeF8th37x/kjx60FucTgg
gn5JQl3RJxKydO/Qjk4gtbJ10Yyd8GWcDpbZmn9Vm0AF0izgcGb2mRuUWozwbWig0pcS7v7C5BBo
RldC/TIEspyfXULjg+e5ThwBvNroHcV72uW0lYMAcZRvaWo2yffd7yLYm8429DOcdgVi0hVCHGPv
P20e9UDPUqhDVaVxDYXtk9afNzx7myA2XL3/FAr2+LUF4YrNHt9SnZkzwA0CG9/Kal7Odc6ZgqIn
lnXkb/mSLwL9xD13OEdd3ceYsb6zJg+CBm3HPN8+vNIruigRZtgJ+ZX4HMP21M2k6AQsJoV6l3mv
cPPOXwhu++RrbWu8wS8jcX6u0cOq0lQjNgEz53Vvsmjd2syMfsecX98Iiph4dz02dpHOTbZnF1nj
3ttaDprYT+7b/vSSrXel/QC+ri98omfdRkVGB1RsWkjgrIWa6yKheEMGDhu0gkAStH6ZhuIOzPwN
gUWovJK+O6UhKW55qoGtY+oSz0oEMDIR7fytHqEkFWW2QmhWQWczFkMeXnLkG0YHwn6tH1if6oe6
J0L4n1GYwd/ZGPI6THiBHFP8gd33talWKeCZ8o89rVfjLRAQ/IF8nia8IV6wyxgzpwDdZeP3ocGr
bLoDXz+Ig71SeQACBP7cAOPHh22A1I+qsHFlZNPyqfoTq35BOYSBoKIzxch53eFN1gdlbwZJjcrW
DnQIV3f8ho4FuBIiWyOo7+fC74IDrMo8EWFWWCZL8DLlrN1XDXWi7XUBKvDN9ic6ampUYn1T1HyB
po6Dnx3HveOu+10SIybCk6e1JnmH8DwMu5lph/ug/xPQQxgqwuSgK6JH444rOdZJtg3cE5+T780A
/irjURkmLXvDfPSrRUMQZqXQ+LuznM0Ti0eHDEuk5+lfeXFbYqAS1zPmTdHOJ3tx7WOlhSrGSmvO
qWsj3kEdbpW37Pe8phjfIeca0MJEgjSwAe3zjri73A3stBTI+PJlyy8ZBU7Y1yc5rRntZHcmzoAv
4mrSObxY/4XOdhktAOjH/RsL2T+xnRtROyJ0OQcmtrPfFv3dUg+Bq2NY91Zab7Y7ISNYFPsn2q9P
pkuICkJCf0h2VIwidcUAXBVmG05QzQNZnE6Yud4VB6gljV6l7taKRqxxOrGEApJm/RNyxlEF7WYp
ibFm9938Zwi6vcSHZnlMGBLKx/HV32sfihK4VQYvzc8A/t00rVzr6fG1nxbIvcyzmqEgUknp3bkR
60O2PvcDhmynyEIHd+h1QMYEN1ua6jRilIMWIoGROv1Ps6+GE9EbCZvJmuXiHY2VRE5rJcaPKGkm
onszstb5cfq6247FVy9IIa9ThbJ+ognA//1ZJ9ykC8wrucLQUy84W85j+d5jxirrMy4OUFEOe/lH
rfSAlvXufV8/pitdHRSurRVRS5pB/2bWnrsi9Qo/hZ4fuCoUwGWKILzTkpJ31cdzIHfWgGSRALtp
Kj2lv50H7o2rB6dWl85wFOI3DsIBiGfh0g1myGn9dAqPBU0qIdZmyuKkGsSrncrVh+yWAegWpsXj
/3pcm8XZ/MpdM47njIM2JWjWo/PhY04APxzQOMuZ/A7t8TGLUK3zcLSycOkXtNNqEHwzuoE9YJCA
myls0Cm9/hpNFDo41YwvZKOxGrTbcfuVG0ewhBnE/enc+/7aSJpuh/GO0qKlNlbY2wHW02Hw5Lht
gkUNY/3J6hosiJRR8JbSXGbKRjrlzqZu7W2flb1J/63kuoxtZWkzcIiJd94E00p8c4K3JEdpucHf
UqoJ1fX7SM+j3QdVvPDrSU1AeavQlfIwdZo0KMwVuTq0VJpus25RTm3X3YgOM6Y3lVuC8imLGQgL
2D+EsMseLnpOTYreOHyKQdxHT9CwIKlGOUPzxXvSecbdcwaWAF9y0QpxnSSZMPR5kE7zVxUL569/
GRELdoqGNDMpJbqyIaq54hzJK7gjYULlPRxWO8WpmHi3OLdzqA6QqkuE73Ks2E7a/fPansYM6k6b
bLmPGAGTGaj3wcTslnm9xOaAgWkQSE9a3WtRbNUeJHYSa7UUE3MkVns3Mr0Xxr2okSeSmIDLxIp4
kDK0G9OkXbaWhFHRX1/I6TVE1ITbKw27nEABWypoFA2eG8IATPUERbRU/U9VmXehxNrBuQjwWNQm
7w3rrpYyQx0CavHKs10Ss/DKzw5t+IETkblcbAAqnTW4+BiKJiFDXKp4+Q1E4HOyyQ5J6H8Km2dK
yKmsex9aQ3p25Vdi0hXWSP0Ly+bRX9/i6vfNmAMxiX19ohde3eDRJjdJLj9kUfT38RSxi2cd50wX
FvknLQ7sJRQlnc0I7/nzDR9jcYzvJ5z57yfzzXXU2GWKWGW9WN44hP0mMbCdOXH28IxVZBvbBRLf
jt3UHwnwKamtkYFjvhGj+PeiDMDKU1ldrSaeoeLlG0+5kuXWjw9NV4UClnOS+2fLf7f0QDiTNJLf
7vIjAyDXceQBKTGTjy8lWpPn+rfWrrF970RnIE8zEFLAILSX0394Zo1P4wAZuHSJWjEOV57WMJsd
eGwYJ/ZDHdIzf/mtxc51ws+wnIRj+wC0PuwfvRHVue+cS46Rq1tIecBipunSAwke8Kzbn61+AE6R
SZBINtjHJvH8d1hpOtnadeDJEdubFKV9Tr9jW1jVhGyTUHDE2JCriWXAQvx4rvOeLsPcHPze2EzJ
hqzS7cKEjbYkDl249SonqjTvcNZ0o04C2qZAw60YBLJZoZiC5szwVUW8kNWYNnB2JQMqUDO8wYvl
FgyyGP4AT+ZE7wEzXdmq+TiwWwAxACl9IfWB6N1Gk0SeqRub8QJ83UiIaOPxtGZ4fQqsiHSaqvXt
LAUN+qRRZ0jjkcgxMwGrkqAjfHyxw0edS3h/8TpjsmFCx91/DqGwJXRxeI9WmOOBaT/fVaOhHnDg
c6nuqwr6a5F5NWaeRYntneOSfuxZJVBqFyNzAGgjWo4mv4jgV0SwqZ2qtw2PqVBVdj3neDDLK1EL
S+I1V/ct2jffytvmAfYM0veKRBeXUoN2ZaC7BFCRVgFG5RxGHq/EvRYFHbdrRUgf1zcnrXnwy1r6
rQ0DuWcAlmXHHz6WH44IvFy4VUCqFv2tUgiiLgExVrEpjph/htOaeoQJDfvFwc4wfF/Z0HG4ccer
jhwSK6/7emRl8dwKGPosRpNkQXQ4zZPji/herLzCrGD8qNsKGJrgnDxyNAS2LXC9+Pdu1kj+f+Sa
FX/pYoCZRBBqwKd7JhpvGla/5Nb5Z/2NkX2M2jDqPP+omTtdf/7uX1qoDqYs2rorH0mGeWBF8/9v
J/nLJQzIqx/dqWSBEaKVT60KgmJdRWmPsInx7BQgNj1Z2U3hAiOgIdxG4GFk+Y5Av9+iC/gy1HNu
PmeMS8xTj0dQ1KCxuNdA2qvwJgoaxo5KX6jJcwk7u5ab3OpvvhUWqXDx4iPGmSD62uFLtaCnMcVK
TqVBrqHWkpF39jCatDnUphXWRtG8xYZzZDJLsVeLBY98CZSm3W9F1VU84z1B7YRonjrJM9TJ8wef
bHWE01dNMcEydxA86sbrFKAvrygKhmSgoYUdik7tNerv1mavb1s6FZGSZ7wYek+mtyG4gucDibvH
5eLmH05aqxcvPLEXoigB7FdNPdszFsjG4cZKclxRIPzUwAuLzD/SBeVFXBe09Im1gibehIM3Dr1z
XOvuk8bvQw0npjuVKXKgDS/ZI1wbgVNfLl6UxP+FfKojDJt6/bvVfWWojDFxa/ElaLnYCzneuECf
dDY7h+pRRr9XMkm4GGocclGNnOJjuNoji42foyvBHR6tqaJdYd60EH88wXlCcDN0ENps5rRvBSZk
LRv2Za0mvmkyNlTlFPv+WyhHfu1b8JbZIJu76hIH7Li/sB60g5sKXkvfnDkrOosEpx5O5T4Y1woU
BhNpUGH1Sgp8mkw4Soqi8zzsq/DjrbqH54yWOnSl1/BJtQrfq700VgQBcWkq+lCJpj7SPNpyHNmT
hE3aSxJPe79jToYPPpJbf8a2EmwfoyZISnlJ/5124O5vNQKE02frNQ42s6sbDTZB7+mPsHjbCsAs
WXH2nTcFNGRjPBIUZx6h4zAgYsahSgYPL8bW0LV2HOGirnSlJBRMPSj/aG345fYswIzS255q9U1m
sciwi01dP9SJLzZczfBm40QNckaVoi3syw+0rsPgM7CK6wXLRNdwaif2l/TjUeponb0rbsv96YOv
VuKCSnZdQcVYhGWw7aZeQU+zXu344nBPHvSV2RnZXOqIcNHs6FKtceCKRudO0oZozOYv8Enhq96d
q+QuMYAV1wRuf8uFkYn4MAMZ18pkZNBDHauUAJ6Z6ZZP/5+8vx5LlkZmlVK4HN7XZiNj17JMjK2c
FhqJw2pxzE4ZCRvOdQYKTkV6gj9ReZKDCX1Cbp1sufR0ChpYL28yjPV0Xwv01Pd6/fVQupZljjX3
xPHS8asLsZM94UaAVKwRWbS45w+juF/1/xBNaHXUM8dPSwC7ON+rq+91wK9ZqPM6CY7JrVarh4Nz
h4JnTQzEjV30RLl8RU6DT4QHs+mkHiwF3qZ2nhluFvTANt7ybHieiJrQL8xhJUpHqSmDgGocPh5D
goi7BXy2HHd/h3WXhWcHpayidusucR9hDjooSAuYaZzo4NZvWISRXbkbjBjAWrG0DwREfzuNtNnC
x19i5tIbVgt2gF19Baw0AgAT8kJQVzC3MJGE0mwou5NaU7XRD4ailV4x4xNkUlPbUT8Y2ZCBgn0Z
ndVWCyFYxgnkzHGIDyZzJ2HtExpdmfPfgMO2FomXOG1ZKCYodGWBZd8P7SMReisZTIBLuL6r4wFE
r8uIKPeLDWi3Zq8tWrxCQIn2oPhCGUtsTbaac6JyH6ToiAFo6jO6q2XHtZDlvPiYB4lKH+gY7b5j
k8L5cUtSmoyscog8CP7sQHJQN2sSa/7WZtx1fOsKcIqwJYijp9Q6maPQFb4D0LTOzXaCI5Q1mu3w
Ea+oExy00yaTQzpb//nFFtcL6wcTex1ntIcPLpjDRmLvmn0BCMQaTLZhVndJ/Ju4TI9McrzOXLjp
9hFnaW8zWcx508a3qQ6IHx9SVGPrmocWY8tHl2C4V2Lg8mafZ69wFJ1kkKVrCW9lMZZszZ5BwgxJ
eKHAPNUdo2Q8puIEmHuZPw8vijfIjYcxkOIJzCMWqhKPbc6ipqU9+14+wpE2Z74EtEktyf/qx6Uw
3qV1VfDIbMaVI1TB+fhwV0UQRNAXCJVj+xWj3wjODqlXJHcWrkYqz42Iihcc2Iz4mcidQr3jKcs3
em/PH0QHvmzGxsn0bzlfaWW7i9jffBNg6xNr7Iu7Vklp82jC4lZm0q7A7ZmuHf5XqmhcD4jSWBI9
M2im9pM9xIJE+3UiZsYDjeebuWFxngCv0lcDN6Oa/8xQamyrmm0Ml+D/LBXu25/deGUgvTzcFUzh
RpYHHpE4KgrZT/22abM5Jldg3dqhSW/dAxypjIHO4qqJmhIMh2J8v78iI9xkBafcCfT5oCcNmhX2
G4U8wnKD9hxhMPMFF/EhmupiHmIg2ArG11Zz19WbKx1fwUyeAfEtzalDvQJ4425HOmpC4SfGdJUd
Ha8dVANSJcswzl3tg8l2vTRP4Kl5gPkP+YerZMB8h9GyAyesNtgj+Lz94S/S1MyFcYYtxgClBpL6
d5QHetPMK4nJhzCSq5hMKUBtRqh3XqN4X+XRU91wLfBOxaxG84e424GUaZ/OqDB+NFiyGIfnR4lr
64c7zJpR6PFe15QgxYMY4vtIgE/x7SUQF/3nqEjsx95Ni7wBer3DFpXYpK3ZhVl69NJLSGxV6hhT
sew4e5HJcatol8WwMrZHq/PNuqayFYq1Hvrvi8vOXqFzTCOjonrhI2vD8tBd+XvA4tuPED6V9R+W
dhk0AHRtddGwONi6ZkrlhK+HN9wW5EBOejwi5o4lgm+MhvPTCmGOBYTCeKnMhAELP/I0SUCxT7wn
Cg/3MUpdZtYzbpgBpE75A/zWKJ+68oRS8cNmUCnOkkE40X0bXMFEOkS/xWj660zzAUKiF0aG4NGO
dAVG/J87q379yEwQCCyJhCXmQ+16eAZDySN3zSKXfz/0zRW5IjTEnOhAVawy71cv0dowpDWh/mQF
jOWCUMCxXOIvq1pW0j+1axXHl+oR5oS7rjZBplJHo7BW90L55YjwQVdXpbizrj2lC/yugGZoZ4fw
+2UVB/C0RGOIGyeLptQZwO0q4GtOiBwbiS1Dzfhys6g4MyyYK98JtbWJ5vQSz6d8JG0OtE/SQrvD
9tV3Qyg8eACTMpjMVZNOqrSbckkLP+k8Z6iSQKf+VkaRtizTmj0Z3X59BOHfq3gNjzqehYo87eFB
1xMoQuiuTheygYJjOoHqpnNaN8yx07s8ULDCVqq4iAtN69H3sLw/d8n5ckFfEsJ7mqrC6vX1ojwv
rmW2G7n3ggO0F5dgT2SS8grXfrtXoMkR5WkYcsABsBUWCp8GF952gdqgKplX7rSVObWYzQklT0Oh
pb+9rNZHyNw8kl7JR+bTV8TSXLMz7uxcJCFVcOiPrwLu5YgptDkz/GuWvRtUwyBBmyW1+gHqbF9n
nVPuF9DcE7/eOoJJSuAlvk7UznjSxbSN8QVYIsTCCfuWyfyEQjrITRZQWc9SHBCURgSiMlQWqdC8
x7MMzMjTZ7YJXm0cgxNfNEITe429RKs7Hbig31OQOvrleYMlPO8B1ppXsqC57Jr3vfX7lE8InYHS
3skGEiKq4J5YXpTkLzem9qyeLIO6ihuKNNU8cs0K7v0C6H6KFOGBG/BNMG3l7MNTkvr6u038hSmm
ecSU9DD0Z3cONmiMQAero5YdyPQG9Fz2xKnPuYczOP44p4kq8Pt2E1lB76WSRexNp1NpPxnL8AkC
/xwAaup2UBEnwAkNL7QBJ0YD6xG0oh742lr1HCGKDEzbUnxqBTtQI2pL51OWpu76D4Sjvf5cwa0G
q958x3FGt5ZF1pf9dtC8I+OkANkxcAZCUny7zTrxY5e2tYesguFs5yae+ZfGfpZ4iCtZK5HVs5a/
1VI5i48/kIL+8jFXwwSJiavEimsjSYaOaVGzyFaovKh8vY/GNCCfDuvqCC8Q3BxYWuyrbeGwHNx1
D0Qe2P7/Is3ctWBK4mnot0uWsNW2WjzsDFYznk5UW2tCn37EA7hQzWIBcC8XwwF4PDcok19ZFnns
DCF1Rzyfi+9/3/PhazEsJrnSBjsKlhkkpplHHwYx2uSivOJ2V/fiCVqZHFeG0mhaCpjp1nXzJU74
NGo14nTYhWDHGbvovwMYxaL0LAUdz8AvA17kaz9eUuLOGalNUhZJ1gBFDz6fpWEzWz9oWo8++Rjf
ChbN3aXEeKWRofK5gpCqWO3i3rNcNs43hLAvhSc5xEH8yGfXYM2ayaspzO7wMDnk2vC872EgNDsJ
zjdNKT/R4J52AR0WGeGxjQaN5kkq7+29Q9TKhu1h7G2z47BPtMoBdhiC8GrkFKxiHiMbGXRpEFAV
KbnKND/0LLwPJ4kG4Bdc4LfyBvC8OO0nx9reKqI0GOUNXMuTH5an/eja5QzYXaV6HxdW08dsC5Au
cS8GXgz4Ds0gKMebmXZeDcyo3TmWFuvdE4/SqT7Jws/vML/uJhRDmeYlFgxo+tPoJVlOygiG3Qez
858BDfmawKudWf4ZN8Kh0sB4gCIIjI3vSdpI6g6Gxpfj9wJu/0oLR2mxfxG6YKd71t5yX9VZ2kN1
7G39ww2AVF3YVIg6fo4JLSARs0j4M5Dap3tzRoQfrOfhEtPGxzrB8S9PzMOs8/8vE6SbZd0kraTT
WNvbH4lClL8CHKS9lnUp2R3BrVII0qSsclmSc1tiFWG8OZ/1eg9TsFINhKieXZeiYhXPs5umk+gl
mN6FvGKatQ2xAe25+r1DevX+J/dRmKFnaZk4e7ZL2keiE372LIFmKcMgzERbkuKFKYvzQc/pqCV2
EYirnj+Wn0EYjDkQKfn5Vboyq3/n/mp7aps4+oL4TpfkPnRgH4N+F/xqhnQ3pNuFcachGERNU3np
Dd6FG4sQCBV9G5Em3S1L0yz1IXDx1NpDW+jFk/aKzJPd7zfh6dx56hWmgnrQ1UagLNY2+c5+Ua2r
r0qAlb1fCKvRqi4AJil8IL4jwY1cE2iAsZWFXQfc68wRh0ekOmQiQ07M74VNoq/ACfs8EVnCCOjV
YZbYaCkuJWJDuRP1VHAoCzXCiwNNrozZdPqNKgWV7EWQDvmGfIBbaSom3iYOqe0+UJlla2dWPRQT
6Fro14yl2fGa/Sstz28TGqHGHN4VclR2RW6xNsHJRBjkd5Z3ISYaW/oztVA0VqC5PWaKG03UJmER
zsyASrb5nSnEjWVSqPCTCEivtCLE0EsuBRmtlyY1rYwW8Prq7doSsmioVF9L79sLSbnmWyn2M43E
07jV35PmiMJQiBeLlH0PZi3JITUEPMWv8cv5FCtUZgVxixXRUmCpFi+uKQb5bF5dKoRXXwJtuWsg
ZP+JKzdw0HHkyPBlu39EGL1rJ6fXyT/ssc+BuluqrbKpdCQDlprON11xIGArd2H92OgeqO5kZQ0z
JdcatWZyCXTGouhr0RRQmffJVK/JWJysvBhUgFMm+GLGubQvnXvz2wP1lSxY7te21J5q32HkNNEy
MvVJ6MZOVLdXGDPJgTylrOwjqskSrXJ7LmhKphQ6mBc0tDmTnx4YhKpQ/58nGkQyat3xhQgOLUfB
Iw+l+lSh5dWT2TJoyZTrCwTqRhooO6QP2uesiKNT8EubyYV6sRKpwPwXidyZf0YlrenxR46STxeG
OD2mt3DV4yRyHbEBQ7XRkYKKd5rxTSQ/ENRWNlx5MbtRIDPBhRTXEFx6eATDq7c9LH9KX0qdVjuN
o8KjkaaopGvUghunG0ADqhoCQTKOVJP9Rn6tiTSu+d4rDh3NPbYsNfKquiCi1Allr/Bp+xL2ievd
hrnZ8JsD01BnrEb8wt3sBXJy9dRTZ9ZTnnyFu88RISPvXIDNmtZjntyXRSPxtouOSbkpNv1MxADG
H4FNinaefJFJHGIHDWQWkIiZ1b8gL6JChRuuZpkebpRZEHTtaRW/zt8z46PXHgwNnOgwOfJ8yluP
/Ee+tbDPAvTEH1d15MCw2h9knG7nhIZo2fN9W/kolysPzT1MsVDcKI93mDZGX8q3POnfTrMv3Qb+
8WHB/e+anFY4QCJLPcy0zDprqIoMdEZVskqANAZKq+dXoUqO08LoWpoNvmt2SOfCG9nljuTQbt9e
SmEx1AvFKj2BB91Ln0UkvR5au2uV8Gfdy/U5oVJ+Ecxsxt2YT5smKgKtqv2QvwjsA/C1QmvmwNso
B4tuuNFHSTDY4cBYi1IPPXiE3oMwAJctwrhDCSqhPARfDEufVAMsoLi6eoi6LrKrnOn4rQ9SFZep
O9ahOANCtskoUYyfNiXPfyc3342VGGmwGrqJ84hhN+qZXlZ+B1zBsRssW/7VptIh7iN9bT8WGNXY
GP37Oc9yRNkNkTk524ch9YPZQEw1CFv/snjIKoXjwlozoDHsNG0t4HucJlU843g1beCnbYVKoGax
cF+E4rTtWNZgge0dijf36jGvky6yp9PtVQpihHGsU4xeI5ZFofb5IxV0wG0+EQrw/+ie7keGvQhL
eyKVpQrMQ4q9RSV1w/En8FO/nYdHQX6xsCjsxK3oHzBGQJFR0vgOxk14RoCkm6yEZgCwZrDWyOx4
SCJJqHqjsDrWh+oSnP1rNbxgWGFAViVzh8HJuhg+983BAyMs4OU04E1HDAxXkvjg8RUM0+URvMsJ
rr8RK8dTNLSBIiI5/3IH6YcIZeB/n+EQb4VN8tameiEoG/XVPyM7hsY7k9osqhhvcNx+pqiC80rT
RBgBzL/t0Cjy4p4UhYEmoNL7BPBsDXL8bCglVNitsx08oCHm4pX2Zzzz+LhY7jlIHTXSEJLULNVM
iDTU4GlztqDGsdyMBr6fVHO97utKKaGVyK/m+yIILdW85UehfmIaEXgl7hA4BwRVJ6HqIS9nkQLi
F0xHQJEiluqgmtNOeMKOt7VeK0saVUplZojEabSUaS0uqafRlKK2YL2TcX4zmVjTZW785v8ZbndZ
URUUCC/n1+GoYfOnO1u8Iz9s1/HpC0/SpxXDSYNF78cTVwAmI+KEpmrldIuKK7OSaKCHK/apUUoB
pXmgUCNV/dTseix5N5CaVu6d2LEP5YPd+WnzDr+kBpHIAEM/gmYY+iA5YbbZtr4fU1jM+WORvXLx
DdFC9Aw+YWl1MrnzrAfk7yUqIF57eLRrpX5NdkHU/hHT+En+5/E761hDB/GVueFaSaDm4HpcBFQ3
k8pV0WsUnSHNb5opbR0mQhu+hxHsywIOaOBHkKhc8N0D7NsXMHonkGRKGIx19wRLJZYXFy7MRaDp
RuaV80HjVADKDeRVPyUrij38ijX8URqmpEKBBDienoEaEsjeLgVzETVsgdhj4SbkJrlEgMCmg517
ZwDJ/wdoZfvsWUlGDUtNZZtbL7eh9Azkvy7UZbDkSzbVHlAzMFkFja4xlhHIMYbRMbj0524nateQ
4pqvm2JlzYu8tMm0sOlpRJd0EOBYvV4z4K/WWmmfEuM53DOB1ukWZPtnqJ3vH/G0yrYu6oZf8D1q
iqs985tgJkl9mYm2xj3P+LvbTBD8/uAsacljD7lLqhHNBhZkvvatfSRh4YYbXIiX0JTZFIcZM4hX
WYnAxR/MVJWHI0zWVi6zNiyrRSGTITw/B4s8mHScep7N1Snmyv1sO67/OxALdjYp4YG7qbcIQTmx
8vKZLwXkh2u+gOTZp+nAtjv32VSDkt6qouMafsEJao+i53U8FWChqggvZfkuIhmgQSo5PYCOv4JO
3lq6vd9j/m2OtiNZX0A8teePAUL6Z+lkWNCji4SHkZxxkjeHTKP/aLj9J8pwcZSe5D0KgRulYf7Y
MFR1Mx7PXRdEoswCNztEl712DTwFWuq8ncRxRwt6UVVAZHSA/yKO1iOiyi1RwukScJa/kgB0lgby
dScMofQItgK2NfXLoQm/0scfnkl+qk5X6r1fiMzU/WGiOT9X+2/XQ08ZtVGYraXvR6zmx1tdt7Ra
nCb6FoLlwTI+4/BoOzy2WWezXGdkBd87ainM1q6ZC5YPLVI60JgFHmcUey/6GEW6TAtu/EbZvOGQ
VAiGy0H5C585FrsHpH4gXOKK8a60uhcx8llyugBjhWi2dS3YRPWwVV0kkhuN/61DFelBXi3uW/ES
9T0ipjRIxC9QxjeZKGXRlLLouF/rO9KRWMnXEY91HAXggADOxX+8X4c9DfUrKOGM15vQfiB6tFHR
LY9rIxyygDFMhfbz/bII1QJrz68b/wI7JBScSTVOiLpfuaUOukGf5rAKKw731bv005sZMgQChTZG
WH7zdC5AAAVctdcB5GkfszAXKqaVivEyTs2ZfoSZnYnFu2+DIn6FpPQnnlghRMIDy4DT7mU9dFmJ
T3CeEVk6PSCqPYtb/bJuZAzpkiLfVf7VWW8vn8Qak6Wz8ZxIqDcHVFkr2pr52j6g8Q7Cx2LFZygy
t9M2GwEJMhjZ4YE7YH8V2bg2tHymssBxYCkwHgfwmFSAmkaY89MzbX3ha7Ng0VbogGZzCIqRwEY1
v90Y+xaNhxxJTzyOfj9ciELcBbI7o1tWhOH5gDQ101L97Cop/AWMK/yFlyLn73Rad5Jle1evGAoI
MXr+Y/aw9qGVxVORXptVU24BqGTRTZlnK5hwyiw0zwyGLfC7xpBdKD/mcIrWJtXAjy/KuaGbXkz0
X8RsVHRrT19Aib7X86j3bIo0udOwNGEQOy0x6cn33UHPxncYKztLleoBZKtrhbmIfjLrhUHdPoCB
ILebxw6/A3aPISoUVIfwxAEVAkZTK2c1d16NiCg8xK+gU5dmn7xzXDyWEMIoFu2uGQrs9/DES3MJ
vcyrBfz1uT57C84FeJFSuzsk73PCVXth4r7AOl0FKiDhbudPQcKcoggBY909JwyCbAgrAXSIuyyS
TQfJQNBEcfIP7cDpfYjrrjhQKecCCjxFf8UhRnCPgpK+mSfffxdgJMZ3ko1nfOZYZ5v+4/T14r7I
+0xLmftHk0NTo11OkElOhcLzoUOrRxxStdD3QMDiHJ5/As6kaZsqIsKtlPIx4q6vRmWs3h1zwcBs
7uMGjl90Rvsr/cBR5xIZL14tOTKML+XqEnRpF2m8hMFfn7nuDuuR9SU9PhFF4pJFRVkMHGor8IKa
zbcdnaN5Y5DagpAL4hnMDJpbVRhkDDtDhYCHEUsLXWGhGIaiSsTqYp6vekR82edYnvDkx2HzxF17
UlVjY/SMkqMiYdmH64zL0h/+1Qz1vxEDPpMIlhDezDqqLM0wyj8uZ1eMJsWR5nuSvp2xLpBfZF1N
se2y0LAZhwgqKiZU239+82jTYSGOCSReuKytwUs2cvO1yC4aCR8m0aGJMifCvTJq3mv0fbpDZrvB
KTuoPfYLMadUwPIA5vXbb0jHP+5hULWxrcWk7nyB9UrtWtevjVmlOqv45g57dIh2MzcJX3JpkRT2
4hWBtGAV/b3AdN+uYf5ZIhdyFNF2etDxI4ePVgnBAovQaFUkKpLbGsk8gNFkICSlkEyouGoQuAap
6cswHSsoL6htq4BIKbT0eFXaq9ovgKD2e5ZIIqkRDJ/UewKO7KxYjW20QSbMbumECRPkK6RvFgEw
7lwTZ/pch/D8c4ls/KKFQrYwtbgKPG27nSixNY6/jlas2RTp4O3We9Vc5U5RE3k/j2hH91U5ZraY
B1NHmJJ3EiuBahlUxMBhNoKuLlJDWjQ8P/e7czViVSujexT5sqqLh7GlnIPpWDV5cd/Ww8+mIDjy
MxQ1p5gwTz4UGBVjGkk5+5Gue468h5ueNdcJiSX/eI4jERz29wLoBkj8bxct39gXQsvOAPg0SdzN
0SY6MaYxL1i4JjnBPMFws4ktnwj+s5UWb8v2eENhS4iWSV3y3Lf4Yl5h3WKfAc+rSAGcR4WvYRl4
lBCYGCpePsKTNn5nKvoLFR9EcoqhmOkH29fEDMWV/d3A4k3ImIzrDtfnaO64Pu9VWWokKFe7JJ+c
4823M2WwCw3XlPvKCemywB/hyTPGlsfdj7HLjo+OAojgcmLfR4ZKqIKPpEy1dEvXvkksYCemPUEw
N5MP2o6YkU4DHFRO1+jtz2CKqsMvMLTsEWfZhLQyaW+ngPTk5VcMgyv2toKFJB9WFpGqN5pacOwy
bMHrSmWFZZOp2fROhNGPOYV8fjuiHfB7pPvA+o21Qvv3JO79KIX0D6K5KVGVBqAruRzaq5do/kl5
K7RGLDCJKYbDEKQ2t6XVc/BAxvTssvyxid4Vlfk43McEXCt3M8vAO8+2PrLXQlgJID5EHV6NL8D6
tKBUx4qx29FrxBiLVzJF3yV6gvxCSQa5xeuRDj4txgeT1jdppw1SauG/eNgBDrGdTehy+zQc0BUJ
H0x3njEsiMYa3vxeAlcSJObyjv9A4f4m0p/j+/6qXy5vXjEBN/5wGm5zKom8pvkahGPJ17Nso+2r
JnFi64uP1PxqQluO826DT0JUaHMr6v9ZWh8SFBaartK7Yoq+UDZMzUw70eJatbXzyI8NZcqKFVtI
E4F0q8V5jBotRG3FXtBR/Gn6asXacbZQ8PzYkfEUYN2eP09Pv28FnbOvRgqk/BOkn+P45TTCIeJq
l/M22cPJ2k9P1ORmDF177Pyk0zxGItkE2aOa1qEzMkD6dBvzWiVYOsrXtr9BXUzxfAktxp57htot
n8UGmYuI0uJHIB0rawo1wVZ3k+dl11LvYzz5REkeJoFPTINeHkVIdH34LiHUJmyADIg0okubLtpC
3T+nUWg48U227lapU+qve9/zpWZqPmhs8PIpVHXpr0vXENXJw+StJda1aKTj8neCql35gBstkhfo
3AQpw3odkHRDnmWmBr3qZepaVzLR+35gXeK/KvNT7139hPD58m7+vHgKql8SCnuSYIZuJXHgIkjr
klDRLmrm9t/00eD47ubqd5g5ntbDV12mD1vNLFuNoy4ic2cJZed0esoU7tOPtJxR9oFDHTf7yisG
pQAePlFP7jdKhFPrAfaDo9HCcVpo0qD7dL0JfCI2bAxF1GpgwBECTLWbruEyGvrYFs5/vGLCUJV9
MrOEUsU++8SDr9UVMYpT4LvdbwqpdshZA/ewp0tuhcyBCjNQ3D7c3KRyXPHavSngoNW1POWR8U8S
5OPhGl+ZOidNPHQ/0B6uvKnBBmplIdGTBOL1eyimWsyfv7If2UhQddzwbZZYwAkaCqBPjxpxXnnu
8iWHHZX+qwxY0KnOnKDpo8yk/kMyUrvSmpfMIgitjFqcNsO1h+iqVG1lzwbzGORz904ZjYv+Ch4r
woYRE9r+ZOZv6VXxfFvRofL9OlIV70oqKcN/63u6hra8Au9Pj6Ux5mAZkV6WyjcrLTKqPakGCM5A
559iTQ0KA5o/fyXkIuy9U1TsXSJGhPLc1cwxzaeD63HGfkkJdLHQ4NGIIJ8WMERjhGDqdlwwSmvL
/MFJlCuPysrhoZMc7o+Yxvi2NxIL1WwAclD4a/i7xwHeUntsxdolldexMpD//cilBTGGfvEp7l4e
U/DLmzknNjbGVrZyoxFxjcGAHEqHnP4Djyexn497hyIykFzDY0A5Nd6t6ttYewBIEvDdy6w0Bg2W
faCc1qBMVUr+k72wfTFleAi96YzOKBkIrnGrg8aoCQPB+LwtLMtSekhRHnBqMJ8juVrpNseCTtzr
TwX09G/N0uM++qPLAQY3q5Z8wg1sgOMbTBiVpDiUyH5p+8bjj+psg+Xy7uNdtUoVRAtfqkqDmrL6
YtfbBgmByvCOPQ0O83apSKLLWy6NBekQdx0klKdjwoeRXT7dTHd8ePj0tKyEMrEkPmt0XlYVgZdm
rmVfKvcBes10DPhsQ23gLnLdfoAHt6COT+Vlkl7WzisugaeC+lTJ5QhBMJfKPUyRNcanmYj06T/B
8WOEKOeYVQKPXmDWlGp/llrU1vsdTOdGJiONmVWKv9Afc4NLJGBSqtRiRnZtFVszEGunMNkhJjH7
zEp4PHLj7kZiWurKh7GFmKDbtWyod4pEQK4FBFb1/DIGKADFKYSaFnFxZy1gh6u4BD5Xru6zgNcA
SeFvcyqZmtWruw+/RBGrZWPuv2bf931vtL3FtVYmWkjlxIUJ4/Vf3Y7gdxwYONtE4gqDehQEtCGN
FC7FTZrf5+Cqqt6EqrCit5MavCHA+9VTkhokwOB8YjKos1k+LDxzP/rYmyehaWNON9L/E301mon0
Wm/FL+CMI3pa0nk4P+DJkKtsK8UZiHOFBL4jhtbHODJZP6JwDufwAqqZTHfelCHABQ4BztUw7F40
oHdScHWwLw/ujo23vsaHnzvX/S8uIHs7to/AUOK1jO1yRe3KzTt+5vDQrMrsKn3trB/aNii0PoKz
h3/lt/RMKR/vmBLtbcjxQOtUvLfOcn4/MKwnEzo4iHVYFlTmZNCMjyFUN2iZ9xGMdox3FbRBd7bg
9hTVIuZiy7VG4G7T4nF/KurKYkoJn4VdH7UX4CD8eKhDDgrz3gsAa6NpNaGM5LLR/kn0pcUsIPZm
nmHL9xGtZTbACcs6OuFTmTtGGYzGuLk6aHFhxU2wuX5nyMm9jRmgQnVF8v347y3biIFlTtDC33NQ
dVWEfEGJbtCIAofIHU1IOtOfDsefHPaoYn3ywg6+Hv3Jn9HhXpEHToP1e2EO2eBMj1fArsBan8W5
AMtTFkm/AdJWN4aOC7t3Z64Q/uhX6PitLG0wRsy72O5l1Bep/LgyphFEW2gn9/ckYw6TGmWQ/WPq
vAzIgwAXvoTWuWsHD35m91I7ulsHOwOI/xdhwArtgw5ReeW63W+anKOzS9pc+4y8l/G026HcbUmC
heNo+ZFWVQHDrazhZZ3znsEo8TWM5VfHmXsi5JxF3A/8p2SMnkorGPzlzjIpfw97zAGAwUJejwO6
nMwqwmb18IbmF3lkRSxYPEIEvUY9GcP7wd431/8iINH2T11dKD+ZhF5mvbOjUUHpfnoeST/xe+nu
31/nSI/ETDJKQFhnulPZyJMu+S3z3FrLvrew2x61m0jVdgZ0xxlIajdCzwhXYUaOJCoGFcLvJZqE
DAeajjUwcElJbTqMSSLfq6IQi22UwntBKGFffU45XewN5oVyJb2W9BKuNE0JrmAUYszfCITu8uGL
LGw/P8SdV7YaNwWOimvprhFQSc3v/7HBUmyflKDAnVHmlb03sqfpRGw2yKTQafzv3h5/Sv9gJ4Mu
+QiZbxrnBBfJjV0PI41eQCaDPrLVUtOVNLLQy9WVeR/Y11kapZRPLtdMbYzrxMwiR33+Vrnu5vkK
OMR2i3SomtSckxVJbH3CX3yA81z0XOUu6AaeTrUrSjCmGSswalu+NWyMQ1/z62j6EHnRj9pO1dP5
+tD5OwLABvl95jAUsirbmZWlKA5Cwz1gQpPPJlJIUOI/jaE0hGKC/dPoFrpgW2P0hN1yDtmrHYuy
dPz9NUKyjYRUDxNb2TCFVNadesoVjiY2xYTUOw+BvIorNCDWC4MJRN7vqhEhIdilmy/kq5hXa+IQ
5d2izptYvNX2f4SuitwTRp69/n04qIdtf4BAWanmS4hoYeo5GHNcHIFV3lhayEngxPNY2UtRSocd
zKHAEWHnas/HzyzdQ8xoVwNIiHqDKS2Hr5EnMq/If1TrHLlcvnUrYii+bIBY/4AmakK606OyQF5Z
/HijSWAZLwntzQYeQ2EZ4hPH1TaQP7k2P0qGsP7NqANAgg3mrfr4idREKxutJxs6bN+lGquNYQE4
GBl2PqLgtcwSyt8y1bQxxfWI5LrziOpUe/WKhNr/V2+d2/eKrtQbvVlylk52kukgwy6cTNxdoA0e
cw+c3aByzNZrxoVmaErFhdWIc4OEHqgMsVzbx/yIX+r1GImrlOuQselaOcP07saJzoCpHVzoeszw
Ypnx8zs+tvLrdNa+iOedfxEYBe7gaFU+dkU1v7Jpe1PGDyDc3Lumu5cmsr//anYKJhFMUhE9bvnD
lmHnQRYH495dY5cTArsnc5moZ5DRgpYi5tRE1UO3ERfnkc3ihDfwP7wADjVBkVnbAcrAsy1FCrkM
AtFqm893TobXs4SvqArWNdR+3wgPluDFyCXthu347mCsaLO+qgwu2mMF//i922T2UyxVUtqIft6Q
MK9/7ywVJ7lxWPUyvoRzFC4xWLRPQyRej51PdfPmL7jvvJHYfV+YCiUyEvcj52Nn6coPZwU6ERaV
1xNcpl3sMaeMzvT6dpY2MNpnAvH7fUI+S1TfYUQy4C/GlQGPonWylr6WarcG4zLWYZ1mV23JYIA0
MeKrniuXmedOBIUBD7rWaxw3KvC29dDIMb+n1HeB/se1s0bcBMYnmHwuf8Exqtl/UwCEA1zl0ElL
HR9VZ7NxZUnxhFLktOZEqN5Cl/8jOO/Hrr30UhRDPOli5nEw7tkKX857UMTZLeR/lcM5DnO3T7i1
X9E8TOiorn9l431kJrtFAqC5zhsO6a4r8lkWBYiVpqZx5JqQ/c+3ZSwQTtnEigolxAUWtg12caIv
o6bzGD6PS3/eNsgxhTfk3kMvdCpQLXWxWXsGPQtGchY4aZJnW5M7dkPplXCDFz8w5vIOwh6ysRwP
9OZwI2pRx03o1bnAxgGS+9+E37lbH0U+uqlGruI7drGxFF1X6gvW5ctjqSmrPA/7yQ0zdw1hLMk4
MZ+y6A3hNK16doxtLrA72s7x6KU6Qz496NFhgq1kKiR1Bd7+p9bI8COEvny98sEhegc9YD1fkth0
vhpJtIH34tn9LMTmfBy7TLJq2vvKzCCY/eH2ooZW/zVsmaSlRN89fbl3EUbo0tOBPqH6mjftvZMX
K/g5vHESohRaG9/mxLxU972S8/cNHKy4G82zCbmwgTZCBuDJ2U3mlmSXstBUKmnwujndwt790Oop
bqfZIAhiRja0FBPRI++uoylqVzA9ZaS4qjhdANvxccJijoJFZXLY/YvI0N5HuXtbZV2VzTsXPs8B
j8JUnt/hSENGZEDXcysv4W14u+VMUx8844HzXykHzo54uvc8pNEa11hfbYlgJSWiBMpN/8Ag7vkS
azztfzX57B/xBWdqgODGJCxSO7g9QVwNYCOYcpIPjESdpvV+dq+NF7pVkb+F3p7fUCS98sFF0jg9
zFeSgWAo2l+7yWJFXmDTbbVCSWnBoZ3mbBLjXA9FR6gfRdh62R2EaB5byeSujHeaWV7b0VoM3Oua
Y3n+S1eKcdxFFox1nNHgr70zMsHCClTPg3NjwTq5YGDtJ9vhzKxTnXADmzyX+hMpbrWQCQ4SvcgG
R3KHngpoZGeRYDRWk5MB19jJUl0Q9RYJPIQJD76bRH5uamwM9piHcZr2CwTgmGmKKjPuBo3fW+H0
TGd05nnxyAqcuU01JC+4wI7tDsh0C6G3REWqheV9x84k/3puilBGbpYcsg2/xwTEe4CeG05xNJ5n
NhoC++ccnGeKCe+F29YK9t1oiSuAuMGmJXhtB61FDNWbxIbvjo+9XTqmsKCWZYY1ws37KCqEaKul
v7rkd57yai7DRbmb2+IJEZ6ftJCtTjuob2/P7yLEuY36zsj11tY1H9tVsn3pmmJAWO/10+Bp1t3Z
eSd1VxDJebuKSLWs+qhlzQihm9xlIIBupR8PdA31cbCCM/7RL6kRSQ8+pz0ofqWCrTdsFK0eJmvJ
YLFkX+KkGR3joNbV4OckwSNnPiCor5pM3n8me7mBwMBsdFOkQycvzAn7soYDKPMaokR8aiE7UDgv
wx3OPidb9bwRJK6zT33ZXZrjBHf46VDZa9901F0LcvGMpkT5V36FKP2IpPHzFxELgBNbAREPUnxZ
ByLFqU/MH0czaIeotcLzTqhjKyVmuGariE6rw7mlcb9An5471ghqthcIfXZTfqIKJ1ARs2Ch0pwz
1odNrl2o5yRg2NyykpzRfL+LqqyYoEb+KcbQ8japJFAZZ/Nab0FzP8Ra+0bHI67dj3JtrEubSH3f
QJPpiZLenUbWKFdX6iDUdbeHKlvIM+bHDEfyTeH0NYQT2NAV7ry6lBxdVNdxT4daefXMOsRnzMH5
nFgxkFbDltozKpPlzwEfy7nzwj8ltSz30L3DujLeGafiozIkee8VKdSasPxtkhleURNYhvm/GGFJ
UV/flte0NleSc894+rKLV3dKbWPREL5DPfOTwDifQvSvNRmkofEFuiR6gg3SLGhDrmTvDpuaLn1U
8yVRbwSXLkP5E6rVXXpZA7/U3NeG8RMBVvx+qpJfF+yar5/nRhJicdcDeDImdr7mQPgLOu0P6+iX
j8/8RZwEHu3enLbXNohWoMjgBIiHl67qxdAcVREfaqWnyWPT0CrTJi1JrhZELFGOCDI2VA402Pjr
1ZLgSj5zsQZKScXCEKFsaEUAkZ+sM+szwBWFilsDLMnxtpKq/Zuw08Axt/cCzJBn71e/zbgWfA3X
c1y0TYDgB4PBWTiBTZNGJTT4FxVWG1kP4aL4gFY7Y3lSf8smzwWTzTj+MB2u72YLJM5ZgtJhtx0b
2YEduh+V6tNOZuvuds4WvixdgayUydlu7RbCEb6U8rNupU3/w3hpsOOY1JgqqmEtQJzsh0NJrgxN
5DAttMnMiAmmXPpyZpAzpLpva03SL2T/VzfYTEKCM6/+afQGfKTZFSU9kKqx2LUX13jIzCzQ5OiP
EgtvmG1gydyinOVfc/9p9kPZ9lHrKdHhnNgWlaAgmy1bvrNkrrOxivV+l9TDXR8fqZjLM6dNM24Z
g19nF150kf+kTkJRxBdI2a/1CVZOLI9r9JFlm6q3g2y0AXws/TqWsfduyIBTsI0PgvsElQhySfB4
CW1acUICN6kUJfrpL8kdHBaU1HxN7QJE5PVUTQLByt+SGLxe3NYV19tBlY04MS7hHHNibXCnRBXW
f4RxXfgHhD/CJfjq4dgdlrWozPJUMR/bdYGOG2sfYSs7YcFQiA7SzwXO6Bw3oAcKDtKAv8DKX84q
C0iRY29IiqqdLYnvorWU2Ejr2EKanPofpYvAAFBdohnX0AU5uPleNOcrw38OYRsWAXHymbN5z+Sf
Iz0lJVNJYqVuvPiU3rNWjMOz1jB9VGfMtee1Nr+x8LzkVUTkSdttD7ptg4lGC90LjnCesRpHKUDp
swY7IE1NWE+7Q85CjdRc0a8IMV54Qe0CwsITELnc/U5/Vq4dhzrxy+uMhycnBB9X8dkcATjUltLv
X/IqmCqWN2sktZ3KeQ62/yJsZC+o4pn4v/l4didcj2OGwEwOYVsLqx8gjxhfEmef+RuoIFcnloN7
VhOUrufTQLgZX9xlMBpCepVZUGlQXNsjAB9dZtGrmMCfCmFAfkPDrOq4BDG1pUR9QQPZqb1FvgV9
rAF8RLnGH/j47WtzL/SwPS40FRIzUByn4RQXUrfbPth7tzOsaJ+CTyUUCzXF/vrG6pbKWp8VeAAP
azlceYlFQP+/FhSAKdYHiMHeNX+OAltS6SShVeSuz6UR3J8b7XkTfeQ4/yY4llZbptsMYz3dArQA
dUINtxTyIE+cB6R2BNwoydWsE432s+ZeAcQ2cIE97YKtT6IGwOW33hjXS5lR0+BCaLq3t9MBkV/T
gezsE4HjX6bjQ9KAJFKSRvGvd7kzQR/GiY/iSjkeb7NskBEW0ee0L3bMrOsSI1phl3cHRjpELv6w
yqKV1880qtiZBNqwuLmHaQ1hXG+hL2dMJOZvuLM55lw6zfDFlzIurpDT9DrOrq0Xhb24XHx0JXWa
wD6Iw+qEN00q83FSYXyCDYWw01T0W+L0/h4lNjqUdnY7HPUvNFn5l9W/sw/wOsTr0UbsU8XHRXPV
eQPC3qnKBihaIhEtPc0/Ouyr+y/8K+2z5m8+ewxEf2qxQNiChYtdCtLxjWD5a/Wo3ohGid1N5HA8
zHidSmhgFOK8KVkz4SGrMXzhH/01i6pohcx4CWNRlv9YGTGai/qNeWqYBc2+qe0pCjAt2pI+6ZrJ
3pLLbqeSP8lyGrc+SbcKdsniEaFJPKwDklV/ETD2/oMm5wpJ4B5tR4cvlt/KPwObttRQtWFCtrEo
AMp8GgYamNXSvF2/TMV8Vsnde1WcjmK3U2bfOy5yKJ065SWkCTN/SXpUVAO2sYuMvjeyPkCqhOth
htbTsghncAK0cDbCxPcrydUm2nKT2sy0ln+Oh4fcvo03WWrz29vGkXVy3clpHsubHbthGjQ64hpt
WZV6b9YsX05H6wJ4YwSbIofY6cujX2J9WwMr/s4rSH7qob8tjl3EH52xHOF9goLGI2Z0bQlFXqXc
69eL+b7NVwPHkO7ulAGpP9rIQJJUtRwEYu067sIWscr4A052JoZVCJnabSr1dZHlKjAEQ/cFYzS4
/0MUkQ3GjaSX9gZl2f6ZKFjNePpJZVYpxdvrqY5WQO31knzKHqSMc3zXl3Io8/RiLctWHh972WNg
mhwlzrtLmS+KIV6m8QRroUdh6onwYwFo4+ijI529GWi1FPYmKZMFnYvabzJTU+/pRUYa9ReNFB8d
nyKmy2wQIUU6QAqTuYGoP09uA6+1owF4T2x7q2chDY9KsymLd8JocrZSrgezwrsV04aMSCM1yDoW
o6tK1qIcYqEqJqxPfhcEFNSN1ukS4AIb+H01rujLfoy3nBWnuusp0WacytrolKlwChutYybHMxK2
a3YMiJZuHKvJsUiL07gGL8eiOEzUMu2uoeW7vFCRyiwIqoxnXqAARn7PscfXopt8rzBMOP3i/CWR
9FyE+DaaJyVJx6euPj16BeWHJsUu0ns/qFPqtajlYy9T0ib0tpi6ej3CrLG/4WmV9fCto//9hHRQ
CnKVQgw/LFZ2e/Y3m13iuKxNeWLeCdGpmdJZMadqHnr0AI7A70NOwBlrDCKQ8h9ior2EwDNBL8X9
Cra7cGWxWOY7kQw2LefFxUCXoHz0HT0KyvgyS3CGKqbZXR/UTtSWcBfXE3HOQyQYRBOsevl10NOV
tzmys72JOmlKnhGdIAsb/DhdiWu4eNG2Mnd5sy87XxpM12IWIkhCKoPIUX74LKJh2X7FlfeXqfwU
brtNCdFsu4QB/jeqhm/7QcZ2Qr9j7jFV783LPWjIz8c3fmTh5pgUr9QqkkDR5C+GUC5RodWt3O4W
NRGHwmRpMD52eVIiYm9hSh7JqJF5PuxgCyMb1uHM6m6PtP55hDOrmxPrAj5i2iIlqGSFmDb3tZ4K
g93ESJjsE/cW22PB+KA8FMn/X8LGnpeeKJtWw4goFKvAGuf0h5P3WyHg0xDEh0Zf6aSe2fSj/qH+
2WMCXtnGaTDESxGG+fvaMr1iypcAUxJyjLtCMvoD8xp/tnmNy8BVkJC/5sLQJRWcfJw9qFSkxdEl
T6kQhWFtYZYrO0aVm0tZAQQT7TwJ7tyAn54oXz9Li2JFAcOKQbQyMjHdT3XL2yQMch8FwXjs1uTe
DZmGQBrftWgj998PUvGunJLXiAL77QCyPSCs3v3XqffzEohnPfjstzvEMxI9m8akjVtcga48egIr
+U10dFt8zKs+rxJFseerV7fkm7QnNQsyKwySKIDxYzZQ8JjjJd4EqgMgewNCI/lqCMP7pvqIx0TC
MtUHr/HFYEYuhvvOS02ftfklfa6PMUZeiXjCe7xic1GIOwS2remRZV+/7uqgObbzQDc4x0rlIzge
Yw/+iIuS5RCZhcWkwlddk8TNWo4XMAZzhDhMfM/mJ5xQfc0IZ+eGCXu/5eQzBrvdu3QzZYn1gCQK
lUsm2PJDqVAecLHrRvsnm2tOXAzHD6pSZ8mQGc5xQx6z44sXDLPndQGJePxKFjWt74Nmbd0HH/Ui
vqYeaAv9RI2+xnYOffiVAAwkkhEog9oJ16LfJx1IhldPLu3agLhO3aam93Hf3ToevgJ9gN93T34+
WYEe3jtrXAQ8KmriMSAwEzVlzuOkI5f5E2+qLiX4AhomZzOc5Jg5KdTdZTX04Yx/JxcDF0bL+2ER
5vx5QkhqUXUljR5xtEKVGrnvReHWEFzUkdX/kStk7mfg4MCK+f2m4GPfh6G5G4FUZ6Zhl/jVRc6I
IM0YdAmDsExeadxjT8crQxc+GJqK5jAZajj2m4GV5Kpz2eMHKd4RMYTadv0MT1lJe1sgc3VZmIUQ
6znlqBVbKfeafeZ6oZPVKf5TKVRKIIzUONr6hfoOeA7nCqkiZokHUS3uCwfIbrE5LrrDsAobAvTk
PQO7nM7Bpy9D4jjyt2eDn7rbI5ifjpZBZ48lEvc7OpAJRjyTPGMrLMOxykhGranaPCX0Ef6j5A+L
OL+cD4H7EnNpRDIFIKIOev4RtYhHL1r0+7K9dV6aNLa9T8mW3ME42OxixbuVJt/cph3iQ3rlXeVR
DFpRB2zeNHIHE/S4W7kS/SN4QiVVdTSpOIB3p8UvChLOzOqettsJmXJrlNu8XzA/KS8ord9ubHqk
9/XMyfoHh0uZ8taVAe/+oB5Mwyj/ivto8XX7LBTIX5lWfi2zFnvcPsvZ6GDadqnwT/9RhHajRd7x
aC6+NBJTtfDC2O+vQ1iBzmlMInKmb3LdtCJ7oc2MQcUeDwsM1nyopNaZTlMHXn1YSq/nOyJVBvMd
0DKos1Z04K8zi/MsYZfHbxNMd/Ox0uw+6nXobc+6IE9JEW6OwGJM8eeJSfLKuozveY/sbGAfPMHR
IKUfpQLkMH6mIXSlIRMdHS5qXpCMvxkxdA2ITULH3bq06T8SeS4PWa+/YUy5pBqMAzt1IADHRy+6
Cv5Jb2L28nF/i9PWwPu/PYWBblwyG4s7dZqEQ7bh+9EYNMe7ZudiyDvKHMTl6EzZa/rOZxm0LGoJ
JZxm9+UaD9qz9YDgyTj3UKkzN90QaficoG2OMaFtUgbBec+8WEYTh66lBKL20xcMkQfRN0C2w0OO
Tat4F9qu+Fh1O+21mLpMZ+fcNW3+GDuX4OdP0ZexK1HLxM4IUxTp2cswSGFOi04aBLNRsN593ct/
wkOkyxxSPMpzdsIgQbcZVS9qbgKD/ryp5QPOd57U0kz+uIjOoV3ytGk65zZ2Yh+TChuIaQA6mLDv
7eUCrx9sWjdwp8Wa+8zEbc/mxvhBKMoaA8zlrcvSuq4oQGfgyjuwKZy7FJhZ5Bmk4GQmzYUzY+1h
vy+a1JUzZJ+go4dUfiXvZ5m9C3w7f9E/9r64UyxB0jrlYuBol6vOSKmjjqSHXbQmhu4OJbgsgV13
DsZj5+7JYem1aNgNtvJu6zejRuAxAceO0ML+2n13T4E0BNGZRMt/YwPxgCNTn8jHQcQ+Rio40s+r
npzD3Y69fgn9Tg14T+PRKcpg4PWMElUelG8HGTZcyjHrnCtAr0Ix/ST08GPCBkUTg1STTbhfKsbe
4X9MHieD8JgX1MsK52CjWkPSuY1tzX10egegaDhW1oxJmsOsVCe8wPNa0WY2gYJRWPXs1fKuPOws
110JxfIeeSn4AAZYI3IfTZM7ZRkAudu/3ttamQwjJT9sPJdtD4G9L/eo2GZxNRO5A6f4XiDTgJwZ
MPrUbuPsp4F6atJOwIss1kzamrxxbj5qevfNXfX7Oh4PRxoF8UvDXzULtbQdx2ffES2qcQcD2TFQ
VFA3dFbDFBxtyPUL0vtaEgBIJlQtLBQh6+tqVdhdkHdH8C/Ytqa7ZdF6DtmQjfFEcjjsz41Fkkqp
JNZTVit2b9qjU0a9FPoevy4NIKilESlJvWuaKvKbUcPtbnsK/PvXoIL+vgDSPGsJCbuUnqjjzqU4
QgqLPqEs19j9/WI+eW3QoClvdCG5ccwLXIlXuexi4nLNVzhCbYRjs35bz9VZJc/47mfdJHhEFUjf
1SJ0oklFvu70Y0cyUOMMLYVDDRHEHe0UGbmwGup5KuxOGDDS3x4ILbc/7aqC85O6zqY7BBwTpI6r
j6y3TnZCHGs2pczfKknhb4LI6A2G4WcTHHqJ6+MmKd4sIOv6reeRgkv4Xuf2G5kMdi+aT96ouCAK
BP7Htj3scdxja1dgaaL1oRiiN40DH7J/DqFN4ydoUo9RNpbsZCHh062ntlJWtlO4GYBQuu1MEsjs
L9iUUGW+r+VM9fabMG6gnHqGfWUUGfPiDWxsDSzB72QyNmigD1eN6T3iX2TLN3zEq6+gmqt8R/4e
CBsRLD6nPFYBGC5VLtfJZJF6oRoe1WOzQPqfTivxaKEpTyRbrFd1bErX01Y88SVWvkzfEcJuMxmu
Upb85/1rDVCjZ2Il4GULiXT8nqutD1XhbLSXhQq3kj/WRk2ogGq29075OzVLuiqT3p5sgXZM/M//
9QtdqckzIu61YqExwiVynJDgfWbUyZowiMdr1vF575RS7kOXZ42iMlgI3zbavR1/0HhUIskBrcoU
p/fw/6xcs7iEAKQWZk4bTLddBpoMv+4N+rNeFMFdq1P4ZBMNkGBZqBDXZ6Ut6xDVVjn+ly7Og1it
3o3bD/YZkCBNiaLemnAHck4c9vRPHE5l1S9SPY1FZn9Jr2vGiS2HZbEIyx+HtCBX6P9/tpAwkfIB
JAX7Jw1svNGYA+p+ry5IV9wZd+WEONo5+foWSjFbQcgnejNfMSN/9iU50gnUEFUbw4sSf0vJkWrb
2cWrENTiwymj0B4De/wJe1oe2owXwNzIkx+UM0y+463i0t93xeemphUpMoP7Roktw4tyvRyAXGhS
VWkg+ER0WBYZ3d+3U1cWCLPka378mAfZ7HF+KWmIqF5zbXPOUcWzRHBnUnc0ye7ZosomWpBrw+4D
AYvUYS+cuxeElqO70KMiobzFiU4Nsfi6NKkDbycEFNJjy7vcXCpATckK1yirwVHu0d25WPjKbiR+
QjsaJMBqqJkF8+nLjrrc5XsSrlwblr/ztNfI82cY3Arft2ilr6rFo0ge33nTjIeO5UNaK0dU9riD
IeZ2jML6x0T+IAY/5XK5a9IP7TkW2tf+0w65GOPnN9OSt4OgLZhOMVAiTlGafc6YOZoERL09/ZeR
Q99q8CNLXzuXCmI9Gx9teM3gMwKCoNq6wev+Pvb46/f3Lx6IzDHj1H0Wu9kHR0J+a08TIkSdGHcN
xJIQKxRdqi4obNnF5QbJFpmXuAV9a8NIssl8MRxvsUnekaR85OhiXFofLfxbzoExefDtYRrnyAaO
PhuhHSFQXyYR93akc8nt8Er7dx3WtNdXLwPwUj8OC7EzrhjKSLrvoJrqpZtJP8c4r5xdw8LrzpZd
ZVcHsujgajx5Jw40o9IshSff4+iKxiQOw/GusRfh5NOHObhxT77lp0nEjN7Di2JsGDV76QThtRst
19YW3qAvFhd2VtN7/s1xZvyqLKxgk17JaDTWeDe0I9VP7KtiiN+6Eo4IZM2K3U2PHWDdOes7k7EP
mNpHJHUNGZNPP5OLbUMW1NQ/R1o7xHpc+lumqnbeoHjO0HRTFzF6PuzLbABLxAHc8VL2vIgorLnA
mC6nvNPKUnkkUYNyA4DjiSNE6LVvZNl+RLJAELt+tmFp60uuu/n5n9tXdDih6qYfT6PgN3WOjzvL
w91Ankxm/ynMTFKFGweUL3NjckU6AUUu6MgpImSXl6uCdaJSfWPExNT82n7k5dVzOEJ4VOxqLjHn
V3SOpGfW/96Zu6qpkdqsnizV7199V6RixtAYCBOYIdIcdRO+zARz96DyAiJYTb80q7/wiosR+FqA
kB2AEQYfSk1aB+iCdQW8z8EpCp4QwsmxHEz9vBw9xF3ubw49LMSbSEoLobqnkR+0v//+FFAtDZ3O
uDSJR1R2WU5dyfoUmc1+3nwjiD50MD1ONfz+8u41o9crMMIQ0y2ZAhtlqBtxwFKcI2xsL+gELcrd
Yl0keQ3gMtv+nfOrGf42uRvX4rMX3ZRzxFZM//yeAUMhf/flBtzfsvmGexKW9rQZ1UG7JRQZ+sg7
KUNIOPw0n2rR3bfi02aqbI2AXupBvY8J1FMyYh8XG+YoqITXxEImPFv3WjShFPAtq37ATtXQef2Z
+79fnpeyc6jlMTlfpwFfm+orya4XsCID4RdRzjihrsNVDxVGG3xOdTFLzFDkE34MCpuI3vkPehD0
x5kgmk5utqArPoH4B1EqEfu3AVAS5rU9j1+GP/rF5WwqTYOhu80FY26h4aSlBSRTbPjbtlT+gG3F
VKkRbply0wGWJvtczbUIPBi+b+0QfSgCdp411nWxuzznfB4kSFHNjXjlgVMe7lz9VreCWtWcKtOR
y7MyhD5oYjGXDascsc+iZL7ZyRec7sBC4+qMDZGoY+icUM0dVjjhCbgoQr4Rm89vvaeN1JiWrQ0E
6dg2mNrlDvF7FiwUtJjNWVI38ZmrIZfm/TidVFKlpkn08xo5sNdo7//NjRbBeMCoL58jd0ctek6S
GTuOLRQWFIhmW3uxXnlbDsp/eMTRw2UXtV/aDIxmlAX6jKZvS65YHBC6FCz8v3g5YQt5QGiqsMnl
JCdp+sapRizYhFV9y32Wk6WwT+5/Y9objNo4pQ2H+Xogz42hknAXpODc8HB97oDtnOFMZsRvzRnN
pumr8jUG53EIUHxJo+F7z/Rxn8bYgw77lHY59ecsjLUVCHdHoZ6c4ZNhaAkx+5V6I9IAY0DSacug
rI2Otsu/NeQCd8NuH/H9uI4njjTnyOEXQVPTUaf1e/4W7Up13U2zTq7KEn/BD3+lgzkdEW3KPSt6
fJsnRXXUtW3qKwbK+qxT1I+DF4PX1POsaHrSrqrnS0qHHZ/9/TgYG4JH+OKs8xT7ylQAHGY2H4FM
dTuNXK9zKsKFIKXPNUmwlZUagiXbf71dLjBVlzOsG5+wuvz12ECrb7cFYyB/Ap0ey0dyMOTm0j1N
xuQbusQN9X6hobxHsfrp6+XJak+1txs7TOQLcQby8AlIqPlowZRGTFMnS31ppvGo4QGbVwz5EZzy
28nCTnfAf/OCcgV9Jhz36m34+sTkuv4obGhM1gKsHD+xadA+4kOq9dvMgXgCk2gWVc+CgAxrAuux
90C6IBsPNqjlssAz8znu9MKOTcOZsu55/4ju6zgFnM7IpR0xdZh54FzUTREWyTHvNM9XURHvWOoN
50aTgRu+XQ7R4/BriCuw2O/mEQsIusjtNB9Q5pXd+E85D6AXoUB5pGQxGBhjIbkdISUqlqoIJG+1
yUJy8n+YX4TmNVwBzdzRcC+kTWoWRbVVrI3rs3zZLuO3gPhiuIYs/aeoYqxd+yFW7VZlDMrCufga
k3ysAhZ6el8jRUHiZUpyR47qBaqxWlux89npDXXgTQlF5IQXaQ4pBwis5jiSIKveqAaNGA0cHb1W
+vnjGavnbH/CFsJ9O+dqDFuApgdgrRAc3+anxsRS5GorcPM47FgFSSy4Nd3deiliqnz7ffynCJJ7
eRlTNqzNLEC0x4dPGr4o6BZcHdayPmglQFjWXR8MLr4Pv96j+39pzO3aCziJxb6pebdRmbANLXYA
ubsBbId+ESw9f0vUGJEmpD0bqfoPFkTDc18KwhHnYVpP3tiKKC4JpaSeWGZ6Pzmga03ph1N3N1mc
S2WBNSlOEgKtHBnmKd9gJSiGJ/HytWs8vVOHyKIo/63tRA1uk6DCVwEp+DXYewu5dScrX6DDxTRh
M9e6fl/5iubq56owuQ97ZA4u7g5BDsJFjqSLvq9d7o0FqPTAaYEidW8/d+skS+lENB0hYvkEyVdd
CMXu8ciEz+LEaPC4QQcfMbThMEk/dMGkPNFsxao8mFXLLD9uXSC2xC4PYSMciIIIyg3IvbmKJDNN
r5DXxODcBixQGPEWelbnUm7EQoyyuZbo79yQETz9neI5TbDsp0bVxJGKe/jdzypwdeIVcFWU630n
pHilfXiv5X0OrvbbNf21JDCmUKt/o0bNJY5RLIsWtQpvNmD5/xayVFx4Leeh9bHHnIeoPaTas8z7
L/ENiOHkfaKgE0stBxO95aBXvL5P59+I0ZbrTfCq6E1C7DusKCpi4qN2r1p3UZVLMAtvv/x93jr6
38qVDBztk+7knFuf1NQNxkgEpYOY6WbaD9AOutDb9vlMP5M/F9FE/cVPcuOWMJST+ZxrnMzK7XFd
VCd/fYQeDUx5ayNQ0Zo6WnWenoiVdMXjKeEcJ+RF/yJ/XPW6UGE8ORxhAPmp0IT4NhRM4T97zuvf
8zrUZOIlMKWXBluElfPAK8kuhZaknlaFunlbi1dFmpvu5mB6vBsvKPbUUR2gm6zVyw1g2mHhEvUP
UYbQDS3zy0jkBByuNbYDamKpyEpeXTP+3Q6SrqlNMxD29n0Qpb+lJFvlydwsTjpFB64NEKBoTnaI
Y4fQq3zCbhIePiKShDSP5JQWXyBx2y866EMHNbQG9I/72ZQKjyANBjjg/EZqNBgQTud7M4mE5jc7
gj2ig3ZFNYlX0H1D2E+Ufs+1Kq9IBh5omw/bauqxXX7eXy14Iu6ixgC/BKNjwKceOMYkRumyIjHr
uCzdPmhczJXlsD5tGmuKtPe8ZxxZqHQyA2pB/ptiPwlJ1q1cVYx29P8FaPEN5Su3ozngLoMw4PnE
6ax+Ma+WyivKCxufZkAMdgB4ut5gmVaLnr53fZ2vR0hrn0GY+DlSJyCgpxXID5zcE1C2b0bhRC4Q
r8wGXyZjRNpgZ+4qReUa/dPbjBoJdhkQ2dSBX+51C7T2pP9JdxCRsYXn4HRI+wImDM7s7l7Hp93U
gXrZxatVHKPneANRJNP84jjhojWJVCTy4MYlSnQWM9RRkVkpczzF6DxQaBY20GjZ0zm7SM8YDkSc
ub+LifvrITmWsaO53I4jXDLaddcIef0apYVwYjy0XJChfIjL7OFIhBekcfQOqpqNFHvNdHYI8kUB
Pok368erlJ9vu1KaUSryW7hTCV1LvVNcts8xM+9WuNHrAAra8y3ysjN1lLHLEit5GbGls2SO4d8x
QntUmhtogsG3CmwIEEw4hpeKdtIVO9Ymk9PyDLhMyoKGgaFSx6PgM44Dokd24s/e14Vhrib/ET46
1ZqPN7GN8j3M6bRjfsPXiK0v1FwFJwaNW8zy2T95FPMsKTWEZtFpOaa7jt7hvoWFOO+IEJtGf4qT
sixga9lbgnVKrcWb9k3OZHJBXqjxmF8i5E0BcDc3tOul/zCmQHQAA+vUrBzaj7edLBUAOaIKqo3G
vGzJpqI06y4ssemdQfIfCdRFgXjMFJOe1FExuhQhNb+3A1nbuRARjndnKnZIKdlAne/GUjPAvO73
bYQiImAqPC8aS9BBs4wd/eKf8DA6CD61T1GsNfQGA+eepFCP14lA/ns4bsuHuFESx9GTsS/vdlx1
MBMlKmc+ghptGjsDrzX69B+Qc0KGC2X0+I3er6u4QQqQNDcjTJSwa65gDNjI1ewH60ea9NQgP3cn
+vCQ03RMdv4Np2LMItwgUDfHMndT9+nJzLIBZOzrCC67aKcLLpvvW9X+2mJXZY9oqWL9Di1wNPI9
yZlg3yGqAKoWwOY1e5OVYW/qiqknZd8KlRqgG0xWbq2IWirndJXvGC/jQRAEIeM531aLVUKT8ldk
eissddF19HQD+w/KGtEmBtUgKxsc/ss9or1+/jBnLdhwgRFXkT2J+XfF+NGWf7rwvlvKjgX/U60q
Dv+KAn1xBXM44zuvEZUkeseFeBz9NnO0VbbqzM7z7V7GTq0KWACW+aAhqtlT8T1FJw+SyHXuGkFh
v2aEFcUAwg9ic2DEnBTY6PejpnkehgLIXEqqtYon5A8i6CICM86Tk5VsJuaVdP4AOoWJlV2ORK6Z
j5otdVZxyzEKKOv1h/qJcG+89O9FzshjXQDEvqdcgxDl0yQZdqlTUGc96o2p9gFrJNsczPC9gwQ/
u8u6Fzkb/1FS4vxSlW6VU9SAY6muB7zqBq5xc/CwTh4AoeWrEFirUwjiZTsvT/166NyGCSEg76n8
0Mz7hm17qOeB7FaFhPch3O7cSzGFZTnEEM+PcotOGP3L3nokzZR4JA/7LpWY3ogrc2eXrGWCVd7R
H2LugzxpsLCxjtO3NgQvFtvnSHKyMyu+CYz789AFlMSP5ZyN1ZpdtkxIgiTPz6fnBkO2viq9l+rS
DtfEh5Qsc2eDcKgbIwzmSW/Gg8fcwncRPvH0uD91tX1lobw8rYOUGGSJ8bWpXAfDhkpKHvPF1/cu
SwC/tDeP5qgGMw0hEW3BsZdpLwIP2zKO9FOIiX/W1JvWiURHkSj77lXL/w8eD7/31kCfWMvomVmP
UVPYflU5ROBclUCJ67de5SLLUM62Y1VWMEQbkDG9u2MC3jgG/z7caCO3FeO9Gd6U2AoMJqSigP+6
0ejJCkdjSutkarDqsNoZEGXtySlt5P1ZnFuHkLKRWXrSBqgHAkRrcxNc/s6Ey6OF5fJ3ZMgR03cF
yaBESiRy4vzwEoUhqfUuzb2FXcAhp/sRI0r0lYRV1WkgW8KvzBX9EYeQJstDk4uOK1rdBRlUvuUR
AfuHAHKntZnUIzzRQZwG2O2bBOzR15ipvyS3yduNYoIEz6uZ+w/1PCBBzHkVCmeX+vWosc4FaSf6
P77JK2QtRZSTKDLedsjprAwPEdm7B44TI22di/fJGkZwFqwvBbZcGzOl81Ueth3w4z61Ny56YlKA
J07eN2KUcaYirnlkDq5iLelRNh+kPhBQ1MSNPa0cvEaIWrbwEsTHDzeKOvYAcy/OQtLFzE+PFU8v
Iw2uqaDT+/9K5bnmjyoLf5G3Cl5qaWjS+qF9tAmv8j8DXOT3zL2LNyBaj1jhOWZ3YQ46jGowdOag
cdwD7BM3qT8MTMghF4j1hOlIB+zETeFS/eQ7oqOwtQHzLRxp6fanixetrRwD2oUDvOXXBQCg1CCx
l7AG+4/7Y8KuDCAOsNK0+quu8LsOV3lb4leF1YOAgIiery/96Z0EU4AbuU/HCFOOlJk625DPyHpO
Rich+A4rqwEzPPWV+dqe/er9fHbjeX4vHBKD52jLC3MyWwYFh31hCjtSmk+OqD44XdfrI5jh6W0F
g/McsVr9N28ztdZZEv8Hyo6vLBDY8qhTpVDK/gjYksl7VVT1ZsFSxIA16HZC7HY8Y6Xflke/p2Zn
xekWe515Ot8+u+mZfA4Te6f4c7Q/7CNeSzK+6hb3PIJK82RhnhgUi6K53YzIgSoUOpZfrIxePSV2
IKbFJmyoAbfbwPaSUWRYfSEgU6DtpPUqTpypMIbS+pPS//IrOqzQeSEetN9XjImCQKndsbMVI+Ii
R/WGsxqSzQkPbbUOys4tt3pJoJgiaDKSt7kCfF/ARMwe0xAR/qCCeRPTJQUlEYygUQekR/AfqKdm
vFKmhzA4HHmfyJ1DFa3mgI+MZnOH1B88xB8AKlYS/2U0qOgasb6rYqcmNEYRKPr4ckjEMdD/aGES
8SSU5/OCGMYpHbcgAmoJ5zbtHn/CZmX0+HFcbtBOFwsds/kIDNuHsNnrtmF8xdt18EU7qQ/jSLb0
uChbm3Z2EI4ySLCIvAU9Y2BWKZ9rHr5gvJcYfZkao0loWcXeHg8Y86T+RfwUgtWcaC2Oz/wcsUFj
T+s7MmI3eYiYam0idrO9E7Ea+W2ymluvZ3ojena2qm58dDIZS2VoDUSPyb4lMKrKUZ2E97lsNXIz
b07JHTSA2Ko2Bdeg8am3BjWrPg011j87CBldnO++zyyZm+5t/xGJjnJ3OEUkXsjvXUbcQD6dANM8
g+1ltd1plmLqKbFDV4ZAdePVb7ubuYrWdA22k4XUMWXVN3lP1PsvVo7brHib1I+IT7ZfBJwCOKrw
+a16GDQI8BntDJTm862VXQlNwyYeUSIRp9oFQqAjCllMi7bPYGorBAAOGrzCpWHYjgbmjn3naYcg
kaZwNObOx4YCKR56mzY7vOeIKaQ7qy6n2Ih7TsqgfT2h+UkzdhLAC+OwQqJuQmgVLnYhalRqXZxH
jUEaJz2ER55qwuJqzIcMwdGN8Fi7nCwPnpi75pi5VCVKnSOSevnofXqr6o0B1X8x/lvYU10IrIRS
GTz1PzotNQRDyuG5chK6pkCdGuKl6Es0RD0GkrvN1Wz1y8dbItAhNUE58JmMOPPk8cKHvHkk5MtS
e0Tb/2tKM42/OCVNAMIjGagwWuVCpWL59nfzhR5syrgF5/KG0Wr4fjEV/3RmchBu4jazeMRNTOxR
N3/gH1uvya3a9p9DTvMoNGGKfeusAEfgUNdM9hiSjlATT2xcaiVIoUpBGJ2lagjBLU+Tc/GcTGir
DI+V34E5qNNi210RBaFsTRa55Fsk/zA65iKMcicAhO7H+Bvl/XVEM17oougvUVBcND2yRA7ykgTh
tjawPo1dSFCVjdQtjQbDpeqnfm/U6yWlwd2lfSAuA5gPqYkSPR48HVesIE3DR6Gsh4lHqY+lvaMA
31N5UI4k/VnZH0Pi77gLs/ryJPkrFOWrkee09j0n1cbW6IRoqEpxpSlDfjbwHpX41BAm/RnCzhPL
+UNAOW15JVm///3zmVJHrUTyHvddmSD/NIQk0YmTcSaUQR5yg3f0amsOuuLO3y5RR2DD5dFaEXUW
Qt7Zc8c3DcZLAoixDjys/gIXJWFKhdKdHYPh9XyX3fALiGnkrtN1Qhi2bnmcM2ysiMxtIirp/6Mq
Rwvl2DoS4d8yigm3VwDhINkwCy3BzcVAZo9v8607jEt7wWPyJRfQH9gn0wVFxk7+mXqFqZLYG+03
dqwaAuqocY9aQ6ofBYH4ksiGvzUhVFbxlEh+xIe5jVJzi0jfQdbukDQQ3zRoXs29YCXtTAuGgR2P
MNEcrwnID8rN30GlsamJ2ZY1aiqgSLOm1MEfWlWRH5JWccyN4sb4/3ULJ/UzhEphil4tsM0N5Nma
W29TFLNIgiXx0rBHWxgSx0DcqD4Thhs5U1vwzKf9w/ZEslch16E10BBD7Jzf0VWKSRhihZWM8j7B
RygBCXXHGKw7AfZxBMV1saca/BxIosSO4uC6PgqCppmfnG0AI045hUOf76c7CRaQL8PMp2R6CQSO
jfHPA7+YU5i6xc0QVqmW7DwSKwNIBMoiN0xhsy0qC++or90s/SpBJx8+ogSY04L1b4DEg7pneYbA
SwxKtF35gBwQDePZOqQSIjoYFWF+ZITT467IR8symBlTADb4m2WdEgt77c3kRaog/C07Lx1vg45d
hBndlXYjbxr55L9XUNv91yHMFr/0Cu0Elt9edtWaKrDNPq+KORLbHOuRsLzn51IttKNwx/JhWvmD
DQObDGAk2rU5hsg4pTq1xKu5eVpVDVpNb9+jjw4ak6sI77xkbLu5Yqtoaw+SIuTDwEFHUeqgYlcY
MdtudS0Wys9cB4+079veOP115IsxAOk7WgcsLDy6s27MLUcuwBRL60tJMLCcxdIZAF9S64NoKZn5
/ZllC2hbjEmm9Qo/YONag60BYir6xhStlNRgcdeDAyk9ydFM2Rc2lQE/L5pWb9RtB8R5+eCHJu3m
oy6fXRlOgUfYjgAvDKiQw0pv2El+vEgg7RfhdL0oEmiCzrs1acy1GXBDRJuZGb+74pDC+5dTgsws
A6DeFyhuOUjjHb7fGSecF2MTvoplsRppPFzrVo/S9Vpz3PJMjyP3FH4y4gh+xGVUD4mvqWC1M6ww
rbgqUIYI1MND0oFARFngrQc+gn8R77NFWPzMTaLiJo0q5PQfTsU04pXkeXHvzGhxfmpDZEuSvbAs
leNqwKd99JtUQ0wLfalvSfRSAb8knJZZLyWOoICqsrUxP/EvOrKRfDaat1b37ARogOzzWuWSHCuu
ZhnNHEV+pLcs6PA0G/ca5NuPxkXBmNNueMQBGFqRLTapRVnhAKRGI06eQvhsou/t4OSMd9kd8fD3
vkit2YCgWfI4aK2usxqwPQUdO0diHCX7dWQxmd2VGfPXGPsS0u+DT2VKw5CZinO/RZj5PjDsSCN8
SEX32CxJqwfJlxv94ED8yGRuP4IwawGovA7pTrWEcN28bzZgWPRfXaSKOPRLlBH0Kwv8BmSwXraO
Hxacvs2HyvMcsEWabBLzS9UrEOJDw97/Klu7xrti7UQdasDyLN5o3f2Rh3ImSzZ/EZz0GCjbheov
sW/noyCdW/W+f1qutuNaZL5KbMxYqbXSMSMEeiHbo9dLFiTGk7mKk2jhGF6I2VZ3gZ7DG7qAy4rB
rdZ9SPD6ytZ4boOTpG6ohXYG4jblMiPnz+HLMBmxbAswuPLNkyRoiC4lx1XfV8fUf2pSrRDV8ao/
K80Don8RJx4DSd1rsho0bzHEkfXzhYTad85iZjasvkQccGSK10lgca3LsT/FUuycMoiyiTLt1TSq
Gj9GgqS+l/J4Oe88dT90ANSETizo4wnDCYRQCKZGeCB2JOKuW5zFr/QK+6PKp3Dk+L2+RuJlin71
2+ZlCRwxMgKPbXv0Jn4lAGY+am2J7lnkLxhZ1L8S0V0zf36IRqql06q3W6svtehL7n5wEe6r1QL0
BzDgNKrsUg891jf+/uELB4alM0/gXIunUgWyw/S7V2nZLWFBXpDf2+ZPVUs9AxtvOKHvLLNKDeq0
iVgZkPz7s4EyEaOWDpnSEW65gl30r4wiqX3TRXv/jkkFzwsID6KSdOkQSDcxfXqab8O5v45Ldkfe
wnIxxY9J5dm+0VcyJzHwcIEqGYPAYeLfVS0iGntI1MmJHR19ZYz3KhVPwMnOEObsgMqBHbli9iK6
yejR/7JLGRjHisaRjyl+HkfB3ht9O1mAzI7TeQv9nztf3C5RytiRlrGvhqle4w1YJruY+ZpJgvVL
mm89wHAkpYQmeWGHLjOn/JORq34w70RmNcB7GASZ+KLufqNRtI/Axdh0QpesTSiZC8XNEJxmjp/z
mZuklqtLARIe0pxaF8zlhOLhLmTjUqhVebR0vNPARZDrXycABnkzcBRMLHsgaxEqyBEl7KpqcHQz
+iJkiRPviMyruVXgomM8e0QkRHPVLOfaTKcWPdRlgUTnm+IrjYebheZSlp+9SWoYfFSjpTv/yDun
iQ85JTA7vkaRT+CY+yvpIGkkAu+6HxAPjtksQrP7N5wwkYxst9J3q3G0FDalcLup1gfpnivLUXdC
0U5NPKyLSW+VGOgWSC1R62fInikYzWAYWBsvMz7ZYbtxWrX73Aeu4wJSR1ING09rScQldrFTQdqZ
Ee5otfHzyAxAYVcH+ujoX5ACaFVJN6iExWl170sdZVn1/1Yngfj0gsicx0ZD3u1MC3yXHOvg9i26
VzQJ/mOwKesO6kVDqeZEvdlkFNP5fhQ33TCxhFQksD+6pjwM3zZXiHm5DkKZRuu5g1u00D01jF8G
zzIDI53fiFUtG1bCjICno1yIb7RiBTvrn+pspO8GA12IxZTZyoTJ/+YIffJeG0wu45B+vXY1rlhs
vECTKM1AabGkCLozImblW3Hh0Yl9pycuT9avJXydNR1gntKeJ18CeyyE/U6w79rZUHKzl8h7a7Kd
1vrg5tFyp/b/Bw8HuBut3IlYCST6roUJkCi3RI5WzdVVfKEzRutEJl9fowmoAwCKQUJa2ntj7rbK
yYdIWefuqSPlBJqqCYCUnMH2ozPQdBgwAbfkGbge7FrllArWL8yvmOCODt3Iz6grFKMRvwbZ25lw
P36KHlm//wnW6M8MwMJfBYW/1MK9c7coiraN9IrJ7jQOzYHJ2JXrgHvHg0gDkia0oRhh3iliSDY+
jnXT1qo0TJt1eIrNEHlHSl+Uao95/ILMbjaTSt5DcrvBpR0VfZG52pM5HvlslF331qcBLvD/sq97
WV8nCKXQ2l6nozzd1Fi0xxrLmUWRvlT/Spb10yv9lvJ9o6QnMpJm5dzGS07aLoLpr4WNSZbCqnlr
A4QNQ0TG2xwwnhzEci8nv8CI8ODDbQqxP1tQJrQ7lMbgNVjU7JlRRbLlyqfjIVhk0qOSwws3/Pzr
pstwRclJ4AoJAb8P3R3MV3S8f2S44lmBliGsiYsSr+iWTUCOxktSqk52LucWdsv4lenTU9i6G38j
2qAjkE3MJYdxitPB+ERi6Bk13SA8adgdSjMdYsH/e/TEYmKVTTEgfzYoImhIcFKUeaafmCOcPJSI
J4UYWbzaTJkQtnBxE89bD92MOso0+wTFiGRH5tjEDwjJkZA4WOXKJ9uQvPsGvZKOwoGC0AjQmyDc
DgOMzX+L571HJX8eJXa8QGfgTEf0lrVoO7R+cetqHRkEBX16zypb/ITrIMo0JrUEnZwbgVSXb1jz
E6Me0TTETsYvqNtKB6AQBkvgPI0MnjH/fdthDw8Wv4Fy/enRxhvTl6EpwsfbqueEZUuTt+NIqtPK
CnssuxLgBSjeu5i+NBEgZzXRtvYhO9nuUN7oxrxSdv1W3yuHPRsd+QIK0JyZJKv6E0KJwsGLhPHX
OPZyZ/w55W6OSfm5q2f9CU4uUjOpc8gPOOVBecIdKJ5nql1+BBHM7b445RAPaz5AUMMNmb5MP5bI
5NsXeTtFTgBkYqv0gwsPSYa2LOitDjc5zxir91MR4xBMAtyFgT3X4M2RmamO6rruco9ryVDW6T+8
NN/QQGXIZykcQxPQeL6e7cOnzsAAH7HoJgPCVXUddGfjvG42jv99317n8igSHPcPvoZP9VLTYb14
z2TdSJWSmiHUbJW65QLDm34CC4CV9ywFE7qlBBn7ix367v7bpsMOgELlAl2P+AVpudnGbuoCIcbZ
uhOeamf966iANZoN+WyaSsDT6+bYvVzppvsfgv7caEUkbITlcR8LqSDgHaysAbvlaTBxEmjkSh5a
S76mWbJauO8jE7eQZ2BJHRJcJJgq7wbsRxMGNMA43tYQ53AKlTaxhBmIOfGmCDf5SYO+ni/vaLw3
01vKctR6w7zdl/LAKiBRlHyk15e1k1n8esmshEGrJdtXz+eJqBygLr5qPjBpHmmJY/2dS86/wJUP
1Tf1JtzQJjK64milnlwFaFy5srdci8C4U4n+tNZxAV/0rZgkIHFD2V2SLktc28OnedhP6y7aw0aY
P6d+x9Oqyd7n1xWj0fOyEyYVCZXggpfnXpIamS44XoLKAAkZu7OKR9TzelEEAou3hX8L0kuz6/Tk
bnhKlN+QDDBR3LjowjQbeFBicEQTz6EFHgcBCeVhCQl0c0AEB6pY+mQHd4yEIXxddz0UNkLp87iD
oHJsCXKIMmsCh/CNz3Tk1uVEIn5bBdpGidFqy4mFAoGEslwkAn1aigO1zuLuVtcU51VrHnu1PNLt
KO2EauOzYO/2LKllcQK8U8crC+0FbrHzLwxPSOSAOiXCvtfmMNTHEVCE5UetFvA1/WLTHoh6Qwmp
+wlDQsxLzMiMD9yPZsbWvg/JYfneIwVnaBtlWYMXnw1rgJtne47DgKveSCcepJu6i0PVT99NnH0M
BfoJlhMXuJw1J38EJ1wwLxYIqDPV1bSDG8Ywuve+0bhN6D3idmbr7mhEN2BQMFstxjmCqngnySRF
RJ3nHbT3ULm1W3Pu1PAYCuiOZsEdYNw5NnOwyW84rsAFJut/DPpBFzDApCkUtV7QNiQE/lAMNq/I
+BvNHL8vmnh+eyvqxYgZvBUtnv2ggfy5UN9aR/lmFNVFWSrqOk/u6t0nk9/uazTXzwFXTttns53C
Qy0pw01GLSYAJtxdc/U+7pRWP0Gu+KybNxlzYWAXHKvGIMGxm32qyZgZlCDVd54it6ytdU748AXt
VnlvsFJ2VaLXWPj7qUBY3SiB/UMMAgnqI3RwpsaGvtH94FNO07ZW6NVlEk/WuB84pBvo+H4RpTog
8k+AUdRSvbZniFhBwVq1ZWI6NHph9SlwEebiHAx/Io8gkdcUteyTSgwAiHjlhzo+7WNewOKOhKjP
IKRdGjSypYl8t6ddHgNBZDUVdHZtUFHyDBgtMLMkOoxg2CTiKjqQ9z0MI5bc6iWJtF72luQBnQKf
40td9QxKLPE4XBdqyHEQZDF/tQelZ3Q3NQp6IRK8jjJj8vcpijVBK0F/Pg6rMaYr0gU3Q6W7P3lN
WG24fyrNGbsXrHvTiIMR52dRvqZ4nDNcg7IYWCdH067mW+25BfuqSvUWF/H90kvV0OicfGDzTKDF
NKPks3dqGCJpIem69pOMh7KcXQ9r7hKSo25JrlgswjPqWaafeVEaDuK/D5ovLaZftetlq7ZHxPB8
KJSocyOS/8yA9pwmvvORlys5DlV6RWZp5O2S9qXlvTqJkCd4m58zosbijr8uv393iq8WhsCAdyRv
SJxCCh3MWBFTK9zOr12vCKGSYXmV0gKajFBiPfM+njYi4ZVhCkQRfVg/6VdQFRWJ3kFDgNhmleX5
DyQ/NvDpNJg6e/H/pUM/OQP29V4VGYEBGQtxYaTU5fviYN5px8Gr4bSYdf6LUUOitR03DxcewN8x
BjOcHSivghHM1GrbsvaHhWUWnKwznbxX1cgl2Yb6C0KU7fEHmS94biGcOenJttd05dunwKcd9hSk
t7xrOqfsL3sSs5ukifZRzQXPgqbvA7/uX8vORCyzRUuF+0m3j5J8S6zUeO1zUtbBX+/llMOTRCcK
yFB8LGkiOzUW9QFpafPHVhs0o1aZGmf7kLC4ApemOsrzxWfUPfgVjolfY5uhRys/qX2qlp/Ulgga
WZokpamzc1H7uuNezXDUtjOzxED1BkvvRMEhH76eWmXyMziJJhYAEHqOnLZuHjyoTq8zUNh90OUD
ZfSYNtq8egMpIWg6VGGZ+N+NSY3c+dxOHgnq9gk/UZPjruBdMg2Ev3hETDNEOl1vpM6S1eBjPgmE
eGjRAjdV8qdkRxZVYM67guuH/GSZsj+kdadvGNEAxsCiyhELUUmOpqomfeMsrqRkiz5HM0jm1yt/
Ick35PBvEeiThSNAmy/VfF/TZBs86oq3+meMCtyfaN6/Xiy5S2Vctem63oCvLP6E/9BAFDF9zBIJ
9EJuZvpLWjXQTyADO2u7K/d45D9iMMqpZY3e/Ei55RLlGCaAxmqfUt7xJ99M+q8hZLnHoPzFfCx9
kV68CFF2v/fYxH3fbCHyKYkwQ7vcDn/z0S5LB3XPUQe29Uy4hc6Y2kb96O1Uvo0qQOkl7S2Bf6Aq
voFzxFSDbOh3Ua68TliNAu/I3QW/qeUt2u3t8U6Mn4Mg1jfjhU4EQlFFuCP+m3T6XjyVnXTfeV+6
gTybuS3JCgcjwrHPX4NnV5rm5mUqPUnnnhn5eUn7N7h6LGRrVGD8XEo9tGHHvMRaqWPA08cL1p2n
yQlcyQWM14Xq/d+fqtx1/jRMuJEAyTml1Y/LZFe9K0WdHq0sHwXkC9suUXKZHIfQ+/YAVyE9Nj7p
UGfVpaQfyaHUbkyAlsaIHvBPw5VH0vFNC7q+FgFAKv09oRfsQu8SonbtFc5BtMu2lQ6Kpo4kS3YJ
vJmmAasHXNSS4D/eFAFfse5CTf8vx0tz3rbXwBWWYZy1pcPVonrGdIG8huW3/v2d62kegN8+TVyp
JlMhAMafD33Ru8gKhC0NkAhaSwaI66mPpNVRQ9YkQ+PgNET/sI5Ju8HurNqxM8yZtCxuIUaWNp8H
7HpF2u8cwECE4OQPviswlZn4sEGPopI6NR+EWkq77z5pt1B5ZWe9pK+LcdqcCeyZKYvvT4u6sLbn
wcopamFCBn4foIftnlg4E9JYXYeQNUiomXCZ+2SKWNdqVhkL33yXfAwU5rLinqIa+H/BvsEhfvLp
zqllnVKWT1n82/2/h0IytZEUVOy8hA3t7Oh8PdStCsqN8u5GiMFoMUDY09a/7Hmr06Xnu34P9eYt
hkx3Ue67MFzqseaivZSrJM2UnJdfDBmC7RfikVe6LQ5iyBvfDRqB8hUOlSBgoS69+TysW3JS8JBC
95FRfEJe1JcCJfvYXEnoLBA7yusTyKazOOmc3wW7CTPoP97Dan6LqriCireOS74XFP0el3wGaCSG
lumwAdgLhd6rhN/aJdimYQrznE7ET73UGFcc/PfKIgJc7eDq2L9H4LPvieYv3tGt6JNTxLoqRDGW
Cx2PBvSZDE1XFCjDNpczfGpO0O4xluXrX895VTvaZYOZJbV7C9xZ0cVEcwn+WmAOXdlvEFbKyleV
8lwOo3yCNSgwtglchgZ/nYZZ1Jo+0Ofr4uMTpIVLfBBDd/qgdn14vi+LXd3woA9oVj9XkPcX9IXN
nvKNinSS3LBBHSVROILkMM7qvs9Ih1b+UpGzQu4MNAzGdRKeji3Z8AYzqJ1JPTOQ6x+fVpMv/j3g
QrFvRKl0n6RtOnoK5/HNrPYeZsZhPsQjCwBwyLl7PedePX08ejB5RAlSGkrz/Xvh+/MAYdrcI5Rh
3b6cdL+ybAtguUIp8FXY/iAwL5XqXWS/QkwddD3w2k7fSFg4LdtnJjuN/3QZJkIFhXpvuEaz9G8R
wOsAEg/7HHLxmP9hvvG2PXx9rBo0fsZoGGnnmyGMxjJlw1vt+h8c+IVeOae18kNpSpp8VCnkyz9t
rYJyM1iCOpXbTomdO9n9ZqpcCxz5gcBKJ6pHPqWhMr9NmLgCAFlbGLTWEAAZP4yV/EsZtam8sT8R
akmh2mVKeANP2G8b06+Y7mmFhGJxV0R03aYQkYYLRypuceefCvVIUd2Oq9Hgupdr+MSRyqKCVu1B
+N8p7hF0gH7u4QlITqPrxJ1LE3cTkZwpZHwEtoH58IlnTPYI0VCfTPjFNYcPiW6L2iBtbFUF2eZh
2HD+uGOhtmWYQTtLH9Hwl38GFNm7Q0OBeLe5r80jZc/4pGCLRL77dlZInz3CGH0t0ng96ciIYOyI
62Jb3rGMWxwly7N1rY4tl+CSVeEKaZ/sSiOrpNn5jK66X5i/zdLHBDn415+USiaRnWtOywZ1o8uE
pKER89KBKaDFBfVrG/yeDbL38g8BPvKH9bqxKNCjq09fWIUIzVuy5ZqERrT8RQjU7zfmAJ4/30J9
+sYbFouDb/0KWIdOGj3ZJnBcIPg7zNqc+GADnF8vUYeoelSdCLvYit3ZDhCO8y40pv40oSVjncg6
DhFLyYmCdsaaxAb2yQAGMPJEr0UEhbX0lmI/PtpXB5fJ50JjnZT9LypUGyidzHvuFHVwVjurp4uV
TqwZnOzAryI+llZz8hJtawUpiQg78mp1BtZsg/ru6zIrITVrRVrVwM424Xn1iuq05YM0swhVgeRn
WLmHxABkpUNLv/JYdNwbLnwjwqnpllwDFaYWvXw+7EPNr60cQkFDi3uS9usm4bhP5DyXEjKf9e8X
mHJRu1WcXq/xYaQYt2XbhO/RWsX+prz7VsxPnLbvVyfHAusZ649b9knK23EDiGfWC4aZxSdmJvEf
2oBh6iniWYhayMgFU0gYodvoTQq7iKwMD42PD6dDdl+wGKclnO4bzVjskQNHnKXYkhZbPmbpEmr7
LQpuLELrexClz8UNZ9PKO6T17knYLVxacxbG2H+y+GpCOFtIDrEafMV4mwYd23B7yGx9GhSBLvLp
p5oHHfp92bBU9y1ZwveEIuxfUspoYw8lUuGrDvQOER3gKZvAI+QoVs90jBNUgXqZGhrecmk/1ktf
dchptNc58Urioe7AE4wAeBRj38kkNfG1SK29WPmDk7evkYh/ySX+t8IqkdqIcdTGTXOxHm7K8K/1
M13AlCJAykauoWL4qwsoWrQ4lQXZQ205k0U/GQ7/OX1Kh7KWtgCLjusKxmAqvflYmw/S/7jgCojA
/cgDh5uYFT8NcrU43Lf20mp4FsYraZ2Ynn1B5g9o8Xkff508CM9LGZUmgOlQ6D7xCa7o/7oxP5uq
q5zjqMW+EClAfkTBR4VilFA89NmCmIi9D5c1AulER9tY3+6zh+PhzRBZam30780VlpiFOEIaG0Qc
j0xrYcFgZqaixFInq6p9wQNkrEzWKCoCTGJ0wtJ/pq++l7n84e4WeTHAuGKnoJ3UVdDuUUgu1dhq
kqNXhJXfhNf9vuagQ7VWJEVYPCSmkTUX8XlquswaoqoJOJjSUXkwwNhAh+sK7VVPT7/J6F25U8YJ
lIEbSmfpuEb3v7yorrKwZdVW+XfmmyRHExNU/3tuDE0O4G3rGlt01++uGv2sQOE4wDQ4+M6S2knG
7BQvMj306V64hdL6LR+qaD1SfFrXpIqQisFQuS2dnDxQ6SazbRkzLtgw7QIZX4PtyTggO/w/NxtH
WT59GeR18TaYyQ1F9ll+rH0UJlCE8PxxbnJgL9ENTcTMFg2rBBmY+V5ycpvLSCsQOBOPLojuJzQ+
qmAVZM3FiOigLBlBPa7XvVtnEWxUf0dZKcmVTBWmTq/Zp+XcjSSGGXBmXM5LdZArJA7YDHnXrSrZ
32PaiyQniyAFjjCk76wiNqkJgiMVPZA5uK2nPxquwnNGwSc1gsYcDlLCOM4eh1keJi/1WGRTKe9U
gh0L60ylIREeaTVVJMU1vd92Rgupf4e2LvSmdcK2KL/0Eu/6fy+sIhj1zhq0kUA5aMTjkcH0KnSz
ZmeB6sN/7s+jYJyrUKVktYuQ4SuzaDk/bqwgcScnAsBHHhszBNF/+sTkqRpoTli3zEPZ67ljMnAn
UoL8UrEjFKXxqRCRo6xdo+q83XsmvCQUrn6XpzR5t8SUXtaq5bVaowoIvQ+ETxVJq9CrGtN4Wlsb
N+4d/PUHTK7wI5F351ca+BnNl9dvMywDb+DKsLbUnlSvTqg1kklq3DbHxwh0WoeCORFCbwkgff0F
PYgNxQJUU9I07Oa2REboV6H/RzSJ3fRPTKGoWCVqlGjJ7cawIClVv+BxatE7V9HQAzP0IWEVswXY
Z3IucwERb4dfX4vYz0OPPubo93LoLhFFC3LXmQMvGB+29qZ6g6rD02GjKrsx8u0ZNVxsXWKXo1B/
FPgoyPFHI1xhDv8PatgGMjM0/BmBPUwqSJ6LjUk/kF54R/5qp3QPbo9ClKGBnEEDsbOQQ42A3kcK
tKB32yFBsz/WQy8HWbeVgIxXdYK5FRw8/qcdSNJGm5sefd6Br8YyHOCDxX5cTJopB+4NHEYkZMvm
F1QtIWFRbJHPgqdNRGEFM5oRnS9U9VB7WP0q5w10/jNIeQRXUpmF11Kx6llH+9QKLf7w/98uVKNP
MX9fmjo3Ou68TLBu00ASgOnMwq+C/iVQQN0Hu1z/wAUM3d5JldBcJzHyVXjacDyzHuuTBwiX3Va1
kbDr/L6ARFEhFqsLoApsFQaNoWts/vmSeB0zUwNrKkTTk2dOHV7sWSKuQtMpGGBLYywTFWABwOe8
1eQkiwhQhUXQLZvi4Hmr8vY3pb5dP/wMq3IInoT0a+EmsavpWnMTC940DkLkKl8LOhOMhGt7SpRH
M0VbnKCbDcgxn3crPMqSDq95ZLtvB9a2ssnDKx29N0odC2wG3y8t5fRjo/+mFIQ3x773fuzfpM1B
eS5Ga47vN0COtzwZh6aPAHUAWhMCZG2SqnPLz1LXIOV/4MnyhKujNv+ClG/TAO1XF+3iESnf7exS
azYqDhZQUWAJVxnKiz/6n04z/cONZLX6jvTM05qGLUjlxTEEySOjP/L4Hfl5WJgjNKdODbtTDsu3
xsSrSHOKAEXhH1bfgzScLSGrIwME949VjduXegq3TUAYSOERxFVPyBv70jOL9dJlXkjRLRoK9ehh
MZ+HkAt3xY/xINzljqP7Jwh9Pcl+828WapQ8k1kplzM5Wu5RGhB2WTrfIEEFzjEtUKG+n6uTW667
CZtC9mHe24SvUiZsUrM3FFvX/0djEDcssDLk0bE/ZIQdKx0JYjQxyWgX70W9XoGrL7c+HfYmLll0
HhlOQ3JCqTl0MOiBNXKlkOdQLkF600/lS+fjgyfopHmB3FZEORQFPZh/WBBnU5fCKsiX6zqttrlH
6DzgICxfOOtsSA56SahXWl4Rq1baEt6U11Ogsc96asIX8QF6ODG0oT+o6jI0fWMzwhPKesxd1sjn
iEIAorq0ZA5xlS3T49wMbTC1lya8ws75BwnUJqDo3H7d6rRYeLVGsMl5Ze23MCkhyUo/pUk3C7cY
SqtcpwRjz/wDwxucA6IB7bzEFoWKSZuy2tRbjGYcW1zFu1P63okrqKvUB3nE301Rd3vLeabFjMgz
pkpB8T34N35wwkGzgA/xTWaITLymKNBa2++kt4A0r+1bGUJK/5Z606ZvhQpGF5o1HPMnqUgIPKNO
zpJMqncQBAXxZdYHScKlTAB9pTP7P0tSMErf0uar5cEE3oESxFvKMi1GzkNiLhTawt0rVKCv6bms
4h9A5JnIFxj6pumlnP3VlAhOT0Ip891nmHVjQ3mfIaGhuoElALJOdFsMyXWBAjhVreYDUVBZ4JXF
+ZdAZNvVqK/cXrj65zGQ+0iAO5TBfHbIQfrQv8A6YKvt4s90cQ6TcCPkSh8VdkYNMToguExrxbI3
ZkGjIiITp5R4qvqVvmzIJfNkJ7F8n5zoDZKXe30Zwfex4pkky3eyvxegKoF/mNN3GxumMkIxipFv
pah84Aq3X/W5vc1CmNTD53IwAAYueVDqWuKWjj8o6YCpg1uIiLbxg85vonCHmuj3/5pOO6RmNwdb
nTcZC92oIoe/fkoxHm9Qx4VqTg5C/B3cSLb4ODE4HOaSPMpUds3FuMRsQhmBkO70yKBkiXptHZSw
zZ+SUNoY1x6OK3LRHJkKODsVU+bB+KN8WurG4qNIDiLCv39+ubQc9ZsFF3mdPZ33+8meafu+Ziyi
QTl8991ax7aZ16UAQZkld545hazdbZpKbqwioJfPU/GVAfRDGgf8KKhZ16+HHtsJcxberWyzvnza
ThOaTAcjIIGDOfPOPoovhE8Ex3iIY2EDiha1EGHSNuW/8/7bGRNSrNSaV5GsGjXtTKiSbnm1IgIl
bboW/fG87xaaus/N9mWReD9JwIfTiMtGRO5n/co8M0V9HD9MJoy4yqgZJUGehZO3epZ83eGLl227
UsMbKvjjbG94cEamyCs+4sUE7nxGxMEzPPQWEnZwDI8TLe6FBe6coYWZy/UrFhSL6oVlmNvrm7rT
1+QMegBQidzI9wvL+J8wKCzdKWmYdbEmdNd9shiHvc46L8BpTDKHYAGWgfyopFb5XcWDeVJxGti8
he2YFwJtk1yjitmyHgTq1iaMonytyUAq9TG8xk3KO/b45mo8gtTZsrVC1dSTrfmRyCgxFWTGRPiF
ryIoDmNVCn7OC3PTkBFhEyvJfo5go3cRCsMun6+y4T/gejtTNsI5/LFFa/6XfgaaqnQr4C1nHBUK
bQCKRye9dAo3B+VLJcVJ80zTRx3QBduEzEsikDcmGfJ2LDIq0qN5WkCZ6x4VVl79Da48maAc2R0D
kYks3XG3DzBPx41s6C9Zgya7GZheva2qL0jx4F4ud66x9oKyxKAwRRTzXCywPldNybQUrBOr9oT/
wrNl18mMKkPFOkoQnsUpRkceKUlJfF8in15BnCZFPI1dDEcABFNj6/PaJvuBzYIR4F17wtCBOPFb
jApqGh/uSryqCbckJph2HhdOy35BjI79fdnuKD90fetLBRriXN3BlytXe4w7QIZgc6SG6rIC6owg
FuVbjU5MOOkf31EkcuTUiDTJ7PyS2hI2Bb07Opw5RuMIOO3Gtm87Z4BEROLvbwuMO8hrorIHH0C1
p01gO4D+BT2rgFyBKWFN4ulT6jkGS4TNcrLR+cRImJAbEgqxLTYzk6qDvzvun/aPzw5ZNkM4lVE0
SEIyLZVOBlGSh7o6/gmAaQp4RvQYpG3L1mCMq03lR9OdZst96hJYM94uDKXr7wvUXsIJsM0HxjMF
u8If2zHWEKWtvYpOdaeoMLfWJbxhN4GcN0b05qMT8VBWQEy1pCrlfEp6qj9NkR9ZfJsOrNKpf/EJ
/Z37TCbkSlGb2RgqAvn/BExuBIGIC4BRMcLR/uh4IAM0iq1GNs+GySoAehVVgCgYgTNRTdTLMOFc
aMOXymHrV1kck57YZCIdQzypxJoqbi7h4FSGg7rMR8fuxiYoZnsOA1SVYh+NvoFtMpgVblmEodq1
D37pm/wbZW+X+44n2vSUZEE+cBwMi7aHUSDaGBuaKmKfq8XVGiwwxvYfvZ5MvyFU9+6gouWoq26F
Gz7ANMHtDz+n8htd3kgyIRZB5V4skFoJiOvH9eONrvGhZsVhq3pc52JzRrkyI75Pj0jvoyDeRP3O
Uhm2iOOU6sIB7aZXf16qO7lBBjEWNL2kSjWrtITMvp/6ZlkiAIeaGx6Lyco4M5tqP0cnD7cOOskh
TfZJjVmW6zEZWqOjaG7bWE3GS8r0yQTpzTncIbKNy+W7Kop9Ylr3ZWeujRGjeUApvadXPkEyR8r9
M5KYLOhDdFFX/9DUG4UsTvVTUw652vcpYpyYglgsQAlucsLTpQSfnViNoTDpbkOKSXCa+Bg19j/r
TWCZ/L3dkmXi8Rt2VLsK1SH3gQW11iKvMf2FsSV2z4+YFBHNOH2OzJ1QhMhFDIHEprFwphPkdRaX
n8kkObxTNEkeprxGRB7rWdUS0mSMLuvMECn/VHaoemSDul0UB3+CpkhMaZixjaF96Fma1j+GCFf/
/MCE6/g62SpvqFYtRFgfO2tr8Hsomn7ZDPqOTGeHaGp5eaLnU//hDwhg1EPL3cj6UDOBRDLE2vGR
OmlY8fPBy7xWjYgraxKe8HlkzeB7KSvpYmpNmuM9mmbW0iov9PpIz/im4AAMGriOIw+PyEzYsYh/
MiHOosrtG46kT4eYVTsMQQQBDRPgzej3SI7ykhfj0oMj642boEMONwaqVW7FsaS/nwceixWKZprt
oFVtrbjkbcBFf3zljTPHhH1vJcbiA770fvk9/unQ1Jy0lfe9WjJNcpmb/13VsWCE1e7hLigklfmP
W3yOXGme0T0oBYuU3cKqo6vWsGGA/xJPW1stHvQcAj0UbkLMvvfkCkppdQOOzLj+d5h9JAf0DGGY
SHTre6mI8213ZGkFUDb6CxUE37x4aBPv72XvQn3SqMvQEEqoq9pTCxV6xsbIOvlTXnF10GmrrhP/
VDGcjPpkVTNOOOYvznbDiMXGxWAF2qF6nV71sP35hC0CJqQ5Qsf2Sml0xg8h7FkOEXFtvVe829BX
lp+FOrda6p3u0JGK8RSyBFNKzWVJKlDRdPdnUosadapBsqajh6VDTawoYgb46FXEqxKSznTsuC3J
jCmgq1g+PPMyV29/LrgmQW40uJhYjyl+0io3hYGndCOB27IVbIibbCv8Ykf+tQ3uOCn+YIJWMvqL
bqIJSVKp/x5NO4H0rC/epQoSreKuOBxCl+DGBf4S3ZGoFwTSiTvtrAvaP4QVpGMUx38GO2UDZD+6
LGYO4SXMucC8cs2sLu/8Fte6LGK4d/Nd1WBr3D/qjXbu9uw1FQZeR7t3yuR4irhUNTIAbFxAWXme
SdfK+kqT8v8yCE9hQ8+GHH63fWoMTOYqlnVZGS/JxZehOw6vSOaM0JK76z82OJLIUX77zy/VUsyV
gJd6h2QS0ebIw7/8p1WspKIuCZC4PHeubXLcXDi/XBnZSVKNlxO71vOo5m+I6BiYvvX/mnxcb4rg
2lNJTYMjHYTCimdSwTc7xn5wKp8bN774Pur7VFXHHX+jq72kPyGePOZGyf+q9OQZbiAqNK5el0zS
ulT8N87G4e0dW+rW+2ONZSfYrx8nrJGxbDKqASvf7LoIcxK37EnMcWEHiv1qe7074A+u5I58B5WN
1F5/6jNRhRihbJSyFYxO1X04wEtAw6a1NmTkD4I+fVDxQSqT+Bi7eC2f2nqrFsYagDjiX3TyReYs
e0mlyO5pDgGYILHgIeirhQQt8k+IqK/gH5+one+Zbo9i6EKozLCQX4tQ9aaqmX2Dyb3XBWKOnmLn
AFpyTc3Ujqf71TCTsInxDg8hJmAAbkf9UCx71bTMGVxY9jXwA+9ggBskBL6d7/oh/JFmQ+hk3Pox
h/UoP24vUb5BXHucg+eAeoXEmyJsNLIRyZh0rqpgeMKGbAoLnvDnuPcetR/ixERjmag4zQOn3Q3R
heh+n2aJ4yiZXTcjK82pR66gKBxexP6lUCljIeIDHTryfuUXQwnLP1ZrakfBDYbr4Gx+TbxvtFr+
TX+5nq6AQLje6XKh96XBO06OFD8BzYxVRQO7VC2WjP0VH5VdwJQZzwTYbi9b27xE2mGiELBfwgQx
1Dk+PMQBYsyZy2dmwX0OQlQ3bQRVGdhB5kcPD4K6zsM+YdDcr8qmcDc17ETlPfHpQraLH++hbPY1
/ZW6cbpsO06CwuHzdsNkylkX2ITT8MGSOnEDh8mdh4cjOvBpNVNPNTC9MImJQ4b3DjYk604P/+NQ
nPaxRmhLW1cuplSpK199fUtEZzTRsqVKN9Ic0xw2otRYuBZONzyRBxL1ScrrxunzFwe5fh48yRIb
xuCiClUmhf2lFZqErDer3/lBwbjfvSNxjp+yMVw0k2GzhtZs546uqGyfJ0WnArbK3Nv7BJ9m0Iy5
timy7TB4AM+En1bYJsUBwbhZiH6Nl5s2uUTBet1yBHFZgHRSEH7f+5jNFUzMfTzGrkHbvjUseDPq
u4fspdk0wazSAgaFYRBSpY26NYfv9INQ8FmlYt9/dtjZj7SndlFAPLYA/9yUx59DFjQhwhuvp7C7
s6UWRc1Bk20ec0e156p+Tg7FTgS9fwhsYSIZXnkjMUiTiYrn8q657m7pLCfXTTGM+c4wiUWicT5o
t2w4taWb6uH54LCNHYCB7mNyxCoBhd3uS3V0TJxlqzecGZj296Kq2UbOu+NEnZk8+zizyy5xTtVa
tDPK3HpRxa1yozZqlTI8KdkcwxlDk+bhMRrQPQrdglWDCFSbyFAzJDtDxSEPbwiRXfdkDteVjNmk
x1PgeqigwMQjowNaNNfrGuS0IKckO/TpN5t3RMxfoFxgUnDuIKJs5noRrCoQKasztTvH0ntoMizC
q92XVoP0YuY0RVMOi2Kx4WNhIFjqpDDp40JN/iK6DBnn2pO+4l/mxzNWzGJ80q7JowGncO8zCSdD
bqZfhEjlSx3TG3QG0o99rYlsAAar7Fx1Eer6slbK0peIZBJYvHZ+AwtqAvoG9BcKA7a8hMb7RblX
//oQLnlVCQ99jHDTUzR1eqVysfdk/IrtVyHTFwL4ee/wWmuEVXuHKwDoxkP63x0LVdMgXPd8tgGt
XLeDtmmSs+7n197tQq4iCvEd9FEEBEMe6aC5DTdj/HhlSi5gZ2J7JbHuoRDFUC1QAgP6CcwAA1dD
9adD/0OHDrwP+EQWmhL9FNsgLRQXCj1OqRM68P+9XQ0DIlhMS3//4utnyYUGowyD7LK2aeeWTMrM
LbtX7kWXF8lhBIztYdaPGEPxUctmwVcNMoOVh5I9gDA2QxjZNi7ThqTGtsGRiQRooZz5avr7v9gX
JJz9WDoceb3ySDsNEDi1OHUcO7B1xsimkcDGZhIs7W+iP8IFlCOz8/ijvQfYgKrIKP13glIbOlFm
YWAGT2u/7A2WQ85gUFkgoH4fAEhkczvNGN19nzXrMdT12fKzymm3pFaX/Z9kDNfmPXTU2DkbhYOn
nkKmtZPEGnMKRf0YhS6y8qYIPIrRgy/acx8sCTxgwndoDO768OVUQCZiHkkRE/Yb9mz+6zG9OoXF
xEtCbgz7sGdRmTZgTsVlC47M6jFCuxvr0HPzBWpYSZPx7zNpiM/e7a/DHuxsMU7a+dheoUNVzM9m
P33zhdp8m8SnRAJ0u/e+JhJR/ZQ0EiDYVGrYUZkDpd1vFBOD2pIYrexIkF749tIKiHYsc2nSyRDf
Ut0dvD3brQMU/alwxJoAEUBI2hO1jxLsz3w0VlJb7gXusGyenfoJJj8l0fZx2a4OMzCcJ/Z7EVHB
Gh5SnsCHfnqixE8eGDqoUysVDKN6X8K6cNDfKz/+qoutT8GZMj2IcM6XkOVylEsv0gs0V26AtXFI
uNMIEIhINd7qhjMK6PpX3Doe5UMB++84DghkKcpTbi8WgumuZExgLuE107G9O74lCln8IqcQNjSN
+U4UOcEWhqnL3qqfAFjBza+PE1nkNkpTm/t5Y8qeHWyDtjER0136SVZAPw4evz3tIOhIc4VrvA+H
Tx7IDLJAqebpqQLAPxTl4ehBpn0Hw1/B2fw090YeG5xYtdu2OIuL6SZUJYmv9dqNw0VvR2Wo0Kl7
0SsCSzBILTbomnmaV1Y8wqskTNRvJdn10iLXutnMMzROGHn1MlT0tVukQaWOs2dTEhp9/+LPTuzc
G61u/shFkTc3eule6GCr9jiKH974+8pqIopNrgAf+8c6vS9TWOw/7+WBEbMwwYiniDPuHCtjZXp6
yM1+hqilFluop/bxtw2hcM9BSwdQtmENVAHL7P0+2eyNE+Ep7Nid9LS5IQfXas0dZTxg4QNOeqB2
BR38KGLkz7dxg+SrxxuYPtNjxJ/J5176rjqRfyBRB82o+L+ud4Dloqltq658RyvRfC54xqjgBwve
kZ4xcpe+tM3R24d3iB1JEc+u09r09LTqbzD6c0w5a9ufLfRnNnMtobINNHi2CpirnFN2AXpujOBj
jOc8nr26YI6XSaJo6w7esBNYhI8Wzaf38o83cLDAlGWUkMbXHBXEQqEdgAEQoJuzZilesCC7suPQ
nCf2US3hRg4UW8kOjHvaFtBxf7EIE96/ywP1m1/2kP04oqDTSp89AJ+wELmsvXm83kNGJ1CrRcFj
q97/QXD9UDYPw92AGqoA1Y9yKRAszkyXY/J0z7TNPbCyGKYmb0s30qKVCzoLrOq9BahdQNeIDLa9
twLM9aYpEJK5pYm6ox/PgqS6XJIzz67A12vlAgtUjXL3L6EEkdE0jpsDLF1WsHjUKuDNUIUYGu5y
wgIuAeytcDN6MtWZXANTal9/loRWk6/pBkM/80YHT8v1GRSAmYCF6UnhvP6eQgi0PT0uXfbX8iKg
cSkdVdBpibcUeR8U7ZKQNZFi39zjJZ70gjn5Tb1wNfPnADtqHwaXp1OqXna1n16cONP5dJmgArOs
27OrIla5A+ulc10aPzYO7zWjNiNecEfwHTuGGm5XgTQoIgdzO4RznAxoYOlTnMB67Qu/4eELz51Y
DriQ+2EWiUG3HTg0h9a4Ea3w6GCNe2ZylF2G1f1UpiHn8b1ABBUnKodi6zP3V7IraM+xh6IP6/vI
9b2G9nLInmmQcqFsBQCJuhLFGK+k9YguRmscccZ/UXs6l4umiUDD0uPnrr7n4vq7Psbv0wWJwXTO
PkC4sNwpyeylDTBtPBnYT6sYH5PnnSoVAZ58ZGPpIJKG3KdZgDcTd9iKJljmyOnZItmvT84wWY2T
73O30uKCQjUs8omPGDyIHQJCnlHAlQleg5b5Lo4DDmLLPlPxFAIOftR/aC5vmbISNrfoUoKOrKbl
tmutXhBK1mUD2JXEkeg1fyLmOLr+mx+9TA7vkWq0zG0wII7tj7UcwDkyiuiTLS1Iolm7K1th5gy7
xMhZArRxZbPEjsVXt2BjpI4oWvXcQVEzhLr48lD5FXefQWVHdDnsilKIfLMmXRMdOLsNY6dZwkms
9f2Ub5XSjmkuSym8GbIIMivXsy2zmYtPkI/kCaTSyKlNpfAtwCS0yrXv3GpxIIXMOSQEqqllioMT
dNs0+AupmrvFdpLxmTM3P3Gyhsv5BkaAyyR4fxYjDnhDs8Ee3NqstzqGCA3XxGeCH/1sVGTap4wk
kqKwSnUqmMNc0ABOpENL2bctJRdGrJU6ViZjl6L/V2PCsDviQ4na1yIMTgWK+NqmZmwdWhN+zwCF
5gp7W6x61k6wLBA4mrmbAyOGeIw1m/EAUUJOlaRkqmJSuxHtZdkkBj2JwrHmV2Y3Uwxfu1d4kmW1
RNg4I0DuOSbNN26Tr2yHR43zUNT8DSCdUdZN6l2F0hBohqjulfP/QQ/6QBkf4cys4qjXHm+scCzt
9o0n0h7wdp+NDO27zjQlcvsirvK5sCzOJpWLWNQGZbfWcNCQRvmaAd+dxmYDG51MJR1WtdITaCPi
bRZX36Q72vWouO+pSIjN9yXGCnkzW3YUn3+JoY8ZjJoieP862QRHBUGsHqktfbykpQWULUywnpN/
6jCadKdJNlRQP5DYzoGbIybhGpW1WIU3QbJvAj9hNtTFmqifeQ1tPgjiQp5LleT289atgjzMqum+
CfBsay3tdHGkavC07SPJkRrRQoSULDLfKRacneKssxEHU76I2C4hB4rrO/2f6yd2wDVQJuUYyeXc
SYAtfp9W1vj0wTdJ9HfAjYbTSOgA6Ib07vgcWOGZ1MKkmGwh7H+tmH+gTXuOQwqW0SOLYqVRQrcY
OBO5OkdTRtvhQHY6acogHZIAE8B5hugFSWMyDZkd+bSCqLBFTLB9nO5vY+pJNK4theytl3jhrFn4
HRr8ggpHY9PDNG22PmGsh506FOAOjzaCs8Vxi3KIAiXHj5bE2qDtXnm39Ogt/+VVpf4xJcqfqy5u
wyKy7jq5c7ED40ad9Mkzl/zhtkA2KRQ1/42s54KqNkKm18r1MqR5x889vip2tz/34llUcnmuud+R
EmdHO+8khE0Z2imM2ulkJNupgMKdl57DatYYaOBknB9GPRBSTs4RvF1mzzbzKgW4LsHSMncNcvbw
b9Agj8Lh+8dM7gy1Up6soeWQ7+JBt0ilCdYTVNTh6QPaZxs1wEy041nkvAD2aRRUOQntWQ8G3BiW
0KiueyFDWjr7LjA6zMjYuI05uc4+cgcp96vwHzP566l28o01BtHE2EUJoWNIG5yQhOd3FxRqpAKj
KQCfSJmurHL7jKKifHMlK/LVSNKMZQFAXHsNta4Q6PkjO5KebUgwFA7lxWekUgtMKZVgpuphqLV6
AcTVxBWx4cGvdA05IgM7G7CfVmaE9zqTwKXLN63/7f2Ka7pOarUOtyU5oyYHozNlU8fudetN3164
43F6ZSTD16K9mO+niAdGemzywmYNWxs2WK+adMTj5GBBF/hzqY7bthHxMteEV+xvgMbiG4lL2sZy
IAI1Zr2HtyZCPsux3xrnDCDbXJ7jmJNKP9rPZfXCqYLkkJDLEVyiat2FHLq119vzZzMKYVO8JnFr
xELyuVBYSqq6oir+m9GNaEocNRFxCDpIVyazB0GXn+6ZniEag3FuBggQWwIdinc6eOcsjfaU510B
V2MXqcJP0SJFHouN5jnxIVUTATEq2fyFsUPkomnBWVejIWV91hbK6qeHEAZinPK69f0aYNX3F+1E
1cKA6Bi/6W97ZO2K4VTI8twbSl4WVSnddi5nncKoNDWkT0VkE7Hf3xtKzCTJbY/TMTx688EL/c7C
+Qq5dkYo2FMvEaHt6bGT0nuX1rZses5ngNh6m/OcSKDuyiQY/zecI6Txk8JAy18cxO5oXB+gJfml
FfqsjzZhQMQhHZMrnjdzkcA7uwon13xPBvtH25Mw8EnyhqFulgLNTUp3RYyoK7kAVubkue35fExv
8DvYhPkHS057PH9gAGhA00TtL9Q0A01+zU6dwq52ENTiAn+Ugq+2T7GLftOmpkBeLKtpRlA9hM/S
wKCrdhLuMar1Dkbw/aeHJnMYnGMFcmMYSFFixgHUJgBawnd6Q3xREsbvxoQ0k7ipFy0QIabXI+92
WaluXkl6KY3n+2SY3zXxx6bqdQK2FL0+JiaCc+rdRx5ftun78fhY/uU/oRY2QsDtcPYv6lLTiR6m
wDf3zija4Irqpv2P6iFlUZwRh7m+RNS0LShZP44ZI+QGyrYmAvY9hhWx1jsUo5r6D8UyZjw3DUIj
gWGA/AWzP9QgIYj4V4Ub0qEbdF3Tl9xR+A1NJNPzqTbEZTczxpN4e7v6az14BwD+evBuJ5tvX3U2
3ADt0VKfgdv3HhzzPh+It09KYw1e036wm5irhG0EjR8bjgcuPeI9xSmMhWHzQ20s14agQSNNLgnj
D894k0Qb6OzFqu1EuuH8QC5OjXATvoDt8IoKWZ3UVyURcSxZra4hq2M5hcHyDAJ9+/jwiDnro86b
la26Np5v69TjK4rq4fdWlXlqMWo3SYUSeUBsz9/Y9u8gS/GQPnUuF8NwZVLDNAau/EjH0k+UGlcA
eLww0t/dcds3TdA3zlcgBVNMlFXMxcgPuzFcFZDjqSiZ862LFdc/eEw18qJHm1c3TScZ9VNY2esN
u3xLMBP4Vg9fi5jZnJ9suOhqkW0wK8Q7o0hi1TI7WfPGapDx+ZWL0SVt6lyy1z2Ln8jcaQGgtb3v
e5JGbcK79I9W8H3Bp8JG1OUBYAv9K47ZSOURNQCj6P/jgOV5j5Z5LflW7RysJFdCYJgiBnh4Y7R+
2qqUFPcTIHUQwjQPB2p25iu9QausRqPVNlnNcu+/ZbA9WKDA4Gg3gQFNwa1GphLWUWmRRsUQkXur
Edt3IXdQgOirZSz+foC+sBKOApg2t+MXPtv7zK/usYq8nCYh9ZE9HfSoUaObJQjJGNbfYKrAu6O9
4rf8gE1S1Jl9r/wuAk3YQJsFs0kf0/z+VrPP/QToMsxcaY+VteBRK5i2Y2CZja9xzOWyTMirMMbu
9zbyNs7O0HrEOyYEzzUMutz+TiuVCSrLsY7l5MJO5G0OM2qL/yKoFE0xiJkjKcsqzqFgBOc1/JWb
iLx1+D6IjB+q+KF3LaUA8HtE87JhoccNQCG0NAL1bIvJ9n/t72JrxkowMQXAwL0UuViufxpcws6w
XlbJERs52LtRKACSdYQfPKRJ41iSzfJaKLnt1xuhssEbH1m7KqcUNWrXhthkIYCS+tUEaDWXPuMd
YXQs5/1QJugBqt+7lxalVase6H9z8yuv45T22eAzn9S3SOqGV9bzbn0UYZO18yeWte5rx1zyXTHV
PfIen1yNsWUW8toVFJPxYLoX+Dnt20ROenOB4jaYiwGigQRnqzK8F6Y5GGZLU6FgSeBEcMM54ZPk
1NKLit8WxPpeXTToXqLH0WOftSpv+NSFMBO/yyj5lqXUqBJxquWu131tYJY3sUHzvZo4lJ275Hbx
NM0u20bHEy+lzFnUinqcHKqFvVd3iiCsxVoRVlICZ6Ap2R4bUZMxUVXRJgw6XQ3SLMbMlRwDNfRk
FEu9pYHHA63niR0GVbsdFN60sapF5CrUGYAyXjYv21cAYhTwCAx2T5M484nc7oF6Ouq/CH5nOeeA
Ua0zCAARFuLNHeVg6KGHatotiNX/hHUEt10b9fuJzm3R9TFfV7kf8kIYEG++aBjXgoF7ze/Iq+ni
glvJQLKJM/ljY/q1YkkSSyRbLjReZyW1DZkHme11OS35Ha0sN/142jIr+o2A9wFg+KpC6zzEV2J5
iSfleoxE62mHRBm2sQrVxlIYJSe46pEbilJXW+9WomoSnWXm/Sx9JEx720HJRqM/DLPljAHvU9+R
v2skoX+BThUc91D8a6L/KssumFhwV1sMVKx9fscYNELzCsU55Sc6nIZtiI4YqriaRrkfSoMsOHiv
88us2wylZvDYbNNJ8NH9puJqIpn8YBRfdBxSdpGQKbVfCdre8XxVqMwhgbKR72VwunNUXvLp+DfW
OB4mGXaPYir2lXrGRfHFEI3D+xYWpl+lfOSphHLIPZV6HlRg0kTYFIpsiHo6LvNQhCNBTXoEjdR4
ODDMxoD8NT4pVMlQrZzSTHIiwunCh5zmAk4lT9M4GuBVrh4voSAik5Sb5PlL8fgNF7F+SiVjU8ma
8FDaf9CW2YEaoR5IpUdthIyFSxd+WCr91bXA24F0yz/Zpw2rj2OCYz++WfRnV1H6NFUtiC7DLt2L
9SB9FBTYB+HfZDcAdWSDflWJyssO1GN/Sb8gZZogPbEYoDHiPwz/L/VI7sluP5xGX6+iU5ikPJoP
gZAuY3SaID1029+beeoVDUPsVWzJNDFzm7jgh96muIIwrEjarkSds64ZFCm43KgKTEcYKNquMUKy
jmPMkFNUAM3+tXr2h93l7hN6L7yUapYuKh0PyIPDc5/udnQQKFU77FYF/XTkhkQYVsC8ZJ86Wti3
xzziSYe+Z+vwuutXvdZtK9JIT/ASmWmETbkoIVUAfWQHoSyc6ctKY2RFlnB81ELtMLoiScpfmoDU
p7bcZsRs/2wuc3BsHU8AxHPP8KyNcGjMTOAZ3lj16QRqBRZWpFdkp60Ep/9lalmo+z/pGZxVuKyS
138HO4xXa5vsK1UUW+mPcIcVrj70FUAWczz1OKnNHcgpsFfO1iBIMJfNZuCgXx1MOa0SoJPJINzT
GK9b/GrV6GIaT3a9MyfwdTzuZDuDjC/TRgvUnSR3rUafYWkAPvROKONXWAe3MpjG3z4N7NYdV6bq
DO1DI0XvKM6tNUcbNdO52m81KFnsb45hm3XIcV+LR8jQU5gyp8Ep6LnduzE+laruFRKioY9W5A9c
DBJlogkexI0cvoiTPOQtHvzGQ8UPoKJ78MUPpYgIvl4pCQZv5JI8rDpS8TwdC5esm2/1UtoC76aC
8POpQDeJzENX/K4LEltlqA3MKjMYbO8nn5tHX0RdtbWXJrSpSBDWmyAL2BOJijV2KpxE6J2L2yC7
o+6SvKTBp61+TWYaNjOTjtTI8Kaa/gRkkYDGfpUiXAIYEvALLiARdkiL/oHUIpfhrMOS7Uf0UrSt
DWiAh7pEEPISwtiaKf7LWrpavcxZ0tMBek4OUKBrSU1goSGgLsjBgBMvxEXox0QFfF9+p5PhG5KT
EdI0AFV9hrgGbJ6/+b0utLFZ8J8wh62hFqgkoPLEGqDfyb1VSbvfcOnfDi9oz00gzKNsUBBT2wBv
tDagES3hanJxOo6C26rhO8WWuVFt2m2wGoOypqEhK0GrpivkJLSdu+6eqVwpXCioqMbzdTK2VDXs
pfUKY56C0JaYMtgQHC+vv6YCUj1gJe+Q+D+b9iBK50PeVgAVE4111f81qPnuWLI69vo/UHhbIXNb
D6gnq62aQcpaDkoco2cE52Ph8JYrHfUscW/JGoFKj+BuKzJKitQF9oRI3as2To7VCoZM4amKnMA7
4zBilxgX2n2yTBiLdbDTUweQxI4Iub4j3gVqIP1Ag7BiEYzJD0VK4vijB7NcWZWvsPDKKrD23ceX
3ZFVy7bab925NcmpYWYdmP1rHWO76d2pmqBfNWZorGgy3g0pB8kvTV3Lui4vPiBxx2TiMmAZXDwB
xvikdLOYSNYW/eVCQQ7sE/IQu8UCPz5TVANKTSBL0Q/h970LwnkdburxpO/sJkxcZsCiT5W79B0C
oVV7qmvDQ7wexQdmo7ia+MX9lxy9Oo6ENedlzfb2XISJnfjqjXZwH65Z8V327MYD1w5FSYYCcR36
R1DPYm2nwh9zi+4yTL2Rqwj47UaM0xEJiWZ9IHfXWl+zlHVff+pVgvwa1gc+OaONFq6lK0jzcNWj
woeTUef7anWN8iKNmwhS9unZMlSe3rH2jFytGB9VTnH1t2xWKlPzwTMYlCIXHGj5gHPQLu3ZZMPt
iVjm5qOTP7bwgR5jnCejqBlUbkSm8T4AGfFMKHTzNytjT6Sa+mdIsW0iWZ/Y9eEUbeJbe8n7SJAT
zXUglxEQ0d6/KSGXgFuNbg3/dE9Ps63ScPUeVZ06sca2GZXAILh6yh+B5jL/hiPK6Z1iQ3vvotqy
8hgS53UO1BEDNxQlHSajSmeXyWqBYLiCBMymZk8nV/IHsBVmJeXe6MwxxjTZSifzQK2EdbXjyFgg
CKCb+7dtmKfqDLn2i2XStios60Uu10bSr/SfdDLxijniQOj0Apv6CQwAxS+rgjqS6amaK1Jx+83m
zrkhw8s0mzGhV7OFWDARonLkvOWHy+YKSYyzF/iT4jRPDFhHFjCN9OvTpVUs3eQxHSM62ptYJqu1
2SCz4DOmaj4FH2upvVbHeqiKsvOw207S0FDltKLNuOnlwBM3PIh1KreHAWnHLUwAKF93WUMD5wtL
9WK6dhap1zauIkMH9NYAnFtlLWvjWQWLyUdfrClzHEjzzsYQ+egqh/DhBbjrF6+qkTheCtTxLP37
mQJhALLNexr7hWOu8kpavyjhMq8Hs65bbc4mRrfjQdrlJDTxbUt7cenoagxYPXJUDh4bJPH5GCEb
w5pk/w9ay++MptwD1iB2EwXYAJx+cXAZc9KPaikJ+f3XXNRc3y1PTnfHSEWm6w2U7AsWBeCWO8op
L/5cLYFp3ilnRMjj93T6UNiUQxs3HcPHRjtVuPCuCKOlD9fpXzWZSJViejcu+YMbfPdVUxPwio6j
43kkyaQJ7JKK5eBNfCdMp9rzLp2AEoCTyq75pJGEsmmr1EIdJ2g0BEg9R/41PL901KQY4cuxbF26
umkpRCvmNWF3kpw2XAM2Qre/dbMeNgjXyOteiALJEi/OqT2H7xJkIvpSzFBfyue69V7Fd4WR5Wej
4u2eTzAUdzmICLzl/AZGc7VZV6aath14XWcSU3VtZNe342q0LznoEF0JwfIjY59HtNepOewnM/dX
/mSRhTOPHD5BM+YxfymdkLNc537xv5GWq1NQJCr1wZwipcdTY08GaacP0NBGx/IsfbbjIStkSSiH
A8UjrfqNMvhV3dVlfSyzm0zTgpPAZZrVr9gbfcwEqmYTe/nRXPPsDY3CLJPq6UXaeiY49ueNo5Lw
sZeE7soorMQALzUrh74N6qcXW4pYM9mCYg97ijirdzzcmSqlfeZuPohMWl1iDi1z2eM+qovGxODi
QBW/VQJPRLGKhYwjGruj0NBtNB5MpP6/rQDvxFbiP56sMJatMGc1wNW44PLmF4NtsISpESvMU6hS
S6tJbPZvdYFlHYzZviCtFzxcpRKMPtdyR0XNWQrHiD3xvp/MaaXEtsvqCIYvs7G+m0MjO8IzbT5q
KedLBi2Noh5qLD3VmgnIlGaHFBUD6b41eixIUYtNDxzsKvOulYHmOEt96CmxdiwaaopyI+ZpCV6a
DTJBj0NljV4SPyA29A5wz+EWYYy2Mt1hQFnf5GDI8xF/lzuSnMInPAEgYAOOInp8RMjRCVRIGkeN
4ewFA5+fks+9kIqfgBYyrhp6KU1CJLaLsw3exbdoe6wg6Nu673VTk+NL4rRvDoBw4yv82OiFyYTO
AUD2JwOd1JuiWA+QMzgAaD8YY6fP2DXsH87jbY6zFTgG6Akb6/jsB/jlnrwsPloUNPlpbMr6jMhu
sdx0Qyz9AmqTon1W89YjlcGhOLANTfOPv3HrsWpE/2gkfsVPDUCBIHOKV5UzKdjznEd4CP0lLP6i
DRlJUzYevf7bWFStdVrGWpZamo7e3kwxw4ykGOeL4xLGnihCVy43TbSvyCcVVW+DXl6xlNtZk7dc
i7UIXWZaAza9XVEFesMnW7rq9q2sLMpoIzJc1sHpRYemzrBrSIvumi8TY82Lx+mD2sKfiOnryp3b
6ZWhUXH/tlt6E4btgMs8RbJFgA6XmLUgAzKCX39bcauuBYTixWrTralfujziqyP4y5JjSOhGyWRS
GJ3n51Mg1Svn57PyiFynAz7/lT71ElcolzZxfnL9hft303jvL8eCx9WmFtXbtBUWPx069nvcmSYt
axCtTTZXYLaqvMyYf0ey+cBzqzFEK/UaEAxG77PhuEmn3DanoxwEdWFJnbpvC9mWZIBeDJGcqCJ1
s6pdFZjUqv3aYL4g95XIRhzJglQ0c1f3AuC9ROv8ca4sSKBG4PA/XC4wCwIHpj9z5I+k8K1ziEL+
A1NOFSDjMVIkn5ueas0rqsM2igJnSyRU+2YDKzGhePzyC6yAnAgmbaTZRs4YfSUXI3a3PuIpbfTu
RwIbMe8Ehrv+k+3VBWK9w4wegfBg84hY0GG1rI/Q4no3uqP2x39kpKiAZmaqgeTwlnAnKtABl8Ds
6yMkZP5MTLkMSAZ60y6XJh4KHLBKy4HEBdbkb15b11B1IAyNrFYFAUFoQYxm95diK+5eO+8KihK8
rKqOThLkNt9D6SjoBDdNO+Q3b4ETKrD4hsLdA5O4o5tKT+GJUyPCrNUCUoAUxwMHQ+g087KcXuo2
5atdnRleqccEhNaPhfbuudyKtSNQUbe28j615ZS+St9epWHC9Jf6ccOqezOC1Z90l4sdPKb67Rfp
keDe+r7PB+MVshp3xb6wgaa+8P05nxyJyZEnnUjZnJ2uSbJYjzQNPqE+G6qVp9pM4v7BHwiDs3ne
yZTDsI+6v0IjgpJwR7sE7cD/wIGddGYQfAVTEv0qb/3hTxay4CYSc4kRtEy6jiMf0UjGlSoAEWxB
mS35D9WTv/HdZiAVQ2PiaLYoz+9XXexGUFLxXPuTGTR3+lrGAZ6s6Yz2/jM+UkeVZtOBfQMq/wLq
gsf3JIs+NAhaYbMyuYA19H7RsNUfeRH2e14dqvTHGTxZz5QmE2qsQ69Uk34rU9m1/K/AQip6o6G5
7Wu6DjgnmAvK3ZAeKShXrVs9nGGe8HYM4Q21AQ19oaarQAX4qrrHmhQQESMUOLN3BgQtOmzualb8
BtqYCAg8AfRsJ6qZSelu6BbSnqN9v3A+vaw4zLVulnA7tsJqChlxkDAGhU9aVwC2TB6yMva5rH/c
gHCmnAQgGBq2SLySA68VRdtS4AM8hi0qEbo8xNx9sagaAMVBUAdnNbNxWiLgGVPZvJgJl4SyPtSJ
MUSEnqRNvA8B6dPECwSSd3RgHRG2+V1YhBuRn/uGrCC7XvyXvSSd4uxn+YEbdyC+qBoKUXDvVByP
0MuiKDWm7IhYcyzxSkA0KSBabmQSTO5k8w9/HAZZhAQ/STH0w3HqvMrgP1lGh7ktbM3cpwb4W8oq
9yuSg9t0mp4UQVYW609WpB7e5ju/a4Y4rlGVBbD+QlluwuhyAd/j6etOFQdMRkqAA3Bm94f/Brc7
lvVgJhHF0R2V+fcqDWE8/8v8r7moMQSQnH+qCRtUCSk1jERnHPJ/QB1nrTXGJ7efJ9oQfGS+76Mc
V66rZL67mO8Ka6TXn2cIoqiT4wipMT2HjZmJND/GlZh2B62DLXiDiiy8PumKC0g0K7hvPumoKRqs
tj+t+0rcicoPua0SH8yuQ4SraIxHVeFVMa5Y2SRRJgRiZ9Jf/N7540iGAHj9ZISlkj1kduY6jSTg
UqGX1Nw5uQwpfsEtd1bhIGqS5pIBrre2B7F00aBZ97BTbW0DQkAa/2+V0U7Z3dPaGeM4/KFGmmc4
D4pET4+u+1wM5JX3tsKcZ+7oTy+f1A6CLSjAUV4sLqApFro8KyR0+cFcDVoO/+JnQI9d2HnCSd/c
vZTU2JZx4ppRUWs78BAqOrUIJSpETOMuvcUKi+uRYb4Q6W9rnL1X/FZoKVIACPLm984S4Z4C1f2F
rIeIbwuADVDMWSA8tmq7yeFoJqLZdZMU0IA70IJLoS5kgXexcl8ETnTlyF24bhILKKSF4NgfZcaP
mk/AbLnBQmvAyl2YvqBpaQGjD0u7tPaiuSoJpOnxVhET3HlVSb+VZnpSSPM0uMESiKJ1moLAP6CW
1u/Qs0NWD+aYBBa6YEv69tT9K8TiRWVhpOqg1XlMrmPb38GwANArxwGgnOH3ZxcVbUfSF5/sj6ga
t1HbvZFk7RfjrG9kL7DY2O2Hbb69Bye3Onhc51phR56MoWPNjhL7bE5ifLkaQiwn/3jWNyppsALl
AYCw0IcnpNtpqUOveVP+SCHPgJKY8NMPBJxNRj+Me2YM/2kGTiDAoBapC1k8TZ8sS+7A9T8Eh9wu
d6wcm1oBACAbjVO/CgXDjKtKBOgs1gcuCWn4XgbF1LwaxTwBkNnWL3IuMB5xVCuvYtkuB0lkEdMF
JhcLJxXr+d87jLse3Psy7muB0WE3rlJfHueCpRiJH5lpi95YsCeWWbDD+hq8l0Gan0QPkpsYNyMH
d76yA+3X4Oiy8Zb4jDPEaKV0TZAcGNVpsNyhxM+8jBe4EUkxz84xu9N0lz5rV4hYCdlDca9LPbrr
3huLIt5xwRuXlpdnycORoNiY/BfYYE+VdjaESoxWseiM0UFoSfPbnRtJ6Q3a+tnEWo2s+Hc6H1SD
i3heg+A/s5BexwaQwhqI/rxt7IznFv4siZN8i4PMbc2IJpWsyveR49S086k8JXbJMZOQ8y9cOApl
R7//XvfgCq7SVovY54ztc/KitNZBKs+jNWYGkM9ipXWY73245zy2iSYuWgARWnEnu5euj3q4Ly/N
I1GpZtEAYXrRbw+628p4HWN4m7E7BZkpbi/5/9WaHVq5qG+81xNJr0d75P0uuPFdMIIPkZ3DYeJh
9neSeDnnzJIMIRnT2WQ3uw40g0GauXhzCOFL8MdmmHampjhpKJ2ssMf4NiI2MR7bwNR7ofrehJV7
fO/d885yxLeHSua0gXFSK6dFlmmjJz9rsXt7dglQ01HphrOaO1z1b6uvwlp2TXS1BWFmjElcQaYs
lkT98E4VG12WOio8J8jQ0s2paTH5pmrgvwqTFaS1OLai98x4efU6mddSdrvV0+NHol8UzuC6fwxG
AgraAencDpvRNACp9VyttC1r5BId4+uaJY1jWFpG+CixSPKNBTIO+rsz2+mLBy0VhwHRj8NfQFkY
K+otO34CrJdn4jUd0xpPpJ063k743I1d/EJs5k5FBFC5fhpmTN+MB4AJJsYxzBws6bLmRd7PMZWN
h3CaenQBciXpEVObf8nraeSGFi0dLAp9EIf/XW9OcpjTELbN/Jg3zoo/bz7sC18eT4rYz8jkkMYK
bJuNWDpkTsn9kHWqr1wfVk+/WB3o1VI+T1IRcrs2bpw43DiJ0w2ek8tntbzVU2LV9T0qPyBSZDpE
HlwppnvpoZjeRsUE9yAAQz759x1KwiAjtXPP4J+yTRemRLNDFOjgyofH3cRw2U35Ch4pHYXDsLqq
UcyP2DBzy2ot55vDdCoIiiOqtGH12ayu3uW4lg9T3FVxDTXmN8xVdIlvNHVmjgZfk0i/yBFoqbBf
pknvfrtZGc8Y0CpQZJYapETe+MScOAD2ZXd2OTsm4CUPTqOPw1YHcE8R3QnRph4LLKue5P+4uCRC
XF0CIB7dokKho0veWtXnisP+skVFOG++lJZr3J7fWPhDzxuWHyiAck+YadMcvkBi6Lbgdv1NnmzV
o8AnPSKfLYvLu27ttcvyQbeqt3IyEQasA0XA4OOF+4EAlZ0+CRmFp5df9dqSizWJvyTKn7Q+TAr4
YcpzwLuMNmIV4uf5lPG+MbUFEkvpUZnbbdTmmL3t6wy2heOnNmlh5j5h+FCOSeHyExR6FDf9skUZ
ShDRUfc1wXgjeJLj8S1aGg3hq36Rd4r39f71hbAgN4DJfrSuhVvVS2/WsTwL3oSQGOddufZjf3Q4
KwQOa2FdBaWoZcgZ/ZWMgz4jOsAodq/us9pb0MN8gWPCHllX1ci71kQDhY7HD4PYXWXY+fQuZf7j
svK6lEBywUgkY2fofxsEa/iOW7bJsig2jdyXRe+Mk9cAnlo1DpE3b5j+u76BjaRdZ6Mxdq8mEKOG
QbN30iOMYHvmnfeMcrYrLHO0c92hpcE3yam9g8g+TsthtHaRjlDX2Xk2h+Hw3KQKlNce0vtsJ6gw
6X3lCSMG75BTkw2/2d0tTPtDCZxR7tKMGYCwq3CF1ydBo5lZXTNbX7z1r3OGxU+wRd/zN4LRovwh
di+7hgzHoVIswGASdstZ4xKZHG47DHNjlXo+BWpd++g9hIgc7eV490B5QzNE2q0yWLrEkQh9PcqX
ytj5rQ2f+hcedzCoUWjS/8LeA/Zq91OFHAC3PA7ApO8MEyGEypS5yEGR+lpccgrHTYliMZmMo0Ky
alAd5j1in7giRFiKeM36o/8Bw6HwJhW9FNuINPZPC7QM9aA9U4VTcsxivLcV8evw2FcX7hPKHBG7
UKO0jNe1LPQZtjI+R1/ZME3Sb1bQiXf3PGp9c3zEBuLBIKhIEmddqC1w1KH4t0WTA0LN60MIrdoh
M9psGIllNZUcxRbcdylSE/fSlS4MdNzwp90IBQNWwFFkNQqqUP1ErbwB3pjHl3FVr8srUefga6k2
T7woNGia3/3QrLBrfX8uSbwmKYeT1vnIwrhc4HraLy1TGE71igkD7JcGqP59lbQguOFd/8fSOEMk
bkXrtry0BEMI0ZEm82ZkxQjyeB7axZtVc0giYfrZpplWtoAfPepRGh9s9uzZiVSVvOUPAb7g2S61
FlyTG8Iz19H8bjPU2GgHlHBmo3lla36alAmkzuCC38C6ajeDcwEXcg8FmiBcpdGI+cyLk/5DepLl
ySAKDRKz9JSsX6TP+Umj4jG8FrUL0+0lRgq2BDNWnH787nFZe+rUQik5RY8QKqNlREcIO3hhNr4i
SBsiwjrGz1+YzNAzgeJzRGN03MYTOsTfMV6M/7TMr2zlSaDLW6XPDonMPW/hErqPtLLRZ2P/h35t
z1RDz10bOYqW2VeJllj0N0/RzOZVp9ZINgdVSfNSRJFotNG71QLofyrQbBsI0gOETYDTNEPqf21X
mxKISmMEpqYhQV8nPQPSibP+klPdJ5XYCyOeDCb6uoyiEO35FJtxKJgH3s5psh+najD4Qlb8a3aH
cuHHUchLS4hjJ4Xzwl0wlJ7IYoAm4ZRZX6T3KK96tE41Cne8f4kA5qTTeSxJC1iinboolL0cyWCh
9QCRH7DUzmXjxlrj+JCvqMo4lilkN1ygR9KmADmEfMoxWHCcFTnM6+oowiC6Db5jsYFday3hulH5
kc6+4nyK63m3K8QH+h76mCemz2l7QX+rcSQBU0R+1tVtDcCcBmxo885vlFiPUTy3QGRzoyEEFDyE
D1BHvz3W9v8lybmf5iC3pvtPCMvA/ZJfhtLb7jOipM3Gi2AhePVEzeS7ySizsCTCELTbSpNbITC4
KZB8S7jArfqedNFLrnI8P2wnDarW5mmP5QQ/nSOzX75Vd3lxhI/359bFNL2zu6euqI+iBwGq7yEJ
wV0VlG67j1Aj96Fh8mYuMzyr1YDB+KOUbXg0ErsBiRYHrFUP++YLE2TStXPVopGd5PY/WhguapiG
23m0qqIvmW2m3IfugGWAVcDY2L170TaXiQytnRTPyQ9FvI2xEBGCN5Be/XnsCgHJqrtOaGnu6InG
LxSOXgjMHC1AT3+mH69qDwYqCEkx/17S1oyxx4D6oELUkmic6u6KN9QSMTgkcHXXHpx+tb4aAa+K
tZHQ/FcQp0WH9fri+QOqdQbxgnRfQM8AdLB3KB/mvD/YXJLATD3FpbXsQdxZpuYEenoi+NGrHJkl
RBPxjkOd91eBKmjMBEvwqYpPSTYbcujO8dY6tDsS7JT46H3cNuI3A4gc4DfJKfb7yjWaolKVcbq9
Dhy0szf2OBC7YomOoQAqqQAkxTu0cTwAry0erUs41+XTd6TYPuPSCEnrbeYPyLTr535pkLZxcc5L
1R9t7/nsKnFpnGFnemSFk/iQXFaYK9elozyIv6EsSZTUEH7LnGQGzv4uIRvZL4k2Q6e8gmRcJhtq
3A2zW4wCGkCrBD5vcaz3pidVItq8/J0jMBD2q2OsBI2XUO6GeLI+BbNoiY07AhvvC48XZweaec1X
qgAl6OndH1i5ev4mgaUxZMKxNsA4YsnKpLwsJltUcqvBoZlOi/x+FuDgBFwNYH7eHYvpXEUGb+CS
PPtWSzP9Ecv3tnDSi7LdER1xn6ZJO0MNc+o6XJygu7BkwfbdBlUY5y+ZAbcdmA70XFIqxGs0SLur
RSnVewMAnFG5vcPO6Lm0PE04iZ0o1u8ruE5YFbmt07UviRJh3tEoy71EoWpzRyJKMGnKNMzuiQ7Y
IUa/1Q3qBVsKp23EUROA+ErEYb+gwb0+whUgvRQij93PWqp22HLaEwK8guwqvL40BFSEBsheNwbH
L90+6amJmGtZ1RoT0dP8jR7m0zReKRsFIt4jATNsY285/VYJr34EqL0ZrBvfYfhwnVVwRm6i/3nH
otVb7+AslMVyCm9Gf05xoBgQNaarKSG0MgWyeZz+NE/O12bqZ4PnCwWZ3xiZWqm0iyxiC4bVl84D
ZlSlyo44KrLgdUnRg4mmP8CxRj7LHwJmfJNJ5iFRz0ixjWVW//XRwfjMP3dhzabDfjTUP26IO/nt
q5yipgxAkwaOe6hhf1nchBYL0ETeWOHbf3viWSZXkzOlmop9oyD6ewZICrVtHgOFFmQ+syt+bH5M
JnfjYFpCui+aqUJEBFamEOo+Lbr5L6enIO11LaBwM0ALwvt1HhkWOcWjCiqTBwCWUT4Dlt/8Fi1t
2XXP9ua7Pt+x3Piw9TEivC6DI2DiLR0L2BGEGM7VUmgJ2RZxZeUZo40T0sWRp8Ig3lxBFijFR2yU
3dakkEe4kpXlVoSbmy86gOGBx+6UsZA4iBWjeXq4gsfu9dtnR13EN3FFa/nHbgytImyrBN3HJrFb
GfMi+w0cod0dm6sZ8K/jtVM6sEw9d2nYMZGlby/yl6ZO7aOus3vqOjZtqDxxoHTzqcdtDj3tFLB8
N0HooexYV+ZzkThdcrTMyHfw6wiQ7d2+ctCIxep3h6ovp2vqq1pU76pFfD3f7pa30dOYwQZHaOhN
WxDXUJkOl0I/3sTpEeNlHCE2edHnBvRQ7tfYomz+rKriIpk3BjkaY/u88hfeBhSFit2JqYKzPa7U
DBfE8LvhMyu1aykRj7Gal4E7GQXLA8UUqv/g62dVR5yGD9N8V3SPJO4KJDqkLjiS2Tp1MeVHzxTM
M1MA/1WL9LNq4PyVD4rU4BW43aGUay9BSWeYarjMJqHyEdrARCtgVOKlcUEjzF9CcavZ0ThlEZMv
tS0I82uykJ9ZnoewlbhdRH84I799FwukJ6OLNKBZtQN8H4OYnOuqdrIxXllW2C0JUuiBTN3oW6pk
yagDqCtXv9t0YL6fBWGnazezU/BQrQqgRGj25jY2iD6haVQES2nMhmBJGcOVKI0IBcy1QSKLkqfO
w13JSfyd7oXp74DXTeTN6zigudyM/1zsxp8oCRvJIjG/3puab7aiwBqP2e4gfZx5ORypeqxUi3Xc
UqS2Fk7oNYEpbHg5JSzTJRn+xyTR4RGJlU0S77ufi4Xjlfm0eH6nrHtvATQsQbQNRlA2JfTNXS21
YdqJPTq4UyZVn+cPg/N0pR8f/HnjOmDoRIlalK4VKbiHpiUko77cbVorEc0Z/Wm2DwIUs2OLoAWj
TB2wBqaMIvgdnYuy5FK1UirOgQESiER2ZvE8riqMITESdPj2QAO9HXRp+Po8gB3bjIkSseeu1ihf
yRnzCucbeaiaND22JJQA8l3PnINt0kf83iBMq4Pic6jCwz2kTuFGw6wUvT/i8me5/7pyU9gYLWpj
AdfiOMonEYIXo9lOvSfqULed7+BCuevRNEkBFPIKLCnP9pDIJYI2k/iA20Di4l2E7y0wf3toxS5q
vEhfnLNBl8lIYuX1rzzpaXp6xDIH3wu0CoJVrkuhGoznvi7090BaNo51G0o/w89Etg2gndDNgQch
DFqI+aZYN2eNKUmThPVnToHTN6RvdL+GsSza3uarHIbFsyXa6IBsxxmh/kOfNCFDSo/jUmRmNYiJ
ze5Z4s69+aU67xtC1xI7agBXahRbzENj6lrWZDK28XRXXNrUY96pogEFldgxF75a9CpouYAjXOZl
JVSP2uS5MWwRTl1iDE3jO1/YERv6LMRYoLRGKvOfBxm1V7pfFi+qt0l0QXbo+lnYsaPa/N61hC0t
kzTYwEiLEib+0SM2kvU+M+V0pyJvzeYz9pjpLbVf5B2/OW1Ppbu6gik7G9lDz3nCs6RQi5gxBGfZ
MYsY/HlFytyfkkUiChvbSDZ/0iudMJe+QSEqtKg1hgy+f+gsvT6hOx50e/gvbqf+0DFeqtRQ72e2
3ldPGHFI7bRSxAtW5Dr0aSYeM6eXSBtZ5b0D1pRIFONlX1vin7l+fDOAzGvcutcc0vZAlSelhvYD
mFGVQtRdN8wTXsAI5Yc13i1E5kRU+AOOcEc3XShecWg4XvmSteXSQHCwBZxVyJfbiSHBfrF2ptBy
7rpg5cpSljVfNKBgOYepOof1jHMoobVEUAoypiJQ6wXWPByYFR5iPXJfFcckG5bVl6VAIIbA2goF
QLJaZ+1I6wDSWLoJbb7mnUNm05i29QkhZOB0Fh+blc3tGaQ2ivfxK0c2Z3Yr2L8ZcSSLNhEVfLfl
TC/i4LcF/NKB0AKPGYVRWpdm3o85gbqNM53SEbyvnuACrSi9+9dR7vGW73HLlylTlGTW25ldHhF5
Klx2+HIqxFIlMdpw1fqG+zyca2fcY7zYBakMRle2DNXZmxi6HgGfA0BAoCzlQJGGt7lRCCaEywuj
5jd7I4BmverWfeQh0Ulr8Ioa3t2XgBhc5zqDTNriYv+8E7b5BKsiASO8ioTG5n640CA1LoG93UAe
b9Qt28Na+yDWag8OdtkeE6Id7FWmItKv9H3lj/vGrtbS5dWKZ518r7xWdh11Kzf0MryT/nj8NHOg
TVg/pC/rvnaG1b3Fg9bLhIAQU0smZn/Qf3wkrsCExRrRT2l2uw63hrzHRIBxMShsiqmvCBClYT75
sKWVWVCBeZPn7DqLGBujJNCYklRui8a8VnWA7QbM8wmvh1sOiV0SyYL6sQvxewGjOO2xX47tZKxH
fO7s36ykCtoQMLquSBcEPhNqmtXm1eq5Y40mQPhc+2ybQ1Sg7cS976P/O3TfrLyMqzTbh0ceX8qU
L0pachcI4a2m5CHx5Bl+Rbw9WJvewI3i2k6dQofxbADoiMXiIOCbqHM4JRYyqmKA9742k71G3PAV
Z2fpjxoR5MQSUpzrNvrwIr40YjjztTtChnZh3YA+6T1EaFx5RuHGmqlDpgm5yKWGd80aqC1O3gvO
iwyXmg6QwbfFA8nDT+zuHhCABRtAYpLvAoO9PsGN70kJP/rGcayfCbIELcVjQENffLKLTLg+XY4t
EAdAC845agowevHXhZGCwBkq/7rqke14S2v8+DvXPFoao9YaWDOA579R4qua5GMj83hJT777u2vz
q6aT8WsSXlbscz7ViZgovHa9fYewRxklfYPG7w05Qp2IVoBQBUflwlz8vZ6JfAlpJJXD0JneA87v
bfBIpJMWEgbutGyBFadkI7tDP+m4FN1ZgQLoQzhWPLuMGYoayqSFYHkH0T/EMCc0xCCsU3AINMe6
Ho7mP7TQyD2nE5QDtCpuvFfVwmC7k8AH3U8/CKPXjVGrlPXmPO3z4LxSId5z9ur+cFPRzCjbRF4a
Lq1zjCww2iQqZq1hISNvDgvHulGFuHVgL5MPVhIpV1eZ8QrsS9wn1jMARWIA7DKJ88uhKRKE08K8
nPq3+oNdHKbRruaD3Z9ve+IB/mnssA8fSmVuEaKsiQmhKICQMcoWnpgEV88o6cplLEml9PJnDBXB
ZnVjMsq3zVuudeQhCr8y+shrEHXklbMx9CPWrOPPZ+NcIvrGGnqW1/rYT85KxmLu5fUxSVTL7Aho
fjv8aGJhXNhiTb5HUcppfyFzYFNAKObE9IazVYQNuZVs75DVF6vaILOatbvDw1xO/wEnazUeZ6Sj
1QD0DrIwdo2TRcd6jR32MeWzd3iZkoXCkqYh3rzWjNaoSOV/QsPK4kxaJlatQDrh496zsp97/EfU
yKOroI/68BHx32Y5GzpSRmuFr9TtbC+tQoxzV77m+FEZPeDigPTmmBoje4UCi3W5jtMebyO8Miu5
Xa3l2sQ6bsQMhIpsNfichm6tRe1YJ3YV3X3l4ankh7wWhMEtnPQTtred2IT7o+b9jNiF0zyInNJF
p425tDGuTSEVk31pCMQqVPSHNWeYNhNSTcYKN6+dTxiu8j52PhtQfqn7wGhED6PnQmtCrWagtHLo
0MhuwGBcnqsV2njyDuMrXGjYrU5P/ZGVIWIfxrNOdnIoTcwiskxtWXMK4oIx+NJAmPgkI6GLHUtH
qThUZ0hT/+/4xAMdHt8o+oELYmpMzEZws/61CuSz65+jFvhZaL8MmR5j0uWxtebrl7PtSEVhuUwH
xmHrGO9VF/GtNNRKeGFdD0hUFudXUOvAiW4tRSEXKCv/BS6x/8EiMnsAOZA/i0/GdgcKuBVfQKyn
tQdHz2KCJF4Dg85BJcSCfOGFKI5+h0t05/sUZxLZAfbOikXhx0jHr3vEd2SC0QqvhrytbiRPJ7k/
fRpoCrp7OYtBjWZsHH5ay6hwFzFLQZjtVVkZ4XOI5zBN/NfZr29vIstrpMQ+e5DDcBqZZWFmEP7j
e4gVdjuJjaMtZP2sByTC0qb8WmOrwINAvIYSU1jvbFm+NZXzK3rmZlqV5f4+hw8vJ/1jXCtO6JJW
DyEL4GLPoBOOMwZefRyU99nItux1u4u5op/Y3Sjo3HxYiCPtkyvR5BWBLubshVkcMokEfY0sNwsG
A7yAcJrmhwhLR48bmlMc90+9IPP+XmmRtXPTxlVUnnpgM7B0LCr8lYjyLN3CkAJLkHEh5tjKnXvF
9tBYUmWWdneoJy2ddEXs2a9j1JUjglsiwVAHnXUogWXfp8VeLU0kPuda/wtgGqc5NGZVO/bx0XZQ
TctKbYcu90QQN0kbQtJxrA5iOrh+VsnQ6ihIDnxJ0dBO28eUKbjJdoPjBwQeCno6xDsYdDJknk5M
yVrCmctJPIuy1h4jac77qHP8dDDCkoy64FNEYWMQfP62+XpEug8HAu4oKMZJTW3zRyNUVishJqit
Tp3Yu+YpqsN/tFWqkJDUpUI5NkO430ttA68CdJ61XXoTYWKRgmZgmZzBMOlvWBOvDLbyyZKtcdeV
PXHEPV7buHDwM4rNDfJAVfPiUHQIp9b7x+KaEPhIA4Tblf0scxt/R+ElkSDAWOYB9U2gqfmpUZBs
Ayeav9+fcO5slk5TMQFkoPb4q5JWg/2OCjaD0oIR62I9OMxUF97dAhCFs1JekzqY8NCegesSNvRT
zLiTbwwM9EizBiw/gcQSgEsi6oWX4rC4rdA1Yu1YabibXH9AGnmWaLU2i+lFMmYJdM8XxgA1FkG+
r/H6SGZ1q810g7BZ0rFMYyGQHo1H8gTr+XthemD1ibfeMyvOXMU9qDaLnxmQuOh/CmbWsCuSAkLq
aoy34tSinWQrY+tJYlzQHbcsG31QWNAW5KAoEkGIrtnkq+RjF4COrYLAY1beQ/Su13gb8C1UYryp
m/MfN3PuZfSaCUbKheIrOk508g+DkHKIkMp3Fp0+gp370kRLLqbHqcRxRFAhG71CTg1cIZlDvF1v
Cry1ZXOPeoh9sFDzk+70fddaI8wT0KX9Irb4D5bDhiYRGtjgly9sKAuKKRITzeGJQlsv8n42NfgI
gtFOd69xvsEERpOLunplfU51hvTLa0Hg8Cor1PCmYlRLuTrlZ3B9iyq+V3B78qBG9nNKPxcoqZrk
5WQGM7Gb2B6340/iCWq/N0w6T4lKoiuq6OLfLP4L51kbRbFBfxjrBKnXcbUOYHyGj+L6nPfAH/bN
Iu2PzAQfbsngwXX7EKAL6yyue6WQhj3Shez1tCJKN/X3VxjjO1bRdKu4+PY9P2g/zPFemRD/L/R/
Qx08LIwTNxKTU4Q8qmC2eJsu/bcC8WgakbWB00Gl2E+DdZOCQL6PMtB9nOpWfIhtkkbB6tq4W9ES
NpM4YKF7cvxj6jnAIv0Sel0AQQXbaoZUSfkxgahP9EdLOmtXHkeztyAj+KnozvIykgJmND4xpvgA
oMrUcpdCodKLmDIFhE1GG37PGsPZyWhjjNL524ZY+EwJeNn2yyvuAGqjRnXs+OaDLXZ7Qqv4B3NL
tBZuUrWiOnCI42KxV389IIK+E7vQ/A3laVZFj6di4Srdw0uAdPVRnb4LfC7tTmG9mMU+Xk/S0psa
0QAA+B8GybELYt++wGMJix4kubBJ9gpp8fvya/LRKDmrHMuabs0tAKkvkRT1AsKdZOeiMyyETfyT
ptFMY03U1d23ljZDpaIvaW4p/IvQduivwPWnJ9YRNfHPgYpwFVmxJNtYiQGa5kaGpeb4jCkFv47b
r1AaKmBW+CzbM+prRdP+tHKV8Qb58vfledQSP8C+Hka+PvIlpF4wD2cmqct+7magUUpjWdRRtY9e
b0zgyDiGMxhWwxVJRLVEWU7piiJLSuSjBInEnsywCSBxwE8TzIFkROWAw9VG+u9BfmUwe5MVU2sP
6lM4poAoN0JqOXYfKJIUqrxw/+/y3Q2mdvTa5b9dx1oCSvJWcx7vy0/XtZKvtMa7c8QBw2Kf5Npa
twmb4hCpgkiqnGxFtRRwX5/zZHg0x+hDFGm/rOknS2yGDNSlxElIDy7IGXfDd5zLnAWNMhcNgdlU
rk+DR6nwdakDhGcI3iBX6HSVfv9kFTQtXsoA6SSJeIOKNmwAiNfogStTUI3Q1jCL14tx/g8VdoVw
zwPzy9QppqdWjbT683XmPBJ3jcnfcQzpXt92OzRqjAPSBK6yxfVccmzJG8e1qYNRL3eZMZO43rAe
/iFOoQ00j+QZ4zUqgQ4/eBsEqVj3duNsWGhEN185nLzTHUiKUIlzwDHK+iN/qJldfZ3V976Swrrk
CNT4XwEzMAQnOiBDeE6OTv+uypmPhZgJVZ04K+N2onEXKAv7caJOjpE6sT8PlpUJue1jTUzUcad8
X/BDG0vdJ1XGR9bp9oKgAA2Yq9HzWMJXsBNcHuN5zNPNRylSlliehO718vVkjxso+6IKDPlNnIim
0xooUufYS3xX6Qf2eGsmqH6TU9fn8VM/Ai/mdzki0lM7eRYx51OrvuZH4uYPYWsvD0QVxikGXyPW
xdt5c4QNwXjV1qwevf2QrHhueDC81mt+lCsCcNh/5Imhd7hSAPfFEy/DKIO/LdgTJoRBatjSrslD
94hfhEnfAZcSxqIoPlcHIANyH/loUPGnfh2lJAnzK919jjKdBXbFKnepVo2o6ENTcNT5Y1oQpT4z
2+G7jo4X9mIcZxTGGF0Yxt/Qy1zhf6/vIOmLWlXISEH/0maoQjd2It6JJ5uDzHNiD89GYSiKPwYQ
B/LcQrLd9OvWen7cgZdn3SmzwXwqYZR5veTbi4JiAbnzup4B8R/Iz9L4EYvYeXjZ38vAoyeap9iQ
qmWnQG0nTmRfgn8FOqfU1e5Yi/fjiJi6WB8x8urQVfZIyxklbdbIOrFpxxryRt3CLZOeFMnasK6L
SL0/g49Lb0WaA3rGw/XqR/ex0F3PDzYesv4s7agMgIevRQfk6D6+ElB+/phQB+H4IVmqTbNBuw7W
cfG7DAupUvgnrjXGRRCNYoA+FFRXEZVpdUbLoiywXFXfv3eJOj3jzm3isFraAzY1n6bzPMcPKpL0
l53REZWDclWZaqZ95rgvShzo+8rMQt5ieo/N/H/6zdtJErgtf8ieWkGbe+5oL/GcSfrVBCxKYwO0
4HTTzp/m4/5bEQoHe+8qrC6R0eE0+RFcI4PJKehoBMPvBivxAHVZBDIOAzim8EYlFUWCGk/3Afot
ipiXU9GjR/8rTWk9wFGVlWWZckol3GXvmR+06LyN4omBqfxDBGD/1zC3Cp8pDUspVGVLtHit28eX
33kxxJqFkNhCQ83YY1L7MrDKD22TbA0ghvodA6W3G1nkRBoIQbzIgzfkroVW5FBI2nI+U41QmVWp
8GIFH2HPq6o5o0e+Fb2Ff5DtYPs2LNmJbEB1zhWP1rEUhRUWIuez6ntJgG5YBskHtsEvVmSyvoa0
dctSeLQngBz8JZfUbYqerpUWq/hUz24vKh1CbbwXYYcQvKYQLKvcBrE3aYMQEXl2cPjT6ctcIkxV
kNKhBMXj9IxHfvNZ6dE7Y+D/5y8/b8s4oGQrPWV660ZKP0dVk1H14CDABAtCQNc3auOXodWtAV4E
laS0JRhj4m8lU0jqY57EeIuqTSw2MGTZXcxLHV+HljMzKU07aCI+imSB6FeX2DLctsL/z/NBel5q
QznxuPMztQjK8XMar8R4RQgIz28R3ZSGVH1hmKbT1TcYsbeQbCeaeC9zCQyrveOmwIYCr8RBdtzr
6t44j5/ZZDsKuUqIkcpIDpnuvXDIUZMQHZLDrEC0cSAxCcGPvk0J1hiyE4Z8YlJ/8PbhiBHrbCZ1
PjGFyRwlhXU+X75+J0axJWbIEfp35eIOcXMyvPi85vofU1bCeJ2bG+5hdNjoqNbnjJy6OXxAJp45
8iY4UmFXqiTmM/iBPohmHb2L8AACPUhtmNwpkBuI86NiQDUEVsDtvexCf0guHTQ9dfr3PHX3Fxsx
kk7EqcjLcmobkHUEmhlp4jk/tB1/4us8x9dzOY7//5NYIpOBxKgAAEJ0PHFgNDHqJXFShAsTt+ZE
aBsX8gRyfdMBBMnpTN3YtrXtqIeGwdoAiudanQ4tNPjRqScTxRpcGsmLLq40nh981nPWB84ZreMR
il3Whcqknp2ZSPdgy0hqH04KGD+P+kgANB7MnOiLH2s++JPBqMAc1V0cIlIIyovd2Kp+rKcsz1ZR
CeD2ff2Upsqu9y3nHWz6lLSqrOadeJN19zJ7hfLneXh+GkBaDAcQ716q4N1yQPYgX9Cw47eAemBo
wRfkmQS6b5PR0mF5M+TLDiX8u3BOGdoytkCkH+eWJ3snIWI/3j9nEQ+PnYLM2VNrphgHlsZ+VqIw
K9Um38MRIqRLsLvQj+vcXIi60atdTGpVRzF9vTSTm7NvoZ0Qr/wqmfvEZHnUVjILorV3MnK3f373
hHHrrU2S7fCiCLTQtUzB8d92u6BcGrHG5SIlo2Dm6HApkUtPjPj6G/J7YJI7aq9Pa4RfPSntmwgk
dtAsz65Xgc346PVNSc7RvodYQSOBQYgcwc91lHvBEvG8dHQnpiLcPfMH3pJhRw94TeBFsPsoV0n2
6WW2Ukas0CibagdPg4g1vzEp31NrPbapvoEbuGcPe42cegmous27BlJ7Sew+RHegJgmyiOkQGxFW
b6nSrYR+/ys4apD6GtZF8TryM1nMxmeLI+owHJbqvk31jqwENR4lzwAaQfMaPd1QDBPnKmE8x0RA
EFnmj2gnDK5TYrgGJqJ1Ge63e725yB6lwts0rtoZ6PvL6DiSFFQgkj3iIp+bPhErj3Ibpvg3rHAL
AQ8jckIgblGx4Y+fVELLBDG/p7HbQ7CZV/fb7es9UOuH70+DUytTTWZpodFyd5eHu7xQ4lfpRQHZ
c6GjmWPJHpLJfMjxFBVmdcxpGePcrYjmoBKu9BPXgo1VIMhHPOUOXKscqfRyaaVrkH2cq6ShB3T1
SFTCjS7Xr3VQso+t9MECB1r8ft4fl+08hSeCAQKDuNmedTDM/3DuSkschEeo7ioqUSnB1aOGSjK8
B14YK2Qxo1icGtbA7QbQchCQLm3MUgmfZpLXKTY1MeQkRSGFVgkhBpFzTNqn52gsrKuacCSEId+K
uEhkGbde3WJviZFObvTiQyptxPrZQ+pGi/G6UrpMg0Q3rpsaiUuFcM+QAvgZgePw6qcVMTn5eLvK
hrbrIY1lf1cpZir7FmkpO+gIWIOtzh1ItDQt1+Xu/3lLCvc9wdFGMMZM53/WA4RS4ox4DzeS3sd0
309N+sApCDw4hKEIF1vix6ftOLvP0i9uOC+Am3RBRR0RYJk+es1TzrgYwNhEiICCbddH1yAKjEIL
vASRXChnGLbsYyM2ToB1PkER21MUZMbTwx/Cmo4BB99PvuiMcaCZKKUfkCXLkg+n3IjeRfDCJFvb
4AP+ur8l3gWYhE7a7Dg2F4RIvFFs382bB4rxG/6Lq5vuLsqEbIJJT0iqeLycxQCjD2xlK2J76Tn3
S9DzBFwfBCBoSInGzji1pAmtvkd52D/k1D18OvA7no4cbCtAbI3JdYAM4n0fFLUzDfjaCpGQN3d2
nSzsJtxqfHM1DndMpYllnMTLJvP/tvtmH32ULAG0GwNl9t7NXMqLnAmipqdi8DhkwGjeUrtabyUZ
41I9hRfEDXglHOecCzkNgH76+bydV23/AW0OEdATh4WiTIgobEHw64N4BG5okZXsbKoQPxNeXPWH
+rFvZfCL5nWqMbQt0k8rBZkTOZq0/IFkrS9wylY+Vpaza8KJZusIvfNC1aNgbgQbCdmyHdr4Mpdw
vbBdioAHzVuxl3yvjhLZ16T8rl2PAcUPkD1r++w7d+wqaPtCSpyjMji+f0TkGDcO74t9VfbcNfq0
dqsLQtvUYaMw4gP81+pplqEVAIfI4jnOeivcNJws/+pz6Qi424AI2O+4O15EYq9JJyPwk1cFTpSg
M2sBGc373cYzlYAC1CsPLBm76yidxKe/wJhE3vsj0XV7wBA2/UMkGAGcf607w+nOkIqSHU+xRvcC
icYqqGTgGzv2YrbHViG0yfMjiN4ktUL52d2pUUVrooVnnoRN9NQ3LCuPkBX+LfZhuDWpUbB7Rh16
FNfcE5lGwO2mM4hQfwmZ9AOueDpSqk8xDVFyi+Bnv8W3FP4qwrjSYUCSU9QMVkzKk10/Cww+/OG5
GwRUq/3OfPsmcojw076WBETKGlLqQwTgA46L/ojEXjvngw8cAi+N+Ijt84awQFqXcEdtcyPVCb0O
mWonIPqqTB0+wB6ujoptPdvfKTf/8SjMwyja5qrcQHHa420QFDC3ospghjPNFha7S1a0das4YAhq
fKCkpgItu6o7L5mx93zOj7rbWeLy4IzRylyF1Q7zUUYAtPTZos0lAf/MaQVbLzV56Leeo4xeMifP
HTeV3Pk7H8KJp3B3pgqBxj4NvwojbNekTxrAC6d+jW/H8pkFx/3/lBFlTdFU4oPzWBlgKBftoM3f
+Bf6Gtg7ZuS5C9HcBws2leQSZ+MYffGDEIXEeJg3OfrVDV71zUldpdypL7fdQpnPXEUkjCpMWCo5
Pd2PK4UgDXGgCJ1tMWP9+JPB3cZ/T7vPLYj573WJL2XuFHOXfY/YSI8ioTbBBuKNRGupGqXR5YQY
96sEUWHdDrj2rDJyFVPI7WMnrPC37MxXiiLSD0qGLUmwOfNBh+QXlY+5e9QwFmazAxizYbqAFZCk
qIbfOXMhprzm0FkBLrn7sxuSsA70QzjuvGS+US1olIuMDYZL86cdSQWhckiRv21LS1/3r1GnsfJo
nylvCVeQBc1HrvuVP2Bj9eIVmwX4NA3g9GCjg6wWomCqZ3NIvBAwZLkoNHXNg+cSnu0UYApUBYWv
9npDQrVFJYesuqdSuHRaT7Do9Tg2/KF06HmD9eLykz+oYOqBx/yEZBRo1if/VRwlDqCf2pIAHSnd
F5lnIIlWKUqcPLkc0danzE4Dk402YwvQd/bPGIgTv8/BeciBoSIRVnlvSIL363a8WMb7u8fxDfwh
A7KESp7fNOXiFAOeMrBXfnje0N3swOzX0tOS7tcBLncX/cY3mj1kxC4NMpDNsFyWaxVSczj26Oa/
EPp0FNj6YOxg1Z0gYA0DfnpImGOuuLxLLPM+JQ6K48AO6mbx5R8AQDwRYvnO2z9kibmXAMXSnK6r
9d4G20KI5qzlGA7GSXQBcg17BEv13IM2qqAJNFE+F6btW988VRuEdP/J0UzmU3hYJ/5LGqadfvmc
kBvxsE2olNCPX3gD/MaHqBWVv+4J5kF+Op9L/OSXulxR8hFqNzbD15hPjsdC1tE1CrezTeOZgL1u
xZ/sLgsNdDHZvAwEyNav/1mLbZuYZoshpAKILIcnk/Na8saG1qg2G7aqWSbOADSfsmRuJIQFT1A5
Wu+2i/061m3J08jlY12sjxPD9wYAWJ55RbPQtDEUed2HG3Ar6jXsUA9Y2E+KMIICEu+5r6coWdiO
TIPmCWQT0yoKewTAKNLeC3cok1SdX6cIS81Ez2X+SmMMK8wpaTldNN1p54PodAu9QgdGSghsHYT4
WfLECDv9puE+D/bueD4i2YPZ6pBx5sC6Ro93RFXaA0Y3gPWhJbJSbCG2IDVQwFHF9AfoLIiz791M
KvIABthrsHPwWWMM+e5ilqEOoB2K0hWBNydS6a1ByqPHvgy+05eesod9/ymrDjoMNzyABfQ/SbMP
eBHGBH8Hrv8pNuiy4HsqD7rO9D8RjwCicHDHE2Dj+8CokmmHaVUMcrX5VlGRN53tcD925anTJ9gQ
02eTRytdGzsowNsQGU3oem7Gy7O3ZqSD3sDtmq5yLZNzlDKP7wIAxiTJdSAtHG5BB3zOteczvMuA
RLXxevMgV9vxF685ZoXwZMzvNaTt8WiezN62rlwwyswXPYpV0Z3oNzxioZFQVypVWTon24jYr/QZ
bH/U0EE2LHuCgIMTkRuFkGLdz1hsF7NWeGr7XuH56dhFX2LYKXQuGlql0cZcKTJOWOprcF4j2XJo
VEDM+k0yyeshQd6za50A6u6WDToMMW9bX1fn7xqFAgh+BWeyp574/XLJY177D38KelE3d0dvFk0t
lLNxFH3v3cG2q5M6jGbyAi9ZwhrK2PREfXzkDAXqpMg8f/mThSXefvU9vOtJeLz4JdvLJUS5rW93
xTFAJRToedEviFWa2YpIrWu181UuFUmhFqWCjrPybmzVGV6fGx/27hIJzpyXQpW6+Ic6faVKZR5B
ckEmIBpciBjDWyuZgTXSH0saitif0ixRROgO3fHrjJWrofFMCwRCX1vMJBCcHdE2htW7kmetLq5d
gz6rwhmFE/vuNXq92MdJrjyd5BW3WvG2mXZ/b5cgUP3rkrFz9pi2hHZ/0au/P3cUbi1oorv1i3Do
OrATWdQO3yY8jsEwCg6mwMHWQf2PO25Cb19MuIBfbw6cAyRrYFchkNO2K6mLT5FWUGzGlyhK35+O
uCi6rdJj9L5TT4mOmrBBhsIeThRgcKMI66KEzTM1rDAs60g3bpC121EqFriVZR2ZdGmaTS/ek+QU
GrpoRErMF4uSiBCyWi0ZZhX5reg1NKbcUJm1hjUiOS71ONYFZVfFx57kUuLdTIKl9htsGi9RHSi6
+GKCfUPzq7Pfike7NyMI7+FtMGvoriyuWKgUJpynj/OzvZqIIXjZkYKQc1OFC6z4DIDdZIdM77XF
vr2t0XNHLk3dqANtO2x/GGZ22BOSsAtiwLfrmzx0bj582ebmq+AaMizSbYm6WeA3pUb8xQUdV453
4EvEtXIo9lERynna+K3V8Mrn/XTqsEL82yP3AWtShCQMmZ+zhnp+Z09lJj+NJ0HDerlQI9HNTIXE
oyUs/8kqYH+9m6YsCefxmZY617jn4ScBSx/T8T9k7qVMrGDMTPyVq58nZWTpzhqPE1vAyd0K1d7P
ohvFmwX1YbQbZLjUal+KOJzjBNOP7BncpFaI/pXRU0S9Cvi1gyQoITn3uHjHTCz5AP2BUXzwlp2Q
yf/ORMxL3PVZo14IZDH+t+MAvwLbDVZmUADeGSFz57gis2zR9dfswbbJk5R8NIGwIhttNvJ7le3l
1qk28wpJn2j61MeweeKrGfQqk+qDm5awhlbhyb4LMdI5yfy1gGOMwcoJm48p/6W98Kos1sTI15Jv
fXY5241yqRs9RqbBwn2BB8+cExsdlE9VK3fAbDlCjCqILsuyh4FyRbNIL5zUhk5g8UXOF0vprx6Q
04TAx3HYFD5xw0yoV+YcuIFwI5RxboGDvdIWCcUZrZLsVVUmKS2Tp+k3eeubLigp+cYmxR5JjDoI
YwDJtYQrbrMIQ2lnu+FgU0vgQ3KH9Y8PvZladKc0vq8srxcN6UMa0ADr99fsE+rcP4R/GdTKP7xi
CVAGJ0r1mncmCsZfK6sDCjQwxuDknqx2V2AkGdhn3WfcXmZPZQ6Q4U4yob16MVsWnDA7nyj/Kybd
bfULQQIB4P9+8XTS6R78zwbpK7AkQ+IR5pQlQC7tx479cG7uHEvPHWe0sAlzXCEHfOLdtLVk1hVI
+73vy6qjvZNiOMtkdtOnIJBLTv6G4VpEsvEfz2mftbRGQUNRUaVi75/xNmepxvLscTbWLkQei6KJ
g1qRTmeAfw8xl4wEMHoJbkiDBW619+QEk4+n7+6lA/JmThUlGO10LloL7NzHEPvSTCM2RYnPO622
Scsd17iSa/B8chsNA3P//e/kQy48z526Ivl6UHQO1zi385ktqh2TyPFZVX9AN9csdxw0WU7MvtBL
zcOcvualKslARk+NipUQF30Hx7bTeDe6WMqhppWkGwhSHEFG7jVh+WGuXxVLvI3Ntx9vWS+Or4db
3HlvDqkQnPdDi9DSmV9TwoJFQl1VMVBpXQsajWElSD7cWQHCirw9ajVg1GD6vhlz5vbOehIGNFzo
2acoHt/kE1Rqo3Ic9LoYKiQoG3MFALQqxYQJ034CLnWCGtp48r+G+XTZaIUX52VhqSLA7P2Lag0L
0UXRlpCeqxctFlipO6cQ3yqI1yOKu4OZUXZcB8AFxIPhb7S3YAP7dJLx9CzidHpyccc/PKxUes24
whZRz5B0Qeh4xEO3a+3p7DUxNNdL9KRndOFZDDOKRQldG6qvqFJ6OhTsggt4MZHrw/M/6ZwzYBCF
5C49OR0aw2FD0leAPTY9IU3YCk+p7qzEs07Q/rzVhDrkt7pEIj1CU0luH271bTMdpLmhbhjX5B+R
H9lLMxuMjZTMRuYJ9WQwaUJAn5Q1VGtAG+HaUOgUaVqEn1Pbp9bd7EDqKsdQW0uSt2eYpspjB6F9
AJSvdU6Apd1xbLo7PhOh6qTVLwwSwT4axnEYqqFe3Ui29GEvQoIvlqvQcpAddtzOIHgvuXZSkKej
4SUpi8R1Dmf74/E/Z1mHS2EjjipKTZHM9Kt8f2EN9a2XUZ5ML00zyq7aPmLoc2Z98EbwGRXEIKQP
AzTmO4RtAnpHDP4+jmrJ1U4F2O0IwojHyKhpWxjgrVGlXvDslBdEwGtvH1iXhO5oENDJY4bEYkGB
8fJ2kLySgXvh2Q2sVMJ/m3cuX51NJZJs8E0io6sZPdaHJVhi8cb1AjMv+4D0Eud2pZo5Xgh3oq5G
PRbVGpCSJJ/TEJ/z/INtzgZDiD/vFAwOqgr7aDEtc0rNhW7zWs2E3BjM7tqZpys74zH/6mTMW3/m
DdZiwiDAekmO/n2l3Md2h1x1AHRAzKpb54Sygpo3dbMeU7oS3HWuBFGWK1EY67QGmeT+/0XHALSe
aRFVWtpFbPRSE3n9hVvluphbFcR88uBFuJfAC6pgPWKTq/bzSC7G+lVGYr0Xm2n1xP3RZ/9OJYz6
m45dpEkhGiz/Ls9OcEhFDgKwuWeNLyOAFvOpichocMx8cv/GfPpxGA5j0ny8Yhhh68sk7fMU7Lyi
7nsT/XlYlYEvJ8u6PFBJY7EQJd5Q6KnLBRtv3dVgILOeTEoPm55fBs362FGLcIYXuOJjqNnYnD6F
Cr316MpSpchBlUwR0FMAbcJq9aR9IpwB6gZEnP5eml4Pa0DSs31KZzMgQ9vPuH/BuLZ6x1gNcmq3
9dbHR8ymbx55NuT9ybYDhYIeAK/T0oisFx/2DJMm87hMFRbCw/SXarLCbPBBJ14l25Opky0uqiPD
r+eQdXHasxUZSwKWco1oy2WLq7b+D7zKY/FSDgQWDvvCOBJeXkYr9Ky9xkyruVuVaIDO2FM0Fi7M
EOEOSmRHjwkvrqLuEWj6DRLh0tIH0W+RVYDSRXLAWxWOwI25UYnbxQY/mB9gdagGw/1yPVapiVyM
h+8gttEXV4ydx+ih7paBK27p3/lxavGy5F+jv907nazoLA3GfM7rVLiMDD0OwsjX2O63k3Xc4/+R
pJb5s1SKp9Et7mTCtrRO6JlBHer5i63znQikXM/ar7qxXnrA4nnwK2X0ioJ433X4PwNxNX+IRsuM
1TYh6UcQ6Pi5M/rPb6+C1Wyj8NgrRwMcI6Jg/16WyFdWjJo5XVAqsVDD7K72twn5X+jFcsRZ+0nl
A6AjZiwYdyfm9jk5kGl76WkQ1TkMpgw7zzqiKzq7pg2HNv4iYsRzsEkX+fMahy60YQNVzSZPepd1
bdr2FVKARpeRlPglMZ7H2lK/rAh+ioTkXo5RUWUNHczJUhKcA8UuvQND8jNgumklBLG/wf3C9eKb
MgMGM7PWcr2U77NVLvOd6SCZGDmU5a0oKat1IP6KCVCzpo68Uzb7CRsIPoXJiNaqvENn9CfYYmKg
1dVXV31HSA5EDSRd//y+2Rk/vGMIkm0as34zqboiRHa7prBZcVRN3k9PgJFXpyd20d540taQkaXc
ZLq+iJf+AM5sAIj1gByrasDKPEjHWEz6bSPuyU4C+Db956Vg7bHzlopeKv7D3EQXByXXxwsioIj8
eDZhHRa1TeX6M1k5HWE8GwA4NgAm5bkc7UkKFmqmVbBsMCunBaTbJ4Z7BAmKP6D1xQNu9e9Z5pG5
8i27mvu5lZxGATkj2wQpLlIyk8WHJiGDZcutrX/MiT1pRSJ6esv2sFdUv/TVhirN0iaTt7O45PkN
JyYQ3/A69oHP77vgvzNLfYv1YhHj+Y0S/JiEC5i45hPFDCZwszJ+LdmLwe8msVN+xcJ7ejbpx9s/
3lc15JtC/9GBPI7cmizLhY3whUaOHtd/bZHzJJFYDV99Z08LU+kGzoRSJAqbcd5H+t2em9rcUi+m
qClSuziTzOo3cKcPF5s/fj3MQl5WLaXnO3BDMC4USBSecQtCEFL+jUjT7xsc5Amh57OnC4n4BmWD
he7RoYI5UQxUwhNv+Bfl2GRgNb70g2De4j5J7Y70cd47GP9seBYZbgsMGS+jhCHxYCZzYu/HEK4P
eNMcMmuVRyzCXW9KseXf2K4os7fVtKgtjRYMCFSyzR8lU06oCdffSzZJpAnUoj9JLspKPC4HOu7x
Ss+Pepuk6ablIRO0Qj0VEBiLL17JJYIHlZp5In2osz+WAQwbEiq22zdvRyjNgtng1dXaAEjvWL9y
2nvXKbT/woONXNzj+j1ehpd0DeHqDp7GTxN2vRO6qVceasSofxqCl115f1HaWfZ2LaB4AA7ms2ru
sqmEbA14V7+YhH7O30cTCLJqmTLV82pxphx2QhmUU7lSA5/A70y+biTlZPZcazs4lRn7NM/bR2In
u0kJLBoDjOb8U49W3tQgsNFZnKiMDDi6/9JBwQSeOTSDvrfvFvfCwaTpQ+R+tbIJj+DPfh52PusX
43WMjFqrzoR6fS+HEKXnPAYxLNYn5mIw/i6z4rUwKOp1aKWuVG8utk3ZqJZFoKDdN8son711QF3T
eki2dW16ADSTQTD3iqU6UR49xlltnHT+AaEFnpRd1QqcT8Y7oGJgjhVSzlIyaIlSM0AVyCqnZ51+
csyMtlrRlZFtoBoelRxgz8A9Ki8nFVS+Pc+nT3eRiko48WH5FvgwcUYxzQxhPhBFL0zwQN2Yzt4g
K6kqj9Y1IrIjPK2UTYWZJWhvP9f2kOnL4AmieqTfYMipw/RysW/PecQMAylz2IgX1yi9OYZof3b2
5HeoirYtzYZQbk+c/poT8unlkZ5aBHHOggQKVplmLQqR0Vek+kc77v3Gu4Egr9GJQTZe8y0WoX2/
rTZ6VPDQyXu/VVPzWkOQnVtNPVBcobzf0FxFFBWetVfDU34O/mKUHQJAONtpMHTAiAc8wXKu8t+u
YVVBCL3My7HEqUZE0stFxHoS+q0bmXQb9bl2Qt2Y+3QzxB/eC52aGQYZ8SUb5oMfg2LXaOebDpVf
vi4+iIrYLxyuj9O2l/Cp72/UvgqfTvg0gCpw6hrq3kcJXpm8FvpNyYfadIZj/UaVumDmBcX4xfCu
QiqFIl1u0xZVdIwR0qS4yRPnqxMRVpIFbvoQ2GHh0b4G/ShtQjA5WTiPoqbFTs7/ikmLL+v1m3g6
DMOzc+zv+TrrQMzUIQ5oCHqCakr26LYbI4Bez8tybKQB5CLpcdcfYNWjHSM9yWv5nD+3tRWhCmoh
P44mnXzc8h0WeeQ2G8RrtWIGXvv4u6GwgOZmmTjFnRMyV/KKQRu+0RXAlE0GjRBFNirOCp0G6jdA
Zas2Vm4r3ECuM+T7ohQC0Zm2ZYIVn53kVAuB89/fPPZ7qzyEbPiDkmsRqB1ygjKV31wwyIXBYdaq
ouAw497OBCWVIZV9F7HEGx7h2nyyTCEdxdFZ3pwQIPRyqw7Aglwb+y0m8jkhpv6jeQ8C5t4XGnu0
rJSKdGX1PrgALMVsLVCu5XFxQsWH1lyJrYzGw39ZaSxCFglt8MQdRwftGVpyvqhtmd8ry6zR/lls
S8Qy4PcsN6Vji2ZNN8dO6p0PvNRlYeqFZclefhO8nTahT5plVhKL90/xP5TgDlpSgJgRu20/P56q
hT4s4QtZbfq4XpBnufBGQv7MxFppcnP2pIuv6F1dV+f/imcudTuY+G2fD3PKxcyXYLdEew+UmwrX
NKVszkn6rpW3iILOpcBjmBQAUCdm3NqpwSmL1/9uVt5i1dRjVPxQ3rJ4vMQiYnUwFPsnnledN4TV
zJS+XbcIotx5skLqLa7X+hNDZ2zoDyAEo11eXzXqTlVsQWKt20OCRUVxx7jZU6WPHcBJc6/s3zU5
4J1Zsy4tFNgq1BG3ThAUWw8lFwkLouc0OjQZn77eCfJU65U5Wx5Kwx7fSEtkwWPRXaMfDNSyAeuP
lTwiz5I8B8KRCPLdzvJN/0/TDCMe/2u1lW3ko+94hzqISi8lAQWPtHphBHiNMbgej8yumWhCz9A0
XCSHU4OvvBg1EbH1xHMPqyg0UEcd+fRitzu/o/yIy66eNrNb/bJKbcKQO27YC76DcpGNBBrZGRUH
v/TfH2L0cQt+54uSholhrRLlq/Ndnrvn/ccwHgs8NdYL5MxlylS0ydCq7m+hjEiNMkmAfrLU/AFl
oHkaVcOF1RVrxPem/GOaKpGL3ZGpP9fMwE73FZTyadprqHor54CDce+fCJEusN6lYnfFktfI/P3n
nllPr9TgPlldbads7Gxp7AO268PKJcJPxigfc9DrV7iXt/NHllrU4VXJmzdVN9a6D6oqG3gAVhTK
P9WAeiRVU+mRonu7HuxI9UWS0+TaZ5kj4HJAPvSpruQ0+OttctscMUnm0Itnnlk9cWLd+a1oHisJ
KEpEVK62jiogvgrPL2BS1a+rkks9MEnW9IGnrwz2U9VkJaUX1jxQ4IENgc4YalD2P+nhvN75egPH
9YFkZQUeZKl6XAU06hbipZ9Jw90V7OgDslZd6ioEpTnOlDuwcuD8Ay27390SPqsBGzt7mLwDDbjf
mivctuW7lUNUmViUwm8eSRQnJpNQ9AtYnfBLwLIx75eUPFaIjDuyjEP3gXdtlrsZ4B4LVKHvd5SA
LEpbv39+FNlo6EN6kbMk0CtgiYjig1bw578D18Lw+xekWgIYBXXMRVq4UvjEzYKyyJ/punV8046R
SlQX+emnviNeh1oRLc+HE60AjJ9XVsSvDly8lmuEgKZkI/DSGnp6STC91+thzG2gQ5h+QuP6aME+
Zr3tb/WX8V4atUk2cr04NN9R5TuDEa5iD5d+wOi4pUHa2EdIsZ2ZdMlxzeyaxTH7w/VD32rzoaz8
s531Wa8R5o0RjNYEwdM6sbBbu5j8ztL9yimMMaUWZShn3CLU6CX8/4Jo8HhfjfqfnjTeh/hTyju6
F9P+Tau5SAMoZa5tj/MaKyOBd0K1Em5O9SmaYAG6tFiFtjOCBNAeSYTFsAl5v4tDYyzqRVFVVTUT
Gnfd0v8+Ko3upt52Ne3K3noyuA7hVKr4S4K4fiCNapEIytjuOUP9OuaW00MX5XxsfJmbEB2FOnZx
GJSyx3/MEpZWUx0wQwxHK3M3v4jWL+m3mL8P6xmnGAzuNZ0QTSigbiSnQ0RJtgDy//Io+xAzlX9p
2CTx7i5f09uIWjkV4hgybr7eqcjkvhYHvSrFAaRtc2hmCiEzuBQ9OqORG5nMi/SLD1sklZekhi8m
wNhaOGXtp1kpsUm6X0NUgQd6GfDXB1Qf1VFPfEG4GHVKJakCpM2tYJ6I1TAiw/ADjB+t5cNzIYrY
OMnhazPn0gChfHhzl3Ertt12SM1v2+HxVN5Bj/8rcHpambGqiJcdv3Lx8l4lSIKqhkJH9Rgc+ICX
EM6qi/wgdrJ655HP8bQpirgdR05uXSnwuBDEC4O+16L4lPGiu+VpRBOtI91YUocc5Svqu223D1za
JGs/ueQUXXUTDY6qx2sMtaIBgVAs5TFPBhc/5pkyeQNJFaaicf63dpZo2x8hldSlnphF1E+uLpgC
euKYAdIm8BQb8UK8JoyRZRIDNMqS55XOQhkjbMdmQqE17Ai16smPQuF02Zu9YO2FwCP+5lVcwAHk
yH0xYg6iRn4JY/b6VPKwjqJSvzkZT7IpaHooIwjdXfmydWCXGVy0PCDheVDfcQbMV9SfkhiD7bQq
ZVjzmMKR4bzY9IjeGTliglVt+bU+RZ8FtODMHzXiakfVsEuMsXqvV2XQuSTx/HfcBEllH7BJxWBG
FnpTDQrumpUxIMEdoyCUrz9L0LOfj/mtNKo4BU8j5ejmOVEcGvDx3F5Qii5M+ZhNvzsmPVTt+o7U
4ezLZAsHYi6IQUeLClfnRFV3/sDKpUcxZRosbniTVNQofrADgM3WHwiibDxtVPPYjUqI10mxXPg1
/GWqbKhdsRLjxOHUpxCll3PMO9bCz5b4m/uvBPOQM3WKLyorgzyiBcEQAT/SCfW5WRcwtNWhBG1H
QrRK6NgcJcQMvoBWFRCCCH9Bm5AP2PuyrXOdV6rXixs8HnJkhZhj7rB9eAFi3kIx9PYjJWCw9iUg
G5m/w42Y3mxumrjU4S4jUx/xUJx3jPCC6a9YHMLSFqpon1dxUmwNcMEqkyT8S1LzVCoAWhH4JDGE
OcXbGIkDDkJCTeyLs2Y559WSy4ztwF4HvIz++4mz2ruVpQFDXn6m0zq4M9ZRZQ+I16VCOr97QtFO
KqR0j9UPWAzW/065R/LAycbjLSSwZya1ft+M8mnhMgSwftbaulCrUWrLZaSJPMuJSArr5AElQoVU
tm0VncoFevEn3ys/ycmX4H7TedngFNv9MoIWwD3QmRgDOg6+8TpwnXZdZh5M5TYYwN9KY9SZ1id9
48D6MNU4jcGxx4f6NpQNJ7JOnBXssJWyZpKpr4fbpzPZtl/KtLWd3IUM+oQPBer8F71VdX/Vu1xq
pEBMos0I51u9QM4moPq5a6IjrxeZFTv34kmOvteFuIrevBuHgVMQtiaatl/7oPBlzdJkLl7SCP6I
g8Wjn7G/risK4R6efAroVoM4ob9fl2+dMYHhK9DpmDCK4PkR58krJdN1e7dYEcLrexseG8VYBUEt
2tf1rwEfxMnWiqaxsoUN7PiVllvic5jFHBAS0kJbm2EGdC5cxjGXdiJOPI2aQ2zwocdzrOTDEcPI
/YZsGwLzelvVI3SFEy8jKqp72Y3ME1Qj+uoauc/j9e9CRH/mD8YbgORmauORYQO8/dE3Frh5q0+3
eDbKf3yLYSdWlLgTeLb7O1J2XSjg+w4QOQvpV8kOj3bAEMnH7B3TGHKnsqBcn9T/XKRiFGg+eo9k
i6nlJTg6IsGI1BaueN7mZ+qfzhODOSZUn2WCnngNreg/yk4bQGMxcETRBKq7GGt3DfuQwZsz2lmY
cSqYqZoDfGTT/RbSEilLDwBaJHdrbY1aGYVUJrt0IZUDNTKwgawhDXUvmrXrGubnt2qNfhCzw0tn
7ijXZ60d0n10hxyDH2gJp2bpkB/7hydnukX4uf6YD902O7U4cF2wG2BolTEOEL65MjFnOAjeWGBl
1HWtSp9ZgBugoZeZTfYZ2yJLbPaNIUFl2fV88c/1u+uxFFHgDLSjeGZ3qBUfLiRaZ+0n7zZ0QfNk
lPG5162i4WzQ1X2lRRhPGRgSyyf82rh1rnOUbNMcx39WjkwUSwGP7qr2tN/WF370nkXjRaAcpv9N
/9RTXyUUUiq17RnHBrfsx2S1QgpyAXv00LcfGu+bLe0++do0JPteYe7KoeE5sosNdwLt2WQl4imu
sDvNo128vmUJe5SuiA2TEegD+ps9n/Se7uqrqY2NVIHRfhGdSeR+pkUS5W1VsUiPgezQLdHldME9
vyN7dRsfpbsJ6OZRyhp9LhF+npl9MhI11flofOpcZKzbiYj8i3rukPYhzn2Unk8gHx3nNLLrUQTR
WjN7dFb49y8x0NfyO1a6l8OZQdr4BcRrS4jC2TPiGrogI2JejPxLuRVyl78Y6xru0ia9PpgZldQR
mZdgDjuFx85rEeaWUYiEpDeoET5JLBgggNC412yCcUjQjOzHidckCqf3HDi2qPHfhfRoyPFivTw5
RRg5Kit4kdhIIz/+UZrbTdW70IjAmr/TNId9nl3h0SyPtj1GpqWe0HJh1vfNFhMJkiLm0hSNyZTR
w/UagvmG3hDdlorNfpwOBZPdEfw8dk84G/V9Z4ns1T+iKwWhY3gLLofp/y8l+Q1lSctjYWtkEuKg
bvZibKHS/HdDIACKZYldVSIjdMt8w7/T3TSSZW78ZCtYsvIAiSn9g/bZx8gIhulZNfzwjUE5rtLj
KDdOwobCS0LZgLA6tMGZiEX3PbWnErH+MzLRebCgbRwPi+KVhmPwxxqPJhUpWJnm0I1MiysgubU+
hWNmTBFE2yD0LPkfmdAk4mkbmnv3aGDMNVXnYXBlP6mZVIfQysQLxaVpTisEYzGRzwvjqNOtSZXK
CW3bLYOEP+5Zns6/IbiRshmvI3fjrPY7tuFg+d9Bq/PEVKnru0KHAdDuiDQXLOCOmXDrYSfhR61f
Y1YTG2n7qd3JFJctjUB9XPpc2t93b0PI75fJ6wLmj2PAim4ZgcX6PyKMgygZlI1cN6cS9Up/smMk
SFUxGSrqlTtH4Xz8k0DLh+djcxQOglV6lh/daX5Blczbub2uDBK5b5GCV+a9QWMkYOSZEkllVgGY
kqv8w7NsEg13MlIJdL/qR26Ia9KnNnrcxRkuQyPb68j4SGpsTIzLVptlTCvNDm0QmCmmEFgkP4Vt
2QavE8bSG+g9SN2sbmvZLvW7z6GQElUY6r9UmLRBAn1IJgFQOj3ggmn1lxAksU9d37N0kGk9cYPW
cwh2Bhh2ZmBEMJSUxH+lzE8LMweSo46HIZJjy/Ew3c1SdM6geSyyKv2nAtRyNQiFE7D/nAskhheC
RaJoJgF2/TRgc05oKdwDtAUokRaYrzFRFx9hnWeeo07Ob9/PaXgabbm47HGCf2juCKL9RC8ofiZx
WBP7qJCzOxtEoMBHx7RgXoTvu/AmRpy3gA7Yp3ohzhEtrzGJ6i6zdZqNLU2jbc3GEX+kbwfIck02
xCCWZSPpvsvADJilCCX5ogiNNB8YaCg+mTEmiLXc4OGBeN0fYV3ZSnEL5SmMiSda7edGcYWR7S3R
HlJKi0nHdGxm55ILV/yRCvM6xXCnZEocEUFa9ERB23gyrzuAC/Lec+lZvZqL8aAPttpM7apB7kFH
0BXeJp7NdsvuSnqjCH7MWGX20zm0E3E7qVYg/4gCyQzScPbMZAB/R5mP/uw3eLfpROrKMnflbBT7
GryGyo3W8rWRKMbxHvynjWUkFTLwHKxfCZT4zq/X48ABq+jhc5KNAWPBYcWiQYAbYCFkK4IrHxV9
AJHhWo5/fCur9c4yYtslJyYEtc4wQ1zG7TMEf5fsyYwNbP3aO2jJ4o2EhWGqjnyhwKbEvntEgOos
T9/RAJnn6TiyL7mzZrSLzCTpmcg74xnvlc3Wa2Lqg99OTm1v1leKAgw+K7GfWkUwRGj3FJHO9bhb
OkMzz6P5Us8FXpCjplInNhExZUFpHmXaBclRUQ2YmZPzf6wolsOi9Jh1397lL0VULIv0P27J81dh
LlYx+cXDZ14EgnKur3sqKEQetdX4PTvuYE/2MS3eB0/wjMyVxiA71r8E0/JTw6b/8i8lzHoKFldm
EiHASQtDm3T6Z86R0EZeo8BqgSUjpBuAmtNrsHAb1B8FbVPjVCvI1WGRadr8REmGEmN7rwAMBCLo
sSYH2LT/Y58i9kYeHVmv1QZuO4Jr6TxZmaSOoide050p0kKVXt0xdJcebScCMAfj3d9jpoIlWhpw
ZogP0Wmp78UsdF6w7xZj/FRGc8lwggAYzOCY4S5+20unwhKY+3qvUEKntTVexISTum8wjlZ6X6Hw
DHiDWn4uU2cDHdizESNDbq3G6In/AlKbr+p7oi+ddjaQdYOB2GoEGOGuV+g6II/MBlYm1QhC9SB0
AbGKxfqyu4e4d7w6V6rAhSqWlkXrJxfLAD6f0Gw8r/+DikJMzfmdnPF+rcQW1NTpAcjuUrqgyAbd
inVXIUV1A9gbhC0aSsrcNHikjnXN0zGxDcjA5UWc3dD/Hks657c/t6M6VsEwnLqiYYEhTuQBVKZW
dRha1OFtZeJKrnvWsADRn5+7hxUacEltMmw+RbTSvKXNSdp6Ra+J5IJGpsll7qH1IdNo55w6xIe3
Gbbb1K7zSZvlqOspkfyfjAwkMRDlyl3omAhuMTmzNHkwA14D8hH7324AP4cUC6uvzkr5NSE0dHM+
9kbWvf5OIBPumNd981hPk7ge95bhJyFU0ZVCjrf01UEWq66G4l8YzR5Tvv+RFLpzT4Dvgf2r1kgu
cJgcCe7x+r2kuzFd6hWhPCyFtWuHeKiQg0FPzNFd80Sa0ZT897ppFzy1PhV0ofkuvG+9GW5jqFQN
k+1EFhV0iIVLbcmeNJ6Ws2c9wCzo3WGvERAWKsgBHkG2LFPyKeDpJH8Cb//xhfEM+aLHJ3lSwFkk
2ITUJKMe5TM859nQt4uCjkiOOdFMCAZTWVP9ZYRYNYzDlNF1u7AkXtQNtHScEo8e3UF6ZT9ybJFv
CMi8ftLZtPcHbkqhyLAq/ls/Egu4WnTJvVGAlnbHIGS6l9lsNyXaZZSW2sQJOLTlIujr58c7sqbn
BqYCc2V/zzwHcCfzhgJ20rMbrBXyaK4jwUAE1bmH0qJsBpxaK3UBj07la2A0Y46MGkzRRmZ8/xlG
dF+zh9KAhuGZyizUaO1MNcJUj528m5P/KLrKwQflSqWJ/ZDKghkd+9DCnHrZXiR7h4Wod4ncDOiA
DCxQ+OtW8mAdxEMEwYFPMb/lZKkqVD3yFgwA1pZzj+hddocIzUX3O2CBHcO1Xny3I5f3wvmvUukc
0FjC6C1ZsH2AgFjqWm59QLlkaOB4DrtnNx8c4I3DWv0GUL0EJwJqROoMXIaGshV+J/VeNPFnzAGh
fSUnDrakei9O91EgTTqUIOIELf86e+e7gKKIq9Nui69EGSYg5Xhe0rclQ1zhiNYpJ0u9K9K+t54S
Sp9hx6alsQAuMGwAzASv+lqXTEvX3G6kwBVo3KOD9gxbK+j6yVJ/VYGCgUVPqi/aRxpgBuuT1uhn
5ngg3KR69EoQvyjK05IKvKQOrDLwFmuQTfgnFIFCr7dOaZ7Fqit2zD2hLM2JT2MHhuyTPXnLU3vS
XVT+AItPa8RMrNlKCHeDP2rDXD+poDygvul0WPhnRBmlcn8LCqZsshO8QXSwyVOD5P6bOba+Oitz
YYNoUrdJdSm61SpKZBim9OFkxIaa8c5UfGgJsvlf6HpN2lC/+Ug94oF258jHwdyE70CDrGrbQwoT
YumHJYX/YsWCi+Hx1ddQVAPkl+Hch2d89btAQKdj1L2viuav4Spi0AFWaIgmKgIgmrkDXXZ3ihZK
1S5oKx4sqjQkQi3KUm/sAU+o4AKmxy6aLT5il9ZMw61zAXeRPeWE24l2Y/hka2khn3LBS5a2mLwq
iOfnS+NYymgSbSUPp+H20HwYRUEr8UEQAqv10KmxHI2mo+E5th3NjW1EL7b8nhYy1vRNaPiCA7N2
csNEB37X/n5YXazopWlhqIxVw2n95/VdGnaQjSrYATuxr0vDoriknOvljq0azQpiUquIk5Lv0lpy
J4owx2mo34MMgQwQv2gTv1gcFiA4UxruoZ54LTcSP0Kk5zHHp9XY5dEq6w4FIzcVsQb8I6GkRRQU
Z9UxQSdjUtIh47iZrDfECMbuxvlo46evrGiSK7dAoTHs99Za1VnNsdDnrssG88odxxOq06lSN652
LFdhIThjbDTeILBI4wRGyoltS8eaDfmHcCnWRlTW3/7x9i+fxaDeqkiTYngjlRENF2xP55eXYUqM
Wa0YsjsTtBz59eM+BT5U7rw+l2zLImkunnBs10nVozzY2Vrbo+sE91UxX4wt/BJdfVOSwystdrXI
NlOlXFDMLofWe9qab1jO509IeYBYzyXxekqbfLhOvR32Q2wsR3XjU1NLXf6otpBdYk59YyCjXtu3
bING4pSWOc6EjYyUPR9syleiWi/8xCODY8snppwK8TTx3zvuIb2x9uq/LalbmFWmfgpLMmlFdzW0
w3UOs6yydEc9aOnCUef57BgJrtNE3xrpsJGTiS+OfOJ2gaJzYXp/70DfD50n2PClzJ4bcO3wiEpP
4JrTbI0DamZVIjfKW7tV07ncDtAtsbtKbwuFXNfPv3W1quDhO5dXxk5XZxngwgRTj8tPfxAikEgN
d2Q5ZIOdq1xdjFYYd6MLkofgeChp2DvvTkTXQhOomwU/3nk9fN9EuN+p9mCELHw9BNOQdQ9CzHnN
jLaA1wDvydtJMrTuEbHQZ1od+AF3Fxqf6QZxyVkwXFSNqS0+pp3nA3dAilmgSUoRAb4sm8yKeWI9
L6TjTwwiGlgUaM2+8+Fv0Mc44F5x4HCdHug2cV+zdo6SCz0UmuDt1+dvD4jDqMnRPCJxYTlZ9eYA
Ah6BKarRGwJUYCNXq86WFEx7ahdLItvbqM+SLG7bqSluI455U4ZbpxGuCUTluox2YC76T6kXGIAa
q74YPm1nIkxOzOj0O+9LjTiGiD9oerxki84VQ3fS9FvQ52h9JbdaBxiNDUhGVh+rHddJLPway4+Z
kzJyxRnvkfcPuqCKY08viHs2QVq+fO+U5DGSAXahz9drfgv/tZtITx+fDIw3lc7QAiQo6Kk1dWXD
fdmBLG9jaYlZh38iUTj1GV3BvvWF0Ntu9CU1dLBQUz8otpefEdj3i0xcSesyvZAgwRP0D/VnFVgI
TC9sKZayLBtOyLYPOSDbdgaNOHzmD+J4DoBB2/ZkEyVFMj3czEzIF0XnIpzsUV4dPjSpof+R7b6Y
BpjWfn/AVV+9NlHWok3lZQFcPfPRqorOWRWjCoPeUgeXdR/7Nu8Fxr5+fH1dPr9pWyJYmCi7NlKg
zKChyyuivst/XBK9W5Fcu68T+RYON6PKHoPBf/fSIrTv1NLmQClcBqyqecDHYbVIcdhqpy76wP87
xarX+MYY8IfTZofwGgDndHZ9TTQF1YfdObFZCoBYYymKPyIiXT2q2QJaluv9OuaP3tB2j3U+Z5n4
NhxLVY+RYRjyrYAIxyLjxqwnonqwC4cEkDZErhGD3Xk3JrE8DhXeWeslFaYkkYAWKWfjAmZBz1Cl
kk1vM5/fjEM7Pkt4lftC+OMkVPemhvVMi/2UwCezC9LpiF7Ydq+KXranVeAHaYk2E2qMtZUCX4ti
ZMMHjmcSkXNDCpLDG8AupRYIDsJeAAWkbMuPZ3vRuruSKBrg/sHjJG8Ks5qYwg3nwLRjEbz/NojW
/l5AMA+c8eWB4yuzawBj7czT+SX7INQlKjfwS4VjjZcUweE36tst0mlaCaBvwGAU3uJwnHO44uwr
EqB4nHlG4jXU+k6Eiu2HxCfvG3IjhCdnUMWXkKfWd2KhII0wm//J9l2cwcSLnTyDal8sQ5zZynpe
0WLWe6qfRA3rnmW9ckq28/B3vihf+LpC4FzZrmlndLObo2XRWRnKD/hG8oZHpyuFA+D+tnBH9igP
DjdSRg1nFc6GxZMEVlIUqW9xw/8EH9mxs2CtokaU3eUDNUJ+ty8GOotIM8+wJmvazoW3y/FKnG2R
xYLeWRh4GiYVIrc/9nrkuydE5LFy23pfYMujfqYZ7vOZ+SRzf4/cQKsPMm2OiBqmiiXjUVLkXK8O
R58LUeA12PNAgts/5V/BKpCIfcY0UlRwstNOWu7h6pzU3NbRcbDcbNVrXAtZDuB0b1Kq5WefH7qt
J2mJALYQ+ElQvWY93Y4aRHJyqqkrcGmRnUW5zGhyf4H8ilsUVdSihodyVU5zRPSo+T1n+JYMEKFV
aE9tZIapN9O/L6+VuhAb6A0DthwAeAsxEC29oYqRhKTWU7dJtJWFY/nzevT41osj1W6NFhWSGp+o
Ou617GaybbDmxoJlTJ1ZsWGLnQBtSsl2lm4ZU4K+jr2cNg+jrVQuX9Jus8FTv2kQNIudIjfj6vqv
jRAigcQHrq+F9Z55RD4b4LarrO0LKKPjeLYY2n4L6VA2gsz+QBJZmT/bUADLdwMluAokHRzJhhQ9
yTic7KXLFbmEA83NrBti9rWWgw6wOSZ7oqB1yNCRno5J0Ky4y6DuHR19uZ2aWrV7IVhd0eY6V5og
p93qittkC12ruzrbbjuOgJz8zVUvozJlRP9JGmb2AHHwS6UD6LoodAtAn1bwEuccryKphh2I/Cve
N4FaQjczeKrEdPkM8zjJ1dH8dJ1z0IIO2vEJ7/BJMsckUAfYPjCnjmR5FkUH4arz4+TMadc1+I8+
jpMOwZ/hrixLhst2f9aZWlf0wQ0L2y3+qz4ILjdoh51MU2s82kWnQjThAip2E4HA65sQjygJnUFf
l097R4dyW7ZEcT+D7QDmv5w4NwfeKz2xkue9OSqlLu3AoHQHUT+WAvJEq6gMCwAbWOjmaWNW2lhI
t1VqwSgS2+xiYv0sfXTTRp6k5uWLfJWK1Z2FHsyA8MxhRuWJ16daYH4+B7MIXO6Brru6tHS7+7K1
RGxGgqbeIGadPV9tvDh79NfzXcfdpRTXajYBqkDMOJSUtJn9mWYbxjqzTX4xpxaJIm+gdt/HJNL4
Bs6sZe8JOz2J+p94RhqipiZVuRJQeugNh7WeLg7nTtANw8Qp04eSxk8BMhzxZ+5NkzaGtmiBcWgr
Zw0J94p7XrgoHonbRTX6QgXOgFSpFlYRbjxE+lb+bO0HppxXatztQNDOfvzrwnGr0XKkpCd4WgX2
Is+Jm8ZYn+K/E9u1u1Y6XpeeHhCPfkNtd8yetSiC9yGFrghtOpUdJ4GP75aRTBb4XcI3xST9s86Q
gUijoegH1UDFqdh3zo9N9/iqitB+/OzkInUja5thTJ4rI2b3yPLgfuop8BN4K9AFgACuYS4d5B0z
t1++OrGa+tkO+2jXtOCTCg3MqpqnWVMuTwVDDXgwr9yWN9jGj66lfXGeOrxnybEmKt4IEaX/rs37
iXhIDz+FOoGw2q/Tdwjq7bryStOR9swozD9fDSzU5a25lnYkddCI30yQnicVq88yhzEDI9f0FsDP
GWpXs0Pj6Qdz0BAlYCirpEJs6YC3IQYiW+K2iRHBBKu6KSPbvCWUp+bLmtgBhhQfOqvvFBdLJXXl
U8RsGet0cWC+FbNHrIquTz/jpg5Q7NIQUYwzHthAqqOUJL9HW4CiiSSwTYvx18SkJRbUOzVYc5CT
dI0eZomQw1aIbqQMJhz4y8bYc4KhkFYdjBVHoYKjB/IAgDCWFDnPaV/fxA9PqPDql7hATBsjC0oE
peqW8xnJ+Y7qAUQZje2NgGfTolwY0NB6/OOsNRCPklJiMzZ11pdksqv7pW6BnmqR2H+T3ZKHbk8h
paC9hSX0+Jp+umNGjAXRv7JRwjmmziOR0bch8R0qAa4IP4lBh8LKFaKCSDYQmMMUAC3FdcVsdAwt
0KdsnTutnJswgHgbQizti2pQB/ruhmL6s7C6KQeYgsGhVHjE59MP1WN6mDc/d4A41ppjNxHfAYkL
fsUsz5e0lljADmt2PQoMO3a+UYvxH4cPep+98DqMRdXsLPPsCfPZnTOgPv8KZTFPcNhTG9pxqAKb
O2tq/z+K6c7T29Iw6SufIiEdLPr3ifXpX+n6lKCaB64gaKbywo3Oh9zqjvqiStEdCNnJJtRX7OW8
sNeys3R8ypdc/NhFlM0PDguqE/SC+d6IrYoLRbyI1HEyJvl6AYgnLJTMzWj4oG2N152cQBeescmk
wVM1KjvjJgTiNhcfEZhceUt4g2f2SCGx6QK9voconna6YF1zTrc2JDQX1piX1fELyqaX+2xHvP+t
Le6/4PkYgPQMCX+JotZoEUJRin/gY6Vw2tzA5ntnBmlpX6+YZ/8rSVP/aRxlpHuokBzkQBv8oB3t
S3tcVS/soNaZr9MR+mr3dP7QBo/H7asHQNVmA21nCJTTFL2sC58W+0nm8o/sNFZj6vhAZA5CbH6f
7Pq/4NUJDZujtfuC74xH5HflKNDRfk6x5wB6Y3kwA/YLFldhFfLPULepyFRejuiXlEfSeUolk82N
PWKcEmCfjHTuWEvxG5UMTi3OoY3rVDRvPAkxw4xLffBPc6EG+AMHkuytFJmq8V+1m1jJgsliojQM
zdEd90obkRwqW3Ppmp54mhrwK2JHGxRAd/Fwk0PlmeP5QS7imsk+R9CsM0umNcZHAT2/iPgOSqNI
MVcALnxU2OELBU+gsshsiFu43CbEyBVckIMhta0AVXn+Qoa2+fW14Z4UOA4Olj7chOxjukC6t2cY
wNtchUO/KFmq4Qukk0mIf4Y2pUBhYEVd+LTwCY9swKhbq9SzbloEwOMple/2zVMo+AQOHT0GbNZQ
4YJzCiRTTNBVM14WIRn0zwwwkO3Mvc1siJ0TM2YTlk+Iz5m1BnARavk7OL8EHgEdmshFO235TI2H
U3Y+NafGvv5yZRWjF1satCSNTa2FXRxpqhKMduJ0jCXAq7ex6JZmo1WpWXVZR8h7gI6KXfnfJhAK
KidqOgt21//n0903Qi4djDQ4+ZKKGVATjzImnucG7QtYfYO+ayIgTQ3k+aLnMgDes/Tdgj3un3Sp
t/oVWs0N0xrC94hHpVwzqynmcwBGOtV6NBWTf+OFzf325DRymw5Rt8IADBRN2EcJB5Ui1Ro29+ws
YxHY8Zze9NZv7C52qV3Kloqh8FG+TaTkwdNEWGxdjS2uGsLSzEH7nKKac3RLLiCq3V7FR8Ps3Q0A
ffthmxpWep5LA8ZNnHWRlLi9fq2EllD6PrUsXeKt8cyLYX8/9/OKjDdIpPBXfUgz/TZfT5VIScsL
/ZNzy6IVUA5MjYvSfINSD0R1j28HRYV5Adp6b+aZTdDsph1O4k8DhHzNbAmfs2ItcR/J4SRpcMmd
CUg36/meW6qFchI2w2+50fk7GuVayC0+hlvhpcSnfi3h3nxVeikElDQmzCvTZDwDzAFQXEx8ukam
gt/jCFvvv8nsuviAPCvNis6vl76v5yBva9V6b0BounFhOV8HAcpeoYJe7AWtJ8ur6WYbNOBCSwvC
wTM+DJA3Y5h9imi2O9cq0xI8xx3vlb4BtdMjUDf1CV3zIbUgQfz9zpj5Hg5Nq57xI5qKAVVuO4KN
XPta9d9EMsjDnB7nTrQ7My35e2q36CUJUzbcS8ykZiPppsPjc1VDm0r0NsvZQPerJlqU/lT8o+zd
oa0zqrX3j8gMISs+LVCJHrbgD2ZB2LZU1ViJ35jFn4RgaHEKfGOGxtJCmVXJwFVBQkB2jQCAWjp8
rW4eTsQTuvkM/SSaHZmH3w1bfNMP1DxmaL8pCM+Cvh2V1vZBLNjr/XFy5M6XpdFh5wVUkEH8zTM7
GTU2bREDM94X0UtemKch6E0wegrzpb984dBi75E2Hy2m+VN9yPrLEE5vbxUwltUb2ps6YGkRCLDi
U15RjDPvviRckaPUQ+HDEh4LvOSQDV7yaElESKdWyHMvjgQx/3A6g9Mi56MhlnkPmtTN87V16AUt
0WywOIOkjCGA1dT1bHVA+/ncmaHwNQEZiRAHALIBwSygRDs4P3RcdqghcS+Vr9MqbWkJlM4uAgDK
qvMXs+5Fxw4b9vvdreT0XeTMsYSFK5kBAa5RbgOck7dInlSnBl3J7YPcZW7aXgvLJd55Ckl9noVx
rNrgctxqjKJyKiKZtNSsHKKFXEY5YIvL2WwHM+KT3mE5Te1CVQRr2zeoHhBBlEUgDF66r0WT1+Lp
izpzVppUBIslV3rkOx5nn8z92W9MkCuhHdeo4G/gsYLbNJDmuuPSt4YsOP/eNcZ/daMjHadL2uPM
8SxSugkReNEu8TDiq5EV5gwBHfB927YBM9i9mumRBJNuHQ1f9dGF//H50vYMHFlTl1ECmZ2Ai3M3
OfCeC9NFEtQgaJY9SEkvPXc5Ia05BiQ1lZhqYY66KE+2H9o6gct+R2UO2en5sPqz0zNSQfNpXzNS
HjX/pf0i8qHifClnNhY8WVOkACWirjLMUXfDnr+Hrah1e5kn7YVGZmcFL3weqMIj4SvNapQRh8Nm
hfnPus+I7RSzUBZCi3m5yb/cevIVD/zc/AvbO2VvV4BB8cdwIefKXX9YoXGyIpgpxQE5meUumlze
VNngYn44gAaJ/Y7aZN3XaVuraiKCAPl0xbKGZN6oQmZucgGCrDdGB9SuXJl09pwe2PG8AOaSt++A
ow/W6tPrWcmrthx3rCBYnn/clY10aqI1eOHSj6sUZSZ6eLjCp7nsNIgZJefK2jUavUBdsLoGyjRp
nFcDODKWgsCbEGRrOMcRRf/gJn8JEQjUXFEsDNM0W+il1s5UxKfe2oNOIEt6TJkS8Jac3n29RKVM
whK/+1VhfG59Ozp86gmFuiU90evfIIZvYTjRvzj9t738r4B3pfWR1qsnaH85XalXBFxs/VtrCdXM
jdrOTu5UmpPPRP+O+EDeFpofRfL7mcnPVimQoRqClcDUU5kR9t+UqnomfaTC9K3mHI1451fudY69
UiYBChX5jWwowAWO4rak8M6VxIb8hotc2aIQdhR8URH5M/SV7r1zcBSuAku/W+wyev7JVsAdXLv5
U7+d+zAAk7BFKtTvlLBMTvDOwuShJlBHZ7DOqsixfnm452osmQpaXQhOx5mUGEV75OmJKLv7e3W5
TPQRHSMVVI3fnc80g7Sap9Z6LhF6PeypHKk46dxuEHgBbzUNg9jT9y24kCWeAlwPC/EN2FgZ4HOq
GC7WuzDdmAqpekgNSDVGzgziUsxGV3Jtsl2RXD6Dj3Z83B/7nWbQQf4PpGS5TCbOrghdHTLomqNV
7XJ+t8Uo11lgtK4CONzOQpaZRYXHaXvWfwSq19qqfzrL5vGnGPmk4h0M/IwIuZA23YnWSL6ciB8n
Jz1RsohLjm70x/4SxJvcqxNdXK8d+DikXbwqiV+JlU/M5FB6OXLPPPe3GOsa0+kJ8eyhHfuFzF2o
aQi+KJWx0pawcmjRe+723BJDKPCj2Le6iC5s917T/N75QuZxUEZn9MtE4F+hXRI0A7dFQlh0wSk4
4uMRqxk9RzHhhy7bIHP97WPnoDs/QD1DjIdKnQ//qKcRgqbKmVgiFiz0mLB8lut+yucrrg4jGMsD
3Kj3MAMOGnYIohv4+985l62FNQd0KMgeHQ4S+wS4JY0L4reHYDy12vaG8++Pv4UjD+vFDQCE7t5x
/w+Es9+WRprkKrx62FVFu0VNTJ8cIRONnZxCVQUpVBqDQktvzA3vNUNLvOK69RAKFIKHt7N7BVhX
JcuSjb5DozpjQ3Uu1MagCVVbd398IbFv3gF8NgizPv+XDlqsh3IAbugWCJVzG1dasSXvku8TrZtY
ruKmq10+kxfxrfOw/LdHyTlvfYpbARoi3oUYuw0Zgg0HgVnW3DItoneBXJSyeZ4x9YUVaYVbAlUf
FdSDHASzlaSuJTLOpgeK1Oqt5xakiPtrF4h2oaUVY9m+WhqtTNNU3JNGiSQzzBBPH3l0q/AJUBQa
kz7vmcDv29JewvWynKSylspos3L0Bt+pYkIuJFcSG/eoFz9Z6kS7u7d/K804Sspdeg1Nqyotcoa9
vMDHR9J9dFFcVKGcOk33N5fgYHO0Pd7f3J1w8FQ9Y701xdkuUEXiZztw3KHTt11MiXXcaxcEnuiS
X0sqDzqLKCiH6Bj/V1L5gt33MC84Cpcwu2IQ0OAoF2FSLjRhAT2bAkrDPfxKud/oLNjIZC/7c3SW
UEDvGNhyJwkUKN2X9l3nsbeos3he6lIZnL+Z+o1q39aFkD4HZZk4bCglf+Pq5voXfDQRXvA8jBdr
fXgymEf1N+wDOWD1Q4cyelhh9v6Wxwr0ppwr3wRESfZJoLwp9d3ffB73nRKWEfzMS30TJ/jy3HwO
nq0i0uumshPMLBi3Tnwk/y6q2DS/UFBGdEtPYZGDxNQKmOtDqSKvhYgGxTID28CqpYOCeW8To6pt
dPJV6aIjZrYGscccL41VeGUwdnj3N+WAeG9Y8gZ3s7ZxRQWFzKxdMfqKsBY2HLrcO/F/dwEuLZob
5NeNdHRfMQ/9hd15b5Q72n62XVZJQHjHjSQHPh3ekbysENJmmxbVCZNnaejVAE3rMwxI35GHBIbI
1+PdV8GfKQOViTCVxga8pWirR/v1g8Sw6fCIfB4dmIcbTZpwYsN72+Zi0nL7ErBqas0JBFoIO0OZ
5FcIDmHfzAC/k90KfvCwdCR1cpGql9DNyKBtRiMEf8q8LdAk/26fBsvA6unqB7pz7Miz6OTJtfY2
pBXSxKrlw01XzyoL2H7HKFgGTpja58N6sBMfxINk8/XI1IT+2VRLlpUQb0yQS3IHwsnEXcmvDL01
X68VfkjxBZcOO810Y3S3Rp0pSYGADEb3BhNldUyY0VoCDK9nEqXGFI3ibkqb7yoaqeefAoYAQ44E
Z7LDNeCbejskd3UuRYvUGu0cUEmR4s4sTteeXOn9OsKI+Ejw3yjlJxxSWups1nk1NVsRF2wEkNHb
gGRGI7FGHhCR9AsPTr1go3TZmhQeoAJleazy/wHUpDZfAtfnPcMcb026FVyUrBNo1DW8riJjO9/7
lEBkcSarafm01T7vXvM3qUvaRFjamon5fe/uoeLF6kOXI6lbbmvrDjPj0Nc7d3k7gFmSqCROvBLq
QsAJnuCwxFiz8TFktOxlhY0FGNn9sKfGuj4JdzU+u+8a5iusg+vPbmVBimfFSkzwT2L9u53ZytWm
6w2nMez8ck/uIswhKKyH6/op1ZUzzTPai/GVBzvZArLCbxkHSLKT48YLN4aWmyTsMw+JgmOXePcC
oLWYiEJ2l75NHepI9+3vafjq9IcOLdZua/v4Skc3ZmPwSd5bJ0KgzgxzVlua26G+h1xyXLexajAu
L/l2lAfb9xk1EQbBQTptYaAn8HZjb/i6+pvtqPMWsVB8JoGXSOct+uprmY1/SuM+14DraxKax+Lo
a+e1WSRuVO8XLEgMqoYuFb6GbFdA0py7iZVZBWEwodIU7TgWA6g7K05uLn/6ExwAP+bTmJLtGWN8
ImXIzKFlREPVFQ9D7odZ9u3729+cmQTVCmomXi2xrVx824tV4XVCuoRMF9a/NfgmsiTTyxxFp5oR
oZD6bTBkxQ/XV7ryWxl6V5SeCUFW5bD32Awnms4NWLlTEZUgZ705biMIkK8EjanRpt87oHw4UpHD
ceaA0A15Cj8DehhQ1NXFGRVeA5uDzo2iGeVaY9ueSfPEw/tmJCn5PfBxiREqAW+SMk4J3nWOM2aR
CQFXyaLZBlEsr9R8w9K9B2uRjZJTwn9r51nfEwsWAcYQBR0oyQQkfb1rOgkSpfqmEJa00nACIy52
UfdyLq+EtjiCRQtYc09Azuo9+3Ulgedz1FWCU2RHF2pwlp7puyj8Dw0fThnCvr5TxemRVLA0e3A5
pFBAYRFFEgDuhZTfL06H59pHqH9g1RNXn6Ff9+zcTvn8dZQG0uhcx5OXDYyTlB6upbfRx1w6+RZ3
631cvXiEm2PUNIE6zoS9iXS7GGToezxuKzlqA3y81MGZd/YncFxBKnuCexet+ptKQxHJ15fKTPXe
pAIPI3WOaAsD42EF2ywairyjvIzsr2jtPttEQIfY8ntF6H5t49XZjqxc5AOKTes6HyM8Y5Wd0vET
rrvrSV0SN+qJzld9Ht04qVfh86DlCiksD9VD+9/uUjGOvXqMYxZUyQ0qXOMv/nSF4l7opHbXTG+R
uzGL1p9sMtZni596ZGCmc0WXiFm1uz0Od7mg/Sz/sg5jzTlqD2NiZ9fYd6HRQKMluK7ojWNu2IyF
LQtFEU4Bx3CoBr7GnLf24Cmf7B1a70RJWuf1zS3Sj3CUk1v5khDrqyBLNmEftEByGWeka8saK61j
s0H5SUbAlwYh+c0Cw93QEsQnB7JmiGEXlCLWYEz5v3l8CtA3xLfvE6U4xadC1Ydh0o7TVodVSt8b
OTZC8C/8Ln1DyA4TqGEDSUIRPK0HLtrrS+pvO75cQNyt1H/+R64l4R9u7/saSNKPTxwWP5j1rLjB
Hu6RgFroKkARG0GPSfWoTHk99VHulgUwrFCbzMZTEBkJb4jHUSuMQyRw2ze3ZWt1cd9Wjw/HwsEe
ZoE/quj3CC+f9Myb6Iu3K7AMj+fbaxyipNhi9E1RQaoEuaYqVhED4GYi/lfWPEZ/AVjcXBO5NHvS
9/BV6KuYkL4iwJRJFTKvMlQkwJ/K68KKKsXej/Yu8wRA70EDhVXFdY3MRgZVBPVxF44+5jdU4IEY
IGe++PXRFqkMGJTST4MxbgWEkGVkAYAqVcwXbp8ADb4q/BIvPG2HA8Z1ZM9kMTQK7uxNEyPwSisR
oBNYEqoY7MbojZ0Yym3qSQYsAjTg6S7+BZQZxuFMq0IQUnHEHUdPCWwu+e1PSGclf02g2Ni++rQ7
S/b4d1u/OTGEf9WZcNrX9YZaCGbbHkgd3kcve9mwe5MZcijj4jZRhtah5GYfVTM2arM831Ix86OM
S00BzF0MSTvQJKum4SCP1Z4V+nZfxjuHAtVSdwLEPA2qbuD+EfY0MifgFDoPzmI710uGj3CPtxmz
6l36TzI1suKTbggYEJkl9tBqv+5KEjD1GjcUAR6bTvN7VeX5fBnF+zOUsEgtMnPzfJzgIbH8SF3Y
vo5ibb47PZcUWb6aaR3gHcxrRNVlbaTZHHeaRdBl4BbcjBziffz/67t6Z9meFEG55QzDBHPkoxos
9sh/906+Dw+YiR/DY4xsXzdVFpP8q0YbnBHcFdvfXzmwE+7+c9rYqfCcPLw9NYb/uZhPGrU+QRDC
MT4cUHOUOHVQUHLiWAnldyzGsoyVHcV+UyoQE9A1uFU3sddEmt70pcLrcxkIARRqymyunS4IASqs
GiYYgyLDnn4NUKpob+Bu2Y5ZO+hdr4rK8OORJxpDTsX2GcSUL1Xo1sHh+3Dvyf9zQaTEmKJ7AGAb
cwZD/+C39N2RXr47fwD91CgPK/N6b8cwE3/Vw1yQBqum4a009pjDlExuPiG6S3wIGA5DdySVCQB8
IgCaMXIihyDdy4vWsMq+mmdQN9G5Ha0KZmBpI0grvSsb4CoTzggl1Xg/Gv6G4f7JSvDepaBOmtcl
Bd3RhRy0Ba6Lcf4EKYhGknrlxKiD5J1BtMsrpy4HKGr9UEQJoVe8PVI7gVGAsCKuO4juCsJUwDzL
rCGOo192dvyPdT4k5lAFtF0/p9T7aGI7pzTNG/zopLXjAsz5XhRECakEf84uQTPmozqeO4ObsEFQ
6s9gOHb8hYBsVISlgTJWrAAD8DtaIcpQjhy1TtizAfVrFIv00C1nEHy2lIElCW+RnyFqTxF+4sNx
N3wT/fWA9ao9t5KlKeQpmDX5iej7Vy9UHaBnR1pAVF4YhAhkin/YMYZ7/YSKle1TbeN8bmJomM68
UwKOrveuRz2sfb+LKnaeKA5fVNgJjyXNA29JTKiBDpCSB8fNkfPSLaHsw2lKdAC5Zwr9dJTqYiYt
bQqrqeW9+l7AbYnZ4817ANRHhwCxWw9wKFoq7jvFU6iv9FSDKUmD/25hYNcAbDvOuEk5tBhU78fk
oh/g2CvZYmMExLGqjO7K3cNpNKF56QJ6AdMRK6zv1I7uTDv2Am+EBK1CYWkroBYxUwu/ekrJ3fYm
gRwaz/BmKGbwEO0kBWtEXvVnStXFMiIZUxn3axsemxcSFMUhIJmFrvimjB+5D3alE2fzXX26m2K+
jj3P8DoqdMx2YIkkQq+yilpfQi5394T67xmkqKetdzF9oMLaU+WWAs5yE05ZEsp8+7q2/6vGgt82
dcCu06zYJs/6+gGwjfy1O3N+XZN/mJo52tOapnpcbqEXATQIgT0SrsPuVvI0mFJaXCP+1bzfidbG
LxV0A1+N2zhpzRy9P2ea833g7lPiW7HTdDxtB0U9fok7icGH1hkF50Fr66IEKRelBybDgOPTOcVB
VShJ8LiP9yLZGwPcvZfM/ub4fes5pv6cHiU4XGGIWZ6TS06kBuoiKc9n/fre2vrf5MLHB2ilxhbV
a+jT/BvJGJxH3lQNRczl681o31rdvkKbbN6yk/2VjmMK/srU5BIp2HLfYRaPuIjGxu19619x5SOr
98i2gA8A0360EBNphSl1WLYjgSpObloomJzzzijetqmDaE/stw+e0wcuOFVxFTVk8fpsehF8YUme
+dgyR8WuhDmpTqX1o8t/g3F3X+ceIJhpYNFvdki8HuvDFtt9YfBvDfYxtSfQfvOIdFuauC9ozUCL
o+ByEf+ECLGD/WKRZ0TDDDKpgvV1Y8wmcMXr3R5faYYW9I8Sw1oBH5oLK7PoedtREXFPzpef/DIT
aP1RCn9mFSZLTs2USd7FnGdVZlhdz/Jvmp7wgUxIR/9aFlhX1kp32W4/Anxi0uJ+wZRPdFzWfXVw
+F6AKMieAXKA5lNgH5TOJPg7jEpDObzntwTaWFP4VPvM0OytAx6ljqJgxH/NiZG5bCAGz96/uYNl
6i+poJlq3QtMQPGOcKIYOVA4mImVmfnRgmdo7Fs6IRwr2LyoB4W8SCTmEodJdgpjVFIsd94G52nN
biRUtIuW71c4WNCqInJJKlqoUxIisA16swT2tbCqecU/tBFQyoBYNuk3kUtO7JtexWT33Cp60ojD
ENnWZPkDHgSGsduOAYiihgJ+gNKGBNjDWl7d6a6w8xJ0Sq4jZRyBpiUX4vZwNygMq3JWMaNxdJ7p
DbnBWZPGsbJF1e5U8SENYQrMCbQCkVognqLYeNMDLTtuo0gU4q4wdsFGrDBJRSn12TzSeqMkq5hc
5NqgRYj7dKxZyfC/pqx+2rRvqEI0F7l/l0OsgTx36B0rh2M7UURK4braKu00/JAdbvDSL6qkBIOt
8IW+ObqFerDo5Biq22u85MXBlyTjsztH17HGOvfi/JG9tidX+3s0kUN5sfkrMEw53MXjd7nclkFm
Lce0po2LdxokloQuZb773L/lWRjyHwWQ3D4dxv+xeaA7oGiNrY/WA4HnDyTqaVrSjf++vV63LLPb
m9oaglKQlOAFMPBVYXa1+6oLjK3UDhrnEvYRxnrs/vs2AQsC8qoc4k1fvB8ea9bipH/XrUir6mxc
H5IpVSdJ1cE8fhMAcOBl4ODGXiMAkPYkY6eJtfZNcTKKemKkLflgluLcGAXg9H86lS3wyxrjIsw7
f2jzFv8k3onSu7T6nCK9OSkLw8sXtV05Rz1L/7/P8Sp/5bSgVCK2GNwo6Usp8KA7UmtyNKO8AEtx
jfUPWq6tiofjPe/ZV6KRHM5pztuizVeICktCqgx0Zzz2166gaslp8ZGckHAMr5Mncm+XZGvQZVY8
XDHSvljUqbqNCrlrdnFQGY/Rq0pYRFYEjfI2yJQqWVpjxrINqZTVpIeTFj9a2D26rkvc69oBZ2Jt
rcfPU88OgMjxrW1Sld36fWtfZfSmTnPtxAL3uFQRpspSl8e70Hc6odmWclUKgV9imxH6sluEtpya
9NJVmMRDAfPD7sIfau85rSzNuIUhNuD5IqOIdLo7tLnR4Y5+Cxy0QjUW0YsYlniuvpA5G6ZGWio+
8iAVfH5VWK02BA8xEVtKzQsvHWT3OkH6ROCjV60+IkJtSXKkwzjK9W1Vf/P3npFooieaxcIWehsY
SdLWPfyrp1UeXgRD1GghuZcQ/zacDkeWFbADOu7f0TPLYW6911srsC3zWNxhfM3HivDKqPC/j9Mw
4SgkjV1pdpQJ+3mcOaBMC0epLzTur84ts4lLUeqh9S5gG6ftKKKyM9xDuIzDl24xdVzSmqyUkpgA
VSOpVBZKndLa2TofaeQm8IQoN/2xLNiQjFA+cFKd7+psN+ZSaOD/Ki5QchlzfuvPY/6TpK2ptPyh
B4J19qT4xs/fDSz2QcVZE6620Ft1cH/6afoiFoDml9KozSlyM8G4+M7smCwOr3an73XyxPrMSLeA
kSuxg1qCFOtDL2ShSrGvgRZ+45EJTXAQ+8GPBiBQi8EOxT4znqG4WYNFRj79Iu4gnNtk4DaWURVq
cO86JH/fLmvXF0J7IGReE3s83bXAm/ITdkjzoQ0Y1ILcFsUjTS7PwM2DX43+Lrqz+5J1CuG2HzdD
K/jPeKNru8Ymzuhn3sj1zqY+eztOHlaJ+EEZ/4gRmQ8vlGaFL40vBxNOITfsApKI77zxLQALhIJH
SQKVTVnnYT0YGxaHUWS0Lx6F675jhXYCAl8TMFaN1lDDhChot6aoMMad+4RVaJz0vC5FKgBNdpSn
aw+PQbqZwvzBFI/c01ySL++125QwEvUM5PGNlaUVHOk0O7OLswYlV27PtzkoTRneefQXFnhFJWxj
ywbfLX9/67miAdkrVKuAlwY18iHE0daF0GwVxJVf58Qcqa5K+mDCF/Guu21Bd/uQ86ZX8gGTMLA4
SW7j9owshEZePwon6FzuANG+BApDPZqrqjotmFc52cZCMcFBJdvN1Lyeu5vYb5jQ7987FKsV/zLX
qBUjw8jF620GbqapdRYc/JU7kx7u+ip7vXncJpy4ecM8cZun+geM+K3ZGsdihcyEfKrUyyliTekG
NgLlQSUkB1OPcWMa2jqoIvgF6buAxiW9jhUgePl0bJV8pc7GxrUttywFuHd2ngPFGN4cTeg7cN3K
/PWV9fPEMPyIkZcK3IgAgETGuLzxjxP/069HVmjNPpwNPIuFIxn5p8jCSFVVpmVw3pOSJA6JDrV9
v6Mc6vpGdepG5QLRhodsLBUWach6Qn8EporB/m/Sc9vEy2bpnbfxEWw4CuWog3NoBZg/UOjXyz1x
c6lkt0u7cJRCb0vcGkrdN7anauz0FLPMmpxpCGAXdcr9A6FHkaQkJ1A8XEDV23LNQC7AH2PzPhkm
zaAQEQ+umx4ZlMvOb9ncMgTuNdPql5kkErOgJUKnw6YyPIQLDXYH4t38ELpjf2l3qVgJdTaOh92K
CqQAUfqWhcSxiq72JKIbB7U5ogaXpeblMX/lcr2DGUs+m78ohAsY0wNJQWnjXv+hH7jlSLOVCSKP
B7GbVMttTnf4NSH65z3PAVLOif/d4pMaWSCtFD2TYaUzFHVi3/r+6IPrmejikJrX4teCzOvofDsg
Dis17SMh5CEhKN5oF27u2LJilmQPxq0Hg8eJhXvnHya/uU6hY9kkQ0dcI8CgtFUQdWgug0VEyugB
Q7oWanpb+WdyZhpeRRS3+A+gExjY8K/3/hE4vSPak6fFq6j69eK4C3a6FWuxOf0M71/wA42g24DF
eX3I5o8RfksLAvlqB9VXivh9AODHih2Sp3jAQt13szJ9L+D9ftm1meWmF1VFgFbNoF1s59xF40CV
p9J5l5hVoIlaApQ/8XllPMX7ucbiwYcfyQokftOphOktnDp9c9b08legFg9gonNDsZEyD5p6mFmP
qYX2TKDjSfOuORh2epOVQHo9yMGp8KYyjzYn202SoOTXwiDHU7Ep2IH7qn0znnFiPzAr0Wlo7UOF
uDHAeP34l7dca1BAYjxHSAvCPUe0ygeDKcWCY0SFlBZI2LpNDR+NhJOXTgXhGUQUCo2thfvTVQE7
5p9KnzpU8DvvhD1yARl3daBUMhF7fnjliWnmwiaXKYrkaC6csbR89zHBMNdXP+kacMYXgWG80m0s
AJZpPifWCy3Inh57rO1SiA/6KtkAnmoq8NeAdXjS1n0MlkbCGZl+qb+Gu179Lc9evUNnpMcrYlHH
hQBzKqbzjxnt9AJX0HcYMd2/49ihDuYhaqNDWl92hfN2SBhrR4Pm4vu3ENtJTW5wqa+ry7bqPvxL
XtFwLqmNdBE+Jq8m+m4AZzRZ6k3Zw68nZMsBGZqgn8LEA1FEn8RXebYDjYpz9d35pG8TVkMj+059
T+eRJ1wdf6N/kZCa0AVtQ2+3LjA10+rNH7ivmkjy0C+lBWQAGN5nEDZuj6C4kYLN0y2zv5bE6RPc
6Ef6Wrw4yh6MipFyi7ZwxXnwJFFzcV0zv/dOFDbxtNZ10vAWxR+XgSCiSiYPOlseMucSd/9tXE7a
9N96xZv541NhWuUbsYA66xWP9CJVK6tMt9L9fYFRCj3sG4K0NFQfTwwbOLOw+hN542vdHkmeCVm1
9mqIu5b5hBA55sCpfRvv2IaXxxIf7q7WtkA2iE7NwBkVQsRtXTY6u2saqRxT9XDoI/H+bYgdUBYv
veVWx4/eI6SYDmfBfrGxSN/rj7V1P20xgy3WX4WMjax0kSwhdFRozY0M6Tx4j/zsqh6YFSUNxoOG
13H2+p/yauAHw5Pnn26wJgllwD3mj8lOLkY3J20Rjjbr+5zAk+9FBh10/5+YYLlEopLTDS4hTMgr
0Tt5NymjcZmXBHPYE0txgWtsnPIVHBOd/9EHTuTgEK0KScAC6rV3Ftf0ZkSQz5kEA0YzSKCWOyum
fNnT79kIf8KOawQk+0ly2FmPhzjlWpdxa7Dtwy7g99jnsfXrIMioB9ttiiy4Z0ADr34mnRc/q92L
r57kasLLTBWsRcPAza7RP4QRMY1qEvZqLzYK2/5NUNdk4cqP3JPgnIPNxjlIOILJudWGAQOZjLkY
KZLzc/DEHJ6adNO+Msiv2BbVVB5pKKl8dFCAWR9gR7Sz+69NoI0pXR7P4opkhQJRgiZWAiVlUJlC
8Dm9AnjN3swf7uvbetL/7FZ7i4eDYT8nV99Pf31CTOvDNvFPT3T/9DOnH6CPxGceAlRYWikJPTwd
iYbWLnTa2b4GQlYSRiS97YU2ujfpWGRLISHgQymZWZQdqU6evpw0doofWzuQFVWDJL9Qayb+PmMA
iEWdgDPVSjw/WPQ8nE5G15pnbqXu+gY/rlwearA42IzUEz3cMyE/RYeHBoFngYp1YvOPrMPrvPp4
QTFhgytPhkkn5V2f+pYhvgOV6Doph/6j++Ycduf+EENPyCNOP5K1WqnWFT+fjeZDHJDBlTFe1sku
qKTMhBlDr8y7oPueenOiqrQqZpJVUYddJ5PtVeQOIlhdUdPXSUZVyDFiFjfY/6WzdNZOPprd57Ia
RNob9S3RjABP0Pjp5NJy+tCnwDoPa9sRntfwWKNAr0WYwfkkQx9f6z6ew8LG8+botqIZNR1v8aAt
VQ0VgP3trYuAXWN2gqQaWLPfTMOdUTk066ZplsU7+j717F6AgjN0775xaJ2sL5K2V3hyZ8BsIkHt
VWnRpOsGM1WsHbAkK7mAmKqK7IYaS+cswflYyzaEkzt1DZ0fCGTXTATfQ8EbPEVIMezkQgByjaC2
9cI6KSgP189N+levJ4EB4pjQsRg+JCGeIA01nyHuszjqwfOBNOX/tufVpBqXuPacZRNSW944Atuf
h9KDx+NRcFTwDddyhA9/LO+IcUdk1UaZ/nXtADR4Cc+FmtFnvWOdewKt4VuLez8YKh715xPbyH63
SimbnmTxuKruMpWL/1VGohAZ45l0898zx422t0c4e0V5vwTyC2sqtIJe08uMDL5IYGc+DQjfraXq
z6/LaC2DqpGGUN6QcDtVIsjjFDxE/5qSkBHtLHc78IZfl7BB3AGkswSX3f8aohKDeQfTS+L8EF8x
YfDZgf2W51C5s4/v0aly1TDO6Ey9ulyuqfG5DiVA7lYfLtipjdk+TJY1v2uIS5KVFvAJrDEe0obw
R2YLa0skYeG7Sq6+LL8s/d/E5r/e1KiXyyTc3IF5t1mfgdQmFEF7kwHp1GvHQyBOcgdLF1M6knjw
U7EeIfNjMS2R4KYIW/PAfZZIpwBctZ7BLyoIN+uuy9h9vaSctBihnSKb09m9HgvdxOI1S60vKQkL
e4ysVh+tezygFuN+zCEOWjg7hRa2oRECOrBkTHJrHhEl5nHcZ7Ty19RUVSvS0aBOMjc+4ANZo1wa
ynG7/8BZy8BhxkQvIRj3OX5Jt3FmTCctpiMmE6k29uE6ICwv4O3jQLK0ypKuEHjqrH9nVb+1r56e
RWpW24zl3LnFmsNd41lUIlfjH3TnSBwRBIZjpBYO6EHcr/9eek8nHH7c/lVa3rH9fwEP7811uGmw
5rpXcVGJA6HtXcUxPI9AHLMSe4olx/rLAGIPLhH6AXNZ8aGIRoly9AeTy2BRm9CVnFpEZ7OpULvf
MC2bN+Li/a0ew2C7cC3y4na7WtEGt/KaRY+wfLU9O1nCBnRlCOUsJhS2P75hSfLPwBQitz9UtN2t
uVwBnfjh1KXIGdPCIIuLcDs/8qK/b1Xn4WOJmbCyQf0AUuMcn1mEn3Jh+xiy0MsXjcS9jVVTA1p6
cMa4MiAH+ix8PDNC0A+dH3AyZoqBeI/P9so8CpBOotlWKYYNX9H18jx/yLUxHM2JJL0VAXiRr8tD
rfpFxZ3XdQxTm/TKDq5q0VNkctiLDOEDau0JYASqoDvLZFC9rWYEpR3WbM8QDj5CLnRYRovBa46+
qN4JO91iyxzAbVY+CQlVG8lVmJzYohQUlhLYmFA+i6ZQFkEtmSNACX6KcAwjL0yHP2zW3hXPs6v7
th5GMOUF6l6Uh05S1XEx8L1+dpqaPEvF5kYGQoL9vEqPBXWsALjLYs3D8RnzGN5R16DEvE2iFPrD
BjB94yz/lD5C7OfbN0z7R+8OemnFS/SQGn8J2IHNiKRskjgAaHmTmTMAHVVjkd578KuRElRmryur
67G9arWDzpDLohG072byq+zoyasA+LOpT1fsyGPC+Mrk/qTSNG2DRFugLKuSfVkkf5MSFnfH+unB
Q2se/fZBK+ejVA1K8dkuvrSlFMrhuwhPxX5eyLHtE1o8TJ0xykVq/fhzSTW6NtG5tVv89V713K/V
IPHhBlK3CHZJIXUaazjqJSwLMAU8MVya0FrPNDY/Y2vHpIlEtF72oLsjPMA5rYSAKTGwATOSetz9
lC0x0542xrpVaNmzq5d39GvKwOt45GFKaKW4OTNVBoCqKLMH8ZtWzexPiawOtHBKnckFntHVHMp3
/j1n/TB280VZQdyV8AuXvk/3zJB54wL8gDAUQOOpHl1VlTFnGm2evaWO5Tt1oKZjM1Y/JmHPr1ZD
74G1E60ufxi1tIZ++lf12QksTnSBZWaGdiW+seidVWip47FFzgc5JF6x1ePifXodutbB83B1DXyr
fJDiya0jhVUIfB2cq0whaKhsqp1nZ7h3Jhesxe05FRE125xGjE0g/GjpAtrEM3ctuaXiUglBtQ7v
5T9sot3tut4UtiRTQ3Ygjk6j3m0euEaYMW4SAgjELiU+zqpI/35HZTXCGFPGrNAGj7z8jGSb7bty
PtO9Y/ccLeq80l0ndNRffX2hPcETTI/S0HNCNRGmARdvFm0Xqy5FOoltje2ZHwwh2jJCAU1x54XX
AJQYjrPWgQCC9tDRzOwOmRE1wKlMqJl+WUVRMxRNaBZ1voI0EqX7pskPGsPieYeAh64yfssLxz9T
3v413jHzBacDzyVg+78/dHbTdKv1RQu41BRAAHtDg0relMLXfxo2ltSNvN10qGvDt/gTzHDOe0r+
9f9BbflhaLiiUvc+JquMHipoN/ZEO6WnzfoLIhTADk12+TnNz4xC83WOzgRufxrVW+VXmpx4eQ4F
shxcw2qoW/2XOHMeMVsW2b7dV62D/Rz2bQ1eCn8WnmVTu7clJvtvrN2TqA86ty9dbDJzYuat5DbQ
tNtfC1IvVPsRFM0Ubnoi6d8UnpxGTkhi7rWA5EwHzMhcMohOKMzCgkUaqVm7LUSKP0uJ9kvFunYc
25Upu53QRXnuXxez60OIDGR4lqpawpypqL73Zayrqdkr4mYvzqbwKwD3egfzN30hJSvWPIEry84J
7EPatilqgKTQQmDLZesaEVDTjbw0lQNzex3mz+KbUAUX0epYBdQixiYxhULmvxe+yaAR/Vg9Kc2Z
Q7Yf3sNJnWa7uJyg04jsSRWznJaXOWYqwl6z/olS4VH2PEHqJTgsqbQyFSJAjgl79nm5cFdr61Fl
SBOjiZhdhOD9P06Vn9byMqidkZsW+VTcaeIidI9s+fJsiBN/72EH6eL7PTXP+lDKYtHd5RK0o42h
4qNR7PItG1lxpvU7dMyOzphfYjN2Xc6BF4w5seQF/b6qAXBB5xZJofteojkCo1nxR6ynQD4fwd6C
BBwvHkb/Gv5PAjMOpz6bBCv4jPDUAgjcV6zis8GtX+156wBNLtuzsjyC/EzKTYoWXIcXvDBMuFBY
jngdPLyBLigpQuD9VipYA3gWoinxlJx97qcspqsEwQe6RGvCoNdIlB3A0u4NaOZfDRu+Z5ioq3qQ
7p0Gxj5hXYnOH7hPxLbYEHzH2dZttvAwrebVyMxcQCiCC9I5modghGpqY4FciW+9Z4krT57F8reD
Efa9S8aeF5ubN6CMS6xsPyp+gH8uudHH5+AnbVfWIdHGNFJYdzSkgxUfRLf3WNpuEKLcqswGIrIk
jbSMn4HJ3c8Kl4DBHPZebVBQxfqbNkYjREaAaSuz+3U9R+8eGvjHSR1Hwp4oH9uWmKPdu6RnjLk6
jPxKeO+LCrCLjDoB8ktu+xdJToQxvf3Y2S6cO3pKMwdK1lqTXI/E39u8xcjKTbuYDcVlPnpVh91I
aGcPZVAZR/8331YGwJ9KaF6HwZbrrp6lx5JxlZs7JxsfEck7JHTzXkaqMKFnBv0tMsfnL6EplrYy
VK4AKRgyb2Y4ayvsBeZEvBZLhrap+MCJqA0AcoCML4aeNooLENnC6wgcoyDjg3T65UASstCZ6EUt
YY5VvgcYxUYa5kShFDSTzeqmJl6+KdyQ6k91GvI+KqUWoIAFH/2eBeT4LVh0M9jE/hk2BzXni6vn
JPUf5gVtDbQDJA0xv61XJuC6th8ZzPaZFOsE6Sox+PhPEF1iIBUP0hQIEEKasBrT0kN6jSRVdTag
G6R/INgCs2NZcx+40jsP6hHZR2nD+fkIGkX1bsC1uK3IViNlfrXQp2M/2DN81J0MhgKKRBOUO/Mb
464/e9ljt34PgOOro5ovW0pILXo7pbD4XXrmjcZ5TkvPRgxUJdwZIkDnnU9hLH+IzAnLnS/zwGkO
xVvTeTQZtZEy3clWSR4XiK371+kd1LCjbV2TPEsOv9BeNjAamfWzloP95KzEYzz5/rjTnBduIHXb
hN8ugXsBJD0s085I+ngTb1ISMASkreBEn4Rf066q9+N1alxrbF8p5cnpzMsEt08uubDpJXbQAzVl
1STHfB/Q6gl4FtdT3M5mneSTp4vwneotzjwXjN8xRevR1ooWq/SfJgsx10FQyV94N4RpWwoNbTCb
/WpQNFhQh7ZJ2Cj+Skouczrm5vr90eHXtJHdtkkDX5CXGRgzI9CDWQjVlQ7xU+lXGxq9+BLeXDQL
e3+G7rG6uspEpLb29hCBEx3KkqPXTZRS29beWwd5NdbpQzPap8N32fnMA2k34gb+teOdXGF5JOUu
Tw0fKGNLFfECO6pzxYlf4+3rKWPb6xW9uBvQpIPrdRvU1ws0XgJd9Z958Yg/WLAQW0NMzj9tpbs3
nMJaHOW/dKqKaPtgg3A1G65ltnyLiUvjrLYZ0RvOuVvU4/wH1kD6uw+ihW2rgO9EuIwk6X9Vx6RN
rdIT2UpSEb6olyFTraV/EAnrZMTiNWSrFwTnYq6Z46hEzKc03YWmTmk1mIFx4u9UDFbn4pjWSAXP
Hz5VyWbreGsReHKMO4tkZPsFznGiBxZr+Qxq9rv3gIWUM69RhraCFkR4Rdz7aW+WsFPDq3ttsx3R
FfIajE4Ynm1AOgUVcDDVMDO02lSw4inE15FPfsR76okcUShq2SrFoskJL8GGFKKsP7pe9+d8mEcQ
gikhrAEgAyxpuRBuwin3T9RAj9aEC8EreZKERi11pokqUnRyuJaa5Lk5tOjFz7uLKcVivuTnvJs/
CLIi+i17aU2T+ywAV+2xQ61wYJAaI1SefMrnfL2bif3I5oQ95RV3uR6u1BX33yJLKUM7eOrqqBbB
i4IcN+ExYm/q39pa2gqJAq1NV1qAbgn7pccyglaFkj6e9wIW2yLC8XCouCKc4pwFoB9/1XJ/g6MS
FVkYzqpF1zQcjZgSUe6SpmetDKJ5yCSu5H4vp7gNtLLMrsfQU+MEv5/wkUk16HYSl6O58BMKKVXF
rCe0B+qDavoELAOnK2F+/1HH4TPuoL5CwEGS9xUVhMJ91H4eR0dq02Mo6Qy21om6YfG68kFBUabW
kHpx5xewA9d9eiF7gRzvBXXXy82ebGLSHtIWkRYpty6GV1+favSsQRjkEMBI+ir7SuxTw4ev7wCo
4Sc9oKJolQsNebqmzvWQdwNOeOs8TNDq4GLY2LIF+UlIQsrm9X7BQ2AkRGVtWAUDFBznhdvFYeon
42lN1aWPAFvmp5WQQuMMuhLx8e34HkJnI0LQvZ/7zX2X46cCaFZOdHmKmgVuqR1NDH3g5opBrQkS
WFd6v4T76pYJDCfprOssZSPosecf+oxFWP8/0ECpZIQIC92nmg4G/ex7C+B653YPUa+/xTOO9EYX
7dYe3KprAaR0onucaxPhWhZ6DwinBc8CurpvTcfZZ5/y/iH5zftv24MpqGXKzQO2hYldZ9ATn3Cs
5GChHOjPzPi1t7JZVLzujtZnctpw3wtJE4fab7pbVmpRDfODAUGUbnAvCV+ep82n7AkmZGWwx1OL
s4U03o+v2rtZpBv0LnAM9yzZ8YxDDpEcTvT5MUNRbcZLneVMvepMAW4VxFlWt5fCNI6S2CeMnZGV
tdGnSv5uTvErcALDMLgH6h0ejG3yDk+hU4W7++oJ6rh2UH+JsSm6UARRiI7mXQOigh/0YmuvDoho
3vomZW55tqiDLdmec0DT17LSjNXBCsvPv/7+v6ISMJ8fXxbX8RhdDOk5ieJC1CzibOQtQlxP0gCh
bPdXnw+VzfkYk5CcFR7lCDYyX6zvR4q/gnzN2yhQAjjQyE11Fy3FpRA3wtEfmE03eM+L5qDvsGlR
ulHIGuzsNpE8i2kFtVPfJ5tbcDwfVGo5FIP4liK2lA9inzBXStP1azTdRKXvj8nHFBRamUo3Ecfu
gjHnE+SrTACYDTqW9IlU/9snJ2d8gIt7SJK1jmAHAtKqyADNU8AKi8w9Iy2qmIP2886gWu7wyGJu
+X36jA57uHRb5wRQ1+2kUzBdC9vhKn6TQOs3IeK68oLaE+5gvO6atkbLdzBFlJXyfTbpahm6CMVK
ReTEElIlJ+BhDO6Rkx5qUqywIKbVwUtI7C6M0tMyHyX+zVE/QdIrGC75SI9QUGwlcFWSvndtR4aa
T0TGyBYRxZZf9Xz+KE/4Ob61lB8yf/o+BMpeirspFlw7tq346MKqOMIJBRhcuszfOFIPS36HzT75
EaSzlFtzuQ6L0TdlJlSG+aYNcJS59u5d+xGG/bOZP0RYAmv9X20zeoxHCePvXSEyz+zZgg7H/9LT
VxS1Y3VqHJVI31jJAPPfBYQFgw8hIbLYDelNtoj3QS1go6T4+XUwml0WHKBAZ9SSq/9GJWylL8Kk
Jmiw/L4Pe+nwzJQC7fZ0zjjq2smqWBNiX9G6qYASTC/cSqKpNWxY2d1CpF28Z0zlRCOWkgxWNk0e
Vl2/n3T4SUfoRImTsKuNdwc8gj7C+RPB2aNU7sPuveu0bSfLBsDeamdMqXbYRfGS/NCEnnKxXeMm
PBRvRPpYome5YlyYuZ51XKmNdnIP3xMx413v/ujkmksFwrDOCAMy6S8p1cp/K36vx3yvmqWsKbxG
YPhA/HRkz9HzdvG0xEHdhNhlHUAT4U8NB5ofh+kuBXFt2bcf/KGmRDzTc1CHiHINjhzrLpGy9VRR
4qaxe8ldWtgx0orOQfv7qFqKmWwr8CdPpEP8VcZtBDXECRUQrAMGGYvN3pkZBuF9mmX97XNQBMd1
Ot9OWcPkkofdWAihzIxGGj8MPXPbeBg9mRZJFbbm/JoJyPjtvcEHWOhddAJgCHLQRJ9tVODR677t
fIowMaSgvD8mA0gVzbgoDaJcDC5iIwFA81KRVz6asBL0peVfY7QaKJWAFb9zaVJ2d6kQ+ggItJ2r
ouXASKGKAIWX7up5ub+8CJcuS7TiYHTXD69x7TjRhgKbdM/Q+PEGyz6Y1Si9M7wCCkHbmKk4dYxT
GNgByooKbR/5fN7+/h2+ZdX7khL6OCF0+R+xg2JvRLf7cJdKd9qUBjkayLsWPhFq/Mhm0kPbATfn
kW6avni4DRIZ5y5eVSODOLwWx2PJxG+NR7v53/mdrlK6UEPI2ikUY8/w4SPKTk1nZ7wZ21MHVxWj
kOaQcQuVaZ0mo7Iua5nHWla7hKrZZMPT5GLQA7VZyzSuYUop5sB10FWcDS4nowLAOqda7OPhLPOu
vn5SyoN44W+baY/fdMN6xjDIhgXkV1tzNcJ7yIu14kQeu09UBU7HPW2Gm50Kgt9WYEbFCwq7U7j9
e2HvLZjSj3Y3pf3qxraCdJPHfHIlZ9wz9TyVjUz/UAV/lvEB5R7M+AzVxOQaW64Z4ZuLF91W4yQ+
PQxvbhyHFjwG9YyyakCYDnsrW5heY0B+hgYreoiJXCojqvwziQ6PahQOnsGtfmp4Yfbmnqo477gR
dL/4ixlxbh3PqxoAK4UqiyRKGqaROoG2jQS+see6yewcT0Xn7kr8RFbCYkHrlvw3vpzDkuBHlRgE
l3EvH1C0gsdqG883JOsgAPniL+B7eGXf0azX3RO2yQ+SZg18tr4mff2rFnUYnmRyom0Tc6fGztEV
UM/BAbmNmMUu9VeU+XB9GqgRqKzZ5KSiBBoVa/EFgNA9qpAbt9s3frI0CUydcMmKzzk+uaLPLMdh
6WCjhMCo61CE3zgNHVNHF7VMqFctOwbBsblOoswNqZx3k/hGMmy3WkcAwonh7z+WcYF8QuGX5vW2
bBD/IFcAEWpLDdnSjjXizlUVUOJ1AfvByFNWXY1SO3VOlP31CiO9X/b2EuGlO6OjdDGd6ZAUQuqC
Ub8MIAZdIe1XpGIL5JDy3ZIeq/z1C+prWxQbjvnkyfbhiG0oCaXicC4s/eYB8EhqXPn8OMJQJo7S
LeHleNsyPQLTI5vR+7EEpdhMrSmw0JKftlvsa1+fW1/iNF6rc1bttKLJUaDx/S1BVqKmWTur5y8T
MsiSx3JbqqHlVWqAYtNpvgK6+Wni9IOgHqRCJu1n/wmS8CsNPUPgb1SrZOu/pAc8z7zm0ToNU8Zd
hrD2H9E4XiYMuEiQof+Ie52qXwDyKXCkTfpF3V8TTMmV/IAAsmosmHcKAjaELIz8tLFxvmcEImr5
HI05osh6bX/wlMFAGvx0II/3EkCw4NqSDuS21s+Je992cs/jv8KHYaz5tfZ2GSBhoMyuoxFjV0n3
AKK48t5QFRhZSTeU2ci6jn7w2XkwOUI/TY17tx3JV3QGP/0T80vf8m8stVmgd5AGE5LCYeaum8F2
nyASdXgqCJwXpimFu+0+Uzs5FYT0myLBOUObTW6gd7T0mScNfRsx+fas03cxJ0fXVTB7IzsSCyP9
ZrFHcCOCV7F8p6EzsmY0Kd7iBLQ/Cve7sd2gBjUNvi4eniYkPfdV46eSTLs/oq5L+8RETiHWge0k
nojja1XGUOdFl1aRiUYCeriIUlUxRWvvGLuI7ScgtaaPe4My8HNSJr3wMjB35lJftiVHfwDMnUq9
7DUk7X+/qymB+JTHmjbK+/VJzDxGrxnRqJuqDcQasBeEJMPI99SjgZg7YuJb2GQkXQtf0ujdHG1n
f+nIoBQtRPJig4iYjQ08nU6XQsTIlH+3B8qkGJdbPNhcAAFWSIrrg08cFFCL9cjJoyEy2kQn0tIi
cFuzL/7jupIj1Z2oW0wxF0Hj2TBN91H8mx6JNLtIuDKEwmEAxe2AUrEQbC3fK+sw5WbyfIYRrKaF
TL33UEcs03IWUNHwsTOxQcx95pA5NEy9Zj7ODx3+hqim2FCnUrWoWJl+adqyDGRQ5EIlS64OUf4+
fRJvsyugAzc5EjvHP/yhzBNTjqzrVVX15fgOj47O16TnLUiXwYojinbPjlp69KDcxxonq++ip44k
IEc2xtCSpat+r2+nig42cIYYs/lMjNeT4vsB2wBeDL2tDXwINf04KeH2QLN8Yl5rl94JsVM9Eamv
eCUcz8Q3PKCqYW+F6J2tWnSWYIkwiPKz0mPBGXVMhgRhexRd8niu2NYig6r4XVv8HvbNC+5NtSnu
DfkTDpqRNVS5T3DCr3lzMJon9NPBNeuV/wcN0gydM/p0GIol6A6r/7Df/F1WEkelLE+ShMNVJlkX
NICnUD3n/+/OdlMuugVujS6/+F5vdvJPq7Ms6abmZIdzBD5TLNN9JEkykZnpoFAT2VhIkJZlw/nF
HD+Z9Y/BLLDPlIMYs2ruBVF9F3EwXcu9Ps3eDJnO7XOcmOXsDWXFXhgxNM3+jigrswwwgi452CWb
B/v9WdvDZMmlBlUnL8GK6z7Lv0Ja1p/YFtgm0UFS5Ft54F73OwnaGCN9aqTqAUv2AXh5N7byQqnK
+s4wyLK5CIM24WvRFced6sSJmPL+5sKFG5vvy32bTeSZ61y0mkRVF30sfNGphf4biRoS3iAqTkbP
c1KjFr7CW4SDGbCFcBUvTH8ZtnUanxX+jiKWY1W1RRcSR7vwsc0dwVzCV6K4wFSrk6yPpTGFfYZZ
zhwcnClpwOOThGrKYl7sFhDvC+EpxB/eMR48/FaZOe3vpQN7ktmiNj+ePUfc3fZyFp+xg4BoEMSZ
L6QaNQYHoh4Omd08Q3YUm/5JC6dNLPb6PTx0vuoTfso+O2pK/pUNqAlkFGRlk/zKk8jytKudbpF0
2Gbtt05TNvURdBvOvkacDsqYHYXBWdFUw/V0kvuVbonzmu2BWUm9vP7L8pSMgVB3EfOeYf5Lvs/A
bv0HK0BeykTZJoGKNI/KKnet6C9gVavumQ40cQmiM1zXtFUZC5hXBoXj3KeGBQJyfrVF7eXfhNmp
qF98OExl9lBrlZhwMOP456mSBQf2Nv7Du3+O7B3wpEGWk08aI5x0JHqsYehmVfYHUgZZB9FFJeB/
5VgPZYL5QW38nEacCzMnelaBsWEX7B715BeFj979pRHZPVFyX6O3rEoKu0s9Jx66yIjmeRSOL/IB
gZzEtiT33xTc48shOZ94q2Tkbh1xBYs5xKyiy0gY+0woOuVnUO2BaNzZXVbBbUY5iRPbukuRaucS
TIj/fqcHVIl0NtuReeAyDVq7p063ympNdWzmuDnlimmqvuLxJ2n6oO6hTDBoaUYF/PMaba5tytQp
Ad9QkAMa1M2X96RlSSDAJQv3s8nrRwVE3zjUqUXrkvfgVBhrCB+tGmvzElcF9vsGaq2jGUnllSRq
dy5lOQp5kSoS54CxTy3xuTgntVoXqZ7qZ2TTB9GBaaBJFgNwyJQpEyx72KaXexRCwO0NcjV485mk
DsIMRCAYcZYueXkNkX0S4Wiv+RD71EDAsqaRvWf04xlivxUIpC/WP+92r1bu90cmqldWnyWE5sFA
amJDvcfU9YhluxrEBXDu42MhLxAisEiilmCiEhi2A1CBUVwP8M+gHvILFfpV0JymBSbMDIVhC2cN
aar/PiLh1oqE0jkaXHTkRtAZ8mpHvQ8+t52mnJMoGG31nMX9rYBo9VNWZvwDelUx8iE72S39RLEM
jKQdJncENbwmWjbIor56S0NpX4+rYDSspgZdo+irTYbmNsLmAn1lqPfaiNw0rXvyGG0fS5GaUkqp
s2s2dv8w1rBZL43ZcivTCtoyppNsIfTqGO7C6u6PuleM0RFsA/EUnNZUA0z8bta8YJF7KTjrDYwx
xH85xboQwa+w7kj4lK1P7j1XztJxoHmWsZACIwpexU6gvtE3w1PcorGDbJ35kFEwnTbLmblrE+W6
H1DpHXAjD6E+5h83QWSc5Fb+DMoA2Yt4wD4fAkC/fyiEuKMTKIJ/n2e3Nm2QFBYOtt2Sd0t6CK9t
FCvFY/3I0+Xe0rGUcM9iZPtKBYk3BLGC6C0d+4yg9oyBChOM3V6aXj905gU70pd3lgmqbjClqUe0
Qfaj0NclXrpMWP0FmNIsAJCIVPvYWM2DvoOVsOtrDh6Ez2tons9qSouiep/u6gJ1Nm50xQj+XMMw
Ek2jxtapQjyxkQv0Rf9O3kLczMN3Pdl1OnNpXXmPLJUYv/dPz/72dOG7zUhX7lm+djeaCOB7/nsN
f9q25Pug1K+EzdtydiPfrimssioyH2i4MEqy3WsQVSE+fAlxfmTge9etCw8LVOR7SqlOmSbhoKHn
OWU0/5S7DQgoIo8ImdjCUGtzA8eViA4CItuZtlMYaE+l7jSG9cpd7HCmBPmD+Ch77IqWJdt8zQDv
R+E5PkaQtchUdxoQbU+1RXllwrYOwWzu/gsMqx9WFR8dJFJv0ixD2dwc7ffFDG5obsX5oMzk3PCM
4ShfFOVyhQuE+1J1TuBv43qqREFydlRR375E0cSDUIMbIDZw6E2itPvYEEOBdNPnIuNPskgMt3yG
MQpttmhLpdNwMqGGAXb6VJyJS3lvXR149atOJjYt+KORtCxbrwwZVQjrHde916/EJI8bCkLMxOhq
/h/++wKtKquSiuS7utwrdQt/uwHeOpvcO3HOpSFdK/oy/QWkAtXjQ8FTexznMayY6zWaRk1wrCyf
4cy+/hLsZNWDKEDnvm3TquY6s6Wr9ZG9rZbpKD0tSf+JGkrskpM+jLS20pSI5o3jiDVIeiUWpve8
lK/Ul8Oorh9WuHvV87IxPkiC8qXtQiwOb9Vgoi0RkttVhv6jV9AETKgDM0Tkmw9pQlM6uQou1UBV
lzW8VZ71NdDa/KbhRmciXEiyYPXkcPU4rFJ2J+fx8kV+IdkRvmMlsI7V1ATVjKXd3mWN1K789DcF
AASrEn/3Fdy1zEI7qmvk/vzSl9BgSXZUgZ4NWs0oPS3ZRBS+70zpVSwEpDlfDoTu/ky0bwo/C08z
knsoOw+p9BwmraOJMuLt5W8Dcx7Ix2lFPQukfEXhUTJepFkfpaZBo9MY2plZ07JmtkJEDxojwjCd
iUhcrj0zkpGlw+bdcjZPYaG1R/w7nI6fCVAW43YTirVbNIlgcRVkbq9rxoLdFabCzzEASWer7+zM
NybaGjiqx0svNsZIbvf/vkHqRxZfJnTUnwCBk+uw/rUJ6i6hcx547LJw6P/M6Yh3F6NMEzR1InnU
lWP8KAg6AtZKhAqKhniAyfuXRf+BfBgXc3xjK+sftHUHTCiXp5v2zbEtVWXPdt6YggqK0qquOGCW
GxNc0U/sp3qUePXwOG4ePgmKum8bHEo5e4CUpeLjl9z1C1Q87YFLLum+C+oOKeyLsV2zFhAqk2Ta
LeyEtmPptILdcJbcV9ndr1m20pk+LKE3XL+qUtCoILd7DZQEJnHoA6mXBaR88lNPS71kcEHUe3iM
NMe6jFdw9CWJRRDkJJQ10l6f3AyfezdyAET801NrGn2T8x15hmSE/ewNxg7JroWNhm4/TEKrwOK+
AvETGVFEAX49hLjf04ibtmR1cU8XraP06dSyq4j1Y+BOfVr2YMSvrt7MqIzg1OojoT6sEq9qpbMd
tHsobclZusoI4USZ8DSKOFdVcSxXNrS5uGhoDXV0hBO9KdWXPcVkZrd6mXVSqyLvFQqmdjH2BJJb
pZU55u6fMydrhSy24AAtTZoe2BiYG+xG8iGbYJ9vlgkK8uCMac1VYEW2vtRxiUYol4YWC9SkHrpm
b8pH31FVdRYdURVRe6V3yi3nBGmHv9LWZRmVj9QzmBMeAENh4CEWxuvW4z7LPNbBJKlT7kRbF2sP
aikUU2lNRXOJ8cobyu/FMpAagQg4rWoIQvPRTc26I/KjKQAy6QqOObrIToC24dRe8yVZqwxA44yu
jkqDCsA8ygU5//+FVjPYd+NHsxuCM2BTp7ZUlamLUQc5jxRpYS9kVZnAlWcuHcWzUZ8l4hfBj8jM
f8aXs6gkK4j2OG7LnJshAtjCj9zV6eUKYbOd2ZVjthoxMP9UND7oakSIJRamhfsg1MqICdOsh4uX
V0Nvb6yCAH8/le0qhyGrvRgjyAdRBp3ti6FsPoU0unkLcdoU9ZAMLsSPKovPaJKIuTDKJHuBhDKC
OFwyvgDGz5NnUYGD0UdBjbGyU6FmX+v6aSMtXK1ZQXQIEELhsm8017TwBXkQ9cvoNthkBapbuSK5
byyvDfzDbczcJ9ap6ygFRAaRoARmQy5PNPL63EIZjRdrqtsOVh3IE7t+IKJfCyLipnuAYUOGb2rA
r8wl1utB4HKBCK1OkuUACV0xESSrXwAsNoeRypKhWeyAKT4+FOx4fTAh9Xw6YbbyD6zfrHQANUwS
tRED/0klJTwJdhUTrQcDFfq/ryQtobnDqrfMuYd8XquHHrT9CT1fNEsF+FbQ+JardNMGsrmeE7Ce
5fusFWooD3VLvZsNh9FTuz6JiBJpz1Q3KIBAOkNxuw6nJL5RgedKyrboba9pNsuZQjLHrzdhGVMp
IDQYgXAvzPwrLZs2eygc74ycrzhqfFTTp03VEepERm9o6WPMyByxYo0svr+IOql438SpkCnsadVn
32YmRPLt0KmYnaLhCzAWmzdsCviGVtqRyJASXTT7okfcFeDkTYKDTbilD6BActZWuofzb8Q7Ywtk
wraS6SXRNKs43YhyUEqoOF/lMW1Cbog3/KHZummgi/ilDaMh220JNZ8Yg/ejWzd50Q3klaCaobBd
+e5pi6vezVHpOQ1NwrUxbpF2nMz1kCdUeXmgjT1uB0+KXsf88V5m53ExJ9MY59JYRklQ6ZTm6A0o
wLDgPCNJEFMcWx0os4UhXAObd89WOIiLzyEJNgchPfXmB6cWnZEBlvlP82XwCijTYdRlNaFPJQ3H
6aresfyYG7gksfOJ9sE3fPxqVBCJeru16C3YYJ3CCT6tG0qMnZhNhKRqNpy6l4a+OugJMYVYxp3J
YKP2s1Waxbfx+QJFubc3Sgo6vZsMIJ6QEnhh13C8eJ4wnAFM3az3YQKNCY8MbFGhz1+D9f6e4Riw
ffflAkPp7kPxv8JAkqK0Nk4jVx6Kcieia3z1+rEAaOodl3eVoYnphwaMz9xiSTvq9ng0g/jmJBRd
gdJpyAk5/wsuEzevz8iyiPTR5KN4nIXo8aXYd6oSwxvLdo96pRilryx2Puw05yIby/7sgxlPPFG+
xaRGMUU1GOeJDOvc7EtMQFt9DPyBftf0f15prx9wCsSCq3XQywqFaeSlUZMk8QAlV4+dK+/jyzbe
jiY81gbGcVyrwlOJaPcKbAfH1brhMJKmQLEwt8wjvfGgiFd1JwL8FlrNEB/kM12moR5QnN5B4s+b
+vAdRrAw+WvsJaCRk+yN3n59zDw328VE5mVDzIYtttGRnkLkaDVRJA/IFmeSJte2MoWhT13wYgvX
g0U9G9VpCuYxdaxLqrPHFwZnm1WXfgt9p2FFP0EEWagItoFgxjFS8xl/npMblqkTsAwJCD+y4bty
enLRY4lD1DJlfTDDxj0KFTmtIhgcyCVaqCFMebqr0zL6y6ZxyuDRMKn1DhNcowi3l+WvfoeTvdHA
tYVaAz6LjVi3i5EnHV08kObBY71Ftbk+vQY3xWmA9EMHqM9miY/X/0wtP6NOufUqbLFuQZcLLfMm
5QVEoUI8wDlXzafpjwDcrpgVpuaB/2RTJP3NTTTa2LKrWDfR3Tk9NVpok5G0zbZfGN06nknO33nk
BGsQq1CuFsBPaqDwf04qUiJJkjrsK5nxEA/bOqD7Yaf+GyYpBLZkibFj1UoBpEAgYER2GgD95ICy
yqe3cQ5y8fElnehfSpOLiJvQuf8EDQpZmjKjSFGlPWIDRlM3cypmc1DMprys6BwkoN2uOCP/l/J4
DD2Gh+XOL4H9Xsp2VkRSVMrq6mNNNB282etvMAdUpv3XcT/Lu/PlaMMa7D5NT++zadbd5Uuif+aV
lnJ7GFAQ+g71hUwvjsl+Z+AxEJy2fIC3ZPcyHfh0iLeaNz1F07krX4PORAqs8UcLfNCDeh+3aib6
7KShpFdv3ib34wg7AAF0G6ze+DXsONfCe9KmzwgJvv+QE4otCym0SGNfeSUcVbAJveARdGzorheF
rFvVdQRl0ksZDzlGsFjOWgHiZe/ER1+dBSQWc7EvXAb2k4b7+ZHvJjEleSJtJaIHoceXJTnVLlof
YZe+U9nA2lQXAMbUMtSVenDEIi/n8mNEGEPz65evX76DemroRrSN74OX6qm5hfldK4sfYEWakQYg
wCWp6PlTMDhA5hvU0rI7+3tSuBPCq1NxVjwgyh12dP3G7Lkadx6l+lm0wu2cM5S/nVCsTpocqGeq
Kw8hJnEDy9ahp4IQCysg/exopqGbwyDXeoWct5NgChwJgKe9UE6wXQ3JQOpZlhVu+jzg2jjQHU9Y
HZezrnYjEtNsIDMyt0Yv20DlnlAdpPPVtmCQN2D7/wtOC2bg2L9QOnhMXLcOScw5bMKIqtn90p96
vbsJuZpT1Q5w2uyXqNSnwlPraMCWfyw5112X3PxA82gjrjobDg3lsiW7rqsl9i+FI+iZ9HT77dt0
ICfC2G7rGUf/U1f27uRE3NKCMDUQVB09zXoiPQA1YOsD1ijyff4DsbT+F9+ekwzZvznBeHiPEniP
Vt+mYoV9MiBygqzmRFpLbjEeMjbgwO0OI+ko5qaQtZQGO0rY3QgNVhYrS9Tq+HeUKQ6F/F9H0dIt
qgwWIoMb8zuiUdIHrYsuMDow3hANLuqunVTLfYb7h/CuVuxNe5EFCcY+TXgksdsPu+3wA+ljHcv/
1qRWoiYKE0ezTO+tOFRZ1wLG79v0YSU9m0IDTYFFrLl+7INsJOc9JpaCx8sKypVIJp5IMZPpKiDA
bLQB0FCB84QkD7v94kuOEVrzUGCOzgDt1It233WzHN8R5HXPm/Jl3qK60o0EvOIj6iKi5+Uzmpt9
HdyrNKKZgAOGKuQmatBQxu2cZtfhO0vK8WPEUZGjlytlZtocWSjKpIqxJ6QmvJQ6/fcriwVKlExW
AKWp+83pVCvE+0AxLHHCfWoYc53OVpL/DXTHrwBHG/RH/+RFlx6MFzwsqLhIhwoLpPJFAUtRUgCA
yJ6EoCyTTCVwZFnFAUV/P+3diX7IwzoKOryuWGV891JTeE5Wqod+usSyu3ToORT5PKQDQz5FlyDy
mn7z8BYpf0xHpq9IvBypdvruElke3T4eK/ND/v8nMtav7YawReDYmM5Bg9qq/XJUcPVAq2lvxjZN
M5f1cWzdcGOke/BsMcRK7+LRcLsJ2y/qDWZAdk1U+QmaK/8JRiPzEVLLi5Z929l7dMy8xD5XfyzB
XdxDQIqmQwveuuNQH5XucDCAik5njBR4CpzqJdgk5v0b4F0GsL7axBrG5iJu9w0sa9manRu0Rfdy
4hKibDnowokJzcDFcd5btpe6ASTFGIrVRBqSoJ5EQd9Dx4NxY4SFdP68xL6lwOjjwxkuRieiRy31
l9IcywsUoL8TOgQx2KUPGk4XphgHehJ7Bn7kUQO3MMHGWXYFeUwzy8VVHHGgnJ6AefW/KGfYq+lV
Js/kLEeJuMhArXkyuszZ4y/n0b1MJbRHiEKERPt3MzjO7bDl1RhA7JKq+LLdxI9FumiZtdZhQsPE
0KHIZRkPBRujY5Tg1ot+Zwjw7yuF89rNlhUN7AeGLPxVU8MZVGzOuhy4zchob/PtanZM4GTnlTDv
vI6pa/1aT9RvkwFbHjo8VufgM5fXWhCxgP6ivlsjrfpGVgspwiFD75d4x4Y6M2V0NRKGqvRlVmhC
cO5Wu4VQzv4N9b3PJfXN8oePMKD/HWwx2pULUPRftIkcHShiWoW5wsvdTjuPJapGB3Pqn44rGlJR
mjetXhA0jpAnCmJkSRgNQiBZ2xZZgzbFUXZYJ0KoFbe6LiVysC6QUn5q4xun6kduOH0Qz5KePUVt
P39HacwGQ5kGQ9nySX/SDbgs9OmPNhVUvaJsnqwjfiIHk1NOit16tvEoF69XM2VXjS2RM+wgQ5qO
bvHZtlaCYnNzvQ4+sH4SSHA3tiqeqXq04n/H0PZR8pr5g8q0H3AKWKnjGOygaF9ELm2I2sqjeic3
ATBb3M9A1CkN4d+np57bXub0iHw25TKOue6YQlJxfUgY7LDkDeBZU/FYRZDZ/8d/+45+Mcm+eisX
Q33CIeIKGB4k7tJM2MQxvPuuacnUr/UKxkhWkqqsyiedRQ5Mn4n/+cfqLpQLpCj+RufrarTjXYmP
7Zs/aoeaJWmmu6Rt0z/DNYD85JU065nh/D0oeKkUvaQHIzaWvaxegHGNzowouNlFAU/hL+Cn0oeN
OWgxDl0GrUHqPP0S7XD9P8T/Ej7TGykDuoeSIj8oXdIRoWDP4NuuantNdCLX7Hb7aDN6e7Pn8yox
iIIIdRPWD8iAdohKW9bo1cWyRk1VYXBq4QKx5ZLRmTmdf5Zp6zJWmKui/XOrZ5TOen3tKF+4J1n8
Yjw7xATjZ/WjRBzOa0kARDTX6PwQqAeIwdxCTNSEm5lhiWaalAndTF9uNTsSU58bzDD0r7b0C7Gb
nxaVwiQobXfctdyt+bCg7yZ9z5aSp8kEcEYjypVKJQeUOvV5bzXnk57ObWpkjM6KsbmsE/2Y17Gr
Mw2ibpmEWBMy+M/EGTTk0i1s8s2QV9RT2hpjXpA18u/0Q6q40gm+6UE/FO0MsCdtlhCRcZFermuH
Zvv8cBk/axPIKIpAZtXkIpOl/IVTprDJ9WWM9uCEbnmQ8dUvR40KYS6bwARKw/qpDjX9seSikU5G
iT5w8wHHUF4Biaj1jz5xKD/kpkJl+uUBDvOdHIZz4AwEMKTIYEBjakkZjwoWBUoUoAHc+8joJksG
/GXdbIzeiYClADCO63DkOJnCc5z453lCielgDg5jUbtADRzoY35GMNn3H+Z098Ct3Wf/L3PDYNO3
vIP4n40/cefVf/7IXrY5waRZ+pFW9OakiC2WibH3PYs7XRkuFPMhL4k3IZ+K8Q8r7yTYXuHmNxho
z1KGy5qaazfQYruj3r8smc4MU9fSuz+XEVXIt6z41fh/FiWkTabpgPczQkVen0IeXTiySfS61EkR
QlV6XNzocHf9BSq9otcnH2I/xzi6rWAELMLsMCCh7ZH4lov6AxaGIHuGGDtUnO4mvlp3X5JPul8C
lJjoArZOMGq5OVeBz5uFM6FZ+qouvMzPZ8fjBha8bZX/IHyDOeQ6Z5fyK6M+YonCBywsiYzL5s4I
aoppy6VmTJYTl9zIlGy/PSKUsOVw6UzjinX484YqDAfwwf4EbNqsKKALCpMAsgVn8wMI1Lh2EW6j
7rguLeH/3WpZRrv0jjO8OztSrhc8DZi0yN+X+9VxjC/W/ap7hqTDZz+B+nwSzfN3FFsRwsoPeYCX
XgGdjC8ydMLgF66MfO+4GC4mkn88WVV2E2W4pOEk9r+r/KtzlEfVBkvW4OyHhxnZL8swkLct06sl
3dBhWo1Bxpnhtm6iaVmq7urUDtfNTC2A2cZTwZRK8kwUTyMTEYz5zrbxSh4AhNyv56PkZstNVeWi
tzmAOMpQG8CyWUK4O+x3K8Vsvgg25HaC+QXlOX17VA+ux3ud3K7heslYjBkRSKMoFf5kGNKYalWV
ftayakhbMbTpfpKytfSmR2lZpp9E+ASbLeAZcxWfnpmawuwEPgXLD8mTdCHJFnt23uhdILXxvvDs
wD3xwUxHOa9ocE1Dz0DzrwqhNuVWrslIhlIKOea1xH1RBGnQ1Ius0lZp17EbYo3+EdB6BcNefEBR
MA+4fKJdm1G9/6sarBGflbzaoSH35m+gCSKSVc+3W/uLvDdv4ZYXZ5gkRE+kYCe4baxg4wLZoEBq
P/+VOIOxkz6A9PmF9qQ0Y0Dt+fbcaUur+oYQ5bLUl90Dq/QDLwiicUVg8IYevgzrNHU/KlMsY8jk
e4e5GLck+Zm8MJr3cmwJbgvGOlJyneO2R3Yq4ZysLo85wpUBTlVlJKXn23L+e94ebpjDWp/Kp8SR
4G1dUU4W/42WWAQ5uHpDIL2+3Hc8ogqRD8SqLYZeyLDH6WFGJgpOcdDrkvf8qoWDMRb+zXD27ev4
+zZAtDanhx3wQxHNJqIq//ZiOj6lkOpYE7Ru9eD6PaRZPCq9ZgkFdiiKAywhm4PBcxWsIG0DBdvc
5dvh5ZiTeehbP8468N+f1Y/w8n1/Re9SR/wFOQ3oZfpBbez+d448W+wnI7i8oEgKhGvfMN9RDx5O
PBKYzUXz5xLNCeh3yDzbXZuuAzlXp0WmhHMewKOS+i3meNIw4g+Ck4w+ddT3M3aeDBBeyvCQv8q5
/ng9hIoYNQ+CUn/AeJIBjpDCZg9ew9ldMkcrJ27SiOKJM8mevyd14Sqi8y5FDXJ6gztRHntEgZHS
/r3WRTKEcbMsAtfQTp+jqa6U/9lAjHXzQQgpD1KLa1DomWEeguCt8T6HL+sR6nrwUSW2tJhZpWI8
ctBCuoP1yzyOj8SdZf+foBc+NLkm2/rGk1FKcRceKNXKDwRnqMQTagpMHR6C2C5RgbUcjGWnj3nB
SrIxDp4KZkGaEyM3/qxstEEd5cuwVtrYELm6cZptGvqkko7030ogBXV2aCBrapiBQoK9SqkzDDHL
BvDzD+qrtxlChCasugJU+2gS3hckst13+hqgPEI+RlFbMzam0bOxIXGHSwoHvuLFYK/cWGfrtbgT
gQeesHSEbb/Uf9PO8A5KCdNspFUuLof4QS1puvBNSuNb/LHMrze+xQRai6y/jAHDK36lsPVM1kJ7
3lnGfAHRN974jLFdiO4hRQtMicZvtKbIBOY76OdtpwgevosydHD46PpzBsTM7dX4n4xOg/xwDSLm
w+yLb2MY4LNnmENtszhXJxoM4LZX2h1t4Ga3rJnWkViRCrfGFGuVYMreNCCif+EKl1NsI/bb/YXO
NpFVIen384/qaVJN6wl0Z70zqx1uBnIgtgh5IOjrL2c0lQThBxQoJ+cKxxTr+Ft76iwApOFagQBv
+pchQVIKEHjzsv5LLabFrLPtpakok1fqgVAJwHmPcvOv5TENbg5i1GBsAgYQxjieTueHXjOz2gvX
o48Cc1g+jHjFtW2IpyWLnR/47vb1shax5IxQ5OnFukAIPfZcFbBQfGduSAB55nKI1qwk7KVBqtSP
vSrmWGJzwUu3k/IhHVwGHeESJzfLt0xvxbeecGGv1jVWluNiZ0dk55J5ZWqS8I7H6yk8w+4bhRyf
dQbEHh0B7HBoO0T7fxC+5k9f7lIJOus0AN2iUldcpzNSIcopT/48/5yu11lwbj6Qmzhwlwkhx/cX
/c2SkYUv82e2iJezXq+dSw0WunPpHv4d7TczYbs+CbbglkbfUALblssawhzcZvqgVhUYl+1hbHoI
9JP9QoHcJALaYLsIKLH1V6unbZ4jj3vfP3Vu8Xwiuu2q6fywBqt7Mm5x7GOHXjMXl651Ch4t4cMm
xVBE6m8lQrwFY+iMcZ+HnmAoXNlIsl1Fd76g2xR8/QsTpBZ5jH5N+ZXmh9aHXWob5kp9GX75tNhG
ZACljt2rTgcb1ULA3eKs+6OExdqZz29wZp70p3KYuB00raVuYhVCFBx3lL4WPk2lN/ln1TorMVhX
elyN9v9y/vHcP8VvlQyDnBGHyy4fmATbIVemMiNKGVTEwtpLYPn07CIuzxYt4Qj2qLdfTYf/r/KG
E5cUbiQfKQdvJ3FYhMTTL9F/spbjzKNKA7tYUMBory6YEcWcYSNllQVpZFHizCl6QtDx3SVuyjK/
SbnbqqDGia8w2+TeimeeoGU279mOeT0WSPGBdFQwe1lpO7ZW6x4OkQSkWhYcD49aEV3470Jhp16h
bNcwc5939tNYT+5IIFDEjDeqMyHGj/0+O4YFp3RjyFmE6wNOLs0KUJxLigjmhulLnZp0B3gGjO3Z
/KNjQ2YFLR4/uHG9e/ZH/i011DLWnDLzgv8zbig1ZdG9S5zIIhUvqcR2XgO6yHDHc7j5PSfMkFJo
yCRLhmZcH0m27w45DUnwfZrybhmJDpit3Fg6HDEcwY40LmToUJ6+6sguXW+33Rood95+zvMrbKvv
wcn58emIqpux/kz82J0gGSVclk1ST8o4OvNbg/urFgVRreHIM7JvOHpd9rwzQJ0jGeL03zdjMPWY
l0EIzLftM1AD8Jxr/xWfI5qIP9/OzKwa5xUpQXZf18ud1qAeSwNe2V2ELCWeTqtIIAxeQ/H9CC/K
l5gMISGCi4IMIy81udSw0Ug9o1ndmuhG+NeJSTb5ShIIEWo/Q+R8WHFyirA++KFBzCbqAdtEfVjB
PSuXDB8wQ05C7649wRzosOsw+ORwH8ayFfdWsnqb7keUHU9P5m9BQ22KWqbEKn1Vgl0sZOzICLzw
9ZQVBXWe6OEnQi/yOKwMnkiRKlyB6YzyCaBOttnoY/W4gcQRt9UB0MM19qLJobaT2wCu1N77PQIh
j1T2xVAYSjKOjBoO+nn7Z1Cm3YwU2kfmS3ci96psKY4Tres1SSgj4WBWupVr7prPJfNr5snnmFSx
TavwysXBkgQnllQ4qAQ59VTI0eaX3X8CWwOj+gkWkin4Med0Y5K0P/2/ytHl40KbbMOe8nFNM3Y5
wpaR4WZw+vGoq0GSil1C8fo5Of9ffXrI4HTu64lKiAThIPhD6h66W9szkU2FIKMna7r968iab5cK
xG+LMdUQ8tODcfo60AzH6f4Qaon+MHu5/Y6BZIZ3oZdXUSDcJmuXUFDlba9Yy/Mm+Yh8r51QuFqp
vOSTNETTaSUlVjHrcMl6o43LFj/JtckN2SgOf6eTtVAubKA1UFqptJsw9JfDylglAGndLqXGMFoI
t0UbKPwzVPApH9hzLTH21+XSNEbOYXkBOeenyMMs/7D+MihoUQIuCQcsW3cbO6dBPMccZ6tz2UMf
GaKr05llfONDL/CuGB1jyEr1lmbnkxYhPzGWtu9yuNQO8dmESAewXQWjFMCULN4ftR+MhkkVaqKV
1cUeYltYKrnrYN8nUBA9NzCMNJeKOfPG/w6AOeUWNhV3mmxKKAzQoTj+MHLARRMPdU2EXsqBtDbu
xzv7D8/BgE7CHWX252PYhBYbp6OA029ZHfASVnSf6jKPE589B0sdQbEbVaaY/gASIh4MHy8fMXN0
4UELWttAD86wKddnd+m598vb6V3GHn2SUACFfO45Ef9LYOKWx9/wDR6i+8t0geoIKj5TRdBgP9/+
AL+BLyAMN22i/a8NkaFFc7S4MPybpnmOzWP8J3R5FSPx+16rP2SzYIc0tUPTj/TbbY2eowrM0Nlv
8Y2It2rrf/JoFNUT51dhBX4gNVCVGZgTM6F8xd34tP2sTwQ7IEyO5pUcHjyDzW21sBHbk6/nRiYu
k86ZyR9LX2bWOGL3wkRwkpvhc9UmBBPj04ZeEE/svqcWwCGmY+88GCI4ighHJouOJGuk9wFNdQt1
Q5OXnF2WgbTj8vcJJahKc/ClgpMpDKqQe8l+SH8WsmCv/HlzZ2MekdE3G4FU/lZaYOxjTNbk79Jc
x1FNwTN34w2nO5Xn5zZ2AXJPIM+JBUnZ0rva3WaKw9ynh72aH/Wxl4RhxoH9F58+dLcL/9hihnPo
MbI8nB9YbeacWmaCCFSpFuxAFSy06gb019dn7oiMrzf0P+mcelXkKqtUfIR3Rg/JTsyTYITSpUvA
r+P4TglpuoFia0weS3znkXmiKAYPyleCVeX99pJfAWUljcHJQOK1upwwdg3HEChnz4oluYPCzPef
me160kvSNem10fr38E2YTf6REUAjUsiALB1Yax7rtxoracGYvQGP50wdxzr2atU7/ASjiwLxSA2D
d8P3uG1LxPBrIA3+JW3AFhi0w7EeZoNjtQKNVveyKg1Dr4QlXSw7vaFFLKYMOO2HKJu7rhNsSzAS
vNBZzW1UDyuYTeEigYgDg/LanyYd0bzMOBXVrBbjr6oRJ+cxrBKfYVRqhgxhOi84rD22/s/Js3Zl
6ENUYBrgQxfAXeT78gTdUI0vWerddj/QV8p5rhmg6DQgQwHaKpKvxjXLO4EKzmDmg1u7kJziEBy+
UZQiV2dmgtgQOuOpPqkM6q9fhbM8egptsAAf01BD/AtMea1/saj2Bg9heIVsiyoy25oOwFz8RqKI
3EjH0roJ6qDtz/u4VErfXJvZtA9+Es0k34Sa7Gp/PIt9PdIwuG1UbOsRkfcgfYngGdWiVNNRh3z6
JYTgAyGyEJ1kADoF8TX0CSB7xtCCIHMz1RiaNRvY0xhSyIXDAn7EPg7fYbjmT8DfNSEEOqAvpe5O
fTQo4L8ta2wHAvULWdVExc7zMZi4BkeV5X7CJpw0JcXjlpLRr80MTqz576hcG5TvcRFzMYT4+F+f
cZ44LooMQCTDzW5RhMGVbidjGutGEr5vuJrQFrlwPKDMvCWVIHNRB9xjD9nfhRSAOnWF2yKOVe7t
FN7BL1lMOCtCKUi3I50JtMHQzbGu8HvUY4dppUQ9qv1qv4oRN3Jw2olHlM/oLG269UnfrgZ16K2o
wqLGyYhFPPPJB9HJdH8hGS7qZEmH6aw5Hd3ytLRD41g/RgVAGe2IG96LLK9Kjg02raRBBPXovQ3A
cwyAgkwLP/rtvYh3oEbT/jFcqlV8PkjrL3tQGGkwrRG0LkXRkJkcVv9eBtYgblxkxptOGzkj1xLV
uAvwplEVFlao+VrKy4WZlKwvt5PbInjdXIch6AoY1LiwEu/mnc6DLNxaIzzVLhMbKIc58u36UNl6
sA8AAL52Ry/FtCbez6Hdvii08dlRIc3YpNphQkG+YUZYVV5GBCUO10P2A/80/yHmxQFmrvpV90PT
H2FBKmhwNTANxneXfAbOgEO+n0jDDesg21sATU2S9O+i+dclgaWZgmfLapvQv3lpNFZdWKiuh6YU
/qcm4XhPGFWdBjNhnLahUQZfuHeS7mn1AqwbwRjj5KjdWng2AK4ccdnmmXIqHUizJQL9/kGoFGKV
VZI4DwPCOw5j5tSrQmgvgzGrIlqelRuhWz7v9P3ReCMBJHiNd++dHjAlujijNqCIvot9Je1yzeHz
LSLsKriQt3ADFTsUSXQjPxzqbuWxj8GDgdZrN+4ZH0+bsSGSmyIW31eO69OYQ1Ka7euzyEuybBxE
AuPYMKeBzDy/5ysG+LjcN39KADSWF7ePWvmyVAgjxp1/ar/BRxg0bZChkCbKZsjGZrNr+23Zv9ni
dVT5srDd5QkBEoSS/6rm2expT0dTkMuYDEqFzA+lqKJyHYaxwDktSqtpLLLhDBmR0pGkCMBrZGXY
60dzO8As3y9JdBiaUSp0CvqHV3umnR1i8DY2TOw/sRrrjsOKuVnbQ+wkRaQvSmnvcYTU9TgRzOta
zC9Hrf4Z4NhUsNlVgAGTDhPkYnBKbuh/kXuB+7fBejAmjqm7IMlpR/YhN+mV2KMIrv7urLfZVNIR
bggzIxQSjA1z7yXhgNZDv+2nuFb6JUwQEgynar6IlY1mJKpz5yp588Odk/+nH4fcPpO4PSqSjACI
TEjgNB6MdcLpnlVTbOgtVMMxqUDq2bLOPZXnj2hjd3vqstx6PxCybuQOcsYD8jAm2q7hrC0ePge6
jMDBohLYpN/v51cvoRDVbHXKHMsllujolTaZlkKylqYfr3Npbl3lAdb1QK4aZIglrPHn4+UqZT5u
CPs4rtN7oj2lXLsKurnmmOAjIJQwaJPpdgiZ7k3hiR0InZdBGCZibPWXMLB9MQlXNwG8dZ7AoIAh
TRL/x0lDV7xESHLxiQC1S6et1LBtoQld23tS8QX+NCElKKxt9BGwIDzN9du3LdjXUIoegWthB5P8
KGQW/x/uumt3qqHHUduJYRhW4Ky6YJ7FHpULasZZDSCUpukJVGjNWfD3Sp2CpQ7IlcOkW81x0dsu
N2uYuEowYn3MikmRtOQzOvB766UQa7AKRGJ0n6IceiG4X0W1jFasBiaGpq1q5Wg3ytZrK8/xb7ab
35Fue4DS05Dzi9hkWdc0CCBmMFrOkcE8SX8t9Z72FKCd/ZtvjxSr6fehB5UnIcSBvvPEvujg1LR2
drmEXr7+YP8Zay5LhiPpxDfd6QHcHhuHhdTG84Z8n4XIHKFzcmOEUrL0M8n1qVId2vkyA6AHsREo
xCrDxxpS/HqZYl18Zg0aBfePvBTn3DadV5VHr9NVBoydtRXjk7xkVxISP3fTk30QbYsdxF5RnvVg
ljYgozTjoPaMfcxbtA5JOX+6flbqd/ggCTM518lU9UfJuXgDxejEnAqlBwl5AeUlhqcVVhxAtqTA
ooYLNvPryYijcx8tFzP1ZUUAxdLebR3iidWbzu8M6LCGTHD3cEk8URuOzTOZHvV68xdNsTHfhnym
Ee9uCV15AXjDBV1W/Gp+3Gi8qIFzR0/punDLKMpcsXp1AyFxWaH8Fcfzra9dR6gng9fEPjwmve41
bzodKw3bMlDezBVITWyIor6JT6Yt05evt6soAzIgyaTESnuoWviB4D+05nQOnUVgc8w/iVInrHpM
mj/hUnRp0W13GvTDByNsuJaUsLtskWGS271sUzm8LoyMSk9t4sLti0wFMlp62i3e6pI/uPk6wQWs
1fwxcYaRufDLy8FDURXFuMGK0r1r97MPaaqJv9MmClYTjUW8h5sAlgQ8w2ER/2sGOFZ1Ei7R4Ccy
ZVAS5BZqs2Ra3RiuGwJPZJ18gVJzouHupzNyV8MgbyRsH2uuBhK/i1Wxsiy2sf5g23DW/Dc6bGDD
KUpO2MEk/gWeLyUogZ7ilSLpdNJH/D4E57D+mG6l+pAxJwn91BFncnyO2iaR175uvVznRcgXQz0P
Be1GYH5DvlrRT2RVNUYOeXvq4TBwB+L8vxJu8QKuW68h2k97KROO7pqR3PvJMY0cAd69WPDT7F1v
DWK6ICB+LrlfWKg6tVmbvo6Uo53/Qon/f3x3yipIo75yziAChU80Ne5MAo0HS+VsEkWwKcwybs9A
LPat3lwII6kjy+9aPeyyfSGACgvCdB8RMt69SJtj68WFvxoNzSiZOb2xxDLpP5jQt/w3GQkOXk9C
MaU8z0Nld0SXxQWMQp7LQYg5UkOFYCA6xP4OcJwVe/hIJzkkL30QtLIkQRneiiSckA2SVARi/74T
esXQoF5Kz/cWTjtvRAjmSEfeZjRO9jXSttS4a9xv+VzaKgPC+QLWl9kuHlxNAa69ly15ISB7VX4a
ZR5vK2M9L+3Yv3b1vyoInpiVfd+mDFyeRaBsWu5cdBqXdByOxwB24yrn2ODWzrhtwyVcZbOomuqj
LvI7Q9XVtAx43FipCaZD92J5uLedll5e98VWwXirZzhF7dcDmuHydtX3O6OnYS7h09JiGIlsHv9x
CbcmfIocHB55rn7TbE3X0zyZRPaO0vgyYKGxJYtPzxtKzN4WFGyU4DVGcRoJ9TIiKLn0h3zC5sdl
v+3fECfoppcZBhsJKiqUWeLAXSr/Ca3pH8uC5OavoitmKa38ZtF3omg9Xc+F0DD7aVOZKvOmpUX6
WEi3nMb/NAbhQxzvAksvORiWwE2FKUmSDW5hHqD8lBShfAAjTXR2k2Dbd4EbItjANltXSXJsRYwl
/xN7WCZKkC8TFwsz7k0WDc0b7lhlN/IOdZypD4qBd+BWLG8C8BbV/JAT2Bnz5NwQcGImhBF7eA3m
tlU0C1VJ5KUabc/XXvLN3ND6PBolqS2yytKyWr1DBhpF6286qVQLs3do2K+kJB6BkJgyI0YGP3YU
UllO+TAr89AgxIIFq1upwZBYVqdYSxezgdYc3bvn1YV0sap2ofzYDOWj00ya4MPybp9mX8N4j3jE
4f7XmuQDjHJdUU6UhMN1EW7Z/1v/X+plnXJdzgGW5XJ708T0yfXONVKktxJSTjfE/etClk5t6d2c
oY+rbwO3mO2tiu9pbH1+jQPCwZFpz99823w3Aus1Q5Xe2c89yN1kI0EnfHbiSaaYbCf1/0BFR1/M
uNwvkWIQpBNlQCsgwzbz9bEFsqi8oOvylZi43dOXh06wxXWnlpZMn/5Qs3dE7pl8fOQFR1irfTGU
0yJ18TnicVLymz5hoJZ/QlNZhAZ+J0ltEKS6vmsyrtH/EW58CuDKGyMWKlBVzzcA8sy0vH7gS1s5
12u1t1rSMspYA/XjquFHewNCgj3qjeBVgMki584GPy6LNmstkunqDG7xpzIGiGeWDGN+W3yxlgUQ
KOlNtHKWxrGRi1uU4Lhj3rmbda1kGGdhqIQPSjbCPYMqpgxjtGXAjp2/HmuXOe2GPla069ia2va8
kx9o4m46QXkF5mrvyruJNpMlpVPWUqbg9ZmRhnvIYmSrEbVdVKV1VKgEAuV0gstn+oY5hulheLJl
17obv4O5DJ1El/olId07Vs2/DFZSZ2FDEcTsWNJ5z5DHS90oUOjH87Lsb3xzTuheYW/hIZh5Akiz
K6appeym1b5AUU6vVz1AGeJaM2q2E7EneCg5DbusdhsNM6kJ+7IBe6YaB/7pW1HtNEo7RLYYtoF7
rSm4Aoki2MigQK4+KfHUn9VocuU9Qb+SkUTWbP6XYNVlUP5HDiXsOK1Mb4JkreEVJSvH2N+Zq2mR
gQT+h9dpzuUAil8NJrPvaGPbzDxuZagwQWt8W4o3VVgU0NYxvi7Jma9TAlOxg356GtKRXGTCRGPi
itC+cUsw3wuJkCYqvlL/idXGs1HGKu1eQ+hHWKbsxCRHkwuUtLwcmXOmNxcvGcL8VXnq+trJuMWZ
8zQTEAn4iCLrAPnphZzSmGuEt+jpBiuyLa41ybtkJMFlqUovRVOjGM6739Tvw0qg+1oOw6qr2Ksb
16QXawfashv3S1JSi4yNfX9y5ZzauXmDkNATqyCHsWbn3fU+Xf5KB/sIeHkvw5HHwVw6ZCDe+UF0
xYu3W1/FTJ/Zo4QUW97iO7SVkCc0CVSl3vmo6o4RdEvaZmkIFS7iSgJ1FzZEosG6FylIVNB7zfmS
+1rfPaiE4zwLsqhu6KqJZldx5kl/5RMzg4sZrTeMxKK9WRz6tBklJpyRzKJz2jckMdrRNK8sWzMM
F280FAnhuZc1FsLXMb8fG9jIk2Th148wlclkjL4egaqgthz4TCy0v3owMVSIUZY+sowTonkBibEG
tyYtPkeDFg6NkltHID52lUMXcgPiVNb/cXMxCmrPlFbUH2Pd2ZiuCHuQXXq9+eQQkN1jSzbG1K3o
wz0e2Wbt39hjal3AmM9bS04yDYqyJvqDCRztrMpEFCt0511czeoe+57/JO78oaE38JwxHjICA/Dv
408CHallDpe1+wDIO1HU2jbncfPXivN7ZmVBQz10TNJdhmVUeAWm417GVq/ljPJZAzKW9BlGn46g
QaqANEEebAEpzPGcjW0QdvS4sro3QFRJBJowATH6w14HIxZho4iHt6b9qt/SXwTH+eaQ+ou15ac+
DgEjcLKyMhjL1KA7earnZDWed/pqiwyt/iIprjaahuQIGC+ZZBaRPVeld6f3tJ3dXgXLaRF7E5D0
TBw/dP0LbJ+lR7Ai/njaQD0gmllSdU7LDlzezdt8JXYa+KRC8tryauD/22bIT93vfa0uuJ0C1ld5
BZBtLuUwVXGgGn5sDmTG35yKmBw5e3/hT2/wK4t3St81AEtCCoGuM24XkM5jrww/sRWKxMMcUDn6
7d+aWG7Sw8HAkhGBqwJ+EJAFkAi/bsz22wkA2wpOM3wBeCzJa8vc2AReM7/OCYfb0MPc+aMi+CPb
Cu8HQyJw+O/UUOI+BF/p+hEG9t8m3HgUdcB7WuIpvR+niQ6/qrgp4vTQPVQc3vA8bxKE2AfSQCPz
cut4VQ6slSgWZZ7vlA3WRksIYsYoloACXumjxUu0w8iHNu8QHGl+b7xoBcJjh0nRFot4Qsclp92I
ffylBVOSn7S+gkf55waJcC6U88/ckh/rtf0ZI8rKqCnko7uJ1mFpCK2R8OeEqBTyA65gyOMtUzRY
792uwKNTd412z2ZunZyqVHkDLlM1ouOVcchAhMV3up5P6fjwuiOs8ikdBThgCQe5fxtT7uE/KcFs
RMiWNyWshpphyIHy7xgEZn31KanGJvrcZ0WCHm0bTffIVq1io16bEwealWkCcwBTIBQkjQeUSrqv
Yr+Ewb3V3B9lVOMG0hVwf2GJe1RoicCRDumJvN0eOjA/mMe6Uxq7SxuMyz8FgFXEDXYi8e0JapIV
mhjqXO46TVBEGLVcTUdIMcayI2YMvZnnGJW6S4gLwK5r2ozlD0Jsic3NE+nkcizk6wk/YXKgynYO
af1NEYx3DUXPK19gHLSIXXpfPtJbDOkgFgzQXFxpRAF8XrPeuu5Se3OOWS5hbP6qk6SKbV5fgJSm
VHK/C2abbVHkvREhrdn6EnoPzmYVu6Pt0uBru0FZ92pscoPa49dxhedYYwd41v4TjkrdPBgixL8j
TveuE4sVIBTwP82HNLzTevywwbgcbywCG8MxcPDIm3l1oUi/faIpiEvp4rkbea/PC7DfLfP5qlOc
o04aS2Qkz4SWLZWVjLeJR77viyTUPVHTJ0Xko+risf5lwbx8Tj4ddZFEKuFnDGHzRo8IS5LTzHzY
aHkoB1SFHoU2TmLNx2yHnAb6NwOynvWmJ/PpdnWF2SZnPpS8NICpxo4ntalwXgPDSyl87QLAh4qy
p5k+w7IjoNd8qG9L1atwyBSTYUYwsEC5/FJ9Jh2/qtZtppZM489MXv+fTAT/nkOn+wnSJyKDfVZ0
eA+p9SaEv7nDhSefg6mz7lknwCHZBERYHsZmJtXKp2hlgVN+RrGR0eVOlCHpOBC6kEq/TmFjXWoQ
U3C3ohdtJ06w25XlW8QJdzicbprAQ1doAAVdsSx3lfKhLh7jWKf+hd6GvYbBu/at9ZH4erdut4ul
cK8u1ERQwrAmg6Q4L1xBhBdEbkEWM3HidqjA/IsS0vgd/lXtTRqMOCI6kC3ut64PLNUHp52R6Ohw
nxcF7q6ThxnRSJhaFZtYQOoq7+Fmfg7KGGrkUeN8sHk00RtWNMIB+GbvqMwJ9JHELGiTokTGdHTM
7pBoXo0T2W2ZPEnEsuOdETgrEXIV97Ex6lawrABAztrOcAZHiEX/3MXqI5Txs1wMEwbk4XeiCtZj
Dv4PXwBX3PnsuF5biMWfRQIe9IRgIcex20spPlCcFhJcmDKJLKcul6InoU90U3UILow4Ha2w7RHL
e37XFHFbe+KmIBhafjegyEUncbFMsixIKDpwyt1fW9FwMl7x8f7ZocQhRHoIHLhKuVJXO3tmDrIZ
cEhCmHSugXFBdvASDw8zVL/5GfUBUTObTxKHuQr6F9caU5OTLJz4BQddihnMPQheKFuym/Ml9DVO
P7MGZjrEM2F0lQRYdRdEbRYwsLR6lyUwVXCgK8OOUrzbNT8SUM6rTq3lJ1FVQrxIcST8nNyMZWTZ
KugEHuwPNeyz+5mnDIMtVoivGhKwGxH9O6vjkGR6g8XRF2Kc++nga/9y8QiZgfGh+MZtdcihR3vI
APvq9uMvA09vTuqFZTgZQQhHjibg3RE5FGQ0GF4aUupyuDvU4hDEPZANttfY3LnQ2DiSJpwAYgGC
lzSn0+KYYpnXbUTGIKntlM91zK3ht3cmOG91/P1yy+ddIhe4HMYVVxzOzcQJNCh7+ghzm5EmID64
Y0vXouD+7boy0VCtgie9JFUapz20r7Z399X7OOUJWwe9sgu7/Qy8X2i3V7/D9t+wcWEohxiBm6ST
BLDkZazIIdVQsSvfZFP4TGnTCCLeD2mXFbHt+xNU6eMf33yQZfBPXFaBwVkW28JnaV27IT1ld9CB
PCFz/jhYWl6eZM350wqLMX2J/BDjyT6SfVWaIzLNX5zt+0SGRGjzuKssx1fi3/Dflh0COSfPArdc
bWVIBsZP93nr1GgPx1oyu/w++D8VZsxoPcZYabBsWkObSUbxiKDOguZ0ktOkRCHUB765mcWm9/M0
WsF4dGa/szBBFhv9EKWolitYqR0JQt6K6dEwse8v50GsogBSaU4arso9bfNvAPOsc+wAv0JcV85z
92TsxMCUntOe1VQ7QncmTlzN702/JWIp0bPbKPa8SB6z2MbdTFQZ3XEll1MQkZzAJ9Yvx76Pe4OG
k/Mw0hhNNU6v9pGZa7Oc6zYtL76/oA5e0WUtrez2AdN+26bHlUVqu/HQ2CruZ/uW8sYhIW7XJ9ME
L68Unv5/p4iVm83mnl4P21N79Mfnlg4Wh/5HiAjoyDF5TDy119OmtE6Lxu5hx9Y+qJ485AdyXKKT
oJ6nEeXWVJPLdmCC1XGAPB6zGwGEWCQSPM2EphmY3PrhQGGKUy//dsm+V+fp1ek5gzXt5/3um3wD
bKz3FPVU8giPc82YFzbBBba0BIiFOJJiMXc0Ei6z/a7ToyujcL3TwpoGf80LAsQysYqOtzEfYvT4
78y1a0HBYaKpacAbzXVa65F9p19RXRFlXkdq8I2/PxDQNgbfrYj3YNU6PDvA+1r5oOyzulzrmLDX
Lgb4Ykk0XHAr3PyANjox7YcIIssbO3kgQBircD8/TkgHRxoOl+NrXTIqqQAtnCir6j5RmwBl6UIi
03EUuVksyWcekmDVjnCQTLBt/v3uygV5I+AKnsO4OA8cUaVqqA+6+9OaMZFnmkCNztNHzeUtrrLa
3ODkj5DwWtma3hChfTgVfqKcPTV2uu1upNYL+vcl2sBtbbMpo6/v30T4zAu9PGef3oIb1oX79sK+
aCf/NjMdi3CwteuUURDIHKvYASeRMc0Hk70HAVI+PPtYD+eYtd6awzVAxaTSL4ctDl/ry2a1oywB
V5375Ns40eiU7v5I92SGGA+awg4L701OxHMJvNzh2HsxEyefdcV6uhn6KogtYW+I5b3Z06Dk08+9
EPtl/YBkO8A8uefKiiVqq9Jzixfj5+Xx21uCIZU95LcowXLvSVjqgAw68ddJ7ahFkD/P2i3Tcw4d
XFK2//0kd1n2ag44FOttHZA+DOrICQwpEPF5RpW9GLWIKsmVlYz7doSewiOQ3SLyyklsXIY/SHuZ
ZXVc06U2tiygeJtg4m02WJhsLnGzFvXfgW66en0Iwj37Knj7zvNBPeg039VF49Ezq2L4B+Gf5525
jIbKGO04T/8TU40YsWv2wFjfKyFNaAfE9c+D+F2plWuPSr0h4UxZWZmGO8MHTAbYYMBai71dfxEO
WzbwZ0Z+TE4mXiuT8ScYMDXOfl6RxR8FxVYut8x4ykt8RCEo0P5AGaUmwf7+f6fxM5Y/PrbrtP55
JINpCVe/f2eGDSwAVKpoBsxQMW2g7YLVwLJBCcoqYJCTTCHTWbHBwCJu5p31NLVhkj7Q7Y5LONDR
odlNAKjX6bST+q0gAkXjmZOernfSEOqLWVy1oobWpEjDg+X5Cs3UFBk3pk0bzjOoT8Y/5hjXWtvi
JmtqJD9zm9qDuQ8mMlAj1SWKJKprlaIvYgyQgvNGvdi8tGavO5dxRTOIjjgCRu8ZrIT/8epfNcTd
VpbHc+AxUZLIJobOBfOCjhJrUEyrwhtYcl3g65xceurV6u9X1uIOwBWsEljVzeQH+FAMm686+DMp
J2vmBGzJMLWUO/8zj523zdU9nEB+2CSOVYN4s92lt0YWCSFzzb7v4TIzQzJmOPYjtL/uZ8xy8h1N
v6vJFl8EP0iHLZ8OKYDflSIRNGQZ01+LR5cRL5tjBCqfNlpiDsD3TEHfm5UFbUJV1UtArd/h3IKi
rlUI/qDh3g4vkTza8S/GNipcS7Tch+fEwUeGL/VIud+uMla4NZZVxZvEHi2FeFBl/1wcTOJlt8sw
n4WWn8UKDnbxbl68gWZhSE3ResNJ1o/AdjcalU66P+4dld42xoXtbkCId3m3jOwO1bwqeYhNhXRf
/CcQNTB5qYUParid84hzPEq5HMENQ43oWAHe6cM9HpsAWiZgcks3iuTmhkJ2uNPxmkJq3tZeeieF
H8NB+Cyg4Lll3XPJUjluyIgaPVBrJTv18afi1cRQBJ7q8LYSRg21VY/Nh8dA9mNSktnLbXvAE2gA
fy7OUVO5+Iv4/H7FIc9L58zs3r3Dii6nBFzEW/x9ngU9VtoHI/xDuYKanxqIGMvBkVntPbAOAoiw
ImzBT1ui/DRLPzoBlYmmPiXakIXm/GaQ/WxsWHGrQz1SWpEdhVmQBs3d8ew1WI6WAfx4h4mbAIDn
JHEfoPmnQDJ/D7hWoEq5uN1uCHV2orFDAfRfKpsQhQQqh1OO8Es3G4tHZushit8A6PBQTbPp9i+b
KtnJcN2EXBJG6PGdBQBDUl29KrEe4tVU1s16EKHK0D5qRNBw7hkF2YKIH51WeWnTfXUfvisktzyR
rI1HwmyKQ7jLOVzf3TDbVpl0oQ3/XPkG3lMYfLOIj59RSQ4KRwRC2pfH4LL9pSLHYjTe6AvdTRda
v7skuQSAng8GEkIcn5+1Ro5fqZMIEF3o6TmJjY5C0JKZpU2/7v9crpYRfHQneGZXx7Mxf4TRJKGW
2Xs8CJNLnwswoUux+Ebc1xKDPJx5H3V6DgXNgR6nBRr/6hOYrEbEex0yDafKflacTVyhffEn/rcN
R6KGP13E/L2Jgk377NzeLwi9oV63ox9tku7FE9sn3J+JySrPNZ4XigyCizDyMr0ULmUJPj+y+QoF
FTXdGDF4ohXZhJv8csbFcgPdVTlqKoNrROOMJL2CS9uwfN5N/z40bj1VD3rXUa40h96HDI4hKPFM
hbmjdzcFb7ubUfeN2gEwZO4QmohEIAOfszEjLHX2wWCGAnvRYxJ1ZKGshHtwmv1K5DwgZ44ihskZ
b425hKIVXwFveF8oEMReJMjoPz3qh3QtyFDF0c3raAVVs3lKFdgVksJdplw0Jf/KhxYAtJyFwXwm
hLG65cdNGtqJ3sF+9oH2ejuQO+L9DAGrsA8noA/AFTVLVUfC4jWH/ebzOOAkMORPpsmu2DIEwe4J
QkW5Q0e0cIZ6mOGgVU22tdkmtvWbX7ljypv5/tHSaY0QID9h+NT5AspcpPKN6wVEPBNPdNRP4tZH
R20vWRm7PFt7t7mPiEq7pbneYuLACU84oUXMyf1ZnvUgdhaIeZUWZOYdDGlPtUDq8+IEln2fR3/C
h+7a6UOpYIRD//WE/1QYAFyPLWrTJ+Vy/YP1F6XKzOv1erCpEY1H3qG0ADMlc6RK3oM2qLQIrAmD
cNQvGTBGSm6xgUzVxm4vnWaZtJbVB/8ST4/bOwiWL9oGaLJ2vhN9P/nUEOervxCh7ZGgMXwsA4df
+tTXbL3mTEbXFXzaxobp6cVNe7qk2ebV0sbuJKk+JEba2vktCTAS0cXcU6TVx1wAu6QRAIgdpBjr
cOTOaCUoVttgSFY5SJFIZPEM7+H6uoqE0eKXQ+Ar73WlNB9+e8n8qWrtB6q/3prCtjCPXwYcPLhw
oqUZ5SaCB+kRd/o8xhozZCMJv7Iclys0f11wGT0baRA9KgAe0pMvSVLDSLar1AFgoxm/aHeFOuY3
/ceH6BnfJgM1r7y33UD9ZntRfSajf3qIS9U4ha0zheaEMLltKMpa82f/i/brJBjnua7U28g4hPA9
nOGlAt8mkTWX36CDa/H9wZQzZGhibGSsPqBtmipb7olgY/UIW4yGkDZF3co1l+zZnNzqFb3u3Vej
j+coZUKCWkiIVlOoH8dPoIZ3D2mxDn2WQ0gu10oSAjKfHVb7KXIMNWatjFC7RO9z2dc4PfvOdmub
GP6aLDZO43pntFXtSX7mkvtPET0mU1Xf+FVOlocBK6qMBKWPbx8RlaUoo2V/O6AE3EdujS51xpbG
8T/tVPVGsJxqtGpLZZ6pW63WsMBsBnSlDIx9MvgcEF5HzAPKAEKw8ZMAnKNJdQ+DnADtYO654yNN
fU6pWsB7P5q6cvv8ubsBdwHy4OGDRWfzpRfmKwp8FCutiWGOMd8L6nW5uGD2fGboqrDJ8OzErWu/
i0r2sScwAf5Y9GhixuEKMBlLLQCSDcblaTdmRwkXqQRR34FPwR5n44gmKBLq51mLu6FtGVDfHFEK
BOtt6rZ3ye/dRlx+SOiz/ym0u5eKQ5jdOGqE397D+OLt6NCHB/ICLZ4i5pkgsU9fbd1MhVsquDh1
aEpO5k3P4utp6ocloK7ERF6vIcU8I+kh8RqRI7t5agrXo4x3m1EMvqCfxJo3CN8bW45PuJweigv4
cz8/PbbJupF0Cx3SoiUfi6ZU6DjdkylB0R+dMSnHRK+A/fQCR1hFsbd1/+uutvxVOV4i8PSR+hqi
Ta5Imxw1oE7s5W0AgYzacadJdY+BUb8TTHp9UI9r9SWOlWv8JywZ4Wul2HyIq32FWZRIooPfTGO4
DbdX0Py0BUeJz/agQAIUpHtoh0ypRMiesEkWDSw1Vou+8sW1eNYc+K4wQpX2Qzf6sfX79NrsmJqp
ZnP1Owe0mL9BJfDbAgVn/q3Oi6SuKsGYPfKYPJb/0uk7i1BzLtgmiQKr+k4TqOvX12n1VSZkQQmQ
TGL5AxAIpD9PyFg2+F49Vsu8aM181NsLLt6aSjm/1+ZCQkvWixQ+6ED0iQbVAao5mvat+xXCRKgh
tf9cxGDED2VuzZAHwi+xevODCk7csD8ibPNUzpy1/M519LXn5Ar0frnTauQ0bLkOI6suV30qITTp
ul9ZS7fZMV3UebAyEeq2VKOcEYK1WKyD7eymFtrXW8qYAM7u+P1L1ourEsAJCQjPH+Hz8yy1xMFL
0POsiY8T94vI45ld6fTO3AR+G2KDuVC2OMZvqDwiKximH1cT28mv7TsiCg51Q3JHS7RsTmz72/u2
WxkIzmXh4kfaSdRv7xF1urBADUIcEP/P4hdLFQysduB78MnaQfup7xlCTciWz6C/h1Yk6p0IhNi6
T6ph7vI1NJAn5ejIIMFdLjmao2y4VfRW9fjj6a88WoF5cxAE6IwEbg28ydvObgDhwLz9w68JIi+9
guvGBlFBkQ65kBymIz2fmMMkrd1phqsEj7H2b9RM/empgm3XraYP6BLGUYBWqAvD3OvX/hG2Oh0F
rLCRZIQe+yewCCL9TiD0/Phlr+7P4jSmyVoOoimjrz+aaHvyKSX3r83inrkSuZ3t0noNTKwQr4Qb
g4sSHYea74qbgeD5aMKO8ongrhxImOlrSTPhiChba/PZoom87ynsVXLiQfAYSY9JHHDJVOsqecJQ
Jt5P5FhXscPrsYvAuPc2qMhIqzQIN/JMEIIDh/QQapkCasS8OZEfiTOOycGK2U/IEarj5sunixn/
FR0Xeg17ggpQGez7KSCfShGaxe9Q8zi2g8tvmz34/KDH4wdVqjHo9gphLoEiCtvAwd8A7L4SYMXM
j9O1Maz/O9/X7mJK368xuWn+Acg6Y9Tw6uM381QqpRBEIHXncGeUCsPqeDhSE+eIRyraM5BysrNV
3NQ6oe+MxL3RjZMH5/rPS2oJAaKNAfJGZmcqsLyG5xkymedhLcBfC117HVMlblSn05hYD1ZCGVj8
GJkARZWuc5nev2oyF0xaVAPIT8v3IJ0fGdDckKwVwm+jZ7VzmuPa7N0Y8x4k3h6YHjGrS/sjdsh9
G/Mo+OGLkwV8Qgb3+LBbaD2/pYqSav1/dhXa28f4sCAH44aO9EDrZADfXzI85OT8/sebHAt6Qezc
8LYV00YFTgesD/UlVdExAhohwJw1tm2iLStUu5TzXcdsgpWn34AUZdg8CzAj4RxvBFqBAJZ4RO8f
Q1BL5UI8URT3Y56YOdfY/T5K7WpfbG0AHDKdAwt1OWCqVr5fSxjOdn2QCVPQb+6EI97K6MsXqZDT
t5ueX5InYN6bZlD89qPWEm8TN6mMgfcU4yrR19ImgWichCBt6CgSSxRz2mkFR/FuadmEUtw/5Pv2
Zp/hfxiIbYfkpWnkbdtho4ax+vJyMUfUYMOL23rnhCz4y9ZxaRYkOwM2yX70soj6VHAI2xqs75rL
ynTTbwxqXXpk5u7/HIHiDMu9Z2hfMUKUuemXUCYew5D7yoJZ1bexqzCwxwDIdcPZBIrWjp4AGQaX
IAZc8LG9oO+3YWAKvHEmQghAhwtRCkNzEznp2n1NK3+o0s6r8/XNl7eny8EzNp8S6JaNygy8pPfJ
nXfgXITOWGTFE6TJAVkYdTOaQEnXDjnK3mY3gCzc0/a4Ejj1epOEM4f+n925vPatiBhUikNYmQ3i
ZFq4TdJMJ/IRPHUl4WhMQLaaHVX8OAkofbQGCTTgYbqZE6NxiJolMxq+GcgymSSeXW3xVE6cDLcc
qUWbySHNnNuJri4cbYD1dHTD7+9k3ZznG2fTCq0FuPlm4juKVi3R2eyNNl2sPWNTRF1nG1Bc7b0L
qAW8LetV0Jw8Ye5LFkWjMbb+YUbQTMhnWpwYSJJSgyxSdpTvw2ohEB82bK/OL+jJIUY87dkS5Fyo
yD9p5bZoQAgDWU/DbHiO96+5uJ1SAedjh0ynij5ajX/VI7STDz+f+6ssq+WCHo55FxXF9chJNrUv
Y0nobNiTXx62oWG/tKNn2BZVNjaOUz6/A7c62poucdNNMrqLjWmSfG4dwgWRXYh2yGDs4rge4mEO
xjhVLyEvcyXbII0Cxd7FcjRNQPl5cyPOf6WOGU4Q/RSST/c3dJbe8/T/hWoAcLtQrHibKFE6Pzjf
H1RPTYoQvtw17w/N1mo0Py4Km48TP+HobWsXp6F5T1pR71rxeWNkMr1jPA8CJ+xVaGl4UKF01Ukr
jpQAPgKakcCCg8OaVmfWRWYBs4Q1yi7z9IChHWhawiItyyolA/LSeHNZwYsoPQGBX9oI+ZLaxJAR
ICUJE8tlP2gTKpK1EfC+iLvOlfOvYuddD3V3LB98xA9PVZ7ZENxnMXEREgJcLjtKR1N/YLhuvmc/
3NegnKdGDBATBnD8w0s1/Ib8mhTE2AHfQ+t7WGgcgzo8risNexAgld9P0s2FbqrKfya6HS2aviaT
paJXHZLg6buzImuDA5FzHxOiJL+ROfTp2jmEzbDXgHNirJbe1HJynHRCtYVZBszcnlJV1PWQuWaM
kumySBUhTplLW66xQ1UeI2dFjQ0HP/bhDVF4sPZl0trF4mDs9bIik7fI3fyaa5kYBAe0NA72hkBA
6NMFsPiZjBqAxoK283Jxs2iO6JDfYRf1BhLbdMExzgFSS1CjG2Id3gvbMSUDrnl9WAt9kqqcYMhG
NWmTfKA/gEdyP3q/QODZn7KBPv5gZq2cc6qkUaBU8sma5LAvbvx4FxPvADSVBqMU7nLD9RaVztl7
gmNjHCQrhzfpPhoCA7ko9h1UsOA2hkY3BaMx0z4Nd6iBwfWOupfnVjPRZRMYhIihhqsRFleN7sfE
MwRIlGTnoOw7xIAC51GGc/gxBey53Lm8QZ8I4I2f3+HUgRrJBnY9N8lmd8ZmyongzfekzdD0CuOA
ptn+q1v95uBH82DOoEWPKXfJuHp/tUhfcEqKKv47HWavBLBLOz62PwxiNfLkfYc1EV+fvtxIWGPe
LA96AWC7O0kjFqshsBO+Bu7wp42Lt6Am1qMXOheIylRowyK9AhKjnpMJfAVcoTciZY5zBr3XHgg4
6/f2oPbRhvxCXdmk0IDbS9oxRNbi1eqaX93FEIWu8pYnCHrnWYt7jFOhx8TNJq5Alq1c0ScsFKqK
GF+64wSQ5rZHwhvM/nDEKxcrK3RbS4o/Dc9I+C3py7UcU+Plb5y2m7vP1+uUABVh/Yr9nyEYB89D
ChJbXX/DkOs3WqeqZBZ+Bqu1xNFVVCoSyAZbRDKLuasptz7jqrwcCztHyxFrzPF0kbio0p7sw9TO
HwERuHrcpupu5bEjbMW31oOB0Lk0OOw5jLa5u8B20TSKEhKXpPiBFvX9QiMUs/JrbPCQUeMUpdgm
QBPxfifpxFdoF8ODioP0ZqngE60Inr9swOH6J72b1s8GwSoxIYdbRhxwyn3DanLZPF2CR176ZRWo
bXIc8RXjes4CtRM4mNyzOuHPVddppOFIWHCzTHWBfoY5jHdzvYGfwvc1WaRvkpzmcsItxSoKVpM+
RjrnTvkWDVIu0Kql/7NroF5pXkfE3DdnOokP6i0qmbVNougmcO9NbImUbxLJuWYvRT+IvuyHf+s0
yRzVPqusKvz0j5vAMHN5sp/PG5/g10mTio1OoP4ji9F9j2uVH7vgvSJuQsakc5rbXg7fcA4j6IrA
h4pxyxU4h0Z7mikcBTHCAmr7nX43EK96tgL/iq7QdpjDCq8JwEp+Jv3SEy1XBk5eKoK/OgOWqM8a
ebDafz/ny3bNwsY0saAZ9ICLmMGZEGvZsUR05gs6DcjJzQXGt68OinUI13I94f3rQ++F6kXTiL5a
fQ4RXvl+dVWwZcauR97aZKeYVAif9jno9S8UdjMYK2y40nPyGX8Cr9zVuyd7TgwhU63fG39f2iIa
khYTLXJ9IIHYf0v4+bSaJa0aub4BblDIHCyG+wpmhTcmYg3VUw06JzOaZxJ+vi9i/BJDWPzcdTTx
an0ASpTS6nnWyCkMU0ukABCzqZ8BXGC9YmqqRl6Q86ZzZjE/8ZK+iKazZzzAACOiLeEYC7gSJLgt
6KlV4zzFAGuL0HiHc+2QQb02d7RgAySd/A8v47BzfXcUOym32jHUdzvYl3PWC9uuxucRjTKlIKQj
uGsKdA+DBEz9usp/5IRPCJj9wLxa00pXBQ+tXMAfmMCduUIvmEyo2xOIbo2XRfFb8UeFEGJ/RhTz
dn+/9X2ycbF0C0vxspaLjKOf6yAe60HWfjmOxs+qeq0XksFgBxFOGz4iExX5HJ3O7rNJ0lDJemCe
9Z2s2LGTveDvr8X6jkkGOEZhfuInXMCFejPlR7sKDpHIH6T7BURTHlVFtSXQ1ijwUHxKbGC6TTej
j+yv1GWNFalpKiTbfIX3AoTlVyLthnrrEmMn4liRqVSYaQOtOGrt7bR+G53E7Bad1+wZvNL1NivR
7N9EQyRKt2xnnLDkuJ0cwKoIiil8KhSkj/lnNXisCQLdETpzutK9WT+t5qw3awtKYXvAUOKgJrI3
9TZPKk4co9W1bbOrjBADBLpiKe9riRwuigrE8CQbRZ253XMjg4oqHWm00oggKavi4yu0Uqqmow0H
qjkBhWjDdh9biARTH68LMJexauECyu3UhX7mI5Bwy5dS38RO+vLgbu5p/kFnNeuvreAjhUdw3Z0C
2uLcv+7Bhi3XzllDhsJ/QYVWmn2g4n6iGNmnzrWbG36oDgiPahBpGGhECbIxsHQO83CQgLn7DndS
7Zn5wVnsWZZ7oomPJaCUfexUurVi0ubvXCmKQ2otvxuBbLKqqC9QDuZtMNO0OK5HYG81cGh9ZwMR
af8TbJC1x+2Gl1TrFPmjJal09HWuxiPBFYawHeaIWHYM8xl18yqAe37P434/pUqK0tM/eZbrh1uE
3x8YLJozocswP7PUX5yGb6QYWezVtDmDYpkOuDQsZLRfMPPhc9UGqBVgXKs3vJubk2ju6sMLzzAF
3gq4lgc+Ps1Y6IB1wMepMhPSr2Op+nJCZvP3x2jhlH20rOSrQNURjiYpLpdV2k6DbznVUGtQ+ik0
M1KNBVSVrXJXJ/qr7wrn1k0nQOmAw7/ix29hvXCeWuIa/JmYBnpjCqK+I0y36B8UhRIM+9Brkctv
mrXjJ6TCKTqjFD7Y8hCMI5TkCCrcKrDx3h5TWtKUk914ADECoT9NXaK8Ya7845E5Ass+/sdQjbvB
0DdK+eJvKXvvyqMFUmDeafvOdUt2BXaAut8wJK+Csj6VVDj5uAyBxQaLeZ+XLXuPp7634tE63SCx
B8jzXWa58RMSnhnnpk8Lb5MwCEsY/OwkV2auDhatlnJTl6DW3vm9fzb3FE/7sXpPsrx1vTo+xNQV
htE68u/xDcwjT3iDk3GKcEqMMXn036Xsq6f8BFRb40MVWY38yA4l+PuulHqtkdp08Ldo1U4FnYqX
nU2rSWViw9MHVkUVQmBVs2WDbsfSrkBvno438KWTPZzsBlsYcM0q8aLDdPidOUBvYZ913+C64+Zj
0sW5sKeE9wAvgTUSXhbUee2ad0UJjB6ekXpSb+bnhIpCBrza8uZVhbqBpH7+ClW3iOvds040O0t1
9a+swqcELxWkog2hHWYcM70GsAGeXuKbtmXjXn7QC1nxu9yUF0lUPwXDi/pcmDo7dSGUqBCbqo39
ykmXqGysnW23v5NRQV3PkF+5a7ogTHBAATJj6LqqNa+I3RUhGTr/oy85NdYzbAfYu8/rYj+DihdR
+xh/B/ZN6VkRmBe4XHjI+b55dQ163TfFKCUdLe7frRMADJC5iVtME2tnypOhOOv0Gislq3WnxpMu
vL0xygNaIMtrrTp1Qcys7dn7mxTuN6LDtkqLXMmNygJf5xN+dpwj863P2eot246Hiuz+05Op6ezh
TJk9dTivuncDNkCiEtEhIubsEmGcFsNE1xuzL/nvIeWquk1emw+K6aJPXpnhVKmImam7kfVFEB9k
lEaqIYTtBZVG2WusWtNjW0N+gGq3zVi0XXuNzTNdkWALTc1HfiUDH50lGF3ENQcVDT7tqGKFuS4D
/T2dOP2bgEQ5FihSac01jNnC6fiqEolQBaYf6ly1FtRyJBrQcPRDMyxS3eRJxMkcW590RqmI1Xk7
Ku+ahJHw+E9rTeubzzJPMu4xfWjUXrViAlmcYQzJKUZlO3uLJWDzjmr9ROx5qi419CxInEombKwC
Fi7ET5rlfK2NUszBgLa8yZr9X60EKu8aN+gqBNUkQGVcBGaQrrgjVlIccrRArR1/Wzeolm4awoil
ytbE5gcxDTOfpVSb8ZlRUtcwJhlE6Awu4DMbycqhuo5IJDmxDE3lmVIPK5niQlIsVEWm8CUXqyPG
kncmuQmNndWQ2nSWq5Bwh7ClfhtcykC7+puldYiaaDwzBEJDaNhry8jAVkJfZ8/rTqcU+JSlOaYD
Ihpu81WVGfNufF/A/r3EGX+MZJbXrKokyc/1aT+1ir3FvmCaSxzxOaj66vW/cQ3fMYW5Sy5/r6iA
yIZ6Nyp61B4TENK7KT19GV1PNRyzlxfzFVXyUYIkVpNvajIR6Zw7T6gqwcync6tyOL5u9hoWkIdB
UPVaAswAe+6GHlyY69+8ZXEq6IDWGfjXO3rZaPaFyj+lLP3hY6YCGQ1hB+zzZYwF3OMPaCss6D3s
Hd9a280XMA9+skl0e6p8FeoGhVOeN5ceaRN5oFYnpAxOJtnPYzu8qwsTEI9m0w///qmpKLupRqJF
RJKFH6CEwEfqbo6uvn1vr2lk0HIqX6ZNzxCisUBrCfxo1sMOPjG+W9FBtLOTU1OZpe+GDXfbWM9k
SJ62s9XuYpUytAw3rpVZo60mRESZ7QK6KxedrJXDANfEb5JvHXIvIf3MgheAtcDTHM1x5DOVCxmL
dQMlDZ3ECKjBqymNx3jypqy/r1Bk/X9WEsnm1pFqB8D5QyiByzEVAvYv0sDU+AcG8eamIGklvUbU
wvmvR9v10z4J674hf+1iQvSQCtgMOMrfyY8Pv1xfRL1XIm1+mJo1TFeMIeZSwqUjUXtBLdJkqnis
cWbAr8OXyjDIv1cYh4XfvTdvxKeCKI43KqFKro6yqSJVMgYUtDZPJOw8Ghaoujt6ge8zEViGh663
FBdyTkaV8oZfFQLlWOXpVyF9duhhtRU6bg/IDDBCet12bGRe/MNhaEKrALEmhSjTOyO+G157sXfa
x95SZBvWcA69JrXbaVgWBg+ZgS3VnqwVNix3P0zV5LA8ewgyB9hYf8invh+Bp/0xPzTjDWfjaeh4
h74Lgom6s8Dp+4fUY0eAqkuFlrv+1C9AJRVH26KDg6ugrDTx0hmULurhpc6mKAXyI8THbhrblrl/
UGOdWHJgiXNaUQQSw+YNPPYnmNiy2L0ml32v52n/jgtlR215GNffN9K+g3LQ3iVahk9JPASmtwcb
anF9Paej5xmMvcRvGkMzuc7Sll/4U2Rs4MPDtgeDdJb47HCyzC/Lpx6UaHiGgshJPkk1ju4uP1Ce
QKzBLnTdc0N6VjUjOvuHDQCHiaZe51fRZWgSha1isvwjvahRvmCkLL7U/aKKgeeQsi+SakgjL+G5
kk02/LZCLHul+kyiPNATcE63Oj8hurr9ytGhHZPdM6vprzKaNpWhwY8iZzCeDQVR8icxJ9sON/OX
CZCqwkyJ9gG6STvfu7VoZrQSP7cSgjJ9WSnod7x4wvsPv54ZSyUqmQ/3PHxbaT0aZexM0lswmKmL
pI4j1zvyH2E9JRUFwiaD7t1kWDhRDJbqvLhsqCEPCHWKkjqCUppK+PUEdAQuXiYi7WxcvTEaHumd
oAUCCaUj3/lWWMxLVSjvbRqLCZEcnFQbLJRflIPisPQD8AS6PqUnP7rGz+/7q2oqc6cWeiNa5egE
tEfE87OLdq47lZVT+TVCyP/bis+i6cChA/BW4q7FzZqp/+uQCweATzZQnYzWkFhtjHc/EjW55Mp1
14pYKF6SBlGWauGX0gxaLQpXip3/PepjPrHs2B5XvQer6AlXHtsHPT2JTkituK/V8QwdqTgJ1m4d
Y21z6zmWzDEesUOaktZfhzJPXOLWz8bcNRCrVvjN+MdSVvqSjYc/+odU6DYnPTnShOj8Q/Q8YpUl
KcZvYRot2Nd/HfXg0nqIL1OaA3qeF3SneGViJ9ITt6o8Sy/Qn78AmHIhDrS1UtG0gNm0VRtjvCii
9R4FpkewbbUxFk2S/QIjQK6xgIbtXKHjSVl8vkpDFh6Zfwi9aXzsVdu8IVFexE7ZSIh3WT9QIPQR
hL1obJ6MZT1CTBLtKfL+j4qhq2M+mHYWJkEHwd13haXgOVcO6GDsv5/rQaB+10GZapsfJ3im7Uap
1HOzHftFgDms5ITEOe7SfJ8zqcmPQg7jt2S828Hp3cIbXj1cFE9jCvp0tcf5szHTgbSrtPoK3n8M
I+XxRtaXKYvApr++W4ZEy3P29KHPoZ7x0KXEjhywPcr8MsEAHXUBgOHbiWT45Lm/3l26H2J5su/h
iPXLhrQNeFoIigGZICAsS0O1KRwsVTqhMFvWOG2PySk1bEDuGZhhwdI9m6w3Xc77jr9JTKscy19k
fDduL4T3Jq/4xF/Oq78SSPO6PYrjToOpsUPULQxgtFBvRJ6ztQYl3ieIsF5by4E9gDJLRg5NJ1eW
ahXWeWwpjurbvedlb24FmUW8clGgP+WuixwTmr5xQzzdh0mrokl55oDghDZdT9sRpEMJ/VD4WpFD
dG39oaIOKp2tmEAN7mK/RYwXNgPgjYhowZ9BP4gElpwh6Bv2g1wjmVCEusHnMhtuh9g1GU3t2alN
+g1Zxc3/WptwKniy6ohPcHPEvdEB7MG5Yqh5QdP7NpukJdYLjIp1RQ9WbFQMlFGdkrob44eUki+O
YUIerdhgfpfqrbSQhmn+MaCoYO3w11d+X2X0I0qZSgxvxnCSWRC93iau68IocWXzRd7N8HxqRYhp
sa4uCyCcBsEMXw30KnYZQnl6s0+/qCXKIyqf3naj6p8vfMpBMY/PHtz/MeiPu9MkMT8P1XH0fUxs
+BZQrvfafXSvuvA67VZl/rFdUVOgjKnOM5sotq2mfIDLzSWi6DL365wtk+2YHBfgukecFPxEBTcs
h0xqPJMHzk2pN1Odp1Y9gR8Aveibl1tXcaZHHirdhLEcAH7/AGLLsRAutjBZ4sE5jEr3akznqPNt
ozvC8cxV3IzRJth66zm2B/8ggWFLwqr2OFP9Hsk5cHhm41BJFvPAZx9yl243OIFudkDejlFDo/4V
wG3sH6K4fHMvFXp33NM1se6ckip/5Ylt1Rx+NPH7VSVzXMysxhf+VzSHort8azg7rZhat1lwlwQe
p1racbqzDHx+87IVyU2NjQAGRab8dXF7/9A6F/9aik6KDx5uuGwEqtZtjW2tsnJ+BgRklrSYc9GH
ftWjWBU99som/89Wh1FFMuWtY0I2cyL5tvOWizF5ARG98G/JArwabFe7OHkqDHzC6MoNvCvmVaYb
iJJaYrEW0xFchJ865wNCdKH38Rg7p1ACWYL7lvmaEGZoyLthj984HdcsK6GC1ZxbFvqgrxJXhOG/
/hGiI382GCk/H43199p5xG7Sqp6qAwbC0ifaX/IFvjHTBVbpHdS8as5tq221H41k4U//eRZ2GWyO
RahJ1ozYjeSOER9hNoZJYnowzuT8lFAPFCNkaZoWeLsTNzSui2dEDYKn+gwwBeUqTdNRUaaQpPOt
6IAxZU7PPgZh1rXO5u9LJYqRmY1VkT4vVMzSeFmZJlPE64ee4UvE/7ng5gkPQLAFjldwelQyubRV
7WKWoTONwqj/N641QJoa3TnEetKRMVGJ/k7NQ3F7O5PwbIKfnvJ6ezhG/DoCft/fAGs8WP/5Ciaf
Vx+D4DwEr3boZA2QhzAtC5t0IxvP8JqIksSFgCHejvBc+5cRDxyJlP//sezPurpz1aeMMXEvgI71
UQZ1pnjAZbZXO/q9ZCAqWa8EMq3luuUC/4uvhxrc39KHNt7HaRqaJFxQtAeZPhG7PGaS/PETPKyH
gPYmsGR8SUGMEQjZOGyvhgZNAaoLz92i6rjATcU4AZaWljfXMH8ZXkNyA68mkXg0nIWRhoCBxVXd
R9D+nAwzpz8WqDp/KtZaqccp5tAGoDK6BRnVuCKlZtLDyQuZIAMQpUkc14JCorna43kY+fbMxTEe
q3Mj0m6jxIsIFvJnxMv2teebEqTZ6xUG7/Emxy4y+Uh3crH0MgU/4qTiY7LX5mmS2NGdGbxAhqQ/
i43q6Brlr+H7bhjLG2CalFwCgbjVosSFK81zINkVRiZ3McQszmbZMxSbOzulMgfc/cTJ+1p525hz
phvX+llgNEHdUeM8dz3QQrzQxJawYTERP7P1hAv/FO2BeSWnG5IMymjrMOfL4PxrV/DyywLqqkPo
4AQ0J9HEBKIZY9CpU3TsgP4XE7QXC+egsWPMWCA37Qyb5YGd3zF+ppeYpa556qhBRT9YLQ2HZ8Vj
r/aKK/N0yWvQ3J7WZIIB8kQzDNpB4+iEs3abFTKzJIkJdBvVZikkiBDwKF27fap033B2MOQGKyAL
ElhwCsk8whT1mOVY6gxcHBZF+jcpKTIRgD44vE8EsFvrihz/3Jqon+GXMQzTARfzZi32/CQoY6ES
MAuLUXa57s3MpP2hz1Blk0Wz+nY6UEkiMODFQJmkmHYJfB674MRFOtORsy4BGCIWd3eolLQ7MOwF
odtZkmrulZqO40z6krXiz7G+WmhmuAqAjvq1ujIxHZvNm5967HsCB82D3S2gbgd+rEhPT7PWNNmo
dKaBAJtT5TTaxnC7jsm7nF8uXbzGre9HDCYMKhhTAucJz9J90W9CYzpYC94u0XqE8mpLVgTF8z1q
VSPycl3WuqzoES64xPAjdovJwRGIu6pKbv9mhFH+Ibmv5AgdXIl18NFwUm5nkhU6T0Z2nHazihRA
i/DlO11MzEhX1xV+3rMGFXwF8y90Hp9KHERDaF0s+553kUMWBoUAqqBci0jP8DBap3AqRapCbvgp
4EttKWXsUpByZKaspeWKxxFOx73HFCZop7MryVYcLU8T2aNljwVWcgX4+U8QJ4UMfgV4pkeFkVk8
PWOAq62pJ5c8XQUlvxjnS4tnNE39YUnARabmSPfWTuOu0ncGs9uw11dl1c3ZqhX3CU2VXcDD29W+
ftTzZvbzv5vfz+f+9e6mAjJMA5jI5uDrj6uqP4UGBH0HJfnGEtPWkTrqtnzDgPvAQvjz03mrD450
wmMLSSFG9dT77qXohIaHjbQ964MDoLinvVtPYnda+WaL5OEAWj6w0brYqOOe1gs1nq5WNEhTXB27
NX1AgVvVaEGmgm1mRsNvRVIXL4G+QYCXs/B6n7lBYRZf1an0bYGg1RaRE0r3CeuKD8B9f3tmnM9F
v6uLx5AT1xt/DP8pTVVLOiRadx9weevDFUWeBAR7+ph6eNCNqd/Vj2cncW44KTAYceY5nvuvKRPI
X2uaY0wWR8B4sD9fOLJSqR628pufpHX6OSZTUgXZ7boOv0Y0IYVtGRdcz/k5C36TqXSSgyd9oxUq
0ATCDrk20mo7d+n1AfLO/Gkz8Z+zVE68V5qoHvREA4C8SbSSdZ940tYG9Cvqb2Mna60AKLvfRQfk
0Pr82szFKg5xhhuweAyesptmAiBuFWpaCs9iAQIDmqmkGitQxsX2dhOeqBM9PHCAAJxMj+4JRxEx
AfvMg9pfUVZLv60mSErTw6edFQZ8ZbXYWM+2yS/F4vEkdUVa6aEf826D2wzlFon+tsxLM0gq/WsN
Ka+tC3qMBjKo5/caIu3NF3EHDQ63wVVdwMmjwPefB3A+vPzgd8iVxky6vYm6Ns6BuWDThVqbSrS/
0yrg49wbtS1MZpNDDPm/oIKeOBdj1o+4WDQTiTm2pDoWlA9FF0MlNvUh4hbTWbaAQBGxcUDbAFnT
956zJybpXDtX28IpFhF7XNwRIGBsmdYzUKchI9g+TzM4NfTmcbjFNj2S11XWZYtYYI6ERptWhYPN
t51JKMi25tX7vefKl0OBT9KbuoKv4ILWOa/TVlndGkFz0XbP1/Hpg53e1PPZ/CXxPAo0wHrU47bU
83pBblkcyqEC1jzPAZxNAlGqeRAKZ/gfpXsdDYbIIuPX5J+GcC7nI4vImj/LhsMp2Te6tQ6ITML0
JCnhR0ImwmFpvk3vCwdGr0XKo8zqNTOoBLg3eutxQjY/eFJzUX9To0/on0NPLK3V5RJEwpj8pj3U
NdkBguco+ET9UW1qJ7G37aQKv/2cChThLP87b+99wWdxZB/s05sLrvOy52iURUPdTBG/45oZAZTK
EsgqDbCUFQNs2YPcUjEafvtn/tXLXST7AbXXl41XWz4PZ9FKHUU0LjZVLeyZ6HkVq1MDq7iw7Awv
fxbyhpU2v5DprtS/QJOrDPjEDgaydC/fdRhPEP7wx6rK0j6CK4JMAXgLqjgDm1wZG1444OxRLoka
R8iv/48BKWFz/Z2DpMHq96oRwrsZ59ZxlzA5V/eu/L2Qp7eJpHjskarFlOUPjKIv7Fua1C7pkabl
xqF0A+w+bv2yiJrPi2BThYL5Mq+/pRJ2Jn/4GW9CQGn2PvuL9ziqeFEdjHH8w7g+redTiGuWJ1We
HMzaVwlme0Pus3F5Mp1m8nEfUoWbnm1nJiBfQUcjQuYinKnsSSYDcEj1SnibRDfShku+MNBHp9I8
X5t5sChd98nUMjArhgezb12CShfBXrbrK5NFSN9TTKPGb7E7DjpZglPM7SSchldCYJAJdK4Nkdnj
3OdVCPqleOaTzrbOGqgVc+v9scf2U/2NhjN7m3U/kQJF+VU95l5KML3o2Bmqji9PbEHuOsQr9Wtt
DLHby4yf4aZOEO24CHJuDV6Nik/Tt1tRI4NJclyyuSyod1eNSHRRl9dvz0OtuJVQC9il6N5wFlXN
kUB5Fv3GFr7ICT2l+mLD13jCCuX9gx+dGlRQmx/8Fn1g67hCpmQoemYqGWq4jBzk9Fftc+F1recA
8R0ZO1cei2OwEDqQfv0mDwyxn9rl09SbyfU/wsK276qRd6qLHBLbU2JjyTUDk+LkzqO3EBgPUVOt
/wwyzAiBFrwbmCAO15QLrx5tEZhJyYcPRMzk7e1yok8sPTHWMCsYQVSzJXuuDopaEC7hUJoYEm2n
oeobDgs4CEsZPWpV9jmslyCgkjQ35JjrHMxdqwscDBeEr9MSHK1MO9qtRwWT99rwF+Gv+77albH5
9iZxMOHFWoUG2NMxsaxRbJh4WCh8LR6B9NUp+YExYi1gr7Wv2I3GO7ozxv65Y2q5QnczC1NdRUVA
k0Oy9VDCsLr1nwAgY7I8AhQtRPVyDuUoPDC2w1BGl9mMoq20s7qB1FJ0i1W5v66moglvgUVVk7X0
+QGzmMMQBNJgFOlhg3kO/pNCUbUQ/Sh4CJZ5eSPWWnhmObQOMyVUURsjt+UXBDS/B6ZhEulClV3d
V2OAdAgDRkKiZDelyoURg+pOFfce6Wxx1Hcbzbm5g3BNJh6GTbGYvOWNc6pcVAhb0TER4FhXnuQn
jB/UgvxPDvAZpIxVjmHKO+fAUzvQdA3CVlJ3NaQMEHS6Fiw/YnpYoNQqVqbSjYrM1YGEUZbgSOf7
ecZWcVGTQyJ/QOUodfx7CA0rRN4oP5lbmEJwaCudHp25Xj0DO2VTqu8dEw7WB8Xm7wR9zr9ijnFU
1wwNOK0XTW4s+ns7JeuMHrXevp4CyHTjOy1TdIOEZzVdAcQu4FiVCiYEzls7UFOabyw9+wlXNgMy
sVACWgynPcb5j093IJcn7BIGJ6sZZuVozMgBl5GzpeoCisbqkxdNtQPDiM61BNQpuRIJJ92yxICW
DQ3UMjELS2x7a+yfcgZGJ/VvAEFcq+UafWtfK93DRI6umMSrlEECAYep5X9gj7G+KK9kdiAMvw0j
eRz08R73lbL3Rcs+vORJiMkrvTnTIvxgMuRrQ0LH2Rw7X5qMKGOBsZQAYSj/9iEuH2bX1Q0NwxjW
UGbpqxq4U9fw7qVO9DC9xhFkI49F9qq8/qNIo/waOoJ6ZqjfCFbvfpWXXY6nV5vJ2zHUPkScSAo1
pqNnK//QZJufc2MbHDy1559qTMdLHHMIj//h+dRZsgnsCn4DHCt9brTrByjmaKeHgSCp95oJ2PGu
FZ1tqxHr8kTLVQ288kSzW1z6p6biEN8AvXT7Ot441H8V7Vr36N6ScrDMJogySkPB9wLQTz5Tgeub
xyHPpcLkymjPX8p7tLpy0jp8e9dVSj9zmZyCdnL18HqdoxQb6G2Y5f8d7OKvshfY3cf5Po3g8gEz
o8k00O3yYPXzQuWZ3g4wPcUA83qMPV1bCZ327mnhR4HFbsA0cRmeQgx6PqyIQMPYmr+1VQsT6DzQ
Itx+URV1BxSP4SkQgJ49AYDCELWeP4jrh68JMD5rEYGTJfEqYgbh56SZzVWqRLUv1mXYoNapi+89
sLtRpDZnsFQjbMEtqjsHACL8t/tKfNBuaoKFP5rgj2K7SjyWHVR/hxt1feZf8WS2VqNypd3Oomkw
Z3Dc9f8/pS5D8510rAWiRyRgJlpjaPJZb/DOojEhAWucIwLu923KGQl/SVV3bRBZfiFuWm8KgRja
y/sgWHxcSfOj/uEyyYHEu1gcy65PzZGgRNLMFojqnLXyLbC9gKOZmsutaJatc8wLsJiYt4YGfzxy
DNNjt8qbrHkM2JQE/Ukq9jRPOhZEaFTS6zgbbNGOeOKVWIuBtRpx7VV0fTUHGusvWlDN98DLjsvK
30cGTzYJP1JMDruSVlXr8q8ZxwLeOmdDzdPcSafQ3oVOLgmsuwArFFlbm7xqhz/9voE4T4bbMeCn
EuADoQAIdSKYVteAfw5gwvVVCir2U7Z4V0Vt9nssI05MuNfRzyj60CcbQv/vixfzWnJkOWrJGrzt
R5zh5/HuCYakWlarepTuHYx3iomkTg3BPNkzBkTzqs8jOwGZJih3c3J/GDFb8ZI90/K71TrhE7Uv
Qd57RQ1M4RnIV6dGE8+AFDBtNxC141lrl14PXxeRhef1vZJegCQCeK7wtnfNec4HmJJ6kFXZZ5lN
l+gO6zdPGBQNlJ/BeloF7PRN1xx9byDY0jqM/ef1o73DY6sXqqbLJDAzr/V96DJbdZtChj+yb9xO
EZzzG3arOHPZx34fDiSkLw0yi7uCvxmkAJMbJ02QTk1p7AijFclCy46I8K0oraEBiFgIublVIuc9
p6kLA/GqbbY3D0jterHnSOTEMsZIrPaTMSzrsWAP3mqf0zM1a2fZxhAi8Ec4ibGPAZBAjYMlWUsj
O0HxFTkeWOx0wWdmAHWh4rGPJ97kflkeUHoayPSCwYNg38Ond3Y6CivtBTkTpiWqa/AuGLKT6TOz
9iSNTKKbyLEprg/i6xOjnP9YKEdH8830Xv3D+z0ulMUiDGnII37LjDIwIgKM8CxeH1gAbU4CWuGp
+YZnb0k3yHDQyfldPF+TWoOEMYhzJH0EXbVcJ3U2IBy4SsqjcDC6FHQUgB7t0ssw3j44dxoPWqkj
M85SScZj4HOBpJ1zKxw16oMOLQExMqVzC472IhMRk6FoiC9VGYlu59WpgY/UUzgpMZQYYFwJTIsP
7TzuS2twLBu9g1+MkIK39jOM+q3XY8ToyQzRbd+rQ5c1A/mkW4PH+b5qZtH9QVbDADMRY3pCaaFo
ZnUmoL2ViJ7hFWeVz0GRf7gPTqR7/QEyj3p2TY1K7n91BgOPIuhi9iWaR8CcSMhUe/korJ3mJ6c4
WPhNFUxyfT3CiXd1u6J6cChmQAUekI9qCbpffPn9vb9hs7SdvEy2LOUQIWNiYnKp1fg4PpUx0l3y
3Ytjek5kQCYpefpeBs643CPI34T3MH4ZNvO0MleYlaSSjkTW14jiOQzCrsJfc5TkeMqxKEk7laQe
GQnqay0LABOcsveH21FzW3wSUc5kJDzkowtE9fpv5wUMcQb8GLSj7fY5eWJFDLYTdOOmb6+M5pUp
T9WImcySzdjC3iNqFCro8QhH2o/FeekJ4US4vEhwKmYjuIw+SYxokdybbv3BJesrSjT6AxAEki7U
hZUMjYxNedN1Jtwm+UfvJ+xvRjBSFmBSsU+494Tu89HkYsPJuEePJd4wew/b4UReMQn8nx4V+Ulq
NQ9jg4PLCWczmNUvDipOZ5ZuhbLDX2OW8IaXm+nQxOlx17mOxzZqDqmAVcnDxZs61bV6aUKGy+Hb
e0VEDDPVirvM59dlZVUfLxwH3c1TUbUKkHRo5XRrrKKdZHl8VEJVB4RoCL1Nwc2Z471kTIz1MBBh
dta3En/0fn7onLQLUrxxf2Zxqlj+mDlon7Q4EuJ/vkGPXgU+MjWMXkTtZJiNrPjmijAn5EhQHz/B
B+lPAORRi8pUD7z6EPNPzHUzK9pxYeBrRQHEAlNPnEtz2Swomi08ATG5bzSWR2vG7hYT4PWAo4AV
Zms3ITRIvYkjJ5MJ7sCKsci2JIR9eDXWFxEz4EdWe4HwYqUP8TOFkY7QKHtSeYvuwAVe9xhAd1aN
HC6Uqkh/oTamHk9+KFdYeGfxvgll8FEajeA7uiK9+CAucd8pS2ZU642+tFg0EwZPgaG8XYBMOSET
bzTxjYfv96rpnWVb7jNhNwNoEYZCUASj6hxVV0Or6nGw/9fTq9DNJUlG0QQVZSImCmFonNeYxBU9
1k9La9djjxWEikEmJms1XO20YnhjgDG2SxoRjbo49IOZ9eG3yNSBWGI8NbE7SMPWDg2x9RY6y8JG
BBDUOdFb51xVlmcdcI+s1D1R4BtHq9slX+SpgXx8hJtr4LISp4PlXqKyOcfmnIJXm9mThEH389Ir
j9mxi1+2l9+09y+AnvIwZeMoidhVqQUJIvwJ14ibZG6eE6mcvSEOGbnGBadGxzEn2mfqySxCen7G
lQfvHntZEgHuIKtDEn1lwun/C5/rxmwmV+act24m+bTfPJA/1fxLkf+t5jSS+VFoivsJFxymyw2p
Pl9TYdCAfedBdNDS7DkO3F/EaW6ud9ZfDjsMCCwcpwO2jzCj8KDCA5+6lnBAzOURif5Z3hmsASIn
rnfDqUK82yML5z6fNvGqh8pyNvpJLj4RZdD6rxQZzJ9kMOot6X5CY5kElklFVk/j7Xffrt9ywg6q
SnapORcsct7mxRWLV91BORhFByiZVQDnICZ3DC30b4DBdVA6R+FU9KxKUXoVGgUibKpNjBeLeC73
wn6ma2In+fyTVEa5tEis6I8uClmvApcSOFNa7Pzxl56tRj+1iQVVJ7Q9VWuQEMEg/dD/GRsHzszE
xWxgdK8thkNSHNqUZdOpDwYJxGk/Cc/xmklbj14/MjwAKHLOV+xlS/D2eZS+l2OaFjF0PWMDOGXk
L4FIWb2sJRf3tH5Em2EqO4Bvq0xXVSRRyxdhQP/Usopfy8gf+kSiZdTunQlkB9Pno9WH2hYr4T11
WiYavRVuCDOoao9LtogsfIaHrBKgs7nB9QK7hvVUSyyEnt+Hi0iWkDV49ZS8X8cAXSwB6g7U6aW1
6ZcjfH9/ug10N3KHTnsQL1ldtQ+Pm2t66QSR0bjOlu68T/BJIXktqwoYgB5TmPSYhXKKKRKDMmrP
LEYmWsdl+u3K0+pJdSSoPeA4Ts9/+WMItvK8KuhUPPibCCMt2+WBKbHnS/hNebpKVjA9Wtxq2cbQ
Tvo/7GXJeEj1dxVJjzcsgIemxuh/r0pMPdpIbFJngEaguRNkuamX/b4jTJC7x0dEYmV1NVnrYWky
UcW8AYRRup/baRYmZktvTLISrHHPjcTkS8dkabkDk6uM7Dkhfl7s7/YKJWYGgTLTqRhn8fQkeJco
EbUfXGFLq8L4N02rE8pE9uD+WWEvdvVFwJZ2tYMeOJCVSv3uAtkLAOxhbGE/Hq9DcnV7LxReP8ON
NZdxTog5VfMnqcWmyJ0VmeG7wBnMzDnpUTJ7E6g2q4QNGG1Zqd2r1sfW1W3hU7A5Sbd/qZGnbIRR
/M3bJY6JHQfj1avK2doxVZpW4Yve2GAx7ciycNCDRir+m+jzR/lMI0OHYWP2n0Vh2aDxGBuJE6wB
EkOrq2E1H5rTtJHIJXP+I1/8/S07YeAs95QY+cyIUUZFOeNbK9WYnv+fAcrjqlhjgicrZfS3ma+F
Ii6ytDVq7rRxfvk20FMMcV8N/n1209SI6ykzw+1WXK76+cTd4QgH4jINBOUgfzg7/0PPwiLQiIcE
9V9LvkO/ZL9SfKmdVGIIJYOCKbeoBiEzS1lKQHYdbYE53xacZCszStB6mcSqUe026IH3XBf2WCfb
5VboSXn63WmvIx1SXdt1cL4Le6S4VgKQUb0joLqSpasZ8mIfHzWv8YHdCcfybEjlh3zFGxf/zZC5
YxWDD02P/oJg/NB5yOJvvmM3ug0QxqMxuFtFTejSur/U/e8/PM4Okk4TN1HpB6vZlckUWpFhjuMO
i83ztmc48gNllF2ZBHFfqNpZkpoAFXyhO/gK1+BeEotrQ8WmEOsv+wudfdXddGAUV+cMgPi44HV6
zU98ZDfUr46O7LSzm9qVOGxQ6RrgVeMmjAiVO4UIGsvZfERKPPaIQd2u0MMm5Hgs++XyQb+Asfll
nqeg08jMl671PM19yLi1drlgWHl1PIGRcShpcIdKqyYx7zbHlnnU0jYUaFGFie8oLGcPrC1yvHfQ
9jrHUkm21xGUzGM9FDO68iilQbfyBs590ROBP0nZOgEI79RJvZsgdlbnJhSewuhhvqzaBs5DqjO+
yJEDSYOEQERJ8ka+tomVmTTM2QdxBwywdjtsMw68q6WVyxNGWBVRoLFy4nAnGhFpBDgrmu70f+fs
aDGMiZjKY8E8s0M2t/lP4L8dwu7kB9xmELj8HvXyQmWd+9Y/Gez1SoU6pX7kliOYHlnCvT9hOr+M
y7rJ0EHrqjE8Y/hwsrUv2T5guvPW8GWv9agVEt7VjZdRIGfozAZmp4JCKJWE+cO3+Q7YsyY2qQRX
57Ro+n3RohBYweFb0ZMLWobWLvDtGIvLb5G7dbgmHGlx60+tj8CShZs2FRJFA+vSo+zTX0c2yJxU
NN/bosS9SYsNaKt3POtLC+8VQMmmD82XfYWk4Y0WDccQQf8s3UHYmppqLiWlb+k1BIxQ1iFwfxn5
50Nd/letIaD8Z3fCdDkzdlH33rUMCddI3vxdokLNt46BguZLYaMumDB3cH+CbT+VOv2KQabdNtZK
Uq3yfT+GYGUl2hDCIy8q9XmmpA+k45lnYFJxzvq7k0pcp5HsxZfYg0WzJUN9ARs7W2fH+hg775I/
pFcJdi3/YHttcAk+DtdGLg8j/MlZmm8HdTUU+9MHfD9T0KH/A/5NNt9MT2m2SBqBzOxeG78Lfjhw
NCDfYeZwsYFZ3xMFheslpmlev62EhqejUtoKeTaihGeFCgKwsnXZseEmTGdORcUCeKJH0isusv06
Pf99YMt9MKtJJwOd00fjchjhIpOVhhTYGnmLpwf77N8e7RCWx74w2Nltg/1iPClwE46VcK/2HfXf
1k4yjypC0PD6oNaoeeDy2byAlYKaJ1ulgPqu3yUlQmqctCnGkjZVa8K/3k5mCjSB8fh5+Ohbe/z+
O2qjlbtgWRl7AQUwyShEfqDSM/zuG8BWokT8cV4bEt8/sf+K+5RGkp1d5UumYs4drmPYTW7qfU28
5sdAr0UWCHyIA2pzLvadm6EE+94TvvlDhTR2UPTb2BFSdG7AirCqpELxYDMlebqBE6YvesGS4yW5
O8Bb0njXHpnNhRLG6IRrJ8my6CcpHmlhskAUHMLkgfvMY7yWgWrJlpBy1naoqG9i0stMFNPdDmMr
jCDeTWSrY1HQLKSlwqnxA4ZovFISKU9qEwqDirkPJt3uIzBHkGKnt5OkBNO83UL34P0Pb45p6PaI
vGoKsKA0f/jFQBtjOG8sNCl4KpzDbeCKp5v9ASwM2PDK0Hx0R4z92ePZ+bcaysrb2fCjZmbnYebb
3ZMldh4mgwdKzsevEi9ZSKRMLjXqgQ66Lus/WSP7HgiYGuEmY0XqpiO3jdZIAA+Mv+YOnVKKtZZ9
icDZKvXOTub5+eazIn4MWDviDNg6OAUGAoO/9IKToVj8JF2LKrM5Js2k2mNg5KPThTes5asISiP4
fduAAqClS8wEak60sOKIj6o8c4/3MqDybDvOMXdaQuGQc78YudCjHECanUao+Lc/BR5sM2Hie00U
TYuGNUw8wsKxW8xzSASJwAkLod+TrkJkocxT0uUiUmYcSO8Bxv2oQpwuWf0YmLsGtyCEERH5eV/y
pfYLQOX2/SQ8/ThCS7nIESRfdTwCKn62iCHIOVsqS+HIjvO0GR8xIOonFPDATuNMIZptzfR0QOUS
xPVJqm/gTdOE5PV2wvVsnax9tWUl9AMeOUqx0Z82DyXgkz9oaMc8Qe5JHzUbfBOwNipnwfFCU8wr
tfCmrZVCQvEOb4ykvX4FYQA4pfeE5xPPwWGbHJqscG17HJTtelLY1mJTwFitX6L/5IKCGrHLTbwo
iaOBZJjq3Za+OhKEX1+r+AEGfuOXsRNWd22B9xMLtcz5v+jUsaN6S5qxFWsh1TCR9EVUcRaUZ36Z
ZyaNsexqHrZ0nPud7v1TP1B7+qXJwiAnP8ejUEhYhQ4cFZD6H1tygFsxxHMIbOHTA9d8rC4Xd2qV
ni86O2IzuW9BqNgqD/IaaZ29HKJ9sklrnFe3WOcymechSopidjm5WByt5FV/W6wemmgPniy+eTa5
6FQ9nMsLHlqw9Ju3U5ahKrddI1KlCvt14vuFG6Qe7MZTo6dtHCe4KPMCtpkAUY9qKWUnVvp9QGxG
fRXKOSxqI+n8yoelQjzxZUWRjhn+pMc1CwB+D+vfd9nMcBbBKm1JfMox9bxMOy8upqFOll4gKzpH
GFcr6lPhDM+CEuy7m8qU3pAmoz8cGD2W+KJDRIX7CPpZI5/5LXNK0cqol4MTiDk5hrhRIXfZniWR
/vF/ZEzy5E+2i1OClQ0vKlNLrwzAiahhe+xCwM4kPGpIn4Foo/HbqEKRKhM7ECDR81Nvg8jX146h
ReTTLEDFAYA7SeHVbvgykwrzFUkJ2gxYtqWltUgvnyOuJXrev7n3ouHbtGWPVzuzqfiYTcf4T5Fv
m7UC3ujTssZetGgXuS1y4+1zQ0C8mdUqBHR8gPt6qy3+9w2lprazZQj34DuRBPq6hbaQ4r9J0RFo
QnaSujR/PQvNc8h7ELrGTgyB8ij0LyBMfcMIKYC61g7dRwSQchz21sA+aFcV0ewIgUzlQ2OC4VC6
Qt9zwL7U4GV9MPkAhijthPPi0vHydKAInCQFm4Y1KsyZp4tZNDzHQp3b/ATH2+LjOCOtnGkz9D19
fQ8CZoFiR3/H0n0t2kuZbDjcXrA8xuxyVXxihjlMBuYW24PDV890az0w46bGN9r+4VISaQDhwHkj
4I6xrZfC275vG+c/8e5PYpIFF5so+xStu2OsbkwWYja7nDz0Gc4jFX11uYCVQsLWHfrhGmrbpOUw
AYTeXXYP8fFFwoBxEYTa7Sj+oMwyrQVRda3MKn69dO7RZl7AUPpTd5v6nlv4Il6ElExYTUDJEOsb
uMAZPy/FColy15B04FupfoXZl7U50txjxKbifkRldP/lgLazgdvKmP3AoxQuAWc2ZBWaxr2UfEap
5qP24/o0IVZoSZpBpmYDfSdiUMHjZdTrF5ExsAmLUNhGS2HXvloOtayfZfu6qmo3JqS/gC78TiWS
NfcvK1FS7w18TQCVwi9Yz0wv5K3FJ6UI8wk3wubE8wfCCVA3i9+ynNPDZlnd1YceS25h2i8w86iz
+aBZqv4VtTmNqbtDOmZDdMFtBD8cx7iUSW9ba5L74kOqpWuierCtU0qjKydh81cMPd+DaV93YzTV
tP1J4ugfdjqTnVrLYYpzUpX+AQHEZglPemcvYyNtg15lxMHT7BuXCFZczMtg2Jd1KCp/Ro5wL+uN
SSp79vQ0IrLguSpa5gTsoLrBOx++oTqr5Q/hNm1jVcwwDIbt8K8pBLYWNNnOuzUDJWj1wp9AHMYN
yPP54LEpDVFPVqtQqQ7n0lbsAIM6uddkd/6msCS7gfJ8OhKvWnEWIaC7BMhq6l8ppx3pVRJ3C9MW
pIpbSf01zRPV7twEkqva1SK7HqWFM1MTetCejX3foAZ9AtfDBCdTuwViepjm+idsBCeaRAiE++NS
F2tlsMjcnRKOBCPPD7uhI85fn1mqdFh2vafa+EgvJSJQnFZUWs1jtIt6DKZiyECvrpeIAefgr53Q
I+6KZZDe//x4aD/ty7NNOPcUMxChdQiEJ3AmF/37lptbIkbmph6z2QK6TqI1wf460vqZlj24lX4B
+piqS/8kyeiXF/kA94v1xLf7JeMS4Vif77JvNQem+lFAi9femwY7CuIP8ltINP8lnK+fCh4XO8F+
ot+zZb1djCo6NjAozUVYyyTmUTnjEpHYL/YLRcZ963YSa4Yh0TdJWZZTLbNh5i8cYRor5MhY3R9u
j8vM0peh2VDm3yXxJ5tPIOC6sqwydUoLAF3i/HYPmgX0SWjgj3A36UOCTG5FiqsGbAK3pUx2/4XX
Zx/IYoYELUHl2VBG02F2z4CbEh81gVfEX1d8aUF/fk+PlE+Q5/L90On1sY+g2EhC4vlNbnWJS+q1
QRbPFEky4dPdEIlQCsOL7Buvfvvg9fE3p589DhcQoWGSesbWNUsv9vMnsqTeO77EWInGjWLsi7cA
EGynbcfxrZx6HSckcMpe9+TH/NKI5bIIhGSCD5NZ9x6SDqRycwx4n5dyFhv0wyWRUhTNqBGflugU
khP3kULWIbIqVb18OJ+IeN1dUJ0kpKtMQ+BTp2DJmGLWZjpNkSKseNnkiQKpN8EixRuzfNn2rVFO
jkqFVjyi6MUOqursEKVgpbEhRWBUoIkVertbr7EAXIkY+q7iBaSsK3V7O1HSKePmAnz8Gqech5H5
0jgrc2L5EQAlofz/mPow0dxScL63skkN8tGlbYDkrxA/zWhOu0dCCWj3xUbVhl8fZ47aLXd2TWYQ
bVPLv/yfPTiOjN5R1hjSPKMMSkBm52Utv8UfYDhzT+EmAZ5Pg9LOFnfsHd5wY9P5lhQ/M8d8D6xV
WvR7dZ7u2pmLaiDjkKT1C1t5pdSyiVLI9b5WUqkRFK2BlXEFk11pvRMQvcrNZUeT8z4DCaAiyZ5G
zq/8o6cOTJLOfPonfU0r097rwIbxsmNdtl28gNPmRpLWSUNHqf51NpuBWFPfo9WxTpbgP80CotX7
ZOFm857XlekQcPuEXXKzpTMWP5ex024jM/2bTVrLYkbeyga3oQ77E+6JFRELGcT+VDO0csj0aSo1
bnuPb/bvVZfjQ4zBRkLq1hhf/b+H2D2qBSFn/ZZLRt8l9LMSV4GlpgVCxRhpt9EYCflbRdB7vQc+
8R0xsiYsHevyrUrlYo6W9QJD3Ssxj+YhxHR5hq0BO5UqEqYwUxH/Snq4OJbxzyZ3fE3yzV9sDvFk
cnY69QVBTbXAh4nCgRPBFu+7AkJbPI0dZnSyRIR2xy8pi7iSXwWlI0SkQF9LlbleAj4+bAj84NaX
Yk4I8kGaup9FSJf3P7NoztAhDVgSiLf559iKlf4ox0mV21Zr/FH/41kPPh3O5Nd/iC5hp1x8+Z1T
6r8UlRhhUFO+NdnO7ANz88buZIXd/KX3EHafSrKKZAp2baJ10WbcwwJCZStXX8ezcSQ2e7NaxUal
usLNwMhdEIuEnONAPoc6sJHVT9jV7Mq/CfPv+YGV8JzHAu1tYy2gUoxwFxBTLFvNBMk4am6ukq1F
B5SE+nDlxr31bx00tUO8muhFSba5Jx/y2CZzMHreO10igT09xWhtWTF3lXi4Mb9iM2OOVH5MNE8t
aOJ82GSOptIBbBCLeD9vfz26HnPUm+jxyOdi7lOcL8070Q70xcd6M4yGSxMnVCT5N4UGxOpDL31M
4YuTOdWivx9bIzOX/QbneJEEb/l+fOR+KunGZV9eB3/Cb2GZkKUQPpSdqudspxHnecRjhlx2JTUZ
SSd2FVGIJ8h3mrNZE0EzUUScxy2k4bCoRcyAClMC/anbO5eeUBn20/vFqg3W2K8nwgS4J/scXZc7
wEoBGgZfwBZUjbv6VfD5J1MUmf5jHucWzseGAs0oAf59RtqzEQF7oKy97I7wNM+10mPnbxz74Asa
mgsaWm+mmiqNVpYopMXQNGtzfXvqgDbYmPTV/bvhLyuMFeFGII/dv2j+mi/1G34RG8jYVfbd0anH
dhiTAFDx3bZ9lvLgYFsLDgJlCdecT+ZpWjWGE9FnbMZY4/QTfRM+8yG26lLs4cRv8tR0OLxREYOV
sFVkR/kyFxj3a1zm/jcC7bC4GIvweHA49c+nczOJoQ+5kLE5CgOA6hDro+8TI/SkDKcRf2kx5lnD
N9QpbtHnPz4WxgDGkPkRZtmoBoJbSQr1nl5V/X+UNgPJ6PuvHaQrp03eKAPpqvBArVDSGNuWNt99
HYLkNKY299ANe+x1Y3SgvRJRH5yhqQSBkilNIhWF/1hntbpgIBRhq9zheWtAIXvRQm9mctp4Iwe1
Z6vMKR3WA0iC9t9dsEgZ8IWpGW13MGu6cCY2OLPMXMiiP0r7feyhZ/BJ4v+QqJ3pr5jKYT5Tn61u
ATsrtgXoUmqVtWmUCwQgQt0l3R0RaFi6HB+ZpCdvzQgeBkb/QfTf+Tsip6IsK6FFnlAmAbgV+XQL
XD+D5AMyy2cLaTita9JVBOuhIZd//mWVxQmv0MIneWy+AQR91Or7orfMcuUg8sBNf7+kRlwSYKzC
k7ijP6GO3ZGiLDc7ayjKROlxXOUy/14F+vjSUSxJeNMOAnDkvFNCd9d2/Ymx2yrLShl0M5h/CbdH
MxdX9+5Kz5hgty8SZs6AFKMbKSrl3Gsb+NG3z94LCOkF1OkHKSfQkgBdH6tUklJd/WvqBl8m+L85
6MKPt3VGMfiuM6QjUJzqNUdUlcXTExluAUIbqzHlsz5YQJT2OUg3SeLuCDbC4dG1imu6BJzR8bRP
AShAMPTsXDZ8RvcT23ToVkFpFNazIo6pU4Di7TCHOsZo6LhbxiJZtJSmkqPNUvVKtJisXJ9aOSCL
f/0q39m36TjHtBe55CZ3FpAZ2XXGqC8MOHRL+oIe4FeewENNOBhim0BQUxPqHJebG9jcrjy7NbE+
AugAXk4sCPDb0ShmoWHBVNxhrH3LK5hBX31tfE/tfjJoy/ea1GjZ04VLv0G9Ug4AAhHXAwcnENz6
i6QBGqfMWr03tBMZ5jSvZO6uCUH5U5nFN0w8eVp9nSqRXZr4ubO9rlb3vLb4ioo+c0wZl6bRNq8O
D85XJ/D/tiG58QAQ1mDzBamq3jZMgJ60klbPlsMxcyu4MTIbHtNRBANkpPEGaAzWy1ronL+HUGt4
aqYVMsmKGjm5A07jp0bolMCQVQGFefBwfUEy6YfC5ObwYR3BIIjfBTeRUZ2Uj30VRtN6UE41Ztzv
7eaqjCG4K0RMgKnkAQZWxObU3QouQLbPMBaDjSguvKFB9WXBbY763vXyfabVYB46MLb/Y3AS0OBO
8cvs3EDLeu27IasRIAKIsU0d1WQRckDhe724cEhKlo2imOK7lHlq2ky+uRxm9/e7QfAMfEHEiDb8
whcG7d/3o8pghsMoUC1yQsCS1RmNbG+UUtbLmQwK03V1FRZsZ/241M71tI2ldXpGbumy9YU0y7ep
C4Bsz/n9oORa7IGec8Ly/zJhgg2i8I597gpVkiqJPNO4so682VkSSKHjQrx+6BsblDv3jKbEi6h9
gy3jS4GKd8b/hVSKL0jmUs2eFQhtJjBZEACJKyKTkvxSDDAteLpn6/1I/jTsnkHwB+S7jTOMX6YW
cgcREregPOSmP8u6H8lUyL+YpBBgd3znlh15m2x4HY1/YuBi4g0TKV8rrg2NZj012qBfWB3ObLuJ
QQmzp/BA+JkUeUTQEMbftc0pieOtf53CeBlroMg4OvxLEkBGhsDk5VaaszaC3mk+Ghz7xx70y75Z
8so6yJUW5ZsaPg972fHx/PUrBDNSc6613J6C6EL4jj0nQU5qOCXcn8sg4AudcLrA4r13GmWyoyBc
tvo+7OCtvqT3hUzyyamGYijt+Agy/MEGoD7hQZ/4uJ3nXe/OJQR7HYT+XmPtWG5AJ1P9Z3wxtaVp
FYuXWizBwKzbllsbRrn0DWm8Xq/mh2DEZyiIP5GSzCIdBuGxNS2X5zw3WluMTwDD1hhknQ2/p61G
H+tiBE8a8RjQJIKBr8GwRqQ4uSWK4dv7pVNVc7bL7jeNpQ1D3j8illflwElGKtSgHSt1VWYzXm+C
JRZL9oFsuKwilcjZZ0bliRlJAyb6clYlZRWToGgal37kraIjO+E1cK9OG3G4uVy5BcE7WaOEOObr
fFA30XIGtQ2lt9u6n/h4Hj8LIFvyUo5SFiIUeQmG8VT3xO8NGVS9iqckxcmXXW0vFrdvVAl0hLqH
QtMGBirJKxxdLad6amWIf4OKfi7N7IDEjyOrHJnONQ6Jx8hFXT+s03zvo1LALXP9l2Gmpy3UcG+0
4ZVQS0DBrgE04sz74bn7LK5pryfQwe/llnTQFbjaOq06ORQOJoC0gA0HI8i5tVJoTgSrAt4MT1ux
LiYGaVlZSYdSe/DGYEDKgd2KePaqhQlC8uIQYmX/8Vhlret72JJJPkAV9Ss2pXILFEa40E73ISpD
w0RMhLAGiRKYsWzUAMs290DTn9A6snQnWTWJuV1gVJbJNx5ATmcMMGFinA+FBIgKQNgW6sPA30NY
e79F23a2DdRT9VhpkafB2YpujGlxw5PrCnNsiyy3n/0hwkDPInoVJ7GK/cXQdg+noVq8ccorclw2
wwWNJPFF8TYGxWOxkZrzJp1qCNxKqo4QeyZaUhJKveMD8PBGC5f/Pu3pKUU4KMBAeUue3CXSj3R9
DtGSdHyKDkfYLk6yOQ4jFQ8IM1eXB3YKqbQlelcvI3PadjSOSePrZ2erGj7Zgeif7JvXvw4pvHWl
iGm7PNS4AH4T6lZa5XW6mifqrqG9k1CFKf2A3xLsLcXxKSFuNSzLQUfcEIHpptWROB7FAi0PHtpR
4mSlmqnNVPCPlE90TuxWbC4tR0SHrV4oP/ueWLwRL0D9x6sCM0Xj+ynQg8aBPvr+SthNm7c2BN2l
5Wd4Gi7DjHFyFNg4s1cSDDjACh2Ar7vpIX5xGtRFNRJgoOAl8/Y5/TWGr4RLW0mB5AHt1q+ad1M/
1aA7QDNqNSfQ4SdStlW+i8795XGBWGvy6osznzgchSMsPFZ6FJWAxiV+b5W4xD2W4Q3it5fo7cgb
3LARyy5FJigYVDzFHNdZdYeCXSZyI2ZLe2pf4m/VaND5VZI2FnbZ7VfEUZbLzyMpnYV1KTGCASO9
rIHsKteXM2sgkl/SfGmwOY9HGQp2o9zN4rlm+oWGDa9MgRb1zilI84a2tHiBKX6e5qQerZlooDCz
Ov6mH81z3St+Hx6/MK1vQVWRfAIeICSvpgvVi8TRdT45cgouMeWExfrmOZMVnCQxUIHt4qr8V9tz
iMSlWCqrevviTLAKFfHVVdIeK4HK3oD8c3G5lVZi99RttcCjDl6tYf2HH4FdrDw27S7nkETkvL7l
WF+Z8mjzp8s0KQH2CjursCIaJJrRWBDy5dWSQLxvQFFNqSvRLXb0hMFCYDI3BpUVMiYOLgSfUg5L
ozr9fXL+nP0Q2X9gEBlKxY/+bcfcpXdWjdC6thMANklK+mJc6eVximzwU7pFd/b7EXFhP9/UmTmT
xshCqyENjDrUs5PyAY04cFCYY61nrdVPjLv5Fp1hHmNJvBOMmPMoxROWcuoE/z9jP8ZPcDEBbrlA
DtRmZk5WOceqIs3NM/J7IeU1boMpphW/VVSHznV5RYfvVT984x9M4fiieK7aWNAU4FznoJKrL6Ct
wZADCnHIC51RdezrUG3Gubcm9+SC7H31/pTcO/lOR4IblvQXU8iyi1WjdJTbSbrI2EJTAuPnzBZ4
RKeh0KZ4eMS3oxOMiV0KbssENc8Ctm5AHajWt6VwTNZnbDm6GeYu0iFvlXe7z4uc1ovNkk78G/rF
zPS1Scm/EW7zDhouYnu5Uhdsj7ReWbif7pWmHt6huNfauWle258QIkgAB4fL9xiPwJ69mhCQ3DK/
6ZB+fO/SQDsS/iGNroXJ0ONaQI/EzZymRZynUqzUNRGseS8iWhH68r7uF9dKFtltI9lA41mKBgM7
ZNw38XiP460U/aDlJm8rF7jhXGfmE2LxlUbgKyk3rxwB+qCoooAljmrEp7Abpu3wzCxwtHS17Tw/
AsnwOQ6CUvDoLCuiiT7uRVtTOjGtVaRGHrhuZXXmeTcJCTS6acqpeBqi1PqBymg0qhJFVPcv+5dT
sqBaFf1ETFAeNg5wzIPtFxZc+UhxrSiC50l/tznGz/paMqyHZ6QeXl/BV7S1KOaqXu5/98E+ASHQ
s7P1tMGxeUn6KIyyC1BOjyM6DDaI1RKfYAdIm0NVGlc6SOur33VCO50g+7Jq2rsaPcSbV66ZAUCC
Pkq1+pMIfNosSJv+Bb4KuWjvh7NvO8ZJQEQTdHjZLtoNxBJlHKPpjm4xcvYu6RIMhmo8FjI6j6hs
hjaSrF0TpN/6vuZyP19CUm9Dhx5YFS5wB1VyOlAadJFjz0y9EjlYZYyEdHbjluSvjXII8RaSVWnz
K/woTjmipnBM9ZRG5r5KxAme1DikJGv3iivpvOifM7D8KK1Hi9Z/I5kit54QCT/OxxoArWKADuNI
xmZoq7QGSx8Mtzpq8LkAJVHIpifNeiKQ0p58LM2hp+JBL0Ts3mJyynJXz5GBdT+dvUL0XZC+nDL8
B32yVfZFpoZyyqT/zWE/t0o45Fd+aSODH23dUxWZ8iLnVY5Ng95y9cugtaO2urDGTwo6gKBBBtfP
VP76S2LF6ELeDaAXfLI3panXBvO0VilrXD3IrajXc4mfCQjYgJ4oWXwA+B5f5fjxAlZZ+8QGuRZ/
k/kNJ/kYA/8EqrMz4xUo28QSJE/uAoUG9sOMJR6wYWbPzzp4x6NhPTARVDqbwzO2w1ETFw5erCMg
Ygpx3OKrh0Wt17AKoK7UcZFhg9RlXzO/GDvttvrtjagNKoKTbTV9dkGVcrWMdmckXWHWbvpMCwwf
dcGKCoREUswg2zV16GaAuT8OjHWf74S1Qs/XuGFxT3JkL2Za6vhnl5j24dUGAExU9Jvah1U1rUFG
aFY4dOSja23B4LpbNw6F6udxRpkJEu0EY6pel9ZlVBWU/WIUyL3Cp51IL6utj0LMhoURXziG3EHl
cKog3PfM8p5VW77cwfb1jMKmsPxw61tL6UTdLVJCXM1uWDWyRx6rdE/CREwdEojTbSc3Onugx1vZ
Zw4ZBEt3i8+tVfurHv2aRChpWNHxXOrU+uAd2ZEwVE6Ez0D++gflC/mR+31JyZa8A4w4mtDz/O3o
HqCecfJ170uAQTMMHQN3IUFLlpY13H1wYQsPZFc41eNkvWbsaDlSlAHOx3QnxOVA7xa1oeK/Mc77
HYJK2zfInFoFoMejaiywev22zCI2av7/S4QpeWanic6uBPcOG5WO7R1JgWIAifG97FwfzDHTw3GS
nzykP2VWc3svllea0Ry4zMcIHIxqFzl7bU2I5CH5ih+9i0oI3IvkBoRfc5MS+wdNiUYfNnAPDEKp
nfAY5aQFY3SJprPpXkGBQMw0fpE7dyKclCdXEbI2xVPkDkzMJfEFYP79Ezt6Sibgnp77esdLG9v+
vPWsXfQ1NhH8m2l3QAgI1otqa7BBnkC79nLsjVfRf2JFe94BVR+b+DiP3nUFs9NoCYgQ/aI1yMPE
yx8mVhgTO4PvgQ/dkftdaiwAKvSYi7/kemy661vqHijQUeugVnkyUSVFG+aQndN5PlaPS2TTDHQS
bYXzpKA9yXi23MgZze8P4/cRCYYBd46/AfjZeQElv9BHkpfG49hEW2ojQtYe45OojsPlNBrMM/NL
ozdsqoBY+LvI1X8lSoRM2v17zaiDB+xiriDu1FAHXE/Ht5XSqPOvYCHd89APppEKdIRupxx/35ym
speF+9tlUhWUXGYGvV28YDeAilhuEFw/tytgLXVcjHnuI2ZJwvtxchnm9QZ21DPuJpvBIZHQg2Pk
Q7kxLxxApzqBsx0qMkpZta+dUz/uS9p1jIm+FzFCbsGMSSikx7oxYwOweuXsbLzTTWIp94hMEAtb
Rex+yWTGlieg+9isQFYvYAcPNuz8m3qL6uNGQT/OpH81v/7kgb2wJ5TtoBO9EiBiwy8xVO8VLgKA
95iY5DyCWQEY6umiGev2r/fAh+OucxKYQVBGqbcbr4q3Z4XEQhPbgbpSnNKZRinPfuqdsetK74hR
nGokXU5tAxav+JdkEV6ryvcf7MjtKinj1lk72UJjM1ugf0k1gotfXS7haouZ8bKk637CPgxJbInZ
nY5e9B6IMEqj2esUQ9DrBnCvOBQSD71k/WcyclD1DXZerYO22O34hJ+WAuAS8L2ODEq7W676yHy1
v6lAi5X4xOC7u3rELPtBrSHDfhK1ys/8ZIexHd5OjlSU71Xvsf2VXk39H+sJHVRRO1sZiM/tEpcm
jK5NaRggdJC5iWXbZFCDHZdzfM8oxVuBzNpkaS6q4Nxb1G/cgICgK5PsRuDeCtI71GkLgJIFXOkL
1kyCw7H9rh7arSnrOD3juSr85NghQbtziHZNINBLGmsLzcVjyo6DCWk776nv5njQ/eda1k+6lar9
35OEUn7SzU6pdFhL9dIoxH5PeKObSdc0nuZgKQHBG/d2GJ5xuui1SINtbo2CDPeGJ2Kh7drYQ8Mc
/sFf2vf5ekA8VnZTbd59ys6fTHq4Z4U81XaIif3yC9Blis2PiS/jf7kNN6laEeQ0Mqy4qyt19yN2
SYW0CBRFMR/oOOy6TTxIco0zjaTdWOLDRxWXu0WZuE2nprAdrwKVlylhdvpaZb6tz+GypoyWGVLN
H9rkw5YedvfkiStw46E4Q6BkWf9ljvVx+nilK7iMS6q65/iRGrYsUVy+8ixC3cx5mlTO7bZTw0QK
QgaNXtIxkhODmZcnts9G2cRgik8PObM8zfIETRqsrxlekkLrDwDTDlLvGtPB67dYrzMdkYVomdlH
V0Sy0vB3iD57bsDlWxV0NTtSmlN+jKXzDbh2Y7RKRNCDUCk0BOSI+CzM8+lYM+zR2cgbXnlWw5Eg
CYkLcsWlSi4cfe2UT0dpqkE69ifIx1nOEv2ZXnKBz9dvFDgsaGY7Ubtv9XnXBDwaGiEZpjtHfXxI
KSG8jcPnwgTRKD77zyct/7rD2TCQMEnKPqmZ6FOlNG0PsRkQG1FTAUCxmRvfyF52xX1xiP1VE/iV
FA4GNRU71HUjbVNcuqIXylYB1LZE44oJ3G2nkX7eySIcE9qIAuVMh6SrMzcGjalZTZd1KYvbwAzL
e6mWg89G3eD1XnDxwe2WV7Bt3mBTtRpawxQu+E0QVGWmcfZL8bh2N9jbgYI7SroznfWkqSMTP6TX
Ce1BuKSptJhu1etRO1+/W1IqZ73GiYW/TpcyM3yi2k2ZY+X2MUyUv0UAkIEPZj+93AzfC+DGsH1e
DaNVd87d52x0qQsiZTFwNFervZ9EDHk8X8UauUDUkN3Ly/wvhi4ONEm9esSoAe72h0u31d3gVR78
OFyd824GQIxkH+y4REC4KlTJ63jjB6u25bUmiZppYl3vGPnvkKxo+2pRjZf1tIwtIwPeZYZAk/eG
43OJkFmk4jzQbsGeuKkM4qVzltayrZA50iJ/HVul26ZaBTKgxkDaIuMsXZcHAXIsa90u4kMnUMA4
eUfneEXdSAS+YcQXlO8oVER/2C8wKWRyhXotvzeIrsHZTTHe3OI7MclJj6MZQQQiBb8kuxugKSzG
CA18BCaOBPIWDttazEGVYUZKjljxhEN1ofEpnnQK9dQt0dWPysgqYgG5AFGYrc6PqPorFpKULJQE
BY1oeJJqXUWc9+m17GyMtu7NvyVVnIyv096eyARK/otABd27P71bWrHozqRw6IT7F8M4wLFOxMV8
z6jUWrWhL49ZIpr7BTcIJPXmEOhk7cSBpVo5vkI3dz+4ufvLv/nf4icC2NMH/V7Lnkb1SMLLckPx
69T6wxGWeC3nx77NkiSj0y1fjarPQb4lMsuv2zfOHLECQHC5r2LN99LwBbX29eLAZMJSiBGg3gEW
UH44fqPUCkoStCkQyZL2X2JUHwmrCNUYEI08RW0piMFEyTpeqjT3s7wWBtusSfmwWCVOXrgMbYGF
niVvCqLJJf7IkZX9uUt48SLyVNFVqHN5S5E9VwZOQN0CRympWA+sHvsnM9L4AO8bSBTYVSbQDQsG
ZdAIEgVf1qw0s3UGyXdQrdQUW2CN87LgnZZdrA2THxwZjtszGvCqmoa3unPEQUO7nXSsHKUoll4S
/YqxDEYzSGDqLFMQoJhO+P2cz+MbmHpnzkplibrNSp5rtSWhqWO9aDaQnzxsvNBqUk+Hfqz7VIiG
d+FIWvaHE0GHw3b5Vs7U3n8RNC+BBO/47NprF9PE/T/tWZ+XhIuzZ3Iu6JQT/WjSq0GJvI5XbLP0
mflGQZtP76Poj9U+WY1L8WVpcKfUiz28nH6ORTbDslVVhZuLzKe7CbiIJgZRF4F4WH7XY2ta6jGw
b4aCLOBjLoMsaA7d9Ye1x2Oue0P5t1w5uDfy2ss4Gh++VHyar+E5QTfi/aqaqyqRK+JFXchIFFhG
wGlQeAjUbJhZ32F2WEKpjHY8AYhPdeEi7cp6BkKo3vVcGXe03JhYSNTgDQBnUwWlbgxUBW9RVYfv
5UFuRc4iiOQEG56X+hx8goOzb5w6Yj/enicJ0CocsavMFEWRS7ly3mMpISLO83d6KuddYqIidLyO
BakXtSl5PTJOW8MKPwr/VJGYfJSz0jk0KX6eACzIl2LRzFajxgNFXOxl1zpHE8IT80QXhQLwT3P2
8RiBRgxapsRvijKq3GQYg3cWrOXc8QpDgcCl04ojupylOCtNRQD9xq4v+9qKLpJUzgJnx3KcgcED
DOWYXdl2bPTn2xyylkwXMP8dhw3cXho0jjhpaFKZI1Aw9dZTdsnB8gyXktSYPcKpHDT/NOlX78Za
4q7o8v7x3ekpeguB5aqX2J7xCsjwcuelwEGrak20SWb1DO96aWsK6ZVE47mTNZxmZc9gdt6K7fA+
xUn8eVG8OFksbqknAfrt67jRz3I8KO7hnA7axoRQ4dp9sG8oeDBaeJkfPKGYeba9PholwokfdziA
MxbOwF8o0KA2+aRoJIAcH8wRc3BfXEAltWBv9V9KXCKxamdpp45GHeS6vrCHmMx/6yHAGnhERsv4
uIP8INPiedZpM+DJiRHvjFUnn6fIoGsH7CF+gKszxY3sfY9zSmm2CQW3x9r2LFwnddLuK8qjmOWb
mwOOkS//BM8lC5r7OAsFWNojIzDZ8hIgblplwLipOBLdRmXWtiu/f2d1skH5BDYyxoBCKMNj8Veb
ZDVyrB3mcr34K3nFn7HKs8lrrPPv/qx4HeJRCEfaUPZJdoGNeuI9m8MgHt25KUN+IgzhLfN8LBif
YeuoW3sP9NjImWblxzt8H+OG5Q7nSsCpKnTexkW/8jdsli2UsCdgJ9C14FxzbOIwFxb2QtVOBQ7s
DHsLP0x1V5pmBPBBmjDJ7RXZTO/qxcWJXjUG9yg8ZZnBpyzj+mfSlVcHRNPXF/KAh9nPsrjAa+fU
jfC3E1SEngaTdgV20Gb8m4UjScwypUwzewE9tinY+wjzv/YCd0KGGuDESp5wiy4ohRkxzcbCnfx1
g3MRuLIUaJPk6nYn3fjP6B0aieqzOCd9yjwcVDXyY44M49AJ8LJETXkq0CzTCG30wMAAb/ObkrBr
iifrn54JYHN0BobCLeWNzwd+dnJAdO7alC2Moe5spIco45UbQ3acXGn+YEyKj+4htg/XnPN3OVlK
4vKP2ucXcRww2eNCcBq206kcyZsuEfk4Z1MJLB+X7gh0CSy9WqTtD4UIfKJNWY6cCcNwrFwD+tAI
iZ3kTGimxa0lfxbSO2ESVsndFJRajwynsyaR7IlEh7VepKwdxSFViX/NFDRpPFlSi4JuRbDbz4UX
UfH4nRLANnsIUOpQ1Qa27GVrQycde6LCJ2rwFBP95XVFttyNBy0B05kmV0JAgjqsNkmez6w95Ilc
Lx15nrVbM4JjvNp0QQm1F96EHJcaRvn9uwClqcLhxbZLOH6Q+FR2FIhw9/AYLHp2pSx0B4TTbGo7
RPr8zf2vtfX0EusyFryRPXvlWpZP2MOUihgEqLUL/bA3ogMIJpUUviWWklIuSmpSPT0tNtOYRXsW
a1qH3aNgQ6QwKujKZ3eft0hwDrpKxkobSzConNGtcA9F/OvBN0+s14/cdThy8gekymP5pZnPGeY+
Zrp2gXEQsWw2qbWkF5AB+ZAVJQuDQi7ypXKQB3T4VHLa0S4TYutr8TA/Y/ViztbboiIAHxF3DpU+
E6bz61GZtZKJ2zTMegZ+ZjYDXzO3mGzuH8wLWrb3+0KZnb2abCat1B4CrtFxEh721Zzv+w3jL1pe
1SqsmgXD+ypoyeNqaD9fwyxa+EBubR0gRC2Vw84xLGjfcAVAL6oUK1fFl8yPDXAm5HsNOFfj5gyP
cH72H86+dv9M/KNmjD0LK4WSzz2vg6Y5gQGYa0D8ItUYZcLrnfbXmyMTwFuyvHQdwbzhVfW1FT1W
DHcmU1Zyc1E9QekcHY4ai4IPDSAPQYiRq5FZzxuPcQN4NY0gqg7IA+etNey/Cvj2rZoNnIRXiRXu
0himIny0LQiDZ/UtLcqNTQkdxwKD/CTCz5yzE6oo1RaN+yrsAPorKmcZgyuRLspj9oNEv3jz3X/x
s04+VOGY97IKQo/71xgw7CscJXHB+QSGpfD68CWDdw4/eYCz5Z3+cuXVIs+JAKigstNWDSU4vcL3
sj8ECHAD7CaIF5AXN6IBVKPLGZWE/BZtOB/cu98uCbwx9xh3rK7rLOCadNuEVd3G//vmzm6riGLz
2VtSqip9Lj9JERpXPh9csim9Dq7+Q1moDEIcQ8+uXu5gOCzc5xIpxBMnvCUBW6WPjC7Y4Sxj/y0h
j3rRKdZRAwfKvPhxySotK90EWik780NUkwFIwJ/ldwJl3ZcLQ3X1RHlhSz9pZk2cUC0WBmnDIc0V
jBdhRu6KycNmKi30MHzzpxUTBAPEGvwql0MEhVq/nrDmYk2LtUzbuKOk7S3M+WUdvok4M6qtw2xD
lVWYy7dO+wHtl8Dg1yqYz/cMEPYSBMA5x9DgQC+Y/ZdDGykSsNpDtRqlOaoKuxvUtkWZhi5ZoRxU
gUkdnS2+AoLnrPJh2l1FqpK/+mVF8Cf6YhqDkb48bdPuqwc2xFAFPt1nvikNfrLgfLDSsWOBe695
8QNz9rSuYX9s/AngfYEPwhWe0uriXxrc5o/7auOWE1PxAcBPheV7vHXT2c3ZTU32FVJxY2/1SErG
7dIYmB4ey1EVRC81sSBzjVvWtG4EadUJiZ+VCSlYkT9B5vRx8C/7HwTrUen87/moXO+U4oDQG2Aa
ubgrQZhwUI1FGwBl9sU3fhqIvO/dol5S49yaVtgHCFhHMKdeuyyBHVvcqqSjsPa2bG0maxjQ55gO
h2WI2lwsN+gOXLT3XNyE+wTQzEI5TlbEcAWOwiMLgWhGbWy3NHNFgr09Ox2MUD9s407+frJi6zz6
F0DMNrpFdjcASinY4VLHkgGjGGCun5cBVikYEoyCI3hds2IP8muLOzfL5Bjqkae9uF7KIpNgClAO
+K9G2+IWeBFCdA+RRlq96PbFZtptCBY/wAsOAAHYSVOk5QHrR0b4K4DhJxhVkHpODit6qBMniYNw
TsYcrn965r5xHY73ysofDx/KVslYljab5hHh/MdDJ/MAnhaIeBjMufv3fKtuGyvsm6PONEZEX9t2
iRnzthdyGYtmt6pzg+gtHjTjbEmsa7bvFT6Y045v6xjPuizcR5zJyZK+78GaUlCMSPEUUf1jdQ3B
Ou9Piqyi2/SEQbmALeM6Q8hnTrlwUpYkn3SdoYOw8PEEeWAhSzYcisyeSD5iFpf4fcBYCu60Tk5W
iK+lEN7LHk9u9oYW9ny97KN9InqCd37F14FYnztVp7dgH4sxWNXZ03+7+fr6rtEqvDBzvmm0l/73
tT+CzVZUsH3csy6WmEEpTIVwZC0e9aw7+56breXibn4yJQEAyhlc7OsMiZIAp7OmyFO5CqRlFI+P
IFaeNRih6H2APeew3MW/txgPfMDS+YJcX2rB/l2cdnZfEEuKJirUO04moTwzYx2/GFdV/PwzKV5X
YYuSM683W3p0nldrX/wEQa8lFWiarz2QFOUJFeFJTCVq9gua5wZ1CaHGjc+jcaMQYirxJrLeiCj7
z/aDEjuxv8gQfYKz34okpn4BLhFiBBrPBurEErXwnaJ698jqpVtEDfCwaeZ2pJULxsBYFcaNHd/e
7STwPjZDqE51SQn6jQSO9+Vf1rApbBXwWpZC99iK7OAOSQTpGgqCEs3JF3KnhAoEc/nuKv6HQmRl
Bx/z0z55ruNlq5nOD++4hL/rdetGlXzYblZr1aCLeDjPVeHQNDeqY0ZXLX7XqSaL2DY0iyZU/oAL
AnrEAvthIHITXabHyoqqgXfXVTyy7FsomoA8fa6zLcqvHEkc6w7npuW75MnJyx+bH2q8F2BUQ2m+
ypDGEzN0z6eH7HYhTp/WrtJZiTlV9xAr7B2PdZHmINn4ZqzuuIC6c/q4HoJ/4ilOb+yld0FLW2+8
AfQwWrwX4FiNGPj4fHksjEuZdbTSSXRxRLQEuutmnh9SqJM8rANAE9nJ4Np05Qv7JrEORcEJdye9
+gQ4m+xAxhnyagJ2jq6zjrxB5oWW1JqPKV/XYIWnYOjNXG3ho8axwJUe+CJ9p9ckaQE1abdFJQpE
aM6wZtfYDbzzZCa9fPGRJzR78kpPIXMOPcBwYzmqtZSe9jiyXWmJ7ma0lB/FnbDBd/AbpWhewsd6
0jRPqJBn4YuuN72z/sq2ZNDkZguqNCZbZOWhZLsF+goWk6rwJcWlaJOZ7E3631vklTmK0fALP1AL
DTtaF4ianpSVA72QaMnMzvZwQnTCTFExdko0ujN+6FYKyG6YBN76Fm0RXr1V4aAbu/NnJU4qbGn8
OxiH86zzbWLD6YtYHrhmjFTvr4TWGIoL+e290zAS1/qtAVUVpBSlOfwkMazIvhqaSFuG85yIBOi9
vLGEK/gejGkHwKv19cnH3nY4xv6PdTYnQtE7K0GJITgbeHAShN0a2Q6ICxUKyg13XZaNZKv2i1yV
ooQszSNPXyNRxmDcsWh7HYjidG4Vaey0poL0d9f1TbC6XOtjLTlW72xa7/5eqTaJEtfXbLDx+u4h
Iw6m3Mt9B5Q3KYlqbAjNtOJUz8SxwA1aCmhvdbig1b1x2ytlXUQmQbL9fv4XGtvac9JJXga//Ac3
uT+v6elunfFnDzZczvwSx8xajFDZZCCgAqFI6TcEJFS9PQm4oRseEsLYUleFZkFqTlupmG4VsdCK
mySAMNCkk8kTN6QGf9Z74SlmIR0d5w8KFe4hg2YdyDkcAesSV8n8SZLeZ3aufawKJcBlRRJjf5sv
k2UD6Nv2qYf6nkbPEHvRh/JOJ+RMgKJeICX/netRCaAA66bLQ7rLctNbVz+Iao7Z8lWDcehbYDSX
4QndF0FanxlIn/xxiFDqw0FWab3HVUQOdxWgngg8KbjaYGpGzLnWQq5CGgOoPdlsoPC/iMoLnG5b
0yoOxlRFRZRgFC1sjj1DDmukHjcoRIGAC1DopUIDpOu7gYbN2jKkedORCF3KaAmjq4zw/qG+bZwh
fQ5/dORBqD3DThz/xAj3/J42vb5T6eWXtZG7U8fdj7csWV8+/VtdvTU0tsN+ETEd2Xj22bSx6nWV
sUuqQ7/ns3n5jfRopzUBiZ6w7AqF4XySbPx2MVsDvWexM8IExlRJTCvcm5erzOEASe3jis2EsGRY
ZUkO4IyBQElpaP9IwKJOqFUyXHxjmYJZzByXZy6eA+GrlrfNeVcejgekE/HT+QzEbKGrYoigbGbE
nLtgw4lkwjENEA2vL6lavdMu2oHkpzn3tsB6Vlm25OjauYpDnZ4NlvhfRam/Emo9Jvob4zH/omNf
7Qdf8d2wijssebIA7ypiszMS01rP909IUjSyMwPYZrnXq9R0Y04BRMdBjVXTmc4+LN5jam0vonVf
5ERaI968brP6woChAvJhTxCChOggRApKOfEc6EGGjPkX+OW+Xbf8KRxHOzZkeE+Xxucki3JQipvn
4mLGKaX9ICaNhpjQN+xBNKYrNGVsFwBdseHg2Dj9OGF+X1gNYJ6YIdBy5kPmdOSw76s1j8eGum7N
1ZqpyBBjOdkHacGPCX0Ll/CHZvWe99YIgEsRymmvNUgWAhnVCkn3HykIjFJswD/nQrnTarCxek+E
v2zp85jt5M+jfLrTelPlVv1FTC8Qxs8SIcSoknbSPOL9Emm6Ce38fJi6dMc2RYtR3zRlfTvdvuDy
NXQ7v08GTHxoR/quqO/PQPPP1RznUPpGyHpkggerAk/cKZWzoYrbq6MNnknL0sLAEl3mr+vqt18d
R71dLhTaCdNrdpyvjGvAcBNqM884JKPVTeIhyjBfcX408lV+pJzgQCe41Ez4+PbI6yHlvnGIdyHA
+0iv6VCHaYRUJ6SjfbEqCNhvJd+UgHsVQ2hGvcLDxwVBHvSnMAdOmDiCztNRtDfYaRffzAe0Z8M+
VfZ0FbXql5nj6wop64OTYsio/peqoTA2CPLUv0RURcmpco1ACEGKsKfZEbpK6RMqwHXESAdDUwNi
92wmgKHmjffNaXWkEXRIzhriQ+rcPWNeNI4FH58DalWHKjiVWw7mwPzFZ/uJkjVvzeZOGSLdw5i/
HA3yFxiz0Fa23ZNr2d1ZDT4wjhceF/BBS3SbHNUuiWD9fXdwe8Q5BFWnAn1eMng5YE7IQ27fU8Y9
J/ZEx9IXdTCTDkMbjIgVu4TvUwQc+V316TBpGow6hVqBgyFhmLRwtPLq0q75wV/W1MtZ4GKQAFCj
6efCLjVZj448OFbN4LEvOVy3WtaVSlbYRMiozrC80D3oMr8falBFKcMXM0+Z1FnvKkeFU9TIpGUz
q84UB87O6CjMh8GVunkevm9dfCF93v2Xa8KfQZzcWFU2hb7+yCeQgvxShuFV/ozR+CqLyamc4b+Z
u2F81jsPY2GZ+PEeIeQkezxEVcesx3f4L11e+YB32desXHCRBCVKXctoQLZKuk52B+QwG0jotx2B
5a5+C6r1wvdXLOFgXqfD2F+yNSgNmnCHbfvz2Ep7OgEJJNJd8xCvpjhxKXspVSTRtD1XS4txsgiW
2mTPoDMqeQ98U/owMn83Vgrd2nZx9dwgQCLeFTk7XN/D8zvtMMM22A8oWbdkHUbeyZ5oZg01CUl+
q8XCO26gxF7RJDF60u/MMCQRy7rh5RJlN3AV7JsuN/qYF61zp4PLM5H7VOUMPvdakr7RmTIysv+T
IdI+dvNvbJjwgHza/rqzl6eOHUCEg2dVLMmu6zqyKUmHifHmLJT22pKd1OzbdMU1whJEr8TCqMPs
AH15VI3Rav+ZlXfrlmbeeCA0YZPtLUMcv1ISZZ2HFgXvWpb3nA1ZWlpr3fWNI0PUrIox8lI7jpma
yOaLdkm4ydRUfngTdjvUO6u2m+0D5PJddnHw1owCOKMXp5CMQ89O8djcexEXwm/qrI8aqRuPaSe9
4/6ax0uykQpQiBuQtsWzkKJMH54E/Nf8zr/FCoo0MxKVCcDhqJ9dnEu45B9b5ZwqSANeVp+3kUgc
fVTb9B6NqOZE1FEQPmxT1NO3cjIaJDfXPp96v/GCYLfnSXksWWpDI/9h8Qn+xB4DdRde9w6wxlVa
PwPiKMZIRAkXh/PsdoOPnTgN2JgSpPs3nA64P31KEKlm76NrWX5t156HO70ZZg/xim24VGqAs49I
UHGIMoYIe0PFeQoM6X9QmnWFDpcM7RX0IjE4t7ZB+cAtF81LROmApYm3JlyKkjrf6Ijx+0hfcEjz
hCzaZDbgbiCHrrGsstOpvH8bGX+EVJiQumqCmZsQnS7LRR3mK+2NRLQ6ubkyfo076C/WfrT4581Y
3SS0z0lMUocboexFG4wVOXEDUGNBBLgULUl7rvpirL9EtE4EuHsy4AEF/uh7NExMmLphmAYQ5dqn
16nftmwEKPre7vJI0tC9RGI5AUHmThHcOwk5le48xRB434lB1Ia7G47N9sfpRgrg0EPo6xKgYvnn
/lZmoZjVU+VO8d8owLBV5OntUISu8eIwl2a4CqRRcz8n36q19/xUVks1McO4d2iBU1RTwaNfUfFg
bfevWSYjQDcnknsX3VA2m7HBNqjPQnM6eRhakYg0+RHI5ZbR+4T9XYp/TXZJspnaqot0sa5ADwy3
7+snSz7CAeFeYWqQOncCZJF3xX23AM6YSG42+nBkajug5iwGzU83pBW/SRwm1evmqf0DU75r0DrQ
qRBOaGQ5kswkMflrkeavkqnk9MPWBVY7AYOTj8ekAGo4NxruZzln1jY0HS1+69oLDJos6EmLPz4R
7OEbwEORJtCaLFFCweI9mw9cU4/4jkbg7DZgvFc8QenWjiN4WH6tE9ctexkywRH0oBHHIHGrnKKR
RkCCz25q5fvkc5g8zkW8IUpNr4VI/0QPbtbzsFdW+gWj0Ar9DLMAE+aDPk3LAe/9+yeJw14rlWm0
O+APp87L+kyP4wPQtMO6BORk89VDoNO/xsUGptKznCfbHgGsSZsI17SpLg7X8YU0rq7M9ha5lVzv
Ye/mrGDSwrA3zHHu6A9etmqGm9vKpR7fr5Gbs4bHIVKX5+LwhmEERtHuyNL0eLVnLEY32VQyw9zL
piPZ1TgTFtplqVe72f84nAooaDDlPVMVywgzMvyzGnm0cfHwKbKemFrg2m3QTAXdqOA1UzXhcF+u
iPv5FP5YifbT9lDbWRUMdKM4QBjYN4kd/bY+mAs0Srs64uIlWe8sNnI9oIpNLlgw/ucn3U74gIJA
U1SfyWkNy02GRMLmutQtHVazryxD1Wga0jwywmMJypa7e2cw3Vog9y2/6kyKbjU8TlBMvGNFZoeE
UuB3LXN4O1XQtG0GMKoOtTqxFcAh2h+/MiVkXj4+iEChDk24hNTIRRKOPWM4i8R9z/yq3swVxrOL
28oKKIh4z/kAdiP0R6X7i/yET+CmyDIVrnRR/26JYWXef0EJbWBO2Hs5wGgETKTyZSnAoeTIeStr
kFxY13ISbgRU4NqGJbEi2VQQg9tP2sJPLqdkIrkv2nmLoMYV44zTDs2r7S/DykqyOfTh0IV+yTOY
56P0wjrM4i60ZYhmAszhJfG08iNZxplAyNejQ+rkEiVoM6O1tJFJ7fSaJelfLUBL3HWnmYR3EKGs
fYL8b2QgVAnysYDQ0tCm0z7J+qTDT5vwqeZkecI79eviOlE9ynD9xWFk19qaMPNqY5A/TC3NwkY5
1ulnXHhNeSO4ecVyja+/G9Ud0F1iYunjOC2vCFVDHnZEWURrWUQj5TvpBDdHpqBBiVYGqO5m1oM8
/DoyG1eDKmI0C5VRSR3zxE4Vktqmw+rq+CV3WIaaOf7H+q+NEhn03kUMKNvhewStjXtdOGIcZFoT
qVADmeDPLB6KEM6acGmyhEm/StwI9trUbgeMFswM+mi267naupincYE6ur56Yokl3BTA2uLMu+6b
L9ExwOF+YNYhWoOKF0SKnnLjuvHWZGssafMeXpcrF2/XB0/hT0kHXygdg4i3fKwk+6bBZiG5aPER
ZPj7k+Rrehv155cEcYV3xwOMhhNi1m+hL71kgxV3lk3SkHFcM10gjqXIQMmMHH3oIMnGltcSlt0R
Y5IstrdDZGGCBpGKrAjWBOEqAKosW0GM0UFjacZvGsrAQDdGiWdbp3z/abmi6zwYE/eE4ZgLvPQn
cx0oj7bpu8ziIacv6t/H5I+egrL9Op9zH04tzaDT8FqPxVRxm8LJuO6VMVXgxJ2kcPGL/Pi82tOX
9y9mXCThy0gk14WiDeJNhGzKxuf5m9LV1Ox3V9knG1BIbPAJKhS6v0N6X+yA6FC2lTvxAyp5cfLH
Vq5psHsVdLvLicuX/1hXheOiwDI59BO7qi8SiBVEYBmGCiHifGmPVcNtCrUjAXLnmNkMvXspQ1nL
kzYedRkmAtRRvqr0+8d9KGIp42Mf0Fyr30ixYxDLs10njoEmrNYiIKuPEpUdV09rCfVan1w/MUjP
Gw9GAcWlPbhZy5kGz0WNkIKZaPW3rbfF4+kpJc+ieXQ5a5gOZBPpc2fMlwE9v+tnR85RdgGywTbf
czcuI9fBCScAt0AD6l4hCKlowS27OTU6YvbtoxvqN5dnM/CwITnm7aG9UO+6cTo5KYjvLKslbrT7
/hWowC1DVVoMmcpDnG/v+z9vQbQ3HfTPSWm2q0w7MYS81HDjr3vcUr4kCNWPp9ejoj3NVKFl0oMm
V5lxn1nVtbpdv4CLnM19k08E8yjrilz1wp18LHyM253/ydxHHxnbNOMJDmeVardKbVwKAEVpBzvb
s7K9wu6WPXLKvFBKkA4JguGItiNo1SzxeqReczFnxUXq7MNT6H79hBLiSJBNeD5UZTk90GPZLNFk
ukm5vfVLtW/9y0uvS8APpGEdE1nls9sB0uUVXZ8PSbQ7GAfjfvNkdvRGqczAFjvaORjDJSRnMspQ
7Cm8C9LcUXZpG2jt6DDFaJekJzajet81pO2GTxU9cUEd/GlOoEzP2xbV6yE2jSZ9wzhiJGbgI9g8
/BZzfXOujoropEJoRlsWE5i527jqBIBuzNi7/qQjJV+/s3IM5C1LrLYCtypUJrmHQ3UUfkaI1bvX
ONBMbsJMgeFEPG6JJ4KzLTP1i9uIye/BfJgSBH100UEsv2g4Vge9MHMQ1eexBf8Tuspl9lrFyh5C
eeszWM0QamHwsAOx+FMo/4J6irtCmvHK5lV7d6dn+J/OIq/eh7TgWlA21tOEYQvMyhpjoeTXvT31
+62BtWUnoHFTbOR40f3xX4LsTz6sxbMRCFYeeCcb9hal/CxGcMgO4RQxiyMpjSVd7AvtsP+N3OWv
EpkKjYqYTFOdsFBSAf9LSxWR4fkdGiHvuKPqS6dV801SISfkmZt/3xyYZVVC+oAauSIPmJm7pF20
IQgRuHYQQ441dP/hUP8/djYnKeaDVmcS3XYmo8KqCormj0K3vy4iflyml4TXo1zU/HGR12LCevtR
1Y4Xco+ohYgprby3arcdOUVsukD83fzznLv97JRBM5DvijkvmxH1gK6+u/1eAbyCKOGdI4doWFu8
GwZAF+dE02ChyK3aL71alKYfCvI8fB4B/AVdOSBIMfGKJ/AZ5LkloGFugrcBD+zQmM7yRrkF6Xq/
oGuXy1SwCNMZtyPwzvh7FNLN0asRClobQ1Oi/wDmwdd/B0Yxos7/8B/+W4VV0QXplN3MhWHSAdeL
TRNOQy81oktxOYtmwuW2v/pc23nuWnuxQrK1mZRkL7ocQrSN7jsgYN58AUdCY/TIS3L9RXrT2hh0
DyrddBenQ7/y1XbnU9e8rKSyEd+nfkKMYhORcBeh5CdhzsJFQZXZAtGSE84Gw+iXtDBZuCiQtn4b
6YQ5duA3+fXc8E6D+U+zrqucHPgssy1ijamfdAr4eKFPT+UGKLVULnITVDb60smyc8i5zA8/9wMC
vYAxLBWjAgcaLuD5Usm4sYYy1+NGkHovzl006mZirEiZ3X+5GyJOI2YEGE00f5Lw+dvKdfLf8GVn
vgOpa6JuENB5vIsXLYuVp+fgY8WbQM8vbgz88IPExWL6s0XEJgUs9Ii/TKLQPHVJ+IhpfBagNLYs
ddiN+s7OQ8pPAOLQNWVHcKot41IkriXrZufEpNGy3usvJwRc8FlnwVVZQlLLXdcxQJsOIZA3Z3+t
X7OYQDO7WDAtyY2JC1oyICgCzTZkCNyw2kNDKGODjgnzcUo2Uu0/dXGG7o2cVgVuriw5yhXfLNNX
i+eygiPxHzioYo65osAJwsffirBoaYYDSjh8vuKK96agKKD8edMe/IIHF2PWR9r7qnG5HGiddbtw
eCzrGHYduHoW60wl4FxUx4o0RdP6M6IlpfPRtyVn5i/BVCg9/pzEXvTdt7e/fl7puObTDUymU2EB
Hn2YgWOFKT/vGFK9FGIHx9U1HEgdoZOMC9xjImNFDLSnYSBR4kbrywb0+bbkkPFfyfmSiX9XEMZ8
R57l8On3y9X1Amnta025ABBTXH6du8Zh5o7kwyrs+7cbhYRvQxbpU1VjTyX9aZiEEqAr+hIKVXeV
9a88ll8Pms0s+pmwzH0k9TLmDE6fDBJM3OeJD4cOAOeUHRtx6uUzfp7CAvD9s1UnhM9tJuYTZltG
JsRQgDXE5U6aYMos5ABLFqSMXomIkVi68LLuA3Z0oyA5QI1+xspkRoID0wQRx4/my8BmOjXLExTX
DTMbMkErkbURf4vkLFOt+63EAOg6bEhsb9q8VOHOPrgAnTyedSQxT5QYzjyU5Kc85OCYzO5g1+Bv
T3vZlbh6BJVlUiW4shq3JVey7MSPHZ9StxCb6nK33PAva6p6AjuKS9AS79GEBDbS9dx1op4/yWkx
qG+PzhuEiDYKDVNwj878kfMDlwx0/3zsCdNskIjdSQHjS/dW3IqgYugyYpx657sCg6MOVyeeGT2U
U162tiS2cTHzTujA1/0+mk40i5McJuAHAEmuOCLU6RlokLhV2lXcxRhZyk7SwT/2ib+5Wvtg3KVa
BKahdMwtmaGb4x+bMYv83gC8bBETsscHWcw4C3IgV3ILQf2PXQ7FLCL8ySw+HGJPLjB9emSI7gCv
tPtIGLFrpm7WawSanPmDMWIrnQKd3ZQrugZZ9IOfUbWSo+1IHFlZOpMf52nikFRaa+xuZgehPXjs
kCZgP9AMPvJjZu83i0LzNv3vqfeKOhl5YMCVGsNt2bS5KkUNDLdTAQb2C6h6Cyeg5X2iycBeuoLt
98cRa84uYvL+CbqsEJ29IBBY3q5RK00jAvCUQ7tngOTV/iSaRNVQoY7WAjsgqEl1Z/c5rtp1y5eT
QTMR6W6/oRI/ijvi+iyv1LQ7yPqaC/JDXbvsLxlUBPXZDhZLdtkucXZ0j/IKA2rXtXco2L+0EK4t
iMHq1ovhNHifO+Wjnvad/bf5JC0yNoV/OxsJrHzUHMQ2bs1OEGrWu3qhiBZHfIbD9kZR8RQ2sYP1
LGXeVQGflv22qBibquoX0FbmzcQxaggi8FHkoQxElfhM+j9QqA+BdLun3CR1crZdo+6mfr1YzK42
u+ZlNSN4RRWpCVb/MIa9fwUPEkgMibNiNeXLX8n+PF1zf++iNV3Kwwn8AaCmYL6xwI5fGvgbqTg8
5UFSEbNyfSn6Ag702AvbwGlOBZLsK2ngmqiMoW0t3gPqVWCZ6GBRgLAk0/MO7AHHAK98ezoxaMpV
gNy5cZ0lJwVrEuEbOqYOMTSOSK+TS+hgvUdF9JZYFqa2BXwzHQLoS/FC8oYK7bFdOtkHiYDm2J9P
jvKzFzxlhqk9CbSEZpR584amARQd/uTtDoIW4WVyoiQSrfX9z2tWnsVTbnU1IPyoMJzxiKuPg7FP
NdLM37ga9/CO2oG1SCy7mrRttZ6VEWCEEWMwDfqfZWF5tZieTl4MMsdwctjqNOiNQz79OimD4v1M
O7kvROgS2Nzj9O6PjyJzb2cet+ROZpI4mbBCjHNZhp6bEXbT+MS5ZbGHMEZU7TIpp8h8RPaxRFJG
imlwbJL6jy0jBSCz2Yqrrsl684gFTbyoJpcl9ByC7jE8guHQCnCRmgAaTH7JYO3H/0u26gExUGNK
q0cA1Mv+7m8ZSO/gV4zy0y92lcImelTyu7W3y6XlChY5geFbCg9a+SBmqwoERVfs+lqUG47gkfjZ
64SfJR3uKWqRsyAKRdX6jLnMrFSUjL5VWDFoGZxy5lrPvR3jSO/KqCtY2Bi6qwk+PC8x9PVDO2/q
egok5vis0lArMZruwlQYXSTUsd2LdTzJcMhSfZdpqAzpgwr+O153rNuz+3AVyeoU9dwsqj73PJqa
Y64ErsXiEGcT5mL+i7HyoG/qbCorQiuoywMaqe+NIpD6tB13uJC2sT4E1BPc/MGIpSt9F5uFV5iT
yHSu8X0We6catb/Cr8XQLGgk+sjLEx0xY9UYxm3VIJpsoHMfj8VTYzkMrjgoDTKY73r8DfZYtwrr
QfGNC0uX0+LthLGx9qFrhnkHegiO3YIi0PKqXx7Y9Y/5jdtOQeyToAqh4dq783CApUYPmO/PNukw
brnHkoJqPKnq65NthH50JlNGIVKRg+de5eTv4iTjmL6+W3TpSl7IYxEPCgGZc6KLBCeSvFIcpdLL
X8rn8iKWpbnqLn9emLDVVk2c9oIxTOoK3Bw8sC/S1IFJ3BorCJpmoMlxboKnBBpWALWRmOh4FRxS
ABPDRtFwRZjbRowZ7hdTqvnl1hr1Fb/SvdyUAyEXwNhQK4mDNP/g4DeDev5JCgHkKA0Kc4Z9sDxe
lf93zoX5mc1GsAUTS6Ya1vgkVJQtA6wDc6HMAql8Na0nrK70E7Voo4EbDVH347K6z0Kfo5xGhb/n
9kgclESSiY+1fRp6O2ZFs77UUibuJ+/JIv4+eN+Rw4pEwIOoHzVyfDbTJyCHRX5VaDlxxa/BEANv
n9s6gdSv4+Y/GtKZAWPXqbFvhVNN90BPYGZkwLBiw5InpelAdE4K8xUPe+Ib5dFFV58jDE3rZMFN
63iyGyLGPNyQK/0zgsAZEwRNY8qK5wMujAsuT3K3uGOFDdRHiBowN63eGgcBLXchQXR5VLzLYFOH
r/M7hNRoeZsJEaua0QwV0Fisv6baF9J5QAM03xCeFsJ0isMeM9kNgx0fshWwU5CFZxXnB8OvhagP
4AXFrK2IWp3gi3FG4bm+g44JpTb+zZYa/pAwGy5YtUjqLxWm71wsVi4Efys9RFICQRWCLzR/GyU9
2vBY1EgoXtytFcFGFAwURhsqb+gbk+ng5ZSCnn00pf1UhyeukvFNQZBQPn8wBAJQGYIOqSFqU7zl
L4a1AIQNneVqgcq0iqtA6xlOa+rtr/fChGsZS/fJkpaKubVkrmFnlczxi0GR3G8ELu12eu3RHUY+
VC6lDoH12fOr4I8owVbcw4OQlViYEiA4Kk/f9G3aI7lDQUHJlMdXpL3FMIU/TNIgqFKZA2zOjf8D
8sf1JA8oGSLIMl6nZxwBSFyWdx12993k77pGw388woK6QVQBH7OAKNSEaQK6H5jUVj5HGqtTgQ6Y
v+TswAQjUiQrv2odYbKEft0xRB+UMLrW8Y0BRXlGcDo6UFUSxtM+dUbNus2eaYoP0XiLv9G29Orc
eJSoxmiH/KGk4ZaOizYidgOl0axP9C+tZu3wgGUMGaKDokiprEkrqnHhvzmGYGSaB5jlQq9JAPTp
Iw6p6UlkpsJT5EANOcQ/7jL1hpDc7j1adZl0ap6u+v7R4THLX70ZhfXgo88uyxvNvbnJVBKYsJAI
wS9h9o/GHwhGxtEaU/xLwl0rVlypUZB0z4W4gZxgc1JtRtYbcfQRAW/49KFuGTXnkfKa6hs0KV3E
6zcKpG8TbmaxP+0lq2a5122lhw3d+wVZgUOSUIS55koxWGGmYc5Uaoyxw9NDYts+rMCftbT9f5o+
1l2CFPqNVELFIXKowTAD5rnjaEa83hX6UAGCDYF1pcPGPRnxtQUL6dYuU4RTpPA9g4Rv8CE8B/Hc
iN0FEcHjHU0xBwWhdbycEen0Hfl3O4PmQzyH0dSGB4NH6KOiQmeTNn/i+6pJ+V/1gD4Ls0FPAsMH
QjMmx495SQn7yZT+N4ftTlom03Ex1i0ZhnPPfOuZW9Mv1XaC3rIe96l1jHW0SnYf6cU+vw2dQPCx
UBF1Mkr5rQzILVCsIz4MEuHDnLi4jyq3duFDLRIQvWTIW9c+oWzGiE7dUStv6VtW2iNjMbnxLhrU
q6dB5Yv4cQqDQtdvB+Umhl8nnJoygaaBeamvLaXnKHeoK9BsAFhThCS+PC5uSFysFWby4Yc2P3Wu
Cca3MQ5iTZ4cP+ieEc+HeK+XUI/W2TP5AXR8VJqlzA7f7k23G2V4QLtsdahjzyziw0Rw93qTtpKS
a9S1LyM7ZYGllrVNqEyju1m+oZ6cNpVd/N+gCbtoDAZMiPqDtWXn6zYT9ymFpEn2T173Qeb630fL
JqN1Op3Scxs0Lr18QaUk+o0fvExv9rXx7akqtQb++eS1yFrfYNmiuziMcw3wrD8kvn3YxRM2aYdD
RC4GY8eowS4o7dsrOoR6n2Ms3Q1NeSRcDw9Qzrjfy6WROtXaSJg3T6jCjLSz7KzCkS46CmaX3cqA
uW/n/jOyieOXPAmtUuY4/0RfkTcX6vqtRxh/iyCQ2UU8D74eDzTXagpc7pklRSFzUan0QSFq2jxI
YnVqUiQS7OLnZPmMH7aWKagueiKVD9IGMz5yJmYhe29UL+uDT9JGK8NW8itj7aPUAwAo8RPIU21u
JvO4niZNbnNGflJSLr6GZD9nRCKAHoPIyHMo7SkAS0pi0D6R0B8GD1fWN+rnn0G7LT1ii1bJ6qO0
zX1RRoAhYwNhEPqr00IaFQeHtqLxX5D0u1z/NDRGZyA61p1VPg6/gR7/clt4kFDQDmlVli5jund/
VAQokX7aM2AwIgXtrLoorEoFLyjCYlzbf99BTgn48yKe0sxE39EdUTLF9zfOY6+PUQS2UYTKuaaa
JmhrL95xkCPytgAieL9Qoe9V2P6+WIpX90owCmpZw2fr7x9EasJVioQyzSDkIx0NAvqWk0VvBu6u
6ZZIErsYH/fbHVGQfslwAxcWKriC7Kvx1JEZWRy31pG/q3stUlkNcaAAL+ian5CrNmcHAgKqR4f8
Xe4CGdImjuoQPjqBlS1SrlTCLHvk9FcMbrKR3sPWCUMf9AqHo1pQV/Il8YO6JpzXZoBhLSV0JLWc
kbFpnDM57I5N0VKL1dvXRQzX0KoLZHUN45pDVN/ZbTTUhAKi/zyGg6EhJ0ftuBteN/e8hvM3HxFo
rCze3NojiVPNbZymoYXIlmZi8qq4gGhoJyrNsBxBQFZCSOCAFRMP5KuCy9xW0N4hkzv1tRKtbnZb
AOh4NN+17B/1Wp8SQbNNxkI2uh6jtHH+NTkLqbq7TBvbddReoo13Ewvu0eXaqLIyZf6SZcmef1pj
dNHJtw3NikFo+0oPhzDsycq0Pvw13EXI+5p02xQVsUAjn05KrqimjLJoXhk4WT6nWfUPuCaBhsN6
GVPFsrKxuzH0ciU6RJrgQDsFpErT/bo3j5yu8uwYg5bj4kcNmBXcU2FTKx9MqB0/FtizAXMAYGUo
UEdKDJuahTTvHApCeMkb/Mu8cMTWAczN1ix9X8Cko0dhW7EpB26ATM5ElCKVZ7MPw95AdW4doLme
h/FOWfI+kOOc6nl0H8EvyTOx+3oH9NEiaJNjEaplJ1HsVDB8zQo9MtuWSwpMvXVTRzI/MuUC8nh3
CC0Aq9v+c1ekzzncc2Oad9cfRfgUsriWESGOYoP1SVnGOvN3vmQwO41Xj4k64KfsTnEskURGYVud
+3EDnJyfyfZh93JUBTbOgOgWgrFGlnCKFis2Wh3ba7D6MlPmouUO5mq0lr34eMPWfuekiATpaFJc
5c7MPnxI2sNMHYlYn0OvlMqNn3TyZ9VboYMK+AhGGAlChl6tFb939t05dzI6J6eCnDC8+PyQryiF
sUVUZb4vIvjO7C5SquZtCQa/iDSlzveTSZNxk53yEBf9Eh0KvJlLxuFIFrFz91vt+4Mfp8mHvt+3
MKb+TlcMKqkx47TN6nyEOgaF2ezYEvFfG1+OScDJoQg1eUVRNU1y7PJY8xXDLkMgsqCZNsOoLmIW
FUBnXQqVIs0eV5Gh7u5dmnOrupq+bF64fkR3NknLOfwGb86vNzmQkAL/62aun8Y9y3GkEa8nvJd7
VKzIe3xxYwTTjfcgrMF6yaDPJRub8zD7diYtplJpMJcFM76meaa+1+zb47BTYMLk4OfxQAZOpI7N
uqFVa7h4OTGCgtDAjSQD3DRBOK7xIBZtZdB49CSAxqvVdrYTpbx3a7E50eHI3eDXwuGztlbYH9iS
w6k1OXOfqpJxOeeDev1z5jF4ZDEsHyE2RKoyyIM1ljOtPeATYMN3ROwBwVE4Uve0CNhAaSKIT7Iv
U6W+GQpSAHFUJ1Ur3ARQuHdbRLSCebxhszTbgZdbSREMIHV2ErPhGzh0tKm8c+zYr//DO6lXuz2K
9g/Xzv6UlNZZDlUKrGoKsWYFeTU8P//qlLVphFyDetTL3+Sn0urP8vVlC+f0gs7ci9X0eNZiBfZ9
5BiX59GxJ/b5u5SN1LVdgIXMtNjDi9VY5u/ZOEx3yQgJqYrS51KCys2nEQRVflpPCM6/BUCwY+5N
gix0J3vygZQSZ/hC7Zbg89C8/DCgJFAiKCE8oBAGfaASjsLGwLQGuSSVbLjPXD/bBhggsJ9wfSY/
DegXNqtFSabNZiyJhqaursSMRS2WQhLJ7HjuQtQoqwPOBFcTh4tBGwrGMB0uzvNvKCFis0jVxKSg
YlgI/2bVU1tbBCAZSQajAW5wEe5Sul4FjgtBwEFmr1sWURyW418/CQXhD/zGrAxA2MLrkRy+JexZ
bwPc5JcuPQSxmnLjr2gE/Y5e0z6Y8Mc4C3HDjzA1pe2+5XMB7gqqa5XSRtIMbv34R5D4wvuwkzWp
RcJFu0gWTc73xnz/ooI53iSvrmqoAd67akSuGuPuKrQNyastc1TMnta07x681VbmWLS02SbUJI32
W/8qOS3Oe4JP3ujk42jYnJGWbYahivkCKwr2WgIdgwrqtdCT4IymU5iNAp+0ezi8YK9JpjLEnyPv
fbkTEP1WLLpZ6yqYMm/HZ3nFGzB6Z6QYjcXZC8NqbQUTs68skpKmKTbL5zasYb3xrmopeU6trn38
6iSCtDOyBzLYCGlvm29K8qMKRjQg3R0ypQ+xFDsPUZTr8wq8S10D6D+UnIskDOztHx9hIlVBA8j4
056QRJfmehnCEA6cwj3mTBL87RVjQNmVeyLyOq4zs1Xm9xj+0dWumdIiXj2D/AV0DJOFtMbslzOR
FZra/7fvrEZkJ/Kw96rwuAROEO+i3nXvvRyHs2FHfgmlRornNBZnuBUrMLmdgvrwX0k/jNvxWkBX
4gSJD7g+A+4XPZdxoNFlRhtbevmqMLWxwzOtVtxsXbqSvjEktH8JKaKlOStVbBMEJwA77nF19Tg/
3FLLQcg3GXazCncX6KebByx5KwDpC2BJL6av15rU6b6SkW1fswdLy58ucShMKHvmzwnxbFkIsJUs
Mu4qTr6vsoepDgS2F3ha1TcPLe759Yifo25UlydHwhnHoqff1yBt2+bgUCmqecjLMwx1JhdEAdFl
uLlNiQZyJRtrLWv4OzOTcboExKARJu1N5xgNuHk62UuQYolxPrQDQeQ75Bo0G2kUoeMsJhy77CPp
FWrAeFnSzl8kSQbfU7Kx0GfJgcwUms2xl3okUqSiItKUVt5kTz0xRt8LQ51Hf9XSI801B9cQwLam
4idy8YigkOr70c8V1HHJIMK7MKJ1oBbRY+sG9QZybKF3Q7hb4OWQ3U1ezCgSOWGaapaMe3eYRTaH
lW0Z3pnUV/1TjM9xAN/Enl7XO2JnTVdagZjgY0YKLvpjQLWDBGBlweGUTKqeODFm1rQG55yMMf5h
A5gcOjA2aoubRyoRw1bcts1UyeofweMb7iKR7IteyBbNjFEnO1+ix4FRad4Sb52nHSFcd3upHnE4
MWSuUg11P1KmYrS8YgLJZIEUC4ZBfbB7pf45aXXm7Ve9DZqDz0SUvM/cESYVZxZxjyw6O/FE4YsK
O5bHLihQY0LsOdl+iyI42trda7OFwnWt3/hMHYXeahD/BzHaxvL5fyfjf9UwSIkIKc3CH8z6t7mh
Pn36zKnA1ARzZWsmbOR+tF2QQs2zEeCS9raqbPEM7wPMNIvisEJp7HVht3lr1lKW3znrr0clORQd
A97HcjumC4Tg8b9/+FmX//OI3gJVp74BGyDqG3lMINW9NtS8VkfPZ4Q42UC/yYtjIMwnYjoFTJID
JmHYrgtoymtnfPha1iFifpOA0uiYxdh0aSWqttmXnoV6QTD1A1QNwQAjrl0yRc4fZ1pq0/jK/e4v
bwDIwHl2BcjRlblIdlpEeyn1XLmYBaHKdz88YOnHLdIZjyuAewzDxEnn9vVor5kWUgcjbPsUU+5d
Xt1BQo3x/nuHNPbQKdRtDlId7QF/2UjwaHM8LcQB0By6Zc7iKyga5hPWwZqTOXAUn5DpC//KzvTP
rz5H8GYlm/7lbbvJMgrhNMJwpKZiWqsQf0FcabHH20wWtto/0M5LEp22A9zXzMQ9yTIGnZZInuP6
p8PmBZT4vw1/gS2ZVAISSSKpRl8LeJVFjEPO32PSxHo/cKtNmGfrve+L9RfNvCQLLJdTeCpplC5b
pXoYG3br5kMSVYqWNy7ij1goJ/VHNd+azZaFDdIDJ3VefVeq79Rf5WqG+Xl4BY9tvvt7W+uli8Kt
DJvESfCgzMlUpxet7HCcrH/6EzmjgskBhGD8rRJOZkdrchH9L71DT4p4Cg84wyzQQuPys3BwC2bV
S+9hrzZTnLIjHw+8L7EBgYEYtPmBGIo6tOL4mCT+neHhCG9ELbCntgAO3CRYhiiTP0Bzok+tNqXd
Rc6M8bh1ZEFYJ1l9HYwPKhvfbIFwRSH3ywLtmV1eVUCkYaXUo8xieHzTZmIg8PIZExiLKzOy/VaM
YTz0ApHyJM10NvapoJE1tKxmQiFGs5V4NTNoqxQZblvEn1xHzI0jDeYg7Cht5c4XJ5YkxUXn4EHY
0l1+5v1G4w7WpxvnRCF8Ma96RF/1VFbgIBJzQadVY8xO2Zspr2zI0kxdF6v4pBFRQM5d7BRP2mhr
W0Il/3HrmgL8Ibd251pKvbtV/2diU7RjW6x3K/Pog5D84Ujop9qZL+XtnpMHcRIgBq5Ec0LilOdT
NgSiqxctgxJnur+8HvqXrDouTz7vbukvMKTKbS8y2GyMBm5hTSZFzQFZJQPwjZzw2LKJe2zohdE/
BCx9apD+xMfDDAtXRQB5uXr5fL5ZnrTIXXf6pxED81rdVGL0Bf071nE75MIMH8Ugb6HZVWFSvSk1
aDN0yoxovQ5COwZp1m/EqyqU0DjGYArZsX7LstVFFKiJnFrfYeafyzEw8jbWCu8/qL9/QR//DDOl
B6/lyEU5qbxVAfrj563+Dhwd+wqGQHqv6pgC2+kr7D4VxKU8mskRq80HZR14NjeW65BS2LN7C903
LTjZGBvexfO5k1kS/hiRpPyNRln/NppaEyeIHzVsjD7JxabT8xp9q4ADcAnONYgfXjJjk5j2ttSM
UzyWyplR0nH5r4P2j1ILNMu4/lyI4Ml3s/dayK9JxSAt8MaGnjdYzUjYSwhZEyFXHP/KD5ZFs7SZ
5Q7ROc2aJnHPp8cMr/Y7XWQjuLW78R6ila8gWYyZrgCll6JuAquaLwoZcxE2BjpBtG+q1Q29YKAQ
27cSaRPRm6HwgtZFMXvzbF/bvX9OS+TZmNv2R2XgSchOR6hXS1iNu+L0PhU2MqiK4F4a8UvsMH8a
0DQjUfgLdfZu9NRltefX2H3q5qaOrlmbhek90/Vm/z0sQDGuYm2GA0YKPgoYSjzllRzNR+Mn3LVR
ECrEVCKblYVkywYPg1STKBktODcOGMO9Sy5yXjr5Qo6YqiwRuB2q2jdZ8jzsKDWF7Ao7la60FV8D
/Wde2TmdetSwPQhTexTnsfKgdv9vwqSA8WV/pf9/Szc8q4WbwQ/cDhA0G+CDq+1B18ZQLRDs4YMg
WbaFfL8kfIFr5vjuwXUCA5udUDLMERh4Z63XwCrGnDaKL8xKpMYzwFOTF9w9/L7tJAc1Po6BwcnF
MXIJLKzGzzYnhTtayW3ByDfigb9g9rJDwPtD2KQXsuBCQMAZR7j8HPLMf2lUBs/8iM3+gLQfFYJa
3wX4EnfIWR7W+SHD+yz7gM3UFDpMzYQ27xha9H3j9vktwf0px3PaGvM3SOuM4zcF7uZqS9rnzXVD
T3oPCp4WtbsjOqE+LS7l3MrtBVews7ohvj9iGlHA1+1sjSeT/POBb7j/M0Lu7bwOY4+TA2hEk3Pd
SdFsRF6Q06t9DM+3mFqoZUdkzw74cWa8z0CBlMrVwE810IJ22JpT+Zve6MmwXoMfcDVVreKHPj0B
9gkUHo03NyHTxTT2dM7IsNJRFh6da3UJO3WdheE+jOVczb3a/HFNWQO6oy8vGXKCZz50Q75vej3u
aiCx2unyysj7DRbEDErZynQeH/hN7WTEbbuh3pHgeTXAmzAbhsSFoAgz3lAEiaEYlQZoAt3Y2lxv
LFchI/vE+CZGeYzpy8UqFUj19098GL9ZA3CclriEJa6BKp1gEsQ3s1p1P/tGoPULFmKAPFwgwwSS
RtnczrNqVjgbfdnk+LH9HNgH2gZuZHdJqawPnQKsIYxwe8n6XMyXwSvYQ3K/dQGaRvimbwLiCdgg
LDX/UMYt65vmkR63q8XO6s4MitkcAgKbOmkAH8N8PZ3MvgCndfNiXImL1ClkR2KGr5bZlKLzO/Qy
1nI1iU5ySIp/nmXWfT7Xk75d7LFZr1q/RctnWgh0S4ErAq14OTXIilg19vOtISrNAIarBMC65K4a
2a5iQ/Jwy4EEMJwTk/u8W2QfLLH/HG1klA1QyqewBMrM2Jl0ofO8Uab8i+1+ofQuQoVvXfBU/fAW
80J50zaqVpOsqiLZWxYn/1yBI9aqVf5Uta4WVOpSpeJ8pThQOAh3Zk0xIB4ptMnRZRxKsoVliN3L
/jv/Mlseds4HFvm7cFmssYGXM87a5NdSMhjDr/IwJ/1NIvROBBi0SNBWMp3aIiySCL0sDDvT2L7i
jJgukJt1BNb+H/hge2Ge2f9Q0RHuM17j0YK9NF7dCLP7znIJshiWpn9PA3red+iT+elPqXR74vmV
KfmKLd2YtU2UM1VBnk1YBMzWCZO+JUL2miGx0FSwhyN+zNQsXvbcwIvTJ1ieIh2hmOUMuZng55vx
xi+0A7sj3KRZ8B6hzAV/KE3GDQxMpPBWIKnGKtgYYfM+eySGUkQp43cp2AdBQzLRopIsXkRDg4YZ
FAGhHxsOroNmccL+McvcRd91Njf62K/CRBYGkLdIB66CRIRf3v9cKxO/uoHoEDVjK54qHy42M+NY
mZE5L9I8ELvZSAxaDShcgRATwSsvjNoh+EEo4ErQ5X3BnblEOH4yPpEJEWICOJYr7z4NS/n7lADf
aT4VDnj1I6Tca9g3Q5rDev4YWytnu/Uvka0qU/PHkdwiRYNuM6CCAIhxMg7fi2ogPnwIjG9zoHdm
/ABwEWxsfuMCPXVmC51LLZ7WeROFzb6MJNpf3V6tGTFFb+o55AZkZVK5rmi0uJOaC83sAfYnywX0
P7nB3GVpe5mjB54ySWmUhd/qEhIlGFJ2c2IiwnobYn88D/32dBRHB6TOUt6Ze6+s53xEPGal4gmE
Cf7ZI4fwB2AEaWhFOIC10zuhrTk/5O7pXk0Y89BM//UNZH+UfiCaQkDSl7e7hBalez7K60Sb4G09
8w7MnJFavCcDBVN+gcnntJzjHAMGCikqTQsxtfi8jpZi84cDP0oWyzZRId3Gmnz6J1BrVNsHqN64
cLqlqbejX25p8iDP7k54OC7nz4sYUW99YUl33CsQTjgtpAmQBeL/ZK+GM6uPpaMEvJYFleeVZFj8
rs0zPSCYO1NiWKdVoVYhZCXKxSqTVcFK706qTsGkHJrcRanJkR3BqbmKZBFyRVRKfPiIbLwJADmA
4SVHZmXU7KcaEJGZvsbMmYulMxtdECgNaELNt12xoPuJtkPaACbvIAWjnEvJNShf+4VL0KiHNwUj
XXcDX89kI5lHrjI2znIpu+TfosFz6P8b6Be8aUHt0+xekoHs7Knb+dwfZfxsgmXaOjZUrL2k2tOZ
FWvJpIw0u/51/E5tqnNx1Caiwbsbc0h/oBRN760t5KvYyts8V7JoxeaR32fbwoLP2ToJPG8YvirP
YXLQF0mLK/s7sdmnxAzmYA82UmhfjlI+u/Gcz9pOkRdICi1Ny/TZddBj+1eerZUQ+8I+LOj/LVgU
5Bren/cSKKwuz7tIYrOdrzBpFVhSgf6UNEW0McQyFsHX0bheoGbSgR7nrBppWFB+9gO1CutW+vbV
xnLNgfzwfwWpdY/XrXU+4yIs5BC2YIsFW25ebsveSmZTCwcFCwqGpD2TUZ5b+j/gJ30bteh4krHi
0UsP7ryuLOHI764ppvuUk8926nVhEGkein2VAnZ8CJr3ZeT1rbwXdnJN8KOFhOnc6NH/8D3V2mXj
E/oAeuL+JO5tVJO1Iuc61sWlUiJw1efbiUG3OQ2mFC5Xij7GxVM/2YL4ddoC+eWTRVelYOupbGHV
FSn59E/4pTavjm8a/UVV01M+HiKlmr7mSTppR03ZXPUH/btgHmfBqWYvurFy5bAQ3VpsudlG3OJS
aIE5moAEAA+Q75dycvjjI9Elk6FsvUP4VSqa5YwlRyEKuH882CsRpgvqqmNjunkTwIVifC4z3xw5
/HSytv5d/WTxZi1y0vZd8s2W2OcHU77PSzZe4SI4jY45ngyDqI+G+W3VdEI2hYdhS6/iq1mOY1iv
bXhW8lo57FVnTiPfbUYc6Ebblhb3B66/LVqRIYsv6VjSsWicAP4EVqyzyc/HoaLcaVC34rrICUXo
3oOIW4HcQ8fB+09+IgvRhRd5/TAXi3QcVevoZ6jHIKbmxNsEpRDoTStAmQvNYSnkdet21sJ84/rQ
vDAMmsKW0rknpmBPT/OkrhHjpG7SOcROWduter29imI+ijMaAjQVHlkcht9OVz1JgCGN8fLlKaQU
sQlYIVjcVHlELGk13DYJ5kL1WeRcy1XxrS/OOydrZZZr6JPC2238WxzV0Z7wvJdjrVyy+lFMGf1M
B7btqY4jJ9Oo2Zaei9UulXcrAFn8a8yuAPWEOB0uSKR12E7wczNq3qS18l9lPiR+Lsz8Ak4c9OFd
JbLw7PyT7Np+xF6Gmi1NP1S3zRCCukzUnU9jFEQj/CMd0Qz6/Quvdj0CVgEpnBQw9A+VVoPsJ5BA
ux3uwB/ppwGThFI53Izp7TEhVLhp4DC2C4qfX+cQFf7ILkGmgCe46UsQjnKc/QwOVJjLk7nathH1
1AUd5CFUEAfNJcbB0bdjMc8uof6O4FEFrLRxN3txczXjPVJXkPHyrR00OfkRfkcyBX8DeOFGvZgn
JK+Qw2D8tJZkfm0PbNfI6IWIe1/hxW2HSOfzoi3rMqHDYbxSwYiTIZTiTGDVpetjoP9eiU7IEJof
p9r0V/O4s7N/OMP6f5KvLpV41r4nYnbOtly2NuXx3ymsW4exgZsJeliDjiY45V6lrnfMGQsPDXHP
EO7uVB2Tz+XBrbF9oXAcADNzHDgi1ZSm68hg8tyFkdJAQA4+QhwRiUjBnWyzd/rKDVfXvAYp/tAA
GzP4KRAv/kvqWq1qrxZT9btyj1eJbFujyBWcgDaLKnw02JVIm5XtvnyHhSdarF5erKG+D1q6Rs01
SJiO57LHwgrvlLwv70UlcgpJcqGGvTl6an7gG6KHYK5by6/2Qd7PSpCxPYQijq8zbbTPeyhOk5/C
dts67XLNtuaynspwXJk4HfEqcNKerkRy7e5l9+oAYYuURMX9e3FEv+kzWsdSTcMAs982B1gwa6sf
61BCt+XRWSt49OnADbzIRfecYJJ5uezNE+fNP0WFWsi1+e9IhQ/AT0R0Qgo4cKEY1fRsUmXAzVvd
8GK4p/Hgs35k4zvkjzmMg4qoOatfUrY2glc7qmZCgFC8ZNlDkbO0WO8BzUSRCyw/V4cPrh2pAkO0
BUmiueA6c+MKRAkQ3AoZo4ONhrM5+L6gn2FnVQJVZKwGO8P5K6FtRufS0gmnsdINque71H9YWJyz
4IX0X2qoFOg10kE7lUAn3f/czqwwKsQIonlZnCf9aEW6hgkIQyfNfJZVflLR1/aKRcmNR3lsT+yi
ASbgTPViu2z4kunwsqp2+tOoIN78pjj7R3Ag5IXNL8ciz0lQZT7OxgM6vKbwUg8HEJKQxRDcrwl3
nSe7cP5vfu7GAWtGUiFASFrT1bWn6YfX6NB2KVKruPOYmzXtTVdzw6tMEwxbDNA75u9TAj/l2VOU
r3ehM11SWf/G5nOOK7JILsKRfoRENVcGQJBz0MeEdVEcKU2efhkTMLYaXack3tzmQhKfkQpcVHgE
2Ov08i25dgmXGpv6HRNkYLUbwsJcAvSyfXkjMk30X9tuLXiJlh1bKdjSyKr0t8aY2VPBUqbFSq8D
hAgPugkhXHHJnKEBaRvUWy8WHHkjzO/+8cuK4SHbOe7TeQraTV2XkeAOuqzBaGYpWCxhQXJtl39a
Kc14W14tK62BcExFYRJxO5JI3bNJLdO7MaFbrJXxctvHBhw6FnI4pvElskzTb1UfPSCjbaWyNx0O
kr8/bYf8sqvI+GF6Sj30VGVL64KSbOG475Dw+tx6yz5BB45fBnKg30quOhVzL1y+RLG/Kv/19JKk
v1nWLntQaEkquu4i6/VcuohqsjLh9xeSJ5gcg5I8OPnZnrmdMmzY1l59TEjRcPYTWmRODIsOtOup
WXEdVK+tAyT9/PhAXlATRmxMhd99C/nkI+RmoKamZbBPKOHzF1n2dJw1KarPpyGQa3c00weRj9MR
1ca6y/e0gs5C3ZJlQ+a8Xp1N2SeeEvIQmaw48HP9KEQ4VIRtbgGTkYduXV4njbUcpA+5Fh+T+dSK
wZ8YRQ4XVnT3kypia4FNP/lduP3oK9cY8mdghmbdLWkJoLa8G+8SfIFpyMnZeTXgh1yYQrMCW9SK
jOKDg0O/tRjfvjvPhLg9mWK4SvUrEaNmf1fgV/7odFkMHBBFcSz5Nkeq+qx0HgSZNgoGEKucDGyR
SzuNC/cz1QDX9tXo6VMIzCls4IaYcBvxkisRN3anDGhSjyLtge4mU7A+C+FY9NqCvqoTLBagJJnN
xMZhKuggE/qjr1zNUsdduWbm2c6yeStG1UKRefpAD/qyt7WwzwTMqf0unEtRZYyNnmjgkqh9C3g/
MLJviW9R6x0Rkz7BLSlPCpp5IYcl8iN930s7mYxrqmPAi20Fgasm+n5e7bPUKkSwJ7KLgB/jgiQG
ZzvCVfewQbwtHxMzpAybX9ta+eNd1GpRE9/fGAGI5PefDes42w0rH31EUdlEyKWchLSb1RRFWCny
S5k8fGELy0JmigiP21PietIaRLw41dKysPDgNvUAazxniHB6lbf64F6qsUY8cFnm3QJAUQ0J00a8
Xwc8YpCu14/krliiYg8Wk6NgppxAmPmm4Ih0bddwPnkbp31PygXMJsm0PwHkdpW+PnDUvRxRv2EU
kEzRPIR8NT1k8NC1KcNnz/XdH71y7Ea/e4HgdL/CT2c/JxFcTO4PURGn+xAv5+tLe1nZuKD43D4t
6TvFS4Hb083H/S5rZ1rUMfhaWdSIPXFkh21Xt7qyXvmqIrexuUjm7h9w1I1tN0oQgI34W8/LHP+p
u/zX55ewCNWyEBvA/HIx+iF3QwpA5VYX3Yaiwugu6XNSD9Caf0H4Zw+jiyrLokKqibOFh7R7jbh1
cATM/rA0L4g05lJHm+4Bzq8O8d4gZ7HCRF346h8R2fLbtRDCD2XHii2xQ8R6WZGbIQR5gtp08VEc
RTtNFaHII7cde64DRyLu/wmxG4YfrCbY14N6gUtfVq0uMN3sLcsaYRNhOm0/hZ6HfvCMwfcIPgsn
lJbR60h7vjfwuaURnak3K2Il8ZjLlBBw7muaO3stnq37B+fBBejM/qIeGWMgATkNmZNIV/PLxBfM
vJrga1NoR2Z8wB7jDGrNIoqkZZW2HpDBucLxQFaN+sSAtzuF4xocA6yjCYlQaoNfRnaqCLJLacpq
SKIzddQFgUr7Qb5wqHRyXRMO5labzpr8iqktazFeEnW7yRYOfYkFXUmi9g5iGW594IyMUfWY+5Wb
eEXoZ7NRHKZgHd0wQX2+hvmAbO9RILWPZs6EP46OXp1Xej1lX+tMSoRBUH7ntr43h/iXw3z6o+ig
/WkSy0/WQzR+8/JQdruXuZ9LsBQtbCOv/ZCjoHdZb/QhHqaR5ss+j8hNxRlJpzWgmxAO6SYUiemH
X6Xl0XYyNlFtNbIifROq2E5vOZXbMMEm6WoShsvscMZnvBuyJSlUJ697VFHmksVr+7tl2bv2TOvq
iLNt4sEt6+rvtTjEOaE/NLv/v9SDCDLPRacUSjb/6rR5KglkvHS+UC7PZURkTXSlRCNnAmLgbYAn
xFL9ULbbCAt/GFw64Hc4UsKlGtSbnofmTPPwL8X3nc419GOzGujn0QFNny+N4ruo1v+yx+DlC0Uc
fxtqhKxwfez/siSwlGIP8FbGC1VzGhNKgIZtQ88X5i4LMv6GsWWj20mCkJsi6FgvgKSTqE7p0cau
v7liGBP3yHA+axWXE9N9h9aYxWjIf8kmgL24CJkdKCDcBC3QFJxQKDgPGKChiftMp/cr/h265K90
CNMPSjdX7NXBvbpc8d/YOlkW0H4m/VkzVzV11srH45VqtWp694eyLWW/o2xcrgfuGP1J0uxSM8Oq
mClQksTTAjh70x0a4seylMTwXTF2O273c2o2u4Ok9VSxlMorrHNU6SduzsH4pRgTudoV30o2TCST
XtBzkDmv6gd7tto290mb5qr65o+ZKRBG/bggvHLAHItWE5UHEgyEOku3gB3IKXqPweFk/uxX523n
wc0g2wYMoBr5UOU/KrHtq6ceAUrofyL31yFsvRvY5qGFyOAAtiRXVMOc4exc9NW/lhqlKvLuE9up
fuj8KYm5wAxy7xZQNQh8DoDBff1j+dd6kLqWRgIh44ECcW7ZC3W7w3PzTJ3kYvRC2g7glaOerVss
+t1J5WplEw7EQzv+zMqduwcRf3YZslQzAPYppqR3RTF9EKX5CBJHHY8cPOalepiZzDrkouZrCvfE
Vk3ent7///iJvQnpjkneaGAO5gnQssExWucoLaaNyDje+W/gN2PKjKAHiNwuGo1P80mdKfBWHEN6
Xq5pFGj9ey6f7mp1CvpiYg7SJD8Hfei6krPeb2kFM40x9SOJj5EFzUD9WOzjlxLXenFM+71kWyK9
g1GTazioIjF9yeyxUYI95MNe8rjEAuurl1AS8XlvTkDAWGzBgvfkVBxnJ+VMionzxz6oM4hhDMSP
ms2pwwObsof04G0mkINv96hI3StvGvFksNLoiz0wgId3oFgYcchkJKyHWfRQpc98IctS803DYNNX
UBU2DikF8cr+erHNMb8az5sKaAfq2Tg7rcMi99awxDy7iBFZ9S4AUGcLPlI/51/PyLRAmpltHzoI
fbVXuvpW58Y6Hbx4S4kPAYfo+cLxiFCVx6Zp1XkeGPjT9R6gd5gEjEUy0hhfXjBpBT/v4IL/1jZk
LRabhJRn02iraUuEEWEbf14li179Q7ST6/ii+LGwBS1UROi2s1c6UobmdorqNTJOf8cCCmQFbC2E
4DRhd3oiaY7JpyKzW+F4KmE8dcsHsspsEkwi/2aIyYfh1AjRwbIJR7b/vuF+M3jC6AFFGe0hmhQI
IZwBNZHoLlVMHyRdBcjrtRM/w6AZC9zMwOs6yOfGKYcFRpV1cLZjLsLRA2FPGFHWDrUnkdtJd30V
i9bkrX/3t8TO6dmdJP/7X4u62H/Ic7HSrsHWid8w0uKxP3H9nQqlqCF8LZETwIE2qXEqXlNotYn+
q0U9lKVOm0PkOdBCmvwbLJY4HcXpVz9Hxxzas1qmFu8vmHqMRdJKp3vKAIssEtSy3GPzVFRWj03B
18OkaK5DUx7tfM3kDIpZmXq4W/JyZUVZiQV4UaHCxGMFP4WxD5oCvvRRakenvPpj3ndhYzfB1P/+
vKOkGwlBdoxs6aGH+4tTbfgkGOzUN5yt5K7wijAFDrledj40DtMDj2Mz498g1FNyN6eqezeXgI0i
BSBFiX86Nyhlmd95qiUE8awK5vCG/yjE9AmFE79hfyw1zeSWNaXhGVKAF6Gy8rdTukhT1EEg20j2
hAWo/2891qOisbjS8IesWo8rG3UTBPRxvl6W90JUdi9C2FDC6QKtdiCH2fy4jHHyH00keMRhkpDr
lnsPztUpWGp0UBr4lcyxO5dp9nbzum94zbCT7Znn7PjRXnT5p7WjpXv9QKrmorzyVIoMmNwPtkic
dpZSThQHWu28HY9NCbGLzjPgYtL65jkMXEx8QXUV8wIlFOQauvkJTjzOg4hcALvXSXVYMY31LAO+
wW147NLu0piIjUSy9Bn6jeFU9rnIlqcY3ap1hn7TjGbmmJ44flIPjTHyV3vdhipQ3ngIa6DiuRop
u2lN9rnRrxwjOSPRfquFM6XKBGopDeSckLF7BcZmegR37OxWojgPFRyEkLUsaQ5vPo6b9sy7cLWB
7M+ohSoS71oa4JEYhG1R0sij57PhhtAVmAWMvbt7/VOiHXPR2y8mUgVMwOlRmHCgILr7UpWHOCPy
e5lHf2jtYgLePZBT9ODEP/37iEPyRLXSXArYWUN8FQ4rC8rQYFIWuQCQgRpRins4QYpwWJn1CYB7
Q0AEXRzwnvCFv3MG8LRRk4P14qRlNUXdZX3Rbs2NxDlSDaXHXSZJbfdYLsMHrirVlVJrxJsr4aw/
aH0B7Unzwo3wWAerbVAH6I1jlHFP6yN+w50MnUaQWT4TVx3GOKFAMkYEGMCV+CFWKzHAAO8x4tyY
BQtmJfrozNo0EB+OqFzggMVQW1saQbbOfiZceoUWoZPy0K0+Do66LVKfHo5Z5L+u/CQnvLml/q3m
rLeJss/+8eif7LesQpY1b7KzYNCFwkaVzjrMZ+ZEOOtnatO3jiZkvSbgyBK+OG+QC9Mqjaq+MgP1
m57jTxMegkv4QdRyuS2JO1Ng8iUivvRuzXixbFvFhGKS3jXwQvCsK+XRKtKDGnIUqTziah4T88CB
cKj2QV6+V6jTntme4V50XrQooz67GW23Ppdbw654+uaJUvlFLkYsDG122P2D84FGY3GhLGQve3Tv
Ok1EwK1hzUSoq3HBxruy/3hkJ4YgnxXKQZHSDp1rfMvPaTIbEPKrHk1+HcQwPSCnaYzGtYh/mgB+
suF5899XIsyvXSQbUx0NF8b3rLf9sk4hNjKY0141/YCam6wGq83e/FNLF6k/PmA5RTIN7w/OsMra
wSxUl8wiky0QxdeTLv9/8YXxOxgY3F+zKzs6oZZlQtDLhAHqPA29osgGHBziqetiHE8v1iupE4Ck
H6jafazGyKFV+29N6d3BmithzCsy2q/XoXL11O0PttwfPHYzdpdo63VD02osXMLXx4YF80K8Pch8
rLe29MEBCTwA3QVZ6x3u0tUmiC/XueY9xyrAdYnQpBzmqfPdbKyow5cXAOh78P8ByVyG0uSQ/+Me
xEEGi1CELv4DVKY3UMo/uz28Q1jsPmXsk2DE31aMWv5zuEqiKb1KNXIZBoM2tf6fuNbS5RV8LLR+
sFCgBzvfxbMMGFuyn/s9HX15rk8snOYQMj12sO+AAk+95HwRa4aXdu9JaOcfx1FbEe/PstpeH7np
9xSgocB9ZBpHM+qILvtVeZURHUuBO0nk+64JRGd2jTHl7tHEgyecTDftzGP11bYWQbd7Vz9JfJUR
KBKvM1zhv/fu5cxxuAgtMhgeXfI/6YcasvnMd/rFPRv1zgOmPUjA5ealFWOLfv2/1buVwzJHK4Vb
wKxit1a0CZxOv3CquBH2/4ntpNe3aH23sSA4yOjub7UyzsnW5OGM7r5zDbjTiXUxeHNmCQ2frFEM
MaxqK0lS65YtvlY7HiIUuq1cMA7B7Xst6MsV6p0Tb4yqG6xCehcbZWjW/WyaDAqrFu4upwS8vCl6
TyILTxs99jde1uCvJDPeD08Q2RjonbJjzVbWMi5XhqPHf6UXaRdGVmPYxIMVmgXHtiFDhsjYUGXK
2KYX1pQEnezQ9ldjbXs65ozq90SD7BmDga9kaXg7Kosr0LNVOmwfQcu6DdNn2Lsy/vU1Df1fGLIN
ljY3uczWbPjUbNvJl13CfzFnffrjV0CD6rIO7GjNjP4ijQ8FMrbODm7I5uUjlk870LfP/5tWygn6
AqQAoyBb8Jjsnc6mfHQstKxVFqn/jN9u/gsfvMKzFlDERsn6M0aciW8+CuD2S/gjMVX2/d1/fFMX
ptlWfbmsMTd1j3FRejMY1rLsojD0+afUIaRzTX1PKXb3WVWqiZU/dK8Ky32iF41BOO74S1yTTadP
ckHLDQwGZY5ca5QizfJUiwDH+kqw5uWMxgQZqQKCcF1bRFYFI7Tfpbt+STMDsAwGMXgeQrToE3NM
VXr8TDq3nOz8LV9Y2DOTEf2k0UPnKGCLA+ko/BlBtlxsTvGI+tNJF31ygbhecRTWQ56qZiB9LL4i
gJSaEIOD9gyC8QHmYhF3QKeLmUr3zNJimjviAmsfnFfW2/VlPPWweEe0D7b3RtZnHmTE64VSktk1
PFISM4SGnW1QyQ2EbM2YXYuy1h2krSIV442OQAgwTiIXfE4csf7us5vfy1NVtphCkH36F8yPTe+I
qPyWePqx1+f4JE4lP8eBDwgPwTku4zAVFH+fxzHNBNV7sKv8rP9s8OH5iIXCYVT/IOx3ssamcWZc
LmGDbVhroFcYCO3NF8DF4olemxq2jTn41wGKxnizyFrFvUfI4ORh3G4mh266lCyCezj1Fo4L4V7R
TjhEJOKHzmshqW3TREjFxlWNDp/fWD8vgRjq2RXbtZtJpiYxPH3wrDrKywPHCClWJ1SlyoVXGz5g
4fhWTwxnvowADonhT4MO5YuwoFXZkf0ZTf+MIKn6ZPmszqG2yf8Ua+eDOyQ/c7TSn9lytzeCOsMU
l5oteNlN2Iub2jxzSE3Jwea4LK+EnEvV8/y4OjbtxB5LOT018ig9xNc6ypBKQtzb4cpylScqHohY
pAolHNDL3t5vXzmvhD6yCyCs18FhSIZlPCW0GHaP+i8viwsECCQO60I/AKfRMgYQqxzfbyhjqBwx
m2SV1urI4he6nz7N7QdRlsePIid2p0eXt5Y7+WskoWN/Y7p9TdEhwDn1wOFgVGZIvk1iFcRJT1Mo
ppa3CiRWA48hUcx7f6+Ai+bIidoemDieGdvxAHFk9OHmoCvdADE5gDc6j52P+gdXec8W7hm1EVW3
kKPRYPKV9YaUPWS+v8SAjrS/coyLbIgCDmHbfQlSO+rsi8hIyE/AUYMcVs8fT6EPuJsPeZxoUU+d
pywQ0y/c6KOUoiscDuiAovSRpTIIbN8FKQh5jvr0bemSZ/N3Lw6I5OtCedowxJPzAqCHKDOwQLYl
gyAR8Vb6pHqvOs9IlXB7BXMQqvhoz4Ay73edcUgT49c9eQZCfZ+uW52dJDYaQ09zKfSwK/OB/qX7
vzRiJ2kBEN8mdBnV4+Gu9pllTlmbr1NWV/M23WD26cVZXfQrnyeGWlRsJ3lS3sWQD/c/hgU747wt
NJckyVon+Pri4MskiVudcLO2htQCmbDHlDQIQyGQCQRFTpPXT4Z2/d/QYQ/y3Ee7e4RarkXp2Ygh
HNcFPnYZsBfojwvx49xVxocgf6ad6F5FL+pZm47K3rvzWXnuxdAAqsM1RPrJF7BHAViF9asNbbP3
iZYcL3U2QYAGkzNawO4VGBzbC8Vadwo3TWMcL0lZA6Ec+OSmt24qkShOqzNujmAytrCzEVamesGc
It+vX3LN0NIBgpgGP6wbGpsNwmEJU0wLqhek0v6cWiDL2ka1UuCILxHzqkdK2oYUZQJdeQ4w2ovD
6KeYZIzWkqIumQMkWFvwp9sMCTK7zLpfBc5FiLZm7PCD14xZM3JUoOEVJ/xeFoMmwScr+XS9XLYV
NsACwqRxA4N3x1cNZyCxyHGLU7LvGsoWPFb5Zx5tge5wfLDQU4Fu8OJ5YJVHztH7voOGKi1iOXqm
rkZuQb960BFbS/Vr8NFQqugGuX4sGZ7t93u/ihIx+fIGpSUjBi7DIjtZpBRs+9WXLGIL2SaAJ9yS
XtSb+Kg+GOXHq2XfT+lcy7cLS3vM6k7P0hiCex8JnUy/ZL/aHq0n5FdVYsBPLBvgTp1YY4Cr9dqP
9PKcu3JZ26YX08YN0YQbQtURZrS9aZgLjo57DqYgR0rqCONe9igu4NbkC/eTHkBqipvskTQHt5tb
GXgKAwmsEZavmkt0pHVjoa0HCcNbIjtz4aefGrfYXC4YQh5pdfJAvHWKzz7ArsL/JMHi5FNu4mox
uvGGLzzsJtDYgc6dTnHr6MB4nT0ABryAetJ8sOtrQnJfil2DymaQQrG1AG2S9GojsxIcQzL5ztrH
l8t3ljBFykeSw4pdRHuIjtDxsMcPop/8XPhlynhd8hLRt1wHddOCPXbqPn11wzcwmNY2PgnkH+as
R7E/o5cPT/7COh8Hi82iaI4T1O7Ik3CCSid29yjKT9c6e14vRMN+z/m3XHn7eLidC8RutAKc5fr4
CbbFtcT2iBIqbXMtboJV7rUuLrqlr2AkqP2Je1SNclqw0if5R5TOo0D4KxtIkqcTyNMmAoa+PYEi
tM54WHPfS5E+PkmuS/5unGL3OEQcxvJIR7MN54MpHo4MJxfYG8aDLZSQ2qsPaABIaA8wBkdT8j5C
508wSMp0yD12IRpWRr4Ozrp5J2V4LGLUnOvWn05urqcvmJu9XhXZCEuOGJ2PHdsDdsWbbQ1LjeGi
2Dp73IhuF3qbseWtuTMkImdt06Y5mCACO+695WtkAKd+4rq6EXVuHzACa8Ps/ablEUUo0DE84GXp
CqG383eZoGu5jI1q3x3wboBJoHzKdpwzd+0OTvFPOW+biCb7PX0WC63Hsnf0Iz2G90UAstaAXqGM
asoWlEnUUboKQhzkFVIiRXjWpI/o8NkHmHOdYdc4Mxi3QLqFBd2YgutSmjDhnHQjI/C77Paz79yN
y7w8U5f0yZdBmn1P9StFa2eUiNh80dvHO2+pnf+yJnvswZFl0ipFJHkIk5JWc91lto9L2+Ip40Pf
yElZDpONmxrM8vCbvF3plVvoP8KzxSeCSmh9KqJKIP8U2bEKb5OOgWQzMEfNhpOSWvBXpU4aQwge
3WbTscfohfZTo7XXiSKkXgKi2y24jyWeFIxw33q9/rTBiHBPJuJJTSHZsJw5Jc4bCNDrxLGXM59C
xcpxWB7Oq/+PtoJRTDSplnkX8l6cKYvUDIKLy847xLPacVeiaMynE6GcE9fBnCOiPVo2GT6maSKL
GkU78Vx/3YGJbhUvElGtBP4t84fi6SGuZTQCxKAytNwP7JPIMaRJipe0gAiOvDnN88YRemfqCyMQ
rfxoLoj0XiKjnink4UXAn/LJU26Iv9uMFJtex/sEVCf3eYSd20B4NRcmG2n4qnc1Kenh4o2L7y8b
avj2F6VP/ZKV5ZtTR+t+IqnaiDmhYn+ACnPanfQmm0x1mMUZyS5RbHwjzweSgoK8+t6JxyLZrsEO
ezyFyk9Pe2mlqXKsMifofMYCnbpT9mWly6IZ5npGPtpruu7qqJfN+1KRksM+oGMhkFlicR/r58Bd
AfnKgmqsReEjTNecyu/1F59EqrAnif5QPMlXrsed/8IoDrk0ZgslaeFfMiBYhWjDfxHN7BVFYVWa
UAiigxYLvMJu0LiRkJFXQ8RcE+gen1K21TlSuHUuTyIitex4rv4Fsyw1wgwMblRTcJhnNb3Hm2YL
eqg6Kn/Lg5NoU2BTQTDZC7k6FtTE7doKyyi94gfQsCWYViTlJ+VF+wKpWhUQmlIrLszg3dX2OyDk
MnnDcf0WbGaaWDcvPn9Fdd9v+mNHDYxAonsLhGdTArnULyix579Jn/2LEqE7XAWLFi+bm+WKdWKN
7x+UQeQYS61bWaZS1XXxpPH9etDgqGq7CjJUyYA25MTTioofpjJlF3vtcz784uq242n5cQ91+xTh
fXPc0j6Uhs/QLA4M6wGfwGn1ts34Ftusxd4ypGTnc+qGxHeaAmKFNMTo0kcJ2GgNIJEnToumocuu
/zX89punC/I6vIFBdnbW5u9xcqI5+qXCb6o5Hbib3/0P9xartvOCk4xeTFNQBjT7KXIi437kgAlH
u99fQIsq24/frXAFJqVbJ4NK7BCPlSZpaL39YIcjOA6yUyEDc7B7+obuhukNY0iDZo2y2HreMyu8
ChfXhjF8FmhhZ+5JLDzhBD1n8Qmm8mpiVsNqoRCkMUgofzgvhzkcwCKuDfcTU81Z+wmQ+t+2MNft
k+mJWWeUom/B7xkfM/zqclWKej25IOt3dlUqp3YA87fd9VUTTITGRftMZkzg6Uo5Jpstu1QP6Ldh
1PRqZw5JSZw9Jc51fRB6H9Xku/ptaDa2mIYT2lBWCG9FwOx0t0qDcIYHD2Y68szhEb/fs8sIVVF/
4jO6GQJS/y0vUjz6M/naC1uNuMwnhdzIWnIX9cka4Q0VSpOSsHnugfmywUAglAQUrDFpTZYgoczB
ImS3TfAajYAE5CkY5+iCuCos1/+GuyCjVisQQvgtZtrQYJ823D8pn7eWUptF9YKk8l2YNkCLk17s
ujlr626cKXHMsM+AHAZONojOxhIdrIcrk3VVloFtzPHQu93zhEMU5LNWx2oVDLkNfPNKFsKKuE/O
hEArf/wTUubYle3nU+QSRKRQEKHVl1mhsVgrPuMT3WLl0ExcK6DTKeobRwRBzMmKRv6raNM7/Nz2
9oFq7hyAnUhSbNPnZpA64FEBTdKDGyJeTA8KlSZqf5qC70WDe3QYE0B/4lrBs86y3JKnHmFwtuMC
jy2XVrjWy6eCbHdaL9ndMpvGfG+xImf4o5Aq/9eA1x3pv0shEClbHecLbQUfhPvjE8TZYSbJCem2
+N7p8w4uX3kn06vjhmzlmioIAT/Lf9/udf+cj2H/l5QMe8o3DKL23b5U9qATNhGBehZGKCLt5xn8
k5xQK/FcxjWJW9oLLVZsifY8JdPq1QNtT9+WJ7cl1M31KoJIrASpt1xWJ+tEF1Bw1gYvb8A2hU4u
Zc5RwPFbxR+lBsG/R8AhEMItOCGFfMDuyHEPcqif6BMPT19q0IoHYaKj0hP8mtRl+qDx4jdoEwCT
5757/Qldx1cv/IQt/49eVoPpvzpJBHL+RmWFuufEhuORrOo4AqqRg1pylHv9B5AGmQOnZw375bnx
ZTj3dcRCXlZ6BagXU54Y8eV146P+57N0J9azcz8f8+hfdb2HsAXQA8bbTZkwuO7yIKxAjvdMUGHL
zrzOzQ1dsetoPYk8J3CyrLYVetLD64xP8ZXfvHyN4r1c5qQqoA3H8zkpFCnP4bumKYejn4RV5XVF
msePhmkVyUqJpNgaqu5ParRIarYkeSvVyPhYM7JUwJ0BanFKBIyUNbI3EGVdudfErd39+A99MeEx
ZIO4C8iutCNxtG8OpssaOTNhsrvfA8uOH80EWuxkPgV8I2SBvgIjCLTwK+1JokjdScUlzL0FPOmB
liiFqztANsXTW1rJA4ygUw/WyETMQy7P8KU9Ne5OM9gYgHDHLS2JBAUiVIvRP8wiUrr+B4bvfvNC
abJWyYh3RM7SWWRWgNDiFWqpmfFb/3MZX09qHRLtwDIF/BjX9CRBHyXduZgRAEwi+yT65+Dm8Qz1
JfwicJw3Dg6CYUOJZ4jCSW+G/bmg9FJrNJNLihpBemVkxqFma0UjXx3lAZvfz1hM4o1KwTDWJAVC
OMM9MzDQ18vTDM7gLo5KuG60WKFga7ss7VnpX8K3EQcC2KYj42xDpcy0TKP3p9msytM9eZVIw7H1
vxcjd2jUwGkFns64nQQYITFzpDFPCd4h1GqK75dRz8SQXtBh0sAKpKanXdsijG7GAd++DXDIQDR7
tkD7aJ7mOY00uQ14AE6rQ5ncvubBeUtGDEymlEExQQxDFtaZ8hwEdJ7PSFlPvuFF6nwRKHPsbcqy
a2rrVPnQYH09cJMgliKZNjTPj417vW7r4iZeoCAdyEHhy7WD9oqMHksn8LL6xRwATO+R5Ap79iBJ
tEFe1EGchBm/PKwZ4g1MY2pbLHfjwAyavNw61liCy+I4YfATNYT2j5SZKRK3bjDjb+jlFf0Kiaw6
8Ov7ZM5BxSIAJLm5MyZacQMHi922w9YzcrhyJwcxfwP+EVSpNeSY8PD88Lc7mkE5u2+bipk6apvo
MsA+h5pP4jIq0KOasKvubPfA7MwBJHUEg038vzpy16LFOGB7EG99ZYKqLb1bWSe6Bxz/4bzeoPVb
4Lt1+UxTYmMWGL1RKWCXfHRYGcf8GPyNcc+ibmuOkDFlzAueONbUfGPlr2cj7z9S0gfmuDkiAgtj
WKU3GdwKxMY52qY0SWri4DAIAjWzAN2kz4vj5VY1HBuyl9b/nbnNDWLedCDF8TAc+RWqGFXxkFEi
4inw4uJCCUvmN0IYyAYRz3gWedziS3xcqgrjJwgPMNRPQZc5VED4i730W6F9YiJepf2FsfkWDsmw
d6OvpWHHKeoLjK87GFfvysj2nycp8VcpDJ2UR+W41xPO+5lvrIZiGpsW8ZszE7KUpVTSIQCy0F4x
bblrozVjhZ5kMex9wGsWkc4Bok3q2PWMX8q4J1JbBUAeJIsWG5txCOB+CR1wZ86BKT7Cn+iZ3Kre
JeZxdlElTSZ39WdivGNcCHzFLdBTSuiuDglHHvYFQP961evghM7ruhvCk5o1DRku0B4kKhoOcLMC
jW5BzLLl5/rDKZTqIUOuLt4E9RN6FSdrXug9iVoMqNbSIoj7qas6Gjqc30Ypo/P3Lye9yEm7jwuI
fDK+eZ1VKswWZ1uqes+0DWaoDa44Cc3fHPpajj5p9ap//8kLwMZFITUPFFNRIS0EYsXQLnZUDLcF
94v32LUC3ls8ZKKlQsuYK2bQjXa5In7huqLsVjyv3e6H5ljZ8OSnqTre1m5SIhKnYr46AVAZi6PU
MZ0xBEioExJKzCK7LzStEepS7tHvaTjLksFQfkT5VkEi8RUyETNWc7HaErlcd96KsBf8NBN+bzFI
FPNZrFIdG0gjdJ5wI0bNxHPpLugpc1xaeN6n6KLFSxcAcBEi3UdkYwiNNtqmVeuTejZpnQn821hN
7m13ukZ+lfUWc+npg/W/dGRjYDpwKMyIdRhaGzDUkxM4GXdKTq0VKyWDSNfCiNyhdzUTbigTd4/S
5z/qht9W3WXrsjpeGDdctVDmUKjeRxtGHJhY6ibUkl3GWW5BN+vtnw6crFicxmcl2qwZ3SxBYGsH
YPbVABCRn8i1Dy16RmDPaU+1pt6wVUYryy3dYiZ18zYPPs+jW0ZMR67vSeCpxzqycnAraWNbdKt/
8eWy6X8GyQAzl+PSMjhpB4UVt2hazuUtb9M4mDa6SkYsOeV49759afPuyYDzLz76zQd+UQgTjfUX
kvBH+mYW97I4zRdTOHEYsfeh1p0qwJuI5MP1/z5pBNujkdqR5DYEXTi0JSXf2Ojx5JqTXm7fIaQK
nygsKaVrA/jtqcLFMWJ3wHvh+6doR/+MG+Rxuztqwf1jWlubhpTs/BubWDC2JP2wmFZZmOE++DFV
BcBk2mtXDbaWk/nw2A8Mp64H0w6FDKLyaydbwbQkiujaFinb5BG2BYGYQjkABgscVAEWJup/o7Mk
uUZyBg5fZ8y2crOnbZ2UEkIh3hmEva+kCtGM0h+Cz1xu4a6au/pECe809IFWrsGHxRM++BavOs1o
/ACpMHhTaEwIeawTU4E/KcWCfw5jyBkOl+P4dMHbq9150F4tqbq7wc/u7ACRipss6Gn8N7KaUdJL
zjKNKQUF1AbL/CC6wK9dKuFmGm2535Ufv8Hz5RJeJe36FQgiuEq8HOJ7ZQVVsd8JDKC+drtStxPf
mptpK3cfpLKh5Vrnmbb1rSp5Hg5tO4umcba57bivDBGWu4KcjQKCRkBYqFN/T5aV0OTwRl9WUCNt
OJRq5ON/UwzvNC+LjjG6tA0tqFJocqLpjOCPLB1T6gGDsMQz1KVIOzmXQcxFN20m5+llFVbnrh3u
Pc305Zy/dS0J4XZL8OFEQ4c/1KXPjyKH2SEZT+ItY1YO1lk0CJCy0GbHdpSzRcB/Y5QTxkNW38c3
tvux8/5hETq6WpMJVxcUQMj8pBw3Ik1oLFC289l/EGPiwwbS8O8f8MTUH0rpPSZwBs9bA40Nt26O
Ddr3AGe7UPE71qiRWHUmuA5zN3+LqenHZVtMhZY13gulvtLT48iAd912wn7miHOjrMFdPfqkwEVR
OlwEtVITOvt7mc4uvH+nnh7pCwqoU2GgjmYZD7k/dkJ8TechgQitZEGi1wHKpwLYArPD4COo+t4p
kJj+rcdeZO98MVnVel/MOxLYvhkoUp+gBC3AMO99p5SZzwEoaHRKQNNw8pscvnPXyUIOzWfm8RfU
NrQUuFFt7YJqaWgGmFu9y+nWPlOsuXoHTLXjV1yuHta85TMFQ0tUjNZXHlhmCORkpgAjW2clXRTE
OjnRNt9NiAvaYLtnHLMoSJQlO7Y2IYiWnUJ9e+3kgk91f0By/VbAXcGZd+lPf/DLHmSBIPedtn5t
tGx3dT0V8q99BYih+wYvxC9YXYFuowD3E/Pjy22U9ygkgdO9t0eVs/MBkbBizAC5YJlXyUisEEgv
aBF7WZYjl6Icj53nBW0K0YyZdBQIWiv0mg2hGalRTMcNOyOFhj1uEE877fomqN5UyKtWN3IaoZ0P
OnbsIk8lS7KkBtQQUOnSxKCf60/5WwJIKehylxFvh6R9Le5i+f6M5RAHzqw4KopGolWM7GubLd3J
Z910JVvSEMXnuWQ+WaTMyBKeSSE0unZvPb/5/9qraYGJIwhNmY6eyZB6ecLae0UjcrUpZHY5atBR
2PSiUjp112pPfufbyNon76sqIB6KDwa+eq4a5UdTavO/QmaNeUHxF5V57MehiR5nkR7CmiCNodEr
oNp59fbEdrqscrmf+715Hu3+yYSz8O1/sU7mo9Wk5WdpaSnWqXN6hZKDW5fH6qrRWeYisE4V3cuh
Y84EZVEpUTXq4w4zFk5EkOkxVKKKL08+nIOqoXWFCUIuFdGjn8BKcVmGc2Vt+znvLQL7lRIcYPBh
9Mw1SnjzX3wUjiriC/7DPPk98Td9EUQD+nnXT3pKW3lKs1D6+yQDchvJQbcCnDRB91kmevzij9G1
8P+hmGkqR3v26V8FWeSyLhWUSTdGTY/Acew5MatT74fcES1eJDIij/ZHvrhlSfrmjATqFbu3axA6
fAKAA/XUi9p6EcIZRsuQgBB1Y5VCURXwy8kASsBgyCNaOmm+UNvOVK3wQIjl3GebooG2aS08dSJZ
xguNL7sJ92uV09SlMUq1ocZ4kg+PhCpyZD91L947QgUoMvNtDYWA9b5fYd/3uwjoC9nxaqYEWxgA
IVtxlSN9NuDk3Mz3CAugMkWUHQAWHfX/Fbv69GQUMrphJQ3YbZHUo52mQhryWfsAyd69F9iEiwlK
h6r3JxBCKBee8irQzi8iN7B55YLs00sMERvjIVJHwzpkfWDkf5pn7Ba7NKjU20WDSaXxM2I4/1cU
WO6XaIcib86/+8N3HHvS4JpZj/DYwNqZGNVUKKz8qnqD5XUOtwDgB3N77ZmpmCEGjfIumVBhsihi
luxp0sa7R49GokDb3+UEubdXhvYb01tOx3lpCa0XnWv+Nmk7myeFVGeLmiV8+X37/jLmNt2BHDKC
Xs0HKzXkY1tRzmATgOOLOx1aoTuf3RWFLvajOVsZjAq8Q436Y9wflu6C5roOzE0LoK6ZdTK+V0eW
EHkQz0nZP5TnZqAwIiBSCIJgQlzxyASe/TfF/Truc/9iPSlSdKil5ewU2lLaKMjf9n/ZREyTNa5w
lLTnHD0HwHuQXG0MKIODQdX04NLHoA+EO4us2/BOw0gHsGgpVCdN1IxDMM8ly91ltcvW//4rVRCf
4F76juX3XjxFYeIOr/GUHLXxrPKPpg3zhYwzUiAFl9hjaqexfEuZ1t00Z+KZ4JEnHAN4KAGHQl2O
mf7mG2/i9ajOe5WJlAFm9px+hrAJ64+QMSFbtHMjTYs3aXt//D46IfF6D+y2V8cKhUNP7t2LUPMY
thRLlOEOFUOmr24hDT9T2q8UtwBhTlvXdySIW1IQMrXOMlyPotWcrWQg2jabF340PCD6wKwfOQvW
ma4ELdOqyDC2gC76cr/i+9InLyt1cXigZGPyEQvEDgKtxuIfolc+E7lsE0Z0s2J+PGy12TWn44bi
YgBFh8qQONY9qDUTOh1cqP+F+brDKcATBHSpDog3wrccJHh9RYbx2KoYzImtyRdamDCnAJavXgDE
eKu/R9XTZQgRcpvS11QhdFUpPB+xmsVQ7kswhRSUx06Vtwu8qou2IlYa34fBQ4DuC2MQcqXb60o/
5wpOYX3T0PiuKgjtfX8BUOl1cIqniMNfG59qHUCim9wfpG9l+J17Yh8PHYs+uW9Fx2MO7aIoX91g
QY56dXgAAx8EerHqiQhio06hYrZd2bv0wbCViH+ToIzctsV5+7NPZMenCbF3DQeYx8agJlQmzTJZ
evo+K9ZvMq3RA15nCLTDDU0/lFBltpyPomqV9wwB6f7xnTdY2xFsu+ZtVl9S5Bkk9ih1rAGSaW64
/TDvSFk1YIYWoOCxJ79ulG+NyEox6eU1hkamzzxlhcYwqyRJoGr6N1UJR6JYQDEloXEl9/Q7iVaE
pTs9w/MbHNjICdHrtzNtSu/9SScLC0uvy6qLbQcTd5qDfAzHrK25qve4aoEznKwjdtyxICalJmfx
HHlb2QJe316Ee2bcujk41BR6BbGJhdmZlBhxHqT3kj65v2dz1m9ua4T9EEWfXGqcYGOHUfXuG3jc
V/WcL20R4dayquCG8pkKoB81wOXQOp8m0pNnnyWJCgc7WQEEFrfjOpXQnisafMJAhSznjaoF4rHS
HBy1x/+Fm/1bFOupI6kmsul/3WVAdiC3Tc2+3jovmsvYwe/bad5Y4ve/y94bLU7FcXW7Gma9Uau3
b26lS39thBh6lBf8QtQMovMczXx82acOl3cgt4saqAE+wKfmyv14cwKa9RbdOs8gCW0L1fa/e5SG
MXzVVNrNyd/f+CTQTL/gfskPPHOoyL+toZtiOPNiLUgKd4NeiNB8+C3W3b0SeHVV2fyk2B/FqRSX
lXlwrL432q/prQCcHLT2CF64HnmBpEER0+EMAm3apMZHOVl5T/27zhxCfjDX3VlhZJj974yhvmwf
CGnKcGRNvWZIYbsPMpauQZFEPYFVcjj281eERWjsVQv0j6NWKAKifsdeuvr/ENq1/EOwZKUAXeil
TLcdZuFdG6LTeSnwwrUv6HkP4g7pq8SPd9fIsyXjsG+WV3P7lLKfJb1/+U/IdY+ZQCHmPwEFwYrO
Q+tqVmIC6U658f80SsTZeElQz8hUbwILAymbOfYD4fG9GGHAqMn7llTPJRyhbZclUuPlsJTDZVq4
1VqZCOqL4yoIXY6GV16P2sZa4+MkyYr4vgWy+K49nnhzlSk44vxEqM0h191whs+IwQ3f5xiI0twH
3i67YLmU41EfNDX2XppwKlaTLSDPWmyrtiTk1/pKBKfXyInE4XPqdeRG4MO/2tm9PkOPiSV75yC0
2T1Rx7z0if+xO7mh/Uzyb3D39gb1oEyoEniB0q7A9bDFRgGescKmTKR4WEwvgG9DHZdcCI+lWe5S
Ynr9auJ6DA42gfWn4kH50U0RMrVXav6xf4jSZZysHejeurLuvHitAqSPC6ttaWdqicHnat93RTtE
2hBv+cE9vF72lADC3pfiNc2cz1dcb9pMWWZ4nv6gPUFaW0TJeX4tJ82pX8AIBsxVy2HrVkqP+eg9
kAxDA1/xfwcrgpJ8g8uVRKd+7Om37O/PsgBH7eTBc0zY759Q+IE10uwsJ2cGauivuwEleBhA/y5b
TJUyYEXBqRWJh6yzx7ktL9NbmzSDmEyB/A57L90PJ2+XiEaHy0bcNgINGAy8Dtixi5gvgxAnwlIp
vYRbaC56d/wdUcsB3AyA9FmnkzCWtwBqcJDgfqbQWtxY9wiwzxChbwBTHsS/r1HrTxpk0YTTjcjg
Xbfp2TV7hlirC2gdjo+cMbKP8pKR2w0rMV7oReBmM4aeCzm44bmjxmXpfljsAGttVWkPL4jet83V
QmZM585QA2PMwGehrSM6/yWGcupJx0pkED+0UUQF81Xq14xPHiJ73BUbWtjRdZNR1xNJ3P8EGnmm
LYlOYavsbrdMWmJ0+Pt2Pcsl66X+SYdQS9OOqL9Ekbn9NTsLp1lQHhnQTnPMAmXZOOlVjjmWDJpn
AFxpBW1AvcWITDSuJ35tsJ2227s46pOaJ+pogBvWW7ZMxEbRcqDe8HsZBHi6ng3fgE/Ev4ITZ69Q
3bIqt7BbWdM0RdzwJlU207rNqIwkZa4OUDoDJSvYvhHRs1Kvtt3lvEL8vtRivkNxZ4IbBKxGanYd
bfzJwAPQToYkEllIGbMeQb4aU394hhCxWkrbtAe5qyYtXmKo9ppljC/qb7yczl7WZmzq9IdtzIvm
WMDOT1V7oTL6lBTnaYZjvohpeFKsL4OIO7XsMBRR2Ysgo4gYQrfAavn63kZdifwX0bRwxdUTfu6p
nyv9oPZC8FBUrp5woGa8Z019OFYm+TVJZ0tVclAkyKgJKrifw77R9Lx7tX3NOv/yxn9X5It91lT5
6rDIOwq4JCZ3HdrP8qJdUtnWwo6/8q/tMUeKjZq/sanV3L5+97ktMYtXI2CTfrmbYgG0fuypGo4y
mKgEbuAz6dAlo1RekEmV0m8MmJhfMZsrIxfRCYqxW3/WlO9N7DPR9zWHnrqCX8FzjZi//8MrMVvv
JfxT058ZAJ/fN/Vl+Em/x0yB6FLOY4d411NBejfW/myvrRPFJ/85b2rq2Q6IjpNn2QwjoLmDEPAu
lem2SAIjEzP0YKXz9RaZb1X84xUwgQ8qoECkHkjfQi7wvwnv7a/oeClAPHJCMcUneEsCEC+bvYwj
vvvp7egnTzU/KEyDg7zp98STLmZTGmvPzuwOENYlNnlOF8qq18Mc0maTodaAty/+f0a5z4EhvOej
IGEMTUlGLL3e8jh8+Cda+gdhVprecj7Hjy2kfoqt/tRBD4W3F6gdMsDYk7NlliAImZRXIJC8Iuds
dh8hYOHIyPZXwHdtH6RNhhoPpZguSRlBycvsBJNWcVlXJi9nZBOm9f2xDxfEA5e1ZVi2KWiRWdBu
p3jXhQSFQquJAmjpwZkXNjP5/AoDq5lDRa1fI7y+zL52VhCEiVVZsXc+P3BW/+MLTGXLVmf8YNGV
UZEZCfRKZeAhITo3S56j9fqKlykC7Jfw4c99MzfcaUCKTjTWMJJdZ7FCibJKPyvHQnQaMu9Ja1eL
MHyF3SyvRSl7XeisNW2PZ2S6INq4uktrm+987SV5nipaUh2yytYcINBXvpyq1+dok9QfViouQYtJ
1XXmn54KrY+8KmuXSELd3OSTsmlGQMa3rLeXkV/1WD6dWTAXogXF4ZGnu/H7fuxc4Ifp26RoD61N
8QiGOqLalQeEgYLCjYK19CZgnjbfNarzhLDuUQR7w6p6korrhDD5mYDyy17Apjl1+zrf4Ad32gPc
P47Y1V5HISYM8dfY2OhCRZ4I+1/PbibdwCn8QhYgriX2mIO0Kc0KH3rblk/ax2OsRCPRzoZJvffu
qz27aWZgizGD1J4jWY7LFln93kQk6QyLtHiERaeSaB5HmUlkOnh8DkWa8Vd+RzSZCruTvJU+ucvO
az3IHKsscQCnh9O+9f9aWB+gPayiVgGE2MnwAaW2a/3olmb3q+D1u4mFbX+Ikx2AcXMw+6+NY79r
pLzaHwjSo0vrXzzUhX8tsownWjKqEbslBCTfcdm5QK3eWeZR8CpPZZFbdgAcyVKEKnjyGm1E91tR
yfnDWOx7ZF7q9iZNhI34GFl2p3K1AgEgE73zjzIuQan/OPoqrUq9XPqXx7aTQ/XpM07oprMkqfqX
rRckE/rmSmMjCtlGjQuwH1D5M/5ZVGkbdryaQaglS5ctnK1CQ5cgARNdia//wXcnrKD3HjPYO0oE
Js3AvVh5R9TP/o/+o2wQNbfjnNfNT3m/bQtt+rx0OIylCrikYlGnylYXVY6dkfjWAyRp59vfiHOw
IY/PjH9TeqkapBaiCC8y/XdWnl5PFZyNPmc+XK/SaI7GgbRCrCcDrolroJ7Vf5zDeWk50UprXIKj
dnZBjau2kPmKtTx6ppRRhejzM3R/2xIAdphU02uDIldROH5LnSWHP635XHkeoyU/K7nvpIWNQzYS
xILT/+i0eF24cV4GiYtAU9vH1KQZDAeW4jf2Fs914wqkQka5Vhsxu3I6uCohWxyi43Rp3NAfGknk
xS3fDa1h1vuKk5VwuxlpR15s2mt7DVFOpPMdWtdM6557oE4aPpa2qO7V2epfJ043gmBojkSM7FHI
kMqKMZ3A89f8wjOa9hnY9lT6EekZqyJsZz/n7iXXVq1lPXIg0XdVavMBtwx6S3Ubw0YryZIo6s63
8eBpARNxWv6ZBsn3++BMqIjIb3vs6oUBd5lJydOs4SeukiWgGWt1hsOMazBTE2DgZqvD+oDw8bNu
AKqIhrdmisHSdBl51xbT9vo4KX89f2eX7WfW6WLytl+KCs0uyCwibpJm+KW+N49+hl8CtqfK6iiC
GiWXKo+J6kduI9AgaAJZQ/Wj5EIWgj3s0ERzW2oam4/FrvHO7Jw1J8yfv15RVnZxnz1c+YVJVSdd
kvWhLT98g+i1Qp+G8LNyP1ZfdNaFBh4kVzLYsLKTMC3yrKz8pbi8b+TdMTAmHIUtLVfdaS4/IMbE
qgv0PZ2mDwwr+axJHYJIhZwwQT4ihQ7ggYfFuRsBXAikP8LZGvs/RGpj5ati7CL/CsBkSAscHKwP
OTHdQAweN4Tf33VtPzCcDanS95TDZODxCkySYmPYZkiTbCBAPVoqk/tGd1/2m/hYm8R8SbcEy6Pb
/C2GWN03ezqF4i00TPblQOZNEp0/i91E+G4zIELQak5KqFWNoWHkEed+9zq9K36cqeRIMBGvsj/t
c+87dtT1HsHvqRdOm4n7xQLD9anO1ECJLKwjwFe/lJBaL8D/tGW1vTU6AP76u6Q4TeEj68kVxClB
UGuStChlbEVVVjR1DVF9XFRJgRjJMdIdljW4F9B+Bx3TJMR2PEzwk55FTU6MClMfo8TtE/HLcm9l
lAv+5pzCCV5F9PoqFnZ8TzVQ8/SN29JRqwU99H/wp5T+RnHq61w1k8sZfb50vghCCh9dJTHwvGtK
OPSnqDg5AWe7P0xuSI3bKmaz44J1/CkAh7xJr3u1UtE3o2RMRn1y2+4Q1y2A7fZZdWq6XVtu4D04
w1ITfrkn9PvJlimvINFusqM3vbaZ0oc41PuhvFX74oZkIjHNL6m/zSBEH2743UOJ9FSiIHherwG3
JbgeUkIvL/P3AarYFinkD6ku6h2L2bp2qVKTuc6AsMvZI2GpI+a7lUB7qLOJABCobhkwUPTSYNsQ
8TTF/UpCcH0WYPcPwACAYiAuWTIB5Y76Xx8i3Zc3BaQRE5LVs/NGSpkSVoji8FniGx0BcEWyKnNt
xufTHsaV4fmQtuukL+9r0TcLQzQfjYZ8s9er+TKB1bjXGC2FeFwyNeoqJNiA5ikhKf4N+FHos6MS
lFbdthw6y5Zorcrqe/TREgZ8pDMGVYE2oinzFVR6E+93pSGOWaNGhdCT9uqv+gkUBJMqKXFMUJjo
SeDEnotaguDu/iwY+UWih3p+exPpSBWW0LN6GCYQzmkeK9fgDi683H2xL7+eNJut6M01jZ4x1A0E
s20PmDA9LqMrVogYZZfYTvxUnT6HVSa3xPxbZ+QWuSc5gd7eKA/qMCoWmv2LRX+PCZv9v5hOwWFw
DcstU3qdM/Jz/yewwSQYICoOuyVHitj4wFRfuuVYFvRRiZMre1mglDF3vQQo2G3+jsn6cdayXq+v
nSfcv7ID8AoSBlQ9OBbxc0fX96l/DmpSH5x2Vwj2J9Fa2LWN3rY4duoTTexUAAcGbc3UQneBcA1t
sAPNJk5Y49gS6HtaComcA1vn5cxf8tlftWwMMXxI6tH4IjXgKbMTvdcPd1o8KpxAOGht28jMylxB
5Pwf5+m6nOyEkvZbJ91gbe6lSQ4caifr1W+LhITMl4GtdZoRhaCRCaOZ7ykvSMmJtU/GUZ0O4ruV
LwbCRuP+k8NWPi9UCX/jSKn8e3qM0V5MSiFQSilc8wJsgkbsixLd6v/GIBDGWAtZ9pKXU+N90oCa
jvK+OvED46/iDopqi3ezwluY8JLmsWScQeEnxTWs0MquWSVd+DUeT6hXbW/qEpumTGUtCNkJUVzA
1ZjLc36z+pILZnrs2ZSA8hOkAYaj52AN5p7eFn2qR5Z3OjyXcrCFJqcNWrGcfRUVOcuID5pKUn1p
2sssVduxQulz51FEYQOkUlWLsM3UJpE5F8tvg5uTuPagxrF0Ea5MxQDbcvb4qHEujT5tHXm+f45D
fyktWewCmbp3IhBsINRySZCvgAHTBFNEfhwVwpc2M5r1DucB8oAO+3CS64BpONR1uqYuH0gZUOd1
4uDDrd/c9bsAn86LeJCDSIiwAZXxQ+kS+FCaajqQV2HlYVo61kpPAFWsGvdEKzpl3gTIJUHYhvVK
a8ngrcMdfTbIuWdqGHhnEXLBvg42QQFwaXQdqWH49nl2j3d7i4C226ns3sue55hq7/25Y4h84hQN
iugJiRwIdYueFZvvIZkTMxBGnVJIb7daWGLn1RaXBMPiS8eFr4qpH/EvMfNxlW7xYvfQnS9OUniE
v9Eefcj+C1sXUpF88zyJPeKoE4SPHYM9ME/w/5M9BEJIZ5mcwVyUCtdArcb1fTgbB+ENxOensLPt
wNNRbMm8ReImiBlZSZJLA/zVzTBk3OPpucYtbINExjMJJPQvf/AljcTSl0xHirgAO2aaEGEUznPO
/kpFxZ0KDZ8zgX2wQw5GnKYDAwyMrYu8DwLedsjPBJlqRrlCeqwJxtVuVYCFvuMlZSEsz22xMYxd
MlFvnI3uqiZZGXeFVu3ko6FbUtcSxU7HR3A4Y6zeAti9XvQ7GwwPmCwvM5bHK/xJ1xvFmMAtdOeL
tI3W/PE9v88C8IBlCEB9eys4T1wZ+kH0mqAVlG9Ifs84EdOyXbBg1dPFHpREHM9WQZenZP6uACEf
megPFypv50Hl25ljQff9Gh+d+i4I1yJU4DRHtTJenGRkOiSxNFNRHpO99CcZIjTixiURiDesty57
wLfE/aEUcTnUFed9uznP3ZDqxX9sRzCkzkUwbllCkx6a2dMLrKZ0AfNOdapwwOKdnNLO5QyIWAuZ
4kT3fCvxxmt3/PWPj0jvCJOHFis0SGz99fUpzHUGh+RfX5bpo2yVmUIlyguBUrJ6SopYiuNBvyPn
ppsYm/NGgQiIGhjSnp/khsrI63AgYNpJ/apKtS0k6doYoY0sdiQxi7wIBZbTRbtHs+UmeoxNIsds
AZsEVprcTrMiklPZ5dFaAkp0ErdmKADGGrjhPL5tqpJYHshxY9eMDqTnRVGiA3SCo76qc57WcFFS
T88PwwJk54xAkWSZ+Z2ar2LNetWEk9vYC5nD//aSpifm4ZuP8r4M8E19Az0U3bvDATaP9G/02CQv
+o/0I69PZsNQaDvTuMQS7yVnznuxEf3gDZcJerNki5sQSvpmRouapdS3FKqAHIA6S6D/oqxys+Un
FihFBF6SNsXcgrbA3PfF1Hp2Ha4cYJJa/UcjY/GmdJO5v/qh8fYuSP9rInfcoEN8Dx51FsCt/Te6
K0gyK38H/D//2jvSg3CNOTlVvBPHzpi3J+7XG/SEKRfpt1qgwo7iqnFGn8gDNttkmMNYMrY2egbJ
rqoUa9brrNq7GCDEjTbViKTnE8bAAMreGhQ1H3zt2pvlBrqILxXVkyqcJXlnE923XzzpO+tH6Z5t
rGImtM42uH0fn/GK2WBp9YGXgm6MxQzNfQWmLgxZdo3YRa6qGIEwbJoS5PAcSAS2KkJPFl7TtBzh
EzzEi0HFWFv/d9YKDZRncwged4K6+q4oPy/S6xKR6xBfmPzBLfhk9L5pmKvGGSAAvc3zJgq9a8JU
hzYi9pzwLWqOyNqWqMbUFqmj/OyEVnSn1kCc5jDFBwVrtKKy1MEznYf9kLAPnPelB6NIz+htrXRU
JWeKil/m5dZwN7ozM5/tHy2k74MiJXKz4FnNUo9F3nrSFMFojhNAlugUpIOQ43Tr4wByR6GUDW4Z
/BBKtFgntrsGG7EQ8fK5Dt/eC0NxZKy/2+G32jy7yCnlnq4orbRi/vvfH6jLToJxAA58x5jj+Nv/
axcymV/Uhcbec5nNL0S1G0plKYEnKFONwJUMGxybpkSKjs4AgwJ0JwUvAtjD9d5S5xorn1tEk0cL
iKOeZAKQPlsBxCslYmha1/JEjoj/tjpr18ntneuvxjEAtlO3kwBtK45yvj90iKfM5AvfDMx0YXZl
Nu6BfkQ47KJOHbhbnx0tB4m2b/OKcKiZqfcRsp2LDbiK4Z9ay/ZNGZ2UU01xdB3rpfOkfmvftRgL
3bZiHbTL+9VIUTv5KwyTi2VRyXtmfvIigyN3kEI6B8bXoTZEErHVpv9q9MwPXNrfxne7V4AfmZvc
6PtaZvhpTo1K1MXtgQ9KNDoIbDjXUTc0+OBys0qkYGWvWUlugCJPRmqSZa9wegqQSzK0GN48vWy+
ZRGpJ3D+R9F+d5aG/DlpEpOibVCiCpDabEucKXL0BD5G2Q0v3ydQzY7Cf/2F1UfSeTj9t2zAAPOZ
amtnUIehUAZafMmeJXnTKttvqqAQi1REwrCxg45N3mcRWG9gTmVLbiZwYq9HD+Iq28Ukwjs0vzSW
5regRBfyn6U3yCYnzmQb/fpPYBu2Q8Xg4iDkSfSa4AVd4fGodPS26gTuYvj+3rGpaAH5A+JUscLe
dv2dX0DdopNjjVFo/gr+KCfiFaTUVfddiJ9bwgj4vET80HmDr6ihQI81XItVOYhVAqQSrQ1Y5xPr
vmJmvwpzix5zR/D8kHHCYecmbXo6cm6Gsbvk0eKG5911FKqo7Sr3lQO2/xeka6OataJ6MXIr6DSd
/3fhCVKrSfCYusB98a03uNAcae4TJXB1DyNsQEXqtdSdxB1A3wdEjdsI7tlniRdCTpaNEUQLvS3C
0DKBqdUD6WDrPR5Xz2KTvlvADTuEQvp3g6qipzXSk8OzvTzo3gbSyFV3v2gs0U9XTNJ01q+PYLeK
hbbesBBCMR0L+tC8/u9/75sq9J1xcUk9A6FCi1uw/oOwZ3NttNJYgautT8eFCHAfobz3t2cwOsQK
NW8qq0ICCtjLE/84xz7fLUEMJKR/N/EK0WHXfCiyXN0ZPWMb5i/s6iFCoaOEqEah4kcm0ywxzELn
3wiaeA3cXnWewhlLikJ6+sDzIJ7j8RMJ3DqDBdGpzjMk7UtKCP2R24MiX6dVIg58ML+HJknQ9b6R
4YZlhRQ7Yb5UeqM/3lwafgqtZroToIkPWoEakUSwL6Z0hBEJgX4sNDGzW/gVhJ2sqF0zmGmmdhPv
N6JBwVZAqW06wuuEgPPOVWWSO7GmOLXgG+b12c8OoWvV/1l9XLI6d//5CL62RbsVg7YKJtwZ0+1z
6quAL2ug7VUE/gU0n9RGaTpRJO4j8fVtNjsbkoF6QlP3xsWGH/4Ssc5wvG/MNrKn5V+of73wtm6O
rDSsHXMh4dOvvcqd6YjfOkNjgK/e58AwVWCHyrOCzLpvdmYrUja3Enf9UfDhTYs2xmmsn9EVaRXb
C8gbXhotcw5tZV84yul/UQm0yLwuUjxO7WB7j9cFIrqH/K69q5mpU1pdgPc6b++qrclu1FrXK2AF
TPUAnF2hkAY7SvV0L4dJbcoWD5uo5KlhkCQT/A0YHQIdINFt6OPL/WHDOg+tBYlPuUFzSNQf1q6F
oOJWrgxnqQolrLd0VPyZzOs015xj3MpKD1KEkEifkCFvuUTFPMuOIWLdKHFvutP5KdJTrLWGgo4y
q9Da3gtjltN0PKLCb+CavCG8fCRK8gK8elNbevcju7i9nnD7BjPMRXu3ED6gCrgpH5sVFdbiks5a
YGr/pDeCSnsNgXPFSg41zyiExMzd4+32WIARgZFlThkyLAZ0PEOJFpZHbtD2kiHxhxAup++Az9F1
Z8kPZhBuhBvTt1j93rCKNkS0yQKQ/jqKz6arI55JfmYccUIdGyRTY6Sb4kdKk+AB+wQBmmEvF0uE
qlzAeCoWdmCaZHeCBd/9D+h1DDsU2iVaiNajBXD3/LY/dwEp5Q16V8P5Pr4mxFdP8N2nWI+/j32E
HYsSO4HBvTuk+9xCgXzzMNy/M5+vAfnclACJQ2XVunJWFwH0o8R958cb5MZ0fgAWi5AyKz96hBJB
fI9qFwPpcf7BLe4OEArqV6iXPNqDYd3j++zZaeXX16rQrkeDgB5+B/l3CdBaHyHd5qkIjedl0s7h
x3Lho8w8A68qlf4YsnrShlkCdsIS3uBvzQLBnLBwKhOPXFTUUsXxSKAri6eskY5aBsPVYSaDwMqI
4V5O3J/mFx0bymbd8TzaYtCa3DyeJQDzHkTDDZ2jD2f6TtBqQ7DVYUsbM4WAahHHgrfPLe3XUYmC
MmsgkoqcZkrFJXonGqSyKsStVPWLAEhCMdHtpidvNGHOMtws2kARWgvJEkSw8eKoAZPTFWJKYqaz
Qs2ALvgeQ+Md8WKZ4RvxM1eArzaMLTk5EDw75XcyWrE/VSqXO1plJuPw+xPYO+Y+Z1jHo256seBa
1fhBs6lXsOZNGR9YT6ZHox7OSQxygoODaRONJnAC4lEA5LT7TyT01E4vx58Vhr0GjfsNYx/8YRhb
3YEfq8zGa0vkNl+/1ffkMKY+O9Nm8KEqo5oXODlB6dOoowEsVVydeA2QtTY+uZGxEYlGDwXT4/3C
mYKSklISf/DcpyD5rEQ0UHnwurt7Vr4G6+mJJhhs1I8whvK5du7sRkFUhbleg/EZ9xUCwUODIpjP
2nSha5whjaTdVi+d5JHs1HTqZePlz+gfktvPwTlT9O5e0J2oDsfk5Xya3UpG/WeKW5DIXEHwLUeU
Mqimg8R8G2cjbFPtefCyQKsFt09Z08Mg9Jc2mPebWXBYm/hXYyADnJKzB03virpl0ivVvf5XMOve
Yij6JJj47fD9uPmZ6caZ1bHz/0GOv3C/psaRyYPfkekvRfNHWBTglrvw0eZSWBF0ZS1f7cfqEAtu
w4Pon8y1dy+q+AOzHZ92yMTxWNfiNdXvwixK2Jv3PyIjSksU8jd8Q2xQCEET5UlihEU80cOn9oRi
W0yXfz1MhCuaYIzP6BI9Mypzg3yOl634/RZcY79D1ibJAeQ1KYqv8gwiRJBBXP4QlwE6wm50yKd0
nwkc9Xore2I8w5LJ/n+y33YxQn+zYiui6dgZU1Y7tY8AyYXZTg75X3SfGUUFLFJOfX+MtfYDkoGt
wd8c66F82Mg2WlObIy2aoeZYHcjq/boYUvVVQjlI6e13s//pDDfkFLklpD6+x2cVqw3dWhejmTFi
hJ/N5JCj5vp+aRV4VrYsn6tf+gFM5laDzG3KelFhxft0ifdiMuQ7EbJWYoaYuJHLEa0MmD/2h62L
M1WEhjskvYFrj54XHxbNB37JF5GvWhbuWSMI/kbE/oM3x9ccwvMVrmLLHfqx60AL9HmLYffrnM4j
GHkhgmoD0PneKxsYErOM1BSR7oPd1MK4B/jyMM+t+Pq5PhdIIssalvvOz8pY+UCQeFQL+IuNnxwX
x1W0zSCGoTcb8ulMaCpfe8kWx0/QDuzgrR37PV69jnIEB6S6eIf9ZapmHD/DKo6I+zoX9suRkd3A
FwnKN77eZB598utlFoQOYxmx8XZfkFJC1o7iOHyCPOdjcBVHJ6jMURZ0vLcU6ixh5c7uBtqZaFdJ
4rNRXk+BZOghec5eBHy08FNFffwmVFbEYv0Lsa7n0xaPVkadzNArM8Hr/AiZogUHP6fx87r51o4w
+Z9V7k/p72otdQTmSY4HgOnYBCM69zXc8StYSnzgFdJiIWHI4gRelUuKFT++8csOsLSd5HDVUq1R
hSgytD4XHFrT8rcsWTtrsWGMKob5KUWi88XaxyBuv8Z7hPo6akUpZALG1PiTL/gz4tf34wXYiMtO
mp/HyYEwtV6CTlH22vOKBmshAGVwphJsgmpP+JdTPsYDvcDkgQcwfEw5NBNJgb/HIlySDM714p/G
h5vuacPoPXjwJODvdkwgpw9b2LMIIXSvC+k2pyy30Ab9KXR2VFhH1oIwYJwxfff6fcv+zmfim7We
QJEeDKetExjsFT+LUY/9AG8gYMy4fxY3yVlm7UuOnCmJgljaQoo+ZnVwOBKp+IPlFHDMJSaAN/iP
mNQv4qcMEDDNG2JZquZgTVjSUryq/kFhEx5ga86gzYPH7/aonXHVkkpsiwtPYyYkIA53QUbT/Y//
Hi9Dxx/nqkRIFF+ItKWd69dEfOtJ3Rgd8lo3iuwPici4Ft960f97X+AyiqWadgyMSIq2KPDnCa0P
r1KPsqkmbB0jTto2De3fHUa8WUEMg/SjMHO9yI0smStazADHxSx+RFTIHTd7d+oi3aI0fdbEfdZ9
87zuJ9ztzAX2K4O9rLymQGprnbzpJrRNXQB+ria9/IWpTTAz9d2KnAldXywsKAHyLsZdPbCUldzR
R8/6CNOW90B6VefZsa1dbK1QhOMbMUCoc0ylKfVLjlzWjWteZrhZBp7T55uXqZsgnGZl3vzEvNas
s6cGv0qthcneIvPwy3FN0UBTUuGkeNr07d/GNcdbziu2c4T6k1QHHBqYeve7dgzoID4enRFbJ4iP
7nMyUAdEUaxieAx5mShoJZFb/aX6Q9Dp44fAWSHdU94NR6tADE1ZFiCqCA33EN7b9xmbBCBaqu9J
U7dbY5B841IMgeOaJ9k3n7n8OC0Y3VCRu8cELGcAiGwNwZsx2sLpECfvpBR4uBMv6WxqDxVcOln8
n1INeAQ0E0rm7f9Vg9J9lWUouj4pnLG5Eka0FW+uY3s07Tp66zucGO5o5x3YRhDmiX9TLwtTP6KD
IZGST2/0I9fzZ9pUvnem1nsVP0KcarjznFUfLXEI/ujEYGZbUNK7NhzkoubXP3J0QDemYQJJzQw7
dXGGIm6NV71xO72fK5RFQO3yY4+BB48ijgvPr/qTpvtwHWZmftLqRSCcNkM3jY8pvHjiLSeErrjb
j0SmGUujfeoX+ZJHHfy2GcYdqDTnyyfRGQ0l22BZgLrRyS//p7Ur3BkSkrD/GCPod28fHR9TJn5d
YtAxA596ADj2dvjFtKrixF0nDONIHJ/cV2vIsmOmBE4j9lBbrfK/XjlWWBPEh54z2YNgB36QphTW
SZIp9FltMAMcl//Tc7VyYFbRosOGIDHIFmLSMD3dPWVybgNcWC6dYHgTx1OUVUlIarR6SPWKmK7g
lfUVTqP45evIEtjgMk1MjaxOTjmY4ixk795PIt+NsxrG8myWZk26d+9dcmsEcaFKBL0mhIANoXHf
x+GQhXvszGxWd/pxfP3Lp6Sf/Yf2WzfKPROSxKDgjsREiE4V96gEWqmUQWMYCKWrr130n7e30jb0
F14BPufZA9WnPFXZRjcvIz5Z1rH8p3TXdjSjtjM8rpuY6Q+ocmhc/WJDaYjRtaT7zHbooCpUxC2S
VWV6chpSDwAs8jNTq+y06ZtyhmOibsUXiMdhtnXhqQzk+qM1YwApcbS00IDodhauohzLbA9P2qV/
iTN9QVhMeg8JedmpRDSaGEPGWYwpyXJgGZmuHsR8DiiYu8aAYLcjizXmrrX6/Tphakq/wAFT8vLv
CY4BtwKh/GPrftoeeihVLJnfmiCsDL9C8U4K5pb4rzBlrmMf+U3pvVmSb7Sh5i8g6A51Vwup2bhE
mwpsy2CJC+1+YR3WKvy/2UMztfu40RcBgwhc7lMtURbc9uHRXBqqTuq08FsaJmOQ0BKgzWu2oixz
PFwRc5ghqLydRHUQf2gawJtwf15xG686SnBT1VlbztZoCZvEu4Hp+ojYq44RWNG1MGY7jQ2bketR
kpRVmCY0DkC3DLU5/ZpeKeoxunB904c9bF+00vFaAzUOPt90AlrmPOzZcj8CfEIdYy2yhnMWp4gS
dj0cCpnFhcCRGXrej7Rle5f04dy/Tv/OCq/j/F6R/34BM9UfzAsY4YZK0aC8PbpMSPRWXYHqubmK
eV+G+mtXLZ5fHyaHX0LHevLazfKzPKJSvcd/mgSvQnpkwEIBEW37PFOmvM2COWD1bHRBXAvBtG7C
dvEbn+0HTS1KhVXqu8okMvXXC8WTkMfLSls0AcB8ZbVVwuleef4qzCkKfaLmgc/h3fgl8yhuyoS+
v0P8pNjZfSQW3RwX6PzeKFgAxIlO8mNbOCRsz4MNUZF5SDNv3vzz/bRddwKuAtEw7evhe9POrpyI
5uIoQWmYjyBkG9q13zxmYMp3wHUdPh3FUsC4hl577qGp3tdlXgkpk+egLUmNNb2VfO4YT8xU9n8p
BoYkmgg/CWwwKuXU8eXH+AhJF863E4TXHMXUVhqq6WMbyash0ZU07aUPHBMId+usEaPauOeq/Mm8
+5Yv1Bc87SAY676yheQRjKxpPR6KORO+mBzYSplWJ9H3M6c7ETveXs2Y6xvJrMfE42VOkQX0FG9W
OH2mBQpc/OvpZDGTOc5gQ0dCx5R7p7Yz/gpF7uVQw7qF4i/JiYSRTwvO3OEJWMK36RFdbaWXdAF/
pWbCf57URL17z/pHELT284IF+Z996tSmvY0g66ae+ueD/8SrNzmwir4fMMtSNhvc2gR0PMKXXQ4d
TNeAH9Mb2pnPT0QgQYX1Z7sHeLSUAzwTAlUqYfAT958PRExwUy273VPRLidyDFYF2e8JuwRrSjRD
hvCewjDv9j4zsW2Uisir06Ldvrwgo0LU6u540mNWer6AC/iZGTjXlO2HGrYLG/Gho5xkDJXumRYw
1898L5Ud2IWfAqa+HmaovcPTk5Yv7tqHMUf/2de2hEXP/RBidvmpI18tfrBacZEMxVpZpMv8vM0G
7RDRoDtWbamnP5hRj8bPtDjW1mAJvmIW9Ym/e+/HAQUInmUpZAw6LVjIOLA9RL41gYk4hj7R7pzT
IQ2tiLtFt9biBX1curzNKLfs2nhLwrlroAIYjCYC+oXERJaWn0Il0Kbp6hp9SRx7mm55X8+xFZHc
F/ArTF/ZeAW7kQBVvOooAAYz4TVxsZvC+Th5UHvdcWyrUr7BO+9OZqFs8wUUmlWgi8exxw0zdw1d
TpRJO2gvJPo3LPIagpvcusrSO5OprjflWdUIiDxu0YepuJ5BJrjMmPOeWFicLizPDSmY53Z3nV5m
tgvv9eLKTzHooO4LWswo1dkU2HzyXqzflXDYs9l31tyuUiHwS0BCaBJXyKp8LzZiMzNXeQlfVySa
1ECo9qGk0DUZ7mBlukNKfyYpvLJZpatABDA4Rk2GDCO8HhAlM0/OZyVdHFP2YS7oGhzcAW/bwCdc
Jx51vG4CIYDI78dFiBVxCnOsmLfFEaFMoAeSIo7Q7soIw/fU84EwN+sGpTKpevQMZAN7rsq+4Ezo
p60+bDl+IOEqjia4772KWW3IqUIVQO6p14i3i1XWEtzNrb3rRRorUSiPV8ZSV0TuPTjDBNFiZPEs
uw3Ac8vGY1/OAfno5d0sDcdRbOM5MXn0vsB3UhpybJxJ9FVHeNUcwpHC+mQG6bBhigeqWjCPkYbn
LyAKNc80hnRtvIsjPlWdPdcfTQ6MWGdqvUpx2NWgruXRn+NAocUOAjsSsI8uFNDFCBzZUtbIiTb7
b/hbwVtVXdx2dkSvtjGb+zO2wG3D9ch30ZXE8/3kUL7BnALcZRJYnHgbkHUho+g7PqId6t0CztFQ
ixSxJE+Ql86CeCTUrHkC/rncSUO/ninHdhctGvdhYTbnVObi92oZRUxwLLgbDVumdHuZX6gl4GfY
kr22POwPL8yd5eSCeH6otNCw3TYcG+Zz+99ODMmreDzDeUEWdPRTd97gqJs9HhQF+yljUpjbqpLr
bcbCLf3LJ0tXJzRDnIoZS0fZP9EO2hOCDKnDvU8+OzD0n3wcerqaMsDD+SS9467XO8JuhQASQoAs
jeGwZAGNsmd9Uc69lvEJSW1b385jEnneLX17DZALu/ydgzZ+EldevI9QyXNSQlRdho4vMB3jd6QI
ZVSfioFY4gRCy3WAVaiLOWSXsiH08c0Zv+ISUKYS8tc+qtxQkq6ZuvbJJ2Ktf2e7GgGhsMINvJuS
CPE0pm6Dyk+EIZXVNMzohGfN+hjsvOxGKr4+xET5qY7eFThPEoVkYVQBxXb2VU8pMIELWi9bWNY2
WU56NAYBroC5/1GHEM0UwhxfbLUEwmPaO9use1x40NUJxs7EJOZTAwCImPF9DF7AtjEdfFwBJ6dz
NMAEFDnVJ15FcOVZMret+yZZNEV56AGG98wyqWmcS3vPsAF5ofZoCvzmQJW4o1AByKP+e26ycbE0
amwOOsT5g7q9uuNlEIZOYo2efslNvpPupAvEoh+KiL7ZKtWXMeC3S8aEnDppTujOnkN3M8DJhqnI
X2OFJ6zyNn2fnAHY8cAPVrKJtGOt3iNOYWO/86DS69nfgyJUOUpcFT4RW8lqtU+ez9wBxRcTYvY5
TzoazxgKh5dJ8wIWPa3VTMIflKVyESPpxD6rTfU61/eDaup14KxokZ9f0Z7FhxaK/H0STMQHOinZ
AA2QdXLQXQzDF2nttQkvF1oKOZEMvIEFvxNtX89CHXr0hqTVqKma2cOa3YRLB5RFow8L3cLasAvo
WPEdDv/VFkFUrKNMkPcY9y316h+XlGJf5h1zZOh5ceRLJ6TPL2hxjU/duyMcQ3n9339zt7u0r0BR
N6e94WRYX8bOADwCxaSeCnc2rxGADBRtPf9JRsjeCVvi4+TCxiBO5naDzG8J2YAQwEz7DEsvWK2H
3jABbbto5MMie09xXF56wTrNCms4dNu1ROgSt/rYzUiH9aZdlQGCrYY4db1HTXGomvtFWoIidpvn
JGaRrjK5qIH7KKId/uN0ny6rEquMFRkn89wYg+Fdt78Pvi1ihUwnp61HY6ELxC0oEDsABRAHw8n2
D8tPhKBU+cZDSF6QpARn4JktWp2G2qXEetj0odRUKga6l/o31kRxVEodtiQJBl2ThoYdKKkCXTee
WwOR2ghAk67eLgPxck0l/7FzS26UfTHJprshxkcpcrVD1ccjITjyQ0QgVHZGoFHVxBpB8eg9z4s2
2HnLs0D+McsFSkSvThyQFUwRRqzoY0zTKaBv3hfIEYMZNMx3hC7zOFWcHNrue6wg/zW8Jx5OM/Bt
9qtzpgNlWRl0SVaZ3VW1F3/j6y67jNbCrG6Req9lO0UHtirnETaieANx3jZEwacmClNDDxPcZtJD
gp26yq5JaaaQBluxGE8kkCfCzfh4qLnrSLtb3AKMA2D9tnfa2CBsHRVcD8DZM8Azukkp+IFWLNJ6
+kX5Jshpx8naoZxAU8vB1OKs+6BsrVYssXJ4oAXbgKclqZ7pr/lgOKnZgMdJgvulv0jSSU9kt8io
Nk/a/EgsI+d7IfRQpuwvpIr+eh6rV2+rm44UIcKHJ10Ne+fMSqwjcU/QgUBqnUhYvLfvasBlsDFt
ObzdMC6HDoYCLCI2Dko3CnteCZxERaAskVokTA2wsgmsIcEccULwdCNbu4sNqaZW1G6GBrbB6MVN
sAX7CnXPeOV8Q6pgGj03Gl4gp9HlCsL2eoqQH8RveFYuwo9kcbriF0ulnb0qqiiSCAuqfBdQ8r7Y
IuoC02JVhYlifgBUJKcGlXxAaSLVLeezd0zCyZR7hBRi98EGF5sXdPmsSlny4kSx4s2zp9Ev/Sn9
mxosi8JiMUgozbjyeXcvGMM3YnUdlB6/9MzeEGViElzf6D/uJsZxg5G6s4ajaytRHLNaVY+Uv4Gm
R7O5/s+4sEvud+UILENnelgtTcIuJAyEB6DuH9wjyfmeun1K/jmbet+ULjsMg/otDZy7gpNg3Cea
PVfVEl5V/V6SxHRB/k/sCOEfMiv/GtG3SSHkf5ziWB7ENfDp31nyWtYbMOS0asqBAlbWvGkM2AME
tmn2TkSuuduMyXwjdKUnSiaHhCaPkR7AbC8lZD2Peye8544ECfWkhnOuNa5oDYSvg9mclrYGuN/P
MAtLRhHpfe2G+PGnOwH4kRw3IPvsyjoJ41v2HsOJ/EjsLdxCMWg3GvPih/Y19RvQ3TMeZFy/kAk6
bizwS3XQKM8UGK61IP5CWQpqyFqG81DgG0/Gz1iEcOABm65GGihCB62ji3rhRBufcf9AfUos/D+n
MeGCRWmbqBUbEm7esGOraSHa9tKd7KrYDawuNNT0kU3eQHY4162eHdOrvN0ahLGsM3YzQooSSPQz
a+Hl1rzJtu0WRdhmdROt55CslBu4G5Q+08IRRmZTVukF2ghTaKLIih/zMQIufjSFj9aryePw5fwO
6KfAFkvXkFsGppR48VjrV52qLOK0/AvpaPeZxpmPAaMn1pVQfifTRGB8ac1yGA3YR8+h3/s+4zFv
uKLU97SU6mLeaLCcg2plBxrPefHgCPj82y1fTHfgY+rhMsjZkQ5QYGCpzdEvvDskvGfIMZmqjYdo
QiDlsfJuiM04TjHa85hbJsEZDXqryPiwyG3FaFDsekeUTOcF53uN+MXrtSZ9FM7T0FI36/Kj02U3
1KKNuP1usM4n/TOPk107HjsRiU6l2L6R4gfEXUtnz00FZUGpdLS0f+GpW845qFPCz6v+UEgNOvW/
C6AApvSHxPIzuXr5Zju+37MZTRY0gKZ+KgqFyQI+/zRfo6ZgxmlR/V3Y+scs7NxvbuWao4ib+CJT
F5hHO4qaSTgBq8WVwDEDpA7I4x8zey8ngRdXBeibzPayR6CsgS4VdQAhrFWo1Mkbu4a98h32U47u
8Q9cIaEwJd/207N0CB3fxuFJZ56BqEz1gjfxSsm6kK30my1YF3EtQ8Cam+0HcjJRi8Mayu01V0Bm
POKP5pS8YYRbswF95cRUPPtvgFpekr66M+4qxv781aUHJYBkkqZhGQLwBR09jilnZ8RFY9dJPUoB
ijtcaPfS+GQA5Yj364IRiX6BVo/PCOuy3v+wQCFuUIe3XuXXOZaF2+W7476VnGw7zU5bGnDzTQ/j
9cWfM2+9qNF3r2C9OC39Pqxa4hVV5wasGBZwT9HoGr0XCgJxillzb4L9Adpw8xfQaCSkhy6fCtB2
UcziRjrs4A6IwhsoVAXVKJIipi5yojCzSqu9mfh1R0puSb4TwktNYzCLxJEof80aXXjUkfWhFn4j
iwaUFNSTCKC5WxgpUQ7gtH5NjAYqPd0G1G4bdzWnFegaxghaCQf9mGDAzl/Zf89Vee01cTtanYFq
umk0XsuRNp9Ak1HLOtGRRxqNlq1CXbC/2XCgKuCxyxPd1tw9swCesUoIvxqiTdB3bexCHjOvu0qm
h/ysJ6uhdk6eP/Gk3P7JpFzmUzXy6k0UyE505oNAsJdIOX9O8EHHSBh3ETCDJRKz5bnV+FkefpFZ
u2jZ2H6i2wn2xI8yoete2oYAk1t5ZMEcf87flN7NaGI4uv6sO4TQ4t+/Qest76sJlCOOdf9fpZcB
UgS4j6DGQS/VCQhqMgiHkMlUKS8rSg3Kb0UB7+yY692AegW/yHxj6U7CtLjLEORw/chlof40YvD9
U28eDq8mlc3mb0E1OOTU09hCpXQp1ozZy3QFt6Vj00JiYoCSR3l5UtyTfKJnlssFt+NA+L7XPvia
n3UDs1bFxbA56CUrS/4STuTyX2NCFXtdGuPvHNt4RX0zGOpr0fYANeseRS9+kKVrud2kl/TskNVp
RThhw3dOOAashz+x9Lc6LvTiwgcBhGgLsiXLGYoo+fb8lEOeJTfvrCiFvaWZypivgquNL8XqTG+h
pYrZj0qLa4TQhjmX+ZSADfWPpfDqPpcz5LWECyI5c8nQMyEcCv/GdORnGp3NGBZ+3V4nPhx34rTd
WINKmgrGqMpkzdm6J9WYDhp30BsNDGPVFI0PLzmvjwvjFXXU4YPblBk9uRf2SX3V6bcqfU6FfYQw
rxn7zPuqxeX8cOj4CVNspXhU6pBAYCVZwvaLglDKL4xyhm2kjByu76MtLCrCqqlCEy8EgJGCqBaK
y5uYH61bB3Jp6ujqmMISw/WiG46zZjtIGYQU6gOn1aQJTm8T0MB6nvMS9kboovk0a2H/TOsJpLVx
tlhFSZFmjYCXeRCB08WnztVoVpCoYxK+RK7zMVtx3qrRO0FOXxIVLHLTgAzDlmy1a9+5v9U7+ZSq
Y0qovuvovQhagKBjl1jxy7AQENXN9QHMZ3v2o5lXsiyQgGifF1ePqohn1NjaOdJze94zoCva18rC
CUTNUnVI0jo4E3MkyyVve3KekGDYUrCDThv5JN/A+bwYRG1AKsoGwkCfZMBLcTmbj3cu6/4y/LLf
cAhkstnjQBAwUjbAy6uVup5xugT3D/2VZnH+PJ1073tuzYaElT6VTB93klJAdGBCpTel14uEwScz
EE0DDactONv3tK6sANTcA4jswYYZyIx9Zj7V2zmEYY/8UN+bOTrmrV0okOorSGug8o/WvSv64j1v
e8vQr73cdLi166y0RQRrdOkJfsVNKeW4N2r3Mn8zyD0jd530crdUFWzk0rLJQchAKgfQ6Uz09v+G
sggD73vsvrGgljj+LlByJv7jjTsOImX7GfltFxQimi34+8KEFnaCajrVjTVj1GL4gcbWEr0TISQA
yj/KlDE+ISJL70uWSTVAibAcCpLJWz0IQPC2VK6nU+5qqKsOQBvCkoSdPWV7A9S3RQ6AAsWcepZ5
5LL52I+x/7uc8ceB/45ZG3KTuoJopDwzwpGXIfve/KR9RJQ3Y9mTBD0g+y9FxNGRl06sgN76UlSM
sbfr1lTpDRQ8e2by1sWRm0UcFhBkXlhLa18COs8R7Rz6SaJ7yls30lMaaYbYUvwi9+d1TpGren63
2hH5/2aiZA8rHJWQ5w43nor4CjcmwZnWEmjjGo+8tG8dD8AozCAhwtBr6Lz9iwnFSZ5BuVDMIvFX
CO7y9ls8OzpcIUl0GpSwE98JP9Bu+C4kg7JQtAFG3UCdXTA5uFJS6LAfh2KW2IfJ3NC8Nxr+CeVw
QEMS7/80GiHT2D28VRAuqI+E31iz4JJZdj+DZX2PKmVq0/SrkjdvaHAyawlzfzjdZB1m0cHFYMQA
m/F1p/E9jTr4nF/A3dd3JvLiI7MfP81oTl8HVa4WVL/QHfuim5r9o+aSYqVm6txXDYfNN6fWMUtK
U0Y7e/CmOb8QcYhNKgol8NjPMjWlIihC8hOND1roa1R4X7+cc9A1rxNdOGEOM1pLIgKMZth2Cijl
4SMWJcYAaqBA0Bm63s2yPg1xE0Yd4NyDwtufpsbBGUc3fyrjNjXTZWIAhMZBUBxwelbmYzmp4C+6
QsJ30b6uT08WEUpLdpmO6RVpYHvnjAOJYpcMzBepTFSFzHis/6IhF9omIGDqNBADHNjxeo7kFJ79
NMrM5hoh3rsHCh8ViAx5Uz92Jx+o96KsAkG/5PGRTw/Zm1I/3jrf9DeblhRu2BLT3C4+nkEMKaFn
gRLz4cCN9PyJZOYVtuAYNrV1ns1++BbKR+pLv+3GfN5d3/MsLcCvEYMObEuGB3l2cXtLgjsDr2sB
VExANFyyzuS8qM5N9KZ+dJQDvHLk4Lj073v2U5gzQ6Sr21n80X5xE4WamIOgNU4FNrLnN+lcr+zQ
R3rLhGp+lC+Idst7IdFqKhEFrWU1o20/DtyDfTbW3ZfPkzCkIgcF5dPk9IWCytjY8GLBorCQWyDp
9/xGh7RndR+tvYIPzOkDT29Ssk6VYzBqznSTRfjZDZ0ifNUmXqH9bNr/CIrocuDjBpXbcxlz383O
AcSglTRO4RibFIoi4ys0nkW92tx9hPLtVds8krK2UU9ByyA+lcyrQC3jiK1T5jDLkAEAy4NGXGBr
qOqfg52ZEEXGvjPQIlVWL+dFY9bD+L/a6+u1tJLfHjyb8fl7az8Oerk80iIJtfEq0rZEGmt6qlNL
A5EAp7Bm+lrl+f/ZOYDWxVPVp99y/zkxhtn5eHYci8g9dNySgQTQaDh8P70vK+HjvA4BcF+n5TxA
fkSm+4pId6mihpE25G5GTbd82ZPFZHgG57PUUSY9mLTMq9CWBdLK3vu607WRYDXzBkd7EczzI/+K
0Br0ckKvuvrxuTqbPw8FB6ur7C3P5DfoT8JrPD3SWGj1lbQ+l2qhA56J1YpcxLRKkAVx6DZQZZRS
HHUW+TO09TlxRmOBHelaXU/Wn+yNDsGDhoAo3BAJTZ60fuVdywVfZm7dMAi5HW5tRIcZH+AQNzpA
aM6geHjEBt20zY2reDQWe4cWV5MgePC+s9A8wY+AEeG3BZqhOgtzYfVOQG3fwCDMEMYY+hu1QhWn
bVnP60QrzDns/2H0/K/NNIorhdanGsKdDnkewPiwMe8Xk4hw3JpdpFiKrLRSMxCTQNIcmY4FKpC4
i/NvZD0hNHt4MaGwhQFFRypb3EqxYKpWXdfpag4dCRiGQljMBKZtF83KfNxtyjSkx/+sQJuI2Pc1
SZWJExtV/PxIi2fR7TWTjwlM8t5bvOdGJY+YScPLXpdFL3a9+e91JmWP/3Ybksx4XVHgGcLccttK
rneFxAnsRfSQY5m8vfTTMesHl/f/pV3bPQG9138rj3MG06ijoaYYirm2gsp2PP3DZqrtenIUHK/L
mNPLU3XAG7+Y1gJ3k3G2v7yacKBPZcG2VDKpuiKzIKzewDILsYFop3OzRF8uY4ml3p/SM9lytP66
1ZD8lhdfV8x4cDU4oUkAlNyd+clqqvMYYxhaYItsHAu3gGwbd/Q2GZJ2NWJ+4KenufZXB7xMolYe
Tl8+1qoOkCGDIQ4/dpkX/PV9hzCoVGZ0mX8mGiVAph0we8pIseMvvKsRvMUebYC7gt1iMAIvqIJV
97/QYjd9buZgSUflmJFDDX2rg7fyWAqQzavDFbDl7niUGC41ErW/wjiTwDtsP7MdGMPzJaueFkdC
ZVYiJUHsiQirf884GOY71dnyfa3hj6Mh49nvXrxD1AvTM0dWJ6H/X3xK1QRiiIQON2qDmvk40zie
IxjgpEpYqMmAm/LeuC0MnA3g4k65Tse0sPlAqjUUSpxCQuZEOkvWmFnYZtrpD7Vi3m8100Yxq9Ud
q83U12yfdLQeCQmi/haInZRqvHket0BNHqiABIVewvMdMJKR5XRTMwvGegxU7cH+lkE7LZgAIDUi
kM5T0SevGAkcZQWMowyLXYDobuopHzcuFdiXztuy+dDCO+2LYbu62L6oQefvAFEM0sOv/oQy8uhz
hshZPGUiyr4SZbfWCC0uJNIBN+zq65m+hvEuZhF09V5qTMbNu8VEYaJ7UuHEnY7cxIfAVmCZyHi0
U8ZE8yzY+JyXK4tj139J6+HdR8VQjdVSCDjpXlRZmqywKg39WcHYys5E7h5SnaDjNPqrApQ0b08n
YfppccUcqwlVRrMNvDWbD2MX5TYUqDoou033neUfMRat9KiOaZEJ0Y+oK4p7ggXN0mv1+MByVPDr
mP9sbtLe44zBBej7aNLF4GfLXDoC/AAcW2wq1fxKSOgb4jLc51zVQHoOpPYq4QRDCMrfUQx8C84M
/AHYzeeT+xONMV+WoC/d6Yn9GhN2MmFtIsnQOjHA9mOvdA1YsIspPU3eDpjvvZhl4cRd9YNrudQJ
foZiOWEgdhyFw1Jn3hDHniLtpsr1nmWkuhfmP7UeBBSaB4AlMNfISoFUxyJrY+uxOYQZwagPK4Lj
m1EuWrnnevLV7KnXbrFtEjk5Fs4QU+6M1he3N9vniHXhikO2d4b7WqJPKbCUcCFbis32ph9ugBrL
z8WY36oDVL0h6FrKkPmeAc31YuMfc+VRT0pgKAVPRp8hXnZQ9OOmODwz/ewQTnggBAnXLndNz7K2
UcVEBFWGeQeaM0gsGMeyJNmvjPukxlEKPLJiBwUKLikW2vWpCducv1QbbMkNNqvpBy+2AMetg5Mm
TtuKC5ZPsDCEMTcrlqVuF51SK26egvG0sRvcLwq+oYPcvoMaceqGGG4GsfRDFd4k6qs4oIch5wW0
0bv1oNaD8IE57tuH8Qz8iytcHcIzPaKBPAHOgO8KgObKrvFAEB1JK7PoS3gOP5vrVB1Bhr4mTry6
DRY2mtWkSQoYZVuMZSQgp2I9gqj7CEis0pBNP7pMwFbgtCNi1C33bcmllFQRlc1nqY8QVWsUhVeQ
kY4wn0cudUzv2hwJsadzNmlbEMI9+TSQpweUm5Q9YzO+39CJ5PmJadD0GNTZrravAUtmjkyLy1eF
L3TTVi7fYESWJ0r204nlhgjMSB3PQBRC0W0f4AOll+ZyAH9EBqWzMNPMRcHJzheqst4PlmzVf5Ig
TOUdgDxBGuNzLOcYev+8+Kt90fI9RfMxx6fn5sO4xLysFN3mSBBXIywLwel519JVxVj9GIr/Hqi9
jOYK4ifltgA9XuMTRKooRBvt77u7iCCewuBSzEft0OqEqloDdPJl2myPfG+lX0v32QNaajJYMNSU
88P7/JIrkmhTSofYcNY9hH5H2updTlZjkzO1zScGqRS5sE74LTHpHFrUmjIFTI1PxDwu+KlMQ15O
rlyG8Ag1C42nbpjVsG8n9xRJR8Lyj6wap2Wg8fLCq43ZwVeh+IQiGxNsUyxG5cO1xtsIBaUpeCCu
6e388bT0HKm7vlr2vsqaS6DZE1VpPVPXXiee6HmgkBxlEH7i78g8g3I8xi/RUUiqD7b/cq9dXC6n
8S4VwjjJO8k101KgaXxDbULNIRezGq5LpOl9pFfsfombUjiKJ5ulnuYnPiFEJrxCT3c80A5I4phT
op4DXNUBCHYnhijnwURqpBMWtxyB/D/vw9pHlykrnq/gufBlj2mIT0aihR5PPtaBOyHHQvuFWxKW
MMlxztA4TGhtiyhbYSaBDD1gT0KnGo8h7+qkTRVpg3cEmo2PbEWYPxn2k/y2G9ldYf321fvZXe2o
lOEwQnQneQx/HCyxj8Iy+36tYIHwaZ9xQHnjGgoZogfjGMVBhJqEWVR2cPhJVvagwt0QuNRktQZI
9vgJY8J6nAUCa7GM/8Xcw8JSOblRQUMbVvbejQ9ChvsWBbT0xQL23oh7KcVrCNv949PAKVpTJWmx
D9TquRH2zg5XKODOD9l8LznhudziH2ljwKY3Q3hZKrFJW1NIn3fLVQOsjcLNX8VPJjVNS4iyhfAj
rtyNotC6R5LVx1CMA3zi+0GghiiYX965BwrjWUzLk/xxJZJy1WLtmlN15zU70JY/XUoqQBLAk391
oMjPP8TJ6O2pdwjCzMrSIX3vZJ12xUrnE4jsxdpCyJLs3PprY3Bu+ReNhrQj2M6za6XDD4cP0uMM
TpiLA+7cfC2wEfURpyFapSCrUhNdY9R6Y6Egbh4z8s0fx6DJqxyxW5JqnPkZrIxza9HZxd6sMI73
L4CZu9RVWAZm3SAKB8Qd0mVj9PXUyM1pOhf3nZ1bEdB9zILv0G5y/HVv/tbTf7rVzyPRTnEY16lp
aZQN2Qjd7LRK0bFNfcKNlTuDIxF/kaaxSnBySJ6VllPrKR84//UtzrwE/OaDDrtzpauitcQw7ORA
v4VzTAhDQCVzCP7jx7eEGF8ldr4rCR83Sxuiql7u5DKxf2v0UK1tg7vW9BaINGVHPfC0k0WBvfAi
OKLVkV3tMu0vdOMLSBB9DCrMizLgupW/1/2A5WVmDNP4RpsrJVGkUAQlK+ZT9PvJBFqz4gOUBJbR
MigXimW9gfrz5ZM7m2w12bXrmSmIbaD8kXbreYCVnZ9XFP590l5Kzkoo+PpxABj2V/Won2wPcq/3
xcAytOCD5fxsHzisVg6RigKSwMcRT25WREyWx/O084+5PYADIw0/yAP9+WmhNRG2kinWNlcIoucx
WaQ/TdOKX1GxT27Vbnmtd8QG+F3e1AESfMfu26uBSMCWATJkhfX0HjyFNwiwMUpX2FwfoEENsoQJ
kgUTNE3KEDfPIPDYqE3RdOvB30z+M1cRcJNDb2nFR9sFSRTj0YuIK6eAPG3xfx5YedpvD3O6EYWT
31RlRSZ5v9HhudqS3HfXzqpZbX9Qv1FG9vXhm4n8Dca2OEVDXlyjfu3GMg7tZ/tEBikydTsx/khz
DK8IMnN12cidjDYewkJuO0xANJsiISuPcv67QKa7seNQMqCk14m4kdimRF/lgYB5KbVF3NxSq66h
4aZgcnuh2b4KLGvkt5JLS79j3cBZDBZ/81a6lg12my6uP3Zp98m/YaGPWDFwMuerDYLvun59LFXk
aAX6S7VVnMLGFlM0I1XBLIFBvV88gS8EFCAYqooNliVrPZxZcQjVos4cKZkzkNZVwmhYl0/UvMWW
2uyNOaje3ps8uW+pdS/gge9z26Lu+zOMxDKN6OqZJu8cbeezL7MvJ3MxrMNHFRhsN34+XXPsMRaO
wksFwqnWOJa4u8zRL6T2fgdJi6QRI7ZeKTRM1Rlx4Mon2alNwX+AEHdU27oRUInMkQ9J7iMdXFKf
/f1XaVYmy859jJ+Rc167YnCWVwsq8jB12GOjoeg96JlN//3Tzq7Mhf5lZ5GZLGVM5ShSG7MNAvMt
TgpPM+l2PF85b22Gt6N8m8EwBXB/e2cSFJYrZ4fmCJlF8QOV5r7NjF2sEYP/k4sXm/BH0NcqE8li
rnqhLscWcUXCv1nF6PaUNkrxuK6hnr3JinXkjgyZvr056jop4oIAlN1Cl/WS5sxCn+9CDbRYGhNF
H4/bCdfoq9HA7RSBwhDLdH/3XTJJp88tFZ+aXk49niUiTPz7hp/aLIOiom8uxbFOtJYWsSXDCdS0
wD3+dw32t2Yao9mvSBtBImMP65MA9OyDpxVvHKdlK5KCossNTYFajNdo7HL++VlAHgwmkpZWGKOk
VR1OcsntRvXH33VKIpaBt98LxL2vfSxaCt4UIrf8zfrB5BVoIgOLUuV4TWLibC9lwpXVoFpJM+GY
V6OpNPJf0g442gH6x+ILiznRK2E6+GtlNjGYuWUfl1TgXKyehLqT2+EscJbXgZxOJRsAGJ5PQmxZ
t8UR4Cd9eH9kne+hcZK/u5k6UmmoQoOUfDWcbGKslYQbH6t3ZLfUCWGJxfi8Ewkvbpj3Ae2cdFVg
rG+Xw6pXaDRoOlSbtPoQolKwslJfEfkoSAtkCmcICzRpbGhNCn/UMmUnuV4HR4AfoGEuROaraQSF
RnFHHBY2k7+a9zRREbi+s4uzNwpjwvUrypPTD2JJde7gOY2E0vfUCE3g2aXNtw/7kOS7bQb+uw5E
yZ05Cyckn1jBvMR15UBxuUOlWXfWjkPoJaf+ri6gpEMeyz+3DnEydvyj41VvLvZgic5SD5YYS7rQ
S6RgGuEDRVnwm0r5UN01wW434D65Mzz7iVOArz/+JEnvcq1bLpDpRGciXNMOxkaIh7jYxVrficg6
SrqpuWs+4rkQcVJ9HIhQaPm6/2joGptIj+FMWt3+4ImGCP09eiF97PDksKZ4CleuE72SReOeOnq/
x1p9HWmBV0efAJp3HoKcHEy1gaAmjCBk98OqC7jRqqs1oZNU44vjFnKDFesAqr+7FZR7m0JZcxxS
HgQm7odFg6ndFSgsOJ9qHSprAOKQf40lztgqN8wnhTvk7g/5IYz9C+roNv4jQOInFWUh+siIH2JC
CWm3k0KXEogedr07Tw/SsdzEfmhna/Ikxpt7y3qmG2aR/so4pQX2PzZG4d5oHLHy2tGWcwQc69+P
r9F2w6hhCQ8v/+uGclcp7ARciaCe8G3zCFBG2MdMzbe5x3Vym1GMHchJrxiawLEm245JzvHjqi4Y
UzBaY2tq7/qt+Wo+gnwziDkFv5Kd4ddsR9a5X/lCQwdmD7S9iNTZ3OT9pC9F9revQkmfkEuxluOc
27YmdecVH6DIyB0eX+VE+hERyaEHY2W8LimE5Zl8SDgBzdE/CUZDyd+kmQY0/Z/NTdSm79QCfE7j
AXcD34Py7TzXuDWlM3UlRVePIaJLgru3d1p94ZU2mQOTc1BKHJ6OV3nLBfrYm3CmofifJyXoC75n
8eiQWY02g7IY+yeW5Ok9ZpmgnG34vm2PHN8b2oG5WXvjDB+Clzyyp/pnzs4k+VzRPfiLp4WIqhv6
oAmDTw8sJpjpxsI+bu5zsgrI/8diulhE7OjL+0F/e5xHnUPXbCfdSDDxxbSaPgh2YzAcPKEz22hR
K3Bgz5uznIxaLrvzZhQwmj2Kkk803u1oKSWOe4csyhqQz9Zxy6p60tjZXVe6QEcBPiLWaH4dZrVe
tE07wXrjUG0Vfr2U9Did0tN23gsKf5nEUOKR0iXVsfkTU4rnspDLxoNFn26Bbw1rcMvUwSqdvvG9
5GZ/xLKwFEJthT76SXzOnLinw+HJVDTDFLnj5GBwrvs+d2fYo13uKUIq0XFxEu6TUdE+DEimtXw5
fvQzUlw6uNYwqLT7s8TLqhGuvvR0O0JOrnBs4BXUr0jaXCzd7fG+P8GPG8baGgtzcwgDQNSboLPm
kNSBEltp8c8qSAu2SJqgzoltr1VhOwwUqUieMVmW73eTUk+oM9/rYlGi95rU+yLU59NfFKQLn+81
cEJTyjxjq9uU+rTV9gHp2Y0X8aTJXxPIS3Om2xFe1OyRsD1R54ZNpN7nJnMhKCCNCfVLaiZeajvk
uaqsKW9drpaTkFrOkaX5RmhYy95zbcADfJbVtPexJS1TEUYNExX+gqI81HSP0X9oL2tBXyyE29dN
sqtZhKC0qHVAd0QPj1Ecv1tOYIWUNkGtZR7ajxDCEtEE5fWiA49rXqNkeSjmh0EBauw///J2d4f5
yzksUwMxYRGXcpOfhJy00iUpGkOsd0cPbOYg6lJ5O/1o2gM2lO+J5gT0V2UH70Btll9eAuBD3GyQ
5lw8jtJs4C87DD2X2tWhLRIfxZgKup6fYpRFpZuyjjtXDJKWhMxa4HYnJMpy8KScKGqrx0IVl3GV
0oM7kQOP0oyn8jnXqywxsblmyrIj2dzwLGFRBg98hzhR5womZloCu3uVlMmCe0x1N2mMdqxyVQF8
n5oKKLnengKR3nHO9ItQqzJZ8Xw5zRhh4AOYkAkkWhEUDRTrh8pySraY1O2mzX2NYeGiRWhDpZSa
p+7Uh/YjfzCsIwtEEZW2e7XW9AMvwwmAb1JV3ufDyjczkXKDYM/+u8jhLxCQkosVMbpaCzfPK/xv
wBp+mRGBqNU7ck61njFGMBiAcOOF0U3naTw3040i/hEYL0ZPkY/rvrLpzX46wWLKRWn7SE8skxks
ZnAbiLIPwzQd5eL6y4C04XVXlrb0lzSBN+GDd7SlU5VXjIhPefZv3j7GE+AAK+UO9ebNbktQmJSD
WX10mlf/JRGhhso6xNPhYbPHMPmG8ky6cIumuvKkgLVH9m/J8MaM5qAKVeBvZLL1CorX37X6Tghq
vGtpUE+x+9j6+eIkaWas//hZrw4YJ409GEAYAz6uBVTlQrIkfnRZNYRBNju4zLBXrVbD0pzavNFW
/HXKyPJUw3biB3bloMFeRWfl40DwrK4JwwWcNmUofjHUzInPAnhW7vUcfH+6UwZM3aWqUhru67XE
yBgKwnRrUAxWTjEhbgKGfycyZaTm4bLx7hklky6QA2MLCq/becJGnV7IPd5BmSTM/n5U802T4ULX
QACidjtF/oAhdynY2k9atUHCzupWes676eQQE/VTTZH2sxDLaWPgdR7c6Y58eMX03iflokTO9snZ
lSD1DepYMm3rVmB5VBF13z3m9mp95gSVJdzi5LPINk0Uzkr5yXV6Bcun8QgbfTxEhA96bS5fUiBc
MvQ+Y4FyOWIK8ioB02FoaJ5tgbcFuIl8YMIsBG9rK+MvkNLV/GAgUssFAAUg3Qz7fMT3AxCsaTct
/N/0r6PUM/NiK5Ngo2T0lPu8mdi/dQc+beH03S5CpOJ8FwV5Dncfi1eeWIGfw0fMSEahHJnsAds4
x9l3RcfHoL0H9p/7d2GIjx+NPPSBY4xIhN18Br25Pyy8T4g/1/Q+cD7mP8bJwySIdIaeFGXvfUNG
vGTF7B5gIJ4J3NDYgWck2ZZ1/gFzQA4wpfDcDfy5YCz5JedJKlY3KaurgRA5E2naKeybXcgxbOPg
FKlzux6WMxseAs5hW7CNfwQ+e4qEEDgV80TNLgeaGYB3ARriUtEFr4Sbtyt0N5ELy7pJ3tBoFxT9
WKtrYV55hcN+npNpZ/wv3/DpsiQs3O0Xo9Za9KcqFxGhVkrTI55kRhyvWr9z2BUi4mfHfnJNo9t7
bVl2lUiuoQv+jM+FXckjMlReSrGP4k6z77ZYgtLY1igwFY73MWf4PUK7XTP/lgXCCxqnavMCJj/A
CQukn4a5tJti87buvCxv5VC+z/oXAliKB1LNlIrk8Epsl/EgLemXctNe+qSXjOmWYjxXET3jJmEz
irnUuOJPjbwp4rMpKIC4XvRPzSyG7Opr0+UQpTQwza2o2hKOEY2ssU0soSUMj6vYZBnZQlG0Dy7j
5XrALd3ZjoPl4d5FJ8ByJ7jKQ8mHQZrMR8FcS0uEU4ybgzfKIjHc9wLjNq/3ZYbN6X298n4mzoXf
/U1y6AuenuJewXAp0ZgwSZ1VPxvih8GPGxatgEMO/dt44WFvTe84bXUKz5EVKU0zEvbvwJl/cDhO
YiWK+qsxXfLjK/R3ADWGXqE9bOKyFQTbztc/Uahm7lpS6bqD8YuCqxcRMXbbvPIqj4zORXaT8vs+
4cM2oMubtxqtvawH2AhtWKcvjySt9lei30Jyo1vpmsjom7v8UpRHfwKPTDwBtGspBfnpr4bzufz6
hybb2QLgft5hagDZVDHsarkV6KFMhE872VdtU/irEPoJ3xlF7cSlvK6lyJKrJDmhk9cA3gnUb9hK
coQ3Ka9Y/cgcd3SQG/4bqanHQy/54CR1/pHMl7lVXp5LRHFJNaSw3z/i8PTZ74aLeNgKxbe2Lyft
DZAX/SY8jmoq/YH+HDGfkGb65t1J5JvPw/Y/wTS6iYhwFCKNszECf9EGsCdzrhD9fq6pcftZZ2Mf
1nn6bhrFrhhvZ3bLRp31bbhPDIQxLpNL2MGMGAhqgmPQnHh917Io5249qVHW1YDMpf8j9w8InoY9
7bDolGNcew/JSDaQfUGJ+rGm/2UKtBomH0M73ivVBE1FzJWLVsqhh16xKcVxJ6yneOc8no+42oNe
TQPIvtpLx/LzyRKQUsT4nDPCC6d3ijOdneyUKvO3B6p8oWNog4jFwh3g5RGTXEzuVI6wkp7MwRHo
zmQoJP7nH1Q1MWz6C6bRK3jbCOa5s6SyuNdmpEl0dQk184xXKWrEkvpv6JzjlWpqGXkZ1t1gDDbu
lLOozXhVCnxo0yp9Myapem6YZJEJY6yL7++bJ0QU+rMSOcTdeNFF3y7kXetqIgKjfAHc5qoIM/Sd
SzUURMA9jqA4mz25fjueWu5eB1kbydo6FRZMycZCgAovpts8grdsx8SrtSUphkUsdIUjIbvkqz2M
VXKNLfCmbIRTdZIjDnY5qVEFSaFmd5JYvmzKJsuoveEzVetIbV0/DAFCQxRqAGDjhZ3Jc020Eelf
c3LpTGttfmU7YtFc6Vzs5eWlds89PL7CIeqnPmzByaEGxUHtowdjJufpRIzq3g36TaKZvig57uD+
/gBai3RRDlLA/sbEryWwxyQ4tEiH1YVWPsM/tOJqYBchqi1oZLaCbV+7QqMPfmzV3aq4Gu/3hYds
yRvlYvuMV+35V/i4DxxNnfnxlez/IO6krzky5S3Oa9aUc50DQiGYEOIjMSee5B3dM7GpLNmQxBrK
Q1HeJi1d9sC9ZwhAI2qYFC0hKOcdIrtPj7tzHV/EIVu3tzdIMI+KhARzvTiKLJvH01pbDzPMfQFE
ZAXC2zJ0+nSiDGtQPqrVpwPDA/tW1JcNbXvMQ27FQ253QM+2WjAIngZkI3gdSSgDRjoAG9q8qVEp
mmz8s/XOusUiJegcpP7ryzn9bOOq6/XSx1zogA4v2tXGweNaWe/PBRYO+yV+y05Js04Dk1smE2/s
gfynUfJ6SC3Oz9K+dMlXQCYs90x44b4LvBMlKyWIRONDltQL6zLKqGl6djfM5BlZ6kLjRWlw8gtS
W7BjWINT2QKWY0TkLdnBAR1jY0mqEQYVSs1lOrcngE6zOLrLtAz6ydP/FDgv3SssXatQJrTFE/Q5
wtmXhbRqm4FT+JJHUBd6HLUGEOsSZSYtGinwLtFOKoWyN8TmtmCox3yh5OQH5AeYZJagJoSbCkA/
vjQHAgsp31q1CqtGyf8lCSADrhABhYQO308vHSVhGlI9tE0lf4GfpVahsXm0S3D+LEbU6NFFEpcB
0SFlxISgKT7bRfxxsHHS8tejxDLD1xjBs/6Bo51vnqOzyHTFBPJlnbuqL6WO+wkdXpWBBd4yF974
vzemgBZPyY7tGYyVfFsahsaZk9SrqN45cxRp2pGXgrMQl3zJb7BzDV3NlcOfIKDb9GnyBLl7gy2E
onqZuKVzKbju3ea84IoTjxYr4BffqZ/l3Kk3SNbGajKx+TvQKowxHemZ/Ygy2xYzboqHf2c/ecPt
fs3u+muV1Da5k4Po1/mFMYmgF7cMlNUiXFx4U66CIDaLANkziQkKwlEECkyvazGuTFmSjxD7DGvK
p81VD9GfHODXWyyG8uXvU2TzF+wDBtgwZkYGMb1hieSNSnaDUcO2yxfy58qXrdj5heSB2as8gcXx
WFlp96B2hxlCgOINT7lwbfgYHL8tJwJkOULCjE96XJXPMeKqiZ8MSsKZ+Gpd5o2oR7eHa5eixX0g
qTZCkl/nq4SFJK7YNElZtTLFDQ2fsBT87PHke6vG9Mikl78drehL5+M/EAZTfNf+8ivCivWAf9jv
C8bB93ICo1VnNbzWWatT2NSqdHCpb04fol6ONDjlYwBdUE4NK46LhiyTTd35GtGRSDdCkJaqDpjt
3iUUzrMtXeI+48P0mVUBaBcAVPut/0br4ysWiSQ1jAW7O5cVg/tSPvvIw3O2WZJJTzuG0S3PT9u3
czVriUnR0Y7DMl/zxj2Ei9knRW6Z5aREyO+aARmyXrlGLgofds4d1dMAdhSshpUi2zwwR+KwOAe+
SrajrnGAXplLBFCAq/jwZDPjJMEHO7e+P3bi+uElT/KeDnCm9RmJQKDSJp11OuvfEk6uZG83N6jO
LhJlL4Yy7uiik/OU4az42gJTBrEy962FPcO2XuZ13UL/7T5TADHb45S0B/4tG9TrXkf1osJAXJJX
A9RH9Yzs2CrrZ+wCUthVXJo/6FgQLNIgXZ0aW9S8BcChiEntB8hyj9irPvPe700AHJY+dI9mm35i
Pt+AH/TvyFFUpugxigZZIvri4PSlUi3+MaTCMxpYE1uD29MdciRhyj2Mi0cyR1tlIYRMXONMtY87
tRQauZplw48iMoSyBBJA6X227eYo/DLWNvsyBEZTgDkqAxgRNUbkbGfjXAQ6QPBUL/VjDI42yP2o
U6voo//tz12zoNCPvL2c6/Ls03qNC6ZTO4dfa1UXfyMNTJdZcls51xig3IkvlujIGOG0loWMhsbX
hj0DPD/Kbmr9Ro5km+bYM1lucPMWx1w9S9JEAkYwvG4J6agYqgpOgJjs3PCk3kSK4BUvt/DdEFxK
alCah47BGd4jBqwYb5BcDey/MhUYdmsKnTCZWzlK9nWXzvaEO1MITTJRTqzeHBRgnQ+Vou/ezJ8a
ZUsDjP8CONwdxqs8pBaNTfy6x/kWeQuTX0zuYaao8/+l+6kiBluvoYR5qkxCSO3tO2d4KVBzEeoV
HakvWnZbDfVw4C3gds4fi8aBlRm17Os3KBz+wJKtyc+viMM5yw1r41z3y9IMLawcstCTYtc/dzus
SFI2cgz6x3jKER53W2wJ+kYRdzV5HH6hoVYN66VPFum8TFj5F2DQG6ekB0Lb0qyXS5bagRgPpkS/
Ud+05kUhEhA39Ni/uWuxefIrAJMFusbkbaNZO0CiqVETmk/LIVSzsKZHRn0teqT2JTA9n3RoG11+
fzz608JdPXxpmGPDVndVgPk4uiTbJbD078EFv8ih7AFHSyU+5YQQYrH2jKTukIxsosHpfasTWGNQ
ofxdhKL0eww799L28xk4RjKivRf1sllbDBjjy+6NTGhkJrhaQUplnV+Xq2bGkmm4X2tr5nelNo+n
uEy5GizT/nSPevYfJYh5NXppPz3PfrzKDR7YJPRbf5xRp+IyYdvG1wH1WBTJrJGCNUfHcvaxhKqc
Pb2uDkaIWZz1pEznMerJ0HqoXO9F/81Eb96h2ux8XfMAqd88qKbAQX3l5nMNgM8LNbGzwQlybhLJ
GBtZlznhsCYF1POeI0EM0NiXR6ci4rAPBvjhkYgmm+Hv4b8HlIN8VVltrMt49R8TUEjHX+soJQMR
qkGdylkZc0Asmvs3Bc6oFT+ip/QdWm/Q8L+Xti355xWzpwus66OeCtuBYuVQuDr9kbHq6GVj6/L5
8G809fwIycMWUVbWSTnujn+O0zpwy2mam+GEWgwt5RYzbGRVY735DC1z6wJB3keXso1ZXVrhQ0Xh
k+HuwI0smqdIKPdhNUrmN4IMzOIxayOB5NHMenL8TeyVM2T5hmDnUElhE1NuMlIqKZnkOeuRk/FV
TPa5417kbrIEWEcZCJd5VeB9lk8yOWtrAt12UOhexwhK9oM/YbIv8DTkhH5N7UTN/D2EbP+bWC0K
CrTyytN02lFH5IabjKOWCtVIsyTlf9pdnI75IWUASWFakSfeRRRwhOgRC8Z2hmrtEzmYbdKdw0IG
xpTpJv0KkE/LhdSRNAr+IrjWYztTWpzUAamRWuTnJ/24VWm3SaHg2W2itGqUXewvxoNqVNrP5KyV
fWIZ/UO21A4nbT9at9Y2ezRTUeqNJzFypc0oQUsO08VgtjNeHIcuiMpI+GVoS7h3FxRn41ugvCMI
7nHq7z6ZqOQtB5dT7mKCkuhTUE5g5X8rVp7jetu3xoCi5FyF+NucwJXeeRdubifLAVRk41l5s3fn
ipL3AKQMGKBY9Zrvn2W0qftoFWQP1GTHsrE0fUBPTm0EeFxHLbUVcloyE0EFqqM6t4+x2YmDcHA3
FYuQ/MdLiqeH4PTLvC2SyVQsilGodnDJ2ov5kpdhSuPXb3azhsWEeQ1ufnNC192FrKAITlKt3UpP
bRNFpwfVA2zGnqI46Q53njCKbIU8aQdxBultfa0vQ3Hv8xdRP01KWWEHMsrx61d8ieWbLKjZHdjK
VkRhPwPl+1ylN2n7075JmpHzVIqp8qjdM964E5Boqe9O/utNNpW/qEx/Yi/RQoZa7CA1JgsmxGSL
mmL9cYTEPTo8hP7ny5vL2UqDwUMTPl4pCNhHEtojdZVQgP+Qbw1aB9htqLl+yxJmtS0Zj4ICVzI2
qRrmIzq3kfgc9o6G2T7JBSJu7VnlhJFSevRcW+dY5MYKfBoWjlMADhS8984XwhGxZDV8Aa5Qrm0z
tr+Q+0nLdHFHG3jIeXf1A6C46uFnPfGtPszuLcqu9ZGqqgQ+GracbfW3TZfgbMQbfu/0f7cCaAWK
G9f681qtzJnf0KzJ9or8Szy1d6cmsbycnNyDZ6iKwyKSy4EYlAMFKbveajXs3b7ASMyN7IqPyt3L
i8Bnw0D2xCnY5BpGlc+Y0mZ7D8J2VGlq+r6Ptt4Z0KvTqtyQpNHBh0txYBl7eijD7NCd/nX3nGuO
uWXUPFEwHFeCm+o0urRQN1yYIl3wOM2+dbRe+1hwNkJneA7lRhZWuvMQHSe1rzwb88/2lk1LN3l9
QOB/EWiGU4aOQnC35Oyy+J22IWO2qigzdqDG2NXjBUnWwMSvn+jjOJhnGBVCI155am+0VhPqq3Xn
6dCyWFy0taXtuH+qR8b/Xh+0EGOQPluJAXGHrwW8cyJuxZxq7iR3DNspTmTID/NeZQ0iUMaZN+Vg
7OrUWMk2XAkmLirwi+yEetnY9l+EvNuCpX8WNxFxOidYi0zDzuX0JAsMzVpy7eXz+q475PPBdy6U
X7o5Gl9ES63VY1LZp2JfPKl/YvsYZp8sysibsh4FvBKmizipCMuCTU+Iq2nqW/Tho784gn8D+2nA
rU0qKBUH74kqK+lGPP3w8yTBYeV+xMBP94X1lDNsbUcAiRGmwKYOW9R0RgM03E+BqvEYFCfmF5J5
PPUtmVvAiil11JCa9UAIFooNifCShrqlUpMGxCAV5WYlFw04czOWtwXi3Vo3yr91mJPBHEPOhXOl
h9J+Eic/M4jWKO1BHAfU83J1qaFaTOhSjuP1v4DOPx9vP8BTC37/3PpfB7yApxS0r3T1RaVPGb/f
FlEmk1J/oc6yat4BW17TJPiTidZuHavmNub0z7fDncWTI4mC0r+yza7okudu7BKI9S6RG3ZKSpVw
yXmx1v3VqLUOWV3lpEmxV6gmbiBH1f7+buicA9Cs7lCeF66mj2Ri9hvUXWqHiQNea7DFNHh6+paA
UuikRG6fa97I9HpSLpN+BDPwGDyEn9pAgvtNhHpkpxOHfHhfsDFgRbBbCsCpRpWxAOnVAfO3qFez
fKDd6q3bXlwWMHWrW29CbplhztrOlBaTlIt/XSJz0GlLI7BhWwvsdY+HIZbA5pN70SLzDJ6+PP8a
MO2SkxHMWEUCSBNx+xTVeqzXHCOMMZ70IDG4h3A1aTZcU5scnwZx04PiBwJoHjxtRKU3+iQEv0Sv
KkiYGbh90oSD/Dr9Wei7AZ/9YYatSdzWOq64q2wZwnIcfWoZXxri9TQSyMaTVM4/qSuzbC4WAlkq
oonpQxs7XeYGhzJrfawXRZ5G5oq+/lsaAzt91xPVaUaKRGl5Jl9rAXId4/DUjXqGwjnYg+Yn49V2
EfbM/tNgz8mUoo+g20KmHXvB6OF+Fbb8FzQeUFV0Ghky9uhDASExihjTzYxO9GqceMnkRiZlsj7N
5JJWyOjmTLrpK3lqCue3HLh++YP2DREDDBAZiOaVb1wIUL747szp57Ui5zXDLCroPLOlfXE7YcFr
tZTXhCZ2Bo0H4Cz9aWEvzDtrpHPVyWquhxq0SS8TVfgPSWdsT3rvP22PPwP4RDPESGig9aunPGvo
BLP2wgZm97cfp6rxvwobwDBj2CTKY8mPNhZQtO4lkuHepXDvvYsdojTuMB5tV6h/MjAhVS+6WTE7
YbZzsY4HV+r+pni1Y6YzSeOrB81twrAoAzNkTN1+2Jy2ZcUhSrzy9E2QU2kH8C5MSlQONOhrJ2B6
KrjMggcKwsilc0Zc/5v6hD+WDiSfKZjvWkrBmoPUfJ8gd8ZopgFsNwMw6GxV6dM9CeMDwrAnhpd0
ry5e75LAlmJHE0vqbi+LGT7wlkUBzz2Ctdp1x1g1w1yIZbkT5ABN5HY18aI0KfchkwiEg13iegpY
9x6sRuLyFUe7H9i1DebrF4t8eiW4eCn/BTCY2qXAn51J/DVD1o67McDAJcCmGrr5Cfo0JaBONI2E
m1asVHLVk4NR/mXmCa/PQGUHSusSx96JXXWbUOr01teRQxL6d6jbHCWvfHKuoK27lcNYrr0noDAT
rbTrx41RRNcqlGZEsvXFjtqXRiaduZ8B6zivFZbfOjMTWuT2iDqZyxvHWxor2fyfYn2NFcYB1dOd
yatnMdrMOMDY0mPmR+5mktauf1bqgTNMfoHcRYnsAhWARzH4pWhvxHjE5gMTEqLc+xok56dceiY9
6kEg82ZBn+duR3zXNr+8Hwh6Pfz2RXSI/soCmtn/rRnyEgbPEB02MZSbRKQ3h5mJs/u5W75opXgB
Ty5e8IYipv79rd/Gb/cy03cB5xZrOjXcSjfMi4HrMkXNtxYIj000EtGaB8Ay/9whbUnEjcBfiqd3
LiyzwcezhC7i0SuH/3OHRi9qexkIKQ9s703GOsRkesFDYMMXgsaK3H3KRRFd80tzbbh4XLX0LCUR
GxF3+R6ZSRbBPMzEtJklBJMrfGa3M15yYN68eeg8CSreFtt1Gfx7Snq5PwtuXNfsfnBXjr/5kjVp
Ahz5OEeZpRu7XGZMUGZF3Y6KGuWmiylaC0NCtYI5bE9yEj1qh1WlKG21xIhVLoc8dEIu82wrYT5+
v+nNdAPmFafHH9qkklNayYgJVQCHsol79E15DRCNZ/Sn0QyW27JO398qzUGwQDynSU0icJTGFINs
P1J0sUdP9/nuKD9DWQolpsQi2Tl7GezvARLXiANfeOEEdAFqPfFsswdnR7kQAnBFQ4BBP5YSuLTK
N0WN4RxvicsfAj2jcQbWeFYOncBArb9bYt3pUROBpP6uyqYuYcwp5hSS2cPzGdhhsbB5m+pXgOwK
lnUalH9phptm5bBbcUxkm9s74DoFctUOXB5opwhlgOqXWcxn0KqBkfkNlt9523jk0AcieY3XpahF
j7KdqooJG6TxMj7gZczhvMpGOMqO4OjPj1OzASbdon6aWXHZxv5K0BXTkOIKZ5IGp7SDcJKSE0dz
iImNSYg1WzBO0pvgo4nrrogztl8xXYfGy1Ybb1XNaphn9KhtYmscoYf+5s+x/G0RevLM89fIT9UV
nJ9d7CIKmAZBLJwzNyOIha5UjZuA/JivBhwvJeB36VRH1iB5EeRxisz+pz/V+j0QdyY9tb4qz4Ft
mvzH/pZJ7Sis2pt01DIwj1/a76hmHRCTxSPkHB+/RrTcOOs+38uR1YEoofwdpVnqRiBL4eVDCbMP
eq1w7BKD/3U6XS3AANWmex9LN/JyTQXa0IE7hdxJEb2iIf72MW+jHltnnQrYSpmVkkir7pzM6eGN
dIZ95SIBq4WUpQuqzVCPGMx1iYtnLQuhiG1x0ligc38S/FPIPzRFTJF/vDw5cCapPdWg6xfJj57a
Q7wUnUKDhIgdMjuLY9IRwsaMaS+CsDS4Xoo06XLSDNGiOpFecC52a7H5V/6c0e4o3jQFTfOCu/TK
/Nz8SRspunBnEJwuC1Q6xsdW9pz5/BGOHJPf8QMS/FjSfqsqFxnQNuIzb/V70oujhFRbNVi9JdMb
BbZeccxKz2sdPXIGDkEf7xN5ujZ9pea4F+GvCIrbDw+P3BQkYlN7/d9hnvbufeQoUW9zDVKa8SBp
aJI6Bo3p8ceqqp8fs5/0jh/NT2Vqf4SvrkdPQQrHUMapgIQCTQQg1nyUPFjbNxibyKciYN1dWc+J
LbzQ2G68jTX7dOGLkfq3p8xeb+lnH9MIJbJWGUovC8SSof9JzelqVBo+aZzfqJTybhpMLO+pZRTY
AV93Fes4apG4zHrs2V8mHIZ2ybU6a+Z3cTpfzJHBwtlo6gS2+c+vWxsGkuSbu/CidXfHlEJkCrOy
un7FhSrYlSyvuhb075KH/mijgtorji7qpRfyD0gJTEkgEmhmUQ/IxKWCzc5l8JtAFRsTg5GgOpNr
uqxRk1LToFrUUFRWsLsE4ZM4l1UzsbW+332nf013TfCyXNdRjApGlqoWflxhBQGZ7Nro3L271+fS
7pdKGUlVcZCkSSpgCQ6iW4bPw/Huzo0E3NwFaGc70jtr87xvgzc1lA48II9k2eOV6IocZBijMF4Y
xvtyv+Ji0himEkYh7kk4crZyqYk1PzTedRbMQbSisjqjBi7z1JbLsp49+W917ei4x5H4bK94nxTw
o8wOFe3S+Qwc88VjA/rVHv+YVQMViu/8Cy8qw9dB4ZM/RJUXJM5H+xYBH9zkjs5Ls/fnA4vEZuRn
bH/QaeobIGGT6hWb5bOzj5Js76kE31xyaQJakrNIM/zcUGXoe3nN0ZEatbyyxP2aPtx9bD9qcvtK
0UW/xAS++YIJyIU11nxZ2ytfHj8Q+EYSCasmwf0CZpWPVW7G68rD99lNeqOS8JIXCdvSvj/klEx8
9LrZwT3cGu+wesQ2ChHFQ/Q3gsoAyegOBJ7gaqjd6A3TWBrft3oATr7ej/4pXf3heKNb+NJXofzD
RUBx3uLJjZX2Xom0mFwlb8FQn/1DYjDJCTPRbO0NFKmoaRAPQ4KGNmL97k4C1ZRDjY5DLzR0FQAT
bu5DzvIDv+92anrgo3StugRBjB7BZKob94ZImiL2ArUTr8sYb2y9JyrjzIBJEcb0mFXGbzG+x02n
WEx4Sc3hQ9XbDCVi3ZASzYHxO60NV/JRyIfGgZk4rZ6e7aOQcpdDfBUSagExuxkyZJlyoRaAZCMq
YLeDeWaxRVM07dvgkRXzWWOf+uR700BR038sZWuGBVsRoWlsNUFmTgzhAF78TqRR5zvlnd+lQB1P
chBaIMIO7n6LtfaVHzlfxU6SZUqnEoXRYhmbM/DaJ92L7h4tI+96Qv2OclaFUsxZa/MBlUqtLT1q
Ny0qZIzqjNYvWokIHyT/TN40WhcXLI65lBY4iDM4aRAi30d4/F66fyZCEdozyh07dj2zvgivFTcg
3Gg5qrTY/09C1ozaUtFKLhcfmOzuicXo9BFEFzbERIKF/yb7oyDSFiGTUHPiVfAYcV09yxloPpE5
zOWIRPnLLydSGBwOMp1R+76an2rZ+9XDtmTe9AYW25SmU37mVs7hNWuUH5NEQkJJRXjALwcAw0KA
tKt+3k1oPvE0RPgBVfRsFciXqW1w69xrxVIZ8ggar/nlniBusdxKPukhk5/SJL7Idt7975uWX2XI
rJ/A5q3fZr6PCUIfnmyqzBT1emXyThLpvZkvht6uBXvU5p6ZrLoAkhfk2IIUE7Sz4tO4GwIpyxI/
U65T9hXQYpAz4CZ/vZNLfsiMMvLp/artIqPZY5IVYVQ+DNmvPVPqM3c4+6i+9k+RlFAe/B/Hcx+4
tTwz2UEz86qs25pjh4DxPy8d+83uZovhmWbH7gNypSUgkFc30DXmzy/H7Qat3F5sCTgT5gJ1hL8D
FYE8dRvvUHR5vOaO/rVqLlMbO5RzCqR/iPmEt2n78hAb2Q8O7UdAjI1vf5HLdzlhDpfEJ4J4WtY+
V3dhYUPePIR1Tn5PDuSi4rNhPG7CFESdqHXSkkDfCw7yL6W72I555vxQKxNaAePxoasQhBX5PkpK
1/8jepyxX2kYPz4qz+HqY396IAJKu7d3bNR/GggeM6IW5Jicx6cybnyeBQo/Wv2Sa7cBXel7abTB
E2+ZfQrgPjvem6C7hzvwJlaXwoeOG+JSWPXVMqNjyUnR2FORsq0fBOh38Ls2OyT94qP9meZp6/kW
SiC0ebYFNABC1e5pKUd8bfm2IUx0WfDRQjgNah24dkoC1a5MuOU+5tiGvBYBtQUiFgXHEIapYESP
8b1j1uDbaaPK+4XlQYR9bKV08Qyf5875N6X5OebjMcN1u36ggPvY86ZXKGoWwhZj7phOvi5/Xtvx
3upJvcIZEyTPPkzcelqYqYWpgWf8CXWTfBJeoF7dDEuBLQAcxDfXX1rzub+VyNmx7dbXyO09O/vi
dXSvn3SS61zwbyelMw7m05NwPCJcK4EKsg+z+WwjyWZZr6YspHSxi6QOVAHPwkJWdFjrT7O/E9xU
fNumApVQQv6SwhrAcZ2grn0HjwLaQN2ZFxr/WN1Iyf5GaKoanM8T1W2xpKRL25TTKx4KCpefIOBr
6TF7LWwKbFepBNzsPsZ9ZyEpype0XLJG05YqeotKA6S62oS5Nn/R/OuDNiHtz5eQ8aXljMYS3jlh
RD1C8MPcHBrTpinn+MNMYls50mIEvs5CJitzNtZJXMviksFkAHJF2Q6frnKfoIM8vpeYDHZkX7f1
wuwEAMOqQ+DmmS2mTMD7U/HplyHxw92iCZYTUehAztaBz85a7Trm+2lWw0/i3Vtl8VwDOXYnZQ5R
6OEEcmepcx5caLWeKp31+uG1gUjExu40UouCOcP51plOdq1Fm7eN8e7fN8LQn6+9NAc6n38QGY0y
xZCx3XKVnNQDfdCA6sEZ7gqGXAf2XvbO6pX9EQ2yxM0mrHNhkcMpdvhnFTvrRti4ezsrpEf1EomT
FT+vhmtC6paDL+cfKe5R3xmM/dPS0Lbvn2lDEpGjSOR0IKU1v9BsyvZlCJZvJXGnpFG4yjFFH8lD
8sVbBM6rCVV3k6wc9J9D49oWdccWEEnWyFJof3DxModG1XHAbe937NYkuowD8gTh1Y6fLCxTEqYL
zpxwRI8TY+hbLyZo+I7P9Ch/Wlx5y5icaXYW6daF+sSdIf4br0u+f8p7n6crt4WljmMMmOzQutqo
qBGHeANH0Gmx1eWfSnf/TQ+g/6fPMjcAw3ivuK2J9l+eFT79svTiUu0DmJcsyNTL+Mc/dQUjyfbw
HkY+DYehMJYliFkjRpenCgS++ov7ErkK+/VwRNWBfOI9blnT0Bj80jqFrP8qQFvX3ZEeuEPDL3V6
aqPaP0KzVPu94pk+XGng/4XKLTfxkqCcMZA+En+gNf2W1wk8Cq++WASJCp9B1AvgZg4AKPygg0R8
7yRhgGgyEW4WucYkhZVPt9rK5DulC+9wx1wh3qMO3JYsuNk8q/Qq36QTPo8kkbyIclB1/8rOgsG4
DYLrrG0EfZRU+Y3mR7BwjkRFzOby9hRrAfWGzT5puE4dHHsiCkfHPRVQoXcD6Z1LhOlV/ko7PW2k
l7wEu/GEhODq8q1NTeRoAJx1AT5WMPlCkRnzItf/mCObfdBvRGq92wyfo6N0V7hJ1Po6rmYpWeVJ
vj44Fo2JsGH7qf/FlS1b5i1SKO6jpKpYB+/KeBTr6MHZ/c12sbD0OOGztTAbfh+I19aIJw3cS1Mu
MXeDeV9Rg4xVRFvjUJesKr8cgHA+QUgB+pIykGiPaJ/Qu6mEeSuGYyJAXObyKGLnhkQ9fj21wlrc
MCO5pnzDd5IbzKjqVpaHZjg3apgF45cBNeT8On6Z5ez903Jgvoi51pvjvNJx8xRuCbmy1n7HPcrL
3+S6cMxnCpDKloacnFIEqyUZ6WVL+69Vb8YE9FCer0lvIPEiNQHvT2EwNCVtEZD5CqPN+ABd7hVV
ys7Fbn1g7fosi1oqOMnnKbNHgt0Mdnn6BUQAJX8Co23nrifiZAle89VvrspmnQa8qx7rn5Fcg9M2
vAejh4rMztLuuEM2vt9T8nh/z4AuUNnlc1H+qZXX8RBRgYOR6Yf8FyGhNoBY7oj61r08sn11eoQ8
18hDiREahBaYPypyDlFZDDadcABBtrIUcGumEeETj9FpN0/sgpCok2byqLsZnbDNaZf7UbFdku4F
pOy0cGUvRYtAvVBs6Jb++sBtoHuP1sXcsd0Ka530JSfXgFvxHBYSqMAuHJJk9ALkKFF6epHRx8Xy
DJlPe5X/lSw84o9y9JhnLTW9g+BrkOoFVNp4CQRORgC0M1Vb/ZMH0DSNvF/j8AYPo12iKdquShx/
EsEG0gPg3Y8eTMRtaFJ5Ws/h4kyIgXz5V+Qr8eaPWPzumbWqGT0TXezbyWBUCIWnkhscpgcdZLuU
ynBQvG6KjjSo0Mv3fhW5Avqi1Z+iCOZZVfwZY4gY9/y9g2oFkTSnnBhsWyi/iCinAh00pU34CDsv
qot8HJArnH+s9jOlnk6ZuvCyRR6+I3x6HNKuSbnoNMNeAVVu4K0vkFtBwANZ8OIFuiWhqz6e4/iR
/tSIGrKanjmkHXxsY69meTlzsgvDN3Ttre/ZihSnwVyjYjLm1qHh5lMFQZUajWAqNdlIv/GlnRnF
XdusH+Rb6aIYi7vCwHM25zc29l77VwJ0EicueyGM1IUBT3bfbI80ioDZnhrXZDTftJQPgGjtPa1+
QzhXjuIiGYGckOYLdijcN5pODbyfIqAtbrDAVOc7umGu0wPdozyrj4Y+b1KZ4FMlW7sWqvkO1+jP
YZj05crY6Z6jCuBeJ4XDku4nT1+PvVI8kyxNSfqSPMMR+FiLo3SK5nUP28KsLzQgQ4oJf1Womegd
hU7ikLCitnD/OGXlOQS4ycRiZS7h/HprVM/oU2zfkmoaFrNiLKWe27ICF5lZX+RSZ1egF8lpEUdu
D91XuSYcAncVQzRZoZ0Hx/JGaegsbDMngP8xECuLBau8AWavcL/TfaMk5BKkK2XSGmE9O14Az3iX
XEFqRME9UPaX1volPkQ5HlmqFtVsyYon8VwLJvTXyuwpBJKs7+dZA7sGshm+eRXp0kSgplH0H+2Q
UdyySBVd0rZBS6BfAz0KBQ4rMA5u7cO8MRnHvz1wEYQcJIdACR8+96+0YssOE/St8Cqmp+tpxcql
obgr/YhhkQE7WsbNIGaQgShxItCXxpAUrDQ3nOVdNZToSXAowfoBNY/IFSBBE0EXN4zXYwG+m2/J
wIYX+qNXqm5YC67dKmZwHQSHbFoekMf4YoSM1TgyvaFUsu60C63KuZKZNKTKf1D4su3QpKhf9dFH
rtESSi9GieJA9R3sgjAkd5JVuYWRHTYGx2/0Hq4ABwTN/bQhIR4VnvztOzNI3fSZgrfA0Gwv+eek
6DzT2n1oCyLn7RvfxZ+Obl2nNH8ZXHLTT/mmtgOG3viy/1bPsdOUiWpKXeb1gzX0xRrRVUbPi0k0
xW/P39/m5yQxeGIOsmvgXW8YgLUu0eHVwt4iHEDSLw8Xoenua0lWJfytIVfXsD46CKnsCKvldeG9
dftCt7BK8brwiBi3l0oOiP0SeNsV4kNuE3Op3GBeUQo9CDwGKKvCAwKX+UFRJR4oE3he3UStYmPN
kYSrw24Q2qmhgQAfRkpW44ux4wWJ9mAnX46CW2SASKYQMT97qrXiPxGiWNSKb3888n6+6+TwRlXr
UQjK4D9OO2BXnCzdoPuk5x6p0sexDzgsKW1ayypbtPCIDmygzIvApRJT1dEbVZvHut05Io3zEiJX
yP5cd5UFWO1RIvff3lPkQKKa3Ng58BtUzPdQEg8hoOhx6K8odmb7JfEtFit3bekLR7AsYdOzW5hU
Xk/GagRI0xQ64btKiaNkjAyjK1K/0zawrwQ3vqXTTP2Ng1mztwyYzEu4OgTYMHiY+8Lrf+7A1lP+
ThCFAiU9yGK8gk6nIjQYee0xO+9XY7qiJfuGSghUG1bkIWJn/Mw1EJ7Gx4qFowCyzgxxA4WimgyT
AQ0GUEYGoGywc5EIszGLlh00p1iKTHaJp6Uh36drtQEyN7gb7IPoOnsLoCIdxdk4wVNA1kiWr7in
v2OGdxIeznpJujDKqlR8k59DfDe+jxvMXUezQYSOmkJCQXiD7gjtaXxlc8hhNAcTg7ltIOvgCft2
1987dXKmzD76jvusUMRZUg/iOkMR3wR+rDsW7Bew2eiodo1FzhCIGP5+crMZ7xcmY1lghPAw29Bk
YdDIbbzwPi6RNNeYoomnulA6IJO4+hmmVzsfMT7iCqV7z86J7/RzrpUP9fg5MDG2fSQ6hYiANgxB
64O8GmCTJC7XqaixHrWJCXixTSHSamRBmjRsuhwXoCxYluPKkCmhXq/jeM/v65pTqRRgrP2/bKnF
wVraRO/c0DTm0rz10T+kkbH3iflX8Q0vdLFJn/GJx61txzosGwQkv5SH3O69cwxBoIrwHiUtc2XE
6f7jTuW4S3yoee2+1Jr0099RwBERmunK+CGdGnkmQBeKyRm/pcK7CPzyzFqwsiyPSf9YgxIgFh8A
j7kYFDVUXhGMUx6EK2l98kgZeLcf9bZO6sNFTYBab3fp2Gz2dfl1pksuFDJt/HzXRUxE4/NyhZwR
8Ry4jLkKM0SF4B98l0XUuFp2L18/NIV9db9pWl04UW7HQU7s5kI3P5oxKuhG3ALgb1QLGuqpbusW
Rvnogf+3XqN9sjF2jB3WpGilseFQDqdQMAgVX8iU94MAzTLMtisJP8weBSjh9Eeg338o98PH2KaZ
9b78HQSEIRXERdONbL3gLkJD0PAUi8naYODbuLh70JAfMeYK92Wnm1JbD16XjX5xPRKFbX5dTW7Q
ws+9BX29PUkVgEHKQcvSTEwFOisSi3smQwr9v9AcaOM3o1T1qhOyIJ6IS9cjrWrOPga2LQFEN6tb
qM8SUhe2/TkY93l2NE8/kB/ohr2oyr7SUmpKb9pU6YIWejxF5P+TD6Y3PSmoC9Pl7DZqNSqBY4uz
lFrrrJJ6NTZXQbXO30G9VNL/yBBV1yJMpdr8HYXnqNOd14KOWbGoqbwA+3BMXA6F6QuzQoTGd+IY
tS2wH716nUp2I4MDetxxvD3Z9lfc7JhEcL13LstD84f9QwXZglFBBDx+dP9uRmbKhA8Su/qJfCLf
URa47aSw3qsYPd99cqZWNkyZ3NvutrYuIN1s73AKcppqzlCMiRV8Z67s5Cydd8VVcSvWmB6VuEvK
rmFCh7gha8tebD+hiq2z+Iel5zByuvCTUq3S7FWYwBlNzzr6iLu2IZcPqZkrcdfzrgFfr4xgK9u2
RwdcgsNotFmuBKRHBDBmUaaY03QylnTT/CkoULBEQ+iB8ixi8ggoMPKwRtfxKvVcMXBUCjsXX38e
s4NZwJBa5sP651/GhytELDT0hYZLFnHTZZqs0hgIzk7cjeInkLBBHbyRpbS2EtFoPNWXC+rmdk+0
7s0YVeKT/TTJ90OhilmUAb7Hjo024fH+ZLLxhQoDK/mAm29IzY3Ack4yzJ8d4XDFTky55zRXG5Bj
IMzhcEQgNlLDXUKxMoUu0Z8smml7FUZEG5lG1DSUWG/yZq23mLhAohdCyIIhQwt365snSTJwURIQ
/Ew8gj5QRgI7KVqDGHkgnKoO1y3xBLsj3iofWxh3TdXvboP+56QJ8BQhRc6xKZPQaidEUQ0jJ77d
pHYeUz/+dhBkWy9IalXuUAzoaxnZG3Qg4obvR4eUrPIi7jlemLI4d9FoZG3CenXatqPaKRjp21hH
WQ3vWuPojEKXPlxrqPYItFlT41FdyB0J2V3lp8Rra7N26fKZqj8ggi11sP5s6sE923hIGwk9dpWi
qigZGnHH1e9wTU2fq71LbXxc3EqDXfLUHhhXl7oozRKqkiC5zwi0pHc81doXtRBHSxEfe8ODGIYG
633+WbEz0yoy1PASoD9sL+jvUCohfjRs0qkiiG958gAPSzl0ehtXWdGAB9nn4E5g0pSnmmklxqod
bwpBRR0OLYB8BcmkSwBzI/ZEg5ff0is4MPX8vAfUTissv+PjE/5szMtC+d38J+oO5fhmnyzsjPu/
HjG5vRjgEsvecwyaqw4Ubj/gx2XaDjjGrlhyW6BQbx/30YoDyC4N11nmqLMJjv+PhG9BGRL0k5Ug
Xzko4uqzsmD68ropv36FqIXTFfhiwDJt+2dY1qbYfIA6ViKqg4O6SjFC1dbUJADKNcJGswaZa/1b
thxvaGM+2JO9FUb8ccIZziLeBYGQXsgZk5qn8h1oqFnwtuSQRbRuK64dpDoX3Iq/HbDRpzfkAcQs
ZZPrq5IX3PPuYM2Dy+v5s5VwnwjpQF4oCSi0gxzDbx5zYIOBgC7ZnwOWgttqk7iG8u0aNt1+X3Sb
fSgiMxLDikV6ifQoIfHYHPzl98kkjYxuw3mLyhyhc6Ev3kDEn2E/yaXZEvgrDrVEi+eeTCiAKsam
H5Ttnr95c0EU1fnKxQp8+pw15zBAMGc9a4ymZ8hygySBa0OFCXgpLw9nDzUgcGlIrhWs7vgAzGNo
EFpgeGaPPmYI/oZfJ0QnSRgr07W3g84w7ud6BGy1r3ffL+AcIHoMy5DiheFIGykJnUmOh0IRPxoN
7fuxGmVd8Issbywghr4nevAIZMRWhQG92LPvDItzMm6QT+QrZlnoGWEDnwXvGidRvpTHUMuiAAlp
sHIQZDqBQRoSqhkHVGsabrFQpbQVS/l9zRI8zWXrK81A5pk+LmfWTMdDE97vHsGpl4a3gu7Rp5rt
b5asfcLEQPS7TfuQoYj8fogR5YCr1KkggyxB7VyeBGRJsvzJhrDm2GcwYF1dauVg7z5mvsZBLRh4
lqEgkoujGl277rAhwJ18PSkJX7rGmLdj5zutx7pjlyYJB3N08XZolW2aqeIyOD8fly7JBLR2LSTR
kG55E5zz0V8rUN4TlZIs158Pi4xXnwtfyNP1thE2I9A8K9WzPfGsEGClJtt5qLnKFBXx8LTOpsLv
G0mxC8iunN5sqN1LdRMifwtRjWv9ldyApq1ocUd3xsn8j+Hfg/eOEKZ5dlraBIwo1jx15sF1xHjJ
8NZ2DB+/6fh7sNFm/AaW6Z1j4Act+hOHbzF/JFVq+ceA16r1w3wNo6Wk1I4ouZ97O0O6SuqT0waM
glsM0P+HV1aG8e92JvNmRx+dDpuxPeBUns8CVxCuSvWzYfaPlG+fSwoMsVRU8hYtaDSquXKJGN1Z
do5b8KsEMNJtGK0QaScYUjds5j12ZXJZU1z+f+ShNvJnPBdreWTme4p/41ZcW4YfV5kkOGNzVkVe
w9yOeguwsCvBkw7ERt9sMc8/8sQ65zLl6cgMSWYPbgmzklSZu1nUUyHF3PWiTXsjpc/AB6ukV8Ke
vyXsK+hWPYs2HDvbRcwL45YMBbxc9VRBvPK55YySIhK0SFa7B8V8sVenyQRhM/PvAMwdXg4v5adk
wIlgfx/es5YltmqfqnIAsk4QQyF+yt3ylJut94JBatP/Ur/vsqY0UYDTTe3of8MjN+pyKKE4FQqX
dQwCNbNW50SBtc5Us4Bcc75guOfoZaDbBlXpQb1Hsn76ydZ1XPcwfJfyxyFAQhOxnEyPu5kK10Sm
Oq0hifYh5P2rDfS/5wkf+x6sUs9VpiWA46Z4HXqswvSGNjur9qo4cjTT5l28ZnWZQ8naDGA2ZqwY
LSCNETiOdiOgE5Yiu+ygO56QomsNCi7n+2ltkS/wrrVfzACNFla38pu8neP+aT4BecMSE7ZiHK3k
fqZkdkVDAQbrJzvRseqg0MFF8Wu3ePEwrR46Ved1XfJgMvr2nFvZzc98BGWHMnU/HoqKYYTUK5y/
VLXzUUWiMlEFZULk6shSj6AoOOlBVyswIpOQEkiQfaNPVN8H5GWE3VJcZWIr6MFrfAqUPv1Xhsnz
AXgKM445LKdqdYMNL7/7sMRdHVAb2GwNjQMNNALZa6H9DeJ3n7bdDBv0G3i7h8IHou2JfceishDD
z36N8pHJbBaQ4aPpJZZu5UFBgnJiZWg08jYOyfs28gRRzM2Eelg/OXjqmSC/pc0kHjCvtrLfI9bV
s1JVI3sbYJj+YnZHX0IDhs0qvr8BQTem898UutVItCbdUmD2a1onnJeU5zpCJPdNtEOKIhZcmOUl
gLJsnchgZIImVIf3EnIKnygrWpjXflkX2eZIRg0mc8YZ0Tj5Z9ZjxhOyye98awGM3kRprcDD3lyl
jYc9t7UK28EiEetbAxQBx0ELT8/CHfCZjyJIOJoZAuBjN0VpWjBtP1xUwjCbFFP16AKYujGtfTtN
8cAcGeh8Vzryl6XBN+3VTQsevteAJuTemWDQ1vSzMDGwCjNCbYU8mYeo4wbQ5N789yDa1SwzytqF
w8wFRmbnl15v1XAJgLiy24gUbsdtJlMxM25og1xQvgi708ZQ8ktoLCWZKCfkw3JefZzc/V1FBTxG
hxFehr6rXL+svdfvJCxFT4KTd2xgJlw2vi37/O4KdMhT8aOXH7YLFjRFg0TosUlD8O5+BOlc7HWF
krmSsf+C5WwrmARNJfTO9gPlTyz1DMGNtM2IhsTQeyqTBGAv4PcZs5WB6mw2SPsp01uhp3wdMRkO
DJPtly57bn38LYyt8kyUEqqXfhWSY/t3yNDBu9tyOkMbFqeupFhLyL4x9ohiVcELLRqgOyk3Q01d
IpAtEpB6fM+QZqE4R3Ib8xCYSADZXL7HjUGrjnawy/Xm+AGHm48d23iIDFwNPG5a2cMABt997OLn
LB50mkylDxJBPvkDvD1tWldScraMFyliHhlxKz+CNxvgC9TuyAfdA9B4uhvGDy6IRqAn2BKm5N+K
uMan7COXXK3C3RBFh0r9c9IYmPfphhdQtsW6kF4R+QeuCwTC1i+BlnTWtV/51lwVkY9pp2YMiEDz
wcAq6AdACnF1q9+uUky5xtQKGQAjQyGbDEoEmFfQ8mZiZVO9WHBpXTGTdy9BZgzbOHJe4sAdCVyj
m9wWKV83ffwToG1ZWfviwJeihOFT0sMbyMPJyNLpOSNys26XFbaA8oTx/xZsF3c5bAJt9n1KkB8Y
t4Vzv7nxOUg//KRvEsTk/xrPHfQ4+b2KBrWl5IfwmaCcdN8Xp7BbhCj2tJO3BaqxTZgo5q2WF+x/
1WC7VZve5XLRLw55eKv+8301vqyH61GnQyCg0G0KO6eineE3rGk0kuXRB7kzjINjPM3FZ0j3Y3o2
WpaRrr9xTj/WTC6so86lGSMfMHjEozS9X6xTERNgKlOPc2MAvavsp2DeWVP8+lEQHFZieNJfsMLG
zXU+OPr5VcNG+STmw+Ray+t+jMsNmkFsCofo4+vtmGLITDBMEaDwkcJtiIJWuXUW9Rte50uMNx2U
i2EDl+9kubfdZI788pwj6iYTfvdSbbhQhABkadDHVnN8Mx5a+scyyttJBP45nQBAOxkfPPJuWXki
LeNEAmMzAsBFt2nvmlIZ6rjrB7jAsJ5MsT7me4dH4ieS9+RawqPgGNX8FNkyCr6YFc2exIlC4uuB
RuYnfsGsL5zvXL9ZoPY4KkLdk4xKduwCtTfokwgsQagWAmFINZtFWjo378KbdAOqfVR8OioxNIEv
8zPMJtnOj7cbntztHh8C1v+soSm5dKMXwWGweJ4Sz7JdqAGYm2DT/KFmlnBfA1Fzbr9CaYkwkVNA
4A4Nult8trwWry9XxjJIhMyKUrXWDBim10PwH3n0ekxPHdi0ieOU+J8ofdfHBObfmRYqt0Z/pYH1
u66XHi/pkbgDSGLqNFFNQLI0spg/p0GtR7zUCV5VLrkvzgLqOWtRvMv5c9iINWDcYYLC5wFAHjuR
5aLZBc8XxUc14NY1T3sSEEc2BCbkLi16l3CXl4qd20l4m1d3kaE5hkotdXtrV2WkOc7LFBO4kUgl
I6Cd1r1fNgjg9ue6ZImzyGzcOZ4PLbt1fGwbr7dte8Rhph5xZ5/dv+f0MBZtia0maKyXQZZJHrr1
fpK2y7pTGTWdLG8P7ALx+oXGrElbmF1J9pgqB5hdhPRSm7q9vc4aZTGvsrkJU2v9u5KW57K7n3ci
2jt0pzwU1VZ5eR1n4ykflDoheMLMCGVh795u/QGWwBUhADADV6SHrqJe0tYrZsYaSRw0mDVFs8S6
n+dXvzU4BmgSf6xP7EvCDTeSCXJCc4UQDB/LICqwNC2vwordkaRcXrYn8v1pZmgFmt2HTQXiApLJ
ltayn9f+rPzFkviHX/ZWgEI2mneIGEa/sibG5iJucpocAXxvR2fWOSZIKajrXd/DQYLnL3qV5bsO
ZD9lxXxdWn5rKF8jwnf6gpxzUcPSXQzPK9aSWtH+q9QnQSqMKJIPrgYisgnZvEuWj4CIFNB7pSVB
BhErIykuGmsfAZOmOjUKTcOeix682CYJuJ2aIDl7T5fDGa/XOs5u2Kf6P7IupjS//SMhrSw/Tvfp
2f4ENuFMbJKuIsnfv27rT9thsELcEEMV/j1HSa+ehB4wFVXy2mHQvuvd3BmbgLNfxWZzqvG0hNwI
ri/Y2yvgLwUPl0GUUiV+TlQUt9MbGL3gu6o6/631jy1dWzuWz4NkXvKqHFmpLi0/tswEJFzY293q
iPgyXkXMkdN0jBrTh+ZTQeszBFEQPQ6MQO7kQU2In45FjltAV7O2HbFgWNXhf1xu4CwUkdPXG7wH
fCLBhVdJBXIekAewXkURTg/wsplZMzjrBmUVnJBpn2/0JpiZTIuCfGWptZe1cw4zAKXioDu4X8ks
6uotgBrUTOeayXdYsTokl6cX3xpmxL8H+UUAH7BnUcH3hy9v8hkpQjMnP6C5az78mCmTzzjx016Q
3wTTCY6L5y1hN5IiQ9PWNMOEmeAN9SloSXYUdaS3JWp87Q6lcsrQm12fJaoOl3jwzF8iaXm2ASoP
/ljPnu9ia5H4TlrFcDzNj5cEWh7jKxwowpB385QXI4VW8k9Hro3GPzcnoeEga4cd/mNOFIVFL/0j
Rfjpf7rMK4PJpHjhFEVpxA6BBdo7ptgc1E2GR6p8m/OCb0UzvrM1nZ2U8JS6ScOTm55NggiLTAru
1DzanpNtlzyuM9Cg7qKFtce/8g9zDuYQ4QOJzBlW4Dj/46sj0oNjFuMCwxAXoT3li7KXASQ/g2N7
I5vvM4+lLbzTeS1zbPMg2FKl9FMxzfnjSF3Wo4J0SXdggwC4yYKKE7/34w/EDfPx4sdtpsBvRWxL
l47YuSNzDs1gQqSelqvpJiQSYgONIYYkXgL3fwnI+TqJNkZs4MnIWNpv8N25XYyVYbms27OPqJ+c
1kZJIN/AQsjQYb2caBo3wp0ljmthAwLF47Pw0OuYYTp5S5OPrOgMeGKeOovT3Obkf2KkhZBMGGJp
uGt27g7ysLfZWmlerEvvnSGvP319MlhTvDdg2BwIVqtw0nce/ZTjiCIrenZsGQN43F4bbUwadQW9
7RWJhIa6Wkm/kAfrbe5WBKF4oPNSU+zTdmLRmtw7apw0/Eea5TbuO0G9BTXQxlGoS5gTfqcKgcw5
cUsHPaJPRQF9bXkct3M3YObf1M006VtD9d6dsD95mH0BKDtJuLEGqWpkzalr3Vp4Q9ydbi1dhugD
ZtcNzeNq5qMLHZiCQcufVB3qntk7vTM6/awG//dc3krm6xAkVnDruM+oKuOGumX48dwmnHAxXan9
NSuoHY8zmf40KVQzZ/hmbcua4tlLAOJ1YqWD9uLvaOCMupewP4N4szfkTHx+Fmrqnynrm1ZS7sL9
PA6YqkhlUShpSLIOTMwcuc0f7JDSxQOVd1MLTe1owxLO96ortRm/8e2TMREQlCjmV4uB4d4IsnJw
Zdi9haRuV7NJbwcWf7InBzEnNTTUNo21ClvwVFSWrsr2J3SXCCZIZZjznqrpC+3cGNRQjDi3SdMG
zFfECNHLZdSC31eGZvyHKwin5bhvQyETQUcaKfZVxx9XU1S4rSsdnmqY4w6fIcc1hApf33g45KfQ
nQV9in0h2nYoE0dLntKKk7TgL+oCRrlhiOpkDkGoOy0ebKG3BmkGksdCtVg4I13zrDTC6ArHJD6o
a6kbG0FM7qyoY+5WOU0vEWVnsANbkZmHyoV1V5qkoqEDlWl8fIBvR8qasJzb8fPT8cMwRLENSHV3
WfZAUjAZrt1b+yup8X9lvEkff+QHGwSUFj87UpnSSyBSFKoX8Z2ki9EGSWonUxkh5dXUN6/P7W96
Gu+cUeLqpODKTNW7ylrNpCXsrvhUAduaSoa8lKjwZjVhsLg1fX3z08bH8ObdghSzN6+iA5REAw0l
lcUXXeWOtsVswT+hdefQ0A9KmiX1ss2ApAr/zaXNCyyvDmMFE8mT34Qq+/0oOW5DITZnXWvyz8bZ
+WwoCj/sfHNrjCYtA5iyrgYSv+GuoEsH9RsSC4Q3TgFOHk6NPMoqwhxDVLIz1BYDsAdxBZFcBb7U
wQxOUI6SntJrAIAN10a5kgtBByICGA/twnyqaG39SCKWHko+jzXkYkObsXKqzPk5jHMycPlBpyfv
o7vnF5V3/8LXhrze/w68GvFLxl7lC/R9mIjzzs/YfHmCWVvg9LeWoIdMJrSoqaJFDHyMvhrJpDod
Qp3U9JJi69CFirA8Hap+++nyJV6pQpElGenqN7HzT728D7T3aNGxvKoKeSzUNCOtG3F6ArfFKuDT
dMKZ5V5ldkaQi8vXDk8B8o9rWGx4q9SD2l5Tmuo4es2LI/vqeDIy287MbtpUCoril5ta8fqFMUL/
FXch9O+Mcf04hrWZmhBjJHZ1Q086Z9xrwX908xBFBAhc5bnpD6hYT+iQF4hvJlnkQrMtNyVmtz3x
Duhv5bopUXuzSXIE/AAutt2QCzzncxysxkjQWOxXukhg4aaHyP3PL/7S6khzio8DD7DGoo6lpUsJ
w339sh/nGGbXqMiTPq5uZv83inh7FZ00fHC6u96VEHM84qV/Bzw16De3g9RpSMFfeMV3EB2SKZEz
LtZCFQ0zXV6qijuzhW4uzRYpk6eyGm+sa1Ilnsbg/N/Mh3YV1BINiy6rY8vZQaTbfJ89gmqEYunI
XPhl/flebSLfWzMbc+0bGiqp73hFVngn3Tag6rYvxwQrqpaQXyl2qviW5EhaDDmgZyMnIz/UJe6p
NZCAUU8+zLUwlgCtm0r/Dejt7W0iIExPziJvgKYh+x+YGAUokUJ3cCXWN1ivSQDzMjhBqeOpQRrH
LdH/6Af/g6dlYBEcD+E+++YPPWECZQ5XFEmnIb/Pxm1WvilDUldPzlvU4DPRT/7ui2ORbl8SZw4V
juA8PL3LzBAiFrSkFrWj/otZRQBQT7HIBkU5EAqxAAHTeuJStON1nXbRdPgYy/vsj9W/SneRZ4al
vMkVOs9K6emKx0fW1gyTf67pKoEoJPwfXzu+MmSqCfuIKArSOSLFywU28AQJaVtLYKMbZMcJtekv
aUyi10k5m2bcKs7UBeVxgzHAcqzJixtpN5PEqp6SZOKQl2lUX1HEXbe0kt/jPWhOR/CU/11CapAw
YnPb3UTSET1rYXP3D4+MmxyrkG2zuh7yXEM5v25Q/xDMC4m75fEyQu2eCu0HjEIpptcl0Dg2uP0K
WjwWNIUOcmW3kqDjv262zqFWPOzHJOgWBnmsbiROs9TX/MEVVTmMcSQVp0oFuz0f2e8exBToArmF
F9qCtQxkPvCG55AAoBQDR2UiJEQM7PCW5dDOyf64f7ab50PXynlwNoK9WpzKRte/J1BNXtfjZUe5
dNZmWQroZbJRNDTufg27Vg6F0MxLAn0wkisTuMwimdaRaX/rhI7+zFgQE1WDIom0FtS746iJl4Ci
IrotzR+sqvahbFMDXubEEAsG6MxXye7yzInTa1zThm88342m17DnRbOC4G8Ls0phjQfAqMiso/fO
Q7d/8gitz5I+OWPskbZImwfOv/FygqK+jl57bGJaTR+Q4mqu3/YkPSy1ITOfnwqSX2/8StJDzXqk
IYEFzThbFUI24xrr0o4ZzwPIGnEuguGnImZDUbPOe5+vwCKNsLeJR2QCOB0Pyq5GKGbmo+sJTmuL
+22MCDNrep1pj2eCp2a1mpe7npl4BCO4bVPDCbHZMaO3oBA2lTmU2r6uRg74a0259cFh05oDlZqD
00mmJLYGC9GSRYpNT9pSvlN1poYnafgEalXBJoWjMe98MQxCeBqAXGvlVjgFpZqSS9R6fdSUZp1p
5WQg+wF7NNifatrIlHenTuY8AhSWkjazT7Lw/N/Wm1jBlXzMYxwblGXdHswTEAxB0zDwWC2dptXe
7lDTac4ASzcrd4UZ7N89SU5oCtIxzjKTglxFuMiXkymrFaOjzyL5uj8Sh2A0kn/340TrGnNhYSll
Rej8ddZ9Q6kSERmk50xLC5+6rhUscyRPc4WC6LeJPv1W09DvmNhLQRj8H/gLQaIPLdVh3QzuII8w
ZT5sZGF7ECgCbRWcgXKbXW2Tv9iEi7fyLL7xyTdj0SwKXqPw4V8yY1nFTjGh0TIjZx1rpPnUsbwg
U/ZdIjqKPGj5lhnYY9uwu5FYGhnOhFKOYrFk3Zao9uTeJwmlJR+zt2xCAgJQ4UDwwim9tS63hPsg
Q+m/K8pd1yGQNJC9xgI20XMpoofxh0odZxP+EJAAHtoAxmID638EJzysj4ittRbKxfgOgtVKvAy0
VM/z0PDvHOUmBGyevlYM9Av8epFZOtMtjCgApOUUj2ksbBJLkGeOfkBGfVsIDd86HN6Bo+Ua5QZ4
1KEASpqn3FDLLm4M8VA8NMS0T9hA8ITjN1STTZlkVj1s099jEtMlZZsAFCAB7TrRD7AUB6D31ByC
Jily/R+5DlMwfKDqqg8fqWSB7eyXqvXyoEINMtX/cWH9Q6HobQdd3ZqK33XTAOR9D0shTHAyGeX/
AXIz/3oRyt+SC6bTrQfI8WJOAGi2bdVsXCjWX0wl+SuJSyG+0nsO81Rj8qqYvOxjLKZMK02sb0bG
ybMOBhnrT5c4S+INuIq2+qlIz1EzHMQnyVTprwmVfhbBu4xPt1ow5a9XnasOMGHzA5nZIy8qfZPb
p1bkRCce2AAWr2HgEnIH7YsdTTj6MARiBkD2p7XYYUHe70e7BH9ZQzW+gEWoxZFj1F/CtgUUsfrh
NMcijesnSImPHyycsrJK0K0XVsETSgyCUQ2QIvnbjNfWLKW5Fx2l3q8f7hEXeTUY8X1QEuFRKgVW
ILAge0ju1PCd0Sb7mqkyZ8ow6SFTAtZi9aN7JphjtlroOCPq+PF2egBCorJYgRyQFRduIb5Vz3l6
WhsmpjmPuCsOGQVtSleqcIQtcCgQs476BQgvTpOAjX79Z/fVCc7E14awVuJuB7R7xwJ0hoUt4Wjh
7ZYigwtssxzVkVt8nyTj+uHzSMnk0KWT7kJvfjFhd8z5l4nthK0nNWr0dswBXtVyFgWj9xwXH1PG
K7RBvnt4ATTrpuMqN0O8sx75RtvGdGO/UcEQSH9ne8Bspy6et0iOwmmb9s/BC5CSalpAPpioSv5G
uOsKuK4FqIbyeiP+hzf6NZvKo1mWlzuEsEYopgZScAzsJnOBQ7PwryRv1ChJS1uwa1oe4/k19pSM
wUJEIFt972YybebE+UFou/yrztXjUCr5qzDOgAf6DfRplAkrOQ4lRMaPO3vzDnbyFO/TlBGSJYhP
ZtCUxLqMAoxlXjzJaA0MPFIjp8OzaSbcmz894AbbFzaT9pZnQiDe17IkAd3/aYFuZ/fPM77rHXFa
iqgqRj794vn0+FZzONTbc04NLFq9tYkS7FFbPmbyc3p3Ha8Nwg62CkrkP3emYLfYVIchM9Jkwxky
6vy5oKfNwD5zDEG6hFfO1UHh+OeS7B/xqgUDwsa/MxqlKTeZAAim14sicOxfGmpFp2C9nhRgxqjM
VnhrSD73GTrmk/xGDVW+VA4vbkNYeFiqbaTIeZCpnTYetCS41sVzX2LtlyMOgNGAx7pwd3DRCjYz
9O5HwOsfQ91PvgARlcMJXwd2ASpbOVvz4jsbzmfbyG9NnYPBNH27VquLLDfeZUn2xtaVcaKVeIfl
bhjlK/602cPOP1JWNSSD4dUTK2oYWpFhkwudh5kwkDICbVT4SfiD8yG+3oHIj4CniYtpcxqazTO1
ETTXYUFV++ZPi17nALSjgMADKbuM3+5Ba2DoAbuVubPub/SkudoOjdT4cSBJqp/Nv/rmw43o4Yv+
PU5OeSudeMWTWA2P0YeaDMFtNPK2Bg5Vcmd9brvtYK9/Budfl3OF90/fRJJZni6IXxO9TfQBF6pc
CQq2uSpCjDZXhDCz+SjwUYp33viSnxiXYt5jgeLp7gMAt3e3sRQH9u4+Hlab/3Ikb6SZQyLKFR4o
Jn5eGRMGsywLvR6gt+Y3jgsWlp8VPXtTFMQUceZPenpqT0gW7Br2XvdlI9x3NKwn3G2A0ujuvuEg
woMo5RefQQVT9pd7RPwJdVn9kCz85h9v5r1yxk0PRC76IBwlu8Ha4d9/tgSgbRevEH8IDp/rmfut
DsNaYnMMAEHEqw5IJptWnZbY+jdUjw1JUlAGoURqpNd4fKYqkIQ/2DoTFkBiE+LApPX6YiyMMlbL
6gimBTeHWO/tYrV7b7BcYtUbwob6v0IlXZ+mdZcT58IuXWVLPibnTB4PxSXAmHEk3jIN05IpXlLJ
SFviAAVLxbjXMd2mrzhzE7LAsZlU/i1bSh5UustqcLNZ7FHCvKIxUGcHc7zbQN9iS9WnZmjzCgUT
8nkAT7m16JXVoi3js9rQqhoeinuMOTvQs5fPXcENHSXkQD8jxZvaCWVh1hMkUCfuKY+rtXA2Bc+T
Dn5Ibly6qhgnEO1+2V/zBoTqihCUCdNjJAFvL+2ov/SN9lOVMC0tYDs4yBO7jZ6agfWbfeJ0k2ta
m2sj3xqKpXKQratalgbUQ5gfjlGznlx0YeX8BZhs6PdgkXmh1VskR2YFBwbnNcK5FlJdLzIF/8p+
SS5fjhJE1LzUoOCCXaqd6VRgcuz3l8mvI3t9nZICCCJa3VnLCbhBzZeP/WLveCBOmrLg61vmf1Yh
4GEZM/g8UGFHlPuU/h0oGjF+dRYg1roBcByFxihtHaetMTsr/i3p1a8rYXHwRGY/DwlenVtG+14w
PYpNbD0oyRVABd2iz5wS64W8sdUc7yIYQpxQY3u7wI5fCHuCKMAojNdUhRKoeR403+NINpntwKO0
Y9s1dnG9XPd9hPnr+t/YzxJyJfLMiOTzvIIsQKPxcR7258vvdiBmqJAxl36AK4wNHgNy29vRjd+n
fpbPxvVoSpxw2cHLxkPl8fhp4eDmcTdR+hjlnxZqpc+vqvEFRBmL3LINuChoUbH38Ay5nc4G824k
EvHDYQllYATDdVt30bBUxlX36AUwABDZ0wFGjIQnqt20jGr1DiOgEeJFLeezX8Qal4iQR4hXFh7n
MsbhabLG17E2qs92o3Ama3Mj/3k7042KTicTiFobvVcMxDm2TFpSTQSukjyxN6HEwY1Np1hYNiGi
vrTUEQ/cSl/pOjVzctwr81wrw69cAmgpRkE1eCqcKA70QyiFr0o5HD2yD617zwQB7gO68deu820V
mKHIYfF5KmelgKuKSaksuuC669ptFIRb/+xzW1FgcwceIo7pgflmFPrAjD5i3Ldv7eiYisw83w3d
Xkz0ANLXpLdzLIo2RdpibGwDilFG/HF8Vz+hxYw46l6j/ILn7m8IDOVmnPTjU2eE17W5Y49LfBAf
tRdIsJzhwsi8K4ufmVR7yfIxUwiEkY0RfowHHFNaxOebpPc3RKavzPIOHvy080NXMGDgS0lS43eG
4hxbao69pMARMmW3NtheMltAViXnbPABlA8gCoL4e3IrEfDwBpNloubErDk7fJLIUFpWeGdBlKyv
2ER0Ai1RueZyEXgEUOTcjkeF2TIbsFumQwIycaH9lPI1pegbi/p8xBXoqb6tRQlJf+Dj6UtPcEvJ
xLNDkK8/sLBbl7xo/gJOH3Ml7lmHCWOjYna03CfPL4pV48OgJxeYOemwa5F0ytY8EimPqdijJSid
2NX8o3hknDN9zHfjBENs7xXs2oysNCzniYXcQtYOj8bYnOrgVppOvPmZBq7BZMHoY5Z49MMQO2j+
2RSN8FMdhoMx0TGGNBBwIUUG97wiSmWT8eUZQ8Cq4wY9IOY1U4UjD/w+JfL9tjZ6J/qj+Xb8nNF2
VwiiNyU7CAzZwwrnYf6FpP4kLJlH2OXPvmAbk1RV8GRu4ZMO8uP4pr6prYcnphJPDPvWy+pqXRDS
xcaz3yP1BHf16As6V5l4BXLNipl+UwY87XULNFYzaxqw2JgSnfBfGei2TmgOpNAnU/ytOvN3inup
NUtaXkn5/vWowq5tQpYHYyMaOaROo5DsgpwK5JlIwjJ34wMwmchb4jCOp8kEQ/BYpi84YaES/lSQ
+OCqQ3IIP24bb5KUe104CTe2qbFMp61SBf/gXl6ZQUSj9LO4PxAeqZN5HJecybWG577Ne+i32HHx
VfggjJwbp0kcZkMEj4H9pA4FXOvrWb9rEfOVw3XKCXgPqwN7K4MiQ1LF0RnfI90deZ1MK2I5XJId
2u0CgBft/v3DGcL2010B/9twqnhE1GC5Y7s3QY0Z0ZXrR26yrS9Ue106vLenJokfEQX5AYv6y4JC
dbtBgSEwucGFyBdvy8p2v2WzznVRivWp/S16GImgu2B7jeu86mXQc46A07dhzMPpGt9c1yvbz7RY
ZV7CoXa/trLVNReo3EDP9H2XqnTmAdbRrg8ROm5J1px99f87H1WSxXehVbw/n5Uh6YZtjUMb0SvI
MrAKoyo/i92OR+zxxbOCFpPc8YImOa33JoMiQHQ89Etk1J3abiwRxqAX8FmrSszbWa2lMzBTWao4
Mqzw7NJ/Vt4NYNlzMGYyGfl6csZiaV3VUK0FPFc3m4Oz+pyWxIDpFY9VsvM59ttFAoWZIuyHrxiD
UO/5j5bmas4RnLPTtniEx8s6lhiMnSvc647atFyWeYZtaETDABHc0oPGKvqbqoVojsldSuPjoMvY
gqtqXHfQwbTHk3DvKoiEFYSooYnI8Hty5fKxd7a8ZVnVR4BftcJ8qqSVAzWeu+zZSB5NlgnxGXsf
wL5KsKqeKg+EV/xqu2nk+uaioSlxuMRHz5UtzL+SuKepSRU5utDdYuj3/dSYFK24vv9PvYdNOx93
Rh4pJGEDhts3FTNg6mfELBJbUItxgrR1IOlhfIq4/KP3gC5FsCBsnshf+3ss6HPQeKwPHAvY0Xi3
OdVEKHeYALlHRcCy85Ktevy6aPOGy7YzdcssgJhhmr7G1HyYtyBwF84sPB5UYPN1Pvqs2NJmrj5i
Q+/MqqH8vX6SS8hMGBOejdJ4kUZyYKvm2+a/3S6MXq2yQLqFaXQi8jMM3Fs1KALD0IgqPhNQzRrb
zJDheSmoa9SWBp3aRIJ89pb3ybSYQ2lb8FibKA26g2OQ/PPPusccCKYpEQ2jx1HkdPqmU79Ijesc
/wToPxwui5Zja3K16Qu2+Kss1VhkcPwdtQsToEjNYPck74HLZi7dDG1bZuHmtIEqkHwqsnP+cLXf
7Ecr/IekQA8nY8KpPKkf1hBDFhTgrv0f/R77VZRquOlaSRPK3/fN9vrBnGNptp3JKg9xg7qN4xFd
fKMWzHPbpKCfG7twCftTODbUt9rZfCItsk+Hk7hGF7wg51gBwh+LXlcUxcs/OaIqnNLVvNjrRzxB
rDFD/x0GYBo/7VyzSo6zwBUehmMYgvq6b/5n1ff+kIloOpNVoUqMQudoGiHdMZIzHlw+vIv2Qb5o
rXntInHNA+YxODgxh+8NCkO+ut2YdbFRFrGOWgnMFTosHg85ZKdvXXqHtDs44o8HIsxen8jttj+9
gkUZKP7zFZVkjYXWjjZ8RuqZRCPjVHj0ufLRE+B2BcnKsvtOGFzCAJJVow3HwojXwZJSJ17GKy6g
sQbXaTDjSkyjo/cf/xsGGl6fOR70qV4GqWhdaYDTkb2+jXzf3Mh+Xf3cnXoOaT2UIM2bb8QV1Jvm
GSZrLx12ZWY0vfKuIbgtcb8frFOQvbv3/UkDCoWl1fWqXZRrlVwsJdnAxDr6t0b1+MbeMRPX10al
DppeE2bYtN1S2ecaV281DPBggKfkGPqbWx7afymRN5Ec9X9s1TCy85R7RW+d5tqGjgj8B6TkUWC4
votsb0UQc4+DBj45sM34CkZe2kHZqKpjsedqafZjYpBMfqWQinnxpX8qV7E9LjSOIvw1Tr7XhwSx
q5xn7PHl5MqVbuUHIUvwRyFQSONMG6xchDLli2eYW9+8YMm1BN5Dbr28QvAZRMGWQmZRFk5Zylcv
UT8xTm1mvdZONi6sZRFRerYe3jcIeHbBxiraibG5mkSX1EUMsJFxNkm25HXZ7lApT30jZx/W4QC4
oZQ8e/2qeFx0BiOmtvsyDH3PPw7dglAA1MS5kAdo5tV3kt50//U0x5BNUArYyVDKp0oxQyGUZql4
hSkzBby9DHMyga3bK8v1NDKH3RMj7UsfY4iVfz+DYGbaDLWDPnFCVuVmc0MlznnXss5CWKGf/cIT
5yVbTYhb6d8BTZRXvU66Tzp2e+b6bw5t/wI7wbR0fgqrozQFBeoxvvWN2nLjc9FuH4NjVXUsCu9a
+Yu+inWYDry2S2gh1rBuo5+6VdOG4oM+ZEuGM6IBzp7jHm+MqD73YZc5bYfAvuiMtzcniHrSUA+W
8akXgTy9COXSpmudR3vYHTG6/pfzgPhhaLehoxVKl0z7y5NxWHY6K0pT3sELggS+ruojVSUCYnhY
JX8EE+Kio5MpAKDSseIOE4W5d+lbya5+zMNtHTDq/2CumZKZQchBPfjJsJW7Dwbgd4SUq0D82NIo
p18wlGC7iIcTv75l5llxHVoH3LRQ9fQxaAZKqtg7ixuXvpfuz2om4q/os1l+qflJZVciQDVHnO9g
znkV9L1q79vh689vgcPCi6tiDahpcE314SmZcWjGiKLJODZWPSnCQW07h2cnMPw3GeY/cNxUKIcT
OvmBZ6yfU1xeT+IcBUbZn4gjoXyMIGITsjlYJSXIkXCX8yPcZz4+shXp2wcz61foh08PvKxpu9wp
Qi9fCniHSNfhtfWtb0I6ip1R481es0nPQ5kO0GIK+3nPJLTUtXS/e+tEaTCmLVhCMgNvwtKL+61m
KuxHgM3KR1VIy0inIzJCnILPUyFU56Eafjw605l+raLX7whISQ9Z6DzC52i5v79Cast8DfDR01Dx
iCh8BwRu5voKqCNWuZ8v6sA+7Zul+HAyRMt0HOp0+m4XHQ4vYikae70WFTKuR/uag+f/YS8i6kRp
z8/2y0SeZuE5jFqpMdaN3rrKcCmQB3s/GKMAdIrvQ6lErMjjHanfQSUh6SMIt8JIOKlOWVN4cRk/
8T8XZIu3oviHD1FmfkhDLhrDJf/9k7D11WYENQRz8cXmTK5DUYYAO88k8iNJpV2ryitQue9dKzY0
yhQxOJL++L25lDUPmY6rQ3Csy978nSUxWeKAHklkmCnDgsk8RTrsW2w/X+nSDFrQaEOl3obNKfBr
xkPhDlD9dUr9OjCps5bvjBhqit0N4Pl/FTrI9mf+531yiU74Ci/z7l02reoeHPGQdw6J+p4nTDIF
Ttw6qEBgcTKxFpotrfCGq8yHyYazc2dUGkpeW1frLpkDNV0GcwSTcPFlT0oFjsT1vPKTs9GtGgUn
h0FTeci9SLAgQT00c3RzuMohZxAVezpFQydYJuhpNI+/DeTDJaCW7LX3KUfi3HGOl4CTQLa8js0w
AefJ2u64mATKrkAy7UsXfaNwKV8ibq3+FFt6tL3BhuX6ACgjKVfO2LaIZcsY4HONH1m6OkAvQNkW
t7v5I8gJJDuvzvfV5wYiTJKwVgFLJM/vwKaNrghCz5wWDFSMYFdW19IAbBkfq7uY1v5A/3VwyBM+
31s5QjBMfSXocE/1JUsSCmuR5sydvr/vajVS4ARGyNVJTQ+BeK22XgnO7yEgCxixNRWuezMC259t
j9DLrZ5eUsdPvdf8ndyk/ReVq7mO/4NzzdMwnNAAtJ54ro2epZIoJ01LJGIQHy/hhiMtcHBVfmWi
yZBo3nlXylOISCPdYjApAKjbniM++gtfB5gnESTP97s0D0wXtvJ9VY5vxaSCH5ABPDRaccA9Vcxi
cK0iWDYNuJqy8JTXWM7kwWHkd89IKGZAQ9rR44/Gdu0pVTEIcxWY6egWNsHOX/JFrVH65KfrBGHU
VX4+UiZ3jSkVhBTMrRu4nUd1udtXGpZb40OQ5sN/JMxGoG/12/r1zNcmCgxwp9gyB9bLz7uuPPtZ
ipWw9wl0d/7Bcw259skZw06imFljXG7lEvpuvtJcMLUw7ngudGEFGlK3w3PDQ63fgwp4OlR07IyM
CUYoF/G+4TjDSNmcVpufNr1ytY7rOjSkF146tY9aGRxaamqJ9dikYcN2MUNOlmVw6o7eLgq8L2c2
ZhUSwSLJT3lfjWtvGxlNKA4mtEDWXq7SuqZedcOQBDMz2sDgJKNyoftknoieTTs7BFB8NKpylfoz
DQXAnrET45j5xcQNqULu/rhw2/N2xGmy0mkoC+OghTmQGCX7FhpZxlXyefXpBrCY2QUCjSuBis/O
pDb5KyJS36bEWFMGjMePTk1CEoXqC34GXS8GwaN7hhIScGCA3PnmI1sX0RNaVIhGDFicYXGlwZ+y
W0AiKyUeHjhjDa1+cqgYvidl8k1l9jQ7MomEJ1YuBRcarjucktsoY/S0sNX79YyWGFcyyJH0Tbvy
A1QeQDXeXTdWND+0YvxodReBZ0W4mEqf9lJEwY8Am/rOsydrNHR2TMuhcN3jmB5p4qt5pJqzRrYp
G//JmCVRAj8Qd6oynOXLXyQj63SDknk7ddDzAugd4mqESlNDGhJ5o/1S0RnP/veSakvOtUHsWqP3
WqiseKqhlK+Qv48Or14jt6/syR5l6Ea500NKTt/w11KV0iuzFJwH0Lukx4urV+R9+/hGG+QI7bop
DVV8oUi+pLmsB0+LOD/C/Kg9NCcZSf7y/mByGRPdI3InNyeKNKg6fXcEEey7eroJ3qXQcIZ2Be2o
mhvMlrhHA3VLnnvOOteOTHX4ncE5D7ttal+vQsW3t7uUc+5pcAezgfvROPufs9Ehmhk0U5Mta9Cj
y24KBIGvA2N3rek07BlG0bWLP1lgvBQmTYWlrVheHsKrbXtay3qFme5Z1jK4NO9WW+QMt1VMONEu
mdFHtfJC1uvgd6XsQzipope3/FDXrHiqwRWZlheJWvOXuQFLvF0FTqW5TH2epAOTqDsbDxbtPerR
UQy7EPmEaJDI+dUDxweLRQcwZJJcpzR9HuKTnBtpiE5vaEL82bNb1oCcLFyupykwK1slT+wIwAu6
LD2IIB2t/NFP65rmVYV4SL1QLe0cqPZ5hIQn/m8iRCACMd+v+HtMpV0/0igdlc8VitJ17g6N7799
8/OrXTMTCSWEmYnuE2vsPLBj7KKvjuh85z+BsWzPit0y2GSeVfnQeU8mBocueGn6fKN228lWJ1By
nT/5toOwmaaEsUuP6x1M2tOsSq3FG+vuGGF+CYNIiIKIIZjuJiLN7b/EvekX533n6Cb1iPai2gS0
wtFU7zwcHOQRTq7tMiyobaV8SZ4ZJ3YqRqfXgzHGGv1KlSR0OPs55z7QVmVWUEL+LHJbPCN/YcP9
kNaszmY+Nn+L6645s1/jqN01YZXY3XqcDVk3MyUf36nc4ZL7GpLJXaSnBLz5rcxd3PnZ+vMAe/k7
rS1ddidhCstFRILxXaS2yWaR4G65yVVS/vd+02rTc5+mKHHcwNB1SPtnTsYpI+d+OnQAy1w6cp1V
89Ql9YnBDT53Orp7RJfvlFCvQ7U4FCgdZhyG0Q2AQUOfiKmYb7EmmHZyFebjQvtVSnIQKTln0fxb
h+riB7CCnQYr/yvnr/lWVDjX7q7iCQvxtEaR5+JTBDoGkrlgduz1GglbqvuWvqef27GiFc0vpfWh
v/9JWrdwCsj+ZgyL9I8JKxTURN/1GFjgcTZB9prFkqCvqeFNmIv1UL8cpuIPCu6srv9DqKTdY7Tr
mY2c3lbRMUM2HflIak/MUL356YwxF9dHX3lfLgc0SNu4TL+Fme7VgoTsZXT+dp+/ANrjPT+df1go
tynueHYP0+P69F+wGPwBckf6tnbihgzFC62p83aEM5zDy2qhOEg1Hxpc82LtpJOPOlHLpKT8k7/8
WRAXC+iPc4Qr23dYJJwFBqXrODZ+Flk6jgEKNlgB44Bp5qvUYcDtfkiQD/UdAmDhM9l0ZD7VRphe
Pjk9oqKUj2xDNwmGuwOjUvyXdTcceZLM4RKiS6h3FitQnl2aKCo6+0OwEn6yxA/ahly3HJAXn80J
lWE4o4zcRu7xIzvUmLj2ZLU7vBN5M3r631ASSrYO7Ec6rCaix2pGh9sc5Sah+QhFJ2xUAQRmlBrN
yCuyu4i8QlGCKI7QctB8gIOOypQKAfGEzLdF2c/fbCHefXq4dZDDaufztlFgeX4NHui+HX+e3Ujl
ZUJBSUwoybhXwttOq3kxDPhARP19cP9kpw5aFKAqBpWCuoDuSKrmrxZ89VOszIms0F9ydThknP6J
V6s8WhXl8y+I8bSel+oD7U9DYc0Q06uw6UfhGNe6fvf1FAEuE2n3uySAL9VEx35HcnaKHcH6chWP
nbVHclSzyZEqmBZC/siaihGm0+ORvyLgKsx8ZfXr3RHLpq6XP+x9vdD/jkMuozT/JC/aN7bLgD0j
Ukfygg2Y8dThG/cWKYb3Q71V3UaIcUt0kMrMxrn490F7MNLMonvKRzGREWpPD33D1YOmqCTBp8uN
ompl3jabM1iA/8GF0GgfUP2MkEDY5+7ZzxMV0tmOD4Ia7lL+0c6q2GUfjQBiT8fZ9IXwtRXJ3Fy5
XX0ogmed59Qq5h9VUm+d0y4OdN6TZ+/JGCLXDQMNuQNkPb8lO4RFZiAVUY1XUm8TANvt+8UaMbid
RzWFwcITIP8mJd4TTacHuEg3yFN4+UmEB25zUP8k/Ur5t4C/BtSrWcdlNFciMAoNJxfIbrYQWucB
eR5kLdKGhxm8sBQ4ogGd0aC4SgkQxqCydpEMESYwW4TZk34jhE30IUfYr1gKzRO9yOm+PckFBzsN
wl2DPnydcS1CmxpWDC39ipa0A9t0l2VKdwnFsTlfkTvdbe5xLXBRn5vkqHfOgdibe3cGfZCkNZxh
OTTfkKp/yymTTxMu++5XRiCTkCLi5Rff97kAJHuHS/Z70NW7Hlhuf922IthykQyTZX7LAakTMp04
G4akkf1dtQPiC0rylEd07iyc2/Y6TeA3csGcM1nSqtw18aM89Dt36n2IDnd2VXspMMZGnEubcZLV
6blVRHg6L38q5uK4GoyLd3/VE9hRBkP3tqmXZHRdjArQhEcqlCdtIRAhYU5j6acdZ4ARKJaT05iH
OsGCuZolZBKyQnsu6qvTFnB5DlxVVJp0woEjoL6mfkREiuvrmCi5bqZGWZKlM2BD6EASdSG7mbR6
pnRlmdJvFryFTn7Ohy8h2db0B6Tm+V3CuqVkH/lDP03WHMGZuj7cNY1M+zzAwj/FOFGWIK/6RYIE
NE+swcvoNAQiUse5INznBfMqrBqKlc1XoBDH6Q6lStlU/u3fXwHB1viWU/drZ2dAjMFbmellSRFK
znc56ZX42ZEY0T7rDlk+ECwfA72dMLP2hXgPOg5oujcU18P2XTQmAfDHHnJ8/H4CGhJhtVEOe275
aNhO7WdUIeaXXCTaDg29SrRSlM2srmo7/qRSU51J20fddw5G+bY5sU+di9DhEPO9I0asYt9FKJHt
VXtkdGJQrfLLNzVXtSGTHxJQloxv604OxPXeVDd/iCCs9yyRmuN9JfWcpQV+uHRHAz0vVcxRpFrb
ZUJwr7PpPH5plQwBael4kkd1rFORwDbb5mz/88fuySQaJhdrnYhmivGa683TnJZBr3jbKL9yn/2a
s3icMWyIT9llA6o4mTbjnF6C8vYak6tbGmEZgOf2rSTPW/AbmKvKeQ0QMxL9L6iUW5ztVvXy7HP1
P2G4XBV7gFQaIampbdZAMh/Mxtoky8nDYTFeUBP0srHVUOR+teCGH/tCHDkSXrbaPCB/0nQm0MW5
NfBDKYrg84npM2uaB2ThfsfCwXbLK+ivCD4XgYsajwavraRqtF0Mqaw5vvFB2zYuJfKpyMFoSjzN
yYh0pvNdeozb3l5ggDHiMG3D5oRfhzQcuk1FWEFo/iM6zDSRvSqVCWgMa1ia/QYvtH0m8GK8pFMT
eLnouJZUy1KXZ6LZcCXquAJqUI4HMMi7Ks9ejJDeb8ge4K1fUIuG8YkWaMYLRQjQwM43ZdOZlh0/
ylTen9ewlpvVMWvuBmjUCn1uGW1wk75UgMK4/dmyS2qMrozNNBIWERkr/iqjO3jLkzoZI/M8i+lN
WRdcnXoieva9VfLi/1j/PeM70ICUDoc/6FIkPf0MrZkPQxMfvHrFjIjjxLqpHDD+ySVvzFlMg45m
x1sceqEH8bwoQc1aLwKJtEonKubskqpShNMsxqB6t4x9MMMja4lZdbM0WPhYZW5YH4ExjvEo473h
H1mzow+45u3nzFdlV2/q7PRkihrin1rraaL5rnvZpUWMS5SPraI9rXJTwJA/JvAdT7bW30lS9LtJ
UED4QeVsCgpHlbeWsI9ay8NGIh6pXRG48mjFOU1ftQ10sDr0UPzitVTZfBZFIj7xsG2wLp7tEe6v
0aPpv9QzCrtiDQqk28QTXMRbmOWIexQ8PCJbTAIfOls5nzD2g0ZaV605YFG+XjfkKtZozxe6j634
pG/ys5igN5bS2s9Qd+xr5ULwtIkKHJCI/MbMSW1auYiHo9IAMLL0lpfgVuk9VyD3DrJPlsiPX4HI
m1ZoYJ70ptKs9r1PIHZOFUTEK1lQChSZXm+9PZii/uiW4+mIfRn0s2MEWJ3ugr2gR91ScY492+PJ
3/g0uvgbYRKKdxPszjrWeOwKIZbo6aaQoYuvQSqaskBM6bT/7G1sGPW+++WHce3BQir1fMcKSeqA
ChOYW+dVirCFYEwrTB7Ox1Kh94c2/JXkNZRx88geMVJS3z4WwFAZ3t1E/Q2Ry8hbr5VFgzXk+9wi
VCN6IFq5rsT7HfZaL8TZS3idtU1aGHJSDZtgNxaGGXBDXgn01ACVEFabRfMtA+xdv3u9wcx+wEwE
sEnzNh1bf8ovJAy8McWKbXK3oTcKv29QbSVE1T7C+114V1NVgoj0CQBfLasKLh+XBS00/q/u6k6n
HzTLcuxXaybSJgXMRMYTrd5Xg5f+MXPEW2ORXWZONMSNLfd/RRAzpjvF+qMeMKZf7WG4n5oUTj24
CHpd/bDDmJbaf4jovzbaW4gUtH0nHIezf4ekosTNdbqGsoCTiCxBlCtMpeGAqVrYZg8+jp68Krud
/tU/XFmmeDRjxWanIKKcO4GNG/eqfOqezNENdjXkjPWvhRBU5+USVm3KCntQzQsvkaIDAaayfxUu
OJpbiG+8d8+59NMmgEMWM+ko7bVcdkgXQwW0xvSOt8wjsSYHbAA5ad98cU02OYifXcqAnumBwkcv
TdoUZFDTvA7jybI8p9NzDVjzDrPq33alZIVDegUlBL+laXr9J02gEacR43Qp4C8cKPc2Krp3Fvqn
WY7vq1O4KVbuTW3HEhkOC/VXVNeNYObc8L1SMkbBruQ3oEvTzVhgb9wTFqQiw+pAMYxmNpuFlVyU
WY5dd03naQ9rzvOEEeseREPSfwzlxE8/eIAD2pWf7GH2+raDzcFqF1MxAavv8aVyWcUi1ioyOme1
FnsJP0EHA6IDdiKq5xrU3P9gbmFEEoJfMkVUvVspUZyenQCKH79rtbJ2XGDuQ8LYf36u5+O4OL2K
PTbQcMwh88R6xqMHyb7dqwgBGgM7/v60BqxKiZWOKH6h/M6UIx4GDffXIo9xV4/87KMw1Q/PtiC3
P2O+GX+EFOF0wH2WBPKzllu4NA/na4lHGj/Hs3XEVIpFA3JSL7+brD3WNZZRsm1u+UQjtvXoVqW9
GB11p80BeRifR3dFe3jLds++vZWzxmP5VTR0Kzo6m73mAt/0NfkAZEvnfFNwIM27+iDGsPCiwS2z
JrL5cLyJ8LazMuPIc8mDT6sZqvfAsd4iZgPS6e0Ghelozmyj40vncE0NARaPhTFiA65MhHyMqkGG
iN3/kILFIbSiiaznB0N3mjP0QBhYuMkwrQRdofJgBk1rtjuGUBEuxaPlFM3K1yN1DP6rxaVaxSRO
k9QF8QD5YJk9yzPUxmg4qf8iz9Muh5aMIUznw/zmTrCtI5FfPFwfBxcOF5BCM7tVzZc2bDrRuLEB
G/qq2zkCzWNB950gfjZtmMT1I9CPGxZPDW2aWAEqoEOfAFX1OFNnK5P7HkVwI3xICzeMwWtvL5Hb
Vwfn60GbTTfNn5x3jhPCouFAXKCu85psJ9Z/aLjH8yUTNO/D1+IXYI81hPLEznKeBTGnngl48MIx
ZpNDyQkvrA7akOHCj7Z0DfnVKl6iVEjxFZUPh9gnSwYJyLRGFHoBps+Y9TUYXqkUdd2SXxDUZRaR
cvgCqg498D7hiSq9O0prVXkQ0h6kVkYtv1OFDCGZHTART/JOKlmJYF69Yb7VItXm0mdaeNqwI+Bh
inSpFyGckHNhoAT9EncAONT+DeQQX3HypSQMCVhR53fwnfImiPvg3iw9lqDBVAHQKJDb2C+GpXRq
dcYEEEyWEBZy0vd56G2nsPFqZ2bwNd4ejjAfSc6B2PTWZMfbAn6fbWsvcdft/BqO22b+PtfvxFxu
YgckKvdMYTZpQ3QIRB0RpaI2+6KTbvETCKu+Ff9jliBmpGdR3MNzj8Ltd0sLQSCfV58v6RipJ7gQ
TPC3pzbULEBPe3K1YGp5Msz619mMTnIcLeecAtxLB0W3YPjtMswg10oRAKrodDts51Zb23I5f3LW
bzq948/cVc/dFmzQqMVehvZOaiB6ispmjEa9gjf+xEziptgpnyc1xCivFM1ZDFJ/UGoaowkSJWKZ
ecLUJQ3R9pVm0I0RxoxpEj5n0+qu2FWZzjJtQnslqPFY1QR6MgQFluOJsDA1zYst6nn3yV+bkEHb
MIcfOpXUoT51+A7s+1FHXjcxYl/QHFP3iDibz8JTm7q0sZuaMq2HcbGxC9M+GK5jGiETJecZdm0H
KsdxMw7n+hNA0by5bAPv+4T2CZUhbe/8ZEqTImbUK9Dd+Kk7oYe1eg1gfkTiLjrpiwYdheO0o8Hj
xPENWfiaUTGtNX0DO8DRKb+lCfwZtxIxqHCJgja2I/8X/aUhouRkN4lkwlP2v6PcFaIamkhjffHk
3nHsJby0UHNlKLU97DD6Ls/3XlQYhw7t9MfegmFjw9P75z+z4BGhqw4gu8N7t+4uzABtQOq0giRB
DVe30c01iMAiylwJJ6FAih2uQg8k1e5ttkhfuwqtdfcDMlwkFK8HsvdpLZEbNNuO+oqIZbAhdveI
2t2flQUvRdxnJrU00Nks0SjoqCBjy5Bk1uE92x5R1bxFgm1unegDmiQ1Csg6aMFIK8eyYN8YQs5r
wGNDOxUP3+hs2jraHqM5+qZMf0b2nry+9CXxKIqBqBQAX09lpCdghWOR76drepCryt0FLAM46waV
mIufo2hXps2nKS/nzw2zz1SeFVXviTVNG8E7DV4NQqG0vcrOu7PnSLF1qusGRFipbXNA6f6sQLOu
td2iMwZOHfdQgz0tWPmguLLRBorHCm/BEIztm21ozwEQXa1m0FSZjQdilEa9KBgvIJtHHd0THJFp
x0Z4hoQc3ewfb6Sp6V5OBmZLVuyEz75OLNy3uWCXziXDEPJo4S5cE19o0UVTQVW42qL5Ddm02TxE
zlUWshUTbYmwcF2EE1+3pqsTM/hmiABeRwF9ceRcE6KQdknb7n3EISqOI7x4GviPxgb5rt5jLRFH
MzgHkHSX45ua7V2Yzh/nPcMVTX6yytsGUuVpplCWAlccvg7gCBEj2uh9klRfstZzGvzNpB8wDAok
P8L6SMueMFctz16S2NroHchRLm6fm0WkRz/rE3YqAf93Fkyw8WhW88ccCkCKmVQnXV9nZH9/e38M
n7DkWs4/odxZnE/FOhIH+zx37vhnYMYiF0gIe/Vhys4Og2/m3PbOAjAT/vBU7Ag6bGKbw1E6i9e8
CYcgQy9pWIE8d9kog6iLwDGdMOj30z4W5rOleyJ9vHTTinLcHlnxo09mcOcqzde0RI3I8M4RDDHk
4qW2D3Tyd+rvl/Bv09bss2HPPc/OsqHekqfkuw7bHthWMWj2awW05di/ntpQVU/sUWMYKT9aOseL
eQWMJ9yQ0q+J2/NUb280wztY0EfZ1pSkVbkazNsaxtUZQkXV9fmRCUPihsbrgUYWSgtisOrmvPT7
oRZNWl35N14sk9miERIi3xtMsVK91DUCl+o03HcHRqd9T3Qz9j0iB7fVHIxeaL27uvT7/cK0vqan
aZvxINOAiWSbGr9Bw9DqtYPGCq/4FVJB5ejpV+3JdnQ3kkhTjWx3N4olZjp+uXntJWoLUUtp/BQk
GPAocIx5va8fkP2/X5QGQlt/+BzN5KiOknv5qi+VgNcIPeVsk/AqbCllhz+R5pQfPXkxcRp7OOAr
OpJjtFhH4SwjsKadUf1nGccMemDBHMG2gdv3wjS3EMLKYbDhkfFNp2+Y59re3EHsxzNLBDXOMmRX
e/Mowtzpy+JVGebOssQNr7Ky4NZ03syLoqNayb9NEYKMEw9WHii6WP4UaXaEPeD42ArmDc4NjZAM
tEHQLtFD2Ix59TMm13laIykyef/FrQhwAvgfPC4znV2ezcVPd+62z2AvCSd9S4ql3Tpk0p8OfAVl
Oqmgrum2wxrKvHrF15dE8QL4/Fq1lwAsPIlEYqq3Rs72X5abR9dduWZrZubvFbY2PfpHU1+TskP6
bDK63T2+O1ezjDC0LM/GaOBX97lRSQCmwZuJf6/F0UzxUzwTfbS7xsy3z/KVTEa4+B754DJPUw9T
AUPevXKY19ZvK/vHURbUl23a7mUgvI5lN/o7EsoRPGz6mievgkoZ3KhbRIMTme1MQaqP4c5NFieO
WmeQEWP9Uk42ldPi7yRQyQlMo62DwCPaBB8fyex6I7N3atE5E90KgbAYabqnqleJwb6FtPvqIhJR
1JMIohMQ+3LJvlDp2EBV4O8c/KOnsjfNaeA9plI9A2GqlT537YawFvlF/PuG3J2kdmtmU0cVhcwK
Yz1Y6wyYTarTkeUVymHbVYJ/B3uXbBo8JwzemKMjHnjtulTmmfRncgFRJIH4FZK5zm1SLmBwIwM6
ULYucxFxbZQ0nUON0QkJHps2M95Odno8et8CX5uwh1Fe3HdZq0R9OxhvTVmv5A7wGt92TikWie54
/Lt4uCsj4oKOx71+0XdrsquzY/XsZe7i4rCpRH3kplx0lV4SzOP29GlycULpc/ee2GuHTP+vggbi
2l8rZhTLXkAVSeM42GW12Fstf0ahbvlQVWIuwy4ZxT6RXtCMHEdD02Bwjh8vPP0j1tBp+xZwXsLd
o5fx1nKsXYiOzFK6m9H1iuIpJ37tWwcv29Y52xiH582+BS4itT1v2WLa2ZKbxpyqCrhoPL9jv1QT
NCW2U30KgzticzSYl4kzVC2n0NPEHm9TYPh4uEuTYszMcPNPvtz/Wp98UXa0yh7TWGp2+7w3Uxw/
f7fGF4H6wurXssJK3KU4P4Kq6zxnjSoipNMRTb0mymyISpS2/sT8IUpCMFzODWbPt6YCGkkIgxzj
G1vTsuVCuDELOJuZkWW+ymLl/I0LdpVgPjj68rHKuQmu67BLc4mj+MF33yHO2aN3VNfcXN7SllQP
e8sHsKXxgqzholfaSTNO3GYy/vz6zCaxg54luj8pz2dpHmIgCRTq4Hy/TzFz5/FsjFKJ3N/HE5UA
rE3TS7wPX6mYsTRN57eapGYWo8BKV7FWxC0S/0EfS2ULgFVyMnNEAVy2OWZ6dVOE6ERnfJEOUS58
xPFqlfkLXn2yNsBBFzk4RnAiKHj5DdhISlb+ejNpsA6FBmPYUOSD/uK3UjvS2jWVg/+tE6gFxehP
upStaQRkuRGY9RdoQBp1vpVZogI/B27Nch2kC6etmjPcL2WDUyGIUhUI2tS2UVJDGifcazTLxuaH
SZ8FQb4PdqWrHj6DGrzOc65YQ5+nRx2hq1I1PKGVDEzROyDNF+EB5Q3H7U9yuqoTpBWz/pE5pHvP
Bfm083y0ei7V1rKCEieFrXjtW77T4WUDnXiTujs2oOYnrRYUTjJ6DfkoiCLO0GgcmF5l5RCbe+VM
Km0Cx1l4atfibnRToTfFACXkjJFClQWhzgr41omSiAUpFrbvfs/JUFjusuib7xfUxE71PyAUdiP8
IIVxuyBPqF5+9/UL3E7+4Lg5y8/uyyUIKoC79UJO06TuasrqT9eyGuuoA3ny+MrVjlpwnNp7v/wf
pD8iLNRixz4yli4z2W+RDKIvn6ZGBJyNyK3/lXeJRO+8vdbWAwlChWZMe6TuKUvd9v2pWxzMM/Px
zQpSrKlUu4xrns+fOHA4VW3F3wvefM4PtHNFaiwhvvE+j90Ksgl0e61mAXLDK2pYYXo8rPPOzmyL
NflVyWqECIGMNa/woSbQ9pKsjdXIxq/mQ7r6A4Lj5xo+6+BJmQZz5SA48HX75Ec17Nup1FXbZy9w
tEFSi8SJgbLAjYWNAj+kY5ei46P2TYzqWW0iceA9aZkfjid8ojoKOh9yORWqExBwBnrEY5Rvamcx
Pne0bv5fYnFv4QDsU5aj7NOlmWViSDc+K5pzsBCbqJgH8KE3tRkdmR8U/L77sRqxaDyXCNBWNxA/
f+9DCl5hXSnMr8bMlouXfWaZTWZOSTlravmoIT+jy3idofdNaOShnb1toJh+Dh0jHvKAfV6Wx4jw
6jPQSzz3gMXb5dAtdIc9W6ehS3jb3aQkrHK152Q4db+w8v0/A5FWW7WrHgiLnU39NBXW+MxdbNQr
xYJ5VVujTAKudM79c4h5LAuJ8Woj1eAeRdkd5nJ8n6YUlCYTjDgwIwLs6rrlbKNUGERgwNv0VUc5
zopK4WZb4ZrhQZySX/P4eZBaRhszBBy0Kz8o/Udc1iHdOIxvJntFy3h3WfFnw6LjZ4TQ/svO3VV/
eFdSn1dwRyw/ockMKPeJOgS5SLt0QRoNZtl2SUvC/bMfCXw+lNbxGhMrI6sooN4WICzg8opOkvAG
ilYNR9ReHmbZ3LS8k2VVOMf5CPLm6GDNiFfLfX+UFsIRr1SwDssOlo41PyK8eBYuVcdckvhYIZI/
+gcfRsn243BRzgVGgr8vwFkDTczbxuYPqaKJyqBG5zwz2RVeydTGaeufeJp/FF+1bBS9f0Sqkr/K
lkEtBMJho/w7I9ntTKtg5bVnS2SAWI9YnIiKH+Xb4uRIJ/IY+PmNt7ObM/BVk23WUmptXrA01EA6
2vffkDRREEjMcl24LoIDPEFdjgnXUHzL4i3Fpa3Mrh5GZ1djte0X9Q+vxnH5T+ecl5Jdn0Ou+V1K
Ui0hS2zLBzjgPDwr0Her6JExkWprPJzHx4yeDLGAO90E4JVVDd+mtT4pNkuvHwBhBDgEy8J9qARI
0sY2t3sz3AXHt96f110CAeC8cE8QRx54A6vqFMtmDKifk6cc+2l1TdifxQmeh8QMEaW8Il5bzQNO
4ztHZAR923K4Vas41EwNMqoPguY3sqoXBKTf6+QGzOUAb8azL7dA6DTU51Hmtxs1wxzEnCCO2wiW
IcpwIoz5KWFBZOuE0eoi2uemuLe/AM8wkNWlYjCn+za4SbusLhCFpRx4kLZgK10RdNJae+ow8Rgu
5/xzx16swMRm0npJSmhYuaFfYBon2G8b1pWd/KGPrubKOJ9G6z/IEDlOPlEkbR8COGbeJ9rrwOf5
VwWntKbke+1KwMo4SlXxSoWkydILqTgy+zBBQ7wPj17JGXN8pFsv1nfayh8c5x/p39PyXVRFji1l
oXpYlL7hW0fwjyPzR9w8EVUXZVm3SvZ2pNG5ZSoWeS0kK8UIN0KRR3CkzsB3SantTuJ3KJg1EgUX
fG+Vk+1cIDgnzRsMtXuX9w3KpJdvHT2iH23CCxzx6gMxRZt5AP51QgLj+6Xrp68gGrq807BjhOm2
x3iL3uisUdDTFBRUc9nfMhf9xKVe6i81yvEg0rNlZNoArHFbo4hItYgRu4chEh/uicAKs8JJmHdL
awas8qQ10ehaPvMhKd92e2hIM/zBYz4xKf5LXA7oatQH6ofYeh3vjG0mN9FFFxNR5purnGHntayB
BrriKfKq/fuMWdskBcLe5doPp708cB9AN9JBbBKaesFH2LzX8zbG+5OR19CM/AerZJZU1tghjBeT
uitmtmDt4upBj9Aovu6VEvjcvAfFFtQAl56Kpes63edk94HLf/TRqmjxBuEJMeP+45IJOVRCF9kb
QWAZFwvgECbvrMERKAJp3/5ixsUDk+eoD1T503sTEhKYHsd3kSOE43p48VV7W1wfxGFB1kIjnx0b
kZkL30+pKEv1I8r2mGO+Kjxlx2viTWv+hwpe5riTlQAAnHzXfM43Ec9EwC8ylHiBhXafTGL/IfVS
46s9pCrlxmWE+PKa/vdbPWYm4GDYiJxV1bLLDqOw0XBaMQflvRk0BO48DWlCUOKmQLi37DgjGOV+
ARb+JZvt8FerVYX9VC5F6oEq0GVl3lUoJ5h0wWn8RcF26PuXtNj79obrdbbvwTr+1vbNsTAqN+xi
WSz3+WjyKcp53mPphNW+lZ0z66LPXmYOxfO/b8433NXYUxMO/muUo/CbNnPTNRn8Ejq3CjeYEE4h
aewbmXrLCDSechcGInPQ2iJe2OZ1SOFmjUHEr4vVkhXY5lT8lZjwzvfNFW+wV+/0pyVSVMhL6fLf
EvQrOhtuPVxTOg0RkeXkbQxAtkexoRCfNFsCNrv4Bv8NEr/9fqdwoag3y7AaFcAap2kKQaZMiBW7
Yl3V6+u+lpXkP8xpou2XxupgDHH6muti6YBSQJme9NlIEWxKmpAIqtFA8PQcKxH+g71LqmYlC/AD
n/u/UW68NJaQjhHTFfTRGrJlzF+Bb7nwp1AXwcYytD+Io0jw0i8E+glEeyOXy2VdGJx1j5gWhqGO
40yFSfUYQB025IZJl5rYcGu/qQsz/EDokEoOj9iNw/B6nR2sqOax/pUH09JcvQKAq5V0ArLu2uI7
2MARFLiQDAwyj+m2wg8/oQhVPtMwZRMVa/2KrpV4TLRLRbb22qqavQjjRy93Xy48WBsReMff5EJK
SQw+N0sZQIKFERWK9JXLBGMzTM0OTcEjQgcup+tuWoZleuQqDdxuWvH/ZIjSXi4cV0WH1nFxnS91
E0kbBntLFiOcBDDbB5+kqqM+ju6h/HXdyoJI0cGejoZxZPOx822zAOaeemxpuvlkGa8u5tk9TXd/
Ko3QqXug6RZ7LQkvCTB7Aqf8RvbWE2RIF274ET7mkzsrEJEAfJW8YZDEjB3rx0W1/KOwtIUmosnB
D+O6yLOsIqqg0+ntB6QPbUB/qAZ26rmYUfuWaoouUsEdGB63TOHmG0pAKbsJWw3dj2zk5QcVMchZ
nL25/jZJIlNWJYjffy6Pali7IoN88GRli9NWNO2ftSYo1Fw5jfnTz3PI4dALYZ7CbfYwXYmMDhS1
Le/2RX5bL4iOVQzM12tfXM8oejCaOrGJXhOXuqbjpUXHuBHhQBLgO10Lh7d7ffaWgVYMPrXGdBxp
aX8V/tnp+mRwLXoSWspZ24ZEHGehZijFlEaHcQzMvmQAZpzoHDEyKYMFaVdIogu6sz2xcEaqUIK4
UkqHXY6CtG39XCN3Es00njROqji8+smsY8ia91WriTrA3rpoD+mQ2SQmuLm3Pwj0vdt3aDWh1NZu
9UELWqRPwNjZYnur2d0aVTClxlEeLUhVeyQClQGxSjafhMxemCHMRm75nZeoxwEn/xOghneh4e5d
MmFf/g/6vYioy6rQXIwUJECs4v23A9GwW0MyErfY4boScK/hy6HgTlUOeM32IxWgv4Ov016NSa9o
rq00Uw8p9Qpx3rHYXes+NeQ9T45abQtykT7AdBGKRUsw2etTx+gn7rz2ALTMar3DgQhY3q7IOy90
S+te3fUUlqsWe/EGEriSDNFoqI48v2CU+a3mFGeUE0kEZffvYraVItfSYifrbyEbF1pa/I1I4Eh/
PgIhKlChQUujMFgHfq+Rtms1VFsRWLQgD9zMpzKzwhUmejmtywpVJxbZImxh+PPsnRX6jsGT1YhA
k6ZWWRtFNbWYjiRCvNyDu/9RGiSbLExKnNmkWvlP4Bga1JSkS4GpYOtwzeDEwMTQXyV0VQZqrb1r
Na2CtIc3dKbyKP1UUhRdHC/QVIXp9sRq5Va8cFhPnR/YyYe0vrqp54rbyYKCMacs+LZ33ey2vxyB
Zh9xmPJPs8tyTl8B5bAmJgXRIcP74Lo9NaDrUUM6qsCA+a5nNeu90/wbwpfdxfW0YD+6mj1Yieiq
dXGDvSyOAL3iCYl1DPt0i/LiR9OmCze+FImOiWnGoLVLiQVmPaQKFbphO5qe5igHJvUcppdHO1WH
lk74Dv4W4agO9w+wO6+gON8dNaoXxvhIKgeuSjzSVgMu69rauoYa4WNMwPv++qlfLuqDJ7SURg9t
g2XWNoh52blchXoyTrAqo/hhlUGYMOM2QZlyHgeuf7o8yjdEknGLmTzRl1Ea55IiwnnW7gxRD/mq
4Tc+IyfRd9f4xi6FpSKFSS4SedOD7G5TZgdFuTOeGiYogL+KoJoAeU56nvwDnlIHENfa+ZImRN4o
vwAcwx28ZFulIjTg6e5WzilD1zlmkYy0I6cGndZtYZOqWFGGhILL33Qk56IDgQwG08w7ymWMzi67
tKnbY7+GR9LSmEqbENNhaKOwwUiF7vdyOh4ItdkjIx7KXmofv4Y3VdqSJc7GYaj2Vl4H4eiB7Hme
RFFnWp3hCy5rWcaep6Oxd7mZz5723PZspNlh/c2KUeuEs1PgXl1bzTyVnvKff5q+oie5VJyhk+6D
JKqaPFyD4h2jCBAAJQ44NP4AiMbMDxiEyKXK98IFZm4Pe+ClqYTE6c6/iQzGOyIRPNQmRkl+Igc9
fxtCxUTsX6tXGWp6wTKX30ODycbNmArp9wBrddbcNpdTMqIhq2NpdCdVT+ZU79naAMrUZHVZQdi1
oZYGgs/0tJtHHvOyKZNhC1NPV1z7uBaKDn/L76UooenPhnj/wlfm4uDzi5ltkUsIYmNmBIYFSfuI
ONAQjufs2hCIXsmgBmOmE/sDElKAKDoESxZFL/Y6MoF4isf7JElo8Xi7ZvPo1TSwwYjoYVnkG0ER
5ngo5udMLj05GhqrXgew6WohgLzTkZ2K1Q5/9E2E0nHiwm3+fwhXA69XQ9FdahYeABB/DWwwXoG0
W6cnXATD65a+2Kw+xYiTwBk/2z8nHgfQMbJJoFwcbytgpKYd7RurQpugLEkAg20WjOJIupgAseOo
6vloW6vVDxBeMUXbjUmTkFANlDbiEUbGgpOeJ8O4SFb8geADRel/34wkYZt/b4PTujcZPpMsXn8a
5t0iow/vW/i3bc6mprirFHap0TXNsm9bWNE+vtWMaiUhR1SmZLBWW0rHOq37qEcrvWnz2EuPq749
v13q6wTdnc6p9vCM+Abx/e1ecMwoNl+o3b48ADT6cKccWvVtGofZjN5RhLqluQC8rHh510tsT3e4
2H68QZOmHK51x9wVnd9WMvabPPv/umAYRN6IDqL1AQlbDvVRyDWZJjV0m4+VQZ7gMDjPXTCO2T7f
kHsxoq/2S8mmV5ngtu2yVGOUdHK38aw8CKe6xM2+JOR8xREX+hdsyZxpTs2WUC/CpuH1lVLdXeKc
cmGj8GUyHjuX+S8MHRRFDaxJI8B0eBw8w6usk47d72QRCQJp8uL3J0F6MXCM0pwCm6KOBHXFPIcK
i1P4te8SJsSkpI6RuoYjoRtdf/C30OGs0lOmUzyMhiQLk55EDjdvZ63/Vva7XD/WJdPBqTu7nZr0
Rtoz5D1UlaqHF8G4Qco4zsA8YKYraxZEB6U3zAOHUDjl1a6k/j5j2W2z3TEhVt0C1iYVzatj+Cky
Oe6yAKXqO1NFYPeSmwv0R/RLGyGdYr+XKu8i5Y3XJh+0b9bb7cp8q0ABFsNl5lvxcpXkW5tBdAWB
COitS6VgELH3mwvyGo9KJ3oR8agu3nWhsMr6L6zigfNlDl6S+whjzourmZUP5gkt4TSHdjRR5p7C
NavJJssUNrZLlDUt3sn/JFlGQIkxTTKrI10xq2YDyfa7LL/S26kGK3AsGeJqK5wVupYs7kXHCz9g
acoPAdGFGBPA1LIdjENvWG5ka4QjNtEvQre5/ZVFmH5joKaAwSdyBtwKRp0laP7S6oQNbdfiP+ro
JeTv1+NQk9Vylv8tVhMVD7xAtQKXcU+RftExV35wngE2htF5780iuzOgm4A6BlTPa89s7z8H5Jjq
oStphqvrDDtP9pZhSHlqTqV/89lDJnv1Bg+RNYYlhHTRvbrh6xZooL7wcpq8YRHlLXnoKEzeYTVC
1yAxE8dcgrVzk77gfXhCyAXjZW8myioM0dCoYlJpxKcl8iJRHstDYfnnu8O6m9jJNWDVOPI0reDF
ds78wTTphmTT/yHf+mEryQc4ReB0Js4uM6zjMJp8P5CQ/6YFtg0xoz1pilaNGOP1iazMXKsLGwos
XPAGQfNJpOXpCNoFUBBhp15Gu2FnU/aq22au3E0OyiRkHQ8IQ+xOxwFljPqIQnTa02NP07l3Wawo
XYHKWYFGXBw04HCH3OQrdzLRjbtmWhoUptNQ9Gl8oxQ44Wweh9e3kLSmwVHoVzYfABIzkjQcLXO/
OpTW6msNRFSEfPeaL6r/9UW3EoJeU8Q75KJ77G6za6MCGJ7Q1MV0tw4Nl9Bw+n3mf4htpBso2uo4
5SkPQa7jhtPgUqWmN/uGNKILhQX2KzVOE66Yuq6zqN9kWXVckWkVS4F9oop2XQmpyCPmfsHV/nHU
KacgoxOJxkcBe1WET4sVmpWVu4L5HUWIqVZ5nqGeCbP2eAxaizjTxV1l118wHMzBI+/W8lpbIuxV
T1bb4dPa0HYXXh61a6o/jvj5Sw5ASMH/QuNKHU0LTkBmONAsNFC27l5t7IopFaxFI+t4lpoMPKGf
kcrKiqhmy9d2aKZx/8zW7h0sTUIDPDNn8dte/UgYWSSb3dL3zmWOrZOscP2cshXIgxDEmnV9k6Rc
f0vjkum86+rt0hxisy3f+R5ggZxJyMGirAK9sc0/m5tBN3RF46jvSHzztdM6T0/fbvl11YJgNVjY
GScMeDYIBM/W5fVQvPvar00jEPH73bab4XA/jpyJJPP/JLwIGk6Atq151DW2rvakWelsYTlYg+ru
OtNTA6FHXajS8ecmtZHkWIDBDnBe4+cZuGsyZPSA7Y1fUaKatQt2A/TsvMm++b8suMlhEv2TH15c
htA8HDjLdZjst9BX9KL177jkMsxt2v8S5NSGbU5sHckD5ENi96NMsrDbMafBrkprNbCbJtXuXLMk
WPzQjJFS+S3fmDF1S/lhGMqfF1amcCYTe/8LIB6/XdFombHqZdsH/1YtbIJq4kJAKPDbm1r/54+S
4zM4ytJJhcv5uD2iqz8eOIRgRjNwCES4Q8My2YrfNtMQrQNEBFyYutTh0tXJNCOExNblY0Kr0Wtk
bciL6rMm6pHeefHFTiR7q5GGyxIVw6mbFOdKu/rchgscoDmX6YYqXf+rOyQe+Y7MPHavtbmlOwCU
Bs8sjF3Q8ifXIJMhA4fGexrAA6W2BcXBl1pIpsGIE+ZiGByYJPY1bgCQZRWSHKV3WnuiDZIIehhe
9tR/trc0VofJYF+EoKClXRNg22DZLc3SyBjekLodJFMIE93ozR5TVtJF54b/X2/o0fg9HGqJUGnj
RfGkQ8D9bNySPXP2Gyn2qLxN1o5hCaXJqiRUa28UERvPlwMdEE6oiqsMemsMXLfeXoXvkRLgFT/f
N4oc68KXg/Sj8KRX0ecT4qr4K5sfrXJoppGHSVGa9rAo2Dow/GeB5vxc7JaoT0aBeumZC1DueTeM
lrem6Vw/uIo7DtFdh6W5Y4QYjwWrdmPlRE8sXCRzV+UeZoNJmgdIy1HkEY+yGYcSVYqetJ5ym9pj
YWSo3dw7HFsO8ijazkK51/XFsfAQ9QojJUzQwEOZ+fhhkxxMqWOpoEPcvy/oM9bOiH12Y1ECvqKE
s2+M82cAdF2wupZJs0MOTz5j+9Q/sJqfpWSeuUC6/9y+v9CtV6t4gZ/VUPa/X0pPPghOkbHF1dm2
u9oM/wOLGrCx1h23TT7f9OxLnigaJnBAurXt9mk6I53gIPj4l/EoSFKnjwB+pXfGj5ZEpu9anyFx
9Il3djGc0//i70NT9ZYUcJpXy0QvYE/9WsWJiY+l7ZlEZpBEkZZhicchA/oyW/cjRP+/J5USfFjb
UA/wqJdyRzFfWCYbLYhhZ2CU9rk115r86oX10tUawE0U6StwiLnngB8CIm2ySVqI72cnfNorkj7E
nsjFlsTD6pApOenZ+/Ur5uM2MpzvbpqBdmfAtEdDpRKNI/gMRG9dIEqk9MCTMjceZM0F9H+DGIDW
kYJFkwn9kGYWYY3KswEGXdV4IkeG9tRylB95K6r7V/+RSfL/4uHiXf8UfcieGFGzyXN9UlF52cCD
gdpDfamEPrOesgNZmz4qlnTP+Lfdm1/Z/G3lJFU06Ucft0s/YSz1H5JjwV3JwszY1ixjLF6wdVvT
b/3aO7ki+5XksHZes3rx4FjxFKEz7NMTTHEnwvwTHNGAabFs9ITf4PQkPY8whAsqxmTf00E7jKnx
WUXxL1D25lY6YITnJihJt0Xx42exstonC8IIvF7rXvBrmdLTfiScw7S5U+ykEFBVS3AVzDVM68jx
DYfkzjyGSSx1QOJ+lAWPxUlZvwx1uDyTqbZnyOhEiSWd5ZIdbbAnJFzvMCJaF4626Q74LmhutyXi
B/jbSAqPPyBG2hWMMIJVv/OZqN6Wy8P/KpJ8wDwV3D2yY6IHin2wnZcY5fSvGWfVtCPl2aGrqRbF
F3O6oRoh150K9jhwD3GyyUuLjCegjjN1iMT72q05SRJ09MUze0jILfajl+PIZ9Bdc2yagHZyRS5U
zb4dSzPKF03WNTPLLOqM6UWkuWtRAbqjDidzlWsEUJc0fmIM9d3Xk8Zz7iMdMNLeMfNcaym5zE1t
ZJRfOtddYHFo8YnUJ9XLxbAensu1VDqM/2pE962ZP7wspaVMOz0x9YpA83RwO/06KQYoze3ZKKTY
SoRUUywvu6uAS4dB7wLfPH3zzvMaO/412bVRXmm8fsv+ZqeQR2rxM4epT03/VN/OM9METNTcHA/c
2iQJsLQ0qTW4ZFyCnBADoB0RETTsekp/wZrtOFv5sM50QNWXKJrK99XQy6EOV4OtXRKIKwDrAb5h
o8+Z0yBXf7DUPoMzal0EdcNzz88Zq+4v3AqdlT34pOlOE2kqLWsGd+5wQn7VQ+voaegYkG93NVO6
gD3O95yG+jzLNxulvNqZJHhy6RtcEj6mdOCC/hBxBc3K6F6HX/viB+Noy3uoZEL7R9fMEty7Zc6+
iKYOwp9y8c3wLHwi9fb7ldnk06aLOIa9nQenDKG1pEfT79XZsh62hBBIzekWJSdirhMbu2MySqLM
4pqhyU0jKF9jCNtWjB8Lc8FMDWIc6ulRgC+A9hr/JUgOOaNdv0Z0jiWFvn1gqMIr6JRd7ODT9G4x
0EL1iuRg2AqVJSuPw/m/5IlGCsq1BXqMmnZ4jiTijUHxPU2OrJ6u9pbSa6uX3NfWz+MuRlazMbrH
QZEu3YSRnpq39/az5T3L7snHCbPEHcZsVnCb4JzQqy5ihUEt1+R/1aa/nOWsiZOVJGXM8Cf+tZ/s
JQ5/44JfDmgLtW6JHLo2gcPCGxxNWw5jOOtN6vZrDfcoAK0rU3fhuL+qAko7OSmKRZ6eu2u4iSDT
ew4g8dK3vqBs/9rwm/lRgvXw9g8tdBEhDazCW5sKhvdgqHLbT1EhGnePJxMJdYCKAJrUt9xuxqRD
yRinZHOgXT3rSYYWVSgO5qAm6Ko63aZhVwuuI1eq3cyID0TA4FLXMvt7XRuOKYt79rFfB0t9I6ST
aI0H4DBH/z7gyuxdtS3d8qw+yA830FdB22CH6z4hxlUytK1hJcs6SzQ2Nx5XcF5FWHUi5Swqh2B7
8YFtOd6u62W0erqGeOpoUzUudV91VvxWHB23Ol6Jk91UU4PkmKgoRhiY0qEvVS1QwAUfAvcmjohK
q5pEyRSQ2TkeDO9ClNG9SwOX6tQEDG4MA34J3ImdRc40fwq5I09CVOSYHQmjOzi0iROljvMJdjv6
Rsq5C5NXbQIkBVXV+bpDMk/HNzx8tZqf6rAC1MVtxIlgoFUtjz8idsKsSg70pzuACd27JkkEIZdj
RTue3ddwZJ+jKNvVuMuSiro8VQ1rrzm4wk5FQCAtXDWJbGTAM46N7PtM6aEnr2TQINv78Um4SugO
c9HSI5L59YDJsFXXNL8Ghporq7IrbZA1lbK2+ANRDwXJY8ckL/TnPzMEC2g3kQkN3rVAcduQQpNd
OM2qYwcy9WwM2KA33to0d8YPboFppyx5sN+Pe6RxqZf3MlvWmupQ/cyC00Us10GsaSMOrbqgrMXA
RjM1hw3AcIqPHoXm4lHptGv7HoOyElyhc8iX63j8yuJICzT1XNo9sS1Ed+FcajIDDhgKz9oBfl+J
bUeV2U8pKQq0JIJrUg4izhOaCgYBevVHW4q782V76/l/pofNjgp7drAgskrE//njM3T4sHlhq/vl
Fj2GDHKhFvakB9cMU8yUbU7A8r7FeZFJhzjwsMsBKct/fOazof1ge+F6rOcP1xW4uNCrh7fw9oYh
LXXkJS6l2Lro0addxFDFTWTCV9rmEc8OprH7cOc6MdWgrI3mCLwm+iB2g8PbD9Q8tKA38/Z1eHUI
6ps/xyHLxyXLuz3UkeUv58L9rVoY/29n9kP3gnk8opK4svYX6LKPvh+UdVJYHE+XbA8GE1m3qiFV
CoaBGDdy4pM2qbnKmV6YjpgkVIaoih2P7PrSkHIlvQtdwk/G2jsLxArVjUla2FtSl7P1VNJQ/yWm
lDrarYlEdSgoEyiN/pHAdExBRYToQxlhBOYri1BrlvdHo1B7ByBnLuM/+CyN6ipOhQYk65m6bNvC
AMHy0Uwt1WBkwbY9w5Cw+Aborv9P4tqsNeAl6ciPNpVVpjmuOfET5IDXWHih3A0ff0KXAOQb7KKJ
OEUCoMPka3/t5G+5I0/Rtigf+WEs5l1qKhor7NpWLsRSucnn8QRRbb3wO3Ozt2nsh1u+VjVFulYX
neIz6Nvsz/uqJeAFlvjGgGcIrTVGAx9FIbard15lBFtaCaAoQ4H2C7tBjeNa1VYlA5fz3rqWDhKC
OxFHXEM/LcHpUxuZtfNmGtjxsYizt/5oQ1Q0kZC01jMTqZRyR+rDQjG4GB/n+qlkjoJj8Wm+bCwG
5TfuvEvHRq8kPBmUU9pibvwZlbiJOs/UwZYpUaRACYIhEcPN1qxgavN9WzHcV/AqOG7FfPaCuAle
pdcnt+Nnys7zKa698P1h8cbDmd5sKgSy24smba5PpXqIz/jOWNwI+hJ4JcrRAo4CkvurgmJHqGme
TglJDx7kDn6whGuvD2/Uk6xoj8dYFcPE13ED+aAKbFTzfKXjkxOX+SwjHKeDZhg2x6vwpgIgf6fv
BC7vuEUhxUyKkN1SWBKne0hqir25yhKNBdCvtRQnDkmWqIoMGJzuQPiYx0eENEWFiAZxk9nXuzY0
O8fkITO8SEQ9wlV8nvmKVmbjav+fwWPF5mvYU2Lz0t7lMViLjaEsdFToLuQUy91fcf7DcpnwFJMC
8N1vT9606G80ojf8BTSnrNHbbmsRdFF1oC6EXtixosvSCk+I1kHArXeGFInxdruoetZ2iMP3Fx2U
nu8vVie4zxsJjQlVSQUvtk2gbu9/bN7fApP81OSabl6bF8L5INRXCEWa7ZDoQFAkqd1+87lHIclC
oogZBlTCqO3K0harjzShwTGY+aJ6SF79kySyploQhTmkhEpnHXsGkwhIBC/RuW9Qb0tXDpwOrTZp
0/dERUWgURHwy3+iJ8pUDJgMxsy4X+fsxyniFqfkXCmYH+Fpvia/IlSnpVHfet2Fo48eJ5qECf8z
3x2nd8za2vSqnYMBW87e0TUgpb6LJS5eEodR1lTV4lqj8PXR3s3boiU5AFYYLJcPW5Y+/ud7rDFV
iosXE7PuZxy8OffPhlcki0bnAajn6a8oO3zrV/c9Jy2Apl1TKWln3RvBg5GAz0zpDgryD31DpiJR
tR4YEZWKgTsTiH1hiniYlgyZf9tp/6/VoOFD0a0n04qVqA3e+ri/Fw5bOadd3V/nvR2AU5V4ZYHT
a1Q2ZxsMX6ovcNAb2tnVN30MxLeM0BHE4ZDboBidFXEq6ZR9Y7jzNXdb1qBNNMkfHY1Hjeky7wus
Ht2KhgdwR4QnFnx4n+iFFSmi1qpn8Uj8cOUi6S91Zg3jg1vwNNlEtjFa8GTVmFRHINSzQn63LFFW
9Yx+i2V1T3TIW+7b4iWBsNX0wSQ+0AYlgirzmcXmYor4t0phHOn0Kkzj9Q2070kWNcKENuZbSCxz
UDmTy+VdSP5IXkJBjj6cihxKRrNXl8luJir5tiHTVebmAoZgLge5C0WTKw0YsJXXRZrqbzEJNUWd
7B9DzKX6KTOwTkgPU5WUBQX9gjqStEcjNIcf3paRsowabKhHNgudN+qD32dW2iNHSbMKLoREOCt3
+vu3mAalrdLxz/iJE1h5dT3dflq9QirNj9H8nsU1f0G674AUl7IVjFZDzvc8wZghKT05XBPJA/Pl
MGFDiU7I3xbnCn9otwXpQUxOqScMZAMrfAYwgM88C/fFRAAFtXuQ0AX7TCQ4vHIruYyWybNxhxwy
1CRkdkC6+QkmiJBvWylakRrG2MOfIGpem6PuG0U1Vu/T5YYpzsmru4go4Wn/mrF/7M0yKU3WpjEh
rsou1b+dTo8p+7zjLCxUEbwYltI21TzVWpWstGCQFfItGEUQLK/cYMKC5Ex0TUfz/P3Hh/7BdPls
soUW6MAzjv3UeeXs5msXXESMr76OqI9VXxqkokPL/G/1XuWQtTeGzrRsbA/ZbRufQKJkyi5K2U7u
aZg+0CPYW4wh3XAdbG7/hbVbKl6eDbtYZqmga7kldjDGx/SpPeHnsMPbDdv2llxeTR0NgltgB2LB
9srlLYDir/lS+QTtuSqJOG4z8Kiu03CbsOhw44bzkNYzQZ+F/DBgyXFOOUZqdUF+iBTSQxpBsMQq
bG3RVa+sLEKoGyZhtPovOJxD1/BWZngIU9VRMM6jqx6F0xuWAqUkzPRbSJwJVhspNCQ5GFJMTwPL
H8l6xGEd7Rbd9mPCdFiYs638WuwKrbtYxcFdjd7j4bU18AeTTahAnfPqPKIS4E9FnwrT7kCEHIcv
x+ly0CnzEb999gPZ34SLGTavTFRzsYYqPDLXITWqYAi8VlVxQ0mURCEJEimGJ9kHMszAJBcKcbWd
2x1k5Mgz9kwZmEsFDzvigL02EPgN6yhmEVtIqoBVMlNP8vYeO2BUubF8swBSsuPSn8KZzzUx+saz
HB9ZK99U/gcWe7ACuMlYOykigFCB33nYtdBOy8LbXueOociEtgu8ndKrwTKxUIq2/fzYCEp99gTy
BweJtM++JXSMlR4qO4cZecXr2+Y51QkEYZOVdj1vjWwVHk4exJgpwPZP6GXYtaadZVTLYJ7LYNlt
GWtaNBROvkh0yIHhzVJug58hLueHGpLBoqT03K4CyN2qDBA1OQpLJwwpKoIvnrBdkAjuufbZWNfh
NLNhXMhLUR5ZWqJdxhG1p6Pk0NKbN66u2moSOb3uXnq6uZJwoiYcvyFk/sRakWhgwRE5O6SjWow7
uZzIy2UCczJ286bIDy+FTJR4rAJEDa99J8COkLzZqV3c1MwMcz8zcDpB2jw2dVN5CvCDfpUcv44z
FsHt0yS0TIFZO0xE+rFHnu4X5cFCDXHUyeUGpnDr2ETT8VWVpyMvbeVDA5Npftuvc0+AWuyl2hP7
pyL8wMZBP28w3782nDcPNokmpMCua+s9k09yUetR6okn07a47NyoPUTpT61JexEyCNEFD0VkJrzh
jhBMOQTCLuWoa7dynSiHkhqek6KHZ2qYj8/Dnt7bgiVEoyWqk4q3+d15vVULOGCWMTdqRD0yyGIJ
E8lGJcTkSEHv+zEu7DWkxW6fjuraCX4lucMwssg6ujJt8fZADPVsJAZW+VRmRResUqy2rdCrW8Eu
QHLZYhgz0ozn1abyqq9jwhoSEFSCpxljpt6V3KJ2yFvnSnjPkc52pqCNV6uWimB0Fmb+tfw09tI4
r4tqEG01rRjqhwh7I3XtuA1xSOW5tjmWQ0vXuBY9+lRQITDDK6T1g5C+cY0gs3MHt88didz4X+7b
Nrj1/2Gj2JUe/O9bkl3G2nqs70zmsvoFmEAsPYy55hsjyOrWZICgE2MKBBmtFrCwOE2uBUzE25ID
P6650quZYmvOJIDZrYG4x68IQEi7JJsInwaH/0nK2Sj3ZYkfvxdsoKs1VlNJvhzwZ6rPOt6yu/jx
wktgM0xwdUfricUdu7N7WD0jBElVPLYAP7cA+dPFuntify3IvZwPbmfKDfY+2ixYrOGQcNc3xjWM
DajRnOFnyy2Hi/gHJ3Req1V1LqKRzyAkOLyzV1SaOtLgnYpTYQc2JIHtCfOS+lh1CkWzkL1gH97D
QMrXCzP3ylJ91Q5NUg/zEgrE/IPRotizah3c0A1lxQ4DkTB0+gtm8XdKykMkXm1HE1mKt/BVFOQu
RkUx6zQf8Vm0Ko7oOvqQZXTwblZD5rq3Sta7JmNgHcd0qmHFCxWPDQQqIh67s1Kx1kiGTDGXB+Qh
olWlyqfqNNfogFS4S19CD1djsoJKpqTpt2OVq8ZG7sf4MNPrrnBJ0/WZf68ABeD7qHADaqVNAZDY
1LyattwZhNusHK1VvSIrR3ZujcrGiVVikoGrEREUDdX+GCW8GcD1lk0brlUPNDMf+oVkRAkrq6zi
v1L8jXGYWLjJ4su8RVsLiSFm994Rbfv5FeSQf5NV/uUWO3hzVtusyPtpQLbVc1Ly/apgdj9g81xe
hDGk1Uwnbc/ms/kDD++fCilpYtLVldNNCTtNPrvMoR9xVCvNoNK9t2d+7rFfxxUadk/HjWpfKAUB
ADmKuPT3xc67Tn4FQo/JibsPtSnkX1Y1hJx6o5lu0p0TH6IVhnx55QAePyq8BYJGAa2CsZa0Stel
6WlR6UFAUteT1NduuQHOirXn6HAL1i5w/MyUyx82Za2CSlBY66qarHYUh+tAQZwFeo+EIPZaKNso
LCARazJTXJsM4QgewXGoMPnX3yDkbwsWG/tGQf/XK2g+o2h4srp7vbqRB4ek2eGE3strnWYlqaAn
IKVOxZhzSAezKxL8diCNbfBRkqUx/5uKexcl76L55YvaxadspTjm1KZhpehCEMUL8lkQKBlX9FAK
FSZ0LVp4+u0tlJjrNnn8VtsdFUq/VqOPhFyLOWX/Jpuho0L9v00OR73BTJ4QXzfhCNJqA6iNeGAh
727w85ekYlf4ohe+kGugB7cwoVMSCgHSUBDbt4NZU9Ku5DZD/XlIOlwGJcW4AYgJn6XKHQv/PRW9
+ug/YhlZbMMK4DZQk+z+EChWV+AuMi6kZXM+nW0B80v7n58IcCyQaqzw3k5CyTcPxawzMz76bM9L
CIfcbqHdI7+Etq4peUetdz2qpTVW0a0A3sWlL7YtdJcLh6a9Ptu6/Mf2V2WXtDZFj4ry3pOfnREK
fkpEOkLbTUHWqHd6YszIFkUkDLG74ac9nSX9NkUrXeMSdRmVytLSnU4hT1n8MFYhFy4I10jZoW6+
krvHKbISXYVTc7toDRCJWEGpvyrr0GgJbxKXDsI4wfH+8DxqdFb3NY0hn916Y/kiw31xr1PwBl+k
Oa74SV5K4LhCJQ8De5pkvpuj4d+nGieMLi9YOv1I4WRugomuXfVwgWeQcjwOd3nPDu8xcE+dkfIA
CfZVEXgwraaq9EwOgcc/+MjvO5ziL5LD1EIGmRxUiE27AS3WTydy4G/zhWkZHk+B2gN6XBPypeYu
XaBsJ0lXHPHx0qP0nF8lprqQbfR6MVN1xK3TwWZbkFIrvbfIkdKCCWkdAXV1caJQL9EnK/CxZma8
9EnAk/pFPqyDbTN2n2G1Eo3WSZveo6JK/9DfPmgfCgE1YJhKi66jM8pLaUNjp0nS82A224K8WISQ
lB7Ln5goTwGDqGzef0wz5HNWYykhhVDIJapGK/4hAOrBry1IMN1D6do6w/Gpy6jqyRkBEwhdi0aP
whmUEVodO0D1hldGuNqX/PpyEkeEZNybJc/+lBFEAouPrxDpsy41CnzYV6gQvnz+s8Y8GUOKGDur
y3F/h0cG7wn2ZFEOUg6m5a+8nJckV+BMhwqQ4ZvNAQhSqbIYIjGMavagILGIig+qlcB8DDsvxlbV
mBuM7FwowYISpRz44ASuWsFA4/tkCBF4SXuDQ0MNNd1NsU3B2EcY2dsRHvIFC02oOKHZjhLYQyLt
ANhtLdE4YXV1ie70JLp/nPXYqk5qXFMsOj/1i/PGiw6udY/+eWtcflAKKiQHLNugSqihl9ggj0UH
ZhXOMuyzeeUotGGn7JEoJZvOqR62y3L3/VCO2vLYAcf+CwQe+BubV0gbMpXPmXxvuqJ8v+YvRajr
m3KIa7oCpQHhtFYKupEZ5cmnKXsK8SkvDNvEvceaThrcpHkGIV+FGsD7+319/H+ubvoYswJlEerT
6upDgyyxqmn9L1T1UNL2uaMJ94BNYDwj//hQX9VKhcqITLzpPjhQFao5qf+moDbz564aWU1dGDEu
GyXItHeT2sI0qUtmS6RUJ49JVI5JvlCAHzNvqC84JmF+awuYIuhIzxZm62dj7o9J0lX+wxcSpEn0
vzB6egvecEYXcGxWVqW5qaCf+tVv4utwoj06BjhkXvZjZPwwVKfPFiv81ntCA5a0+rMpthUUl/Z/
UUiguo8FzdcbAndCSQ+HDOlRZR/52kwRsAS5GTRy8ztTE5JW9r7KSy2WC3K2hexdKR+GwpEkJxwr
Lo5JtsCn4Xgy3/N74/GTy+6Y6h+4zBfTeojpYMspn3olVt1dqFc/IGCmnNm8wsvnSdmhpLqu+V1x
II5VJ6WLZAAV8AWtlHFMiHPQ5V9T9gWdqpdDZ1l6hgVyxYx7jWJF0RQsJHzejfKIvQGCqc+hdwV4
vrk66Vs6bx0B53cOWHYuaHndZM6KEkQxtgic+0UuY9Q9JtqQ6YvcWcW80GeojFuN+ctjt23bLGta
Pi6M5z3sU9/UsZW4mdZ6s1ePd7vT9Pvdg4WZLDCfOcrr0Tt5yjJZT/JNSPKpiiXSDguuLrHFZL5u
NS4GKIV2/LEB/ISctHKKJKCrbXoMRI3uRgIKVxmoSkY9lCOJMooycxli5TgUcaAKLf5tFMB8QnLQ
2VufE6Cn2zKPWnTRYRkn0643UAFlI4CLO3EjZg6xpn7ZGQx/NtGPH4PgD3zvYglGxNF0VKiTnPTU
lk4xpmULQ9z7b8ZaL1SzOl8HYxmmjxtKnEdH/79+0YwrsJyWl6fLh26axcM72sE+mI6hmI2Ee9u4
6Fk8+Ys4obGl45pDAWMMIPtmdxtcCkcKQ3MOCsA89Ikc4Pr1pzRnZM1QgbjhcLlimrAjsyT3EKxy
aBkOQEvWW1Cj8EvAwjkYvRpiOhjtivW0AQa8kqMtE/At+jWKpasFbqF0TDVtr90Qk3+w59dFkNwx
PBycrawmASwYc0XjfdWNrd4m3CDBWn8Zlhu2/JiV2c2tieVEPQi2O8pmHkqicdu0/Wtsisnnj1hK
bCQbteXu+Gw71K9XAwTzZUWkLVVuC3BjcRRdgJNgdzfvoJ1QdVczNXzqvJbbgH/leIvpN9lFX4Sr
GNglExWzDiFbgZlB1esQUrK/cfYLbGQtr1UZHbeRM7unqmTDbQ1fJKAOyDnG8kvUixu4/jrQMzJ8
TNplWGh3CxFgh91rgvqc6NE+doHCyqs/bp88Q/lAnoNXRDbuGqpMuMXZHG4kyt+IpuQqRe7IoU/e
UkFWB0XyXYATLRImc5efF/B9mGPbb8A/D8WNEn43evVT4TTm9us0CCWbDOQMYofdna0rPg9e3K5W
Da3g2O511Fe+cHNZ22E1gwFtlKaOwMIeqHwcJ6DjxGEDq1nfgumZ0TbN1+pHkVZ6qcKzb5SV+96+
1BpH+HlSYPriwwbJ+gJUOh3YbJgvOaf0yL2Qj2DDR7cIcQoCFV/Stq97d7K8NpxqTVdHPo4wTypo
9CAJmg5gfRaB2SUImOwGjC6UjzlNO3rcacsbfB7j4bnk0oXLsyc2tCVn7JtyKljT58bBsexjgMmr
5qkwuGQbU0YXiWTY41goqML+sytXJ3DXk0QQsN7hhip31x9LNycKg7r26C6x4ZZCy1vNs5GCbSC4
4Ts2OnDiW3jxPH/u42N2OfbwPTVG2sYqWcsK2Ryp7D4TvosgAn65JHaghA3F8Wd+MkodO9OdTxdj
ibZ3Zww7/so4Ex+7+vm9yQTIfpL4PuqWaJIhJJTycjFzOWYlLiL3JFc3jwOqqrrZqg6Yn3KoWxM0
c3pAVlsmsZ1m5L+GGiSC7El8xzto/4HwptBJs90bFNYbJul6lNDuRbBzJ49Pm5T40NDq5dlAyepc
Xv85M7NhXpTJIqrR4aHQ4k+E7wxmGFh4tjjWIz2RzGN/t2/vibQojyZ5dqIQ1AEQt35VbSP1MKr7
xT32sSsVgIV4voMdORSsekU1l0T2HaAJ22R9tYKNumNaxhrPMqysYPhHM+TpcXGhyftoHC/x1YrW
rMwFgcKSNb2TZcoaGI3Ge0KMmf5oHs88TuR2da0jAI7K34G/tP6xZDurcQwZGAKsJT6/miqMzxrv
Pitdt7veU7P6ylDQajBb+s3YE92BwHpsfqircsLp+tK05qCHe2sUEN7WuQZ19EygW/kupkEm+5ec
FC6725BmhP0H8O1grkrH9tYG3xA2ba8UtCMDy6LBPq7iNV+Wt6xZr0KM5rqOfoScG7Vo2n5WiTB8
rA2G+zB+674mcrbJVzKQ+HU8Ly12E8j6Kw87zB4WfB+Yq8sVvxkZdwl9hRkk3ATFY/oh9d8V9s7K
qKUXyyOC4RBhYtHq3v/QqnyF0x3KhrldKumUkL/ow1m0aj9r2pIDNQC8W6JbWC4/L2oDkGby1arw
bEUYs7xsUOUSjCGkDo1MyVLn1JOddDRj5BVApVCnsBkdwnn4+rk/S53pwu4M+i77ZWzdpgEgv6TN
AFPLXLC63Rby6Uxu0IPy2A+gFGcJ4F07YAurNgIkrYHYIh3s+KkKmAJrGsbEoIMY6RZUI9CKzYIZ
5og/xbdgYRVEQHaQhWB74nhdULLCt7IOoLj4fbeAVxyH1gN/bDGUY78LJFzcTEUSjzmkmRbVY9Sq
zA2Ft1G7NeoU7/iLKvkN5IzQj8C8z/HGbVwjMAOjK+HhjHUMMIQn8CmQBJhcWykSRbwcI5B7Q7jL
jRqxwXlhSWPW0rzvDifZcyELbK38V+rcrAlj2BAsbsONZXa2n8Z7c/3CcdIcQHVcdol0wsjqxxgq
FPiPhcwkainACOE4qj6X1JrkSmhWpjyrapq5Gq/TQZmr19oV43Qed4gywFpJIdzOz6DU3T/Fsxnm
3O2Rj7z5mv+T6eMBzFiGmyAbYi8yabAHrtmZYSxLzwVUEhNlmvoSffNC4cA2x7OefJtTejrRqbtg
FCvmGvVBY84/lsc3U55w0HS2MyW4bv0JXJEI7iRWUHCPepZvQNqGClU0ddJ7hRq+ncckbgnVLyXt
6lafWELr9d65Dyxsj44m2abC+S6lhGCRiSWRFt8Z4rcAx4pd8Gk5MQT+heC69lGROp2DUSnR045w
BuGaq0Vr8UtYSc+Kg2iICy4GqCfazTtXfWvYZ4HmqxEHY1E8zC+4NuG1g8+eSlqD4J2pQmY7KOes
/ggdW4I7SIjLiJlq3FLAZ0mCNc1/Z7gUou0DzMJhMMtRkMlfUK13OVSI/xNEr8M7Tq7J3Thk6Jvd
BnRvH92pY0Vhjkmo5hcLlMFJdynpC2OzKBjvr6fnFPzvXAo+rSI0Xz6GFlQSa7nZ6ZrTkn9XzjDA
wRL9QmAbFfxMw6Pgy+WCFnJrg2pha77I7X9bN8ZSxqAU/qHW5E/0Vr6E4izQd5joLSGs6kVo0nhm
+yfkDDwPT6xR15RBszInxSeZ+wmJ7Kj2RfCQm5VAoxxNhmY49eEC4vxehmwjgUKo6y4KysIRo34J
ioJpQB+g0hkgEbLYMzympf40DereaUXej9F1g3YNO9g1TSWR0Qax/ho54abpcRrneswJKvxteEpV
gSvjIiwEjAj4ai6pTDOyFlzWMac1eyOMD+hcH1ivIFZGQwRQ/7hJG3sW+AishyCEgg/g7c8nRsWG
ULn4/e1tVx0nM0JydQJX2cdVZGbddNuOEpCKqzwsGQjzCu+UYC71nq1+3Y11JYg12bEvsiHEut0/
OthfQr9iWQv8Xv2jtjEpbKTKtJexChe3Vzz7PV6HUH0J/9RjnF7EpTp0JLYcXW5PDaBLmLkNVm7M
2hkI64CtAldqXBTNjg3lOrSIb2EIJDZYanq5rsX17rxJS2MahWtfZy+/j/lK91NkBXGghHBV3N8s
xL6OnuS49Kk2Djy3HFswIX6TdMadeEoYLys/Sx1X171cqj8kj6amgQf5xiHarbMdqPcCWHJXsA2+
7Znm8sf0COKcM8MflhMuT48il8GxP1FpBKtGsGYiL3qTH73mJfiJmSdjDvNw2SbpHhpjVSrN9/3J
pMP+abTfjxiupwTrT+kTWHfYPNJFdOdyNzyqQ8Dz5BB2MxCmp3S7hxy/E9KgeSJN7fM8Ctr6HUrN
IxaUbN/cCXdYxDEhO2BQftQejRLWkJ8QL/U7M5+YqnLv3/6EQS6A97A6Vxo36+nrrfCIkmfycHj+
BEyO0EOycM1RqlXWq1Vc1iU+zzb1FkM/UYzRPueclwDlowUPGhi6lq5LjlX+WzbHO7030Nt4V1+3
rOxDfaxKfi++f0bTIFBMj++edfvAkSLvwU+FzWmLL/mw/aA9qaBVUpqCakWiQeeIMxexnVFfQyKN
eJnbuweZhFM1OVRC9AOCBQ6R0oV+XfHbr+60QqwdHywpiqmLfJSE/8zlLA+U/Y6iVAAXkS26ReNQ
NmaZXABJF4maIZwTKLECZh53csqwY4+etEorE0/injQCP/0XrrY8RIMFEABLznG3tPVTLmE8cScJ
S75UaWWY+W7RVStU0wpFEuUrfQEMfdLoCYcBR11Y4Tysa/cHLdtarOxo9b0+aFFF38jMN0BUI2Nh
V8+F4EN04LBGHaTC4Ea22NbQQhJFFHxGEUv51IQHJPxm4mV7eKQlU446PuQKlqUR0eIXxnw2ayUh
mDxMqgXzlPkwufNCvtahJ/iTEipeiBfHdSmoOyEhjP6G5NCayOiDUTT4hfFHbZyDRQTkQM5YHWoL
ZQgtogApaBfntwg9t1hK8V6eKOJ44Mt6aUi6iLUvCx4Vw+jDkdHy9L/HhsUjF621cJwMfbFWk/zX
qfo02YDBM9Uuvs23nUmWvBPPCYQHBf/CZvNSM684DCFxyu4UxUPblcAZhQq2L3og2m0YjiJg+tGY
EzqurcQpkQCEZfdq9cUyRTLVc6hpuDhR2xE9KyGT/XNMPsXTYCsCDeLqIUMBO9+NKhAfMZnnphZ+
mt64lW9JZlfZxE9dTyQ7BRJTzDNumzItmsU0xvqQFjYjQqotEX/+EseWrOZxiMmRBf/ZJ9C7Ip6w
Zu2HzzpgmK1T/1VrtGNAqFWlEnF9B5UvZqmDPOHli19mmturSMaRfr9ogxyhJLjQqxKjFEbdLXVr
6S4Bsg0h9t2phcU9wE8ze0AMXMXXO+VXUKv1OxMRR+YKUAH7eZPhaSKCJovnW3dca5idwU6LwFs6
LIZ0gAJMPYr5tuYxUKF/qwJa3oJ07wfXcS9Bg20kKwbT8jkJsho1Z16v/rNhYLQuwAp2IZxEU+aB
Hbu4IVWNHhujH5DgrIrdHO6Pbyvwo5XrDuiUIeA4GSC98sJTMnAvQyxGIClLS162IAh6QR68VAom
YtwY2VSLPnrQMvZGRMCWZ3ChWCRbll7enG0zksOtoeQT7DftHiwG159ZwZc9l7ZLSuMvOC++LtPO
QUgdxsD1jmN5kbefYlCVepy587wxv+RbEo1HklIlOwevx+1gnT/oWdZdwc6odnpBWv+Mh2Hb6tI0
qPUhqVN58k05/lXXWLeM6MH5c4xuKq+kRU1OxCgLjdQ4qc1E6Cx3fZJFysyCnsUo7LoMvGnnH4B3
A3hIo0KoshIqRYhHprII71AVXCVF/rVuY07cVp3ffdtQyCZCtY6yVaCHxnEQ1xGo0++39iXG5i/D
immpQSRZRCzfQPmzC1LEdzPev3RnYtz4ojKaPwnY0xtYCc82b+1z9xcR0PCcyos0NFOZCBMURiWW
p2Ur5KNgXahQ82DrAk7Oy2hXkdNmCBrP5tAVz0T4u4LtOX5NK+DCO5aDKiklZB1ISHNvaWtI4cVv
SGosuiv9VaxdgBYxYohUCmYAKb5DogZwCNHezzWdfkpwclAmaB1cL1Qj2EyUyNbeiyIpQWdWGqcI
1Ci1D7VlGAQBD5de2Ouer4iXMbbJsp27zkskwa/bNDaXqbmLXtLzqVX7LOyDcTEyDrBmyzeSW4a9
XkD7QP3lOGil6Sf1GqRVzsUz8+OnX1ZO7zrkst0HDqGMzlm/h8Zlc81fqnOQgKZMb1hfNLzWQwJn
HSyM19XuKf+4Knc3Io80+PvF5WKZz8UzvIoQMtpaaXL/lhm6AGKP06CQwCI1FfJ42VofIB+3ebwi
/TfDmMhE1sGrw8NHSada9hPD7Rfop1GmRmTiJGXSxYT1PCQax55QbqmHrtxrELSKpU3D/FekRBox
84QD0qQZPujwmk56OOGSHMVwqxvR8GbYTqhR/Pi86nNaY0iRbEI3AOPgc6U3lgLOVTl7rsCy8tI+
smavVKC42SjWk+4ny/Se83Bgez5SvcMhKcitb7hx9LHjlwg2EMTmuMi/8im8H+NFJSfynlFbA9mB
5gqY4NzUc1lSkI//q8mzwi4/Pyu5my75ortJ7P10gz+aRCv6j5jW87odvWgvXCQansZe2qyfrevb
KG30obiScKgsiNu9zHuVAzLNVcg0ge+zE7ab2K3QdyN4pO7xtnNlqW8kMHQxVSOY+ik8IordJ9Ab
btlbd/UXp+3T9f2Vm0Ydva4Q+YApqbzkBybUYiGvfbEqA/mz4TFVnTa+rYtiCda895nGOoD2gMlh
mU4KSbLMu7x0Eefr+baP2+tFz6e1WiVJ8Ls/K6wMxA8hWBAVs1kPdHcMuLqG4Mt4/zJziXvMmgtq
WIuxtN6N3R77wqWB0bDx4x2eA035DJs1xHyGERe7zA4T4/HYSJlWv3gvTbmxvCOkawHLYx/GZ9oF
1jtASbHGqVUt/VFT7lyFeq1cqz6JXZYrYLonlwA/Mr/uIdmH5lntmAR/2LNtmrjjuikoe/KoNM05
okMrKcFRQTj8CjO/U5MaxHQNmsyCmZidrU+WcE5tkUVFKxZncUpBA1+4CTikiecqB1e44DOS1tBm
J0S4My5f5QjjaVcGkNsb1VIUtd1N9N/HC7ARZb9jhFJ1KmVua+DdoTjf8r/R+XcZ9Gng5NX/tyNS
xYJRrbeVl44s7qCBe8CwcfIaF35NckOeKzM/SvPfATACZn2bP+iTQCg2oFd/Iabh+Wd+YDmDhAQa
E6uuFY6ttr7N8PNhM4r2g+ryWfxMizxg15e3Xn6twZMVAAFhBMxlI0DLZWrzxVkECY66IwGgFLts
FQlPevFn2L3KAlVltGJ/PHmbs43kwzqCRR7fNXCugpEnXauaOon13bPqPWfcH9npn09Q7AuGvCii
HZjtHepZ/DxNY+7sHEmIjWJKxcfKl/XUMfKsrZb9vG4qHhdqeNhcHj571J/N2uTxm7HGl30SIeB1
JYxawwaiAUQ50BEmUFUYeVuDns0302U68SdMXWm2LVzjOd6j+3N1CHfgoUV4jJsJepl88vXDYUx1
x123yZpC0NIUQttuiQj+voUPUCiFIMiltoFZayB857thGHBaWvxHAQTkYMJS/svkiZmQTWaPFDEh
ZTBCURozPxx8MAlYHHAxT2/3hOhM5kAJ9kAOQ67tV1Ph+n+qbaXYdHRu9IpVGsiL0U6GfbBFS6tE
2vwsO1Y0mMf4PH88drmd6eZJ1+Tz129S7Pb2tgsxtoauXKYE1Rn2t82G8veX+iaCmasd+DcDS9aE
20B4jeluplpqqDmRoQoYIV8uvi+SzYngW/D4hyU7VFrOhvDwsGWu0tzrTVrnVTSH6bvlxZ2W2Mxp
0CSvncdN57+fC6EyPYuR56RbaXRPf2f56em/F08eaHifPhmWSFJt/EBhJj0F6kLQO+lraceWlBD3
zFZ6B7phUQDb/mFgSWa1nTzoiGZUo/cDJb6cQ+BeorgzE0RqlUV12jX+vyTSJGhUDKSfxY5NMPig
PDLchSh8S8mKvtAspGGCdfo7bee6yvb57DR1LK0x2ndNJFywZFKDXHbsNZIOoTIzYaE6ku0QIx1q
zEdr8Ibr9y/aoT0z1XLIeEestXxEk7xFl3xVQOagG7Rb8yNNGMH0XWrhnKeEL9gUCx7Ye2WL5nW6
ZvscItu/ZHu3ytgQNYDPyFohf2EvlgStHMYJiAsxD1zhXt5zCacfBe3kwutf78lAji0hyye34lwu
58WurPHa20RxAIJtRSZv7uSh4ZIovkVnwpJyHCkae7dNz90oy2lX9B1OKwpamN5ZCHBUuAL9Ox6r
ukaoXBgUKxpwksG2qh9+nbZzJQHcHNsvCed+0Y7p/zdJHsF1QQW76tMI5tZh41mWAgKA3MNlPNCc
Je202eVU4khGnXfsciFgSJN7WoA6cOXmiLKGf3VP6xmXUc5pKQj+PK6PVE1hdRV+HjJyZg4Max2u
imdPLhQmvzcuFFba/xBnYxwk40+MH2x1d3szHmLjSAiIAlTPbQbS6h0t0jisc/JMJBPA8EXNEVQU
EYLGu+eIPt2BQjVHh37pcsUTUFeKKK1gADSZEsA1WXxVR8ij0QD6vL7VW4aMZs2aFse+0Ujb0Yfl
I2vbKalWEQyd2VRElPkT7jT7xtWD+l89vOq3C/MD0XhxuSWcmfh8m7/s9SfXDMTNx+yt/Qs7qIfl
P2ET6JrtAULyHHde4paK7hni/+/5PwAq8TlgFWLwwKuLJoqr9EEyakc5Q+1FftSVKCA8etbEUflB
nkDl6Z2LfRGCO79VSKxIIqhFVc42dzjGvxGE7c3LrLAHVKn+fM4e80fvpWvHf4aVLHDtqtSb4DYs
2+hJdJPV3AQORq662DUzNtMceMqulH4/2SxGoTkJQhQUiAXbZ/Hj7fFZB6NJwnnBIVc4dMYwdVrL
nb8EU7Pyrro8wpPix0dcker5is10HREra5jAr2I9Xi/DL7w5e8TJntj7eRrmYijBKOud8QyrivEd
Yg4jUmrz7I+VoeMRyDmmx2AjuCikcnLk3kLHEhPpxV2ZFUFGPFc4mhZx2h6TKiu9bvUAJdSYX9n8
SFNVFfRV3hnxu+wwiDE5yd6np5OHu/rmOO2QR1XPnID4vAgTkRDg7ykqAeDfnF8M2+Xdsnvskfog
ZwIjW7Sp5uCALeSUBZ5CLN7MUP8R5PKQiDQpOH4LUmZ1pVyxylbWbSAmtO+AJu4xkxKfQcI4l2oD
sH0QDurzdvarwKS7bx4qXkUYFUBJT9pUy70unF68Ga8bX7CLY+/qcCFU12Vr3YQGTqNJFWsS0WJw
YwnTC7HmyxbbnRSfWjYnf8n04vQQgK6o7OThJxGKK6mvijVzXnNX5nbfkWZPD2+fYY/FmdBq17I8
ptmL2Zz9K/SuYoOqEHv++0mSIhCJDYvyduNA5M9ftg0T/+Z0WKsDZw78iQrr3KbnkUa2+qwYvKpC
eq3igh3VHFAyT0zZhzY/2MmrvAsDMirzdicVofQkrRpUvkNVEgGapre5sp9Xgus+Ji9apSwMm1o+
8hjdef3PCTkJVMXNekLFUyg1IdJladRMAVa9guYhzC+4F7TloaHr4KBOnkIECA2O7aG4BgP3KrMA
acLLEo9uAbWE9JORp6QXmPHYtpNE0dJR72FBo1JnIBJ98DQ863Vj7TSYyqpaPLS5TQuyy4igVT3w
XB9iBwh/2+YYkJioBeawygeiCL6KCkQYNk9nXNDNr7tb6SmprmtwnmWwvLUS9+GFuOP0KHZEpD58
E7/ZgJPcxHIao4LN4f/rrZ8eo+rHWw1XdcDN4Ujao3C2/9ltTjJfhYqKQ6uD+8dzBCRp3QtUiVLF
R4akScUXkf+cn5ysaHT4g8/79jpQrgcxtcEo/AsGDAAIGZBIylOI0t0NE3o0VMxoJshhZ89llNjg
WZng4ELVPufj1asKKQx7/yK47TlHzS1rAwV8K+so7XB1Z8XOneduz2+4MlpcrYvlDtjJXR34kH0S
FVCMruMunw85Z5Bz1TNppqOpP/v17+QmU10yetm7MnXDt94vcb4Y8ACijxNXSIAsm+uuro6fWLOT
FFOCJ3fGicPiybISg2XhQrKBIRn0Eg5cYHy7sFVMNVpAroiPnRApe5erQtKElHE45qirSBFXEfob
0SkKBdFYrHnsrJu+dGplvJEvN66GKLMzzB9idH8Roe2YtKpba0mqOoolWKBnD97vEHkXDS87LyQ5
Y548xnakXOyE5L2S6zMPaO9gIdORWRVhC7vnF04bHdJdWs/qccKzG07H1eSgrn6KXeduvF2UZByZ
mqbtPw0CdtogxXh/aVLwYfr6lTq+6MGaej8NLjAQ651tYTiCHVIlGkv5/6UesRM3DWuNgQD52LzF
/IrOxIq1Ufy41M2UztASRjiE03wdVu4ZBQTO5PXLf38KlIUrgbChxxP4700BkDhUqQK9bto6+EDP
KfbklBaMy5SYxFMeefQGJm+Q0Bz8ybPLooSh45mtFRbBUsuPHjkkiD8FyKGJe6nlAj3OliHr01vh
Xi+ZhbMT5Gjm54XSi26I8DmQJtnTGNJfRBHdn+QGwkXDSp6vrKDWSq2tLrmT5ShlfFhf3kDAVbeN
+84yLRz7HQ6CfXWrz4t1En0LRzfcqnjdEGts7DhsOWuaM//+1pNTJqq7rilhSBsWKRdCz9M/xwPn
EoEJNyzQvi/iuDH6CLaXL7uwoM1/1fzIy5ci3M5kQGyc88YGxklSlKIf+X+7BwQxQC6NQqt0Cn6I
pPopWFPfgzUKw/LmifxojoUPsXIKMRCg536mEtsN/gWnysxz3nL1uGJXol9NxYIpojyf4YDgcBbm
CmUBzMzXVQl2iWF3u1FBlufv6djGu4Irs4AuEfxQC0ds8qMhKAsLgfNpK58rMzxyy74C1gIM4GYp
y/bpOuPchfXQU2EDljX0p3kEgE8Pi+Lt5xdeHmNyNNF7C/BVrqTWflGwYqQ/wXZZURXxu6mmfEFV
cflL0UpbirqNTNo+hxalLL2AQGE4eTl5g8IprqQPpzl2fsAqOM3heGB+XO4/45+LoHmrzRp2/KEk
NUgMJ34FtD5e2yPlz1K9QJeQI/Eaidrsn8M6k13bwymCdbYR730jWVpH0iAWt5MxqsMiHO8wRnk2
TPbFqiKFheZjRQ5m494YnQy9U3dZ0E0KS63H1Qfn2sjRw0HFGKpQ/TqhF/CKETcxX6i5zp4VJaR3
aJukOEmXxVnul5bmR5cnKuuA2wBHCy2692F1cSMCdHvZp87rJe1EYktA+oqBS4xZl8D+E/OudzRf
7UhQl6yCbq4lvoLgHkBBXGgMk/9nIPji0spHEo11e6cOZOMx31Ui3n95bdKDSsKUFVtTu8+bbuAt
ClNmwi7IZnmreULmUtaJ78Trwdihr5VcBPUD3UhPdZSoalbMRT8nD236GOwdQ+G/npWTu5CV6sBk
zxXHdf0EP9/OE/kppfTyRshyqvL1VKpDOAbIHvFJ1uTvQtvGkwphegaOLcz0p87MNkm1GURkkVYt
dyldbM7354t2ANJqNjnfM8IKDQv2Knkv2y4OFg2QvyriZjU/uqvkImbqBGww8RQlq+zj86G2//DE
n7tFXPLvwHXsg0NHHoqR7mSLeZeAXJ2a/R5vU9b/NNhsMHTHr5jf/y/a0oChzSXGc+C4s6xb5DrA
KNbO6HDRT0TPyaWEvy6w1AUzIT+nhk73OEwGUPTBYyuyA4wHXb9Z/IS2Kj3Jk0tTxM7Ahyo2Byfy
H29ixyBK5D6tJlcLkullVV+g3sxqVyIliXxxz2FgJiGnrpHXN/7WJ5r1aK5aOd9vjDyG83niZgFy
2uO57hqJif7HC1zTkZZwNGg8OQzqU46l9XyS1nyWhnpwU3TXDGGNATjEKqNgKp6nv6au+u2etWtm
U9R3wKacTNEacK830ktoB0HF1Ruu/N/aak30QekyJxdNuDW31pODZIttIyqjEeNuByj4uCL3Dzqk
zQDinSa+yeCx6tG7N04DVqJ2Hgk389T1f0nPStGa0GNohtH+yR6upMz2Pxs29M2bvcYUKPod2GVy
7g8pAphymRyozCbz8N6caI0n5cc/NXgEmUVd3u0WFZayc2Cl6Lg3XH7IgBXMq6ct21u3Xm2zlrwx
JuNKqfy05SMhnkouOTokSesEyC8k5T+z4zgK3ODDygUEjsG/BeSLqj/7MgcXy1VBI7dE3GR2Lei4
6CeA7ZopLpeKQjiBiE3nMZF1CAR1yDFFjrYZLtj94wCujix6qgPJz5FIK9dGZHZ1RwZ02vmGyeyf
ChYp9VFKhS3C/OR05xJe5P4tD05yr51l6EXEswY/BdHZvh1GXc1fnZQIhIG64FuIgxJtRGAkoqHn
G3uSRbpyi1GcKAwpZfk7ZApLGT/PYXLUNOY3g5y7FQyPOog6M13HnH5wx0vfIkm0BXnB8dNAImQJ
NX3xRGCMQtnjcLIdy9XvRLRIrUGQmCJtgMfS4U72CotdaI0X+n3Q7gNKlcYMaMdG63Yn41ZcPNRK
s+8AU+rQ7SflsEqNDCRjxmEm+3saBDQ4gQflsKDKvMTMsVcLfCHewPUsjaCEelD4r1Ccup2xH2wc
WToE2Modc7CXrhdezbxq9gAqgetOnkTYjURwYja9sxLD7qK3lTkugmvSidJ9CRSdCmt/oe1ezw8w
ppzQ2Owl6dxgmxcE+pnD4KpqqG8hxYigfdBd/CQJG2a/96tXN9Z+0rM9jul+cQ27Xd0xnj4VosCY
7OCDbc3wyMgErc6HqkzLKeJcsS95FN6VokPG0cjjqk9BhMeSZyG2KT2XeODLgT0yDH/UtvNc8Wwp
ESV0F8pCciQq8EqVFUVOIxmIgOL6etTxD2iuVSNox2IVWxT8KB/Mqn36y9YLn5EhOr1YUhjkfHjm
Yo0yY6IN7sRTrdi7Z6Bvh1OgAoxKG/ZBzAIXhBSZRYPXRKzyMVChnlWKpXmppp6j4w40ir0ELc35
cobr2ChgJ1Sh47u2JU9ufNNd11esRLe49meYVOKDOlFLQqi4LVxeeHSlK7S5GnEyxK8/EBCKkNWo
+8zdaSoi36Np3JomFwhBtibGjWhucc+Gb472j0a9s2bLhG/q/HzRWTYXu2MtL5heHpVZABBww3Fo
PR/w07YPnmR4Wx+Kuj08lKl+zjT++9pyOvmSEW3SRtkkSWQ5FWXn5eSroz5CLHPHUfWVk8EeLL43
ug9NYqu39fhuBAD+sc4wjwTD5QXP09nYwwoTdqpA8ghmAHGhh7I55MqS8k4LPyMgxySUVP8SeA0Y
4D/d7AKDVPrN2dWjFzGt2JXsd88vGy+eRJG1DQJk0BXi6medFre//aaU1HW2NaMf+ifBFglJ/VZa
58P+Lhi2RnOjv94kjGuNm2P4Lp6MBG/bqj+IkepKHoASTjZLGG+oZGF1PAE8ErYs+4T7B+235Wj6
R0xBPvpeiqlbp7zzQqi7tUO7XwMpyYsUaBukO7F82Nl5fpJY/7UNlvRWb873GCGFbWSCgICtzkR1
hM4ligfRATtU8nBNeG8iLWkdUcYM3OaVk6no+ltXumZy3FgaJVLfGYwqvpBFvrrumuLjm0jo/v2x
Xj5qT9a/xk2jTWlA0HgYfKT1JWYZpvYoSD8nSrkbM0cD9qA1a3gk199zWepbDHH1BFggp/1rRLUw
FTJMutTCmLsdKBMlxmkvmKmPhzVtqOaxGEsX9tNBTrp9i82VXSp5G9q2Ig0SjJSsYs82LXpibI3r
lfZOU7Mtl6KwDnvZkb251JIZVFAJfETfD3M7Wq/hJ+St0oAL1xXyn4nniNmwaSiIhtGDKXjOLNCC
tbR2EuxbaDezl++Bbs5qZvGkm40p2X4mc6eYuivLJnAc583VQFDs1mfKsI3mjKdE5Anqgb8IuZZ6
8HDpMBK3rQEZt7eyGyFzzOCcuHDqwpVJWP5NA3Lh7opI+DDAFGEJ5X8CWFT8MM7iu/Q3ACJfsdb8
hjWVcVRGlXZX+1dN8gzkKF5+XQSZwuBExQI9ENDfva9t5krJxDf/H6i38GiXNMGnRXNywBkRUITn
24UOu6N/VG7/F2exjpw6FHK9av2tu7DIdRhi7iacRMR/D6NnRKVe5IgPQg4mxhNZ0EAl+iz/rajT
2bSJp45k+NxFY14D47JCE0qzXz3NoaDZlWWyM7V3wbYCUz2ODBLQ4bd3GCPPHxeFzPk3FHjm8jkv
Mib1/DTH/Ao/fZ0YqIXltz8aZ04tOKBs2iyeqvRDq8URMrLb9KfD99dLpvTQEgkexcnZPIlTxeZh
9QM0bWl8/TLhnjb+sN8Is1W/hkSb9Zbd3zQGX0I6VcTbM6IW3H4TfYfgn91GtfYlrfG99fRVfNNV
jmW4ltWeuRPSm7KVMXFYCRKmGQ90+2VYE5JIHGvbD23LpqoKl7r3POWivOiMLdBWF3Ur/8OhHTnG
YLh+r8xws5Hob3l7OuInyDCaDQik2o6V/tzq1I8lIqsVpSQ2+DRl8EPlgNx0/FYbZrcQlzVyun85
zMV/AG0biTnxYK9Oh33yPd1YBeDTpcAk67XeeYw+8zzvrzRnnvsSGPT1MC3FVBDtfnOY7sxKr6Ly
kG2Qw6SQF2tm8xycCIXGTqpSJ34scH5yvzD0/bU1GdNZSdB77KFIbvSepI4HoOuz3dyLvyGW2pqQ
dREnI90ygzZ5IczdG4VWXwxxfUpc0/4mnxN5IP6qVACegA8HWzL4ESUuka3AW7gwh7TJ26j5JfVS
Af0wUYZvhhzA7ABH93uA26hmpKuBvVAg1u6sq0EL/NlHrEVvGiEancnwkICKYIn3Nygz0m4jHgSb
ToSMXVc7bRW/z8NOVhINTaWBr0luZdExCh6ot1SLFPvwgmfz1EzYR7cOE+boR8/6PE2QyCRdPBkQ
VTblc3BAoBsiaZChoL6Bx89Ph0Wob6m+K9Sp8v9jOR33wfe1RBGOwy5+LOKbAdzqD8AOoaXgYDwm
dK9RKanHvCY1ggT0nk94HmYkGLvTEfufVowFXdum7CGQLee2q2Qk5HHsA9btTsMcvWvp7Vwsd6AK
HE1h3DR9LM8vfsPuRtQK58c4HTufZyncehAcjJCCCn42u1y5z0XK5HKzWj15A4TVtKruubkIkqVX
1D8CyckcYxl2u+oMeM42pcY94UI7rFk50Ne9sq8ekk4Rs4QSTAh1qKiA62e3EXqd2KzlL26oAXbk
WRpGRBfnmXWF0uo5v2I4GSJk8iVystUryiuu4JNqZRPJVCadmPV+rK7vqe+YprZxcE5ajMEfq+gI
fJ5mpVIrM5X5v3mftO4K7alIpzDzCVTzwR5XNDNyO7Iig6E2hp43cQwTg261DEswaTslL7qgYcpY
y7hdjlDXNzsYAtQTFX5w2uaF16ZUmmZF1dD53oyd1N7FlPhECAct8RjMveZMKgyEsRgRWOo2LN7V
O7+MhO2PGbWv48F4EmKP2VfIrh9EUzJpcKTQn+SV0zy2iol1Fd2gh5wxnX1EzQ4otY1Aqk3yhNgA
USVlW48AeEW9/IKuy7Yggd+vRD2Cn8O4zDHDeLP9a44bkNDNqSWfM1wXzv6g5J9bcEEaP/xiXNa7
fhHkI4gp/gGa+Abvn0sOnU1rJ+QOAZnVIazeUlCRgCXnAPHXEVPq4mFDULFOxS21A0dARcwQR6ax
KYOzie+ZUZsjap12JcvFtftvBnVNyGkP+fK69iTUu4x40nuYKobqOG6J9m61OQ8d50OJ74hhoEXM
wFF5rvA27EuWISDo1uxvUQL9bZerJy4/0d5yQZqBwKg8VtxozYv/8GSJb/CnXNuGPffrbkbb3XWn
BI/29YMl2p+PJvss01rmD+E6eKhiIs1G8S2MthPzgRra0wYhiptXRDZp+uYxxHI9fy58ys8+nSh/
mSkc96SW2bnLN+YAVOiMur/ZppLSerAYLaNe/k7Piy1fQN892UCRTYKmlvV1cFPRxCW36s3k/kmr
Y//GZcY1elPSdK/4NEOe/4DyPDZlFzwK2ScDKGskNttyCaThOKqAEZ+7lEFp+KyEGInjXi8/AKOC
8mDiF+vawSNVZTl6a6p9+AEtJ11H83nOV+IqKav3NdyufAH4k8DNt3Zi5Gt5Ga4wmq5wCoVdX1H9
yiQrmCEL6DQ7dSyKoAuxDqicUsJUXrvJQctQRNO2QjuvP9AKE4TnzGfS/vU5+gcMomJdAjNeDl0P
5cDbQuyi1LqQJzP7o0V7NSnkQVm5s/n0fLtLZYoUz3tZP6dNwsLJAlySkfH27S5UY2kajIuuMnYI
z8GO+AO9LdjSnu4LQBVM8zj9cop6L+KXGtiJxB6AxEwWTXIFMRJ9cz3eAAR5PI8YxwGJVFyh5uOo
RtHFbepNqy8scvwuw4iPJbEynI8zo1e8pDYujQl26OFt5dnAgF0t5IxFAD/+bF/HX8K+Tnl6r7D4
eCq0YIc3W4kca9SXsJFonf/HG9FfmcjYEuU1ySczCj88wnYQxNN1vQSJ+nAH16IdlIjm4PN9TJpk
4nVkpOzwVLJQhp+BKeQfHL4Pg0f0c7SZDSY8tgzOE4idEBAeS3X0SojhlDHrIQ0Q2OwpaCyobMwo
pzT2rr+ryJogxj+UEf7MdiwUiisVQAXzyJsAizC+gFR76KG9g9M0vAidwi7h4evU306SG4HJ7VLs
z5MPIyKGlXQic5hP6FkGreqZt/0LrqjN9wYitteXqjwfPLzmahSc5Y4Ni2m6ikJdV8LraUI+HnKX
56wj/3+yGYjxZwu+5oA7EgIGwpNBl+Xq+SBWQNeXSSks6HEKNl0ua2mQYxBBanDl9Jh6gwdCivzn
FObwCYa/LuY0JD5FrML65aVr4fVb0TelhdSRgcpl5kFxxwKKxGAv9ibyUc5sOCWBNqEqHM1abpRu
UGU00jX9xMKK9GDab4WeVnPiZKN6ApIVoWhHh7sluv6qQDY/S+izZ5jlBAFDPimjxL1xh/h1Syc+
bFvVCcibQKQk6Nu7BccY4cxet4M0I4swMp0j+ZAvEuNubc57W2ioiBVghhA0rlGFRoinad/lT2jZ
c8MY3sMVN1dAho4wSgsmUd1OItNtJywGvdGASEK1vjkLUpdx3gUAhn7bMMnFfGaMJX/K/Ark3ahG
D/Ns+FCR5/+vKgarzhDNXmN2X3un5g4KdiSRNCuzmPOrG8kIdmD94dnaskzGPtM0rzlNa8yrNuXF
w2HMO/iV6VvFob2qIP0lP3pp5KYLPG+tAyu64HwBhEl5eBbeOBYmhLUzc0iGqBGNE2RZ0H/uZ18a
zI3hrK68f0FkDfaqYc+pg6ZGnlthHYzqULtprUI0DnpbjZ6vrl92rbH1Xt6s8S3esBUNB5sNbUS8
N5n+ObcsCImqLNXyMeeb6oBFoBHI6YguiO0GvD0fcU03cH6ewNyXyyxvQONgT2dBHvBOf6gzZTnq
qTCHXyGIuQQ/ZvI0ZYYhkWydOjTxVreY5UPzoT3pVQfWJvRmM49Lw2Wl+2m9bd6zRLtMyxf2Ebnz
o/cebLrq348k4sQKkJcsoQn+Ae+/rSgd9wXYuvhn8ySahx/3Gz02vekwRQh0L89Gdx7rXT/Sottg
rzxCHp/JhnGqw52JNFQAbJwIIRsRIXl2NE3R9f133l7U4ThaTEH2DA1ipvTPXPkq997YN9Rw0258
yVWtQ+8c9rl5lJzHzL5qCUcuOY8BKwacoP/DeUUyr0Ekrv0i2UFVuc/AEon+xLd3//IQcx9FyfId
Bdgh/AbryyY7IIz7GfxQCOzD26dpuynrWNisVrSEJ6QhJJOSDn2QxvGTHahoJ0pV8OW07J7FWYR8
DGX3lMuthq3LMNc1686kUKBtN5p7bZUUAwwGtk39g+8ZLiZvDF6f+CVPZppKO6/HFeF98T0NvnK2
9Y6bGqwx/QHM+2iAxWVU5Ivi6gJ0x3dTL1PLij1bH3pObZkK6gEol5WsIEBV3qojFZZp4zuGRfJi
sRz7N1V5ypny+emSGG9LuRNVYqL8w1O1ClLB4CAUKsLynnpA9TtiJzJX6bu2Fu3iz6g1JdmAzNIU
EJGTKyWMRo2vQ+hpRsIRNZlHqNGr9ExUP50vemGSPx0hIGKIYET9KExgJ+mSWC4MQHIM3wNCNZua
iKKk4rNkYFc9VIpnHt5ulsrwssY98UO9rW0ofcHxCafYsuEvUph8KC3BNc6hew0GkDQ9S7odW5ya
JaomfWEcHH+6C2NhjJS7z3WvJj4RWNbI4w1vdvXgroSX6XS3B+iFLFfhQZPwFA3VMB4UtUTOc6y6
mJ2K1mM+ibv/esGflSd4g8Y86J/VmVMgxCViMoVXYvbq+AosfQV2g5wha65ktL//9lY4/p5M6qBC
4Z9iwszEbiKK4XglfKNt0yNKzFni03Y9T87318/m1SQn4p+BeHi9pYEWbYP2T/4xOhfocojwS0N2
mQKmP8DfBUFzeHM8/JXpIgGlLXJ0ro37bcf3MPbFKfVLbN4iGzVI4lUpKx4BF/ESwSwxCrCvAb7f
4HkbwyBV9c5vsz8NE366SgEVd0tKEdu7Q8S6Yw8ZkFg6kHQqgDqc3L6ljJ7PkV7yBBPYrjYIhueb
a92kVU1inERd0Ep579QkbL9iCIS2x88KbGVWWFFevBmUDV0ehnf6tnneGOHDipzQEGNAVNCEW3MD
WHKkvExFfeLKWxMkv6UdRFHMSA6xRpTP4t+c2pwPLEX0bBCDuUtJuxtYWPXrE4My24AF4H9xys57
lgauFXUydocX6UScoITmPTtXu9uwTung8m1xNccl5S/L4jJPHeVWhb6vmkxuhUh30Fv71qhxC5My
8Co+vf65G28MyfrJq4efdL8BBt3a/T1np0HwYnDUSAhRZtdCFg2Cczm1di8fO+g4CgcwXQBqGehC
I57O1iWFcS3nU/PITxkb1S9nipffkxM1Fw6zeQD8Hhsu0ouRXcAiiXL4tTszbA9rizw+NBdfAAtV
8L9E0ZZL1v5h0h6BMrvPN8pMQf4iuFi7zkvxepYHVHZU6NJdPk0Y5XBXfmTenPSm7tS1CfIDQEcm
tTjVSM2WOy/W9J3Zid9p5UCrmJdEzIY6JB25gYlm8Pgh6XRgGzMQ2wzB4/Zy1efI9+Na1RFNRQvc
eGdMfTgJe02/5aQxeR2Hmukr3i4NJ9vMksQcmWt1LzyEcks6RUOaJap7lj5/0hJAYx03509RKj1B
9QDaxN/6t3iv9HByCsJTrG7omdxIfEvYXhqXCytHpfVsD83J78O+zEc3RAKayqMwUAzgcuqWHnWe
/9zZMoWs79X4Oy8BTiBKxfjSxW+0L4ZYJScJyxnpjDrwnrcDr5rYtq4zigJUzU2+rNkEPrhAHR+r
RDdR2ssjYM64FlWVjwu3z2++7nPvDwxoad2uaCT1P+nWmX2Pc+t0I8jpufojNF3L+fSrQ+EDuo+d
IhwbF90MLidBbKNLl1yP0b5/I2Funq01Btnb0xBLYKzLIuddJ3rALQpCHuquj3YHDISxu53xsQ5b
BvdePhmZZAfRPu7ZXR9ojqGFoLA3UBqbd3r5f6UXuyy6GDPkZBIzO5eS50U9phh5ebBdtNPD/2Ml
BVtlyLnY/omvuKggWBGtOYmgNfmbsMBol41A5GnvyF/BxnggMTb9Br84Cwce+MjAOgEvLeLtPfuk
EJ4rhgYvRt+YrUYqEoP47RMMakbGUntxJWTO64sJz18F1kfNhNRRZt9nmxHu3V/bFcGD0ZxE4e+V
09ho+wC9LhU+kOmrp2KHnfvWqJ5DX4MPhkNfk8nJe8+6ehm1YFQnkf8jagSba0TFeb8oy68ilPPX
Lt/1LmZk3HNmjkmTMkJjWbbp/ON/WCcHvscanq+sHQAqcB2qk91gDHowmEhWLO3oDQRd6T17/KSh
HLwToCo4qbt9SkYOv9a9hzfhMuORKo1EGD75BwCYvwek0zGafl2MiOuYR7XxGSwYsTkOqzuog9mg
K9P7VX3ZiTMKL/I3EV4Dp+VSg3n3ojCLR84GkCkLySEForO8uPrKpl+HpAlBHagEkfA4KdeEkuXi
iP6ON1aAFx2wS4f0cx2JqUOkEHheeUOFJah5cI/LXctlHgDdwmOwTAkkNnJBg6tS492d58rXgd0A
b6yXwdlCHqORBrkcBAFFURNimSdlew5brUfSqp9/cZ4cPb0tv+N7cY8uGbV/ParUY5YY/l1sVaXv
x2qCydzDhVbT5keGozmKbB1J9LXENIkFeWaoZD3d8MPEsb6O4ilzIUhz+03vs3i9fuq0ueZ3AC1s
d6R2N1w8jtCjcUagqqLiOGvwIcuQNTwOfHT9sgkB48QLy4NAsz8n/Li0svXMAufi3s7Im98enb66
9tyDcy5fv7EkK8F0eXlsciRvKvAJXzZFAtAIO2tRuTqe4Wt+pSOEig/4G6XCadCaxFvpdxWNiOtB
t08cTJBhLOMGYRdK1S99ZB3jnz6t4LKKZqBzkIuG0n8cAQdKb6fVAjpAbfKI/ZcNn6SkavOb5G13
cp4KOemslwqHklvsse+ZhCbybLqlHw/oTKmmW/XbMFTI35vSZsHxXviEB263/Gkqtw0M93am18lN
N3zDYHjlHZNJapjkXf/gK+FNx1XJaGIwGi/9aonB7yjJrOKDVjL1S+v6ckHblvStX1h1Y/Ns4ggm
vS/rKEfKGxuho7l7VuPe1oCp8kjfOjm7VIj/mT68xpjDSdG01xK0JTWbNmh6a/RpW/8VLAt19YYX
4/c1v8WvmgZCgV8m/IIeaRfLvGYtO/iClkOuK8w2gbSz7kvNHkhxA7GhL4HLrxzsGjuM69kZlhyp
sybj1YUHnj16e8EOibr9rte3suEEyrzQsw5NDnvLLQ42nH+HlM1+0uB6OvSNnybS9I+VcorGyGy1
dCILoCW/DmAmYa+L15QlU5zmqpCRa8WmPcux4QnXSMV0othi3mKNO7aHQURUSFA49lg7ux8SETPq
H4sSBo0kGNF6nFeuritBJuMXIdknsYQcQki2/jLqoSr6wu+X6K5BfTNCJkzaPsO+YiMqvSWjUtCa
rp0NLTygq6E6zRcCvGyhLzewb/Uh16KGEwdtYQkbhQJofcAxbc65H1U3DFq6D+XjgT0lg5nVCwk0
966i3v+DFxyk+YbXp8nE6RQkw8wwheNytdUGQ3YXerqk1CkGcLidNyuSdTW/b8BlhAIXX3f2HkFo
k77oJM9JCgebumwP0nPExeJ+nhirYT9gsZWP6Ds02kUUAc+7dTyEzV7CzdKKVlfP2ysyIAMD02xd
aDt+j2EK6ohb/oG3q/KWWX1OFr1mQukbETWkS0+tZnbuzFhToHLA0V8gasn0tjMb/HFGH53P5JTU
+8utrfDG+J5ydOYpuO+qvH6Rr/AwlhFeFox0j3TVv/fvmojD5sCU3oFwUh6N3SUz54niDNSKBB4r
jxGmsEqQBvXMoaYZN38NsQYY/Er1uauvEXqtPdTcKANHvyEY1Qg3r0geNcs/H/ILyTskJibQ9aVg
tSKeAHUWFPZBh4/DKSVB36I2UvLULb0qQYOUx7b0XToLPrddPMTY9NAnBakaRHfSGUM34hyeux3b
jg6smiPfS3rFV1InnIBrOioLCcz+mVFGEHwFEBbCPtLeY+SWmiFQbV3yVQFnzRhmXTgP+6IqM1Gr
dguMWGtBx2xCHtxAaFVKXKoe4jtpUa163x3BZH2uy/K44B6vxqEIqRumooUfZ7ItPnLaQxOdQD+Z
iujOAO5mzqd1Npbt6e2xm1Bs0M24ypICg6MKWFNPdIjP9jWg8LN+kyLiUSFz+kAls7tyPuet8nPo
D0YqjssCgYq1WARC3VqJk+566hGznZcgBZqpqy/sF8bn0aaEYJjVuUmJ1D5hi1Nhmdi12TfQFf1K
QPRVEyjcILHr+fdGnK8CphUs282O9/ctILs6mgud6ddosOVwFpoGS0n+Y+zPW/92xpMDgIwfd7p7
Y9qljbX/hY5PhFiEh0jKfAEevbE4UHJBBC5tWCQQVIMYOCy9G0Qyxp99azRhaODX7w0yaLXyQPhU
VBXDMVKlYaKX8sUrmz2Gslp48M8FsZm39QuI669s4RVVUHdg7mSDCtTkAjWAv0xW+VmIHBlR1LCv
vKjFdwTHkYxFh/KREqR+sn+hq62fxK4vesRzYNbrU0q/NyfPfQUvylSLgzlPcFaXCrM36YOvQv8x
HIcmBo5O+nwwFqOxdSMVWuIBg+VOE6sZS+P/z13SydjsrX4TiwXleZTIL4niw/+QxwlTWgN4Ydn4
2S3RLI8caKmrEZ/b9PRiR6MGcBcFesWHSN/i2BwZRSZCs6WUovCKW3zy/vWjPj2CjFMTc55pUuKe
p0bROHVv22ufZfRatG1KT9ZAzrPH1at9PLK6hKxllFC/UTde1d1Z0jNMAUuK7SO3Cee2I8uAEFXD
6/H7sP5vxINveGh+ptnNsfJS05mej+E9JujcWCMqOmIvvN8cbwxe7/bwwBo4DPke18m2b0Sz0TQO
5dWd52cUeJYOMwBeTF+0BBrQeLgogQWjcuvAYq2jejWBDEn7szSB4GAm2K+ct4nt5XzO3xleM+Bz
yL0l1IAlwBNz7jDDR6MO2K8I3gxaqS/IEAgatasrCWX5BoPutoylhHKtp1oibVTmaleAkmFxU0kg
KkFJHD4HDlAx/CvHot8uaFKIpVhLpwsxZCod5RVnnxKbr3GJd5mbTqY5/nc6c/5wLCAKYRXxg1lx
sqAZPDt+2bcBSGbBhifbUlh6i5K0dHKUMRycupiJC231bTkuiwagpKFKNCyU7GeOdKkOjVaaSJwx
Bk7NlXrOs/RqjhaCNsal9S+7fHeNx6m9tQ2OxeL/0DntPhfn4mhEstkfI4XVbqmeA2cpnDJHcVuC
qHECS4FxjEMUJTF485vu53uhCk+snC2giAF4Fg1vJpzomdBzTghIsuMjl4WVrIvuwXEy0NfgsbJp
foOXiMM18KcvLrDYYAUwsdlERJP3AYd8xW29VWhIyt8EdrFq4R64futDb8+yhe1qA/km7TonA7jF
T4e4YNPE3UiqupzVr2XFz/p1X1JpF7pj8KRCFC40vtLbtXLAl5T3pYolXdX6vD9dmBTB00KXcFWX
XdrA+Exy3RpmEv9plEqoyktG9DA6fvBGL5uhSETbXQMv0z+lDlg/mVTRfNccq8+BDNkedkGP5Qrt
yu4aEFX9MGvGMl/L1LH3/WLp8F6kwnO2zkkGcOCuJfFIaULGKIPlw979kGNku0kx+8vdPd0X/Gm/
5qOl7vtuGYBlans/jHkjWeCr9aPnHVAhcHzHZfZZRilnLMUG+Fp62oPNb+o0k15TwXqa8pJwx5CT
cGjUbc6z7JNBul9sdTlZkua0xAWuz/JY4QPehdt/SWUeSnVsX/crSfu3ZPiMf5gGpPuYldpwxQCB
fV3AUlawHLXL7HQwnf/Z1JBEOl1fYuRTEJchLmvFO7aZhXtLbJM1gr63Vu7cmFN4bw26EgdXL+le
pIZuLse3PhKCdvkojAW/DiJNiHfJKPsIjEs2RQVSZChu9AojHNwKT2y5/fQwifU0iAGRN903MB82
ltedAGIxH1ELGrcQ1Dz5t+iHHgNFipotMYJONNMJFKkJ9GX4Dz56SmWreWA1HrMb5CLxLV2rmQsb
dctaOLee/d5twtWWki8UxoKyokzXBR4bt0OxI05BHjAK3jcZQz9YKV7KTlPQOqNcvCHvHaXcOv1g
B4Ks++OWSYYiLLhedqD1tHBL6HFg7eaAemQz3YhLyCa1zv8/u4zMvI0Iz6uIp6e8fhKtqRWrFNYd
PhZsDZxgR/rRMUAuQCWTosi16QuTyr6lJdGUekB4X0HkmThfcX3qk+pftygHfAR4MKYZemj+w14D
Y9fIiGP8X7nNLwzZjtuw9HsSuFvG6AO0QSVu3FAokQgbvfu/01GiCkrdYFs1LY2mawn6J7dtYmbr
+n/Y2wTG6AF7BAzrUAFj5PAUYHl9dnO0Azb2rwwjjREg1aXQclMfI0OnRJQxri0tlJ8bRdY9+o2+
s/+MX94vOCFSOxkrt0POWkxc+3KP37a29pPSqmfPTj/Kn6hNPwOogdw/BeNjsbiouvBnv4dsNOLa
SwYd0lJVon3qdYCww70lBAxVEYfKzs8v+FjnRe+gQZnoNAApUJSyqdp3STT+hR0rQsdhyRH/KRcE
ofdaqs7VIxSoKqhlxOSiIZDLL4A4DGOxiaw5vhy50JRtgnaitOetiRsV60VAXTEcf38o3ZY7rmTI
++vlbI6ODYaUv8fPMOYEYQW/A1ao8atfkWOgFMZJa8bD6/dJqGp2SfjSx175bIwEwjaqt2vTsGnL
9WvMS5muASg2PyUjj8TCqdAHG66Du8HrjztwKjp/b8bKU7ckMj3hfXZQOWUBZ63JmC95wmF+e1qn
zTqo3ehrNGLH/Nl8pVn3uYUSpfyvnZFAU6DKVJXO8V1UeOZx1XUbMjNY8HzDgTU9yu+/06WG0edX
GONOP0G7B3yA6LssEP1P2AKrtIXwkxMGuKi+FidHsSwcFQOaGS1/YPLblWbGbr1ilXq5KYfgAMDJ
NPZke/o+z/GaEpl3dKCxCUuJ8O2f8lXiKIRYOg7P4czl6sp2B2AmRBMOMIPNFMHle7S2YeuYTDnb
RWqQgNt550nG8WOa9xpidvjq0grHeUSnwFYROBin+gEOePcDkHd/LCce7KFSmcVTGXBq5W5TikmT
oN8qsJ+QUWnsflxIvrRtm+SToRRWqQACDzPj7soNrB+HMl/0c8jn3BE6reYElgIINiRO47Cf00EV
7DI3Fpg6kRzMXBh6ZHhpOZWOGQegmcIffTdwL1WMYhI/+xjVfeZaBxkb1lA7fUYT/2MTz+XXXwNR
B08nbFLnDzetxX5maMB+URV2V4hLqFqwS6VHrRgRNvLVXt6GzQEadrpd0FICYpWps4n+NwFFbHiW
P2k4Q8cp9/Q7ChrdFr/aAniOCJ6VvzTAjfjwBzW2wvZSFDEe8E2PN+Px+R4Q00cCkIpFAemaZZ1Y
R9y/ANetqd2wQWCn25zjkG8p8iTUDAqg9OIqJTE3ixJJptD17M/zkeQoKe1HdH2r4ZNpZ5HjEh9+
uyRrNt4s+DE4F0XpQE+phxPyRLQj+OW+WCCHj7oYSrYHhBdbY8Ju6TpFZVj27xv7R6Kmaa1Dcxag
krWjnLpIssx9UFfT+bgZsoOjRQWxetISbKL0EDoaKKfM+mrZ3qM1Zx9EKaT2Vdp7mDvPsLSpLIGC
6bJDIGcc2ufyuo8XyaxJwwaEcAkw2tYd6VMuoN2wT2PV2rQ3IvjiuoMFwR3Ktn9s0bVETc0GIeHY
ahMGcj0utRXSsy+Aux4+mKgNrwGKV/PsxmnY7RbQ6ufp2ezyr9qh2GtZ+7bM0MZn+s8EIL3inihj
6HiIy9xAA5+aVzpskDMEFMy4+1rL7rfC5juPTumrUur7pgKCOsH9gFKvYoCk9GfeVo70mpiz5bKS
ol6g5RXLC6YV7nvsZUzMQMApaFWqWLjmT/xnlfY+0TX0VEerDNwYt0oYCXsvKnqxXr+1LngN71m1
GrYsUkZlzKpUsyHW0tLMo9d3JFv27pSlzfekw6EgbFtMzxmutpdOPFO5757ViwbM6pEthI9nEmrc
ZShb7AySvIlSZkUEW7ffroTtaXp/Ar+KUNR+3EUuKSm1WnbQDGRb/XzUM/c1k0UnShn6cVn91/HA
XcxUSTZUoStyVJpzJvDLi2rLYAd3+5+lp9RoEg5nj9MtcHFG3EWpY6enWKTI/RoqYDpF/488yL6d
dk4oLOoEQFIlJI6CiYiIqKbOcIkjgTmW3S6sSX9uzd9z7PN8ta1B22pqzKLPxth1OAEtQCxy7rc3
2j6ZkfB8+KygH8j1QxkgvAHgRWPt/Cdvd+u8MvYIFQl50tkbp56padlXvKcU73iA8rM+M8aELT9A
1F02wrwNKSfa7LfmyifNLDdvMLFm2/oHbvsfWZJarx9bs3RCXdn4F22+9MzapHjPbx65l9kDGJXO
HOVQT6C5yYsGKpmpJ4P1rLCTQsfz3Z4AO5tCzB8Dpzh8D/NRO5jg2jii5nDHndziWrjRMV6HB834
nvX0ZNWQi4eXazRFgE7U49JSemrUMfERnUbCkT+qbAduqzwRicPMZJZAmR1WLKrU60p/7nnsiW9d
bqD5xwWV1qB2p7/ZJ7JPIBVQFU2GZ8qOJhsQJiXiw1mHECnWLE9TRAGCFsiVbhTgkRc178QmSGUt
/6pWu2yoOLecyf/cU3C2qSDCo7pouC4kiaompwvRFS6OihUpGyP6I5y8Sx/yK9MSomnx2nfHsoSw
7zwchFaZwNc58ocx9dwWG6PHHtN8DRNmBYZ+nmX+30jWeI7WKrZTqZwan3wQ9wbfCiSFY0rxxZU3
kZjASpisMG1tRSMQwJjiq+pIQPeba1of1sYz9E5nu1ujm3EXRvrZ+hqvDe9sI7ViiWQlLzjE8P1a
UzIR0gsEh4SHycxvT+oYCWU9LTeF/pEcw5wUnx9myljoM/yye1GeuS8pj/c0q3AN4Nx7/9Dkoken
yvfAtV0RxWQ6oIWWNGLJfR+dzzBLiqHIpNEG2BbgH/z1C9WRV4F4bNflDhcd4FJyyHdeltJ5ZScb
56kFPtfi9ZipYf28yIbll3KjmL5tZAhsWcEZt/HbYFJzOHqO9tSY19fyL91xfy7lWKq5WaJ3s98y
eQQZ1HSxqprK5+8uO3+G3KaVrVp5Cq7Mo6+etzzQoVSiH+R/41L4Rdv/wl7dR7fQeup1e2n4Byzq
kSObNphrICEsvyyKtKlhn46Yeri1QktzdzWC2gw8HW6cN328PsdbUd6BuatID64Itq/V8FSBWxjj
bJMHd6IUNmeIAIAvta5IbCO3Vm239uuOLWE5qyL97NdqwVULe/dPKEDVXXiXk9pENdcOeogGEj54
7Wihq1haGwnJI5UgyqCep4dwVeECaMxLWax/OS3CSpsHOhKNJi9A3kJsz9HeT31UYqO5TSSUs22O
0O1I/f4bajOOrAZbaUjSyup4ylTzdAVtkrnxf7eFXiHOTc5szOQqvN841keD9iiLkW1qj/cpJGw+
woTkoexT435n111W9nwVJBGTXmDxFnRXdn/OlbyLTNAqh+ttaZM8lpi+GsqeAwqvPM0lUXZje4Io
xX7/GMlTnBGFbla63DRfJp+UAv9crG8zT2SG01Q2c2Vz536EeCPTaJl6aCeRN/pQluddNirOJ5GW
GbDeSMJXVQb2e7IXhrtNMoGiUVX6J0RvLZCiSY9ntcU37giDCeI4FdVS8kJ42N5OrzStcsjY/EWG
WLQ3K4XHCUUHM3NglDdv8hIEr2pWXw7725jY05Px6slWLVmon0ygILgp2N8x/3dMN3i4HsVoL6Qx
/y5wdMZbpOx6xJzOrfNYDF+FYjrQIFZPVjdLekmUTjc1wJKnnSjFXnSXanuOhgVxSX+8278cjZvy
MsCl0IvjKZC11u52eycVWfibZGL7+L43HxPXnODHiHofV3TafMxzoKoKx4zhsss3wfJbVtqsyEfQ
soRrCD3+OTvIPFXPTY3iIvTOaGYAJXx8O/B6AKR9G+wwEs10bJSIHkivdjt/wrknYnuXL+I+cFgO
TNwqrMsW+fdnHj59fsP+7u18G3cYLgQrbkwGUkz4bQdr7T6ah4pmKp6UzMcPGr+Omx5DUaUAapY6
X5VXBIcxSopAMRKbo0B1AOZQaZ0iAswYBsJnxtn/OI8/s6QCFmAajyjZdaWNnzhar0NX7NjljwqD
QSIt/m2A9VytwFNY9SjSVe7t0zKBiEXvjjYGmFbG884pIz3d1DctZfmcNI/9M2Bq2IGHI26MLWXX
BSerL9d4+tQGNUY/nmT41aME0/qXpgUXDlN1ZCLP7FGdEsWjWZsXIp4tLJeGmnKqbm5oKMfP+kTf
iUquuSOhU4ShH/xmtVLQkhbF6abV/giMRRjYpRzYdyqHSxRQ7LsuXdPNRZib1yev/1PQlAkEKZE4
v/+2o7Romh2be9Ce1jhVhlG5lEx5w1zcDWiiJcHlUxNmL76LEUIzSNgHR6jfbztXF6fDEPCTCJ42
QnZQT3iOqdxSfnlpg3ypaJ1xJc0d6vtJW4+olXtkuenpz1JwqNTHCeogol/z06K/CU3uhkHnvpm9
swAou1qTqPoH+8QU65ti3A1GLUf4cdQo32lhlGSrwINHLls92PdiBml4o/OnOBymObK9kD459sDp
EbV92Kr6pm9e6PD7Vhsyj47dhB3Ut0yoYqN365JMyYygD+mV3WSPo4/JK7bZ7j4Q4kk8mcMS2y7F
ZurOcO+3mKiFnB0xF8E+jbj4XEhvC1fkaPsepDn5FfuCiV/lbhW31OC2xLCWGlLDu/M7omMr7DPr
vM4bm6SIH8VGKtPDMTNv5ZSrtu3CDRT7jI1MXDuSGnIjMPhOi963cHl8mNGsJ9MDZfg2M7oUBh5B
IgM0wgT2vohJUeRGhdaigPyshipyYWI0m3pug9LrwkcB2GEiDT/psSCDEiaP7xBQayaNo7J9R+bw
eX0gjShUZaG03tUsCpQkGWg6Z11uzFEemxiXeiZMfa1mN08658kKhx6cejJ+istZrOf9br1sl58z
X2ihFjkQPz6po9l1krP1W0HX6Ti5ICmWvyOwsAMnEt9X5aFPfF97GEtMPdY0nL4Pz8+nzgT0V57K
DRIoSeVGildMB9ei0umhh5WaDHFBu1KLuRSDRK5bU9E9m9iFdxGIDJY0KpkPq9TEjP6CrLSVZjXe
4+kFe/kHdcyRzqm0ZI9sAXEzkmN8JpS++9j8Z0Bnqo3s9HaHHuzutEnP3Wjo7A1/A9nqUk42/AvO
JBGkclTflxmTMt6idMpZPqVdt7o/hRN/5f/dgL3HtjIzzNf/HcLPmJnkWig1T7VLbFUv4WUyT4Vg
6WHmrAXrP1etcqEHUBPaAJbLjFx0xov7mYSYvGWd0PW4P3oLT5RZO72V/kDiDK5Tm2wKVPOMlw2z
S1rzcmMlS4vtVg/kEszZJAjAwxIllLW2gQBfV9l7xi4KLyxxXXhorFQfNLJFVbisP9rsjSiJdbR4
vguLKUyG8KVEzdHOgyoV2IyFlNtqzdB+H7qZQrmv+LU7R5oCjjrUrVvy8ZOXBzt2N5v4NP/GBCmF
DndB27YZroMdLq4OGmtywwbvcLnwixigHuQ09L9LzzKKsZY8nUprjQSLR4vlHCcbXN3nJg5MO4mh
pagwfzHuthGHAY2IapM0xOX/oRxNLOu6/GxtmewFLkZfsvLFQ8Pjw/9HlR7BtUfsOqLqKxsCk4+A
3ocWH+yhDdl45dMvDgbXUy81iFnFAbiWHZEEajuQAqKcMOb303llE9VqAkNSdTJXkgAz2PyXbCxL
KHzHqLGbo0rdfWWxufNDPKQJ7GcuBdFWY7GDL1RBsUvQoFHbM4H27ir8sEJ9fLBmQ91xQe0KAK87
gFOljx9oh1oFmUXSNc6CouICHg/oyRGI1u43pgsaXVX8vBHoY5RZfZcycYdBeVPcwBRJVGjZddIa
crqJ+UP2vHQNY9cuTNjBlhKn57D8P6VmRbZN+eJ1jto8dZ9pP7GaeIy6g/Y+IRY3khZ+DgwzyXT7
aw0PRUhQ6R6GXD/gBPA1HITtqWgwjcfqlk5pPN7SOPx987mK/jhAnCHuM6BCpQ4l7hoOq7dwc0i/
TauqDbmDG7c6mUXgeBWznixkJ+HZHcQSdmb6aKXPtnSkBCZuBGiudF5PXZFolu+8B1ZvkjrXzV3/
n8Ah7sFZHjfKWI0GzejPgazTsIBHhWQIiveLQG/ESYKOHXymcYiBHOgbE4qklvXKvkw13tfbkZHD
cWSasJGJcLzxfETJvVOhRvYy/ZINw1mSeKcmrNLg+qf60Qhu2kYy2Wv8O+dLzwDf4BSQSdQwsb4O
bTIfh/DdHvGrf7MQGUq2jQWdlHK7fVUKpGtGo3UheuCA/RavBB7qkuN9pckpycrdBmHXDUHeO4Mf
Y88L/hL7Vv0PG01lh8HMgQBa/Ci1tA3FnbiIGJXnPyKi7JDJTOiHMzi9SPA9445f7mO1v94US7qS
3dYhSCz836dYMqEr5bzG3jeEzOnfKtKjYImaCAqYlrmCGN3mp6eU+oEPzC3iF9p8ubPqOjM28rs4
jFC+shQG7uNQNLZF5hisG5XgLpDGmPx0k7J8IovcKMLbMbHBPsjWWtIQG4uSmdagkubE6BWuKAjV
XGRoDR5NJcZxfZ5pRLGpQYkuhCXnP9VGeVjS13/JL5lCs77ZKskRkltIqoAQbcoZ423G7pJ1FnBu
lbGwEGnHyLZ1gUStsd9JZUqUejmla1zBufDbUbpJqDTKp+mKTuD5Fz84La0hXn9C9Iv37WkbnMRe
KS42hpX8b6rdONQFe5a2KuZl8Kk6NsDUAtmjevXS9neuZ5ujPXAZCSL4NTHtIGxS5lAj5kPMxdxy
KO8d3II763KThg0+ljmgi7FPdK7PH6T21gEyzDrD4bvVHe4cAFie2xyVHGE6q0TrEMP5LUqxsLSY
uoti9vEHC+JV1vr8+l4MdmfhuXVEVF+ZxmxO3mD4aw73ErECCf7ZDKuSO/1V3BiApOayn1GZJm0f
YWoJUalwFhrRF3M9/5SmkbEh3x/IlhS7IG0F6+joOhJnpvR4/VRxJ487YusH335zTJhoU791R+MO
fuRf+vt23+m4X3GZBMzB2DeBURt6gQ9anC8XqfTg73BM1Uk/P8lVQefkAQdbtHZTsPuZHEwS6wIB
mFcmrR6iY6n0jYzdBMV0biHRYAsCOMs27LI6qn84dajVH2iwfbzscZXR1lys8Zcvr3uOlLiIURQY
5j5MlIk7oXoxixt7pjSoIP/BZTLhUXOA7s/hhjgD1dtLX93xIqsMdHEx6NVAnEiaRRbGTWJgiAoV
ll16eRvpQYYjTIbOZhBwKGp9+5QBEQVLv8LF/HE9J0W8ZbUiIIPFLEdtH44/aWD1tr0uqaLlnD5O
8an3lNvDLrRgsVu6jua9C/djgPcTm1Ww/gWJJ7pQFVnMtTAKW7os7zfbiegAy0UZSscHiDCb9QOL
Pm5BhTA8vGyODmJTIEhaxXglSqZ+yyLnQt5aIrn3HqYdCHjDboAavQLCGxSCxk2QfjFhbY/JUGzp
q8YhBj8STOw3bFVzoFIWXP5g421WPYHpgBRbr/2ig4Nm5mFMjsI6pXYTeYrVVrpIhaP6G6yvlWTs
KgwIBo+KkOEhMhKjo4cZZUpPDM2xN5co18wrd8JBSnX5Em1eXcJ0i5EMb46hrLQ+HqUtPyIfBn3l
2ZyNmh+3hi/hRizg8WEjXEQCaZiBu1M6Big6rMXGXlJaYgCzqMIUUr5MVxvs1s1q/vckU1qSkf0d
6coEsSE8CNKW0FeE2nCKkDLD9h9EMwRYmrG6Uio2OQa1hOTogZgHK48/+SPRg5BQh2svaOf4JriO
VwZ1xUEZz4pzSY1hQFOVXUYEriWtR7984K9UOF0pgU596YNRO0pSh/AhdkZM6l5xIr50vfOz5CPx
MR+BB+a1ujoVADqDWddAZCia9UVhHt/kOTo7G864+UPAHjhUZH8VDW9R7axCSbogVwovqxoR5b/E
5+U4LaAX7J8cyjzB93rQC9N9JpzocLiJExHUq6DG5BHJ96awqGJ8Jfnc3FntHb25YCvTACRLqbxd
gVUZSDplmtdDlfCdrOYP54aM+ggq0NcJqXHz1v6VgmtRPexMEgwNb1BNJnu5Qsv1Y+B6Sitley/a
n77zbGzV1HZQYWdHdmTbaD4RYXu+oRt0eafs9HD/Am8JrrDbsoE+7ECXHxvMAQ3EXMGEB/aLY+aG
9yRNEYAaUfa8xyMSsatSzhwvOj9Qr57C2cF9Qh8uEvnk3kHCLJPXYTs0uiWGyQG+7s+6F7egt89f
VnuvtNBfY3PNb4cPaC/RY3FCffxJ50WYyuUsRFImT9w8g6sPUfytXoKQ9GTTIkc76ttrwxisKgut
aLs/pzvj+h+QMU9JMLmE7BHNzwFb6CFC77vOdXT7gp+xukCLV0GhEcyV+NWscLFZU/B2bn3SUnCG
z7PWIdqy3io05h2MmgITgnkNQLwln7nmBhVBAzaSjr2UEi2XO2ZNgRznHHrzraBgTBDcBq+PSMsi
vXPtZuQhTdBz7S0YvAVhB0OliId0HXaIr7F1d1dYAnSCwowoWdWAaxwpiwPGs8FRQcEpSvYSOelz
Olh2kIfvhykMDR2NISVP1kc3rIZ3HL4H76EPXTdDQaF4beSJBLx71NSHN8BVmxpgS2uh9abiMBoG
Bz1TJ2mBM6sv6y0wpagZCLQkjG51M9FYBNwb2iQq3okTF2uS/r4URunI+vgSmeWIlSUUsnyRwdur
UnS17mfonm+DeyEdiFPPoL7LtvYfZ+WMTawwsKWRd1/QhH2TRG8IzuQ9Iz9ly3mDO7VkdQM/dDp5
y9GDlpxmwstr8WLf02/BioDCzsDhi/RJnVCSekH/Pr2qUeQShenkyO5/8tF/2vuQ3vrm+AIc5hCS
U9lfMc6pOPdxT8mMbbyxghrfS8olTIrup1KVuNvKVihzokyfYqIwjtn7x99f5OEYjgcN8A9ZeW+K
c1oHXAsXetmBaix/FiwoiBDpyCxDh/ZQ9hk8mgaNH0m/4Bi9/EDKHXeiuIqIa5mQLrhebit6GUIU
aBBF3qPN39QJyyG1obS9WAOF5swxLOIqIPhv8llOPabZDLD+aYFnIE/IhnNpxSFCVlt6iaPwOxpB
NHVYJIeoTWWm0mlXa3X6bawnEosj5luPOVKhU4f58gAPfFUaXPDBrabXdhFhvajYH0Il0bKpHNGN
0Abl4PHnrpAThnnq9gA8dJhdik3Y0qWxIiIZD/ba2+P2HNzDP5fQ1ys9Oz8fLu+rq913163fQ1bI
pLgcnSqLKfG3t6VAG2Ozc5izmJRdbjoQFa6vJZ9jUPfdVmP3eQ6hW+wDuzEL3+G9WJURRrpaWz6u
u0QK4iMYQ5YDnzf4Qdn8eUzXuKu4B2nEiEz3P1Ktg0qbDqur2MUsnfCmcgr5/IDvno7/3W1rLk6/
XC1/DGUh7cWOiXMvoZpUxaxfZ+EVycd/B5CLjy50t9TVphTUTSJ8RMjasbPSzeH8B4SrflW0L3/H
xoL6tF9CsA0abtz1mvAePaCoBYnh+pQslIq4xA+kLyXd9tjs1RhCuT05JX+2+/Mll5dH02UXxrhe
m5Dc+P0wo6XbXaKomSQff6Jkn9j92RSgXwkuW7Fs3SsweuMq0mGCZfY5/ShxFsu3TXyyWOdLOdnv
S2iNtMFF9ffBnOfvIx8b6mPKLkb/KPhu9e4AncYFTSXE+ZzFze2jYypDCLQH2LN+BwqmEQ7qSQ2e
TcljXBAyto2IS1cXxPHD13mPpJ2KULiZtWkN56kw3XksyGLmSN0VoeBbshqCZhVOMKmbGGvuHMx4
mIFRYCTCNoGQ+uIZBx1KvA+WxgmBf74QHIJNZRcT+e19k+YVT/zY9qainp/EnVHsduM1qnOC9bRd
IVw4qQPgFpxtHudKpPuBWhhQwCZweFvCEcOi5fmRi11sJAuVzD6FPl1hwt+3UE7hrXWgAi7ND1AT
7ebJvB7mkW8lRycG52UAWyX3hTFCEBsABZPN9MnQa5ZFyPKbX+se5EJNt5S/3rPEmwtObjJsApRd
NIyJleS+GWa5nOrXS2519tIcEtClX7mK4E47qMKBxcy8NWfwRJXEX7JCa1qhALdKfzDKKjgHG5Gv
EdHlpJd4qoUzvp3Hx7wGUAQSboWFso1rRMjSAERMALJCLebcQSKMsZfZzId6H9k/0Y/DESD4g4OI
ZW+RpLfgFQgjHB2KuOjEPOmmmPAF2NjVXSicjG8mMPgafwdqpBR56N5TqDciGMH9+2AXq9dtdnSh
JjZlrG5ovrrW43xgSVA+Tkww8DLQBsReLUYpzkUJ+HLNzbgC9WWuHOpZgNA4v6c5FJtZ7y5I6P2s
bsMB4zq/6ZvvsJ5/KfHz6Uk9uXr59eByObORrRsC1TpyvBtAIT2ZI99xc1thz/bcUUhKf0FNgh4d
1Kj0ykmbfoE8XdO7Qtcl1WOLNzuoIbNbbp97Td2j+4EiEgU6Fhw/xRECjTcP4Q9qk8f82VeFkS7P
fITsH3Vy/sERVhRI7+G7tHhipHYA6olULm3esZKr6jNPVZIBDX0xvOK0mibNbtbaA8laJVHzuR7s
5G1dPq7IP1KI1eOlKQHflDsq+AQOMKtY/WVBCobNu4w+Yer1OLEgvxMbxtYVaMaX1n3n0h4Z0ukp
mD6t7gjmdMnDXiz8fAzvdEI8m8u6FMwj2ksoZaCNKLnUpcnr53+yVXvo71qWWyteyP4afjLyGPng
R62dYTdM8M9dGHViODt8AB07lm/qdGhQEyKLCdbUTNHRgTL8pyCf4UsTuY6630lQfimeJnWatE1w
MZjG6ndo9uO/Ow2AgWfhccUWMASwWaEU3Vo1z0URDJ6t7+oU8fh75Y55x8H0Mvmm4qnXlaxQbxJT
WlVm0fMEGfwM4By0LKIPML6Cnnh8yLR6oU9u6h5J/wZXjN5dV6fkMg8rRM4+Ytx1DzHsCZ06wZU4
6CoFmQQ+gy1aXytTXY6WeI+wtA21Smub9CIpjt+QwkgQHshpRzGehlJSo2lUsIiKKwTZ2NnT4xBw
KzZ8etc0qlmxuduDFTVXX198PtPC5Vcw/eHwzHzhGN7Q3OAgcWI+uaNW7wNflueBIFmkC2Zk5b8y
I2ovhcBdWIcQxX1sD0AyA5v1mPytjKq+xsvk+7Y9VXrYOTr6X7GgtnEaVbuXe7Lr6BtG17yHFmyL
Syi9Jhl+8kVFD229I6EInsgXxJL2IMXoEilwWM6kTAVyvQyGAODd7C1o/p8D1BWsn88xODhP/Omx
vkAgZBGpQEuKBsRB6urJnApyKI59Y1t1+QUliOwzqhPo+8gb5zO2Fv2+IZ5h0tj/KVgLiJ30tcLW
DCqT1AIK76fpLe+XYj9opOYJHSGNaOMq9+oXudRNj6jO00KoFAt9t5qLMbnRsn5mlHm6yHglbI5e
GrjnWGH/F7KIn1OpNyydgyDrW6OaDpBNeaurCXIp/r7Jd4/pC/Qlr5ug5qKbMM/0skl4D2PM2yxv
MaIPfuTpaWpZNGf/wuKkyL9VnXminrGLfUbSstGhB1nytt1EpnSC0HwEGja3m0KDkX3N5IcypIiW
GaTK/JGqu8+uOOkdJwPQymzvY9i3tP7yUaiZhBg+HJzVg1POUtFp6vs9VxrAKy3ZHV3gV6JwDge8
TX4w9lwMCbSqFLM5F0anNB9D4IVHKBo/RAkMzUVHis/ug/1D+0Gz6X4u9SXcZKZCzNN+7HoaYhrE
lvn765A15JPtPGje8n2KyAKdIsJB/iBaCQNyrs7bTZNw3N1eYe7pBqx3RY/ckCamU50tnuvLIg0Q
9Vme54asy6J2nqNrY7zxjm9lH2dFbkSt06Ywl/TNJn5ACFSyzOtadaExFIRogpWCRzXOgEeCLzdM
G5ZfjgA9Aj7LzaISpOlPcvsI6DIBz9u6Ge4QJbyuslRpHX8QmbBJH4fvo61+HiXTmKMaJMUU3e0w
G86rxTKI4yiIjhoImQ6tf/3eDefLe0BTE7UYPFM5KLk6OVYB3nGIgSM59W6ZbVaPWM1S3OOe053i
1EmJQZrHV9lMMLdPnxjC/sOQRYos+gKk6YvzFQXkUqIwloT/5iuP+NnXZnpcwEVjpxoq/At04Ea+
qIwLpNnsSIsWjb4ENU0vuvrwNbrmXA2BylDsTw96h4+1RyImAYB0d+rJXYPrpRBTmLROWKM9qCwg
0DXphrUEqPS75VTtIhRhrk3lQZv2/MAIVkFFg+W8RuAvJ0i1rEBf0E0DbWGfMjVswaPap7gjEOjd
wHntUHVlnkGiiNUbout7sCmyTTwd97iUWgyrdeAgxMk56KQwcJSf337HxJQkcs3MKB80+UKt/6Iz
n5fMLll/fGeH5Vo1rp+mFV4CsvzA9YZAdkfPSGY+aIj+K4y5M2qO/9NN0zH/2yJZ6XiLzPrPKREH
Xp6OPOhrBJR/+Ih4lksxCW8dJn+pcbtrv+A7g/Gvg1JD2dpPDJec0MDmJDn513g8RQVOX8W3IQfI
gc68n6a4rVofIsBWJkU/FDk/KUjok/YlMupzhQtmu2hfqIC2hAr0gizqa5h0xYjKNu2xtZdIMQ5z
pKpMZzLch8AftoQZ0ACExoxDXQFj2qrII/Akb3ybzmJZH4libmpkIukha+i3w+YQo1Z3O6ro4vK7
9gVigeqIKf/pvhxkNvccKN3xHL32lOkTL3r7bq3dC4InqOSQ3YcGu+OatLoOsfuv19rr003s0l7E
LwovwLMoNNvZmG8POERKMNFqMKq5kMYvkt8W+kSyn3iiL5rgNInFddGWfS1CXuLcWf5buGeK9PNx
LlcFGj9k6tdNB4L1km3bbU2kqKElz6KU4GhMJGbhGQg0Tm+YgaWoObHvIIL0TIZ6qwM+XxT/bhD6
1znXg1+azprm/veieYwWM4ebJZBsLXcUzfmsyL+UT/zNr2v1r0Jr0C8toRuMajvg6rOVAstjLdZ8
gV/qtHYFWwZJl4DEo1Mkra5usx7CCuLjDB+yUbaTZ0jc14Qq2/6ibQpLH87o94OKEQB+YQr4Of3d
/MpZS6nubF5xcaYRLJ6ufY1trPh+cojc7akr2BUzNAMd6ijb80KvrowC5VZY3LZamxWZEtF4RJKr
pPOndGAMwzgWOSfAPGdWGX+xaK190fPlmhzaBCOx6KQNc+jpNFpyt5pwopVawNR96eCfmQTl/pjc
XzDtnKMM+BNDvATaMJN9SwUg9OjJlVg9yADF39q2rs2aiJDjpoJdX2Kb1KYQInuHjtS0npCzjjxK
wZiYOnEbp8Cgx45uz0ycXR+i6oyLh3O60G/sR/wdSPShgDOoAyOv0zD2HJ4jVLzb3C+tNpGgxHdQ
QYGedQ4PCLK3gP7bysaDr4FONQw7O9WhRqRrg/+DRXw4RAk+chRn9pxCYuxPX3bzNarDtetKmD86
U+vSvLxO1l1vRrBAl9xTj7DFVS/aqkA8JdkWaqyJ/3pui0+kbZnyBW/ySe4iK/jDhiRpWAz3mPo/
RFRLkRDJ+/AMFXpN+I2p91Ci5RelQHlLNsMINLXxZMb5rooi53TnQV4P6gm1TIE2nZSL3NmR98u/
AfsgeBX3kvZY+WLYeXjrWz5byMOLCG/0ImygYeNQqhozLDoRe6qrVP7l/8GO+qe2bnZpNZFplyzj
UIJbbmSViNQDxKinBYOiEiHELLFBl0m6TE03SBtoRC6wyC4DTESuu9/hItT8ad/xy+FBaccd0v2N
bIkAXVCIPgPx4w/thAYUh9qOZN/VRuwYsD3PmuOYlTlbzRPAy3XSbw4nwvDRhp1kQh1PSH19e1s/
7yi56PlMklVCZKqabdL2PBmB2Dw6vy4JMj4nSpIWBi1tHb2aJDFczVcxedIekUzsHiSPu+YwMZk+
FXE53BR29LH/yHubo2UAbjGhB6RzOWv3bzxmlKDUXfegGK2YMBU0pF0zCgZKlJ/e986ELP78cgmb
1wlHHsMVpSP3cEufEDGmNti/APzTZ7cpSbT291hdpz38GrW0qu4qVI5m375LzDwUTryh23VumBor
ihqEukjKD+puT7d34etwCeJ4+ml4KkqowDuYEvD5LTL5NlQssO/cjy9HD+EbOjn85AlFcEhsn3h+
4bZiQiePMhUiRrEEcIK/n1pGGALklEeb9uC2WXa04bDK85lAIEGcaoKSdqWxxOh/8VLS9Mb8ovSe
+31fidQo3dWECjK9Q03y6WlkAxA4tT+N2p787ebV6CBI60ww8nLqUyKP6sOxHrIHgsMvbyQmSKte
D25gdL2nR0v6tdp+5px79w5GBjkVTcP17h41n/XM+H75miNzIHAJDgzo7oIP2uAI8FR+g90pgB6a
3QqZf4yTG/YG3MiapExFpJsDPisS7va2D6Au2kqZYMx9KR+MWkBpMChFjLukV3wDxnjlkTlXHXsv
/ZI/PZREHfd6ie1ZKbXGsvHjiaovPxOBTmBu73TiMzs1DSNngC9oDdhxznFJL2d/ezQBc0N4Uohn
IRXUlQO+zMxe1sjQKMwsgnCBT1gVSVh8d06JeU6xqKKWGzB/jSPr+IHOX0ixjl4MclT+mfPNDBVh
qWVQxvjFjd2xX4CgdO090F9hLBWEzFeukJFVBmAgmwJBeoByJD9akxoiNvhn9g8L02usanmAjRMH
zuLC7T4s1Eyz+KTGTwvmGhupSPGHoHIftDKopOFYVgDnKGEBCY0JoqrARzCcZKOObtEf/G8VYmKa
s3OPCfBcR6xM4hVYtlfLtzRfvAVtrS6IdN1Vt1E49Cc/XE+gPvC/fxiIk1IngowJpxFyblWytkma
4PsAvqpyU4UQztWvG8bDLb4vcVqMkeyttnfDc2WUQc+C8j6ABeQpS/S8Cax3DE6SeizDo973bFo4
8aud6P4GV9906bNoazlX480stoEjw+++gtiryuCu74zYWikZKL2BPNG494sYeSsRTGZtMgY/6nR1
il5r1tYdK57D8XUrWe7c5r8nPu0YAHYUMSicr15CuMLSxyWU4jH+6b0g//wQ6X07qnq7bA0gCPxu
DByplHze4uuqpb8QzHm6TYDHEafHRPry3us0g+5dLkrz7SBNlJuBP1MEHLQOwNfNc1hFlHgO/0FD
HVio+akfS5e+EQMrhnDSEaZ5DNFhhDnbOZ8HUT2e366z+i+Jn4eXRdsb2OImDsU8GHu7lzHgITr4
phnNtXFjhJLCOabknynmED1YcT8JupPX7AAnEnE9i9IaYwQt+LNLxH9g/eWiqim3xb9SuAi8Ro/S
l7HISB5rFaX9Bl1/KF78i9WwlDr4Ius1qbarSRG6SJoLkkhJ7LduxSaskfOCFEhU9oj6BxYHHfLy
9uIYcBC8VzmvY0wlKpgk/NB+dwgazi0cGm96oGemjerZZNMI/rpckTyWlFvBN0i4YEuEp8FoR+Xh
3Wt7ObpyqePVY7v8cAdsie0wdsUZNPYMwjKJxjtR3cXGudzhHSNtOA0eCPrY/NF2zLxUai/5DsyM
gY5K2ydWg8D6lPxrSi8RlvpqH5GWipSZfcNDs/bkUdglEGEbJvXWAI3Gz5O5YBRrl/IRD70Oor0X
tVstaFin1I3LGLGUlLG7z+JJysoacb10hsMXdsZNAvi+2ECB9cIxiThrPr55GyIDbYtSzd1RzdSF
0yIsJjiiFydfDz0CAj6t5q0hL/7uo+8UxPr17+4OX6Uxg5LHuchmYYWtccegKZ4Z59VCQq+3OROY
GqzH4e2FvOjSeYPpd1h2LG56V9+4R1XDg7y5PXhmL6al+mR+DhSon5g/K1Zk7DzhEnp6eids39pw
sSaE0TyL1FEhC/5aZTMcPablfVbTBOG/uHNtHGjSdnV58wN/4f14Ixr236rChuNoobZ+b7+pvME3
kpu5tzPUEMnIe6QHzH45+eBBC/3yhJhOn+F7tGEkPnWHLrQ1b69/DmBX4x1NrvVdJGBojSal+aPR
DfD2fSujwFg5CFBet6YCb3acZGVQ9BFfH95dOmxPjzApOmrYfxEqtM0ZSoybUoBIt0UBXBDx8nKK
LOt9yD4XtJ8AENz1ezP4S/xU8QhVCAyVOr7kgwMoUQQx+OdKouZRJwnVZQcJPsXCHus18pP+Nlf1
l5fjFRT6R5ynvqJZdq921+IC1IKWo+S9V15b9gm44LB3ioDYHIygS+Pgzu226duPJiTbAJrsTkMF
9EmqTiqZjtoO0dAPKSAzarqZZCmHTbotdT90z+mZijfMcZg1BOIYEAuD9W5iLiKKW6y/0l9iletQ
lXm6jQgpvfLCdS7VpJAHlfs10vuSo+X8VqPtpahCzQJ87mk2qvT5O5zrxMkDPL+D/HDOsh+XwUsb
OvjFrlk+63n4gKGS5/UDEgtLW/zJl69w86GK0bb76TyB9lODmzkA7ggApJRpjN1zUE/jTFjqsiKf
s8gvbDqM2czgKbfLaPfCgeIWEuqMPy7r/RqnejUS/o+M/E8mZ88uw/HzShIi6mH/L4qX1Rj9IpfH
01PGajnh68sV2NP5UcrHk4a9ACvzOrzrJZXTtp6Qb7RryQJiOtBWbKP8LxgOZ+A53OuGkdgkaEsk
K1A6/5oq9tyszXuwEmKZV4AnbwNOXXQWHhwkc7B3InpepxhcH1K2pL1y8EKm8j1gwjD5QNUCbAev
RL5SRLGkbAyYAnIbezSn1as0Oz1WMjCFwC2JDNL/EFQOFkILoDdvqo8+BZbSrYRhX7r9WFiVbmgf
9KtuPHrjAFfZa+Wv0kmeTnA/mDaPW/uS0fOpgRqg30EmvWWMtwwmuKOPby53MVTAQ2Y/m7puWmh+
a3j+u4d4CfpmblyIuvsIcOzBQBceEQkPG9Y7gfXmK2w1sgCG+VMfB5vkIFHcEFXoLC+EH4QZZGGY
9I8gXnX6TEZhwzz+28pxXIgOtZ/jxv7GGgZ91Ga9SZmxbrNIWLcPR/y5p+Ygzb4iLHx8+/fdfGIj
XbNEo57j+cAn+BZGCCI5qTxgXyiPYtcPEjrjPchXL3bmlSK9beGJA0+Q4Bby1H+uiNuHcDBYjlnj
1qHMXmlirAqlpxNr+f1gBqaCn4JeRrnM1cNdStbux90Gev+aDAX8/ELYpFZYnTlU6ZQFZr+0DzvP
Fesk7z336RbjKFAfcB3lK2N6BXEyVcRfuL7LDuhA0h6Z7BzU5RMBVJeyokyv6Rrp0GC+BzpExyG7
RI92Lyr7wt3YOsNcbMinL4XSEMFjJUpDLqkPlp1TBgm5wTWrN9knIkqR2ujNfnW7ybWJnJXUa4vK
ugKnHjdiiucD37F4BRtvSFKa9kaij3cvuCArftZfN8cLmDr+xDbw/aN0I2JrgFNWcuyriq5EujsL
ZyArRd9sIg5a8hrDXPWBN4JqHIYgUFXPKfzwMS0isUUpDo6eggpsaCIwRGR/34PN53q2tEccmCy+
gY61PZIQmXni1XFJOuQMeHb8BTIZf4Wa09A4gchui9aQUx35EQl7I9HXpEpxbjJHXIgUaMqeck9m
RKZdZ82rWEtB+qIbeuf/nLABBe5VZAWxjz2MR683lG2OEflVqvZZIQ/PIx0R7uQYm7dKcQdnQYe8
wFlIP3hVHIx+v0FtRVxb+bHcJ+l3IIzyRgejgiEdQ6SyOCmdbby5zQHsU58ST0oe2SqvX/omQCP0
WCEyO3dguQAnmLNq9n5wWqOPUGXLnvZ42sBKrQtFC5pNm2LFWHgFPuwhCFET188f9PlYGZRS5amy
ZAJPYDNTrLaYBLMLs+HxXX/5ICyCsG1mc3uJ/CVOl7KQ5eioUyZ5XUvz0hRUnGKYqOBPoFtW4klS
Ml1RkUbM9l4TXkSjHqUtqDnin6qllIU9GTzDDtpHaZs1a37oZS+KaoCSMcMlr61MxBwWUERdg89O
N9+3RrdTjSHqGi2naX+HPgXo0HJDM0SmZ4kXut/+1loLyeHedzcHoMweAdqLvOLQXUEyAT5ESvOT
2ztQrdKdxTjXab4a8BQdgkPnxv/i540G+qJ4yirG78FdMZzW8XG2Zsn+xh/LVhP5p/yMQmkcLbFU
BOx3JiSu39z2ZyCRCNrOWfWa+EG7Jkhre1WHFtEnzslEym5rn5QsikpSjz8hpfhY+6kTj9Q/SLBq
pYRXP1u5seMhxwP2/z2QvHrqpMvOe9LQvFlPx3/QHaad9NgBP4KJ1cUHKqmF1ConhpmhpYvwWJeU
1g2a0mVc72lU5H+6X3/bPnUxay9RqMi3BFlcbAQ7j9crEjy5sVnIemzpoa88s1DwQqj2k45MMVfI
loaw+v4JoNLhs8Ohlt9WSH1Z4HpwZ9TtrnjcZ5K6WvKRL4Efu+lmaaQDznfmJ5hUWUD0X3tI1apw
/JzBa3IwsRTSmunHgNGCrFVfS+FrfQhYlLakhLp+mPVOJGyVfQ7LjlOpm9qXHmAYPLAJd6z6ikO+
0MF+QTyJh+KD2weVA1Uk2X9O+jFIQQfyg0dZ2kL2ASXHhebBJEbA+YjfDAyNVFT+g1AcXw+ZjjGu
jyYZ1GFYTPhp3d4qsKSulCdaUqxRIaxJtvpYmMPqP2TC8waDTiQCiQeYRIjGRGAJFEG89o43GUMk
n+pO7DsxK/hX63iFiYXyuC3r+kCvhwpPyoy2EufN/D8rrxQ07GCkTfLrqV2yOsOkteqJoKaBA69k
Bxf40EhcDzH/HzdPcDgCEXjqixJvFHGllJXXDKmT3DxBhN74MZFvbZlu3K/L/WpAlQqBrO1tzmAI
0Ha+BVCMBvyAgpnYH+VeyOq4UkPfG8iwheX+wpOmnf+/rG1hnYkpKcPiMJuJpo7fyPDmp+eOttgP
Bf5avs+MBOolAoKidb3nlAmLT71OGNxN08m8+Byr8VXFnsUIWd3dPu1WiCGvuzU5ruzWCvbqMuvS
zICHSRNpkBjS7+SF8QGnHaDADcxa5mZWmJkT6MWk5LNvLAS1qXsl6ZROsk+cW3W3UqyJ8w3Q/u4+
yB9xSKJ4fLoisnmFIMt/paqSN3Cyeaz1gUwS+3TOdLGq3a9YkMfPayfpJN9me12z0lQch74Ckntt
a6jUcVhcyYTf26cF4LuXT6ouJf+YEMNGlzX5mrM277USLMwgLOZFBv825kXSroRW9sFFex1ldwqY
qRJYbOwhZVuEB0PEpEnkA0t0C4StrM2DeheuGNx1pYxvOkxJw/SXzLIf4kDUD0ABxCNzkZRYtXJw
uZXc2CzUxOuVLTsgvY+wD9PJVX4GbjXC7KcUnYUOKNP+/o8+ED7ddHnv7kH96H4ovO1pHD0Bejcz
XZs7ljEDw7srA8XEKbpMbP/F04TisEE7c+A97VcIo5syctoJXkHMhjl1O0g8jvsaQ7yb9b5wBSZz
tpVOfv266zDwq6ymOFcEjbuzitbDfSQtjEvz0V6c7wViUq0kX4i3k96p5qqUENTdP5MNSCB2ibXs
amsjBn2UWtU8GhQ9JQvEOinfhG1gBNi3uKIdd5XBQhbc8rWTMA6V8wjFfW1pFsxfSw7c8WlZQUcu
6TeQ1QFtTVmIAT0ci/4LfUofsNoVBzY5UtrOg8V+e9kGyGHUfLrYdIuz7PHgDNC+x7UK94DndDY7
RBCBZ2NSFeI/BKI4Vp/XY2Yl3/03Qso9XfZqW3rTCHiwHpgajpTj6Eyd7XLEK4TKDM17AAo+ON5J
hwosxqU7Tl7Pnam18F0ahS22Iz8X/bxaAfVImIt4W4pEyrBfqCRyUtK7rVittK0vSYvKhQJ2EeWK
3XduMVF5BOxNBfCNBKQEgTuP8ulrwgNb4b79lnBQNW0E1MmMC+eHGnv6XifzjOsDTnVTAR0UcE88
MPq64TF/3iG/XUvBQ7lz75Ofb/qo8esdmRiM1V009Uo7wWcH8EjRa/9mTKZCInCJjd2ZAiBT93Tp
y4ckeBUhgzvdoaAjXyOAZKoIkeLbCzjrimgQiC0W2YVrcUWAhID3DjHTRSVvSFkdyYI7sdjJ3hUd
2vwkiI2vH+SVN0htPvnkgIj3I+7fSzdPpKqq+Mc3odhsVOyX/8FttoX7xHEZGfyiu2V1wsNq1Al8
cw6QpiDV/rT5HWpg6YlnNfQ9bLdMuarr3kWb/iF6P1QjyZBmwAGL0SwBeazF9nkFD1vWzJSqrb46
a8p3zThBSfY29i9ZyLztnVk5oKzpTBcWXt8Wa/A20/VQKLsnqPM1CzRrrSGrlNfaIvjRs9z1rjJT
XydtXyMZOKAChCGvuOPwUP0qomps7fHFH4rqbc2J8fO02zvKpNq5LPEc/0ZhB2lsCXhnJd/LYbo8
j4aFmVIiHk1mBx38t1EOCA6L7dqOj5NVqski81BeTJl8RrYnav9gdiHupoqSzEPaWv134x6ajw8K
vjz6xmgucGiJpP7wzi9PGFyTN4N6lH6MYtr8HGncOsfgvNxOQRwcZVJ5b/KtyBrHnoGCCez5Iu+g
5h7bGT06Ax4Tp0XZok+Tmb9QxB4pH3i/0iYm/FKQ4KsVB+U3ntyuIZe/vUVYUeCwmqTzJoH26klX
wgRg8WmGBl3yWdjHSbqxibIA0lu4Zkl02eQLcMYi861VzYxGWCVSxYqU1hnZDuI+bAtn7dR7+Zt7
Lu64ShssUXKrjjF74gtAAUGPgAe07OCPpP6nO/7u6nSPN1414S4OSyPW31hXLNPC2XKfoyEE0b3a
ZScVLFGPB1BfkY7mF9SVZ2C1BRjgk1yzY7jjKURRxzgM844G1BoE3P7gXG+JAjXkGF4qShn5WSl+
1D/tmXdcATcy81pwAftNvycn2YPhYUw/Kr5wq9i9GX1J6l8EMzopUJQLRUwq4KgE8dxSBlCjBXzS
maA3LAmF4qpczM16JmkktqAe2SXrAcfZIZUnjtWj0aSJvFerrsdmMbSEG8GRSiXJPDvUzYdhvWFS
jvpaMD2Gto6UfcMuVXQzLKhYlZ91Ri5vmqOpbLfe0vTDOf9STNzWsUC89iiBZLNakQBU3w0mM3Sy
VqgGAVc+RJK3ITe/c/8aYTNUhC2xSAok/JPB0QcdzN17DzT3aN9tZ7f9WKOAG0f1cTkglVFg4u60
9zOKAXs6stAXrIeEZhBIbn2PCY9TmviH0G5rfnq6vsbDuKwqGQ4wOUcOhqEZGYYXgUIOXFDqalD9
rEpn8b9/zZM/5DHM66GszZZZtVUq+uvIIk04uG5PrRZb/SVEytgPIdvm+84JZmQVYhyLvQi4rmEn
dXTfqsqbfZTwmdNUMSGcfDlnGq/Xi7zlou3WAbehW2Anw1i6+bQGNwo+1pnAiXOYHO6biPdVkaGm
SJphaUgO9pgVk3EKkyHmZ3W5/D5NZDuoiWeVfr28DnT9x0E7Nr+ptn0GqS+fyuvzOwK8ikig4pEr
2H4fn/OYShBPHbIaIQHRsfpQvfk5tDLoSkyUWLyYLi6l0v/1un44TEA0XEwHaieCgI7hD+YpGqnD
WYn4Pm3kmq0pgmQ1eGGY1M+9CJXTs7jyy4jkguKvfAHGp2LZtZ4e5WPENZTsuxlrSepqxV/gaGsM
6M2rSLnrsMjeH+YuUnUEJzCcI7DzYvB2feaI8pAlMClRFkdiV5AOMW023HhSxzTUfGdXWLR+F5bS
qiUFPf0l12zFeAkBxe+siBQARxht+wlLRdEiDKIpWAwVYBnqUpq7glorTXFhnmFVs2EqBa2L1cN+
wWqjlTX/wPRgBgOF3hmbK9T+3xFds3Fx0jo2bMf0VXEPU6TODG7STHYPomjH5/MG1aYyS9nOYXEc
lDeNVezWvI+j+Fez6alYRAxVRVR2M3CAXuaFjXx/v6ifRZMGcOy+jODkKto/qPCxyaLttW7Lf0pK
EwJyckxmjeRj1+uzp9fITL+pUf6sYA3VZYH3apV/yjhbD6FIEEZTqSipmOVV9+0r82pdj5E9DcQ4
YEKOPzaPbxdZd8Da4zssKoXNYI5u5116AcJ0TW5NWNgJ2OhpX9xFjUeBvSycGMIWXs13iC2vNQa2
Dgo0KU4YGyHxvuqcZ/oL1GpFSWvynZ1PEfFMTbrAHbNFR8o/Ni0pZR39BKl5iQ3gpWyMnOu9Q7O7
USymiIl2INLq1AjXlxolruSP6EYOwaGvS9M2Z2R/3U6MVgsNx9/SWInjWMJm+fhfPzusBY5fTr4q
32av8r+nkNqVXowPJOV36+SwKhtynTr5h6u30/ToiXQfg1ErRB+6eoZCuqWViC31sYXOi6ztgA64
yOBrj7LqfE0AWwStcNTnQH1YfoCt2nQPdHudLgMuYcUsM7O4vFIr76NgX6dhKMpyylIWcOE/3uo3
tygFbaKHntJEmL+uW/UWGalVAnQJxpmnoBi3RysxgubxUS5SB63Rsuc/JTBAuBOjL7Y0+wc7WSvE
iMvkKKV8j8ZQo+LyOJ9etkL2kgF9djc7arMQuOl2e9Pe+COkTRWfz3DDhjH6kiMij2qvKDhNc4wj
yqBCJus1OZ8UGd4ttaPyskFdliVzHpvl1JC6RTrLGeRJK6r3HheGUhLoikjAJQH7/hC+su2aC6Y8
uwh29LNNMxaS+UMVr/Fqh0G87t2gKcBNzQbeL5ugSdvOL1I0Y+tJxU3KFsXTzltHHKfdp2RH5J98
yT54exFcx4aXDbuWqf1kfOp0vZ+PMZCVmX3PfCeP+YstiUfR/f3xhbufyLH6gbkg34ra/u3WpCzR
nevOoUwma302IE9tASqnE+w8vc6tgtfqbQ8S3coFTHcJzFt6y3+qYIA3TAHXQb1d3g2rSoIuz+ST
aLbE6bo2k4JVm/O4X9omjI3bEOPJ9lwoQTn0wwlYlV+b9AWHHYnn6jGALlgNr4+yqRVHChl9Ml5j
JbldDBzzVljK6E3Ddj22t+xU3G5FYPhzj4C4mGzdOLG85eg4bgeLqJsHP6p9OGwK1aCO7Lbizul+
qeoYEiM3LZRePPJmpzodFGQ0x6ZsoaTqmPh2WPsBv9G48T2aWcS+Y4kIZp5QiI8p2nAZdudUAV0s
Nt5/5zWMRSboTrzCE18JH/yXzDdcyLKJFU83iZN7uz+39EgIyRzL17D6JnWYOf5bbEEO0KKnN28M
1N/MXaFsjsFN+zALljDLp9XFncHaI6a0cLmkVynPo/N5SqU8AZVEpYa0fSKxJJjc367Z4Wtnrrbz
pwo3PcHHVMmG5y2/Them+o0+lqWCGSke+IZ3vC8FKbXZnyD8mdCENrUhQJkUej0KN8BJVrme7kO2
8TiUza/4qYApr6D54TIaZ4IlKYKU8zynuFoyz9u0RV8nsdtrkPrfWeg9BO2CGjOIqif9DblBVAki
yhwYNh2jH3su5hifNCEBSOL4P9binzcrmzO5ZsUfeRfhcY+0Ywi4UHPpxdgOLo0ge38JdQFjUNxl
/0iQP9LHKyqQN103PTUCsDKzGyRWpuvYg/UNkpZux3tT4Uhn4dFDBwJ29DXdNHO8GzIrg7EbTQ9U
stdR/ih5la1GLchTQMnFR0sNRDBogQc56CkhWIpMq64oqEPJR3wV6ih4E6IDiVLN+4nsbpbTqecq
Vcz/8tLT15Dzk6XaOIPp812k7uuy9Sw6QTXbK7jGmiB3OZ7L8NjMS/DUXx1hDmbu5wuCJKvcTnC7
YXWtBmkKrihvnnpN5uZcdQ3mgF6ZsVP5HTn0oP69g4awVXwxdlQZDeOAF+zMoC0rLDsPMBGxBY3U
mp5MF4x8IbdkWAKBgETAg2g7dyHUgcT7iH/c9ZvKjFnCUDoG7UMef647VhSTWWlc55Sggb03B9Oz
qwHWyVa1dmsn0cZy40FMAOym+Miy3TtKzeOP+ne2Q9yVrpa3jTi3su/Ekd9GKkc6/VuX1qVYtdVu
Y8TBjENCe7+gFEc0i7PdB4xof/laFnKGUxxx4eUy9G07tEeTY6ZFBPRYTrepIwmgi/n0e32Ak4XU
jK1059eVo07EOrcRRlqG6wGiZR7nqXRLoDyn0fFr6ltMdxuSZy9SBCZW0f80Qdt+0C6LlAhZjqZK
oD3evWgRRO4AAn75Ky8h4CxNKz4Q/1UvrqQqTwIRHub1dZT6YyygQBPcCX45e7T8HlCq+dE2w139
3x8CjxzSRvoZAuERs2SP5KgdPUFfdegpBI3h3TKV82MfLnbvHPOCCohIfgABm+AIt/q8gPxLkpfW
quP8SUMc+XUvnlaJFm8QLSwyhJg/Hv06iiq33DBwzEftzdUTRaf1ydWyBs7M5aTPwYn6UoOmWG6C
wm8qv9hROdmg/HncwO1xvI9lzhNVHhHSONuvfEzHCCzzKZUHIJWvzc3izWn0EAB+xmhDeETSrpC3
NFsneSEngZqNj2dbYhb55kAIl0Hl9nlgvNsR6Rl6QJ403V5JhkVhPSeDm6esZZmUxY18j1ifTDcv
2U6t0M+eqFdV1mrHBht/I+8VINQu61VDi9r3drQeiAMiwB6HFAdqcXhoiA2XG0hLmQRI5QN3hCgU
6LsNcz0vA9oWENoTRi7xGyYEbMYO2c17RHMC1bYIgSquobEySzwlTsZNCK7vCBeRw+TLpQWiVub7
FLmqfgTglFPtI3s2dwBtJvrJEEwIQtGLJOtOq7InVzL0iHGMmHW8Ned8YlWXiYde73VfPVOjM/ul
aLo5QAIik3crcvSVqKIUlJY7gsgqrNqTXgmPcCfnpH2Sj2U8SLR/Sd8iq0bIJc8mco8Vt2hG2iK3
rcapYDkB1bp5QsStBmfdHjHuLUb3KSKZl7qX2DX6oDUAl2sbC0mOrgBmmylrTtmZPGBCgaPc9hkI
0p8HHDwyjNb/5tqIaRlOP/Ke0kIyx7TooHd4ZCOaUzlAUoj/7Q0YEIM4uboIJfRVZD30KYhfGu3y
YgzNn/eZSJn9Ibr4s6XDfBUhesVn57PAh1JIpZNn6PUhGe126eoQ1EeryJ+sNBABs0UAWk5rdchf
eZf2TvFGJkkBkk1cDDyY7ZJeWmWEIyDSRBI9csWW55Q+MbRjPlYiBeeCa/ujdYLehtK2GlWavKil
zR24IBNTABB8LjZU+Dnts7XbrcsQOIQ2zsONLgHQ5A6vK0QU2aKxrCpqBW+dxwvhEsZO1eryiL2r
i7+XroXur5ISKd0qdn6fGzON/7HAmzdSJ3Qa+2dWDExF7tVSHds8yhbN6u+MdURwkpkTvOGwlpnp
Bg16aQIkOIRkVG/Gy7meoSWCtbgQDSc+Ml3QAwcwOG/xBrC96StSltGAIJJOD5jtxMvxv4vVhIiF
8YVBmsaCV4cMLTSQkro+sbTr1mt9dMFCfRuyB4EVOXJ7iAhObJ8QQ9XuZ3Pwn1dOI2VKU3HX0mIF
TcRpN5mMvTFm8qwyI1ORSOZzWwUGmDQBv5EGZLMRAEGKOv8210dzRBhDb1MA/8xkw/vbBlwKayH9
L0UztGsh32D+09w307myY9x9UYmcRGSfLzM3gS+Vn/duNENBqdoWEKUsKSHOgyaRNj46tMXdI0X5
OC9UR8CW18c4GM/D2FJs7Oi9CwssOUdczuPPssE6k2mCR/LB9xQLxeExaFx7Br7sVjbqcCgvYPFA
9U1J6RId/vfq2rNT5wOK/SIwPf2kIkFW1jzi0ONlxr369iq1PJXn+eE+ovipEkVJvw9Cy0B8IfOs
SZGdBaOVN4LxWNvLbbv5pFk5GzLTtVK45mzecG8lHwW2E+RCWENN+wW97po8AQfRRypuqYWeNpWq
aOZaU3b+hlZVCKJWyepsNgpiLF0tDVExvS3JD9tfesFT8Ka2cVAkSZYWWT9PO/EtOm2aa4Jn1tiv
bR/nvHVDSaqqHNk1yYrIDh0AboljfoOjdciWpi4qWB0nlLvtZJBa1qdZtJo+npanQKmCe9aYBEZg
7D0vBQVm6t/r+7rnkywhTjCc/tmSO6h3xp3HcUXfwk5N+fBx5NMz8cr9FS3JYXMnczUjS9zjQaJO
YfT87bjXvnzBTK/vIYz8C76uIy91rWPvwHRwUqEDLD0YSpao2W5VGfd+lfCDvKLBm9sqVy4rsjmv
IA48vU4hTRhia6ylNi3cn5uPAO0rkzlZ4G/EKRpqQjW3pW68jiZrq2SglrcJ2izirchgTO5JIa1M
RSjkVyfAe0M99rQCOPZXZg5gYraHB2Fou9RSFfDQMV5ttOENOGKQeQM9bhCVBY3NCXGCGSDU14MA
wkVHofwIkllNTTyZfOG1b/Jm/kbpq5OQC4gSWyhs/8tR69XPwy1xhNmP7UVrz//c7fxAdo18y98i
Wsa2DLYiCy6EkSHe7Z33SizH18XtgrlQ0KTHec/Ko8rB+EzntGESGnf4nZiIwhVBAFCI8ObXlT1z
IM01s4oLeApaAtyDkkgJiPeinQMJcFg0D+Ellw0tJwMTMaIaCOVXjqVgQIQDhkiRjUPFMLq7YR9D
PmdhTePp5j4dAvAJ9EW4zoXL62YssB8W5lMza2TUcaCWB9dJUTACOYvKAdxrZPK6QYLLK3RVfkqR
PAYXgtQm5rMbMOeFrMUzZOQSqaN+CHpvs71QMN+CslyW3jTKyp9ODmYxBjXruFk5bn6HQW6cFmkG
/fpYnoy+zv3EpIkWbXHPuluMT0Fwo1e1JTivMHzBqt1kcR7ZRolietlWqZOhGcqBOazfYtbPQSNn
arR9flKaaLmm5kzXC4JrHGlfQgg6KY0fnx9q22X58MsOBRilYGhF5USnsOiczL/TQdybwcY/+rDk
4QG7Q3sBGVS0xO7JO3DmlyQzXu7ML/vu44eUUdYyFofLVuSROfzT+qKvShn8+SdX8y/0IyIy7bJj
ByWouwl0gXsDCtfwGY+16uLzm+QDhxsNo8T74TQjY1PBHv47Tpe4EKp2QUFNEJFCfucNK3Z9faTT
IPlw1jd8rT4Pa/JAFcnGLZ5woVyoimjWGQ7UoSH2GCxVG7GM1qX6O98fTxCcv7TrPA0M391NUL0T
KbkUNtosCrSRGXI7d0GDdhpFkvS30zVwbIT6EEqLnVRwuLNCoy5c4iRAV3bbNB7ASPxb1HDNlkqD
IP1siUYuQOpbG9QLeRf0dLXenr9jHfkJk3oWTomGg0iQxZ8TL0SF3m/J6tLHbW1xms70y7WYaog3
44EGwIpCJFS9PpOjcfDhZB5oTFRsQ9ltsBjGjg7kRkC5OaFvZ0qkNdT8QeudYhEYo65US9XfcC8Z
j6sch0XPeB1W7vZ/hlZx4c2qdFmS/5kSMxiNTP9KTo7xeNKUYjJ92EeEIR21wSL7ZauFmJXttuOx
gw/sdFI5c9qWubkreBmlRUgVXaVpN2kzIKwh22oEY9vGt2sKvLyNUjVxDCihOsvM83O0mvyFkChn
n012UB4JAiiLe7oDlH/h0fk4nh6LMaoYjK6MZxq04l4nescfqakADf9LS0uFpKa7u/sTxUAlTWVt
/2GtH+u95fph0AiNN96e8X3scfeNY4cyAlUmS02gKOuSuGWsmmTXa56v9zCVfKVVlfxa1ITwOM3x
k/7EI1PDBFg9ibt/c/4LIwt1zaSYjlbFf8mOYDIgtB2W34J046q2abJu4T/A5oiPgOuqw+RxmNst
NLK4N06myZnszy+OcEznrjOw/NuwYc119M2sGbQzkmrMWCUXZ69qt2qlL4Q0U6XZfNSoqBVNITt4
oqQy9qlrsRhwslHsubbZBC1OLhuL1zwqvjo3/tv1tYgfqZLDonOgBbxLKPeQ+lTlyaL15zJ1tUyQ
/fUHXtAzvuFqeTNK+66qdGLNiCf6ARDaVgI6Rt/hw0wxkDaHPNxE2jCi++btDCfK90CylwIUmdIF
oKcYRSr0suaXQSvVQlXFCWgyJjs9prOCNCcr/K36lXFjhf6WnKG5dWZC5DyDwnN5YuIOF/HNSPjt
ZF7hTZYXSY0+F/sFGHGC54XtJfKA4SEdsmn6SKhma0xIbSZmDudnU7lknMJtcCk0S2gFjmA2YqkQ
O7I+Kkpndo7x4r5NdlQ4I+Kq+zcbIMda4Ehaq0p5Pj+OIncnRy8fXpzcQToBp9amIHqc0s1xlD7n
t5LiqCkBYVRxtYiDtratR+40Pp4FWSWCVImBFKmd2nMeNgfg+sGpgjkg1z++gzXDsjW/6a5qBTiE
wtlYkGaKrO7LaSxghEbslSUpB1MTSEC8pTfKVYVNqf6Lb+Rh+e+h6rPSmBKRoExQSzMdSPgD00Wm
yd2FZsdCleaqQWc1ui02VvfnoLb+v07eDtpR3LXy+F5k48pWW8NNY0olt75WiOaiXOrKTtSgrZX6
RtpmXiQTWoTbQ9wjO/FeDlFCjzLtlnJlMED70qgLK9dVhZC4xfdY1Y4WXnJn7iFm/sI6vwXfd8qN
yFXJWBudBUWFqUbKZj+ZZABrXI6jPhRi7E0Bs1lE9T8KQee95DbCv9n0rjz+KEedymuUkcqS8t50
jTmwl5E9WrCMry1Tpo6gzHocMvOMGWdKumIAr7UFosyf5zW3JaV5DQszMaWRYdNoaVp6HsiuZ0iv
7I1yjXaW3XfCxV+sIVWG7cpJfx/s1DQA9IOIVnhxlehM8HkxQXnxP2PVBj+CsylzEg33gq8g2Nht
BoUhlZfFry45taTSmN3dlxUGQjtg2EXa7BQiIGbwt4Rr6sGNt+1Mc6i10TP7PFNH4DnqVyMIQmxd
a6BIxLyokyOeBvX4hsMyC3nc0eaZfL9cm/PgJBtHQLppPcMWaoxT8BKweqpOl+3YDh74Gl5CqUbU
Zf9YNaL3XQ7m3yO3R0XIy1ui1LaRyE4K17nuVi57O0jv3mANWqO4VJ9GmylzuNk6FA8LasdMZLFg
+hV/sxwdT+bsoxyCYVGMDySeV0CzjbBtH2Qpnq3qi9Fi+fExTDrnIQTaRkgAaf3QXjqKcdO+abiv
JLdetnyFfpm8VpRr8uSkzzwEBIJOqL2gAEa5pq1e1WFcnvifwq7v5IvgldzHS+2kYHJga87Ca+VQ
PaKcMuRJjKGWOdAwqVzdi2H3twJLHUpmYBbRdhvP0QwhaLcsGUV0kn+G8gO/boNOCakUtFGc9eiO
vGx6AEXhDAcTZCLIPtVfZ3oqI1PZYu58FnN2nJf9dZDP2qRyLao+of72xb3h6AN4IJt4rKi5fWq9
B4BjeqeA2X5y/2X8ntwPYaalKGR92OYJrHj7Tm33AEHyYGK3XySixzzirF+NzI9NtgcMZ6ZLsbgw
Px2xn22RcUoEEPYs2S58K4byzlAYgo0RpaZGtB+/76ipZQaz2D11Z6fmDucmeeavwEvdxvyw6HEb
JWEBUjf3KHe/F9vnr7UgLcQEfXdeGQ817w/i1PPteXXlFcYCssDgKoyc5FPU8A1wpWLRA/+WLRKr
PG+FZ8yO7yc4vwgkFRC/6/y3nMFf9N0qH1S/Cq3mePnzQ7vwnVqqBKEU2sx2lI8pmZbtBPymbTcj
sWo2AP+DirijRv+Y6xggyBSIw+C4hWYfy2yRF6YPyWN2jU39iJJqcmMPmJxjJketac175AkfqJ7Y
g5FcgQgcG0Afsq1KiK/IJMJ1f7e+H04SFeF7fkCNrTO1B0AtbgJM+VF6EnhQWRY20R5lMWGlHvem
72buqbwb1wn/P+fakVcyB+7SVBqajQyNvWNyJAbSSEyRoyBI1wvWLvMBpfiYpMROCB7al0LH5Q3L
k4O/gWRZIPEL9t96Rwg51XiGmIi2/mivwRIWTiS9SD0WpWfJqPHQMOJ7XKVSg6PFT8PKZRNmmWhs
xhqkMxlwR5dJFxf6EV/e1rQj7lmgr7LaWbNK8BjdMf7XblxhFjm3Is6j0OyN3OMZm78KRLivuJNy
mfaYDTadixlNDwBuoEhR3epykLKXSnkA8U6c5+T4ra3zWqCv876OX9jrqF+5imh50VgL72xDFF3x
UkvIkEJBvg4QaxFtOPrvsq/ak6H9TT7cjBITFNTPt9JdcPWYua+R+heB+x2iSDKrj4NPo4b6zuTj
6nKGzstMguhuX89bsUSCc15j+gxiPahiLQsPSHkn9ShTZtynpvb2VannXwxbfkhObugzZ2fZNqQR
5G25dGgn5ybqfITy9xRcJCB1ifqZtul12JQH0A4U7ZIGUYKZlkWG+A2CeEb8EYru4BySF04Y1YNA
N3TZwbBEO2R1nTTcVr2Ys7Cj6JI4ASUiz4ZiEa807vWBbJRYZj3q/ZEWs2fa6Z2ldupNqtf/Rl6O
5ui8bQY068lL5hMD4Hn5fQeLvhqGn950md4/CJuXXhYnX2GOyngKWcYkqiDIhVf9CoSX/ZpBjfM/
E0K1BeD8RGbKKhOW0hIZpbaWib0/ehx5fWRVtej2r0+IgCDz0bfArmZHVCJ0Fcgc6YivEm7IYG5n
oTa/255eMkA+A63SKhNuaFkVSdLoqYXHhsdlS6QYEtIR4ykc8SlJfuhJxKOG5agMgNFwyH37nsWS
12wCjE9YxknObdL4ImAkNwwflWX0Xf2JOFRKEe/CqSlmXFVQQWtOl8KZjNJAS7JNvorLPr+/5CSM
UO+VpV77z0qWNycgW2lQUtDvcqFs1nH2ixXqIM3mlO+9tgy0qjkHYXdj4/JVSZtRau1c7nQRd0Wz
3RmUkvc3SV1PPHu7AbtfCKEUjozgYATcj81cbAPxPflzorsJMFcHYOhI6dl5nF66c0c2adSM5xIi
UqaeM55ivb9M+Om+C1vVcQ0Fx7vHwn2v1lzHth2Mgk/qjGqj9qOQKB7CbwPSDJF8zhoYMq7izyuo
MWC49IivoaUWy4YGD40LboL4WPI67aIy9fkeu3C6qK0roUzSWSaXqTTcMp/3eArmhPukAM78Svim
W7SHPP7tQqr9mBFolIsjb2G3ObOXmO77zxOpHdx5U7ashqFrrhdFB6UTSA8AOGQEonl7whiz24HL
eSNJtYNX+PxrWvx1W86FqEz4vRc5LgdOhUF1QJpQPxC07WkxaaF4J/uSENiBvTFMRmv31p67j1ot
SbdnpVzfrTA0uBequEyEI79E1gkz0sKGHLSi9/ViBYNWu/5sVCJ/7Ys8alau0TjJQ/6XhGGSlf9t
Q095ZK0YqLOpdteH8h2q+yLHJT74zcc+JpOBTC4d0lo2ImIBFQgq2O4GVYDdYgfU69g82LaIOXRu
w155ooqfjTpUJDZKVfju2BtavenUFwIcb5JmdDZGdLLlAwiDYRw9iUdtRjGgpEaDQIfeEytq/6Q6
1DdYFGaY2OacFJssROL8NtoBmAC09NcWtGSrRfZgOSOpTnDuSyA9Ny/wR7VFGeFoKyCZ/mCCVcer
1QHAwLOSn6Zt3bvMk8i7TzD8zMSRPrORbtYI3sEIR5XLQ6BC17Fk7IEe+UTJ0RbV2bE8fDjY49MZ
krt0+IU0NCuLvth11xBsT2dJl6R/vHdZhEu8d11McK3IHhHLjFWNNAJaUbuh12lk6TWtKqA868I+
dA3g34xxpiB2NKrUo4XOSoso9lro3v3SPTtwtYtZ0rWrVGt+TlKC2TeGWPG9GZD7aT7DYCpf3ZoR
DyFXoXwzOHGtykswrklvwpnp6HbXPrwmh0rpvjIy5hJ5AE3H0b4Qc+7au1BjuCdSeH0Pe2Q5vHYs
+1RE+ksj3tBt5N5RQ3WSx6w5KANZxfpJFFo/1GfcxGTPYiYx7a6slvvoJoee9Es7BBUSyoN4Oy6M
Q0tOctVBA04aqkixFmu2gi4xK/xo3eX+mKW9Q7PdOjAznbHa9ujwSOmkrHGIWP5jkNgGtSH7dqlR
AMJGLk8+RJJEW1srSzo4AuK/ZzXLe2xLW8C6R/StG9An3dU4Vh3d0yrULszbvWtnAx8khsIuPZWj
vSdiTzLHjDr5Z8+ZexjE0+ffh+hKYBKcAT+zTm0DTXQqQHaAEgPNWkCNS9ba9t5z52Ez2tt7JrTq
niFvkuzh70mu9oZw+EEPqKDH9ASRYeC3OgnmNODTd5aurXcY+QS6XXtLSGbYRlzmidnhjYWdU9Pc
MARxqnkj59jf2nnBf3SMmCrFdifTl4xkGkeEak9JEFYOkEBLTvsAPVM4kI6qlBPQDfjFJmvHWMaj
OGRYlOq6qB+qYuM5oOsjFrQvEyF6yi+YtzuKqUzMIlpCL3JMN0hSfaDeFLNf2cJP3xM9aLRn89Nv
GkdZTBscm4fqVyVLUUJVxkFkd9UFj9b7OkARGnty3icnJtTvXYtB7xunEPLcZRYAIR1GjUMUICth
K006NRmIa+mGDSjZg6sfGeOfaLCa1LozpP6Z8C8RCaxphbk1so7tfkLANO6Kxm7HhmHzTHjPTygq
nmOk4I1u22yURmsG/UTKAtXt08eaPyQxNsEYKiD1qqyfjwBtHG9yUDnHE1jwmPEHqiiwJ5l7DbB6
opDq577rzrYZYns8Dl9HeE61boGl5vO6bgzys5vpxYvZKhTs8I6KS3F4Pg9QtGc2dZ0ctx3Qw1aq
pMrRCFj0yhW7p3eajkMVhtWmCdPFMTrLSl1qpNU6ov5m2vkgDZ9qxk8wfi6oLGKIPPFwOI2OnFre
VkfpcKd5lwGsuqGI0UAk2eKemM98EVmZI333zbZOb4FHWUZOlzTucv59OKh++SKqUktlOzc5Zmw3
KGXHVwt09BJZeDWwADuA3IHbResC5zSYBeBI2gXZb+yrGuYgxyedgBucsehOfOr5R62Y1EjWXYGO
ClKJ19/TMuRd9M5X/DG4gDumRentpB90kYf54N18Wugc0peO93FbodjqwdPKdF+xQeCBxtXHmjlV
neYvj8YC1PLOP7EBZZ9i4EpNQ8wYr8yxTAbUW494auYP81RZfYPH5H+umpKdjAzeQtleIzN4X0si
//0fK7hxxCfTEADvOuLrxXRKv/Dd5+6f2d7w4nBVnUWsTi609LbpBO1G7hWzgZ+rjQGFMUnYn6Tv
fpB5K+5iL928yWfQb7zERJHgbYDkUqSauOeGOhx5RGmukGyrYaa8ULO1j3Zoit+FBIWoFlXeOliD
m1Sa4423TtscoAz3IzbAEeVGepJ2u1yyo8Ze0vdHBPQD5JIXbD6jFshHyjsd47uSGSgefeFapv7/
05/dN7I+RQIkapbOHAJI45X7KJTNlc7H1M1Flg+tpAvR3iLvP5iIRhIh8jKWcy8n5I4KrFW0ULE1
+WhjUmuZGEwqaKhg5ENAEo6+3OMXQbgXWC8c13io41vqwwKEA96+yKN/Bz9hRmVQBMC1nCJR1ZFA
GfzIhOSlLD2JratflU41x0d/Ch3NXzDepvuzTl7T2lTzW8BdmOoo3uwOXt7HonP2nsqJjVsSXtG6
+Ca+4gXS+4iD6/CXkUxeLnFG30e/CKkYbX7D91MNwbKbjEoC42GWbqI38wjH9ZXxKDeYPuzs3zJk
kyBCHVoGUdSXO+l2LdkYIyFAzCprJim/LCwZyJgSAH/FYQvP+AsjZ4pg5IlEbw6d3Y0h2RD2mIVQ
si/8WQwB2PDBBZOH+q4iVklQ86NnaL11p8wqOt3uGkcvwKVl9rwy1xaYAm3j9MxKjVGhWMgh3Pcb
l/MBf0mvFTBtg88Z+dUgeWKNMkqmwShOPaR9JMva6tsvG62xwBAXdxlevE/9mzAyX0SjM+Kqwycn
206BWu5xRqYnqytKf/GfmaHTMh9rWS+Wwva8KXZKfTgCKqYi8/cRLsDwA+VDZEY1XXWVN8pdPdRz
6I0A7sTbd6TRhSUraNLKnSR5c3OrVY62RWcnsyN5Opsf8EjQwHbz0lHYWvlmsQPlBANLqMByYbEK
KcHmIxRGCYOM0npND+T86g6TJSn5fzhFI8rSodHnSkTVherLLcOKXbsTOzcvoLNnKRMt6qaq4aig
09VDVLG3gfgwL0sVNtLum3GxmnwkEfUbhr0u84EE7npiX1rUlJnveechJP3w2uzKJ0RP0JL6jtNh
EXAhfACQg7p+HcSEtUC+ckZ7H/EWktw7o7yPkArufeZLZKynZeHhwKW3jrNnz9O9UrPd2GnyLcRD
ygwdgwh2SEsBXH7aWeNnRkUlD5J5QhXzx/UYRiAVYwNgPhLw9cvBQDbojET7WdZhDS3yQalTJSyj
D8TkAn6Me6QBvGj1cOnsH8n+bNLelWok/jKu728SxEXF8lLaPW+xsFYV4kIGiMgVe8AIkz7x8CUs
ua0UYmmw5mt+wvrc457ImMPXvnfdJ7PuF0DoJk8UWjf6Fy1gIkPTbrwehiRW2wY53WIoiAofzsI5
w9VBTHCZcq8XSe0HK32BJJB3/+rH+fDVS6w1Kc3O2FUf7agHZSCCvC1Pc+5U9f1PUzUWTB/4c4RX
JiSqtuAOyR2RYKgdJ5x1TU3WMvBpIPlAvbnBjHMX6asmvWtA+ZqB77kTvF2EkPknnFmmRt4U9UG+
TzDZBaqYXlwEsBmAuf1UugD2GV14u0c5Ta5dZxPTkxdfaPN9smtmPk6XeEektAdsonWdCpR0mOTZ
Mc4W+ekqcz2cpFAOtqTgKqDPrKej8a3I5VTZNYXpz6LLm47595vyMkJ5VLezyYWjJRjyvjx2mja7
JHu5wE3cw7X7lt70ybfqCWdhLClBRLSfEYbN0h4yWINey+Zxek9y8/4l/RheLIhWPcbtEqPUrOO+
48JunfEFO8YkUWjqqLBFOsGSVAJ2PdwFnpD+fvYp12wmtRjGSCFmDmRSqBrytGaPqdYu52HlFsS6
pM5LrZ1W2Tcq9jFRQR4hWWWqhNJeIwosFtLMZOL6KolVfhJax7/fsf/RkL5sZx+S4QTy4Wk3VPRz
9YDc4Pd4qsOSvIsn4FZWsWyEzQW9DU9rrF/5U0FkHCsPuSCeBn5rwzu0dr61C10h8K5LXB9fHfGB
qERAsS28/hKaqC6UaAku+l+7AvBkmvrDXgx6tOGgp2U3AWbSe6fP8JkwGSWRchMGU9FGTEcJAxHG
fF34cZUpGSmpuWPLKpvnpgC2GFP/CBIuF5qpku38Px26/12WSkwwbCd+SWt2XNJheekA7y2BPNMI
WnsJHA0x+EV6YiOoiBRYjmeQjhoSaPzc8e87bkA+YkEHKGAFr7jT+c/jezzN9mQ7lqRygXwqrDeY
G4UrO4/LGabtRWaEjP2WZXhOsQZ7Zy2cVfSSohlWmw+0Llsc3X7EeCjB6FWqnIWeT3VXfffbfBMW
cmemaarhjzN3OrGFexp4q2MjfydBVxKBjoevQLjN47LflT24/j+CpVHtKDZliWHVzswpCZQ9xz/S
whM21VvgJvF6vraaQiIZ9np4l0wf5q6afeRGqKalf3r3l75vu+XgOX7MkUi2VDVDqnl+0Q/NEY/G
SpwNBsZysvn1uuybLVvFPorYprAG3UTjfJE3cFPCbpbHKxojJNkXVt1Rn+sg0T9QyYhOp9bjfOHI
FS7cawdAIEVHG+yzauFwHTscdLjQ2Q+0Ic0uZ2Vr5Igoou1cayJyIvdm5vmZhcPkcCy1W/wi6stD
8dU0y+/fFZBN4Ow2QQoZdZHDI6fkeRwm7JVCxF1ueOm0jaLBMOReMScq7/2YVbLo0FOmJ5pCYxUB
sNTs6lf6btCk3IikPE6UBl6RecLlyvQKZrh5J08WAizIh0ajl+RoVaHwkL3yZ9GKmavz5waA0yNx
N03SWpHrVh4YpqGLbCZwQHjTxxjHF28P6vdjVpvWkilxOrtddz2NZDumoFPtI2VES0Pmnx2g0MQL
FPzjE7sdtVrSUr99OcgodDGT+2dxxjx4ZKV5Y08gYI/2O0yfzf8IpQe3t3jZP0tZy7Z+awo292+M
a3WU6Q7tElmcf0azBxcrb34em+jL2BwTntdDYfe1C9bZ4Sv+y2PrGht5sJiZfVrFBJHVsAwx8uNh
9aQHvuzgNowo1mncpkJ3jJLDF+UsNPLN47jC3aot0IEORQjqPVEpk0nsGr2JgROSvVkHM6RaGfzi
t4lPPjohl2ks1oNWB1+2Piche7fr77DzZdWxeCAPVfnzHl8BOtCPhwyJNer7iQXceYmdBLxn16ef
RUTRXVqJkkWbOqEPAaZJl+3+YFjV3AhI5jp5lIm3K1yjO6LNdEI4/yivI93W6C1gRxchgNLstAS5
oKpCl+2k6FKuDKQNmdeSYGmBb2wb8ixPTugbcdHfAGfcVzMdTK+O3PeprG2V2Yyxw13qrWjymMzE
C2ygpyWNaZIg7/V+f9PV6AXQDMjHboE3UD+qdCMdc/3cXO0PvVNIKe1bonRvzm7+sPuQva0ct8TS
2btDnIy1LvBi/K2hMTgeyHciXDkknUAHwEL+ATiOwu7rSC8d4qVNKtEFrgnSrsiJIxLZRD+oKMW0
RRXInTfgBGv+A0jN+a7Z4SoeKOwNGcXdPdXd7NROBbQdWs+a9YaI2mVVS4mSFuRY0ZJFDgyrR3cc
7iA5zuW7VRSuJ98piMkOpDU/hIrDgijOZF1qy++sSje6QDa1vBwOwwwCWW0uR3px7ZBkSiyIp16X
+BBMQKhyNby3Dgoywg7skUjIBZ7pLXYJs0uhyQCgDBl4uYzctDO3d0e8BpaE8mj51bcYhy9jlLNb
a+63KNpqRzNwbAuZik+ICg84W9awPAfxzVvcInL3/cR/bOhXUHwDS6oKjR4dYHldLMEeIUFL4K1s
SoAETEZfdp0cHZmmehTTnDDwyeRGK5KYqHF13M7gOWwGWsasTSnD6ziTrvBbkvfu2ly6ZmRqr8aZ
24TWuPYLTzN6niYcInPBCQ61LZBT6aBdG8iBSRDWIZDwwur9BFmv3ZaP8/p64KkybgiT7X1Mm65z
urlwQcYKtRIrPFlzbcNHmHvOo8Adb87VXonw2g/hicaQqJ0bDlMJM/bmKFIUCYs1JJwElMCJd7xc
pLeCQp0ax1lZYkQLMuzLI6LY6nF8dMUq2lAiFUL4SDXVjYcilu9AJ1mUn8k9/up1TLNADH7OpYG4
6cUptpm04c7ubo5/+b0OaeFAOH5Bz9VqRXJjPV+br6Vv3sppNKKdFRuGsItbJisKBwuCgV5aCVm5
Yzx5vxRwSEefXBFjyAzLvBhIjEQlA26XgcIAdFgXF46MpBmuDXmQZjUh6c/Mb2dO6icfcQY11Oa3
EFXiOmemABKw/7RIIPsZuEGw9vLlfevi9dnmIztckgUM/uxii+EUd1k2CnETpS32ar+RN4llwwRO
nnOH3vAs9yu/6AHj+K/423D7pz3/gnaEs+cFReuZ9K9GIsHcI4w7uQJ28BDl+o10d4qqQH8/1gml
xb6b2JMCKluA20fTiuZSTU/2zySFZNt153WLhUy9JaJAkcg2yAq/HZorV2rspWcK7R009YhwiWo8
7/2basNAU5iKr9qYj7u069lahPUwNu3V4/fELP6KLGwPX/fmm7knQzw4z/if/h7JsJ1XhFqTc3xn
gWoJXhwvMG03xAJDbGPZVGGnS4YjeZIdejWxH5uLT13auuNV4encSG3g4MzwFDKp1oIFCHzOMqH3
mAK+qgaHPVMsfz46GFk+1LT5N2oL+6y6YQeZccibyWJyEhWD62WQS4dxuv4wh4ulmF7JzCYDHPaX
5T1Z2gUadKIISv5T5OjkTlaH7PnHWylVrXpTfLwZ/pKMUEWlAgwP5Vy55aDfZ370oFP7qMp08sOM
UskTBeYnXIcyyUNw7oARn8p1+WJu1uhcQK30wKyC0XYsOCCzSDlgxMTOnYt1zkG3vZvbvre6kpTR
HGDHblfcdv7V71MmVPwnflJjWXRHmQr9ZJzyUBhAgxLfExhkUH6SnuiYGLvvqR7bXl1g+6MYFLfn
b1muC0OnFqrY7uKX5o68ta3OTSfQ4lmgXK/bxNLeBx2YfuGOg8AAHCMFTrIDNzsJbn7a00MByK9t
ATPIPZoeSzuW8N5+DY0uiSXorRdy+uhyU4E9FeF2YWzUlaOyCkUrk6N6ddaYBcCzF1erZXSfR80A
7KaS8jDZhjnBKolDp4msYgYU+RwSp/j1WiQB5l6d6egnIK/bpIwy8SJbo2xAVBBY/7bBFf4zIjjv
bcWz9JBmI66U4jWbxGW3nLZo6eZSTUIG61W0+BD0dTIjCzbMrVA7qf5yVO+1LwOoW/qbHkxCbhps
iB3gwbsOfg73Osd46W2e/zMIHPCYEwdzuru1mRYCG4YC9hl529qAEMgPsaN/RVj9k1ftkiuX5gMN
2M/fufKQLYGxXdM4asZ2YPnFSgWYNB+hBKWlUXXTMTMSOccqkHDjMuKBA8nlwnfAlgRgd95JNNre
Pvj8TX2VZyxvv12W3t1C245dFjRNiHJ7pM5bTkCHXLpp3QPmSWhu5xCrCnRYcoovdBFfkM5g1FLz
CMM7LUIFlvdNctqoQGcR65qTcJ0nKDAG8UOSGmxETQ/c4xDFoG9rlCl8pTy9QPXdrLTEEOtiotSq
B4StKzGJzdq2lDA9aPmhRvAbbIqtosZkIPnbmW0fCo1b0LY21iwN3/0Qt7pr/EzjyCnfoZxcXBXi
RzJjkMcKlGJiFnVey1hYmInq2EnTZcNH1PDQ40rryM1yy5mUfVcQULi7nyuFmqFdGS8LRLB+i7di
e+HEA/f48IJ3z48MpXaglOIT/E5XUw/VsDJ5MtY1GlXj9PjAX6QrDoCrxhCQ9tbfyUatFe8Y0ZES
3lTSMHdiATFTS9R74IRx8fFeMRPHb2STmq0eTICZtnli78T12JRsSvHkh3mus+D5i8+wSfW5K66s
S2beKtEH6WYwdhT2eqQaQqCmLrDMipv8bpHt9b+Y9xgusDkaRsotvPFnG+cIBv33Zr1jfhNtGr6D
LV0HSmqCfNEpqCPh8yq58UY4cYh0Uwo9eKdl7BYBztXfA9yWHZMz+HTjbElbYMEFzSFj/7gxCaZa
li/y93P7xRUjbZhrNIukuNXj+sxSuCe351CKprLf2xbUv8e79qN+ChmzodQzcnH8oRv1CrKrOSw2
66Jn527W28LxjZ6ppyqRWQ4hKZMppC07Y5sgseCerM0kKHEodwinrhUuYA022fZNpl+crOxzTCKx
V3ypdnJrMOJXrDyde6YGjoFYroGMC7aEMcLYRYvTuKctMJJGlQHhBS0Y7Kf+2LT+EZBENleKZkXK
cFtRpz6RE63noaoFuYcHGMNKn/+ZWpdiGSLj8TfnqBIsP/Tqn/D/CSIs1uLvCUVkIs8kqN1GmPC/
zYCrXnEgH8n5NQS5BMyEKXCtbPdN4dvCNlWNxfqiemgiwQT9OMnceK7Q/haLNI/RMCe51zQaFur1
mrTIAi0Vku/qp0tGgawXRKZx8D9p1kvOoi2fCd2xEobDfCOIpBqYhSQn9wCIrx+8C8i6iEJzwTAH
O7N5u8VElk0PZDXosw3ZFQ888Hynz71Q0KIP3RBb1LsuCblzRXMqmJFUu/pmUyeNuOLMwLfxszwn
+KHUuIOCM0e6+iAskHTHxgBXFNR01LwKjlCQ/BQeIlQWQuWAk0RjLRrqhvpj5R4TRdUsEbM5Vuds
eQEClBlwUvl7UNrDiTe9q/USdKh4q8FDl9OWJhpTF2T17/HkvJXDmcEHn2kho6YNSDGE9DBK6yEa
eOWJnCfm6wfq2UuQCmJFxOjAw9BlmgMhGwpLJBugrrYM1/ZYqU6xKnuDr/tyijZa86qkTpWbaDjo
k+WNzIA4hlrUkxzXATijAfT+oMlNOk5g3W575OnqiM4huShhVgb6QdI8Pi9AZRAKYfpvwBSrfuj3
rvhrGEUys/zhsLT+dwvl+L5Zvs8AtVYx2j7vr02twyYqQLYKWLD5Lx2kZix+xpcVh0wunFW4YTqc
S3vMOsePUupbLnruRR4TrGPyX4jTbuAUNqnrm501f/0obrw1rdTYYJHVdvcJaNzXS4Qov9UwmGYz
9ZoKV6rdp1U6PdLoqS/AFe1O9Q1T915Gyvt+KPvtcRjNpDFJzs5kCV5MyvgDa7MxI6LtI3JLTOtR
xdKZ0siRH2ADDq+XcX2y5S3SKk9esZVuhzGNXOZ933whUJxH7y3fvbsvMjV93qi99MvUmftXxsp5
dunFr7H3ncS9cSwws/J2zLnCt2qBTaC0RgS8L2bPIZlFTHcbJtA3gi1fn7byWbHdfr74rCC9rA0C
H+QUoZ74M+Ml5OTsqsP+JhUMyIrQsuD1Cb2KqhX8J8xePIvs1iJo7MPLr9sfbwGcs1FGPqPbBZRH
0vWqBZpE3LVZGrfzIUosUK06t2v/y78wofW4BhCc2O2IFF9UCTCtkqLI4VdIa9nmqht7/hgKCba5
o9gL8AUES2xYR01X3qnOwcWOMlNXifKva/g1Vzmob5OvomkG++z5UgnVJrunixGT/U5GsZ2ccXcM
hiH6cenKM9f2XZCriEF+Kh/xRNChwrbklmiBMVrg4xF1MkLLlOgtdxRKJVhiKG2gKv7ri/xT1LkY
/Lh5X3iCKlk1qz9FbGv8WQ5v7jx3AoRGiowxZ1g4fO9LTk8P0REHbJWdt+CCH9iwwEkgN0fQipkg
4KIi3xydkTCodYVFsc9aUtrRg5rDJt0DtYsy7etWd3ksz3fH6F+as4kazfqQCDTCfnGzwIqlVqmn
Q5kqMRT7ZY0VRdx5Og9xwAECSCQ01ndCGsqShqo/1o76fF7w8EsoTKtaWFzIepbVLuuE2FwDAlvv
1A2LFD6xVUoRfrF+mlTWdwpbRvvmNM+43DusbqnrzugqvpsX/lIJdQKmP7eTP8FegiF83+1bI3s6
Km4YPTd9/8JRWxu0BXPyOfFcCdM7On0xTNYi3k1B8hOcR2ju/dcUR5g68ZBUMEcqnqad6/dGccfN
yPJJ6L4X+FsWCs7numhaWH9pQbCZpzEIFNtMnXY0qZmUBuAuz6qV909CRmCB+KH1WMJDs+4wclZY
2n2W9Z7pkBBBtQZEZvgbAIxt6zi5T7W5beSfjjCL0dTqdnNS6fdvGEz1Aa2QOEv+/6AXwOR7FUhQ
sr8eFsrcF26B8y92MxFB7KKoMDpBdwKn+pMDPMacrdfSpL8WxHOItkATgjdqtu4YlvDb6XPCKHHn
Uy0on4o1BN+YfY5VAREWuHBUNWutGYGPVbLRZEUGbZl3PAh7ZxEz+COjWTlmRsuv2U0Cb6MXohJy
hD4S5mBiY7gxC/U4vYGrm2la2EOyfXu/b+RblnV9mhK+THUDc49JEJ5heQqyvPT7dR5v8EPM8/+x
yby0dhLFNKqrGKL26LHv9z6HNKb75LhJwUKFUBVRhtGQ0xiQCwQqbXSTjB/v5IKtcU/16YUMg2DL
Bc899c2SFl92WhEREuLgqp+2HkjwR8paNtGynjRwGEDDQb1yQ80uK/9zkmvsWrEmuPDiXJ85P+iy
4w0Jk2XiNy+lERrlt7J7Bd/ZZqNmk5bBMM5SdZS9SW8Lb/HDLyurlMrsj01UrJM55reT0maOKWl1
qZ9FKBg4EBtUIigaUi5Vy8UMBbvM+1iao/EEHUApIazOUENJsBHJNCAMJVi9VVJQZXo4jEfSwnVF
3qmuyPc9EPWvCzQNUk9oucAWWibAMgcqfsm0EtuzgBFEyUJyns80xLSnIYECFW5u5mFUOYnMw8k9
HvGizJVDtj10c0MucEa+pC5QSxvkyBPeAsmzLRmAefkfOECqgBSK2cvXnjd3kJPQ3tF/yiM44kCT
bqj4ZToMnQ2ylP20xFcfjoakvv53kTi4+Jo1RvsJVUwu10Xxu1WCqFxslFw4WvkGcsvTH1SN9zi4
gFdGJ+pKXfqdJjUvWs/WKeHU4ncfvYOE6M5/ylZOmMGLptAesCQB+UOkc89NdshLzVtQhwtQKIgd
9qY01H2tU7XJqAkkefJ9RvXUGqWzRl3sqCP/UqMxqs6MPnSnordJb5DM0pf041aXrseJjFaDFFlX
/UkAQyVkDQLPUASREcPyWwFyV5CkAbbTXYI7ZKqma1JeMVxtvrekaEGglT5p3ryOa9ZYAUOvN8YB
E09gGkKD50XWbtVOedkbcKhBzHf/i0PILdPT+VEhksJ6AixLn4VwCHo1hm28C0LWriHHsCj2bL0E
s1x4wZpzIy0T/htslRVKrY/uD8QRxReiQuKywr+mcqO/lwU813ZhVoFi/cZJIj481bsaMCaIK9Gk
X8VB9KWJCXZpgMXkoraS5//4cTAxU8MjAE3R8w9Y8yDLK4znEyU4d6XNYIhnxPrmZ0V5rlbbvDWe
QNusb3On9dbZsw1cxltipRd/NdMO9UNkF1Z3bTrqKRccw+aPKc/4aefaPPIdf5wTND252+U6TvgB
WO8sJeHMm6NLOaEs21p/li75EspBYhLXw7mzwXIjtKOvwhAfv2wmssACKMJhnSr9VtQB90Gs+61W
9S6A18c1/WQVe3Kj6KLnhYGppdMfMlwwfxWkFC+VBdOkGOLUg3Gq9Obv+nRTZxh7TXsBp08qrywz
2wx6ulI+i/smElpPLCXD1XFYnIK045yQT3rKamuNNnJmZxxkzSeaOTgMvNbx8IDEJBQDCsyHTH/7
+PAuaoE4QXQ+85SW06lDZSgm6Ry7FI3DX/Lqrm3l1ZVO9zfoFrw0X0XWHkpbJdelJLufAR5xSA9c
b8b+CSUoTNH5KYOA8cNvl4qCvwgMfGrvBD1VBbw1A4NRw/75yZ9hKobVSWoqjmGKcb4dulSzDr+J
cASZg/Na4/h/aUQKKlpviE3i2+ipaS72fU9q70rL17sW5QYRgTqcxgh5WsUWik5yS+LOQU+9L3+v
r3NBdJyNyFge54E08X6U3fMNspwNsKOX+FHUc1mmgldjxx9Cms2frmvUaeKTndFemJFmlilqjUsW
sOfHdsSs1c2a7MBperjnywc1KBCKbWXH79qo4OKqQbOrvIXOVYp19LXBhN5HTEFHDdLEw8lXXY1F
gqIoIgEMox8VC+CsJdElWAs+yAKz/iWuOlDVk7bJZ7f+Exvp4ycny8Ng2+ZDR5iKG6+NbRUuidNN
sQb9PWS3kTn0gCJDMeDQjyayIp8U0/gxjlro1iGVY5MjoMDUDo/KTnVFkJDmV74AtvF0MPKygiaP
dG42X4VZKdsOZLtse5SAaSgExEccfWOUMnLedPQavMmo1Vg5Hl1U7uzab2tAC2E0b7kSm0OiBXpY
a0DjrEoYU/Wno+zt6Zb9VfCoZjyWjpiaOlvDI2j/VizDkcdxUvzcFAWOpL3X00bchfeIs78W+JG9
qXVVAwclTdvTEe8w++cV03jYzMQOnWoqA8Jb+97nmguMVOG9ZarEuA3ZGYUHUy/RHOYNDEZloSNn
M40xmBrbAUhyHvV4nL5kMEEhtUVxslxDD1upRFOnZHG6336O9LZRa2ToXwDAWH9wyLMFlpAcODY/
XwsNzudXU4NQf1SdH54U3bJGwJ2CVAMXkbwdibxOD7/wSCKTGAMIoEiW/yV/cKD4fOXk3RXyI1uu
PE5C6Az6JVWsclnHYjrnOjz9SnmXkeHW08EeNRH4Jb0VCt45x4aWHVByqLh0jYrdJcTP6kCMZ9ea
rmAQ7X+NPPPtc/z8pWmX62V/qnx4LHvOojdZSnR9ofPydHMrQO3RlEyInX6SEzne6RvCZPE9T3TJ
TaE80snYpEzzwkZbC7JQBG/GYAjH2PkqWur8jRrU9luo0WrxaC+uF5lKEVZAi6Pl8Xz4risD3u3E
g4nO4dBtlkhdA08B7gPHqWprkpHEerIo6zYCFXhl0HkdZ65i2ud1fVXOrZgl5Q46ZDV4BI9tN9Kp
Y8T5Q8O6K4gScVVsw+UNzr+ZyC0SjRHAPAfmrUaSUK6cwmu2LBGtx8tmWV1WHYasaJpWphrbVW16
PSlpAKgE/qpDheW1672gHmp93HymzZ/tnplVnilSGp22q8YPlIzUo8raCpXCrjNNfjWzsINxZsay
H3DnrHHObA5pwl1cazuhqtnThxKhzn2L2pnans70bvISPJXw7FPgRVS+FQZhH3sSi1IfA2dK6MCY
EwsXKMtGMmSLorfJOOyG0Q1aIHynyZPcpLsPNbZvfWIaqxT4XDdKlUp7Gl6Dt4EYNqaMcNs6tBSK
OxFmJ8MyYkhf5tVeRdEjynrCBVvRAHX9jY617UepnWCGcaT3LlCto2/3LCdXCpEX7AEjn6AQsNpN
BZ0r4UpKKVCyi6pD5MMCMWJBn4eNjX+G8jaPA+YJGDkyacYQu30uDgXuRQ8YNg7TaLpnCviPR3bR
sYufYmcVN+mjnLmzl3+AuNANRW3/7JKXVIe3IZGDPzO4r+AZ6DbGR2F8S9cxr4OPIz/qEMRb3t4y
yxU121ZU2xFpeb0pmaMHx4cjqfxBM9BrBL6jKLPhLWBQ5flwDxKZW2xySuIYW6aJxysYcD6wauOz
HckOGRwkhGbFKq/M0axPUanFkkI7k64cdl5ypiTJQHuGmbR/7umMzPF6CL9ZaTn13vpypLWU6j5G
CZSosT8jQyRSbLpLiiXEf5wkrHUsXxWWy7UJBCX5IMmkNS4kdmfjJH3n84F9uTURZBykP5m7Kb1e
4ErlWhBzXKlrTh09gHPD+jWq+zKZS66lpzlQ9VsBF3BaVFfZAr6zd0gdG3oBjoNaR0R4/bnAU6Bx
c1jYryqrQzCMzYWO7n6Vf70t1jArMftf+iGYVEmpTPaqP1wLUhmWM/ci9rv2hC+hXr8psnw0xqWK
yo8OvYYAqtcleFhhUtzuOj1G2bu3FbfAMhXzMaognAa8/HMjNDGuHn8h7Ecp3jvLsi9EKHbFOkNR
4UqdPFj6lv4B+z4uKLF9AlJma5OipLg14Er4A+CYtqGDm9rgFxzi1bjIcqNUvUtHpdSB/1eOyMtF
rxuIMQpdK0OW1b6zS7CgtntwfzGDvaxQeo6Dn5WphPgQaqrXw4La0IiWHc4NushiVAASr1WAu3pY
YlQ/p8x8tczcvAU64FuIp05jTSfpfaQwDWrVX0qBe8aBK4smIuskr1nMYjTdJLEo6f1Yb30a3PKc
AS8+6r5t+Hs11rh1HOpMNs6w2yhVPMA9K7yrNqDTnVNqxWjx7K+BI3CcMvZ7aj7wqGreL5MlMfv8
kgysWaSspMSFGYVyfjnrpwnfnOJ4d1b9US35SA9tXoZENRb2Lr6xeXmBqxjgdevEf3rlg2+5rciq
0a9mWoSRRF/zeCeqQ8Qhy4WvSPsfp0mD/aRAfZO7CfoOF+Qngg5tJ2y5/iSwPchdrtW2Gmyv4GcA
l+yRoJm4ITKZkS8ZJaWuS/fAJjTTMPpFkq3a6lZNH2k08GIwYuWYMIK7BVEcGlOJoJmKPjqKErO9
vGbWb273j0+WkInx1VJrPtyZHo3AJR2Gh6mm0hveGO6h+kD3tN3AAkpF+KbaCghEh3J+KTaDf7UV
qUJe6ynqPPhcWAgVPoRhvPJCu24oDXE/qW4iWRyNpUY7NWxM4Zz3avFAqIZhTdAuVbG5+tAxHmOs
KhIGfbkSAgE5a5GTOO1LcsNLe9U+EgVsXDfwi9cBXxq0mozSphSrfS2cvApi5BLLow6gDTPArdiP
sh4r2uijV046X4X0wFou3BQpMD/m21oMLxA0FnriYeQ0Gr98IwZxhrXKf474pqCgmhL7K7fmFufT
m9Hy166fgp4788MDsGZLqyDMTn1fTfnE2+7AA4UT768M4xr5fjUCqJyG3rfwV2np7jzwkzg3LR8c
jzWf0NwUcNw0FdhFIbftyZk8RTUGegizkfSXddBfJCD7W1jOhIqs4D7rgd8Ahv5uLJ+OOw9cNnWW
qhRXcfErpEXCVOiBKe+V56t6YVD26Fqazj9MXKD/8nvjc4lBePBZlKxVVgnudaisFs0rZ/Vwhj6t
N54UgjDZwULU92vzvqqzICmBlFCfhhYdbkDlG0nsTaUsavndNyWwVaSAAVsMP65L9iH2Ut+MHCMA
JwSxA1wr9aNywmFhoGzqhV0+s3kvVtMjauNvAx57P8veT06iqZFHob58aBfWcL6v6iPPVDIRrSX3
9oMpocyj9VKlR6oD6fjDOcDB+kSnghdQ0enUp6EstBtKa3igX6c9Hab+2vPBy41BH3kweRTUXfJz
jO2eQA01V9xNfaxCSayZO0N750TAL1X3S5V4+J9GbhkcdAthBt8hvKVfaIaoJTTNlthVOJuhzt2o
7ZBMF/iwyPRpgsusDrWblrU/eqgfdkYuEzDwzzJFzuQuXWkXUH+/dGai4hyB7YF1NOfoT6B5fbEV
2Kcuy18ls7cwWOVyNcGanF0dhWNFUhFUW+mDX5iYxhgJcg+kkDCfgvTA0e2qEUC4ig7yGL0fqyCr
FsYZzrB/BAKVkvNzx2i2LOrfqbyXiapCJR27iLxEjtZlcUWdQDrit7N41fXriJsWPebaDLrDFQ0n
yha2jXvys4eO98NXNiqcKTWznNeAR+lF9I0Ik8HmOCiRntsvijrAhnIPBjLesMoeH5csr0mlA0CI
7QA85tuD4hPoR+bbRCaFLSw5piKNd+VPe/mkZ7tConFo27095xPz5dHycR0uOW5UJOOnipSRuidB
uZ9KjV434K9D+9mt8bwowJ715oUEnwA0oS/DTfC5lAZMJnLch9Uk+9AWknCi1Pa91Hncw5aLgY22
VDEFBLVxE3h0aBHVaWBICE47yQixI6X9yHpCqWj0p46Nq18tz7h6APX/t33RfYHZ8lZTzdGsqygI
GhN4Ic6Oa3KiIVeWwqsEZWpzerK8997VTHvDZWKjrF4Sg+97FRlpuyhCBQrfis8Du+Z1hO17x4Gy
qe09toTbvx5xwUby2TpftflQ99KOv4GpYHXQXc5AyonLmIdAf33M0glXdya9K2auApFif0qyYFYE
i68ztWPeI7EEyK2SYwpTj8YFugRoCHC9hujqEiUykFELNnenGIwsP5AuAHWlZEcLZnmeJxqd0gLt
MUepojY5uTokxvVToqHU61i2Gw0eMfggvSXx4MrjGTDDb2Ned0maA5QrZKbtb5EB+U27I0WkY34V
hInQPv3bsp36Mf0drIJAfepNTDiU5MELNsn8a3O67O1UmWVeYQVP2x81sSLmlvS+Mu7qYdvbYOlj
3eNDT1EBlbxsLYJNl/nZRaeeMQ4NjUngO3TIWk44bJz30Vj2WT9TY3OxdNfA3xVsqOwvTBI1OZrH
57vdiViGj8WTW8y+iDLnxEmTcKXeHYX6uEC8R6izyuNRVIaV2kkFYIrbQNzn/dJFWjXYIUDleOw3
slJId75uaaCOncmwx7bSj826NDvFuVZZEEDCU0wzGaZccpzvxECKpixROvbDR4fUQLI+G6nMHJ3e
EuA8+H6eZhtUNeFr+FSTCaHtTPyiPD1LmSG6AGooiaFWNfKnNGLRCCEWHWuZ8yqE8t2brYSRPD/x
Ro2bXBikYr/KB9dPjhYjjVTll+2ibYpjRFGNmvgqrXp/xX5S7QZlYtjTtymnNqxMO2r614L4lTgF
Nzoq41Q5yIeGsshVReU10oK33uqRWaSAjcYoane9Dh5Qmzrg5yip67GaEgSwqZgAdu4OBca244Q/
5GJAc2dIM3WRaPJ4mujj2egOZ/wA1Aqw/P+NwtibRFZlx7cC9jU31AfRQLzqjqumuV9c/PhELP80
RCGAYONQVgfHewKm6XephA5Dy1iSV0LwsD7oe2Y0r9OFCO3xuOTFlv/EE6q0HMompYte9+KLh00X
4SJ90OgwUADjB9/cpDUKZGr39QHxFqn/Sg3DTzfTDvrge06vvUXrJgCpV0ZAUypesQsFkMRp6T13
g5pwtRl/6WDq2auSCW44bQ//TR+FYDp3W56zkb6VrPHY8RLnPsodLpsGAnhwWgkfRDD0gMD5epCD
ClCYt7VhU0eo6avPH3OxTLsplR/kRVH3/+PDgag5enn+c4oAzaZqPb04pskF7qMoVDRgaDw4P7Wp
FMBun76mqgfF/oj0IoP+ikGdg2ySsysAdKuZTuRQ8UD/LXe1Wid4sr72+SJGRMd2a/lyqWoNPRUy
l3quOkV1Jj5RNJQg3th7YaZiNAill7bfjXWdJ6+QmwlppVGwc3kJHdy8LA1lAGvYDEFa/dNU/mMr
ocIDwFJnFkWssJQ7weiQl27dbV5DAMaGv6fkwHyw/Lu2KapOx7153y6ICpup+lGEJrBYV8qJFYU4
77SFehw9LrfRY1g74pAAmFyR0yXryZPUuWF2ayqW/souSKJLpPsH7npiUFltg3xSHxj9nAg7CSj2
dJ6G/IxqRwVrQUQKny6yfRkP0Fv+j+eQYP+hMFflXd00IWf49SISt7b+Ey8lmTvl49rOzIVU59SR
OUP5tBSy3wnRdQ+b+JJpBoJ3O7SpWvi2QfoOYCXPlzPK+Am3PLzK2hy818awFpjfqqJV0KbOVNLV
139OJub/xMGkOzOc3zItKX/ERwCyEoRa1aOyD1JKQmoRkCB2aMcTZj3d9Zz8alDy7avdEDZJKR8E
uHhpwgt/W4yAiV6JULj23vCRQ8O1I/LW2avPQIFpFRwnOunL0wDYIfSl4QSnBxi8yK/f4v/NEO0f
pvyYcpRrhxgEUgO8EXoR7u18vpak05hrcPTljaM3f3DLfYza+0QxJsNvdRMqaAt5ahWU9cGRv0VD
XHI+qPNuFQv01gMIRUTZ8UyPjTCFpE2FbKtpGkzu6my3X1WzFuTAyF+VQZROKfI2hb7l+bTHL/av
7+DPJw4egUlO1O+CtdWt86Vs7cEuiwvuOzLq+/QW05ZZnSryM1jxme/6NPBUnjvVCZkLoIr5mrkl
iidKxmxFxbSRK7j7YQZtbgMjUJDcrBjAs7j7AMq9uHVeK6L2aMzXbRjOZQBbxYtgYnKXRXaiBLtD
weYfUZxNmqwNLNt70nOhtiaBNhD8T0jAAkQ3A8OLT4tNv7AmSFoZKXp0N7J+3zJ/XZaURyjiEiu6
lUD4gF5NSh/983JdIaNKUEJm2JHd3Etry9NOiLuuMY41V4AOZ5Yly3AJzPvTkMkfAgwVEr6VNxbo
OVbipM4Sd2yPfL3jNUsL4fJYDPrejT/ICKV6h/5sve01oA9vCssCguWIANaud5q2VmQ6C/gG+md4
oNkZTdJrqCZnFif+6do7Jx/EFhagiycDwbVoruR5qv17yb0+Mw5BdMh38jpfpZWuGktiXJfAcJtQ
zPE7zobQznG0RglJCyTQBZlf+YwD2yjM7pz5Q35p6Rk22iI8eRzaXZ9L1oIBz/YGPktKzfMohKfI
O2u1qPYhs55B333l4jtjAoTP5QBdqKupB6a4ShAk5LMqk+9dZmP23vsgwsBDAOrny/TiCI2yIrp+
mHdPpacHEXezfnaIEKYCPI4ZtpTq28/3DrQCA3/ypoIVs8ehqJBlaOqia//fNvpNB89hHj+XjKgm
WVHkeVx1T41dciO0cg5nxkONbShPiu8YjAyc/jyxZPS7sVOKJTF9EErE+ixPuI06ma9ES8/plVSm
ZgERQ4tAcvIfzfKO6+jxPEzkDh7SU6YtJdEq43YPGdVfUEJ4xVhlrV9cFqpnmyQWdRXmIOUo6jag
vfB5z5XDhQI5cqpDGYahi0jZCdnOljX03zsjXk4IgD2OBC94zD74NaORplIvlckkZzkAJHXC8X5t
YlTK3qECWPbifJj5tVEax2L/e5yznFkQ1GZ4bJy1CTnYg/NH7UGvgc5EeemY8ZTiqCZ2E+V8QbLe
ic+PmMjeSaYY5EFt6aFf5RS+XMvZnIaEZnFxszAteB71P0ew1Wv9k9SP13mjWuazMX9zRfn1QQx7
2OSToBawH2uOzV3YIJ+NkzCZ1F8vU4gXpdGhu1Y8mvvDZRS5XeYQQJsa71nDTAjXlC6DRyPA4hCp
q5XTDZ708wIcjPo1S7FlQ8xi3A2md6QdDPfrCZEgxJLv4QwcghbDlxrNn+WRA7VbCNhlJNg4OKxp
0DwYg67+Mb1j3AjBM6gi8V90sqDF41Xn6TBbpgER+05rjm1Ljkuuckdnca1U8w7gMvvk6ASM92qR
GQlKZeDEUwgDFH+Loic8CqZGW/4CHKU0arS6ASY7/WbJEbb8X9ldDbr7k1pBzX24xlIkTyz32nag
FZTQ0rpdCiS1ePtYwe8Si5moV5Sj0WuDy1ltpXOluDiKqNalQCVd567+dHRomS2Cm77cJQZ4bEx3
ajjiVRbf2iep3UTQ8ib66moW2yck4GufvWiZJpdODJ22Pa/EC1vw54ykOpyjwe55JgOw6q2VU4fH
WwaJf+aghwETjX4Q6qSEIrKgSg2V44+HbkmFtfFPYF7ZQzXLKcq2srpPdt85HclM51k94bXbK/o2
oVwRlWym8HtkQKraHhgFrsP69Wl3aCqR1kTWeTiGgExRYTqKryFTFe0aRhewy4nvnEHYnLAp/2cf
LpnHkKUzAMOBNi2oGTEWw3i95W+A1Vm7ccjxFsbw7+up/wlw/ZwKT1/l/SknSlbxy+RFqMLfGsz7
o4Fg4BN40pCMofiySjDh60OB44/NgLsaGm5alzVj9Y+wXHJOrBJNI98JHLQPMh4sPMJ0OMmaxGqf
TqMSZG06bawCBNNDEhV/Q7dwPHGQ0AhB+yUxM5+W70may1vtF2Zrp8jLb1k9d0VYNl181zi55JZD
wKFf/cUaxPXgEZCPgy9ONamxKjzVBMnss0vWUpFfWBrq11MQLpvCvHY+bbNf91FRvgrtYSCH+Wmp
isGHTBDm1+y9cUjShu3Hye4n7PU9MCfoqqYLe/sPtNCLCDPUXyxHAnV6P3xVAe1I09HaciKkS3qj
Fk+qdz072/9tM6i84K3DbuoimiIWn8G6/vIHPamQT5Qxzfj+tpha/l+Blb9qH/qhPIG+LnvTuPtF
LF+C6/1fmArClYbQ5pvL2ZmNgz9qrQsu7kK/LZYsKpMWaW6FJc7o3zHa33sRSHcpVdh95qbiZGns
+IvvaJbU3TkFfElWtP7wXqgGE1I89jERoPJzcSNf94Z5T4LSHxR8SLw96xcmbdsFbO1hW6z/Uhlx
z8GZ+IaTi0B2JWeQU1iRJM7aRqXySxCq9loUWirW0iXoHGA3+I8P7FuQ76qOfdQRDwyTaSZw+tGD
34Rr9W8T7oW2D/bqHYbc7gZTUba/Sow3zNDSPSBLkqDUTxsm+T30Q6RBBng1DSXNd4rs5a5VjWtR
MoKOD0mxL9ylhDWMkgHYQszi1+ML+w8vNfO5S8ZcqBnGtGcFwC+FY9CVh71UPyoMEiXjiUnT0rsG
9aUFi2uydd9vaWpyTy+Ec/o2fsAEEJGQrKPZeuDQe+cyjHjlpEfXmkPohhtdLdMWwGvG5pWd8xbn
dfqdoKKIihX0LfXWjrqATJ8GAj0wUe9Wfus5AOj+7Au0t5O2l9uVpiGOCOMWUD3il71aD3K+AjPx
6E3niOR7RGOT0wNh/DZKZvNnPQfpfXdrIJnGSkIz18xpqDapqU5gaL8DAhKay0gd3BWUFEm0sQlB
aM9XwKvWgc++XHbs/OleWj7BTmPlza6LRVNwUtOOBhvS+gsx9Ia1e6gDef7LWqdUYPqywvH0+QrX
7GZHNUSmhmDriBdOoI3hQeU1uDMNc8ysw1awdubLOV+id69oVxFa7d5rFMkRbeyNQCRPTq2Ksl+K
T4snDpsd92zuw0iu0Lza49OQmA1UjgaPYpMGi/sSC/8ugW2+J6ieEmSC4FJuWIZOlMB0cJrEHrf6
y/UAgth5lIJzhhCgw3FwKw8XMN8foPJJz0qGeouX06s5GNO6l4b6fizzl7f7gkOZsFnQeaSVUfGd
fDnLb/0V5f2BNTyvKzl18S7aMiv5r+kSPXGDi/WVAf2846RSGiaWWvu1me+3kQcREYivfO+mb2CA
YdqNVIdd0pmM1Jqwto3IdZah2FSWhojg4pz9Db1UP/A8gVAs++sr0OqZPsdV4yhf6niHsCQbpRa9
PDyPsZBrOlSkYp3p3V3QoBmq5/HQ4NhUmktuZpyypRcghQ4hcgxp7yx1QW+Af407PnG7JpN8TuRH
OVi+txcapi3QP3WxB7d43Q8Ihc9GJrbJUVwXdt+s6SKX5ndUtHUOR54/vK9G/rlOL0iNJ3dkrdpk
8DOjJQOiymofrbzhjKiTe+cLMW8o8pL+xg+P7RWaIdqbmWtBT/fXQJ3Tc8/7TmdX5oQUmwEqDzDn
G2K/CvL29fXuGNGB/8nC2KYuxFC3ENEjKHJMKaMwkFe/nmKlWZzPlULicptX5yogwNGBGSon4tzx
Cib7htzP9AtQliti1YfmRBEPyHHplyLCZ5bRGEh4P243Hm6POgtxzUVSEekAqWEixt0KArZwlUFW
vivSdbpKd6OaHlmBMR7PoeZBU60UHIifjcttl33pBOdGa9ydKuRpY6VNrAwOCRUKJ0Wq0oElDm4U
whvc44ioYcV3MoTMnwmkkumMIsvFE2xd0GQnw7GhN71FkAmnDNpxNcY3b31PHsa2/78B1xF0J8nF
j+7vYU+90bXnDnDOguKjQGF5THO4w4WMyFwgg6jVbPZQm3kaWcGng51hkQbzShnHuqtyhnI2kPFI
OlCSGXaWWSbyZ6kh0hsXrgY/woRLWlxoDvvUy7V2ahkM5r1tO5HE0z/mAlU9bF4L2fYpv8gFn5/D
jJ69I62r1J4Z7Gld5bKdKGIzCJTZwwL2FFOOfakY8JWplWK0vKh6m/zIkqrN4Dgw+2QYSkrsY/E+
ytmd47EmAlS9/eZfmNJak9z0v1E53gmAwFpWdi9N05I/bgH0Myg0D9yvxk6MA3O+dCqmxDPzdjSP
R+R5jT3zfiljLvbHinF1+QLDTIJfPhpredTkKV7ctDkEqxDj7dlOgVcW7BzmNrkxbWrqiTqLHDmi
b6F+P7iudYNuJbEdsiJ/MwmFA11NFt+7tnaM3mXzDAM9/1QnAkZZLvtNEwbZQupaXbTYhOo7TDq9
y0QKtc4FOyy5mwy8Dx2srpgfy1TtkR9/wN5OIZE95GSDWCCi+uZZupwQuF0pxncqCer3jxIMYRVI
xGGqx+/7DhAnTpaxx04gdk9gX0g54YJsTuWcnf+NM1I90/jDz2iJJKn/aT7EnWnowOQkO6afiaFa
6oIIv2NXZruev6R4kb2EnWopx/t10V7+2LiN7GT0YtKj47eZOfE0C0qAgyJIVbgo2M5p19SPWNCh
XnM+C3N50/4atY/GdNvqHiLiGAI20wxcJPeXUBiCt8WtM18DAgrw0k+Hgx/L1URwKcUmNIQ7iGo6
K23GPcT+NwYkGVY3poJXKj9zV+6W/+LIvDgtyiXkUR04NZQgb5YDcCOsXbhLe1XyNEOTzJl/LTGG
QXZj1NfpmVyfWdQ7p77sIGJYhjRZbsc4XHrAfXssi4yD1GRIdG2+0k1agspqkRS1zD3eF/p5Dp7B
yR+TRasuYxFF8RpSzlhab90cR0NljISAdKX6e0VFFHdidfWLC4hmfGy+fBcApVs8VFpLf0IggAik
U0dj7rtxg7zaAuH46VMHexdxMKEMnIaR2yZVyM3sCgnY6i5v+CUVJq45rrsKAUKWdZiZAhHNoKB5
x9RtQ5OYyeinjaKZY5ZIzKNMK9CCbnt1ZixY5o4v0ouoFxPI5q8sMP3cEuBk9I9xI+mgj8PisDk8
pj32OoIvtID0A/nGRG3Q/GHCAH4FQ/VA0hdRQCbBAdlueweLbh9UKsC/AnG5b83ZmNRJbLn+59pq
LeX6O3ds5uSGOXvSV0WHZu75nR1yZwktvvazsC7/eCnYs9hQRCYGQT0HhqZKTcUCgWR1ArvUm8vs
HVsPVMo2krqkeMx+4oxdXNM1DYnPLCE9QYfO2aH+mrXZd9CY5M1m8/pVKKZc9nuRcxLvwcbzDnv5
Xao7wbEu4umpOPwdEUjiENJWY4bnPdkW+2JJA3nyC6po+rP9iG4zutYEPNtC4Bo8PJHHdZ0XHQDV
2PuWR2x4qkLrzF8GX56Vb404hnohj+O5biLmcKljamBE2nmwEMxjssyLcL+zAnrDZjzlzSEaPncN
SGYilGXCl+Wzykdcl0WWMLHF/hmcpqfgPr3m4dDfQJnGPu9PnfxdWWb5OjiJ2a7NQpjRQWQ5Kwh5
2N1u7sit35HixIZMKbci8CiEpMRyvSzs1DXY75VoOgGoUyOCsWy9ofYIMyC0PMbXyuFXc7DxzJ0D
K3Y6WKHbbPW3hY1TkR7t8+afzrASMwCeCj+RdnIPNIm3fyjmB4B4Qr7AiWwzbVbIPz0hHgs8cNE3
HGIuP0ZeNIbPQ6uvv+dFWXtAIqLEpqY3D8A7bC6eKEjyLULlpuvuls0kdgQZO8vPde1U3YTpUDGU
qoc+3QZP0bY//uoP2Zwt9KU0hWnAF5LAFfgdXrGsXANJ7PtjvtMxKa2AiHLKpOH+G6CxD4xMluwi
5N19FMxnhUpZwoFhdcVYEFH5OUd7w2kN15FS77Ei9ZuXhcKG+KljN5heG6s5HGe3IecFKRvFHRAS
Md1D73Axe11rXkRm1kmC7OhG4hnRgQ3IuUWHp+MwGZBI4TL4z23HRhEHU8WnCaXjsaxJhcKx+VGL
Qedwjv4qQ+8+QVE3qnzOM7S1QDW8RvDxcfC/i4bQHMvzGboaEszZ9/TMhCDN0sDwEcFvFouQK0Mu
Yo3+awGNEEgbAAtOek7wN4tp0c9rvKOL4bdF6HU6cw+G28kW7XDiqRjEFNEU0/jBFMI3k2hm8/sm
jAObc5/olLqin34Dxr6U9BtHjEyab1zSJWhVqI0sqHEnaHiKYmI7WwgGoIKWQgGJZUb7rZsGzcgY
ic7KzmyA+Zva6TTPzuozDGx9gN7Yx3X05WiMiBHGi+EQ9hBGw33aSa52FH+jF3rZWwuhhFIgImUf
sVRq4rH5VvIVqjEcgm+GqYB+sxyJ0pSyDwzxX0TcnsfZhrvsedQampyXml/N2P4tLYm3No/r+4F6
/C18tAuXr18XmQZiksSyFfoCO6vNEVIeH1dKkdnSiEkl5qSazjhybm+w3edTsOmqD2nhHDI11aSp
S23DR+pT05d0dZxKoXinobkLO6X7LxlF0SBGKvCtrhNOS4zd3X8+J8FyZKwElRxbRAdaYCsWE76j
lR8g42daiJK8WkT1ZCRM0EDZsX036VcNayruLKUhqRdhOtDZ7UEYfrErTGO5/2J52ZkHVEucMihl
Dk5MKQIpPnkgkkJB056+VvX3GM5mOm8TUN/qho0qXDVC9Mw1rlLVYNqg0emnQpyjfwYdOfGHA1wd
9LjcyiHkCjyDaBR1wZNc9QmPNOve16J7eXqUKoYmyXOEnelTtATVGQ7I+oJSrWVzxIffu4E99ghZ
tMEZjaFAdfVocRRLwIwqi7ow/Pz2UDD57vnoqB/NwbqQcAj33i/x4NsF904tWPox7zIFiR8RJFbw
by+EgMQDeirfhgiQasR8nr3+O2i/rksudhOhYgSyWgGNICt7rlSQeV/Gppyzc+j/6R0lTIBbJ+no
ZSNK2lhIlOdvxlNIGwxaO+MYMemBSQPqZXMfB302cijMUQaicVWFo+3A79nLUlvCRugYVZquE4XR
KY8XeK9R9V7o4KVptJX7ZpJ0xYtHGpmjnLHrEdvLFgkLizFfhKvreKr0pBWbskxpAJ+BwgrCMg3b
1vEqC5OKjmgLx8rJTTxHsXI2/4oy5anAaoQTUlfphbNQLr9VZMFfG3l4GPTbgwHKz0BvOqy/L3y6
/D23beZZ/Y+p0RqPNlqPl3lasd78f8Ur9L3hw5L2FlpRd0eoB3JbkvO+JSJTS26fEbz9D3uKe2R2
7/vIRMtUkqd0w2gH+LIu7JcWA2pDEflJdRInavQviR/vXCfmU0ETRsOQr/NfUGWwosZxkI7UmqpD
zO55rUYek5jWOxku1TMy7pO7Gh92dIDlGW0lD6O3IpUlmFq1/vYGlub2uWUFC30DKfxqB6e7mXc7
AKe+9z2vZxeXLflbxWQ+dUXG58goWkGCZZmKy6W9nwmpn7nM7vH+SvkBPxn1IvZMb3pn8Bj5RZT5
Ah9jG+K+S+5PVE1ICDix0Ynyte9CC5YYbw90jrDL6RzcBKGGoamjfv2JhyLN0fVjHBNuKbsgIMIC
Zg+VcTso9T43Ov3i44wUotVLEZ2AMgqfU/awEHnnqK/pG8lXdypw7iAXbpSebYdyzPRbvpZRWd8Y
8v8v0W6BwTTS/WPCJzbk8SH2UeGOcWyWAkiUQHEZXEjeAld9WyjoksytK+GDEsIMLTJErxScPsVn
jCMndyBCkMFPHKRuL4D/i2GGSqQj97S7W1ncXj34Tiu2h7GaDYs5wBxLFNSxyvpTj4ZEsyUBEimO
qCZiJREDfAD0LvjVoQInSx/VtSnG8PL8R09NaaZ3HqkNJVpkD4WrsoxZg6vs+RvWUXJC7E5EVlpX
pqB9qXf7muKY7/8e1Utc8tw1OumaZpUF9u+gGIBNYjonholK/AykeCca1umSXY+pcRIRlbiWjmb0
r4iZuyDdSEfrgSjuJqUyEnSje6nXEPf9FqzneNhHfgcMeXswzbvjq8N4EHCtbj80/7LIcu0DMAB8
HNn+PgfiTmebN3XMjgQ3UI/jaNzSn7Db7rUcOx8fh3SydN61yAgERQ5MeXDtjbPYp7WegnWBtnXc
eMvs/tLZLa//za3DWO00cR4OdzYKwQU1YawhayCP/JymSrbvKXPhxf2DVMizH67aVw9mju7QIVpA
+H+Ty6/rdOkCxsDD57b2hA2yqw7K4rR7ikWyhpZbEEGcyn4YFRHsvwINCfLHLAI+BsaNjja4u57c
saaSSMZ1lFvLmMqBg6M2nRi9pwIs9NeiZ0dtN5I56SYbFLF/TrUI8TYoklyqLnhR3Tt+Qypwfa5e
c5mr/5UGE40OjpVM9JLu5QBBx9UA2CXXm4BficYOAOZsIODBJJ6OPxdPu3WY3HxQYKEPjj61+5vl
X68kpq25WOWD5PfBSWyKGHhEW2FfSgdYdtjpWVb8UXfvTVrhE16SQfTpzz5d1gkqQ/FNFdZXTKf+
/ghaJoJlhtSmulvv5MMv0NzPYAMZbRRpKLYuRT7QWiK7iFQfrKR31DHLeJsQ21V/7AV4LzWBVpq7
/xYZNE3SFrRiJ7wBk7Es7Zaz7L1n+EREfnIWx3JVbTfIcbD/5E3jJWNcTL/wuAzgO9etqb5fDjck
ht3mo6ztvrQ4QGOVPaSGQTjjZYCtB4zOpY4S8f9+xsHIp0iTPxUKEk3VbPk2GS14jnf5oVDR9+kZ
/TptsV8KvRmsudlJgqMcCZGGo4qYTU+3QRbd6T3rmEgq2ABmJtNYKgWhMcRERE9ZXK7lHHKJM+hg
aq/tOECAzSTP6H4csNjBcrkJ4ZTSWQmaT+S6JU3BVBbCSOPjtCyKzzh03Mj3KP8YktIpPcDzXuYs
+QphyOJFyYZsvGo2wq/8KQ6v9bzzVO9CwC6NL/5RHOO+ap0zaXc0GgAEsIApSDnxvdCdJDZQlHz+
s2lKXiffzYLZbeEtomD/ZYA5RkZTJbiOamvzR5AbDlwQPM37eF+kKhcVpz1KpiE97PAUu8MwUt/S
GOr4mylij0LOPa9K5/6BnNnt+rucvEVLgOpFlCRp2lwoZm3Wnx7onQ/yhobQp60ukLvXp5SkHxg2
F5xtald/YNq3uIBg13Cc08L9qk0Q8PKerIYyojwNCkAA1/xTKEd8fTMrgfDwMKS71jcdcgsqApny
xvXlCbvlfI+m1tFfsxL/7ztHafUvqeFALA8CY/0PPWA8NEs/uuxEf3Rhw34SC2zt3kdOdzzXG/6T
gqBzT+gEgz0NYsGxMHtyLeHFz3bD5SjcpxnDHWzBA030u7uNBTils2tzsdaMJYbs1lJhI20hVTtt
BdEGAm8HT6qsF/820N46RYIW3muc779+oFvFjmSiadeHrccYg8wxTZ5ApgUbi2rYPWOJkjSvGcOw
ecDlDVFO50mWhZTC2zzMdjToqktlpgmzbqeEmdT6D0F+WDh4m6AtWp+KOuQGgJs3fMJnniA6Xs2c
eGCE8RIKKNOA3q88ELMlGEtfyZv7tfykGOUGn8Rg87D6mqju5MZ61g+0udD58HfAlniR3sXtccC3
VtQp9KXN/0z4L6WYiFaFmM405oZ0B80aIIKDXnqVi5eKW7ixh7d4JtqMIXYTHfENMlyZW7Wywxfw
Twp4w8YhxQkPlsdKEwVIa66LLpHxV06TU98gUHZNjKrQzH3pppD8FqbognO9HSfpNHALPUH6nIe+
SAM2ddsRaYENToYbU8Ooc9ab+Ho/9xiRJM6hSaIr1SWPqEML23/T1VF4ThAvaEKnOAOgoEbwTpAx
6ur2o54/PeFmBeBmqEZY/3fpvx+6gQe3ZJruTrTTSg4H6AvOnl1uZiz9/TaJjOcs6VlHL6SEvMeG
5IKJy5uhn6eegJ5JjVAJ4MJoUk80acITAKZhQ92kIx9s9whvdQVVW5Wj+ODOL+WSL9+K+3grgXJg
I+2cf6ybM8VcAh8eVWQjEMO5ym4o5xgqSVBDl6KcBuzLpYVaB2rSF4G+t0hXuEMwqPupsgsh4neJ
2YbqCeXrHckcM3Af0HUHoSAy+cCfG+VerTjN/oqX3JRXfS1r/ATHY/wx/O+cFZ53MpTqYsreRxZj
0acD9iLlhKJuls3K2q8lbUpl/o9iNqWjGgp7TSgYsBtGtqV6aM+xlUmilXy/XoIRwRWGTaqM3JZ6
2yyJ98hQJ2Kq6GKPPTv9ZhNbVxdBz0Nl+2cM2WDMdtVmpbSjIEfxx4nXK9dEfUPiB7822PRKfVGg
eUiFkyIaWfotWqCJSi4o+ga7WfqVZ4vftSASMQ8gj73+hnytFBCAGX+LYHxVNp8heaHL5f7+x/dH
qdsW2VzBUXV82ETasLoy3nQfBsgAumsqIFpoKSp6Hg5h2/yM/dT9YZthiD/T6ktm24DaIxVHaeyY
qwAiRa5EEmj7QfAZTV9KwAo/ZEHkqO43MG9FcAaFbHY70bFT4uOPUkf8m4WYi5s+xymfMtfZUNSo
D7zwzbcGXZOSzp/370OllxSK4bVR2qnFyyy4rR5AVP7F0VcBt9Dax8FiyVhxa4FThPC4pywYbAay
8cGT5Pgx+k9GHhY1KkIKvlxFjyZ4uqMqJmzqA0PN9IvMwaksKkUW6gUzykJzcndQ//iyqBbt4CDy
tb/IUtIBx6+GvnDOSrCQW0CdHDokVKTV69Bh0rh21OskIKjSHUG57UvfuX127/wcaQDPLzBHfFS4
Z7C4kqLsO0vSLeX/p0V2s8+72SvwQTckewGqoFOwLOpg8o0PDTDr9MYT0hXdBBxCAA9jzkg9pQWo
C+jyprQx2yrownA+J/t9BQVtvuMml1w41pHsiyEL310mTJtrTi7kEyU/auN2xcfZ+cgUV8QacwXo
H9YtHGqn2Wo2EftGvhrIBHj2WT6OjUn+hEpUzwJ6dnZYpbV7QzsOUPTBy2KeCOImqkOzFrqPbNyA
vWUNnb51TxOqmZrcAYMUnTABCgZeaOWZEhPlafPoRctZ3WpMpL+QBoI6PCqKX4F53/hN30DClBbI
qGMWmk1PLOYeoERjQk1dl2PtDEGO3LSj8RfPyXNuvvaLKJhCjQu7qRvArR5NxShbHQMfOO/lxUHj
CJqufjyTihaL1Cx1zB7avI/qZz9ghTbT6/1PqVKiYwH0hPapbtIUdItzCdYEAoQGpfixJw/3exB2
e/fu19C9GRTLSzbJDVhGBvFqTCx3VwG7V0uk/nHrRqr/Yox++PogEZacMUQsiv7uz5JTYQ4SznW3
IZtks0JepttcA1Bhb1ATR9SXmK4Qml2pKV7TtqP5FwsV0z2jrtzE7fC1i9k9XIah3/fHGGPjUcGE
QGtIqQZ/r3L4KBpVK70j8ZlCzD3yigp5Pcm/2BbOxh/oMO1NvEYg8IqqRa3EhtMYZg77gnrrje3Q
+cziOWIfe7cVwDpPEwez/wKypw9BnEfGwcKL6LxhUSG4xyOjW6Sfs+D7Co9PAZQxvny5HcVK9oLp
crJH1N34h/KkZxyNiaPjZBBeeuvyyLKDbcWlaNxRYgfmbio/u0dOH6ZORsoVprRdcnk67yvMecYi
Xr+Jkdc2QnO2he0gz06JAs1BbaKpT/4ZOh0EUQ45OpReW4QF3oVv0LVjRsT568M3H5ZqfGfj5DJZ
pzYI2HkO8IGwcjmkIfDXKv1rRDOLIyq7ekcglvt4IGB/j6S8Rbfhf+e6wB1vaMcv1k3JSao0Qwzc
qIBnpFhm2Vb4emY8ku+elok/dfBRkNdLP5feGg2h9ru5//+f/x3hNyy5hsc/pTLWZ+nt4pU13biZ
aFwKEROZQyn4Zl58TTGqyDA2JxUJ8mMjICXqSv/EiNdOYtVBZOpZqGxqD7z2cnuIhqeXdcAHZGW4
WG69Coj4TRuM9PirN/DczG3HMTvWzdonOTfKnfgjfe9R5fhQkxYvGtAX3XJCjhouloSYRzJUOUkB
d4wf+BoqxF/bFKiZ3riLktdMQBhOdUAvQPe5kQ/5UHxUKy4EYS17U5UPjcrlYiH2bR7/fCIh/t+z
+wBBSrkDMP4LNiVelt0GywMLPKTEMpz3Qf4ntUyqB0iXJvjAy3sFq+W8mZU6ZYZHbCCQ5NmqGmm0
09sRpoPs8DHZ3ldjdA6rZFOLxnbysIqmdLZutnLp1eyaAitWDSEh/A5FpnsqNm2up8+Psx/s5MMs
V0me45DGxeBHIVf2WYi1BXSfNWZjUuxBsNSHRB5vH46RKnPg68ExBJlGQQZpBYwu74fT4XpYUQ+E
VKD76BMHVs72ncADK0i7Mrg0gnfpXIcWgR7d76jI3xogsyo4q9XgCF1buuo6EEG1+M4Uhvo2NlGM
eu7vSdcORZa6Xo5EOlxyCIPDN08H8yAPEK2YP9eO8u6LSlb74+i7LEtvxzfrg/rLDZnXocgxLiHS
IBRuob6aM/sIbQl6I65FzB++TXeyOYV1yxzbYcqu5+xJpo2NialC7dZZMBCg83YpofDJD3raHBCy
ok+zXFu4uTnjIabZ9WG/0QdetBAdAduDOQqs9cW30cRfhUa2pOq3eTXpckhDHdxNdPHWCLmZMP4H
/Yd6VFWukHscHTx6PYnZWW+GLmcf1C6QC1+GoDXnEQz0wVfYBkMeBxoUKLy9LTFRW4yR9p96XOE4
Cw+ZU3OjUUCfhJUZrJxL4ljvhEEigwrt90MnY/FJCASl+KML49eIl0ZvVe3Bp1mNiBmJi4H+vo99
xfPEfMICX83s7x2SUkqNaBRQngmlzyx82F+YF5iaeOfVqbGA0PGjhmHr29p03vYehthfUV3+RIWk
WvcIuGl8I3qWB1Tm/YW5AK6j34IJTh+prQsAfSNn7IqOo/hpd2PZkG5x6J7hBP2nWYsv8bBWJXww
HrQ6WjKeFSQQaRZwvQ1SJz2DlstX8XwSYKrnPEV4qig4xHccN18sVXxNvJ1X4op7OQbGJjBnP7HO
QqZzs/8y7IhY7c840Nlc7bn3qRbYr1SN859QRT71/orlZ2/mjeQthZFtWzLXQKyiDCdeNDSvkMlT
ydVJdmgrF2S7xKxS4/82FUJCo+tcQ4D1Goye2lGvVNfGNvoSuiVT55C18SicHG4OFNJ9FXv8oTL1
DokOQS3bECBPCDPrkrr/72Vq3LJbyJT6hNlu373LcjSmf/xj81/YeTsNaSoE1kiu2LzyOUw+vdcy
Zei0ogpzCjnodaJtGFnz5YcZxKrloi6SVjxMrjCxFYSBXyUC4Kd04gAy2ZoBllzRrsXGAOCIZ/s0
X0XwVPH4jwixPREiNIfW/pKMzmytBx3pZTGgSoOtZ324R7w6y3i3T6tceFpRXjJZg3MqaIrO5mH3
BlrFc05RPVKZboX+J16tosoqcHj1Of3RMT7yr/9o3NTLYWB7BPj2ua/kOthhkJq75n0+6I0P596O
qiZz1fc86Joteod3LgcCngrbK/3LeuOi8bk0ikQZCxb4nXaptUT8eChgwMJkwHNiHR9CBuYYN6HD
QbIfc5OwD50NBY7FdIWgcLMQ7gynrFF0donaaCrxgEEH2LUqXzDxlth/G3XsuvTtnHhyQwqvjndW
gjC5zAicuOr8tkpyc250inEMrFx2tMcAFK1xgUMg9rGFTLm9dw2PKxduV93rjqcaa1iW8TtiZ0tQ
ZeDtndWtM+tR9sbX3DClU8gv6twlKhCU00BlcVcsoVlQJ1xKMPD8UyHFF5kSi9mXCgO14Y8cWGrQ
Pfix13Q/1u3rVN1UcoFB1z1Mw8PdHONnbDiotElWnVvOvVjjDmE5IgC0I1Jf9D+mc7erWiH4HbSK
PQLR9Prxr4b0Y815npFlDOYeLiJepIXWzwOHwBtX67NWXJo4xnEAJ+5CHz7bFlPHIsKDaGRV2S4U
hnZ0EURxsWao0JkYxeB394E2M7WvP5nU9MD4q1uAXuGsx/yIDFKRgoZBNiDSQFzaD4XgSZkkNgDG
JGRK827eGg24CiGYo7RGjSg8gBOhqUYczins3yNJKVlhvafU25aB7ouxxF0wh5iyHA9JBGP9jHGn
+ZN4t/oZJ039EyNsgn6KtfmsZnPOP6t6JgJFRzKho5Iv5wZEfutMZQ286O9nz/qtOYdri2O3crzV
ab+kBE8bi+uytRArvmKOmyOQ6XJelcoX8AwV87+5nmq6KvTYeVPK2smry83XBdw7dWtv3ySnVbDo
t9Dm5vGgvA41Y5XuMLzj/tQTRXuKu1WHrXp7Kdh9xHRR24wLIu1YFURsB9YTFwQQFcXIoBjNqlxw
6UlYHsbTJcEDRf6X5RrDSnsX50GgXThxPr983u8RkeIz8rRBf13tLyqOn6zsAg39qd83WthwpOZq
6xeRAEG+wrohhE1h7fSLZwQsa5Ib2D+IqyZvrgn7prmJ44XOCgm7NvS49ruACouHAOfLCI/z5gwv
e++JwwNWUTdgb+AYbgeRq6rUrU0HqYu4fG/LDaUy2FXsiq0KcFe01eGqVu7CKGANRmkgI2xCAQRg
oalfRP1+XInT3AQygzdhqQC/xCKEl8ZfMObHYN8wiPH17Rn6r+YU95s1FjMFDp0M1ZqRZJPi3md3
omWqjhPg17mRMV3g6UUW6dkbg2MBMEJh/3IV65MlAXYKDuYmOVPlvfWt7skAcs6yXW5W67q7Hax9
djoQi1eZZumPRxzuzKV3zHrSc6CicRcWrVB1c5FqYAbMdIRBaqHkzXe082SLnG87RZ00pHCmcDch
AlRZHDqCFBHuaojrks+x/GntYIAGyPK+HmJklGrEz+fRuhraxaw3xOEXDcQe2Ws8ZwbkQNVJG/JR
zqAXinyIA6ynQAclGSWLiwq/cbrcvama2wrnh/jmL0FutpT22BpdMg1l0IVPcuyROmTzqn+XWbD3
A8WStljzxwYaRvordlK8vW++MkQHFMNQ3kFQxqrYTRV0vVAapU4TfaOATcCxi6eAypSw4AyJJO5c
pu62YP2O079T9+klolw8aK4ML4SD5D5ebRJvtt8a7EO4fwlsOoOugjL0/Inx3tk7ow8GRnuMezCb
H2cXEA5sxK0sdatR22FTFq/8zKidxFsfvLyBssNF11fBCiqWBdeZRCGWahavAgL6KZ/6dTPunFs4
J+N0IU7H0Pos+3m37hXm/jDucM4jUubpFNtBpLdM/uAqy4pHgLFpEYVSQMGPMWfeEcnX8d/TCp+7
7UwteKGIddwlh4uBcEjL3wHqZyCNTj9oUkdFDWnYTjCIbIbRf0daPUhemahrQr9myUI4l+7f/kNX
prMhVOFuWOS7BlHQMtDW1duiAVw6/qmzdI94ml62fguN+8DNRo8o4Kf0EMXO9ahJVA38oIB07IIY
TZVny6PZ8htX/28EbMGL4Vx0L1W0xubBaqARxHmkmKx15CfCJeoeIqqrQDhyv8x04roSpLlU114A
oj3PsHv1NggQUW6pZ1dUmLPZzVjiONXoKr7uc6Lb0MBcWio5kYRgR7JrnTBDpj1XGVS9hP5zAL/X
m9Yw9taCURX+GzuVXcXmHa90+TA/w51vFVXh8fitaPEhHpuHkL+PXyr0mhf1MsSCRplbXHWmGKUw
nwamI7RDc+e4NWlGooSbsjtbIvvngCF2RJIvGonPno3tk3ZHy5/fb8m8aU1STzMBFxqCXwxzIogn
adVN3g9Z301kj6uiYJznP73+v6cYcDDVt3lY8yiGCOU3X8v5+uLIfz1HtB4wo6Mq5MerlJaloJUb
fezFcr3xv2IXObfowXfbbFFYsV3YspLBPNVHfGqsP7K3onzl9r+dzQxxmZlBiGw915SpiWjYzok7
uwjDL0wD7SP19XN6FgEej7sgWeRrRBH1csWxdmwuy6PgmnddF8hnNaqp3e+LQL04abstHYAvN697
3IGMZkBArm0dpmATI90zULyI0ibGSQJkmmJ7x4MzmIU+tMVKASV1n7LwxMWcPgJkvyVyn1KBuN24
WDg1X8SO8g6Ptxli3ok3TXrFL44tP6X9dPagadEZ3pIAdqZXiMvYMg3Utu/ANyQSGWqF8lD03nGy
bkcR2IE/7ttYYoQX3+oG6Ekj4OqYCClTVuMryga1N/dbtzk44R0JEvlN5m6QuHKu0tMwWgcv8czj
+18sXUX1nCYn31/fSh736xdLJem0tyg0IG1lHND4VJCgj0RIiScFeYZraplUQ/UlQTJQAkS8WJDI
KlawyUdsLuWN4TSD9maFZQaeDY1ymX4C3IFf1r1frxwL4r3m/QdhhXn1Dt6X1laZ1VtuNgc5l2nR
0cGs6IcjVjxhuwh7a1MsRoG7JZBtEpeVy60rJtPJ0g2ARAcObnKhHGYlGSOF4WiQSJeXtPaV+U2j
DRB8ZcvICdIQtYog0HsDcgPJDUqEUlQtBLZQ6TdEostu4Oh4DEmAb75xGvaJ+27KURrB9GrFEHrU
otejv0ISK+Ya3WVBaPUiAn/H7ghRh0vikzzZpa65/sNbNecM4YpeWoeAhqqjQAnub0NavoUBJ7MT
h8dIDpQ0U/4lcPdtM/n+m/bedHXnMxIsBEuHfiuSZ1SmMJs65IN7/souBPsDzXsvYmbtwQSKZyxl
QurMZE8y2dD61bpCbcIihzVWorAprQAjSXdxJ001Xp9A7rG/BblXB2CTC6JxARWQ3nQl/E14GTBh
3NxvWQh8uBmMVLQLL2NzVJW7lEFFroHAJJc0QdxcL515Kl8So2+mtcr+PnB+vzEeJBVfH0fY9eeb
inu1nGYooUFsF8ELaOMMmPdHEBArbEK3/NVL9YNqV0WY6ucWOkl3obfJhMaRBk1pd5E1QJckXBPE
DmeNGwPJ48ZhgF/b57sJfBAHSFoyL1uTu06gTmPE3n0NCMHMLbPsG8NjQr3XskX+TqYJwaSUzHB9
bCr14eDeXb9rTOX9MJ6MtwSAaebqAIZsjIodDe6ljDqfigzLl/xgpz3Cz5euld8zkwDsVph8jikE
T3LHgyuHZzc1VCxaf387pCotkl0phjHk56v5avp3rce0fTXqV9epdkQYgn9Z23HDbNlVEk51U4a2
JqhPYWZTclrbDm+q+H8mHFgkK7zHSOq8t7eKc3Nh31SPfg7u/FNY8ii4E+bi+yxaC30SR0Czfl77
/ixRSe9e8hrjvpbbcZNahy6xCIaeTfVbyHtwuoTGWwciR8fMtgKbekryH50/01XMnjhzD2R30gea
xN4BF1O1DJsyafNYwh10kQg+p6XzrWR7K22FODTSS38wUE3rDzP8Cpy45Vhu9a7WtZoa07peYbLU
r9LYK8Ka147d2z5YkecUXxZC5nQroVFakgymKggxa+w83JOPiIpgO6D/tKJepklJSa22JThWCGFg
60CcLaXvGovdXDBqeY6VXirI4g5dRkPPerEGuiuoaJdMmyEi1WDTnT2pPLMkvF8AnZ8wl+Z3+PPe
eEYmLUBxj3qTU9GW+phNS1ANRZArN9Up2FelObHf0RD6hCC9v7+j7suYU1CDSgaAZHL6iP7dsZR2
ERoQ+czx2ZOd2U8oDXKKUOt30tiu/nEGE5i5mj08dIQgvqtfe6cq2EpFwkfoV9GgfMJn0liCToWT
BgkxTgFQ+gp+CYYENi41lhQdrlNfwJMJ5wHRjssMn8NrKVFW7GD9N8Vk89VPztjBqClgQPtb8ZIz
BDqAoyh4AMK6ugtHZ6+C7MDGAPQlfIEF0FSDsgvFOK8aF6ZaGHMG7h05FvXeyCHu4srBe3x/edOf
q7m1ekpWnkL0hsckPqcUpPZ2lqIClOcEweCeC9wM4NCIwjLTUKv46y8iL3XpSbTR4FCWMFGUUcih
0nq0zN1iLeZZQ/B8H2+EMc2fO+l8k6KYLZlWAhvyjoWG9xt133d80JcYYoGVs9wf7txyUNiKgPgX
/un3n09mjCbKCeI8/MWNeadLC5VljG07znbwzCLNRm3I3HqTatFs6+duKuSmN1F3ykwWQ2cbKQRP
I1B17wP0EHsXwoFboqe7NAzuMurFSnDMVj7eRKRfxZj1VH5GKmHYpuAPvG9c228TwfsrhwR7cJWf
50/dRlJc+sz9aKOFonYJ9bKf4X9HwC0MgzOH96ERRse+x3V1FAWcn09csKPGj4dLoZ1mo99uqo9y
Xtiq8MsIVdFAaGl521jKXUg00+mKE4sNv3Xa/RHFJu68oStNstFSaZZv4sXBYVHSSB+3qdsM5pfG
2pX13EHa6esOUGdqqMtLybj/63M6PUcUmudlxxNiGbsFMs0StyMYX0kcxK15FgzafGv3g+QbTgvs
Ak+mX7V2sS1wM7XXydHXUQEXAYxtgmoFEP7jKdBfmk1gH0LitDK7ZyBcaEGdbeC8KlA7w4T5tGEY
azuHy8D99EjqRutAwlrLowH7nzkdMHLBsHCvsdTPIYBj3Fqy217WkWpwGgj8+bZwtFO5GLYHWDI1
l9P4RLQFqCvq8ucaMKfXhALcArAPTRam/AshEah7536sLBdPCU3tqlSGoRSb0mD9OZcfguFsiYOa
oPVyOhlBQxtCxDddU9Rgy+kgBMBhV2of8ObFvpUrQrILzYKU0L15M7CO+uzFbnjRa+egXuXtBRkP
H1S37tHLFNQLPDkETGHgKpuhUGFx05r21YfQqkrI7hCAX5TN+1b7jHveUF9VoV7BI93SsAothrDx
2a+T0vkYpb7O/Pi5DbiMok3+ku8OPYLwkSttWoo7GO003DFtVkY1ynEHjEgJmK+BDdnA5RLQED1m
QERJzHzQzCTTuUts5wcjjn5K+zTd+fq8Dt1QYbVkDzqjaoD9c3enORza00B/X2BbLw7SuMXjps7G
kizn4+g/a1WNmooYsy1FZ2IDay2ZLmBKW2QuuENOmEwl02CoBYwXGF4I8WLqGar25wQFi6gD3iVY
G4Rk3lKPbVe28kMiXjrOYmqQ1Kp9aE6lKd1mDYAsr5fT7XM5UTyWtKqOFEX5FzCXitVCOo2shHlj
JGPzV1JmLe1Ev3lzDpP9RQp+N9MM9K1nDuBE4RHJ+c5N5G8Wdgys3A8yPoFwjRr4uyzjYpbDhjvN
r+UPj5hnDIxsXVv9+xKUiSWIRuVf5EzC7DbNzPcXpfjdi64nO8l0bjc4wZ+VGtJ839c2xeCGZV8F
sy3Qb62wJGXKUUSoUcPK6ez+SCTNqlbSzFBDGGbHCLQf47cvSq0j+GpMp9Yb74g+XD4M+BDOSo+i
06duhRhseqoiLnprm5/k3mWaRRQjEZR393Tvmc+UmrwvubF2lF9QbHvtprm5KH2rwj2Wpjc785I9
ScY5wQp0+e3GaHx4LpVOOt1GnzutTDz1xx5cwEcUOptjGgN+WKeuNiZnPUZA1tw4H4WGEznpV/ix
tkQGvslAlN3uRX7j+hShWyLLQPxkCvMlUb2VJeoKDieN3WnjFOnZX0qiwLzMbDxiWRoPnnhjAEiK
GvW3LvLeqRZF+yz8oRGu1pJjn+LSHQT9ssqr8jIdJzTA9KhGyz/mSA7oH5wXUADQVkMQTTKbfAIA
V1AdR06wHEeukU7VmwLVClp5YD5V34fLxMMuXrvVSCQjeZuv4BWKVdH34aFpJ5OtYlgXMYPMQKxQ
B4Ze9SeZfPCyCX17swemNYi4YxrZ8nNkUcxjARzsD6RsyjfgHrUMrFvfHB6DFx5EK4WCzzbrmqp3
WRVw+D1E+71mH8B6iZnM/pSxNlwhDmo9Cp+K+/dwuBlRm5dktPFxF4t04NKyx7RsI1tLQ57i9plN
dhsz0S8SlPkoNR/GifDMVBx2mx7jTR8c/dob+QZWBpgVHsTTFT7+o4Gp2z1gLJ4sCiBxWmRxotLm
RrmBNCO/LDQtcv3RkCVBQH5iouYmfm+zNYmB4XWaJpLWiuPzsfbmjNdQeOV/AGHh9tBYNY9dx9Q4
Adhqw+TZ5jVfYaBSTuFU3AZiMjKIO+lPY7+WrWozRcHZnhGfxSAcmPCEfbINTWrLNGd+qjSw+1Fl
w2U2e3qgapMmu0CRe3ejbcZmyaugMRMMLYQJBLGguwgBkugWudtWShdk313F0Z/HajlvxNi06WAc
7gADY4/VmFE59VgbdLkC6iI4QTCmIMa1LzgoGdEJaIkCUkOdjQPew9W4CFe0XE6f0VquArUrcM5G
rRCm2VJIFkjupW7CvySok6P4ns8a/k+GbTXdcpl00vXtmNgf3+H00zAImuCz+Q8zpmq7QxB4VUd1
hA93AFNrPuRl/2BqAViyXdW+zt8/CezUQKBZOb4zkRWbBh4zKqgQIjyFc6rp2uqRmu92gHl4ndE6
nNd1kh4Aq4F+62YGgbCe7HRzS5CoZntRfyH8lq4LcBIpeRfkTGCcTXwUsiXWOokJi2Re5W4+g3NC
+EyfrDuwCueTQFnD9NF3yzhhcIkjqfZs9hTT6j5V+N9GyvNxvNxon4C/+tnhzZaXWqytM6hYSBMh
h6pu4vKk/gSSxyo6tlt6OnZ/gchxf4Bto81qyBZc2Xox8GpjLyN68TwGcqFJPBzGJ4Iwqv8kWxOc
tft9O321gx9krrulrhdCooEg9TlFeQb0al0wytm+vwa/p2mwQWTVEuRlRw3/YuIYDuvvDo0QYqTb
gFH0mPIW0g0IhrcWvxP7ZpMn5ozvdsHPGPsRx8nVj06UttLh5SlGeGGTDs46Wx8BDTf/Us/+r7Ao
zaqkdgimVVQu/vLVkLS1/JiCZERGi2Z90JrDbi8hQ/sPqyAzeaU+ImcpYysyAR8eruxqAF+zV8/b
1bnMwUov+mn3wlC01CqQCzCwiDuDmmjfIiffI/+SXaPs4B2xssYbS1+6X7Rm10xr5kpoCvu2dLUt
1onu9VWNL0K+gip/7V5DYJ+CPxph1EgS/EEXr4QiFt0mYKV50DyQ+IkEQxDw1rp5VVaCQvPtz0pQ
AW5NrAlE6kqC9guUcibXm7UnHrEzzPMRks4WYekFr2vIDbwX2fKeMGkdtp3bG69PmOkv14k4BZfY
v9za296Z5WeZrsidVmkzDpUmYHpDviRtNADe67j0KpsD2pJHtVDmm1J5cfCdKXrBcreJLveUrfsl
vtoZSMHg/1/yGDcepFkxzxO+fSre7+g6nI5uLVkxv4eeyZJ+q0wQ2CNb0ncf8RVMbOACdqWxYn+5
rWhOj1hF4050URZ7s+QhXdwiK+vC5CR4TJjtidNKSGrTIBd/sSrh/pbN8QCKL9S8UMeiYfvvGKvh
jsa6835G6GARDr67+Vm9Ve7nUHYeU4MvKABXPO3WJfP/AU4LwlFM85dBJwFApoSUhZRbIsbVM1bx
86qDFJE29jBU38G7vJn5TUdmc5k9disBBpEhHD6c4ETl2uZ4Ku+CUc38qdS+w9jG+fzzqvBte4DW
lr5BQ1o4oEStZH4aL7ap6gScEYvudmLVVPf77fCz85g1pQdUIPyq2KM1Q43Oo6cGlSUAYFuwcx5c
JGd6yJt17cV1ocqCFy7vbFJm65ph9YwQC97TdLyV+kgrjmFYweIX7lIBgZHXnJXYXSRW8HaWowj3
z4aU71Y4f2hS6T7BLpxgY2EWb8PvBU2etYgiq7SGKVVO83Ut4V8V9k9NaG89NH+vf90S3r8kcDrn
yeeWqg+EwJecRHB6uDMt8MRXW9W4epXnhIfodUbAarVWq67R/1d2dNjt26pjgCKH6BEsh5VKUeMp
z4IZQeFo0epgxznjJIKw1QOs5itc91rruryIExT//oFJzInVxh851Wfsvm+HMpBE/uGDqXcQfG6s
9bicEOtCG79Z6CObI11k7yn/eVkweHtxs74vg+n0WQ3jKaOMlDd8P9xHM4ahamG6r5Q3gBuYXNkD
14g6256KWLtc0pHBA3dB7EwiDbt0VCddxf6MHEWglC1Y8TjXOhqjo19kjuK/WpV73UWoIyXLG77E
McOobmrHueKXGNw5l116YxTNn7JM4IqZsScfOJl9gSjBcGo3HmabX29zp5F+zd/ZZEB39FPgeq9n
buqcdFj4ZJ4QUUaNsxLs2BPH6aX9EyhFMKl7RFYox07eSVK/GDf2S06rI+1YpPtYmmEo05kyh2BO
EhU+3k6HrC/Q7i5r1D4Bwq9hM9mVvMLh8w3U/c9xNNtwUyezsvWt7jiH+ioKMhKC2DAs+OlVFBCf
wSiMULxEER9ZjomN4JZJ8lD5pq9Ky71Or/R+MhCnJbAwR6uuHUYe3kclZbGnIU2Bs+tmgju4WyVa
VTf405mhAkG0wyimbXVq4/4eFHSywuSsTQhhSlEHRKP66UsGIv/sri6ZJQosSdd/AJUgtTPo7vmK
OeJIvrrgVbMj4LgQQht4tvafiCaz4IA4Ch+HfMQRo0MdvDtZr4rL3CNh3yiJ6KogwQI0LzxMH8U1
H7mIaOeG6OmR7pUvaTi9w2w24EMwbdW+fI3Q+17Q4Txhb6FkE0QxdKvQ/KRB/CzpcA2m7fv8uzRa
1FjcB0yOEY/GX2b1PIk1b88+ihSQwoIuQWYjCiCp5HD2yDszmRNFVGMAon28H7kMCW9Jsy/ZWCmt
ASSCGsG5x5+hNyeP9WQk+ri4uF+U/6f0rTda6lfJDrLTX+CqkG/HoLG/6rLX5NBiGfny1eMTC2kM
xDHWhCSz38riKc6AKYxqrrfzsNX4/ljr2CejI0KdKbp13KJMuk8t5wJlUxhMuKNKNmlx8KcUZg9Y
xg2Xh9wMtmDtq1VgYIQOVbWbfUAMok6anC/mKJKsr0BX4T/F1aWw2Di4phm/SWajDAxJkUILWqxe
zsbo3fOMrqbKQ3n/YAJV1gr0o6rDTDaniqhsoyjkOkIBnoxFkw3DO42XlHK8hAhhFYwYIgwW/zK/
YcC9Sh7Dk6urkoM3gen9B8rHiZazn8fQBXfXznUT/lN8jtv/9HFLIgKa3gDKf6YIQs7sXNLTpPSt
c9cjFQB8SiJvjeVEw8akOIIpEJwITN4sh+7ATC3acvlYnDBpntVVRoV733lajA2QB5IiuPSO5+3T
pISXG86LC6rXjWJEz+RlgYE88X5pZRPqma/MjpJWLoHJ8HLfgsP4r/TWlbVrai17GfrTNdtrLdtS
hSf7MR4VaoV/hCAqGPH6/+9Qhn1PgMG21+tmg+GJyDglkPivHy9xYsLfzU9TcIE2aY80S0I02NGF
u+P6MNTh6kaiqXbVJfgBUbrpu5+dQsbAu/8nd5qkztlDfcgjD4l9caQR5GWbKA9VMO0n1SAvoz3p
oAVIbRQySkKTPnOwt5vRufSzr4l7cuo3USoKSiQV9Uub3WTM1rxDDYQTDmYkm0BoRYjLYJ/uCXIh
oyzHwF7VWrJUQOVDcpBCdaJTRW8dePHqXoF1p23kxv7x88779rGgOjZz/g/+/ZhXJ2AA6Lzwzeh9
tsmsOnHEraoiwYvQjspI11PWP8qgL+ODRWaRhpuSf2g9UTgaEgggkUsyo6aulXOOUu2qHg/aac1Y
ei1Zj60vwAufrePj3wvKISc2LLoNsfaDy7LgL8zvSr5Jgp+QJpSPuWmf6FVV1iqFOQe8tkmsDgkk
0/9Sk+IsYFvHzhgru0JndZL4fSfSrfKfeD4Ey9VH+HlKov68vvYu7OKRGkmPJNwWGQlwOpYHcG7/
G+4gsGru+Pst9sX1nDUnukRspoZNa2ljkjSUbKVMT2BkD5fareniZXKYpMvC6F7yZjXNYk1RctKn
jz+Hik7JsOvL8DT2ACyoNremqwwnxneXMf1hMRuVRsCBEPVQoXwsruXoNVkc0J4HlYz2BkSiA6a3
facEAveSuXlDiVcDWyyVmH2C0CyrqX4wPTwPIkCBcoSeTB6tWXLR2bGlat7nmhEBecKQtF73Rzxa
ZhfpAAgxyvgxffBKJsSJdWlGgFUvT4uNgN0KH9E8llk3uK0ZBLcYQr8hOp5EP/8rQHsVipk7Dgv4
dLcBY1u0sSjJKl17teTOvu8/TUSUZhSit9tM24c/B+p5wfVvpU53ME376yPQEFCjpgx/mlZMDNBp
orsnYBqEHG52/OkxJCySvGiwjgEEoKaLxbQmKIdnZ48ZJ/5SZoG217Es2mwbeSRX9U6odbM91Ju8
4mYs8Htlq2MmNqaB9CDjVW14bKrxrWEInUyU6zb4v6uuFydtseSnHiUUtA73x0A+y8PqtVQou2lo
e+owbyKCNiQeJWZITlssddm2WeIKiC9lq7T55il8DJLEdEHBs1ukFZxRL0i0GI3axHju1Da6ZOKe
OuZrVpMypQYdu0afvplOoWk9twsnCZDkbm/w7E9CRpg1OVo6YzRtrBRfzdB7luoYnI4EDNLxdW43
Gr4m522INS7W+hy4iWIgYazFnvMpY5w4E86u5NPTC6Ej717IViAsUT35C8y/168vvCtqw8dgpIx2
jTUeXjsg+BagCwNJopOCQ/ASWg52KsdjlV9vuN4sc0wuUtXzoUg2QGBLeF8Ur/pEGt4iehuFODJM
Vz86rXy81ixAWsCQPcbGxzdF7qa7eKuHNOs1+F43zeGhDZGOb6DcR3LhH8vg3NZUO+HGV2g26OcE
LMeWdmNlCLN92jB7RoHBqlcO34tg5DR0gVUaCKZ8ELYe4z8fGaqUOGQWgZyYwPW9DGcTWQf6+zim
je8bl8T+JKslvUrg3kXj7qMDOSjsHrq0t7dIQuP1+B+UNhqVkZdsKgjSXrQXeGBSzld+AhmPzr+f
ymQKkJ22hfjsgG2aeTzHdq5S6ESHTKPR31N5aXFVaHKRmaB8bZuZzxneoNTU9KprNccgkAiR+dyf
+bq0BAUpoi5LRajQkJzVKUHHUshUMk3AhgQuHDw7SWv7xGtK83t3schAb1Jga7z701T9aPcSi4zP
I/UdufDme1idIqeet13O1vOJUHn3jYYfaOaPxtwdCYuUHESOdb1/goTuc6+YZT5y0dwEQDX2iOMt
DakktsRs8X3Z9w+oW7GVmQph1SJvURXNpgjntRmP8NS9mrKwOMs37a7cHCck+Y7FpigqzHqAOEKj
2z6mdKPUocFN9RpwnshrBWFG9AnTHbiUMROaFQtG2bnUe7c3PhrBDryveS/u9floxPKD1NfsQMdD
gg5EdZfS9/bj/uWhYJN647rkUXMSfUNNSzrIwJ3tGhO7PQTmB+OjYG75q4mjCkbJfj/lf8X4ADa8
z1W+/zVdUvdkUVoqRkdV58DI/aCnvEmvVYRd6jsPg7Hl3Z0bXhLJatv+zMxJuS63clv5RR6vGFW+
Ekktjx59jyoJFIDWM4UYEK2a4qnl6ee1KZfGNX6V34iL/cqc8AkggO1ZMJlZ5RH5IOEkVRcBRGfY
YwYhf7CSSdMSsV4DzO46tMnyTdRhNfbFTSaGsqeDvaCYj9QTgPCjj2yw5DfsGtIgjV+mrDrjNmZj
rCjgMANDuK3yGF79N7SsLbrEg0oPQujhYeshTcMOH3KTuY81MuTAjp1nHv6lrtGxyq9yw5siaHzO
4pXLGWzxyP3h0dC8d0Gr842gEZD0JJvlNmZGckrYmHpqq1cOR8UWfNl5/4v3a1/Jvo09XylNCoYQ
MVtiGjmeoKdZEcMXZ1TL/Z/NWaidtRMtiHTokOBsDT5p8sbmFryeD2tUYkXxxCRt2xVf38BQe9VT
as/ot6RusLFI3EG3D2jlQGNOaAU7lnvWZHvLVIuFGuY4w6Jtea1qrul64Lge7rvNFTGeSdlS1jra
2aNcrraxm1fCPW4CcW6ohR96GFq/NKS6ZLMfsdJ1QqaA88Dp0ZdFMkVR5TjX/h5Ej5jN57plZbuW
AgMx7+7hDaV9spD5whu1sjDNDf43bnSLcbMq4Su3F2Em+7rNNZppVuQRc+CsyfgJsxlxsXSpF5r9
jaKQgRZ0k/pApljoPx5N9sPmCzxFQp7cOjPqPc9RXELktSsS9X2fcnAhlbyAVqhQw2ea7/rwZzTO
PIHQnmZc8wfoeyCR4P1xoiXiosfGpyuIgYtK9iGHjp9geVZQy+sqMXrdZiYDRWbbmXa4xe3Rl/F1
6m8zLT2JL+ftj7M5TCpdDGG32YfiNkaxghQxKgsJuY0sAhhQi26QUknkUJ7gviIPYNxO/cYCG1ie
uUkjZXdHAO8pb6XtzsnuaZD3ohhOhvqUXkyyqducCcVXGZCewpMK7NYq80rY+8v18S4nBtlfXAar
E7CCASS2QxHuJsKrUkO2/hxCWrZk8IkLnhNqCh6EbOKKjF/Lv0c2btXHHnxGtB0c2l9wm7Ldb3yt
z8xYksQiTp4BrxDD7BzOZOPXU1aRQCb4U3BSZLyALGjuHlNGp540I0Z/BFKwYJQAkssAUmW79puU
zK1xou2oGRP8qqkD2yT8wjP+/5chWSn8RwAbHS8HpIi3+z9evdjt+b8fU7rn3ZMcjnF14RE9Njrp
wVBe3BvpG1MzBBDpZc+WSYRuibFJNRMH+M32+bLJoxkfViC9NKkV0ZPGDPUCbnIRqN46EBqaxl9C
LkS13jS/qlphsxJKifs359UdN1FQSlNMKKrzmOJwuiAJtRyZ3EpiZvvs9SZ6DKd+enUYX7RIHcM7
t8yWwJI1QLt0PyDHbUTfgodgQINrWSyKdmadweU590saNEwBN0k/dgh+9OeMGBqzaA7EMwcJ8T5L
5o8+4kZk0thH3poDiggNFf0cZ3JNOuOEgHbROW4QkL2XW/+mjvEQ8lJPV5yNUZxoZBeXouuz738t
lTNPJl+zVGagCQ4MTXs19BijzaGPZBeBs297wmxDGCzqK1dwOvMDeRM92tenPEycKuukMk4bFQWy
34U7cdXOMsnWYTB32bY3BuiO3qz6KBuf6TOlNnk6lawlyMyuOeEIoqGiA9JcpvCwbbrtuZeZair3
LTV/fawmiCQNgAozpZUZUurOeXSe/G96l4WPyR7ma/oZ0XaxoxbvaYRAzPX/Fmxs/hMyQmO7LWBT
Vs3UEeBgoKCQ2PX98AYybOFFISvlNkXPDwpeV/kPMbCPtyrqr10WpjNhKda1wYhHoGACFMzqV1ra
+XNW1MtoK9OzUkEBbtwGhrBJ7UmUX6bsNDacy1GztOaOrQ4vwr/OvoceGdV7a9eiywB+RJEAw7C+
ldczZy1xSCRnHnl5f1e7UvR0a8tAizT0onHfWLHPW+cotklWq9ntv4P5kJ0ptn8LkjFHw37BkyGp
nDlg4gvJift3BkL1UtJJ1vW+Hz+a7fVTqkn08FHEZF89FHWnGeyw40TmpLnliPQqUuu73Bk3i8di
OV3QqFcwTjucxkzMcCpfGwKoE35D3LpVxZE6JhXR0WKp1sBfG0DNYI5/I3u2BsarUvrrlTTlH5/r
IHSLbshmtiY0xmj1SNzP0spTHkfe1LFjmfqWjk0B1EZP14oJpGMQpACEFHrxY0Vi8m6S2ByHIQAx
XqMjJvUcU0U83ChlI7MoYgb2PK6VHxr180HYgorFH5T10QbiNK26srQULaCQzAq1wePYp98uiBAO
8JmrbtwqzpbUGolSShhtOGJ4iYjIj87qO24nH04D8x7k114mKbOxS+vV/PQCoTI60D2WxdveYgAB
H3KnK6TAh4FfahgHkNOtsjXzdj8vJPtD+dsvfUbGP/9xd+ZJqzCQwB0lCOkLvTRwaPL3cjH1vLPx
+rlSwmTzSWr8f7gG7h7jTTKSXTM17jTJqXEHtbNMv3MvZuG26Crokd+G+FQsGTz+axLLrEnhj9ob
a2vEtpdVZIfoYY1Rdfua7NWvDjies21isa44FLdUYf1o49+yz8ZjFQlgST6964rzuGlnu4BvgT9B
ZCo1bpDGL6TJLi2YNSwiZDqDElhYtVhtmIYrXDrX/3M0u7fR4pYvWEtrWgM2pOPCas53YO1OiYvp
Zrutrg5+sV0qYdgd6WNYEF+xhblMukIm9tsIIuqCWwyc9+G4BWkuoYgV8LcnOqr7xlLRE3rGjqKg
FIaO3NedTvitTcmaC7RmD67vHIvn+eokjwqHPBQ5h/lymBlMrMB8ALYlnQtq1DTaw4+IC7LNY0cd
ESf41GVuRY7iBCkCjQnRJALrhFn+ZJvbQhvmuLfyF3ocehdv8HFq3sH0qZ8WPCllfkuxcal+VqNM
CaIWeLIPYiNCYSClBTLxHiy82NHBgiiIVNrwX2tklTgzMvbViMa7zmU+BltMkgMP+IgxLiQVRetm
FXbwvWznM+CfcU6ywjk7XW/Rn4kbAXpFXLWRhdmW0kbdIvx5SfUvLtXe1S28IpY8USMZ62kJxw6w
KhPTbhKJviXcjCRJvu6fbikYrXf4caOZeen4uXycOIKQGU4FJo7mPrieEi7n4H+SJ4QZPX3wRd1+
yu5NsSLAcwYQN/j1sRYGaWRhqUxDiFBUrTDtXzZl1GJQqXwDsoYXNNOUnXGkoSgl3JUpTbSt9cNs
0Fsf8oEdEeN4ETljuwxk9ZygQD8hy7UxtsWRQqIqJV2+ab1mIkFedh9Z0tpy5TJ9vWDQXJncOkF2
qjdaX/j9u5wBiEpWRLZCtsn/miwnrqXVw6JfWWyfQ4aQfvQ+2YbWsBD5OXxEUTEn+aUXHkeYw5Nj
GaRuiEmFcIg4nrffyYU4d85xKGOgh8FJAnDc5HjBBw8zYP5KeVcxh94sZqpD3GyV/sRHwusN6WnU
AZok7iv/axrHFCMNuLEhfQVxLMEu8g8M5RIpFlm5L0y7CL1AkpEK7HrqY8veYJKUiuVFxNVCLZN8
MkBcRW5eCbCU/L1AAj/ZCg/JzbgFmCCmG+CYk6/HYvH5om8efs3MtWb4wfmMrtzXptwcYTdzDmm1
qTrShndh8DP1B8CrSp1TXviUopVaQZS9AwODvc+xmPcQcN2VGsTi4LrENf2FDswa6zzePw3J0Va7
5AvziyFxUctXxyf51pSTO9en4Rqf1U3nyPrmt4fuorzPBlS/PwiYxnJB43awNp9yig7lQvsABqw7
/FHmXqVJW5dTrmcUzRFvVZhBb+Uz1MIwgZZKhu3zCoqz3bLcK0D+TQjJSxjV/8cioUN+S5SUHYJs
tMxVq+oeaBVh8/CItBFkgJFvDywdbmL1NU60zixJhaWY7Vc+Z1jDoBx2hADfTCRz196j6kLXgpUm
qbFZhWxmaxJCOTH4sguatGASVaJHAYRaRUk4Q82BZZRjLYv78p+dPtXmSNg+u0k1MNZXJ+JlAxJa
63gbgPKHxfI99auBWJCePcozqWuc93eJ7xE332l+4/xFdbIW1rEy9GKIqQzI8UkhzspwMwww/q4T
IrUi78K+VtNUs+i1+iemqLwDhI5EyjJzVZ30AuMLOIXb0g55GNMP65l3E+0V7Hn6XnShyNMEQ6gr
ghnIKcaXNqGvlQWp8dt8MV4pksPDx9v1fmUSRrSS1NU3kFlqAJRKOJ/KGodCKdQACyC4sRsW8gno
L8+cg53Xehry/qkx+VVabFUuo6gmFtQGFJ2yGIGun2HLqJ/w5H5rYeAG558CS3gAx3ovMMw2Qb+1
JcL2bTTexot7k3o9x4gLbt6kMoBjzr0jTt3GEL0R6aofHZXVAnxrgoSLpev02nvhX2cw/JBwOcht
oC6yapR5EWdNL3MPOkzJbWAq/2MJpMSdZyarXraozj943QRqI9HCcRTZp8161apuU6hNg7neY4iD
0y0p/Dp3QRQlMndznHt9fcd54+oXZSVBauCxffp2AXxS1WR/oYvUl1gLR7xBmM3+Vlo0NQtxWX/F
gVjz7R5w8sLNUp+YPvToAXZEmU8M6c4F0IS9VWdTA2AvxC7RHap9gzroGgEbCj2mSY3aEvAsH06R
58Rn+JNh6FV0lQFZLZcmXBvrUvSwYjfDyUwvkj/hJxUqY+T9LS9a9zQvi3wgrfjcju4ICHf2zCfW
fBA17G9TaOuc0bzy+J6wYHGWu4NymwfybTnHZytLLzC3vkN2kFiPcvkJLmQ4k/bMsMhnbNQZAfhH
lTWoR8Li8+cyM8Bfh5a7+rWpQ0zYmMRDw6mohiDrGp/7LrMOzKdubVxnpIN7HuMiDaaeJSEjv544
PEQW4+MU/iXSBu7rxKW3vQXkt5ZkXwSa5wDsL2k+BHoLkHdEfVUsFWKe/EsqzbSSCU9WixAEiEgL
+tSJqHLVh7+GQrVGEFPTOz/NQQsNYGmlDrgif0icql5UnfakWLTc96UnHoOc59fGkmbDLLY7+ePc
TJn0hrszIGa3P5mj3P5fig1oV2oSafNaRBEkYQbCBrvzJ35NwFf28THTm2NUKGVyzCYUnmZ/1Ind
LYs0LrwhLuYWDPsJhK9Yaslf2e4sc2uxVfO+EFOiDDWsNRKIyJRqTjJEtD72A5vaJOZE8ZwU2p7T
mFgiVTaFNgTFgHgzxVTsi3peHXhaRDTOG861l6ifpcDN0vRa8iEVW/7Ppu0pOuKLERN+6RYoZNu7
zNbexHUxNxs0W6PohJDgWMWkrfnLXsA+6ywD4URtASPzikdQ3hjTSOJRTQ8ORQO7hk61hBkSBZv4
rJ/4UaYYeYIhFv+Lukz2OhK9XqkgTGUmcHwuyNcKnybbUSbOfHpHPrlQbsEwb4hVwY1FLCdZRqbv
tMiVQQlWYMT3Fx6V5PmKWufPyjudFK0mYHEy8CDKrCslyrIpGQjuT7M9oP6gmWDqiRiDFHgsU5Fm
t2PZf4xBqB0FJfAAxd4V9imo53pdTjAqHDGhdcrKqW7wrqhZAdTHsxu7Jdcy7b1BvwtUcJm/C8io
TE0md82wDfhOvsc04WCIFQGCPgCLBpxVuDO8IynVQB2MDK5tY2Z1pmu3AzCC+AiSxLwT+uDryTad
2VGjcezETXefS0WLYyxnLVdsvdF77HonWnU08yhMD7Jk7rlhmihXTjgFKS1dCJvWH5L8hcbgqG56
hZsrK1wxgT+yQZaiC5vPhcfqAntenGOT2Tfr+IEXyyUAD3RyIkT1EMT7Id4B5+S+zPuaz5yUIZlS
ZTvOC01Q60yRgv6A4SkWAtKPAVs4U8UYlQ4Jm/i2Muwlqisoepp3eTRb2/jxBTpp9U7NxT7FyGhw
d06x60cP5TqkArLydQYLwGJslx338MIq8ur0aIgPedX60jkP7z5495fjIbFbnJ51X2B+DS6HerNT
U9ks0AQ4LhEXAvJg6XwKT/+n3A4sMCCRKhgc7kd0LUw4h9JUZ5wvTKV528OI0YMfdy2Urp79Qg3K
QOxs1GrbCSRh+QtQxZpXq1xa2kbNDWNVtuS3nBjoTOlaGjwoRh03Wovz+oOoq7ITXj3NSYzvhk5D
2v4FqJaFn5T8WwsRJ1/RQpNBDK9fuPBDqgtUYK6L3cFXmSYU1KXtmt/QBPgBm/xBfVVNvs6tZzNR
ge8qvRDkoDkzGIRur8SHz/AGX2GmN8mp1mxjKjGc72qzmNwvP1NsZcYEwqUOTwSPNAipbiMir7UR
BcTVP+klwWm3HIUEe+7c+hOUZv/98MD6Hue+d9fQHY5gLCcAulZjbRxuA6GeRTjjccFcKXZo+JSM
edtVxzldVDFOuUG+/qmGVX8Lpr9ewt68SoJ2Ma4httVHZ/TwBwAGptm5uYI5L4xxPlNEe7aJAzOj
/U8IPB/S19wsQj743MWM68Lws8c7RjYCzEgkzCHcnq/vLwO5XlOH6/Lv2KENLo6Ut5kNBa/hJZmH
8pWgyiWG/U1l952Z1N6mMSTWwtoSyxYdpXwNCPPh4g4XdE5SN7gcmG48rvn4IPlE2zndFasiBhFv
GFokGCkAHs97c6RWXd6ZpCpaYnpwxvNCDSOoJLlqoMQm+xZoUtlLP2YgPsTj3TWsfEcqMoFaqVxI
CqVgUbAEpH/GGm4x35RfINfXsVP+PwbEcS34YBxHaOOkmwwDqCvi+ElYIauKWR52PdQoV12LHZCK
l72mIZaxLv1qqk6apBbFWiM+uObC5De/44MY+0qHrj3rw2xSBaGfqb1i+hIrP0q0pQUUVFz2lh5d
0Xpe1dzjOtdgbVgdOF1mt7ZiCk165X0b58GEfK/ll+Zb8tm6pSCIhna8r2hNRK2wp+wEJZ4FwJjY
ST1nGM24S3uiSDGBVUUQYZTHdPN3Ebt5EwFsIPsT/VVtcn2jP8yYlqzgRszlMlUIGfI9wPVeHwWf
2EYXwBJZaZalDpoZr7xgRKd6Ni+V/wLBbKaYKBHkJxQGwmpriwQPuXg2pXazzFZrzNxR8xyi4nAV
XAcQWZbD8JrtWfgqDKyMWeLk8V+z3Okk10wSeJmrrppvIqOBsP920OM6R/OtwisYvnnoKLhDWe9y
uq4FU/wSN4arPxEfL+vhCHZV2Y3poqkAL99OZdOMSH5sCogfloEN+3b6wmP63UI+E6shGdxZB127
p5ZX+8feLwScg83TBJDVN1Lfyep3NG8WLeUhsMfWv7QuajcIFfq5ZrPCurgyzPX2rssOiA6tyqxd
rkLxum/PbubD5BY50lYWiHQDkVFa/zJXWFq0+J1sUoiYk9LuXmA1x99dFqqEVtvPzfVK2xwQOIIw
j3r8/O2eZyUXlJ9o2vQGRY00Zquj23g3RyNSHrqLGtXfCBJawoU1E12EI07NVMgyJERIn1x/Z6wP
kZA1YonJgxcGVS2o6M3V1gCMDaE7OeJH2NWGUFs5o/JFXD5udkbvVlOOHW7WP9oqCzZvh/NDw1BR
VYksE2FgJGrqm/9uTlZgPr7ejEQ2ZArMD0uu0Yh9GeHeQScM8n8pgiPelqufoceoyQk7LeazCnuN
vP79I2rEnI6xnu8g/btZJbIOBsZlSgD1wJzmgKggpSY/CoC0F2QxqfHHw0rzKEyh3OoBYicsN7Th
FhgxEvi6QTo0oz/RfL9dQOn6/jETVCsjQNOIa/W9AhWffdY6V2I3LV3/sIC4FT8xxkDJgKdLs8Rg
Aw5aVUg9LOoboc+IXV725410Kpc18uRmK7JQrUhSX/UhsG/wIpieiX/G66ikEcEwwbyNXohscVuX
3Ck2mygBWIjkcvPk5BV3De60QTLYFlCwGQi7edGRzR0OrL7P/mtEJgMhRFsnT3lkBX4hp/Ii+QlO
jlguV9s/7sSK+yVc/P1MiORUTZCphsn185ClAQA8pDdG+Hyjf/4t2zj933m0WY0i7pgo1oNi/ldF
0L4OgPT3r7PhOu/VTlDt2pAKNiXa0WC5HyBUOxs4WkuN/UAxfK0raKEtZy8sS2Kjqj8529TanI2l
IEsSseIgEivitixw5X8qWaTwSgV4tQLISlJ3vEmvUbilT6wDyox4kxQPW4+vqOhrSpifMcsuG+HK
CIzegzMYliOGQ79HZ/vS4xQ0McOoA2Aq8FF61Vj5x85zdgoSsdV0XBHNByLrNDVsNrQ2DJcVJ6jy
011rIBzWb/eEArHizNNfMjhOohC03MCY+psG2FTebNxvwQcLv4JHlfP4OuU9/gkoz6adAUxVqLFs
2EEFxTCnLuh1SGcQw9uRP4CWYtu7yfuniY4/E4fx3qRFM64n0WtgM7HRtPA473r7Xf0Al7kLvVq1
nYktIlQYRW4bcnibggiR40VOQVQ3NaNHmJyZIK4JY0qt5RL1F3HKYnclP62QIMDkq9+HHh50xcu/
mgnr8nZPdIk+/JaZxuXj5n5fR/4Agf8Ys8oPlFAVxRa+nix2QT1JFZzKkfXo/sUbgar09Jrs7d0H
FQTarwBuYi3CeULAVTbMrHM1Hcif43gP8ALAHR2HU5OB3HvnkW2FB9u9qm3kSkxLxm/MBl/FCMGt
X97OhbRkG9s1QOgoLbKbUhQJhl65gL3uRjlnMHODMUcWS4j3s460xjANTjkp6ZYQ4D/ze/cJ6xVI
nwN5mqJityL33EY2Q4iH+ZUjWDybs1m2jI3PmkRWqo3GfjRI+yysWQsi4GWmS6y3RnDyft4W9/na
qoLxIo2KPNAqXqBCOnhaBA5Ov7c0uTfK8SiJbnDF0k0Q8hwyPnw3xqHsyiLJ+vmSj1o41ZGQNyh6
9IOXsHZcPfLAbHeAfcRLkY9pO0bEoqiU7cedw9cTRFGTcu78UB+UsI8tTCrDaI9B+XBYKFdl2XWL
3f+WK9NzOUu4SS2F2QahugEvNh7BtKpg7Ts87eiiX30lxLRrKQwKaIfAzMcRMwVUmDZ/ljLEiS/9
Ax7jcwzP0Z/SQjRLIRQdK086ZL0SS3/ESTV9oKiSUW/tPuGKI6RpPpfu7LqxXXBWUcDE9pxC/tXs
HuwvWZgT/1y/e+C2tn9F1sz64uv+P+Q90l1Jf7sC9+z3h0luCE485MJNqETwq7RDeaytVBWX1UiM
YNMBPt36tb09KgMsUl+ALjlKfK3L83bDhzreywFfTpp8Bo9zUPTaIuFewBtuJIIMPsUMPJp6JMYP
+9HgKnc4AFw+6m/9Bg/WcpJGcJhBiMUUW1/H9y9S/GsRzj7i32hrlkS/INqENA3Qsd/WLHVBwtn/
brwIJ+5R+F3wWTPX6h8iCYPYVnIgUBPIfhaZj0tNz0EsxtF+wVUizKVnxf96VFZWFWqlvsX9pVRH
iME0tcxEEiSbh+Oell3Eu9insWUWlll0IqR/pnGkyyxYtX/h9UErYXE5ekBrPKIGXdZ+YOnx/NBa
1VtOglJ2nkZRLhDFXXqMBSFErxsO/cDiO5jatN10n0XWr7Q2HdojKt3sTUComNKSTtVFsEY5JPQw
dQKTpYM2KqKHJhi3bsLID2lDoA9BbtWumfjw2MTdDrfSpjODU/5be4vIxwCowCwz/S4BBsZn1XZ/
+9txVkFYdihpCS5r+52kAA0sm3JZynDlA87mOKvrbDRgQ8cFvQnwRablh5wCf57M3IruJriYRE7q
4snkffDwBZ6xCes4Fg/isrZrP0cKwv+j2LNXnecKfn0ExoV40UFTCEM7QQpDQq/e0H06hvhxjkCU
k1H2IkmiXZqjV8rZxkIA+ERQ14Ph3wDRa4EldvJ/Hb5Gm0m6mEVOPrCz09wEBH3wlLo+n+bEsl9V
+FH87XWVU4vs9QmpLH90yDrzgeRT8BOsZdbRowO2uU0fhzhETv57cTYTiPOSlztVx83sedypZ7CW
4Ou5PWJSgaBjZgHMkq18eXlx9cCDpCV9P31nPGyhAo/X5qS87gyMcXTAF3dJ7oW6eWC5tJQpi5qD
yP6bLuMrUf3lTEGzu0ftJWOwomIpdSWvBCZa5RaTGyKeyDRNwxuRLeR2og9p3lfSLYLgez4r0mzO
tmDBLPKeaTnF8aYxzOpZKqI87MSYUTATuZVfD9NitmRz5rWDfdSCcZxACcLVcVZYrNvDcJw97iZe
UKR/jaz+eiUarilnBpTbKRU4+mXn9VujAV6uI9Bve+QjVMMh1RgOc2fglV165rOEZ52J1voHQ16A
LhOurp8WyoWwgsjE4n4RmXkS8QJHuV690cNsVDrRyQ80AtrFRn1boFuZ5Uxw+6P8HSA9X3HD50kb
KyOcepQuB8jNtvLqtb3vPVD4u8zoSal5jPr1P4XG5gwjXT6t86W/2sTeoC+aQNDzxoZH4iYfGbiu
/h2P4ORE9yWldnTBgH8x8ZtaCQk8HlYTYJq8dIyJ/QpFZwVrqO+Cdavz0F8XtS9I2YWlaff+jFp8
0KNTm782506kJRlC/JcC5Pk2cvV/6u/EvlJZyeafMTTQ6oHUAIWdfisYNl7/UXJ3zCWvpWS1gbhD
jrmGsB61maq8Pi0HiLec4wIGipRtCGNz1pgw+42hyqr15xI7gu+UWqo1LCCrR/r9ThE1YnDrjBvh
G+3dUd/AmO+6ueNcXcYF9aRn1ZHgNsAqGe2sRr2WdCTow/t56hhh4OPhNLaXH7O7Kq9UcePjDAeH
DNlHMzLiVjppyW1yQsY65qTTE15XBGubzmbuowJjvEPb2veh6u94fg2KK9bBXsQgVk4dNx3eyEms
VV1cGKGKBpCtwcAaO/idtwCj0/s0o/oSsfrYMGGKSw1sUQL74Q5zbZFsTp/vXB0teursGz1th6ko
nZJQ0+JAcmEmodtBEhT8VhXKVSms9odT6yVfy4Bj18c0xol5hF0nJQ7nn2Lo6Ur7bTJM4yL+B8AX
4RU9TgVtjsUqN4UsK7A0xZuVPEV2QU71cctxl4yPzanNZoP1G33Cth/z8HuAZCi+W7JYp0s0VRzh
cH3ror7rqZ0N1BySTQ/evhF+ZN8LUafeJ0KmE6iOuTY7/9GidzSnogLQo3rVLA4r00G6NLc8kWe7
N3IpBmk+A6V30AAjacSS66YYbe2kXBp0Ys77911Fe9wEcD160Un2rZu7M9WPq3fa2XC3GvGT3/fG
uVRCyStzCTK5v5wD6z7IB0LKLmb/jK/Z1DNWw/GrnrkOf2rS0dcAoGt9KWoelNIZ6+VtYxeEHgJM
zDHfY+xMe2z8V0Dpq0y+PpwQIjMft9YrFQ2Yw/VntdUSHn7zx889WrxMMOmH4mduuWl36mvl6Bqi
DZUPqA3jh7psElsFv2zCquPbCx+4tiNYmCA5yB3FqLHTMWV7aVsMxA7p5OzhJt679QWOCnGGQven
KGwkHaaVZ4AIt1XAEHNaKY48u0bwqOI8jmBstp0N/HtVAj8QXYYJBpV8fhnE9388oyYGyFUZ4J5c
4KHnBU83T8+aPeiZW8gv8mMNvYS4o2E9s2HrBwMgn3+ZOwaEo1yPoB1ywhW2V867qf3b3vVyVpqO
/ac8GWHk+zD4GsexNTMm8jkueMx2/CSU9ShC1oewZ52I1868PlW1kitEwq/rPaFhHJ9MrkvGu8fF
lqeY0fcwHhkmQo5PFdosZH0T/6jlePFBeDy0JTxUSpln2u9UQ0DZXmTn+2mWu930L7ULdz9Mn7Kn
YnlJbDygXSEKB3J/PuFTPe9W/q5ZZsiIZ6DhMJMJ1l/Ng1w37yAXy0QNAtZr89Ltu8Njh6D9rSnZ
rpq2YMk/1XP2Ai0NvwPaFVpVVz6xmnmeHYLzDQZUGi65yO8Tu0fydonOJjO5NYBZOwYuvzCXrbEn
Y1TIRndOzkWJOKDKqyddX4bNhAj9LPbbvlOT7UHhb3IZUt73fv0FZo9Fh5pUV1Xj90L+7HH0IU1t
FOswW/s3cteYH1tcVan4BF4LwW0INYD9VJgexGlhK2eyeOnaM8tP63rMl/p1jkzRs8qBIOJe8tF8
qfAfnOY8ciz8TlyN95dONkDcGb/awTMIt9+6rr2vMXbo0qWWcTw4x9TnpIZHwrBzodz5JMuWl8A4
OBEkxPe64BXxxBwGuR/HfJCQavpDNq4RSyHZrM2uqZyW1br/nJzY0tPh9nFv928smLTatSuMqbhY
pRRnvgMeFZgw7LBCGDbMS+zSGFWipmtVGK86RAz111Bq03NBAc+5I7LUQai4Lr+XCv4ifSkUEbyI
e1RqKDSdYDp2O6UjQTuRL5KqBAj9aAlwF13vLsHJCR8Fg+pCI6s9CcMF+OhJUiWt8ooh9rjJSIfb
vDpmgyspoQghA9u5lIfJmxUHUiAg3QRH6hdcD5CRj9R+HO9rRu5D03wjR7VkPPjYhRy3txUnmhkn
1Y1LOx14IlgdsxnCowVoo+0sBHpGV1bk3pTzIl1UZnoJfLf8Avb2LxZFlTo8p0X3dHN+W2pPfR+H
5Aoz1RLDfa2QV0VvHfU2GS8zcihuCfDakoqWfkCLYgKbMqmswr9UAqxp5eDREkeKWvdQ4qlpUYmh
LjJybfea6pWHjPsf1R7WYqtGHQx+qvdYu7rRydkkuYGfrVVv/W9nd/HDfN37+KnFtZS3YNIYllks
6ou12bQ8uwYLCpUcm/hCAOB3YHNR0N2ANvCmN8q2tjV8FdS2ICYTsZOMhgxUwAY2QxhS00iU7uoO
UKiMSq50tSArpiJT+Dr0X4xfhoLvFhm3VPR6tUoASNHL9lJMqHJUoFAi3slvn21TOPLGioSclDLc
UcTLF+KUDtnuxuMwEa8Ytm6HQbeREXF9/DVUuUYZlWXhx3l03X8TRD6SFpl9dO3rY1k0sPMyiWjL
2FHfRbjveQfbLFXT9dttGGkOxW1VRZ8+ROwwDRm4NjUBOYcoG785P+qpAGtf56F6P92L50S0x1x2
+yXyFU7NluHE9v28g6KpWIYoKWiVa6QdsufxKDRqwiOJZkJM5Eltls8zTrB+1ZyGway/3lvqHkv0
5WVL6ZcOs38nvTFzCGFELugEvN+wqWEtqU/HMCsPdDZCkU2Y6sleJp0mJxK7MIT5fijYKhiw8D7l
ecWMjsRN+MuTUuW5K9swCb5tCIci58w/uupb7Pnd3KnCTns9K8PJOkv/id3SFlE4zQS438foeXMY
9m4w94py5nJkFMUTRLumL1kORDeAb9c+NORJWia6746uQfqhFOyx+igocmyNa4OUcBFleX8xC2Xt
s+yz7EvnMQtYTQk5VxMTXvhSkXSm6dHBbn16t7pJonpGIycWVJInq5HY3pzgoSlf7o9xnN9p4kyp
VPTbhQvoTSXOqRX4UcW7AqrCs0oxZ5kWH8SIjFCpPYA8yYC1n6OUpHrYuK36fHOuSyAXnS2GlhU4
aml0es4x0/CcUwewjg1xP1EZew1nK9Fqho80IRclrzV8uu+lvFFygoAuFQeyk2YPLi6io3hXLs5t
dO/Y+/QGIGlOqQKRtYCUXytXccd9xPX27KeStJcS2XUz8iRri8DKvhZ/XPlN5r9RRCHlyqKzlqHS
FQECUAo9zino+ErhjAMH1hoJgnnKnJbJn6d5+Z4ZcwqhbhKUGdDztbiL8wATj6lmD9S1fWxwAEdL
Uc6bJHew71t1HGlVfPef2qP/huxF2TX8HSpZiecv65XyWDiC2zzoY3fx4pcvyL694iFcrC/KRQWe
60S45ZvaURnjsZbP3RBu/nGoumMSthVOeYQoLsRDzDQUT44yseQf4MX+oJd4cPleoh5FienFGKA4
Xrk9I7EDc5qDxh9sqk84UKjg164xUZEmj8Radoi+kDlIBMbO5VOrBMJ97gfynGa9yfVXstztLeFF
VLfWyI1oUR6drfQvJU3zzBQbCN/Upo8CMV8WkfhSO5UW/mBEmDbHAsU4XDpaOSJymyzQDa3eJ52Q
1oB6CLY5ICeBhbix6zjjjJNE6fV5BouYQDxrUabojIU2Lj8rXmVqRIRvjhsXYNxUrtHE9ErDg2Wl
Ovx2wdO7bMzsQ10ZZvci+fY1vNJwGbNgUT+QIv+Hl3/AKNoAOEk/OQXLgbpkKhRs2pML2hLbBd3/
DT/P2DnYTws3xgLSKPtS/eMDgdG4yY+5lSngMTnOwyPlUwOiUvRk4VT74QlKJiK2Q7cNjbiUBks+
wY4P95rlTOeFmrWNEBlLOTlBOeK/kvrJJ0ob/N5TGkWD22m5VWQhQLOWSludqkmQzIaOmC3NFADA
H46LTZiYkOCEOdBGRjpbigU4B117jf00mDvZvRJEahsZXlJdeLGgk3IxjQx9i5fzwil5MsmSEyeg
gWmh8ZoSZT7UOZpXUTqSPL0/dgynFRngDdoESGpGdXLhxAjCw1XGhqW4bJG2XI/dYejeBIFOeGaF
QbpO1OlwaER91xerXLp6idJ5EPYUsokIqr9xOJAGBa2u4x63+2iGK70pFyIt3iE7okKi1L/3KZce
9ROQnyENm35J4JjnrBNXR7G+5vVFTADfmt11z7I1BVYFevrODNgW4VOXzIB+jcPw8l56F11aB7XW
D1Q+FSpapVKcdLPvn9Md2hhrcP7u7k3fwQx/8U4ZS8g9qJjBq23sPtciEMNa4kgHItrvJEh2JW3H
7jE/pGUUyEGHBvlScDGqx/IpiJrD7j//HOHMQZ0FFqLi1+/X9Wba4QIu4hZp1bBSKHdAtq7mdg9y
8ZMRLc0YopL+UAe2E/UQUy+5bXyu6qg0PfyirLuifJB3vJDrbO303glyYRJufzeXKe1UQtvjzVWu
HJ6WMz4wIGw+gckMRHwV6RKrOnxdnoWYI7DfSv0+1xV2wn89JR6Ha/9zDTvb5gGAsiCrl4qwCN+W
YVT1GYbverwMbRiIA308KFpvR05ZPUYtzDFuVHuX8IBV6Z2nFU/lLLeWZXhCI/QdL4FRDrDD4XB4
w1jCtOFNr1y7XvKTkKky0/tzb/tIbOPWRCfEEdkMqjnSvkaLH4QkBsrlyJB8ognM8CVzlUjuCOvO
RFy5hdQNCsp5H6qcHFzyqk0GDkPFZsczrsyMIfT6iJ5IvkiKjMNh06f25ghwFEsY/4oaTylZSEst
XFILxAtgugLTd7x+kIc3ZC2LifAGQAWEEwrZdeKED21Ux+tHLhJddGZol7866knzyIAYq5lmsO7x
Av3Tnr1HnfHMv4CGiwYE+vBfvoSe9OANPe8/c7p5Ao1KCbTGVjCZIaDkeObOfJxLo0SkNJMUW0UC
a5uTyso+sUngyhLcaFR0hOji29yQF46rS0BZSvlk831ZSYCFZakS3pdGRZxI4pOQyeFAyWfrc/79
hsVs+1JDrJ31cNMYWtk60U0Boyc71z76uWv3QrKCiyR9mJU6AQ6SGqtuaTEEVKo4Y5ld/+Ul1x9R
DM9cFzr0u7vpkxo5+QigArRKPrjlZHk3KBqOWj7O5MTAV8y1e00PTC+vTkwSR583PAhzxqUAogKu
4nmSTFvh7r3x9A5ZBU3Dz+KEsigO+v2UBUESu8xxHKAY/gqltLqIihMkKBEkz4FzSuMzTDVRvaaP
qbp3VbAkFRldMb6KmKxQ3MOGYcAmJaG6JXjtDP6PTAi39LMQfgg+B4pMOC3en9qQREhgg06kcPPJ
gN6Tb2ZOfWKP+KjZli4y3QSsFoQsiXNA+yjv+rWiUoN/rKN6ycCZEGgfzLmU/zjyBr6Z6du1q6OJ
E/c7Z58qazgoi9neX5YJawZvNKqiq0iwK6fqZ2+4hEDktzH0pBEwm75yyDwu8ZFMKCXPzeQQwmND
CCxRhxbqFuneGrLQvQlWvHovYfeNFbCMCCknTeecE2ppf83EF3gXl32setZh4v6cGxvMSwVFEQFp
vb7SKS+UNCisE/eGzGcaTubBtEvN4Plu9X/Az3Wkl1uMtzmAQSopX+oPDu5ateeHvQsQSSXyNLd5
Zoz7+iFO4vE4XkxnJAv4hsGBloyGBuTAVTTTl1y0LPDurMknCbrd7VJj+ioiL+NkdMGklB5y4h+1
Nl0xnz/jJ/GaLKBFbeuS1ivRhcbP4Ww9NFJADC5rQa6/82P/KuylIxVep27Z5/XMSzuryujmRzR4
GK+dxOp61EB9Dv0rF9q3+gII2wYQVQffw0Y84Lz+SRnk8fuuCWEeSInzz/EOLrMOzOlPuLCZn5Fm
fhFGruuSGa42GqPLaMtuNGhFZpOgH9KDRyRe8AbwkF39ta5R3+SPgR0pbO4WYKSjUz0m7XeJRz2v
kNJTXRqsb1nMtTsji2+2PYYPZL7fjP5BfPxI6OKlsn+tGzMRHpX6nl6+Sb4lQKKDaGwoWgJ0X1Qx
y1oP7+7kfgbNRa4/vqqKMB+ZCsiV+bj6b3yDYcMKa0GYpsEsvhVmjp4pel9imT0yOTvHTDIU/xPN
s4Ur7NDAF6WPwCgYf8r9cXsgj+p+iWeFZNBI3B3ePx6GSJEOjOhiTBHi/ljoI6Q5V3akKMxgWrLi
p1otizJCrB0k9MyMSLE68T6+0ysj9u8zl/xzuILQZ38AbpU3DprI/1cXWHgvmj91ThapmC0Xp9ch
DmnV6MLEPjnfKQgTT118L+PFWXKEhA3Zi8Kueew2EEukhTbAdOmaOhEaEXUR5hbeWnBDjfgmEkFB
u8isShXhh+KIYyBfxuWmYGLhwpr7JGs6mwwsxgjjzz3eyooMUljaSyj3ELIlWkveYsUSwcQwD9CT
wkh8DEQhHWEF51wri4ehPWg9Q9NEVLFc3Yy4o3aVJQxtBBPhYDs2I/Mm6jJlhjLraDEJ1F2CVuSX
/Ni8tq976teNrdSvOLo1HKFuTC8eXpe27+veX5Cw6nYtPObSuT+MgFk16bWFYcxv9w3vc/yHTkKh
7Np/3D80MNlUo+DxMVJ0DPIQImxb5WlxKtcuRdA/dNaY+wQPOmkvoMbDJeZb94wA2uLgWuabPpyi
2WUsafOmUNIkjQbSM5vYbl9CpzP62E40bxkZFHmWrilyu7wQTilbyulU1UENEdAvgqMVUoQnfOEf
oDb6YCsTqb9QVsuKao+cgFlev4z7zJ1ryOb9k0SAC/5AIgXw+uhG7OGHi9dzeWF/GFXwSevf4wUS
gkez2BXQwuoI3whGzWrqEPrLyle4cP7dYsiYEw9sWazAWHBNKP+VUkri/YLVwjatgy4qstUGoOXe
OtbVmuO2JIYCPr2tKlWGdIz1gWzMlql2Z1nmFCGxynQwsypsZpryoKFZo+/nGseuSMP4OSRhGmjL
FpyY2Rv9cQn3Gn605YTffAGsuADQM0S9kMgLv0hMak3kxBEWevwYRWBeTLsUgPY/X7koH21XyrBm
0ucZWNFeB5vRGjTaQtzK1hBYxhWvdJ4G7L0+xBu1y2EOMHaC55trc8R2cRFMhWr5EQojpiI14kVd
zy2IcOxOaBW7zmuJxc8nKk68XUC2PqJuOb1TBAE0LpjcrtCROTz0jK6mtPL5V7Kxp/LjzEBcisj0
t1fweUbU3ekz5wl/oTt4V/UkWmK116zwMLkYGoWcI2sqJp6QcsAGT+5VIzt9ARTbuA+xxbpPN7mU
q+wsb7hX59YuCAxEPq1u97fA/CZa8F9SiUqsG6hbePNDq2ApfMoDmG1EslPUu2dkda4T7ORD8Mdw
xZJBXMKKQm9VUI+mB/hQ2rPdC+3GTAsq/UY1MSD2x6owLLS+pW76JO3/N9fdZhWgvLcUgv8aTgeA
7n4Xmud9jD7F2rVQ+Fou6P/vZdzRD0vtCFS+ZQTPJ8yXhXzEyNfN1cw1OEGxI1RqvddPMW35YP1B
JUR0cS7Vy4oMarvF9/1bxXYHmnzd0qdrvb5UP9yCHxMQV2DdZDIsuF0dwqn8ChpRcxhu2wUXQILX
Y8ua1boULff+yYSNzq7Gg1iY5EJVsBlNUN07Grn+v7fnAiISEy9jCsibOdIm2sUVKcdHJOP4qC5V
55RdGd3yFW1IDuuNMbNdWoYFF1ybNgv50deZr2Y5UTSK2rE5qSOdwc6Ti1pTpMv6kVtbGdztY7f1
kVC9tIlhXl+WgDbzfTO8LY4QnhynXXj3dZzBOCrCOmlbVoFWzx0Bo72O8PIO6zWuPAX1uyru1SHU
J85IN5PetImXTuTqnbIZfbgrUsmsKpHLIJl1XlGePwSZB6bsDhxJLzu0Q1XSwLFGmjXBR+jR3I+6
Xxr8upjoiaQr4awUoYvQ5ophU08IWoNpCvgBEj2Hik7nrNyhvEmt7HNcmykhf8IRKKkp2YlSuHT4
wsIVPQ4L6JdIMol5comfOmyds+tpu+WnyUM9/oGGsHJunl+Cwiwh6tiE1R7yzOS5MPsrQ116BuZ2
dUOtuyqg7z7u9dvavAmthDUyEJqhM+6vYfZwnS3EaEcup/KGmnlZWFMBKnMs9uIiGxXMmhnGepZF
WvmzwKUmKF/KUXOHGkRVE+nPZKjnNAEgQ65zi3gKzEG5JhYZNQxiUdIEx+DvM2B6vk+A2Yis0Osj
QUZG/QkhWPmeGYpoXboO81CKuWyDNT/16k1eNngkKEx4UVVi3qBa2l23EyerzezTSKShxFtHMUcV
mUrS0uwoZjHXHHewrD1lAsIIiSBNZX20VJtCyYmwbq7WvGdeFvEuF5ST0CSXGCWR/CdmnhhDo2Lt
jcSMlodjFF698apoi1sibaBnpRSHsZ1qKviP7Q9hhLbSCQxn7l+rD3+yhNG68hzbo5vDThf4vhvi
7/MXAONnvxkR57mpemWxp+COnUIqp6yOLm3GTGR1OPd9+ko8zt4QGxoX8oTYKBhM0gYWcNATown5
OkncSC0habHKuaKce3SfVQRVSWjSKpQnXfFpSYdjt9BsuY+a/VHnAn0/YxTGKXhXOEbcD+j8qXw6
mYcVsm6a0qvcX2k/zbHRfXpGg6JUHtp+YTyJkGqRK48CpBQl2i5fQtrThMac7f1ZdnKJYY8q3ZHH
d8PooNhuPU6D3XNb/8huPbTsbuxz4sw6Zvw0YpDRjSj1jZJOE4Y1GnYYGZNkqm4xJmy2qy9100Jz
x48MvqNk2Y/FWoDaPkeeh0P0YT6Xz/ycRqJRYQBBM2ET7gWm/QaGpC5ei1y0ovcDPmeAq1KEMbrr
35ca4nwaWKRm3+Y9AaAkAxK2rCNulld9x4p46HakWCD2raw/EFJYsWhyMkMVyfsRUgzBI77ul99H
OwU7qLOuhaKrvzAy+WF2afhiMK9XudptjOUwf1YaYe+Wx4kb+nh7YIX+9ts2BmnEQRBsrbfxcmDR
XOD4RupWLeIAGnXLd/53aw1Mzkh7A+aCZDx3vz0i6H9VTxT406EPjMLpXNj5ywZbB1D0EMo4soDM
ujzVRk9Kblh1fPCSpucEx69xeiuHKFMMJXy8DyTVdscxj12Uh0S7ezc1LAvZ3pEl5qV5Ms+Usl1c
Zy2HN5D+71EJnfwjlDF7TyLYbM0+3G51FkSebBL6wZAm2G/EYpcG+qKZ3GhbW4VFg+fXHFR0oT74
9AYWrrftJU0BB+gubWhnf2s++krW6XKi2MkAjNXuqTXhC9o/62l9FaLS8XwxJNqk25ajQ6JhLw4f
cbTm7yNk5ncBfNTy6DJCgIq7lxAzf0U3WeE5df1HdX/MxpbgZEzVWc3+kWTrnClFam7tPuBCpd8c
1OeWnzqpG/HzxhtGrfSem4EF/UdIgbdnBtKcrr4sOy56dc8vIv2TW7Q0aKtGSFq5waL7df/iuw83
EaJeJGYTOvsfrmoJJNucg5tGY+3O1EBCn1SD+PbX79K/Fwek+svE1JZUu0DA84w0bhgnLi4egE62
7HcNycffvZ//z7LHWzcbFgqdeb+OfOwb9EsZsCVKZQM2GIIOjyEErzYiR/vOjdRjsDDoEZn3u3n8
xi3ZB6Zzy880rsYnn5jO0S+3ReZ9zqnxJmHm/W5M2MLsAHmA0pmZiwydPhTphgSG96MdbxwNZu9z
qlBE3Ca5c3pRovW+or8RVY5C6p9LOXiHkZo28QyNzFeN9JGBF/Nlonl+GLT1CPZriPP6CtnKa8rZ
y1C3Hd2puPmBiC9Lu2nH7YLJicQtm++Ls5MnHY/0QPs9l9Omjhql15UeENeQGah/fauZUYmIl5AN
881XAsQ2hvQTHyss/tBPnMpz4CqA49ukbmEjtpuc1RpRbmQSeHMYwi3Eo4G0P5aRKbC7YQAoZFzY
ld1FqIg5t6V8dLyCdkMhnvA389opvL8xlrkoT+/86lk6Pj6v6UHFBI4MR6vEsZLf/6gmEFjy8mWr
iPoe2pbksCJiRj12dpuCQzqYo9JaBJlq0Y+kGFYpI5PlxIpdwJ42YcTu9wDjZOYltPmZkHdwcNeH
V63c5Xi2Nr753MgnHziXeY0ZXDfAuiRMD/pGzVUhCu/XszhSEpKxrkr6ouY8DFD3bWxZxfuEB5+L
ZfUM4oXlKVb7OOrAsPvDLQlxOQJyiikOHzrYeS/t5tbKcLsXrJOcp4JN+UQKshsAdJeuiJpy+CQY
0AFjvQgDbg3kLkwyx10vk87hCQQmJOAcGbEk1MKRfxUB4B6S5OvwdEZ2OEWLphhBIfEcnTMxiT20
rDnvB2m1mndMq8/6dymWk+oFWO1wfaUbXpGgrvAYWEHz5NNuw+5IKKX8SylNr5YcdJiV+xmatVPN
iC6xIrOjsXZy5yu0HPgBMc4d7r2Zcos6QhgqKtZhER1P2us99GnYzaUnVAiAq4OQKPcSLggHJv8t
SIab2N+N5BBdJmLh5mxuAKL0x3B6UGPWrl71mcvKYe35U8C+79EpG6T5WUPmnrlh+Qn1sNOki3Tq
muP4rl1pTeNaTScK9ah7ou7uMKh0DBuXO+Sloa7P4VOtt82C+2ztdHujVq1ZYBaxIkKSLB3AaqLG
Nt1NfWcuw9J9aDlVANuzMRb+MzYyhzmcqDoy+n0IJQe/3ALvMNOzDInb3YR9Rg3Bo6oljMEfYCzA
8FAUE+LZDz3HT7kUdJtgzwYwmzBgdBhxSEu85M11H1fo6rAVK50Ew1/KryraO1BNaSu9kvSrEiol
9YxMa08b6fS0iCmw8+fqY+uZNJcYeiPCD0hBBcRmhsFRubgHUmjkxYIeoGCGCjeONwC6n5IpQ1tg
VIeAtr65Z8aoa1GW2FeY7YqV8r7CGueh+1EcuV//mjgvXy0fsb/UUzESiM/8ksyT3k/PXGoJ5q4e
4H6zB2y19MU4FqEyrTc+WZiM/skucNMa39VguIhtz7ZkBfGNzV6wQIEClhlDkkhYXn/zlA3dSwxC
PJ9YIPo1z+qIHVz5Y2cF+2b5Dhr8vcAOt4vDO1GYPtrQBMfhTBY8FNM03vwIJ0Khh6hIJ9c1MjRt
Z8kFRxywGJcsUtzPEkVDjvmZQUBs4/U0bo9GMA+H+u/+JJ/anQDWgAAHpHICwMYHEQrEB0WPgkJf
qolIOBW7gbs47vnie0wKpEvsong2AIzuk/l/9r8AiWeDyY3gib15Sl3uwIxrOSb6UiThH1pgepzJ
pNz9j8hWRqtu7SNPCD/NNP25gg2xRIeHv5IFUVB2GevoiiW9FxRIm4nF1iUnNGH6PCQC1+BphXBg
bajUCBkmt3S4F8nWPt4Ut7GFfhcp85R1s+gtVNd+9GUqpoo0U1mzPg8mQp+IxQwV7aZy/1/ChAwX
1PHuPcZOmcum5lunS3i9k4RisISlnTbtTPvT09f79iUl2nYPeLEJPJsBX230Nt4tkEyhzx3XarqV
mJc1BLyiHf2nVjEU8mkjVbJjirGCM83W8l7Wje/V9+lq6aPxgDMnc9t3ho9mF7DE0ixgXGCyvS+V
dw9LQ4A3y2fbQ5892b5F0TUtKPn4IGLAGrVH+yp8411KkHl52Bu0XgvAzPvYmMNs7TO6GFzybv6j
rAjdhhiB+nXcH2Fgtv8uMjCEoW+GEhvlo5F035rSHtxfD6c/U7iGSmlF39goonIfFMLjYz9dlICX
Z4zRu7RC/9FpKi3eY2IBGDcUix+nH/EfjmoR+ETeklUetH2V+9bzOd89vtWiMhAXHZgV2tIEINbB
gTr1OBBBl42OJHPAJw/0O2KW/DV6JMrFlH5Usgr9/3cmcK0URP1DWsRZOPLxomTp9TOr77bYBLLt
T9JoBEAJsMm02fJqT4GrUvN9gXt1we+vyCMt3j7mAwoktzg06hpJ0dlpuZWEkV2pVIRRMVQInwOq
Fa1Ji1GerSyDoYYMu6bwnZSNwmpVTQzX0CqmbRqtI9NcmCNKks4D9DfILZT9idIcN1N/Z7gQnwV+
fgFHzEpXwoRPdZWH5J60ehgKrqIlLYlsGZjFLz1EVaAgOvF6BiAHlr2d4ADro1iididjEYT3MAgw
Pn5VadI3AxQTGy/KI8zvH8595bUu9ViRJTxLQrJUIwOfay9Tsl1WpwGsxnBor5oaCDXW/oNXWyOJ
++Kkp1UhzDYDm1/vLy0zCNligHoMe9cYx9f08y8AUvrFSuHth0PXWjjNJLqV6PFAEKMwcjKWUfpy
5XzgzHyZG1QX3OPe4QYbic0svkT7RzX8WrhR/v60CUU+Gj2AIlhp3wF+EbRd93XAfqn8irQKqA0X
nEbGvtYMO1S/iEaSzfV9/rj61ZqbfK8fFHI/9ys7lFMtsulQP9ImH2SUOacul7s4b3CK8RltR5IC
/pHXYTItrMQLVx7Lz5zx0QwqefFLe8DIpJK4Vx5VZbWxAVSj/DqJMlOXsJps/q0Prqctwd3gZkwh
Vtvcc8FywI2rDoH0w4mtvHGg6VKAUkdfMCu/ecOfxmupgTT1HVHmM9VqN3U5BSHn6LmiOi8ZIDLR
lX9HHOqJPh2E9cG6BM9JITJOYX/nRZQl7eRAT+8lO/GDup6WUTGcCvtmdreY3VU0zOzreRLLhXlY
04/FAA2KseSAum743vh54OYQDtHrPINSb1RW3/KVzXE+QNcQPHnSLMT/hHRs1ZvZGGK624J4J2if
myLXytWsbjuC8LXlNqwMV6WjCo9Xyk29boyPOavhQZFquQ9OAWZ2rGuALeCg2pOYFPDF+kdh72rn
fSetJf7AJPqeeie4Uu8D6nMws/PJoygtxSw8bwfXJMpoYAnLF6Is7FjRu0fStcuTCgDXdnQ9c06U
YOI7AcctYjdoqb3P/ELndfppxGLCR9yJYIxGrWh1gSNZX6FzfqkaOs1diCkhdwspu2T17E1EFEu8
yg1BWVZatbJab6FWUG4L7oLsj81sSp1aODN1jw5MhaEWWeFm9laDO2JvCpaSM62C+HVV9a0gxbBI
4iwLGV0sOzN5ysWJPuetyrgSYcfBUcuBxd7gIMPNrNV33Pzwtxea7bz29KNyNOMdxurvjE3q8CJk
ASmeqLwFG85V1o1IVdjOgRxEIez1LuSqAMFuuY+ntPOiwOOGnYA8lg3If7zultGrhWbiefH1Oh6z
YuenHPmItx8rZQg4d9nnGRyKV2M9nVCHoYds2tTsmTIVfQBgyR+d068XgDzc9BbINkD5n6TBz5X1
1BLWDfwHJEPK3hNYyVNGR5BJfGpqdoDI2V/BlH9tLFlaO3cL/b7DjgssPeUPgQkFu2QW+U+B/p4+
JqFSJHo2i4eeIzXmR0ZZHTTcmJQQPl2Xa/NgDPmOV6+nyeOuqT1DXVcslPGTwG5uGOcNNCmicBas
fGYxnniTnf4/DCka3Y4v09uz7wKXpW8TNk3M50td5OiMKzopaLZHVp4yMlzzOR8TdD8D8NJupOwe
ckF/VSj4QH7A7k8wbdLaPL0gZf/OiARW/Gg8eOn5vePdYQzxFjW7UXr9Jd29cLjtHvi6iZLg2f+J
Ko06c+OvVSv/mSpZcR3/ICCGEpz7uBS4bYjzhGlz9jGL7t7mxkfgn7tGVW0CSmKUOwF3rdZxhk0C
RpDFinZk9Egktfk6ZbATlg/WvgoQK2gFkL2xdfAORDjXqrC0bQVhfcSK3s8K41kb7lCr36izxXQH
W1zPgFSRpXpn2pG7YkvQlZwDfl7gpo1h0rfZ/41Gmoaiyph/PpCG0zxyqlz/Z9yeileENsRTClEy
9qGlW5JAvOupe7V9FLZgEyluUhcMgeslnPKIm0GkjgBFa+x82ohp1jVCyDteUAtMPfjW4TBgfeNx
QjN9jY30rMwZ9TUPta4T9VNVps50+Wpv/LKNlT7E+FHW9MEsXxiGwN7iTCggK0i1klKVyyGn+Gt2
IVoi96kCNq4TZhe0Dbsnqs9dl/BYCmnlcgPELpwiSDfaBpAMyqkjYI7fWKJpqjbNtN/sPNHYGrVy
7UWiK27yvgeddSeMpw5hFpsShxtsNLqSrnxpO6lyPoN4Ebr80QMBOskG2MnsBHpq1ikMisa7o10B
Q2BzoPWbzQR2FY+5wpBCz/8NASZJnzCBvl7kKcnfbDlBAG/lH+C67DUHTlTXMYzTtKf9AP0PSDKw
c2mNzDVv3eYrhEVOxgEbsEwTPHhiJDSvFci0gM0cH0yc9d7bXpwE998x+jYlQHCIVIvthj5xLDBp
tSLe3uom+nDDF2wDDp5tceFGVg/oUzNLkPzhjtavVT2JZF/AJtMmc8dDLn+5hLwUFaOgyOGhCCXi
neePr6++ww41TQbJW5WVgfO+LWnolJCWGBGWDn4rMD1D9Z9YceeP67gDBAHGVsZldaHNka9rOnbC
NCvZAcTVD/1fy31cvbZFBTjb2n6X2f/af3ADK8XFo7HfASwyLKwJ6Fdw9XvqOnIxy7YtyHmifEFe
kXmRU2S1wth+WM748WIqrpz00c6ZcXa0jh/4I2U8qFJKNtyqlKGowPBmdYnvrYiGPUlyo4MwI+2v
NxvbWd2EyuPh8RULYX4+8dOcJu9a+cp0xYN8WSetvkiBahn/pPrgwHdv08jIZ5VZF5z2hF8+iY/A
7WdL+X9S7o7RQBJra7wdNLaJSC+PHjSM6zmIdMao8D3lgttnCSJieRaA2rWyTWjYOBrLTfVE3F15
+++GTOO11lwLznfuXBK12c3Bp+0mJVjs2s9u6QxXkfNmOnWfnF1ftgAJaghCH54XTSvBZ0Eu4ggw
v8jjR4RMyDJS2TvdyGzEOH6gr34L6cEMdHm5cgw14JzuhtjXLnuoSuiLap5QLe43sIwWLF/q4PXa
xLVQFTcDAX6QSOxO1Tl1QDPA/Syfu42z7Xm9wVZtG44BbTpp/f+INg0WCr3b9+z/eW6UYJEYVeGb
luUqj/A3M0xSK4No2VBXQv7Dc6MS4OILjAKmUpBC2gYTqeI8QIQUFtl4Davu5vsaCi50Z8A0E9Zn
ZkgNxizmbrcOd8qqVcsnTF1NQrUmboWqjRvrnv8TXIETCFYtVJfd/4sdc+CCB2E/x1P287E3GQQJ
900YmsOGuBz5NQxVZpUuYFHiATmW6sRaHxy2F66bpYfq2ealZHUCEgtJy9dV8+7YWU3LFBpFlakF
ydwEOuKX3uh0TNMHKhuq/UR00pqcRhTuAgx+cNGUgPc6RbMP6h5DspdFxl+UYEDu1VZQ+AmuMWlc
m5yanvaRlDKkQik0mvt+rOedpNpqHVPykJee/R1leTM+NPve6+IyzyFpof7yPXA4wETvkIbFHTdD
yK6edWNexIygsJquk0UApODPzxB4c1vMJbsl602YXIlAo+Ua2KBpVXYn4C/NVM7SP7C1pW3m1/y7
xrSNQ+7tvfIdLBQR5QlaNDbqEep0KnVrI76XeJuWmhQQ9aMa2EnRwl7hf2AGhD/Y38FWZlFEyV/N
UQ8bPHpXxMSmqHifSgwmByJm/een4sAo8eZGajWhJc8ITr39SwOkiECjbTbVEOSE0PUUOpoZz1q4
PjeFO1hhuLNhGJVfrRWlotyZxRdBgrtiBYhVq7SMGg3zS8LtxEN0obZZ5ehqyuP6czPCZOYRXRTE
Qzr9t74ksJ57IejNSFn7qVTPAUKK5WTYu7YU0LF/tiRZn7gK1k1CPELvCxpRBoAtrwL3pO16o6Et
81Dkx+9q3XIl35dc3sg2MVqs5bSIhm8YPtWI8HbcbtIijglpvCdEw1JM76yd1k0e7TcfpGyCz4zV
Em38YBimFFlM/uvBytQKVvZjY5MSHvZacp++Y1DIpbduyRDgotQxm4q6k66lJaCw4HELeI8TZkcD
h6sKMEJNNTA/cXpzV8dNVu1eK76HxecBnqZHK0Zy6H9f8lrqj2QCTxfC+pTG0gEncY2Gv2MqBshT
ORuocfnM064k+Z8McdkRGuoT2KUo72ITk08Zwks4k9oiHfQbFJDJI8UgfILdjLemdhQqal9Xoi02
NR7MR7N60s8pT8F1kG05V2SyrCnp+JBZ6oFUyte+fX65qGnSC8dE9dl6WMdV9JOXgSWlBhsyv8+j
7QW/ptc2wvn9XWpFagdLMZ2gEV+qLa/AL5rcRqFvdQJOF68S1bRUmJXqGajdCy4jWtxuaORvdz7/
W7o24mUQE/2PxBmR+fE13if9WQb4pXyYHsuU+4pmb23av7fFDcsrGaSHNHSoxouA46QMTJsOhoPH
PeHKdJQSnfeWQRDNvWz2wlaX61jSwXd18uReguxXfaCTvDkogzA21yA8i7zs5UobAH31ulBmCneF
wznmg4PT6vtkemZS+N2xK0vMMkdhSba6t5skYWWbkf3WA+9oa0a4Yz56cuMjZmECDNBXh0RM5ZMK
lzAAHgpy6EVSVKaGIFcyOOT1vsxCYOWmGDhe4BvwJTQ7afNBfaIa96BJP+aimaF6URM8lTM1/3fz
VVhUOA5KasnSZ7dd9ujbWTj1S0kgZG8U/oUN8PLunHiZesDzJgnSyU5s49DfStcJD4gIvISHilI/
xCwq/cYDfGtW0Ky2IGV6WX/LGhnYjZSDBRlAtixF2BEeW3hRDHTQpCRXTt8TW6G8nq4K8cjB+Ibn
+r0DKwtFTYbwRZnzGoD2m2JSVFhM1AWmIjwILJo+5EVqzbtQODVmJAnOOrWCdXY3YpFsr6JXEX0F
PJ5N4rrv+3Kcv0nsEa2bD/x0KTVZp7R5eR2/GAPuvtjeIO9BnjtxkxYGyppP5Rew9+M5IMb5VzNj
1kUGj2nGobRLXtC8BZaqj/2ceh7XLDr4pYbW/vygnQFT6KF9j8WmNb+Lx10G9N/ly+teEnXXoOqn
mzcSSWLKmxg8AfNi+M7MWwflEZzLP213sjlZZ7JPmDhX4/GohDAYKBs6qvDz+nGnWrVtWP93T6PI
EQCcYFJAO76V3sAwPnmZacAs/QrxI17gFrOcI5ifz5zvYLSo3aRBsgHuLXgyN+V0f0rrkgrIf01i
ZW8W0z+nYuJZgE+MfvWIlWF3ONF7n5/P48tfWat1TUy59MFK1CUv48fjvwGiWfOV6dRf96gSxp1e
mfqHJ8ho1+00QcDLJUZV6Z9GK02C3p7QyTb/CvqAOf32YXGtA35jdY1Um3veDOh6NfZpRXxpDNod
QZjiDtu0+KQIm2KCep3JQT8xpq8HfNNkKU6AfAe0eZRHXy5xXvweKo+LGzYQkYNBCku3OQeaGdD+
R16gcZ4iccypFvPNQEP3Baj/L85xE9oG6NFDeEITXuZAKpDDdXULOlT0Ak2TZw02vVDrB4d4ujG7
JrEd6Kv2y4HMahLQ+4vStbRVvlCzSUTdGVSORfoiZXO7X+vdTIz9A3lISBPyURLVMg9WdFM3iyYS
+tBptV8ajWZAgRD0xhqzhOZeqNOVEiYB8Vw1iFOZ0+kSXEoEX2yEA2VfsnTqNdYg/dD6/igcJdRJ
5qIWiRoU616EH7e9flnd8jmcKhzEw9i7+aO/+DX0zDizdb2urow8Wo78E+CdYj1m9wdXmIzLal83
qbUkHFAxpP59xS5DG3DwxePIv1zbVrkgTnSJ3XnCCxNeKUhEGwybv7rvkjZ8cVQBvUpWR+IxpPv7
zqUxNZAyRjL5eZR8/I/owvD0PRI2huRXIxy+7oLBODjDBnVy325l+fxIilm9qOJXaWlVmTVfvSKo
RRQjZLZub+pC960lYL5KNHX/ZbO2oJepRHNh2TnlhDJ+BnrZIWKCvAI0uE/NaeWIJ2ZoFeE1geuV
FZTO5jmL0TUfsxGF0R7X4ZSSXgO8ktKlVHyALVHByJuaFC+wgIW1+DZLOQfgZ7rtaxbQRflRpryl
Q4IhMr5+z3JNw6WjDynuB4X/4zEuBpcRpKlxjNcijL4fj+8sayUJj+mE5/QI3EOoJAImY5tY2xiV
6WfcGJk7ZNIQU+yHUbTJq8vjOchzyG1B96yj1al1SCytLK9zpj5idfDfxzdR0MhlLGXjfocH4v9i
9z+NFgp2ifAzeGu3Df8+DCd3XXY//JPl/tkognWWGcX8vSpfl8PSONhPAGUhX9jO5lsJLEjVcI/b
LCJxJY2OYGzXxhWBkDfnpuSZcs4xI29rAQHogAVqwFa+u7dN4vL5k8wODWUg6FcKt0tzz/lBYkrX
MS04IMnhPrXp2Ejtmz8W/mYElVwCd1mQkiW8usbJ5x8njX6ug7RY70XRv7A/mlzX59yMdYFlEKhU
+r6fGKbtdoQcuhHJ8VcGiD0SOqY7M/uV3Yca7KlGgU7gGnGZXmWXjg3ypwKRlV1A3pHZeTUWH8jk
abfO3jbaUD9cI/3Snzcow2jk2RPj7GrUHhwKbpgL5V6dH83VGRVsISMpjhqFLzZzrX7ehUEdT2nZ
6eGFXairLI5xax457hAr1SKM4LFcLfZ2Q+fiNes/onfjl/VJoRvTXvWyw6b6hbDzkNh2LPSWdlPz
SKS1bo58/WoUq4q8cL5svN81+v3Lpzup/bRQj+J67obhVqIi/M0zPFDXgfjuq5HWIS3naA9VJVZc
WIvCQM+HVNkVEeGBeVFPG/E6+P4ZRZomEU02MEvIZYwpWbdy16+7Lz3vHPAHwBtrRYRmOkgYkfA/
8Tope9HW8AYk8Mgfd5Aa79+ctvq4deo0dt0jBu+KTznbcGTOolo1k8w+a5p80AvabuexCd+hPMPT
9EvxrsF70YE7JCWEwwzW1aunQ0tUQk7Fizg21O3kI+jLAQPUgHVpND7uLBnoigrXo084l+81sxMv
ay7RQnS6rtOHUzNlNrnamnyC5sjUssCQe2erx9CnZassExTaJzoq9CCznm0+DOCkyOHQVvlpGeAH
wrEMnQ8+lUsPxnHkZX7VDZxshcSBXweCt0mCdLZx6e5m21SFVkbOno2Qxa6wTjzgeT6ZOQAY0Iqt
RR0oj6QGKndwdLbO+pinC6ME4FaVNem1tXDtRHooHKoIlFJJX1sLXr3SSqtCvzHA1HxI0GIbWBhf
HuqEBapOSru2S4HtLEGZLIVsFmxLNeOXZEso+SSgADLBMCu4RBbeDSM+HMc9ch03RCmFpyQNiZ+p
JPsZI4xV16e1KFoICaMfTCei7nXtTomtvza+e4GBnIlnuPUehyJ31nFTPzESyTr+Uf+917RgWyNa
0OWXaY3t8WaN6G0tGEdN1nYsP8ee/8ZSsVhh9kG3NNoubd8htQ3Odt78KSm7YpC/27HVCmd/pQUU
4Z7vQRmsFJtEKvflLUSoUxTLoaZ/HgbxeK+u8Uf3uZymN6xdYlEt59dLmkE6nL3JI6V5jhoDnQKD
9KJRohdujc8lVvxr0x34s9r7nI5x8di2G5nwWE3wtn9Aw9iAvNhVQjiLBjIq6rRLStMhMOSbMQHD
1RdX3PvjHetHgkrfALoWjfmMg3gLvEYIj7g2hKnBJigXt7zyxKvjITjA3K9VM1+eRBlwHVwLtTx/
6RvdwRt9DGvMVhVH+MwMiTbo0YtR/ybFwpuug3YLMRG6mPF4r1QKIxdiZMQKjnJGqW/ippL4ZH77
8mggMQ3Bo9OymyhiuHHxBG1d3ttTtfGh4dOpC/YtiVhZeWqsqqTd6BvaxRwhnGatGeO0xGPKSJV1
3qPThIUsKZc6GuZH+StcJNus7Ak+DFjKtMzAKPz8AQPxEnTxbzOhw2dDfaQAguU21ZDHfOzbyXkb
xifMythaT1D79XJ6yJA+bP1Mp1KcEraSxS6lRslK8hgM1o1EseZWzOR6vK9ES760C7DSN18DMCUm
7er62EVzb6OPpy7gz3YK32RgueseKKU/Yrq+9XMT11YI2Ul14NEvstwYlqTJcvdsQwxZGq2ZZAYO
yxRd+6TUFqfsw28P2aF/jKNM0out/p5FhPj0iUNKywEMy9zHmY37RKefFFEpob/4Vba3JfS82udd
pCnttKnQrccn91zkPjdcMBgQ9pJC4ZR84CpV6B11rIS0dfPHmy1fcrcn3zOgMfOuGXX1meQ83iEa
WmARNudpHPaFwpLdUozjAaKE30t86qCO4ba2fV1qSSiZLP5BIAEKho20EE8/LDE0Fz1VEzsdou81
6Z6gyNYzO0tdEfRaIWNMMXaWphTY5prfFhf+3GT2VpzoZ3aic0fSCyvm/Vu/ahRc2qtFVbe5B0mz
5emyM2+y2+09220fro/7oQRn7R9VBDfu5JKs0za5U6/EZC2J5+8YDyeJyion8AGTTbQ/a6RfJWGc
zhBS57fzc6FRoZh7aLgsvCZIFywrueXHNGWCle/BCx9vv8mFTVK+lVd3n9Mf9JR/QMb8+5/2OaVZ
pjPKWT3aKcXKBmuBcqQlcDtyUC7XYTqHwW9u8gunAF0p6zGD4+M/bGFFj40rnZwFkdIB2NCxycPA
KvmRnIFS99bZx97UU/CLO2ZnlnpPhr1a+9bugm/83GpiVtXX0Q2sqBoTblqLFA0tC7aRv2Xkq/lS
yWmOlM4AQN7RqmYef1xd7/gVMEaju2FCOFN/STfjMTMajw084QgYtwiyGDmazbQYgFflcExSdKtN
cW2jY2g8L/R8ItuEnsWebN4lvrnkfgeeZWvBGmx6ieRdo9Ar9XmTLjsyQw5YrDNKDopSSAX/8h8E
fjPKXs/1JuQOyNdR10KrAIDwUtsAyYm4/dN4hX+iLeennJvRt/o0mvCSk5X+VXfhSYe87X8QMOa6
v3264cuSlucUefAFNcgHgmGETtttWNKIjIFidzuNRgdmJuudUgrCmQHPOnvAL3vimMGmx7kNBza9
BBKaU2y9lEp/SguIZvtcrYhJzC+8FrnsNFCjozq+Ozf0SZm45poCsE2HHbVjv3/mSMmeXtYrncyx
acTaQ7Rok1WuRFwngVSxsAC02VyT4tu3Jd9Ofdk81Qc2wtDJ5G7TcmUY+5jx2yWWBm2WjClZDY5B
o3DhnIa+ev++GUSh8HudhuZgkfdUXGjvhbSNV/ASmubXEhtnyyYFJLqy5urhe/rivlX1K4nDAbNX
mthx0uJ6+GZOyPdZUytQef7MEnK3gAOnNPKOvpRVzme2/mD/K3+wAj41t7xQMt2v8HfG122C/994
2WaBueBbh5qK0o5RgRhG/Wiak/HejBfJdLylfpvmd/WOmQmmch+XUZ7eUsRFJ4hyyX0f2047qeF1
Ou/EmNo6ifRzTPubQK8FshQv6faWL0Aq2tGRCUCBSX0jOuU0GjI5JSi0t3FRA3oRDu3BdZLAclvF
jDx77fpUZwwKs933Xa/q+pLJlouR46G0yj/Gf7xK4OTdAj6TnntmBFP8+MTL+DQVFcoQtbA/6E6d
C67pNvmq26VHQSLTAEHLIYueh1+iHS1fWyRibsHS15lLWYY1Wr8kpUGMqVigjUiYoiHMP4rAcpYk
Ckxr53T3k2rKsFCpWosJ9SMjeCWqkhkFnda1FRL1J77ZBryBF8MdRap8LRtuPh8el8gQcaAeJLx9
3RZVz2Qjvtul9jvhn1JGfTtx6rYGGpFOaPw4k1KqrTN4/HM4dG1AsFZWpfBB0naZ+sLLfvqp1gRs
qFp7Fq+mMKi7fIWvAgl7+A+YjvzGQ6luczSAtve9GBOKmyDErm3LtZ8dsfCQ56k0aTF8upEW+ZzR
djHz92xzC65P2yYl4IW/MJX7TnrYnKsMZB/++wQ1BFFC+Z3G2dDFZPn1FN/X2wyA+gSgTgLBJB1z
+hJ7yE74WZulAMAJWYzmkcCYEtt9r78kIxLQTqgDAZhr9weAqlELkG4godo6R7cyhwMVbB4BYtw9
Uy4D2FmB7H0NB3GGhNPPcqaadI2rPPX0OZTpkPOYCVbc9d9/WVb1mt0Er6L9mKunIMUfxnVnR110
sFSBwDzMqscUKrHWXH1z0uBT9LXvt559ZmouRAspgzY3aqvxjONtHA3xjUsOyTvZs1YUOKq3lHBQ
vLpp82g6BL8UHSElbQ/Z+9kMk3ynROSpsR0Fhqb51aHVBUTD6c6y/yxrmMnf4TQOi5sXItcwEURI
N8rni1YZZ+kLdwEhtNhy8s1PKDpv9AYII8aJzO2ezW1UDagQtlcXVK1V25H1u9iG/cZ2UCbABceU
PUx9gfeBYwECibJfrEB4GSWAQFQMMWJjQhNi7xlPvYraIbVyI1M5OY6hQ2fkFygM+HiGxa729B32
FXpjyoE1k1DZlzXH+VpPDAmrJ+k2HfaQVn/d29rxyTEHVGSJQwcpz2Qm3eCU/qtRS4zmUjMHAkTS
zAsY1HV8PAiksTxlMR2VFKX856pOwrgtISFMCWc5xcSEc3CMd+1UU1nwO+/EIEHPzW4bOnA4QAIM
HtJ/ZzV++CDYbhdKoscoyLdviA+2btP7vexVAcP2lsE+TFgSe85vEHFepg+JTQlPOa5F/PqIL8uh
1+AsjqxIhFZbg/FDPowjxuOYcijpVkXDJj28n3G7EkW3ib75eit0/uSZl4A055rqFyqj1uCi96V5
SMip81yS+dCOP219WIThogUetqYvjpo7zZScv77BGlCyNSn2MFgrryMlWhdr4qYYkD1XdqlF7IIs
qmrqgyM2m12cACASgAb3oNzXETa6YQEnhNApFsGo3rIkuRrAIxFCnULbv253ErelcabVXhDNvfR/
vIbwbVFYyopc1jUOIAN4gTETU4KSxHTbXzSbxB21jr+T/aSLqmMO3LkSzRXsrYQraPAHKSPt5vZs
V6H868deuHMO6oWZrP/ke9ZsJ1+6Wa/obAEBOKk7KU8al0TQQZDVlbI5j33dLSNUgcSsDB8ty+qi
n04+Hlb6g2JzTNmPubMrWNzsE2CudYEfPxmdOeRWCdB0gOR8HCxxDHaetSYozEdxvKK1jXzIhnLU
Rrxj1hAO1xcGmRh1shBWUG3l55AlCH7B1yI0VC4CV8CgskBEAKrE/HyJC1FBmlwHJ6kmjiO+af79
4lxkxsfKg6UDZU9JDotWouLdg8mUNeUPxGBgf/bB5ulfhqZXtAzLArtqfp8CnpmELOFPa9cEjZQg
5crylDyMSQuZg7NK16NnDlVKwZ9xMMNlZZJY3IuqRZ/57Yz6EQt3Yc6JUw3c/17dPCm2OyoUJGRy
R5mLuPf8+JZS52Du/K4kcPx6+wXhsBgRsXB3X6wQ6hPJVFyxeITKpqOAUxySW6xesGuycNcu8pFW
i0fexr+5r+UPDfOmnkbXjRBXlZqRaFmMr6cZ+6/Hn/zQnEGamb1TUcuydtEoShVc7R61VHijKXtZ
0zL3Gms/OoQ380MlNh4DLRt/z4C4+RfaFRUm1FVALqUptnmz1meBQaAujs4miEOjka+Em2r0lmh4
jTyYrHyE9Q6JlFJJH95HwPEP8jVCjuPMsXGOPhML2G1vLND9cw6UYk+RMAHKgIUfLWaC+hCrPLLh
uZiV5JTpPbcBsurjUkWEXUQ/ux/Nv5LdrNENQ/1J8bnOyD8R9f8QrWgWnUyC0BvmydMfSn5DXlis
5k5xioGdT3+WE4KXuhreAgONodh1WjJj9PGDvIp/0p2QIukHn7vyM7KIZxUwAbPqIvTh6d9T8XBp
l9fd7SViR++4x5Vf+uK60t/WFiCKfmnEYCe5AqXC6BWAHO2wYpkf2uV6VufMO7+SPthmtdWdp5Iw
6WUz0OTXfL52ZWcS/4NEzxWi35NMVYfI3dqDVVezWEU+C8g0+TcOm64rt8l+GZkcISRJru2q+OCl
JTtD2NrLvmZyQ8kkrYy4oT7+ox3tFYOCg5jJpwXjoeqdgYX/MuyleC2KBlLHjmDRiPoZ0GzN46HI
iTq5ACiOL2AK5WGj1NtGNPUjtwlOsu69FOc1RI1wi0YVqBwU1li3KgH4TDlTXOuPVEJkuXxrOhSM
7gs3FTw84GbMHBiSuVXMWfMD9uiuUvZL1GJo0tAjkXm7RvJ/ovHNnqAiD2kmcTfA5H4mwMYBajsW
AKGbbD/PyDUDcJ4GREwHXbG/ewTho+Gll042eCueWrEcBuNx5cTLx2VcjkISyF0UWVQwyVTveSli
X/AJyqIPMQUbWDotEqfLxdOQ9TcM7OMWgjEEFiNvC7PDXaxZ0nVfNVyGI7bacJT4ugOGGwZZxjDz
XKOSvNlTdFmy6qW82zvfb3fZ4ESxDqOrEa3XWqdRaTkRR2Hnp2LNzUDxBw88d8JAyC5JKZaSog0I
Nd3EGrcFN+MVd/NjSlMb3wzUpWlUow6CPvyfXlGKup3aO35xbisZWha4PB1bJLOuEqe9FIh1tdXE
laZR7ZbYrLF0ZXM3LmOyuB36RVw+dLuqg0i7/EOH73dk8hPbNRLMrc/Aabopluavsw//SV2e6Utq
0RikNfzRpBdkLsJvpgCSwuYXGz0rNWvYhDwg7zn/NOtIz7Y+FjIVSlrAEla/bn32fSSDTiDILNMB
7rK7BzZbUYDtKwyEMp5v3B/SStRxNJ0rolFwf9CXpuv7dQRl52kOuIB0+Or6sftmFDmv+zCj4cox
axl2RdFL/sK8I3Vvci/qFxnSMdnEqeZB01RIba5NsdSzgBZlri9APy1fVeqpTJVY2s/jlIxgF4x5
wx0cpohBChyfyfv8ASug/RxyydXWU0Nw44WZIVydxiXdwIX0lMw2OOWMwl11TInK2BVw+GQpbtWb
n+xCo1p21B8h/FO5MeuM0oDa5UxtPT7tteU4xYAMIzJ52taaF5Z50O3FEFt5cIC2zw3EUyiKygCc
HAGPSo1SgcPhqmFYr7HGuzdpG9A/2iUNIsn3IP6+pUepF+iWWxR3wOOe09Lu93VvNhQEElq8VbLY
4MwnGQTduGD3VZOiiYyg6RxSb8K6SbuQRcRYZvaZzJPvmEih1LzevRjX0iUSPirwuMudD0sKYvGI
rLUxe64qYojGbX765vl5Awl+lhTDnWqGkL9T4a2oDPHEQQ/5m+LRRodSm4r2GxMPktoglyw79qZk
PlegPlWLoCZUvANngwyDw8fLHE9edDUlel69qYhuNSZo4g1niedO4FO0w0qLOl1a52axiDQHp8Ao
UosR1zIu+VlRpGdSGreraCi2bCpIMCJOCGkbNUe9ywr0OkIrF2zfmjV4HJQfLhg0urpFIFj1VUxH
k91oaDOz6YrBsz4ONdsaX2uso+6+eqFoppKeejiSnDPKA7F3oFid1XIcEHNu93DJExVs3noBXMfM
J8gHbqqkSM02Jzf99BuGuMdnKL1Swj+9fFnyz6XU8lhpnnxxoToV3Sdx18AWXlGpHP29+ZI78nUU
u0x4YLp6KnOz3haDymPwpxKmmas9onZBZzs1TedAlxV2FJqAqV92lFXI/JSDtJ3edDNK6v+p6BV7
waCXRi/g3PX/c4DvircFmK99qp3pBkhVEPikeu7AHo6qnka9hEYWBJSWBVZSshn7B16SxNH7KkST
pQGyCgBQrQhjuvJjxwhItzJAWkxszsvK+deWgxKoSUQCKHEqXgEvEHFgVI2rtY7wvHVDpOtL4pyl
pKYYCNtT0411v41QwIZCt9p8PjoIiMe0BD8mxWKk2Z5efJNdLt5x2YOVDRHDqjbCCB2KxFRLgZHt
1+POwY0KPoEXIPcGMRaAw5HbovlZfLnwomYFRUYNwi+vxX11Zd6PCGijOOjVkE25B+Pj1WkzDhRB
foYs7rmpyeS5vKJwRrzp4ESMRpzVI57hyTf6NMOtVFIGNH/lMqxtoXnX3d94zTI7rpfjK9Lmqhk3
wDn5G5+T7eiNXE10boYhBsctnQx4f4Awqj3EDAyw9Ev9JKzGj+nRPWJyvayUCqM8KwWeKeo2fnQj
RrQBkDPElrDA/zGjGsW5WliRPYgYwTak+KpJbtQi+RmkCy+MM6g6AoL5S3DxToVDv65xbu+KbGTn
eE2JtVzstMsdUo3EeLBTZOLYao2mkLKTloGkZlZC95MeC+/uWzINd8s6FJc3E/j2oKDnKJH0NkZc
+/w/bIULZPs0qbWY6C/fUKa8A1sTHbmaYPH1N39yfTzHirbjDuSdljIPziu51mQ/ypx6OOS9rd4E
wzz75muAWvZJyPVn+msqCW/csv5RRUOi+GA28vjnaJAXP0KJ4LD1lpqiZSBcG94w1YwvdMBWYIqE
hNzZli43JHXDXTBfYyhBoqtRvCgQ0359FnTVHm+oAmWGQoQSgDiNwDwI/s5e4u3yCO9SonekUcl1
3tIsOIPD4gR94P7XNA+r2u+t1alFPYnS0Pn9un6o9otWz1miQ4OtWnXVYFmPj9DUnGbOAsjfKlin
rXhuoU6lxsviyUuQ1fLUgD3bsBSN2SoC8JyBrIO5R/KKAUk3PF6ukxFVY+7xitcnhObJZ6NpN3dH
fwO1CsdtpgPEPWtVu4KPCfU2ag0KR3C7a5QS+WVC+WflzxeY+vLkJAq8EjIp4vmwiTaJxwyCwWaM
rZIboBuYda7C0ZhxydUxvGJOQ4sV4xa2N5+evVz0/auMWacjVqu6g/5XOutOjYfu8qQD/PydN9NI
BCN/1OHOg3yu7gHefDdd66vY17oxn1nTQNt3AIfjsUwM8sYyLFb0JF6ej/blYfUoXcJ8b5cFkhGQ
WaL4vNDk3KliFsNRXO0iAVh0VCvwKcR6SX9dGnQOk8Ldmw+C3mvAMUJdQPuiR1zil9qN5woPuCzL
Lnl3MtjLclbwbtZtZ+5VV0UymZB04oknB2edRqI8YMsHfrT15/2Y+1db2x26S4b3gArKSzUlvKpk
S82GptTrxJ3S8NCaUJiO/zVqj+ueD7zZS4Fx9qun9Ys1xlJILZVzrGkYpQjdKWMTvJdqm2QDx1DE
7I9X5V9BBkadaMNpJUXWmdhrYGSvNhONiiHF+d21nAaC0AfTzZrjD6wXIFL+ZKcpoNGDuaKBr3A5
dogPdnC4/m2ZjREng9kJ4QLO9WkHUyOKtI0Em997tWflHu6JuUvxs1w0Vht9J2Lb4zHl93Tp67aN
dxUVzYgQE/lWEoT6GdOPtKcjEVPG45D4Xu+lQVjOskdikI2exKBe7R3yylebAvrh3Td5kW2ptEUp
hXMFZKtyeRt2tJLibB7NuwP6F3/Elx6sOYadt/7Z6nhIUC9QrXElF88JAfVKgBZlnL5nmxWort4r
7CX2OFm3umFqhHGtsk7UjZ3EUvgyw5OapCLF6CGh/IRHHOVPFxagH4CGaYQpPtUHnKH7InIxoKKJ
HTD0sVX8QsrpRYiZ/fnZJA2MCNxyf7OQMZmewg/J7IjZ1wstL65Xy0GVxt9DND2p46je4AnOBMVd
+mUB+MeB4gTsCjPqndJebo4sSJCvqt2t0o0j/GENuXgXJcPh8eq4twUEh/1Fr4T2CNiOKKnkGu2p
7SGjA+oig+WEQbqgzvR5GuiH9XHTYpEeuQYHd0kVlxMhMMSxbxACh/VSAeKzm9+CRigcxb5PzfHd
X2VU+XRCG3+DknkAc42dofdgvxlFatJUobj4ZTHIri0ReDaYXBJZWU2BaJL6pYhnS8V2ly/+pa5q
rLMAXl2269BWxWbgtg5AxIfk4YoGzpzqIcrY3AUvix89dxSD1BEyTDchUpZ6a+v4KCV7vN2i3iaq
KaNoDKw2Lay0lq6an49nyA3TjzA1fyUxHnUjf7AgXxIbsDzOFVdGvpBj3nnU3JyGdcoX4Dr33Zo3
zZW1aZS5r+NVcWe8cd8Md+s//4/FLL2yJpNpgJK22qPLRJ79Al4WTf2pRUkQZrZw9A63YVkSCm+L
bvmbytU2J1pEornWumgY2QPvwzeuVTAhv4XTIueK1lc4eQ8Cxpu/rRCxgxGXFKDtEbeQnG8iJvoI
p/bkwuuh1oDh/7/tLON7WJ2h4//jYIkWpXADEv8rRF3l6N2K5bUIzwfQLIZJnTC4FKvdSJdyGVQ5
KlAiZR2E/4IPCWY7MG9wOh7QHqyxBbVKBZTcU1XEJXvpcyoJCJeiAYqRZGJOitGEoYJHbyJ7m+xc
jVUNp7wl9jFetlZ8mbJEPJSwX1eQcxTUNK/keIm+OBGk1VZKxAUSQE5U1UTxPcaF+IjdzasLWSID
eUZhRm0OW7TnGgwB7ePYivnCDPPD+J5HfNt22XB92grQpPkS/DUTIupgKKNBNSyQypyYXt9YpSJi
d/aRK6DFI9N2PMs35YiEcCdxBDBQtN6Zpyn2A9IJud4mF2qqz71nfsQT8Mug1owR7vDOqo7purLd
W+4tklZPPiZL1qgkxU9q2LE77E6dsOy7F1Sz3kcLG5JDPLJsmOnLVY2IXFhznOUhZcegQmw5yw0i
yPldwq25vc8LxozGAdrpwKteyavSPWfaMC7DKt5MuUyrSonN6TcH0eyUV5y4ORfvp3XvvGYJkB88
WboeaUw/wgm30AU/wmmBRHxJYL9s7tLpypeFtN2I0yEu/vk9ED3DcnmaorEEDbaEvXDyNQOhbAHw
2re4KKQBLT0N7GORJemc1mz3mSzEb28jx9yAdCjMs4iO9X3eMEuVV/T2DZr/OEiyRvCELWJk1Czy
oKNnhfxNpJG2TQByifw4E/fQ+HUf6DDDhUsR3DaCwagn5awfVn+zOV/z/UQm7gS5aqXrea+GXenc
VBTVRG7bcUKYPQYbIuh76Kmx3uGuibh+pOSkWG1vUYj4YMeBXilH0pGjg6D8L+qOkUkAMJVeNIZd
S62ZnHRMDv45NDEjIIeHwL8bsZtIf9vfoU2WQ6/4gncJX61CKSIH6dbVen8wzblmlZy2JUaDNJXY
kKyNOuETBssDYiX4T2gwRSZSePYyXbo0QB0EEW2DuosKcdf2yZ6sWOuP4ZXUKTWEotjTH150Ybki
2Q49NnZSnJilB2akgbv4KRS5bvOvKDBrF7lC7BligKYDj2HsUixDMArR5FnVz1QEh1MK2T9H9OgX
uCEE6gMwQxrfUXq943x0hjqWrRKxDWlBl4fsgeTQu5u+7Ach248rQhprjmLUa4+rh/+emjwMss9A
B1lEJvWElV9Beu5sm4HErcsm+aIMU0RPnaomOpTNbRhcJbzDwJTI6FC8QFKDFnE46ZwifKfY1IPU
i30ZfJtdCaBdbGfzCFPeGruO4ksV3z2d1ap4NyggSMMKwEbe73gufqSnJxKwpcN/ZgbXiI5N1t03
6V+jGtIlIp4kSF49O+ZcC7ENAWkr5a5GHO3TCovPJdneRFlua+uOx0KC/cX7SsncdLO+JTaZah24
yQz5gCe3Vfvuk1h/W4GWcWEpBLZKJZHjW/3WUQbpgWZR9hCBs3WCCcgyUrjvEl3vhrxRSfJrdG4X
FTu3ypS6kIy3qNKMZY8FTcQlcgRZFsDvfSEvJKcf3+ItrkejnSyzJ3ns/yP2UIeA+Kqm8jjNa8In
3wfs4TROrscw6UMsoVtmv+yrSNX2n4w9bCMgSAtLcR+KjgmtQ8slSf5ni4BUkyF/E2Ee8YUCQTzz
/londJeVlPAg9Y5s407A0TLsTXuncerLcZo3ccZbq4q+Ux4g/pxiNY7Y4PSHMFVAjbx3t7Bj5mnA
qp1WJeTNyYAcGwaShH9ig31wYsJbztk0St1F5U4+HOE3HI98mBogkp4mTR18opjOcOt2tmJ+zr7M
4Q8JM0PQmF0obmePfZQCjMh9it56SVIa7x1Zal4rANUM0LTwAyV/0Bj5pZuxGnegChH2EmevfrXd
V1cWUd6O6PeEsyNQMys30Dp1RXP2WwU+dEwN1i6rN9rXfOCitcbXZbhOmtDX4XEE8unwfsuyI93L
Gezs3dJJ+maXaCYjkCVyeQ10EacN+QDe7mDpnFVq4jiHfAjsW9meTG6+jrBnI16jsMOoLeYZCfdp
OqZ3ZfOgzw84L3VtgrZXYKbwlszp6FYeON5jkVQ15LbW8gx+SkhS7WD8XTVRQR7O9qbKD+HuQFAH
/cmnFOkWD1R1PQ7cV1rkjBor1IRCy1WE0M5LsgLOedmFe0c6WcmIEypTbBXNlLV+VleRA6f8JQT9
9+Njgt+M4n04t8CSmjEOig/iq+hgv5agqOiCu+FMwYr73KjgvGNpETMV2Y8gbjZJ5HMovt+83/VV
dHr0ONUWeOKfw6t3UjdjQ3NhP85CgdR3ews5CGc50MHoXNnfN18E+1vaqdow2ZhNfKgD8xlzpEKO
ODMyQy4ZXDVAI7J+oKTfCOgUWsGQuODAbT5Nkr2dM5yc1jfaoj50GhPzp8zIT7AoRlrSsd050rM2
/O08cxvfOhhCrzZ8iyyjZyAEY+ad5E9e9XuNIXOPmlpmfPEG4kLcANrMTUPmPL5zE0tk9or4BxuM
jWBaqdFDyqbYuR/ID831fuujYl8j3SdI0wm6eQYE9WIKGI3ePJ212aImdnxHU/fIDEejqRj5Kios
fIZG7T+orbMMrDlSrYDnQO5RJ806pf+2Z/RTvrVarXSxKu6ff/l/3H0Ys46WvA5KUTgKm9jCgHPO
BdgN0ql0QbwNrzYWf78YVO4FR22C87l/wq3fG8M2Kxpf7b+vKCGZY70F6dJ9nHusf5yeED4ytPJ8
OQB975zPBjtQxVM8u5uokIbXJD+og6XKU5bXcrE2+h3HXby7S+Q2sEIMaxeToG0n2MO666YKEa/B
m5nRzjbzM9JISiZqHqZ3mIG8BpZGdxtr57fCtwynUfsrZtLILjH9cr9VM7OxrRfgdMO/maXAuSFZ
+MPTJjX3iHyOgqfBmUk3NWU9BJrr2UNTVj9aJe2GdnCsMSaJVE4ICPGidyNvtX5OpRkUrdJSgnH/
Y5gWs7esZAXYhwx4pq2+B4Z6CLXsk78g26Q90Uaof7Nu5fqqgxHI1GVUpmYIrM46Koxz4vqv1dsG
TimbgCJlI7Bf4UmGlgD81cYxw/+peSBP9VC3hMFpMJYlfkdeTf+APk6NhIdU8qp72f4nyQ32Gr9W
+gtZ9vZyKHHhImuLb9CJZ+yaLDq2Gw10ALnhv9p8+kmvJnZPHutPOxU0mmUKe6ayNaNHv/gSDLMD
L0es9ImkQsOLHD+egeUGjA2ZswoTo9E8jW1UvxerDQ0nu5USHSu2skgZNe7TlGEgCYfHlLfUnuAK
Z/drJatMdf0GEG03QDBloBFonBTVIRFKIMt6nr+9TNLae4ZYqfuRfSrTC4S70GkwYkxL+sdtUS0D
eap+zsRsfAjd5S4uq+pZXpoGl2v1K8nw8WAAoxBE3VmL+irbqBUz5RWbTxFcvydwADYfEf7Vb4dl
4YEipQ9kzRFsFtU9mUT8tWHuLD5AgZ12w77HVTAKkJbrq2UK+p6z1pWeYGC1j2/3bgI70qhnnsuA
MpdBIhCmJMe0QBtz5wB2Lr7gRXVvkNUFWFim/A15h//fUoELnuMnxQhaREZGtouifBy5WXfcdwWM
v56FdY3BmMIFqssV5GLWjyKstEJe1JpQ+uvogINLQubGm50GX26hNoV6SDmyePfF1QsjdIKj0bd9
y8p/ycMatOSueZlXeQz9Q/+1GuFl4G0awaq3i52Pp96/mloWAzB2HDd8ZfXWyFsmMy6vQxgjTHGN
jMULMYoIfauZ+K7fas/ujvg5/N6L/nhmYPBPMTrRzXJFcKgttQSrgC7U+lhhi8lpmn/84/YzwX9Y
GeXNC/+ldrryhhTrU662bH0efCMm3HnKsnJLynhFDvNRLCnV+29JLTI1TruBphruyBZYvI4YI70r
f8b39DH0L62zqvx+Cshk1zoUPd0I5+R0LAkNdl96CSx7/2NQP3y/UZJlyP8JLk/ki7jGW37EYeY7
kH9/2ki/NZMjDKKW8ZwN3LXrkIzGDwV9wi03edg95cvhk2SN5XWTholX4NMDpScOqNXnrQ3uuB/d
OeB90UrFmpQZYCvnvH2SvL27yQoFFbzfvYoojkmfLzWBCZfg8aS5Kha/L+7z9SkVF/x6MKhF13pL
b9R+h6UViGGmfSmkqSm9PwWpwpPSzqpXs32hnnUdfEayPOHbmtNV5LTzy1W17bBh9VmhSZNwMpx1
XmP5jp7/SD1sv+ChflJcbPylRSvpx8YH1cA8++tvj/MkfpSF8n7k4UdMJHnF+KGViuNUw3FD12/U
JRrbjDvea8EWMpGKZEhTWNSmW0a4+ZFqReiWGnF82z3inZCoFKwXnF2V0PvB5CUpYFFxBSV58ne2
Vl6BRsV4vkgOJN6vwBjPwba1nCDZ9p73+NQ6sxf4YlVcDtgndwy8CP+TY9+33QhLByUOqCC4mknp
iMMI3PKGyol9AmAs7MA1oqlrVqq7bPnxb7c2bw97Qt7QgZDfry0bXT99TB2yL/PAwOo8CaaiJWI7
+s+NqmWohGnVGVhXkzUOM7Jy58gwuJBLrpfPUBBv3zXHFmpiquwv6kcjB8+dTTHYSow9Uo5Tlby/
VFPzL0N/UfuHJ7SJlfHV/G0TeEG039RDjWv1FnB232umxlvDGodAfVM8SLZHhjfMcDAkSx3BYwin
EyLZGtFWMGaUkMkOTENap54RNYRkx6enFsY0sCW5AxuoNt0b2g1ow4H/Bqrd7qY3P+QCXNzMIIpA
Jf/vU1fiyH9hK07DdCy8+BBobFEwJ5POg+HH474+ixx2Ub3WuU8Md+/yKkJcd7iLroeCUsMhDh1/
q4a0IEkjAzO0m5QnKM85KlL/fbdXNFR+SwUbki4Hn0FWjv/4Evou4ELH89ip7uGT8cSz7pscwFhK
uHLOMM/HS1UstmJU1ZEEsR8UtgdJJUPoZB5XuxHIng5gAFTORLpNa5XlDV2yy3xxQBBpmvUgO+dO
LrsSgkRWL7onB2j0YX0/ira95Aml3cJWb6C8DAC2jWZYIEregXwRY+61X8mkS3RK6EYJOIvF5n+R
xEzURgDZN45ODN210zJLMtWkqu1t3h4kYXvBFU1pefqvYw5Jsq7RZWCwjQu+K3vl45jofkc/iijx
osZIqFMTbIXEk8QTHxpLDVrAXcASSy6sEh4iPggo/gF5SNnBdlfUYzc57ep81rlVkp26Nz4uGd64
2JJUim0A7lAnyHwMqKGwPc7EQEF7pzF43uhEGEQN1KglYbYfo+kxbdGI3oUicoRXY0y3akP5DBEC
UCMB4Ihu3c++S9e4wbDQyrBtkRuPJ5ZjFTvhjftZWMAhvp+SN8IW5iYMjn5fVXxOAyVTaIWqL4z2
o9VQHMLC2AZvr0QMhvrvg0BCPFuoMf+3wQFGVHOU0W31z8ds42GGLyE/z0VMl333yQbi4wDWSrtf
or+uuypE26OyXFrMzlRmHf3kYMPXSt3pR/dAaO4OqfK3jPGCcXw/nJ4Aney54sHUUp5bNGJoUrHE
E7nxeGBTQ1SJzQxIExKIwN3PHWYedpoayo6SNZtOPKnRYIJCc2ROB8v35v7JPuRrpbjFnIpsIxr+
yNPPSMirK3BcABSzNyuHp36C7i5agM5LrFKYN3XptWkZoBISda1Cqe6PBU3cbRHeOHbdP1++fLfX
Tr9j8Aoa4L/MSLjmkOaahYyHVO/+CojJMn9M4OEBAdZo64NVtvH0kpt1bufakMLepW+0kYqtOHWq
yVdi+N0xnRR2jr6Xy8MUfJtfADOZy6fV/PywAz87VGkXgakPqYm0HAv4GPXEf97nqD0qZwed23Gf
ETx+62TKKsmY3YOCg/YWBjDkt1Li7OlTaXFdXsjBg63qX9l9YvtD2/mGbguBqinwJ0Qe/s7xhJQj
Evqp5/yXF2I/k23mDr+QQ5Qlc8WBtaU/83IlMVA+b6nrkAaPix2XT+GTakikHGnBikhJVI1vBL97
AoqGPThUmD97d83anqO856AZ017zbgTXM6cYcbjV5MeqcUvZVArpQgawrOZZisN/oYSPWhnES3xe
FbiGb9T3MRIQQGGnvXu2o5PFhaCx06cgBa+0sIke9AQoiCmj1iOmV1zuBXkQQETFjgp8ZrzMJfUj
uK6Z1kHwbQzVb/KLRgVjbBe3sIGl2g66FNEiCfAVFI8mBXzK1FnhsqwXC4+nX1RSoci9VzjjItP3
MIgq7/weaTaFOJw+NKtmG78efzEDwlgngX35G/4x86oFoYPN5UA6C675jqFG6Amkfny6Izh8kxpv
nwaNF+ydJKw9a5kkM/YhKS1boBcTsz62acQWyk3wIo8HpYbT4nszxgBeHqyp+jVgVfY7x3Q2TnOS
KNT3PLDnfbLFK/jM71TdY/O1QaahxidR0LOQOc4qcihVpCqAFwMu8Ow25a2heJen2c5w8q5N/IO8
vrICXy9fn5knuq2fr6rAnR/KYx1iYqXqz8UiZgmma/vbJ0rRnR0Yix48KaczK2jlbwgrvjoMfbNf
cpZzLY73lRk/+EZFjPbhqqeny/3sPahGYpEQPeErzrOFAwUzbMzm8FhFHUbJse8zfXJCF9xG8myr
7OKpJrLgksco3pzaNrThB4Lk9T4WxiT7fhGmS6VvrrfSPSQuEve0FHvvJ6HgVsaGoNnuciIbQkXM
rgJiXk5r2IZbN28IL0x+B5NOQBOutSBaQjz8AkHLbrsnZ+cc6zc4LTxKwDn5GTpucAEkCogsc+pa
21UyGll0njxSE89nygZegTj9RPq3IirzHz50h4becP5Iwwi/EcAAk84oza4q9luM6toULPuS8DMy
Mx5eLCfNERIG2ZxyiXBaHPcKFRIbeOjcNDsYYmS58Jediv8nGFwiQhArpkbDgwm3B9pTQWrqEdYL
ch1nwM8CGVsCXV+z3rK6L2iLz1QCZsKz/4J7Y6pckQpqmzvCl2x/sczLONocYu28WbgxZeO40hOg
a/wdZVtZx7uako/Pg6Lex8u50jNOvUP/B5x5g8Wyb9eHygVz4abqfftw8bWSD0HNL4Of49dFlqzj
Q8S7RAveyc0oRgUpT00/oLlczN31dq1GbBILuVqWhNEDUzIT/MZQ8Kbd/8ez+qJpNNnMFe2s1bM6
YNZgzTc2Px83T92SHxNljQFBJVPG5347RE34c4SyO31qle5bF1pPtdNBLUYNs2yheB/UK7lhifWz
fUOksMcN5XVn2HCOVoUEA/xJdnfaSKjXRz+yYmF5T0okzl41fgP4h6NQFFHLx4fsoZ+DcdF5soFx
Qd464N6+5ZV1eNm8W8c8lnfKAhgLOyZCsfXRYU674uLeVxV0yCrBha73lebrB5f1gqtepfcOo2XC
8sWrCXAa3b3K2ujmjkdO/UlQlIAGOaHCmwEz6LQ8F8yfNPNywXuK8A+lusBpouLxF3e9CBI34yws
TCpgswh2T5AyLz3CJFmnYWyJhlz1/fx0bE5u7lhbpo9wE00xrqWN1eURNYDfFtXWbjkjdpaSIaBZ
qcY0xFoeEz4wNfi+eMHsheUQC5Kr3oXg8mo5smS09ua9eAMZeuzjkGBXXVTwDizLUJEV9xc4YGuy
N0TkE57fhdc1XSz4T6UA6lbYXNo00kLcctCzaa7icbS4YQBfhnQGD9URkmUn2hE1CFF2WD5dapa4
mHEHKgKoojB9J6sKpjZf1kZ79UOUxt3kJ8jPHTQhPOcYJSS7cqjrXu42qZlXLdPbMqjFCucI7X/7
+5v0RjvaSCFfXkYPZ10Pu/CLd+VMfbPv3WvoJGTp/dHYrfhgf4CUaQwu6pqUE50otwd5Re3SabPF
yGWZEPBHrdBTuUHJxcVNugf31usAutPvLwffV/pLogMjyO+bNUKOxjRDREy0hlsgwfhwsE3/cMkq
Flz7G6rHSHNIZgTPw45oBJIZoX3YMQB2sRzAFVjA4SLR+UdYh1jW3CM+zHgcm3ymKPM8Kpy94dea
JAFpX+Qk8OR84tZICiTu7gvtxEPM4DWUD+8tKlmx0TCIWEx53eXKgV88MVnJp2wZKaYEDpVsND05
vd33THTUedTmQj+3nF5MGLqxiKH0aaqvV7XCz1/S9Vf2R+OgJBsgdnHoAAdB8CwmxPN+5nK39+yh
8/TXcvRLFzHdt0xRx53LmE57SrTrev1X4iOdbYvR4t0nRyZMkg9clo35gGl4y7k5voCNGcbhz4f6
m0SN2LJo6DvJ/kIGoxJxayhnmkBuS5IM9nLpZteHAQdBCgtzVG6PCEFkCLFqfyNvRUaXe9Imvqhb
rAnQZjT5yUPESttX7hoalgLYpwBtkKCZuhwSmMA0tpJmcgKBYEqp397V9ltKVFrljqbl3CAZYCGS
EESJRbtnmmNcyk1y343LmEXcCMlyz8hV5/AswMn5flA+PH/ZT63lP5eFv/91g5vG+K4FXWsK0M8s
EZJ5S6yeCcaMLiZovZnU8shlvyjIK1zUAf5bQMtLADPEilCCGuHpNEC0W60qsSedqA2HqBuw2KRk
JvyGuInvl5AlLX8sPjOjKGCAyh72hc034rqMRFE4hzyJN2Y2VdaeFRFkzEZiiubQCoYD+SF2WyAS
Mw+CJCrW+yCAxc8uCzXNoMl9w3SyENXGGAN8uUFvXbMJJtaeqzRQpuJjScBS+tsBAunUk7RQkLGt
0Off8GbEVocT79A0aXQoQBiV3h2Dxf0gDhA7dvHNW1PoOQTlWJiRqHEyzH8EH3QzW6V19vZ8U+O0
0KsXZfuTDoBAR83wBTKHJf3kCWFCr9VBXAn7x/YBYccP6arS8HVp7syLjOwowZsn08LIkx5x0ydx
dB9xhf324BR7X9Ckg44i0wfio/rJd74NfowqnDqy941qF/pqVStDU2QVwXZ9fHYThBIZAuFzyqA4
XbunRTUVvYzbQrbXH71oDGLDMxaaL80/+6TwGl2fANe4EOgEztKIAAcXOA03AKG4TFn7KnJfgiwR
L1FqHH7JGf8b5dOpJWlfA/fQNSC/HRRoy9PlNd+qBOdq7urfayE9MH8kGeCYYfWsp3j0t0GRX6Ry
T8xwjW1uz7j5K2w2VHU8dmQ6WMghWa+5k3SgiFdgOxONkSW+NAAQoKJQ+K6YoP2d3Uph8LBS9Xyk
t98CUAtUCtQVIR9Tdgqn7PGNg0FvUoCxCOahKuFJlja2LuZFQQeNWi9qahJW+IkYU19EW+Pq+BTq
Eq5Pcg6dCtDdIPfmTM7qeKKkC6wm5MMtPah5WhsVZwajdaEwWJm+npciAaUtEfQfTG6TRwQEWI6i
E/Yz/WAfV85tTpRTCHkedd86uxlYqsJPW1gnFoHGvNpLMJuE2fYr2cC4zG6ZQF5nOwjUfpNircKZ
IMjI0l9TjUwRBw6YxF11WIXnGcn05g6tj558YsyZN0QWfdi0jF3MTmHBUvrSoPzTsBnkK/+jmC0C
qaNVTT0jMQOWnMSuPXP9dIkAoNMDCeUaNWzKzi7cu3E+a2OVUTbCNWkxtk2ERyIH9D3Di9TwFkZV
DUU9XN3PhAslXiywoZ3E7F+pZ3YraEqyA7iz6b+r8lXTCdOTMUqMLjrT1NpIp+e8CH7YO6I4b+aD
LdfVFJW3Hz1wrygEG31alWNnbInIia+us1eHdO15VAw7fSc8EMCnkeINdCLodqhn5JvQ7UCzfdrR
R2pFmYcPODQPpmf0y4Wbj6F2s+PwNOqZaH7/xP/PE6JW7R8mhn3io9bM4hycqd4oMRJaDMjDDyDl
kruL17OGwzQ+CN0BCHvZamjvVuZcuCbuLbu6z+B26pJ6CUmYULLhxA5+42KaUQPE22NqjOtldDaC
iokwZSZcP918w8FW+27xbAMZl9xWlMDvbOCwY/g+0czmoL2UMABIYKV5QSvODmfPbbJ1nwXxzbmf
sDiopsmBiMllWIFRaGUysLMzeSK1rV4Xu1IWqv8GYeI8RzOWWKsykUQGI5P1q/L/PgHog8RbWsWq
oiRHJuRn1kDGHOenhNuTsddj5H/S/Czlo36hxseSzJ8AJzjex11QxKWhMxpfa+SJ/ydiY+k3XKWg
Si8TnbGKt9zBWhuNs7iTksiQBizWU6ZPTLGc7IkGbSDJFQKd4U2+4hIrSDUJ8bsZw93XmHh4NWes
gUaE2zc29u3oBKmA3leCbRCjYdPLpIU5X2btfHogVELGFwrBLeUm0jl/dU8PSsQm0GQ9UMG3nfBf
NVXQKa2o1GN83WgdbX+Eti1QRVGSL3GSgbSW8rO/bUlulMKPPmpsEJhVh9HkhLSHcwPk+FBfvCT1
m3keQXGBe40h0kWm6PO8wYIeRxLq4U8u/7MfD1R8ToYvtXtnLLtZHy8I8MPtrLyjaGgjh8X+e+3z
aoIwdmPCPLYqBi5SS0Ib2DRdcN9DwoN0gygHL5D4WUmvyXPFRrrBXmEB2qsDZ5dVRMMOAcj1MkI/
1kL5NsPwkU+/79q1xSj3nBEsErdXUcEnWDD6UsqUnKdbMVrU41qT5K7MnGVvkqtlgtniqL+rW1c2
D1q0E63921nP3ZM/RiX4yQI0nGZlX+HcxHVR4ba3L0kSXlNDJZQIXVwdei0yZRfdx9o8XfyxMw6A
mpk5v++IGbFemJWYmxrYCau1/5SLBIGwhgTyLZKrZj0+Sj9cXGJOeyh3EdBzVYFE630OwS6XFIut
aCP2sxDFcpqzBUczX3dmUi9OaGk7Nfl+rqzOocF8vuOOO8roOXBdSnS3GIR5Hj8guC1E/w9dZAIY
dGuAfKDfRRgPG8I7BbVXV6NJqpbb60GcULQSaBdepKzdk6NU7TxU8haJMfTIcxHtKIRZN+HT5MGV
pU4DVVcIlXKSUIB1IrZwRzsIsupsOenGreA63eOVoobPkDCUQ5uoEy5SdqMuAcKOQPzWmdkAuOS2
WvLBA+5TQmGW3mI7Tbct9oSTzC0TR3yW1KIwhE219946X5tvZs9XUUM/A4qAzCkmxCSwd48T1bXq
/hqL6SeUsn9xYVhyDE66gEs0gQ85uZRcyf3snvf+5EJs3a4BqTINsqSQced/IRbNlEeQubOtwqEC
JyApkLMOhOMy6rht1M4AOO8qCutQDGa/K2seLmXyJvjbtVJYR0nGnWvdWutJDIB1/I87rmZowwVQ
Sf9k//n3hBIHsvjsjh8MIChzJLvpFY8tjT5ZNdfGcE5F/E+6+eSMRMYhUuZdqPsOQ0CrNdMUl4hQ
5e93EvNu5VPSITQVCFrlwJOi0OKryb/RUg75IaCt2sb7ap0ByYaJ0uGRahzCKz5auwexR36lwqnn
kT16eQDVpHHlub94nEUPxDWUmBlmpDLnlYBaJZfDwlFP1YxN6CJ2M2JGJVXUho/0tgqk75ayHwEZ
EsgmxBc95kYvl+AH+o1cre6h5F2aJ4TA/SJulhUdetCcy7wdIrnNDiOE3LShpWJ7cJagZ7LC0x97
NZX3NrOv9YkffBT2f/rGEwEgE6s5n2ezlfRMSkdm0hnfBSG1k0PnYcrkFKdSDon2F0z0pN1/VTmT
joa9CniLxhzjCTNnc1TB0HNXV/BaY/FrlcFPT5D/nMFDvYdDGPUO92XVR76D72VpGgPlLVsrO87m
//GwoF6+jcx7XfmITNsvRTiOp0A5rl05YdRgVSA5VEYzO8X4VAMEa5tAWjQilDomSBxkgjCPothO
WH33NdQrmpLIDqA4ofGHe2GxC86Bt7l9+PRefu19Ju953pdQNwWlAcVKgQlvVwGHvWGgtivxr6U0
qFq8IwrS3wPImECFPc24kG8ji9g6xjjk/GGYaG0SFwp6wOA3mTmWIkIcWvqSbZobXZshh6YuJfr6
S4l89KRcCEQIsEkJgLBra4a327ZS8DFAWiu+owdHCRE0oQICMMWtG0+v64sSz+00ue1xlB6GZEfk
btmoLN9rmGpoj8dAJM5zEIY+tQzpNXYXcFOGaSmG4SeiFr7g7m78Xip9izSxNIPEN5FhtUQmLy+P
y6/Dvt+G2YJGFSOVcWzsd1GL5Ic7xFWP8jy0R8kF4qYp2wXJkWR9nDm7c2vWGT3oEpGNDvqj3N02
N9Z0NDFpDwX28SEFqBcfcAGPQsc3i2TvBuP735Y2bwmBW1nODNRKOYgv36+sLRZtsP44Be+hH4vR
hI60jxGqs8eIymyqCw8eKq9C1JjA6qG1xIrEix97btkKDimhmnIkQUTEBa2iw0E57MiR4gbf+imu
RzlSXBwmCW/qA2G8fjj2VcRbfbe8DyIxlLnYAvxlw9XwdZTftJHoE9udYViySUDCxGe9BxTShtle
B4LD8sWvkpRyh++U+iFlOLhtJAMdHMxLAE4Vt/YqzeRRFbH1ULpkNNuPcQmxePumO/Ed8Adn9vBN
PRB8XjVkwBhhuo37FpKZvuDRhE9hnQUfG8iV2z5s6phxuBkk8gxZbSK44a3WkoyFfYAkD7R2OiG1
3Mx9YfJkG02Ozl1Fwm98bIkPUTx1BuIu7EZbstzUb0PexHr6IxVlIlEhWv2XuJkRCAR4L5+DxGRy
uW+L2HFmSG1g0uUnLk1bPs46wew1swUIgjxt8IKLicd9fKlG3t+/awMZCkC8Sqq6LgIzgdDuna9d
m6ZevgxgJebyfXaesxdAZtTU6S9moWnFTCsRFrqeQET6IdiPGRr1GZr7vuXXeEIEBTPu+yc4Myya
FRzoroV9qdcJ9tP7Bw134j8k82+jb85fTp7BjEWiB7fUt3HUj7dnG1OL22GAPB3quuhWCdA1hneZ
jo4/a3JwXpPOUA1WJ4yFENPFOq93YP46wIMsYaqPbtVLWdJ9x4uqUUgNy5dDvbUF8zdmNEO28krk
BfEG+FeAjonAZbPnv6DhXRWPAFbKppHOtE0cX9BRCmJB34mXkSETpzrxP1EyUCq5dprdFPE1w9Xj
bOIVmM030ZM5wyUVGjatVPXrdK4AvQihzPsrxLS0yLBzlCBn4xk/SDyRFvz16yVJFAAZxbmPd8n+
qVRZvKWzMXzxJdfISGZyvAczt5ChNStcWLf3q/z0kKfC3dXR50m4CdcUvZWplt7oLgw7YT0XQAUF
KP3q1j4gGIwI1MZW8A3N2Y0tbF2PkRsmX+bF+KgHxcQujSiDUHN1r+mPxM8EcWqJTkdbYnSq5H05
btaQkj8OofHJfRHp6Fznb/arWLHlACiYc0F2KfQzNnXeeHvHbeRPxUmH5zpkDwVWZ6IvG92vMQVu
P2ZtoaFJXkq/OrEnIwbYGrN1rpRRmbxNn4TrNxvctenbAs54dCgBCuPdIkIywm6e55qYmSRnL0yc
2/22j+Hfm+ISZXSjFCiGkaxrNjifoHb4UenOxRpDlJsXpplAYQO2DU11a1KREWBhczuWdCazNny3
eoEupPA+ylTQZlNKeumu++jFyotvLFyHQHbNEE5+OTR4A1Om0s8dMSbO0c3MumbtM2Vo356mcEz2
j3ESgo+LvutVNz/i1ARad0Vdzgs5TMU2pCmSNDhM8Z+qr3iVfkxr8z0zw3RTtB6smZYC6RqwNO5V
wGq5x6h+799amn4BWWhC0XM5Le47Nxq4vGXK/UK/SRLDtgUOLjZWGJZo7mV4kwaM3Qdhf2gyOK5n
dj1zd/Gshq/UPqH0h4Tw/zwcNJi5wzuuhmGwMgl1Jl9IuiRyHdtDaYrzlyPokl+GVnw5t+EXdSnL
gnyySMCaw2et5ogWEHzxBJoibyHKE57BZbt/iqH5ir4mwQ4bYeRDeTlsrjKcS6VriHwIH0zcK7B4
4VUyD3GxPs7j+I76w0r1SrTPUap18GyCBvORHtkQJ9N1QNJUB1lRb5gM6JJLMJKkbOSWlOrjr4vR
mf40psnS4WypU3yB5GGfJ/BF10CKPv04L3qrSYVFQ2bHvoyg73j/K+c9GmKdAKilVrAJaaZSJWs1
KKMI8NxnXjKhjoUYwCdcKCBz85+ICpieBDy2ByZavwPSZN5tVHApIoBij5S06ZoHUz/OgEcsuS+K
0Vsr2AMabEdP+CwUZ26dTRnNyK5GxO/P8LEtumXyQEDbL19IC3r/vaPfZhdw0KQVMduLEH4QqDsV
8BC/mFSCndbGk/j3GuqtRibmWj5s4MD2v1KwD+Tic6Y0o7S7vEsHuOdXl5TGuzfXTYbZsQSTCr8w
qgw6CQmrMYFud7Jfft2JtwrpSoSXs0qlvNTg9XXMr33D52EGt6MJp5KVokY56eGE+mSyhgoK9aQt
wb9XSqckQECathns0VRWp9ZJDlauAKs0emmgSU4e9iRjuewVzqw3HMTGoRyBUn3MQ1IX65InxzSC
dJ7s3YZTfMh9QqRbHwDAcue4PGRrIjyMfheHxrQiMOr40ZircMIn4TZCO1MfYztT8pIzh12C8jsA
4X2nWJTKq1gH64YLBkamQmfia4JOpXl6JoJ+ATvKejI99cqrQvPvg/PFseaIkkz6I9ejTGY3kK15
r6nnMuYfZl/8s8N4KsGuRQ6RbybvM/INzwGUlAgoYGJSBqHEp/7OKYhPg2+K2DU8KKrfx5xttprx
7vzwhUQlPV6c81Bz6gz8MbIbXGDqUVH9KdCcpCqAksd5hM2ZSYiGmrIsreOxL7GyONiVz/saaFTZ
dnwKxPXNQKpCbcI/vU8daKj+jXZf45zXzypuGnnxYxw99c0aPhct8Gdz/C41L4wrcHdNlW5+i3KT
kJL2kz41rqQO3QdQILnsTE7u2xsEnjcgM6jD/cgCEXfPEft99fASyr+NoFlgFXWFZjcZs3Pq9wVe
m7PPtz/753bfwpHiYT/pUKfnrHTH2jWWOX3RuD5JuRISvBUyVQ5viTekOSXjItTK2F3Lh3rvN1r1
bZyZ8b0V+IVno+gvBokCya/0eqGdV1LlstJ4Sw8b6Jp62JxEVpAsMDPoMn0kSC2m66Edx2DMe1pY
T3OeEQud41evqreAAAePwk2Q3Cmk1Ip8dkwYrrWh1GCPhZcr0QXGvRs7jUsQcllJx+D2AM5XjYr/
TLxdh8IBsWaMnWC4dZ5bsI0ruPlO/luzR7ZbzGy3IGVlWW/yMFu2iYsG3f3Z9nfjaZJlqaQ/0Nix
PLdtkjO3i6ab4tj/RTkJ6Uf+pa8+E3sLAlujJJd18rjLlj4qTL0LLGkI8XUANjuF7tgAAXePERti
cpHCq1rNOYBHbTNUHjPhDkDPBALQNWIsHhIWXqLA0Md/uUJKgsRxW73H0bZuGAZKsm3ufma2b0LP
9XH/PpRUGRMWgs35RGa+H1elircHT6mydkLvGvUFRCVXYPFGNwlmR5IuHvtwja1s4kaW/FYKcJPW
dPhPBVaq0SfRrxMF0c1YssqA5kShtb9nWD6HtJ2KkQcIah2VQD4XywzU3hhMt05++RQv/rwaeglH
ZTnkaslnpX4siqW57X0RMaZJj8yTGRkOGQQanNhMkjaGx1rHa4ptArsQHvRrejIJLFFszvFPIZXa
u79EyR1XJA6CqdIrVZpiKa9iOGBJGdKWpxsGd5ggWRB+/hf6ppb3PAJ2NkEsXD+oNOquFimTLSmE
+qjSoJrmz8LfZLYdMivjgLnK/jV8LQ3V/s3jN55bif22ocBAFuMUkwC7Kflarh8LC2pgelvF5/tW
Sf2XmPASIBsFJYYbs9E4d8z5/qXNRGfzdgtNo6dCPO3rKoqq4+5Y67iHbLTfZvOQy1qi5LaNHpUC
JXHp8nUm5ZL6iGe/aWO2MWLw9OKjQJcdV8B/pPk3mBFquU6iugSNldVoNnNAQd2Vhy59gmb8FwyD
TbhNcEQE12D7Z3cSByvH4NGFsLiM4/gZHNAENx/zH4CjoY3oLCzoAt3xtAPE4u41+iaulLeQW+kE
g6UoeZfuZBUbLH3YXaTH+LojPmb1U6qDFsB9YUFMk0dsXPf1IHifxYcOrpibqSjYtuIuuy8co8Nk
TZ+Sgil6ncR5VLooiJkus2s+Rz7m1kF+itHvf6au7HngBebqAzvvlTBcXr0qXShBHCLHo7mFkPYG
qg7y4JYIQZtiEcIkyvVUK/3UXpU7X47KfTweqZcLAGBXAPh+tJlQn+s6MMOG4RrrzygG9MG0on5R
coVLH9e8DjONKDDNgCOR61BsYKXbcdxDlhFh67NPN93vSbCsbtF1XESqtVMG0zn2Npp6uEqHujnm
EN0QiA0/dY6W0rpR3YRGvG0kSX0rqfzeyqlgcIt9gE/7fC+Ouubsdvg5NHPBRNJhh+tcU8Bqe/CK
UWGuWa/3ozAjCIzVQzTZ4d05HnBFK6kcfn6Z8FUjEvuVErnFqWDSr8BYdWSxf049oGozhlZbGsCx
0pmJvidFAxYCyd0x+6X2+H1OVbPN8XLyLSvUeWtUZrXjbRS5bgT9bFa1/KK8Gt/2tUVzjvknRPKs
nxCSNwbQ7+sUOCMC3mJA7Wh4YEFR0bZNtidV1YcnkNVLrwX4LM+lltOaU33LyN81xjNbGW0b+mra
xZBZdAqHGTZNmFkGpAbs3MsfBatyuJDm+0XITjmxoyAA75FVgPwv8eJXgnbo3a4YeTcrrklJThS2
A9/2zLAXAjcWDw1pWJsyxhmtgzFYdqf5G1un2+4XiBNX/uiHsP7WPa/hHq0zc7Cx/Z3g3hOFgpv8
k4xroe7Rg/xdxGbnR8NlN7FSFyYnJ6fBY/CM1B3hhA1iU2IeYFuOmzUVcwHO5E4/RsweIVDu140c
Qo3D7Kjnyk+wQtfaPtHacCz9lgbWfeq3PgIiZVRGU5Th8CscaHRl8pS0N8u+8UTGQwX/En3P1eiz
rl+OFeyb0ScqDtPVPQZA3DgnVDnTk5wGbbY45X8ilEJmAcVd6/pYp0P6LzlgN3Qxy35zHutnGOlf
TyL3WYucGziHNRkabQdG59rur1MLL3Nr6nwGUxJy4aP0xyKVOdIAxJL3I1WQyzxbItVUGXtgTb9c
u+/OSZPjyye7BlPU6XvrYPjMOU+WsP/2AQzb17Br6UN/BK3/lKo/qmT2LtKWhwVIwXYC9l91E5ad
I719aAJln1c28JPE5f8SOZl/DiZlFVDr3+Pe/Kz3Q0tu+N10hqjXrDgB/SiDc5NEJeIjc5w1eD6v
ELHB4ZE/S1trqT51gzC6X8+xcWMWL7ciJ5078+ShiwawGPWfKLp0V/wkcUtpqdTVT93u9q8J1SbY
1Kd/RgYkSsr9dE5uCy1SGOiUdCGiQdnUYpVtnQ+0M/u4UCyTJ04qdeO7fAvI8NeOTriYZhu3ZHlc
+2BNdLpraOsF6kdzSUsvgrak3LtOUwbt25NB3iWwGojFCpAcgGtJUDAyy0zYp3yYwCr63bOi2/Ux
hpHKuXHeQGBFqxJEvQrA6J6TRH/irF0A44CDjw4ndvxpR/4r0h+JxuEZ/rn1+/BgaocPlIj5x82W
hc7gzUEmjfUn6C0SY2c5oMhFG/bGWZl6mEgrsZCsLzL3JV9nfgX9AY70mDdHpl4WEewfrkRT16/c
JBaD4seuuQ0NQLy5bAJPVibH2MoQ0vyRoVhRMhRW39pLC3KbRFpputAiCEAdAIcBlIXHIgd/DHbS
D2kZ7yHsSDV0ewVYVoXWMKu74LOWGT7zmXu2lyPkjNCo5a9na9+IkG49vsiC08biiGjFvkxaYd3T
GAyVJkVjApxLgEx58rbH8sbE7Afqv8rTqc2LzCnTaP88XDt1COFOt2ehVXat5heuKtN5I+Nbs7au
72oJY5BBHcxXD3FJtPyVaopSJ6p4unVmndINtVcXOrQ3xqNh7Z9xQAfioZbDhVw1u5JRYY5cGu9i
wcVu/05xAA/OPzyRr34VmgqyEKyTz+lZZuqXwUOJUrnRV+Ry9H7RH0rXKhMo51TqW0UTamcBB/HT
Osvf5+CSdLcqIw6m/CyaD19tUd8ccSYTtAb4PI0LZYPgt0b2HjnzMkRE4gCPYv/xmqswl/HOc9aE
NUEaLvcrnTWYR9KU+sdJva9fKBAsati7c5VJkzC+1xXIC4gnFyc+ai1KBC2/DFV7M9kM7dYpU1pf
2PxrO2ua/+NysX5AsZquh0X90g6YD+qiBU6EPN9/3jOxeIpuGZsXc9IQwj/2fyEvsYUDqty3R7Jy
sP/BLeA6X850++tB3JJGrUBTDiGOjQ4ApPtj+39EI0/y/+QtbOC4za38kHvFVdvYZ+B8tt2LYraw
hZUHVreOdKNMp5EKydDwLzyUl011PTF5wd8xCNOgvyA8iVENQgH90/Ty+RZWhpSy0JGXza0O9JTb
MD/6XEuoXZm+7tiOJRwQl2+Zno9u/NcEBKP6uf68gvcPcwUWbG4D4CWkjNhFanMQdgk3wWTnv2MG
kcdd3BakRQqWMq/jzivViFGOLvg6HEtKw/iUmytNu5CGQr4B5tQRvUlheVM22nYyanb+Cq3SQBxW
jMDXTEt1fDxEwrZycDRqf2S/PLGZXBhCgHf0gSA4bINSZHVDM/TieZJg/yeKIaVU79QhdKkl+FC4
rBNt0Ive8NG5knCAl47XpAiHjRFR+B/CjXEigQevqPCfglOhl2STNFiWpoKkT2k9EH78ZJFkKE59
qbulDuI8LO9CdZp/ORFc2aYZRsB9FniLrChxeW8DahKErGJYW3SngEAJJrmarwKmIylCAXkANIol
n/0rXPuPmJaTXwnDeTUzvBBIT8QA2kLJEfblgK2PZjUnne9BKn2xgt4EqAijzfNLm8vkVdvg/Y3+
DVcQFuXb6SShg9N2mr75oqJvyUR4qUwXd+tj4FypOz0d2QMv3+uZK4jFfojUq7OqA+jVY1iWbqms
K5rTMBiVDj4gs7POMEcxU141jhIcz5bgcKTDW5vvPRybhPZ2ZVa1oeeEjIEuSVQI4pBtelVRtz/R
BDLoiRG5dzBkA7ot6ZMPnBRPGShfUdTPTbOOTw/3+FFTuwL0JHCNUrjuXIRw2glJ+clv7LHyx5qG
tzOHa8R5d01urva1nzqAF0tkLTt/ay+4AwVf1Bd95nWzAa/pXcyAKTCWebQN858fFOSoDFGAScPd
IYZNRIGp1L/cTzSfE7EatGWgjQFrXopEd114/NJEvj6Rlvx/5it0WesGc6eZM3FAXHJTzJwiyd3O
zzLL4J3HPyF5ASK0uplNMgnMhq96hIl0aqWQz/TmMR1Kzn/tYnnc7OJpeQcG9bQeRjN90vZN/csz
q3vQsqax6bCFR+L6PZYbugvKj/EWsZDnvQMc0xaBlx0VOZd1XAaGnV0gLsJsgol8sUZuMYdhwNsO
hBrALVLNLBVbNyWl7N5OrJDs9iUL9XoF2goXrspKQq5GcGclyFWBH6oXcYsNGJCYCLXNqPZZF5HW
gxmUA1GlyUrc5T8as00znbSZIKqyDrSOHk3wtaeBrB+Ezd31Yibxb47imkgE4AOILw9R65ttMpXA
IHvWifREfXReyaQZdUfVQpHm+CHxFEZ2ZvlYta21GKrtow6EsBp79YCNLTeX5COu3biR3HNf8zWt
QOh2oqYGOwPHc9FbuhI6VzGHWiNn11NjvZfLnSYy/+On73CmgxyQOJIUQwOkVMO0hNhRdwpibRxw
9DViooWNMs75sbPsRVJV+cDHKiQP5diheTVTs71o8eRm+06pYzqaMWcOyJMF+Lwldp7sUFAdI/su
XGVoPvl4M3XyTyUD9blbfKOuV6TApS3XZQnMRzZZ3+UEPSj4DyZkStQywgJw8UHQtcs/M+fliqyo
3Woo8/sn9621m+uGbsObm4O3+//AmTYK5dk8yE7KzsCOCMBAiU13xtHeQB4oLebPl9K3Bo/kvPJr
hCrdE+xXHu45HIWZ27rBYluVlBD75XlKwrGRXxqvEuCtYBvJ+vZlglyLf+y8gp/mC28OKbxS4C8y
jKYrwG72a5NPPE7hhIEYtc8vY5SUmBIFjfMclk+j/7qc99XZXalBam+qNX+J/NKI481RY6hW6EST
yJtkNS8Jnup6Bsx6bReRgXeypFDGRmySRd0i+Yx3kaZZ3ZpyB67KiwuVb6XUmk7CgmHxOMt0nOIy
Y5yZ6jBGBxp40krNi7Iailacajx6uKWw4Yz7pPsVw5CtCpVuvsyMqaeiy+eEjoILk17x5KF/krmd
SFnVTQz+A630IkkfNafLgjzYhfElyCpgopJL+chxGlxokt/grsIzfErqpmhsPpLbAK2um8ZFepHH
g8hen0R4Y7lVj6WDRiCbbBMkYs76+mgQJgzQxJ9yTQnbE+ZcvD5SsOXWgZjjxAynfvJ2qDn50W8F
96WgJZH+elod2q3GyKIoOw3P+aMMIJwnIN4J98ZeszYuXmgE8OidBpI+dRiibmxUN/qoanNm9jca
6wRYvQExcgrB7px7rp4a688kGM48Bg4q4u+UJANcm2nCjsItkV2zlhJsT6gamNmDnxNZBDHgd2sL
HYLEy4n3x6MrEBOFPb1UDl2xhwL2PVGy/wivJjFxhHWNRVtTQuqfdT4T+BAbXy4lveg9N23IRSUt
mC3fHQ3dbYv36s57M+OJEfuTPVvWlQsVx+gp+Ka7bCjGirjnb/0w2fZB7ead4dTAl/VLNctLnf+6
AfLKspqxwgcBy7E51X0RfqS4AA4gscdkxQiAGNCjZLGXFKvIc8z+ymLvymHU9ncJdytCrnK0kOF2
P5fYqF2+6R+TlG0+2uviVwjzwPzovAlKAKBCccBPVnnr1XvZDu4OjSU6NeBX4XCyJvRkBHiCV4J7
9Z4IAvAMrGQmG97T/sbRj3TFrxi2zF3lqUj4cCeQkDiPLkkogW7/IuqW8Hy/X8QzJsZrPXnQxxuq
y3Si75lTw2Pjfu18onvRAODa0Y5psmRohBtsJUxU1v5BT7td+7OK0cvsPZ/rnR1aOiIU18q726s2
NBl9KlmCFE1mHcFRMQ5r0tla3XgsBtZ9hwrrLShvp2zh3kV5c6rUvIvqDgh+ueNQer+9vb94i8re
cyN3LFpAsLGheARXN42I+0OsQ8yEiZsLxzzh+0P0569cfwRIV5yJWrFDONP+K22AVOnNr7uYtezC
Sq6gtaHQLdJJphLt+C00UxQAlXUsLOoW3nN32q+ROUK7U4tHdWfoSlu4JrvzM8B4FpHQH6/TrD5e
i9OMRsxRbD+bbeSC6rcBeH1BXjsqOnOv8pn+4xo067hC/snFduJtE3DPXUZ1FkW5seC9HOOTJ4Gb
UHR+Otk1FxyLds9YAVc3OCakiEM2ajijlWUh24ZuyFYMbu2K6Dt7WQwOYuFzVUsl8lTuAP7JnwYY
BGkLuyfzo915ufyZTbaGh27lpY21VsD0KaltDcf7Sf2Q98GxD+U3+6kNalCL0iECcTgnYIZkEalW
BXSPMkTi12OSpqzoqzrxLJcQGlxhZr9fWxO8vXsfMyCWVPaUm9WjE1xWsuQtdLdQ0HtxDTnoJfJg
cevMbxCBVhXQfephjwIzfYSYRNoCcRQGHUkMK2OX4W4cC2LnPWjfeCvye6D6U327uS/I1pIDqQKP
+X7KudxzGetsmcyaoOngba0NfXWcSYYFx8QgGYnzs6XvXPRxgUbqbZDezr6vpLZ1dugC44mkGk+H
ON6dsiWyJ09SsKiFXEreJky/a7TPoIF23mK8WNtWedi9F1hIffvmuxeSxjpd6iqtzf639knnHuNI
19HdOz7DeM69f8ZIMtxywHTE+yTPmRumhq8fh5wfG0B6XjH26HWaT9XuGrL0zGqWs0xAzu3J9oU3
deklvhzNS1s5ow1LyZ3G2qExo54rERaK/wKBhCll/RPvGm2lYiUTHdiKepYquDzjZq5dBs9+zN8V
3kYxyjuF6sVm7hWuqnQbb/GQs7E5jqjQKL5e52lVsRlbXIOFYPJBKA1Bcf2Og3yFkJOJlZcIKl+1
pa2kN0CIwoeTETZJ17WowS6uAXQYg8EXfgTOZQkSSbRsyp51Xx5sx8I31rpOJib62LLU8meVrOPZ
zERqS08NDNWqDrZ3hU/ge2Z/NH85yjQdjuLfmbRapv86qtdyuellsHBmevnviQn35Mt1GWzLKDTy
fO42Yk+n1y0m3VvBK80523wUCX9xEfq9lpHRuUE1x5aAbmfN55egfRIkLBYMfnhnW8dz8DuefEJ+
XkUsZz7kmZ7AHPpkHiEfE6MSuYSBqgOpORQLNaY9W2+nuDDRflxP+ZvNtBWSfvBegXYg32LapZcd
KnUqkzSnPi4PXyIzamA7xdy+ckDMxM+XcPtpQDzGD1h5ERaW5KDnsHi/xMA/flMaf0TiWlpeYG5s
lQHJgQlzwKjIO09G9im1HV8jXfPtCXAUudtciTRGsOAxBVFk+EhqYhB4Z+yWx5CgNHnBWkYjecrg
N9c/3HfY7ilXA9jl36p0bHs3VPMItJ3nFd6AB4vZF2w7nwIxWlpTkJerSqzYF+OavmZhcQWlXDj+
PkhwLMpB+8Lq9Cu2538SUz3MrdazaVUzIEvnbdaHELN+7OWl1vtFT7eXxZfYE/EZJT81Fh1lCc9J
kCjg+087sBWKwRJPAWy2VQOPFXrh4zn2/C3bOaYRO2sf1IDGCp0btOqVS0tmYKbJX+D056RVP3qP
oTGgIrQbODvKZ8pROLh2Kcnfmc26jWHULa5rh38/SCR1JLq0pkiWSH002Oop2NfW2WZgXwD3+wKH
EGMuOLZ4GbSr7vulwG9CUke5fD9QwpyQYRDBAXOjcpybn1GSzb1jvB/ggraS77va8uB0LZiDeBS7
qf51AiE7RneeUYRrkf97AkoXVgNbnBK8EMXHLcvlECz4NMuUfyPcH7dFxzxkqsw1ZT3NXkXxUD0N
JzZDi+t0IDwkdf9PSqxI3eOWFJPvZhEOGhbPkj2tZIOnpZGnBqiPm3Xs0oCamh6UYiAeWA6pRtqp
m9ZKxenYxalt8qjJO7kZ58Q1tLWEjkucDHmj8J4Qbvn/n0TnudFubQ8JCPZSMqriSa9Laco/yvd6
CtckE8fnuLP4EHd3PzrqxEljJX0exWq6qzkEYoqIac3eX7p11t7lvsNnQ6QZIeoJ/SP82vCNCHk6
L2G363UM0gDOcLlbz5p3xZ8HdYuB/xyzZ1o9R9JQXBHFAdoRXK3u3Wsfnse+GPMKVUylkE3+iNT+
SqenfdhAYVe4IzwOF6L5bQOQe9O9qSklnez7wc4I1ZUftrMrg7bXMIthJJbYxgqioVq/i7GO1F6y
+HwqjwFj2nDzJATsNNxRBgvw3TuJw7PbYqPOWCNzTzjWOaPrvvGC0GRY9jFrXkOU1fGqLNCwhmtl
V7DPnKr3XI9d7y5FbbVVkacdHbcitIjxkmSNWwMokfOKAHDcSSyXu+fvwjT/U+bfO0e+l/ndLazR
GnU/uUiByCefIrJoODYPT2IIsz8LefAQMlWr/UyyFuAxUpG+ZhIlpDM5FnaxsIQUSLe6AjDcuyjO
XLrdeuQm5exPhy6UR6udwttnbBdEPtCMMo2cFvRKhOfUTqtTD9QPSnAwexqTnm2aO6cIK82rpnee
TrrtoAmH6OcYQxtxRtBCVs56TVvob96NBytX9kMFR1uamOs0rvS908lmOsDUiqPQAr0UTWZCpeMe
wP6phaE5zyU6Zxz20187BWilO7GDml+EgBAHTAf5gf2D0cJfUPT8W7oz0P/Q7TXZV9Xhop6tpBM0
xzcGAElmU82Vn2UN8C0LjlSyUarh0xrW+XvGlWo/BjAnpsU4yzADW8UP0DVtcwsDcZgE3qTxbzfS
YJIaWwVHp1adeKBpru9itLZKrYuw67ADNLkWlBB6HKlw8iQYIWm+9Mr987aEk0AitHl0ZcGFuVO1
l1E7SFSXUyH+4DIKquImgNB60Pj+xojBoYh8lw4FZ3yAhvPPfRYBGA3d2JiJLbsmSofm7UbPrRTg
XzxEU6Tav/wa876DD3Y9v0WBKvwBSQAhtffm49GodQ7u6TvqUCLHlryCaGhZ8lwiKfm/IIDtJp/x
NqU5H/ze6yxONbtiG7FPciaK6FoA3NaGhqfaPFXuObXQYFFJI41CRrWKLxVHUqV1CAAsGB9TklOq
bPvcXR+dKRoOMH8zTjuXiDwPi12fq+uamsFS5eXMiVNhc5B1cdjYYmt9QoBmJetZtgQ5GcTOHe51
+AzI5n4rVhqudqoyj0UGXJeV1Fbhh8dsxMm8AqjY83cDsNsgCqbfErNXZxzikB+Uc/KvgbMrxd5o
iE7HQQ+Ja7F3T7o+10BpZOLxlzIput5sjVl3rdKUUCczgs9X554jLVvAzimGjhay/QWRCttX4cyE
BWIsgOPxAIYovGZuiUWPG5uhOlxMy/kY4cr4OIw+EeskNuXN+cbzVXUkSNapw4lbogynIkbSnHys
2pC2AkQ8jQs6ZwlcBTROs2pKz+S7QGVzw764oRUBdzalE68rrs/tFB+Sl1yis3KU9VH7irlJFvs5
EvsiaZKrnli/JPfNaah650/LqlAu9QNhqpl/+va8aeezOwksG5215yiSlVzc0mTHPI1a1teAy0i4
qZs5892EABv+oxjG/mHAqD4wc3hN+ryyGzDONdMQYAn8Dp/Na9IWcc8V1heR6DIqIKgGpSQLLlKQ
flwXY+J11wzsSKrVSSIgVGBtOBF0fFcdwf1VXV7TLSHFlvtUq3llpYS576XYXxOupt7nnVf8rvjN
tGIrKH84Mt3TcCWMU0TY5HWNYz47rks3a+HraZK60ArM0QqsobzP7cE1BPIvSO0nvVTY/M86kmKk
BK/X7oCBInUPu9aNHZ1SxiDTKVj4y+Z5dlmRBhslbok06dmjPZ5NdUwvqeV66RO113FBXswhyawt
Qa5G1eatPVco031XdHn/Yc8Ht66eLBEZpyWM1hQskdZk4EUveveq1Hmy5mRieFapPf0yhheS9RDS
rNJdSntm0PMpe4k4SSWiBWnbwucgi4s1otlsHzfsEwKXZHp1XNF4Ws5vlNoDGffcnT7CzZ3dso7h
y6tVgxAJjgWwuLRG1s6i8NHdAtU98+amtPdKj6TcmFV5UGWrrviZbnb0TLHDitZkr3v1haR0/Ujs
Qew1WXfLvuecYh+GKLyEbjJX+mgj+73Fn9EROW/eOaO5q3T176LwsRirUnV+/Tb5WXj1+Dc4QLIL
biXbxng3b0kFo9Jttku6P7wooLCYkpRdvrAZWIeGj2fQ+CMATsmUjXe5yz61qnbEkNKFeuvWsSpz
cI2RTQtcNrqWEx466n5DpnBdo9D03VGDcnxrxT3HejJmpKsbRpBgBnC291ItWhpusYZMWr0sjPW7
qGGR7+U+nKRMH4Qnr9Zw4jnSzd/AfzNek+Sz8v4JcmXj2+r/hzjx4AdXxw1fVSLDZ5cdKjeF3bxS
8Mua5wKkMSQ4Bk+Koir+UgPX+y/f8MxOMAw8ftntTVOIShJj4R7UJbCx0Hpeo6v7G3L+jJGXDEhF
uu0+KdQp8QW9CNdmFrVfVzLi/0ZGLo/ZocrrGjPpA0N9Nds+f0UHO5MrUUC865NJvNwokQR0vw/w
bmIATiIi1oKNnH+Z8aokEHyom/VSLhVDmq4wO0wCXpxblirKSnGSLnjyWFueY8gUrKJ4si6kTutl
nwtgm7KxP58+KMkK3FPKoikcnqDEhGtFQv8TvLg0P1GJdX+1pkUEmxn/pNBEH5cQA/BxIKRyS8JF
wFFE1wYhcA1rwxpzK8OhsmE9XZDsPlSM8Z6XwLiTtLSQuq4E1QKFq6Qwv+zRh240I9opS58CZF/5
oYgnWXzrsELPmpkI9pnxdNKVa6H4GDNvMaXhSru2gHPjuQIdF7dlY7axH/lfzDalsNRviTUmdnRS
+vWVoOr8/5gKbOiQP/KNy2yDnkw2Bv7omXojkiLIrWlustNV3lO/ANVY6mJzkSJDggRGzTk261Up
OEGE/AUbknP7WlJnv21fkuClfp2f0u0F3GLMom+cSb4dhTX8QS30ukH+jLzfBSho83jzz3gp+ILF
D/GGGWjcWOPiUonJHmbIpnvS5zZWSFtZ+MSdwqFOVUb12k92e+DRucXxvq21+ycaJVpKS7Iucvoc
GmU8duqbKY315GFZ7WCxE5iIMJ4/GS8FaYPcZr0aZVPfnnXO6yFvkcSCRKjRD48aGFTBEMxFGGs+
Kgm9rnP8U/Lk/fzS8uS9NAHCZVbYtQ9/LApmjx6bQT06UyIWpevIFPsAu3dqLYLD1vF5Tm0hfDvw
IsQiXazU5bvucM+M5f2xhLaLUcpKOiBoA7o6XtDgJWQvJTWufgeoOUJEPZS/qAdGF7zr9uw9b9iK
diJpclN+wDBj5MpnFctPERgiWH+V+GWI6/QU9olny5aHlZITpukKCO3So6bfsy/PqWqJwQzNTsiU
8EYC6vA7/5NOwOCpFWxjrOjS/hq/hj4wLidLGlqpbZwwUN9DmDu97X2N7YU2JNKr6VyV9xe3SWoB
tDyyhb6iNizFjEWRWQm2S7HtdV6/USnYcvQ9nKKY/hIuqDhdn/T27UV9Dw+uGJWcm+gFr564WtUe
geC/9xeZdJpT/a8FDgaRe1FkTRKWfs1kRjUFhLP+O+BPLW0flGEd0bW37jASQ1j+JMMb0ydXqEvT
Lqi9U/moosQdJ1/Oi/E28px+fTeYF7bFJgfqKufvW54v742lfKDAfwXLcakl7RMjgLTSEXxBQVQX
yK764AijR/jTVc8Qyud6u72CLBL0X/O3qSDkBlWYz8wt7NRDJ5aLzr4cTkO1us2FuSQ3RSpP9BiG
h6v6prj+/PLHeFgCUhdagEV9mnFbdvcCxO5rh4ZIbdKn+Wp0LOMuLx/fmna+o+N5LhfB4hdEKEef
FASdohoG95oor0QDIRKkxDJbrWSftJSyn9aY6ZfHjQDbCQpfnxeUot9MXrJhblDdQXK285ZRT8XN
rQ4gmaHomqbbugMUdaw6mJbMXYVUVej4f9sUDPX6bGq1FU3ECK1m/HslRoHMHfRGvxoUYealFUEy
9XWO9KvuHCCd+mn+2DTYBXSwb+C7Uj/D2/59jcHHg1WF+8nVFghvzs1ioN2zdb08hwdowRd848fR
bWI87+BwPb3wh71Zuwa/etn9mq6FSpAZN57zSmHU+YawZtNUH59Klo8u5ROlJysU7CHbZPKuHioK
4VH22fFLRN4p1uPiyycu+PopDl6g9qebEE1/CoJ1LduMIfgr3JqBd/qrCkIzgdapzp06UxLrLMFY
5RqVSVtRiKM3Gk30hQHj5FaV1nQCPkeji0jStesPys9FAikDQQqjN6Hz2yIZMhZrovKU6UUbhG6E
dnyVGdaO/jpTuaWBBRsiZkiek5x0ozdXro4EIwRuLvj5rKW/cAOkRYESx26VHMU8aMY22xBt3lsq
5oVlpfEV93/iimE+RDqC6CSYsabIsFDbVa8a/2zNyJROnyTwI5+AFAn+6fvr78tmmD1hyu7zxjYK
ks8089H+UBQV8Opiqo6WrOf83puLWLKGfD4S6bqcMI4T9OI5kGotxR3DLS0bp3uBGiBdzSx3UVbg
2ofnTow0w3vccdYqX8d32OKkyVyn1EyEwaaazcuysfHweJIvdsMVBenERxOwt6X6U1tt9whsrD9q
LZMBh28C06nqSoagyJV8BJ+qXrP9ofMFZgCfRefZaMVHyjmwzzkAQj5OVk08RksAec7ymHgrNFm6
5p2jrCths7/aIFhIksHVGQSiImdyqX+rDaZHDJRUSpvb6RS4yeUKJhtQ9tTK45p7qO9a29qd7Epi
3aWaOCLeHZlGCBX6OCpWWHV5x6/QI97ppbK8hbdwU3uJS/K7U/S6W/H2pBk/JFzmOfIJnjJTyu0l
MZDHVqc4Rpj/3cnNGAVaPM/D2CbIA3wgMbVVq225PXljisHr1ykZHsGpExABbPCCTS+wctFy6ZIC
rQo0Rq1wsHaLjLU1EJrUB4th0QHxPFEmrh+MhGTHZnkXvwqsTq7Y71xP4Lpa2ubrIW+C8RbonhC7
YOkDrgOdcJMRbqas89vdAPyRqQGrWszx1eOX3TsHWCJ17uEkKcgVX8QOAtIUO5SlzOxBLtiOQQKl
9HEJBJN0IK5k9pbUiROV/M5J0LZKATA/NyCvwLm/3EI9aRw1382+dTX7vdUnpYW1sor4Bii4YBuM
8nsNnsJuD0+neKCY8u+MFlqy98pSMURRz9kj6ktDrlwFYZBG2hM1A0XILHBPL0asKW0/gswgmKWN
4O0tQl8hEOVgeFS+2BpISYbSKowt2+vZCUWAyE062Vk81TUZF+7OT1pkrGPKO3GYTiHpnQxR4cja
Yhy3ZN5c6N4XpSswU8M/bAROuIKPf0HtJpZe2+G+X9h24yNIt0sSFn+UzoaOh5zAMIQZQ2uHawRE
nR+jAvzf+Qzue9KvZVk3nFLkq47eqA24IsJQLEbjInFoR0XKMsd3KIQOvbcm12IShLhcMGlgI9qY
R4Tdv+8bynHvDuOXnI+5vs+l7R+jsruXsUGJuy1stsxNTi1LsTDVDdyvXSk3/xZ+gThxQ/IEAQny
5MYZijzrJP3brZu8nYjOJixKIMBaeyZqx7yNp2A1W449Qt9lDODdkJYCB0ADGh1C8LMDXM+5Zut0
40N1+7XqAPlc6vLfks3JUuiinc0Dc+Xqb0lGE43SgMoHAxjjy47rpp/k+Y7PbrWR87bDvUvoguxH
Z7U7XfjFkf8KHp/rxMNFcPZA3aZpHcq3Pcrd/+QLzBljcBwTZWU2c9ut2DCoSM/6n3/rXWMuGTkk
TnXkK9YWn5NApr6Wo9M5eRLMePCe8O5oj2K/h0fbs0su+DID+R4Cfg3EyVOJeGttm6+6fsuzF+Qh
E0zZ4p85VSNGWMU9iHvxMN8oaSiqZKm5zH0BzJUfvJFgH855olKH1pPpyLUIpK+D/WNK572cQkd2
a7OOijqKtSmdFRKj05w77/jn2IfGy1BgJrOkLYORRIpD1DZHOcefwlLW8CzPhV17JzC+I7Juw9aB
az8/LfxfukRlRfrCVPS+94m55w0hE470ypvgJBg2c9aLAcNgXfZA5JiocRt4LVu3IxY60He2CUka
1Ypm/Fy6vEjtxm7aABfvaEPyXcD0cK6re4vrzT2o08EyEiGMagDiUD+1T+4/DrvUuIJrJ1B4QXkT
yFo+ATuf6P+brWQGXQ2VVW1+NtOoVurvGGdD+8BIw9F1StGBo/djsnq4sRYQe2tsI6UK51MtTIvQ
3OJfaMFznfnGK/stqwBBWcDbB1CBLCVxcFuu2jbmQmLN1nfpELQJGzxpe2DDGNep36CcRU2J14Hg
Q4fJleW8B1GP+x7+/VqCCwsMLCW32/GO8+u16dBjkMzPWJogBXhn0huOt1PkQQG5//6EYhAECR//
4107G8EjPNFe5MwcrHWIy9pNs2+Upe1ylqdSq++g00E3YDv9FbALJQmxdF0SBVLm7FsQdNIqyswS
C9epKlOJkIAhzApPLG58H3Rbxbl+7UMj2FXZIUe3DUd5O8jaV1RWNBXPrgV1zihM4THQzPkFAMG7
B1IVggbqMuK1bu3fOhH8763vavufK/UD5Kg02DLJyx95R1fhQBZnW/WJPmjQp4I9jbU87FGFrBQ4
KqKb9er+d92iHYmK0rl7bsJ6PBaCoMoa7w8ubXrXvFjtZVL5TAubih+82APeI7jWbLBGeVf5mNQg
jMeKMXm2MWxxepEQk4ddliK8EdoTEjw47carSG7Hhv3FhSCg42+NsAgXdHgcxx/0TttCFjrbfNA7
kWtC16mY/dxpPYf9f2NzGZEo/+mqhFDqJOYI1bIfFl6EJEQ7PyyHCPkCNoj2DrJLJ8J4UugDWTF2
Ut2PhO4BFtd6X1Kkw3VtKho/QftKALAw621xC/M2WmlKuVOOxF9CDMpTiko7N13KwF1eu++/Lf/C
NtcBlIBge7oiT3wqb+L7dmOYhSf8O6+ZzJ8VOHWX27x7mtAcOYIACCT0XJIdg5WybNqA5xNqIUPQ
OE97/21jiOp5uc8zPP15+KcMjYOgNaPZ8sqllVzhwAR1GpiwhrS1gnPTCrZP7Skc9f5yi6y7pH8y
ZG9Mf2TjMp6XwCqRCMPVukCgKprQuIK5t/ya8KDysO/Jqtpp5/2knWtLFSCoD9I8qnL9YGwIfSOY
p4Zq02EKEwd+NhbFZhu3JeX5N5+Gtd9Ou83Wt1ISegfhH1iMNp3+AEd/mfdbO/CLcGtpyhpiURby
lPFXcrDy6+0uKKZAJibJMAHnJPB0IwKEZ6DpSJRYZpC/uLxZEgsY5eFpVHeoi41alLLn3EtWGeBb
f6K01+SeBS4pa7z6zj4MqzfNoo+uwmP/0HRJsONnt/ajLSc5aonzBflv8xch6GDHmPa5syk4rhZ6
6Ky571uCGBohEaJCKNSHBt4ge41TZEHtJo3AkM07dJ3KcuutDxb0sGFcScUpoXSFizSjbz10AxYw
n/kZxxWQ066I6/ngUMTz7OeEiIn8lgf6J308sZhVQNhdn7uZno79ZoQW0PpIrGLadtQFD+S0vaPs
6VPsAU4MepDBg9Rfromoi3OW6mFbqmnOjcWLbbA5szi1aYlc6n9ZX4UtUEzwCh8+xpyob0sDYz5t
/YkbRSYHVMpvKH5hszft9vrI0PtpfaYrlaRTkAyO7vOdrW6RkpdQAh5+jCFPx8bsyXVlCOU5rQ/I
5P9Tly5gtpfXJS3yAY+E2MD2UDWQlZbTTYBFvN8Xj4+Zzw1yK6sboKqZtBOsvWxXaGMQldwzkPtm
r1DVKSX3iwGS9oG3JLh8lQEiUSD/6oD9V2BeR+kMJfO58s1uSkHi+OJP7uT4jfBobN/vpeYSl/Z7
FCvYjMxMY0nv9eBoH4aR6PAtPOxUM2ZU4wWeekKPEPY4NMU1HKM7+zZB9CKtQQwqTEk3fQsGckCC
dcZndvLvwWIU2vCk4Mx98VbhZJ7mdxnOGSLk0HPtIqxagcVZnyRinhyUACR+xwCgX9tl7/1hQNDr
3EkORgZ8J8fTX15tqg9t6nBSM4SAXVLKs/p3DNMmz14kxDhIpjCVstbORXPOHs4Ie4mQmtS7ZxPg
N5IusSd202eVant12l1MQ1I2PDv3v9MrBFR8rpwOfRGKx4VFcDmfmj7ftLIY05HlIUZAOANEPVnh
RL/Q/4YHlQc6M1Toyb7a1hirNpLY0aWGAHfIlR49zUIztNZwsbH6KtOFECEyxeInwGJN9Op+Yn//
9bWaoGdOhIy+DbcKbsi9nJze/SHflyJ/ZmROfPvFuikrmCSWcgHH2OZBpiARdm5xeeqPjFq9xPjV
HrBhlveRezoY8ToAiDdL+c3qix5XSg6TxMeLQjMQ180/j/LUCXkU57d5AAbg++3sMjru1abU1Qls
Oz9L9XiXiK8iacUWArhTf7TXjrvh+YB3g5iHZDhDwOi7HOQcrhsc5kOebf1xDlDAxWIk0lwT8k8e
R0c5KAuWp563mp2Fz2JRBCnhScajylK62gGEPZx5vqbnzyFbZDouno9mfl+r4xVxrog0BAP6qWYy
FWCHVCRu+hZ69iqyZ09ZDGtM8v7EGcRcB4un+XsTToimAY+mL4tT1FnemTXj4K8zMazPFAj8vAtD
YL69H6r8qJC9V7/CNd7S+BLaLFtMgwR/gy2vOhJFDjm7nJcd/kUSFa27HRbTKp6Rxag0MX0x+4fK
JsrmNpAYLpBWQfzxCB0r/IggPNBpRsov3720dBaSNYd7K02LVKhmj2g5SMduiRiPpekl8FDGt2jr
Km+LXvxX2cCCupquc+laW+oV4tNX1oBovfV7sYmXGjI4bKHHF6TKoZG5sIx1jqeSGliqw9Ij5xZz
9CCnx3PPRrRwRVn72C6Cz28uBuS2Y8AV4FIMnvkxFpjCaCp9LMjzBdtQq37ef+4TyXu4KoCdmPAp
H9FQH53p94kyT6XrHs7dwsE1/6seK7Pn0XBVwdagyYdb86pHnK51RAdGMa9KBtFH8n1aj+j07XXf
7SdqhBXavjfTLHu37PfTAlWSmqKZKkelowDJwZDIzJncDqfVyuwKhhmEdsqKSScIDiThBL1rcyT2
R3UDleJ6SadvfrSJ8DO7G5DWrhrCsvIKp5Mu+xk5lbPk+sVzlPthRM0ozMwsGWHNkPHrsajB7RwB
lPL5IfjLIH0/N/KihwXY4BtKeZyq+WlvY+WXibS3Tja4oPiHdPS7h69D8U16oeYY5CeO5/LE3RSE
Jqt11ms+sBxiNcehmMWBWDyRuzYPCDchcp7x85mFK6dQUxyqmvh0kV6QFalFevTqy+fJzb/etB3P
4ihxyl3cBfcC1mNx5kMjz/Nl7OXeEVJ66tEscaq0BTs1g19BTaufeTOKNL8wwBCRDxt0hwpUO+JW
TKWDoRseMUTLvZFBqOsajTssm/COpv1L0minOuXRjzPyT49EqiCGeqDEnzIMzUy/IOr8tvypU66c
eQgtKWrl7dmwLTBNCjxUVUN8xRCg38UNvU8LBmn9m1YSio6m1JEJXgyMUHrFaiVXiTjxUfw87jdN
c7I4lBjfY/7Ie1mVCh0DyPF8ca8LWc8Wi/ssbmi3RQTVulPjM/xwR/4maC9sk51FET5e8p10Pmzl
bfE1+QGrjA6w51v/SotozZGS/z+I9soZ1+LpZ61fc1e8JmOGem3gWRqAzrXSy2VQLW/loJ0V8lvK
pxmFokzMvy3s77EQ3VGVyKA0/eD9gsrvJcX7ubyBjm/0EAfhHUYiqL5z2vAtELV/X74STBRBIThD
lOY8NlYxeIXQvqExhiOyaPQf1kvQ/w7ZXN6IoAaKjK3sZvMUrwtMwWXg9GthjV4TqorxN5Y4eZ0g
diDBz02M9hHwST/dHmagN0NpZqmrJv8r46Gg6b7oVxdDM4k31F5xG+rAScC2PPb/T06gM4obgkoq
huZdk6B8hom4rEKk1uzDVm6MOqULHNehgCO8+v7mBps7VW25Ws4Qfej3UlwiG9ex+VW2z0j73Lec
OsmoEBJUmGQsEu4YFHo3GjAJ4SxoyjYgKFPxCJID9hVIdkhoWWwRKFJSJLdUHqTFNwnWKLe2zK0A
/KMeJMtyz32Q6SoWXYgclj/E608Tt5wfZlh3Ql9rHaC5XzHZFugtwma/wM/0BTy6Za4ySt6Utjb8
AuSaBDMRqIikHDvKEzJgPyhcE43xUI61nAN46KMTTSMGU5398bLzZN3ZxSfxWLz0vpyzwtJ4Yh4x
UYuDwy+jHnNfomFzjsxr7f9nm+E11lElW0juN23w1VWrfxxFT4y3RPe+BtfQ0f8SeNI5oPfsUaYB
QV2oXF4nEDZKUI4Tef30AdNnebROJFr+R9VrKfeugRJB1uB1BV8yKRVLzyWhxy2sNqXp1e5YnbPu
1hyzaY459J3nO/dk4AepDc3ChASxSpUrwt9+E/cCXXHtCmPrj0rqj1M7wI1uIrxe5/b+K+Gj7h40
QYxYW0sgbB22BfHAXBZ68Ggddd5jtfV5Q3jb7CzdFzsPQQVLINMZHv9Lps8rMubllvdBYzAajj+3
y1B+iRQFRh/AZyCQnIhva7URYfxKS7GU1mmmA6kRerK3KqVRmwz6TaVaNVfLGqYP1M75IV1Rj0MK
IFVTBLi5e496sd7nEezn+kqV+pfFl8flGBlq2IpGpW/wvrDS+O7KHD4LBl9heiGNg0guFSID/RxM
Mf1DvWJEUNfFFIcCXrFPuUg/fgG5ZNj6yZMogPmj2eFupU183bNF4GVtN+NqXxiS9nRdxV80TFJM
jeVttmuX4tyGnM/svm2u7hFGJXgzJLNN69r0wq7wholWAMqQ19dDRMEZ2CgBFnYbisRHwNA0b8lf
huGqzb3EL1rcwLTDo6noAWiEbiXz9Lb6bSv6FkGUWV96Jf/g3BYpa8h8+H67vuwLfHFpoWkaPRUO
LAGayuzLW/gq3fdbM6gDSgj/CVrss7sx6c/uwF5YXoeGZE8EU+vRk6YwzzCMe3Go6Vd8t909/nBa
lYUoLqGBXp03FB5WEBLmEvdAGv9OETABpX5oQDTvRpqAgHteC/bFMFx3DBgN2S6DJwwgq4c34Pqa
3dQ1Tx/a2oI9l350NDbrM2LkRo7gP1PmKVGTpR+6Dn4Flj9AEpLNn2I4UNjIYZN6s+5FWyyy2ug5
jqcC8sj08dXu6pjLUa293C8TFbXEJ5uDXtRKxaOkss0ROePt7qZplDKfD57gYdUS0WAP9NNsW/Cq
DstQNhPBjLEZzeCChqErhgg21FkFbx4YyyIH7MbiBWbPNjw9YxYo5Q9chU3ZLuBX9A+EdUW585IC
vTU0Y10SRcG837Eczu9bTyRhO7hgU/Y4z88OeSpaoVz1crhwHd57CzAGX/Xe/4ma1KSr9+vE+psg
kH4GCXLL6ckkO0VUdfURk5fFLbaShhyQoRPdq/IZabLbYfxktiq2IoSp/QBrXcQT68KbZSDwBqZW
ZEJ9F2o0FkdDCbucRCjiByb6MppHb897bgkbFqt039f5AsarY3ysYLTX4Hc8GtO0HNOIbpekgZDB
uB7Q/TvCRGXM2e02iLuGOOBmHkjzTAp6mjdx+BEFdsXabgA9SJWB9GfODvHLq8Y+nQIeVS66nbTF
Z/9MjjzynJX/0Dm4iMsWcIIBV9F6pMcONRPUzqWaRvelis6TWRoFUY+iPWcoGwblqlL1GNF1qHYg
TVN/wz/zldwo+9gm9XrBLZR2gq9pQ7A5fC8JT3slEnXbKbL4XhWfvWlwr9tbXXzfVZ1zsEEk3bAB
1YbTt/gGLS2Y4BiFKdUtG2YlV8dj6W1r4D0650wegFKOhKwGCSaQ8alA6Oc5MgIXhBEg/Aiv9rrs
nveYHW9z7u7gCYSdoBJCdQUeonP0nDe0S4E5yWpwdvpULd9E9F1p21FalFfcngNPQilWWtR2Aytn
TKqORzWs/H8ENc3X+Za/YNShGP31zOU/iid4AyJGK44XDWzD51PEsZbvhsiU0PVjkrMUsxaZGuk8
y3dc3uUqdukOoaqvr+DeroNAZlDLBm+HBptsxYxiKa7he0jy6q6SNw/2OmPkkAupN2r9msjblkzX
j7v9bELlsKq9p1E95c+7rgEH9wauRoodKfxnXWf20zN7LjWBYdKtrS8yxPJxKsnbk+AEM7htnqV+
bJ6HX6upP2UnXDbWpwsUsXJzW5stxWl0mJdVmY70rzn2IgGb+YfzGZdWO+HfMgIB4ujNiBRYxB6Y
VelUPnOuw/GzRfmrHMIhJtDMhNvCjMKcUQRP+0Rzd1N5Sk9C8wIKIKTZ8y7AzzowLenq0XlQRVge
E8n2Xb2vcPMmix/U/zRPB+jMOBV/D0ib4RqeburgeX6+lK5WUJ9F1HRPL3RyQmj6r1dkrLv9WPS1
+S9EcDAXHB3VqNfCzT5ypvBuehjn7DHDMi0B7UoLFRpb2ykUF7FPxhHenWr05GR98qkLDOuUqty2
2Y6nuvvXLc9TxGDNnwb5Rv1NLiYUifhfz8T6Tp/CiwH5x/tgKQXBYzyj9++1vpP8GnZ2Pw1o6Egm
j/BvJ/EDcIYJBzs6EzeCx3uJWtkSMX1YQUXHigdDxhRhSbXfuf80uEULlvMaSZIopgimuVhkDJkm
cGwWLrQUeo9u22TabixyEeYomknZeDgvpSZ6OTdDxmFR/Tek5D0WdyKz62Vo6papiBL/jW2M650m
TC98StRVgFeXZefdQ8GKHn1M66UMOUwv7XXiNmILQapaak/sBrPUKeO0/jWxRB0qVDQGQq7No3Qh
54eQw3DEFh9FLXyrt9B0JJnOlra5uS01iFEMK5nRJdVytg2dkL2Cmm/PFDHyqDjWuggtLC8OrNDb
heIIcF3tWZ1lpZ4mPM+HYQOIClrzLftjwQih6FsGkk3xmxgfpuS1Fyme+I/VlWR6L+Ry1ZskB6zo
PLo8Q5VTTowyvtx3R7xfaMwiriALuY5ElbuOdCLRTNbxi59rTzQcd/EJKyAPLCkaxxA9BAk2+kaZ
waq+N3ZsHVOmh+2rWM2voIYAjIzV3dXfuMLu9xTBtbDW52ig6tTW3sQrpyx4EBH5qUzMANt0G8ge
3EMS1sx4gi1hphzbpAd4KY7mq2AEZRO26rNplV2pf8Kng9ymXj6y27U6Ebj9Y4lEaHCgWS/Eeddd
bWEvKLND1h6Dqx5QGiFsJMVjOWX7WN+gifaiSOASdt55I9pNr6zxQoTe6WN3i7R3AN6h2Is2FJ98
argq1pmLWwKx5A491pHEOyTllCEOvNoqyZgKAuhr8q4/0iltta5773ZnZwd5gQAVoyGJMiugeY2v
rVvOE3GG9hciZ7/tdKSecIb+C3ncj3fkHTzxSZ6BZvcSu18LgRmX6yGK+G41ZkSlFga+Qb00ucbD
iNdTLR5qyd/I+2n4vFsODpT3Bf2f/m8iJ7U3ceBqwf7fi+r69ZvmLJkdBHM0FPXI814l88ldaphy
/HoQ1ZKFknmgWJcxZRGKrnnudEfLJEK0it+EdJdEMWLzTl18r7T2t3Xbp//ke76G6rsRHFoUqN+D
UQUJknkFkJyzHyfGQi1LT4PtNor6QMvx0yqx8WABWVDUK95jxsnLxrHGAYAfquG+xHKdUP71nEam
EufSN/WyRYlkFpw2xJrtcQywTJgXP27613swytoHNHZPWgGMg6h3gxwp3XbiN43r4OkLorOw85l8
By83G62k/1pffDi2RwPdy4AxSUARdZGUPNGAVKTfDb2tU9Rl//IE4ltYyUVW/1GC0xMDOkVJItDJ
f5LSQErXNJjYgqE/Vxh+yXcrjosdTXkkoThrq9Isj4RwWJW4DsUCUqaN4RjOIY4lIIke10rgF6Eo
cZ46trfVvKmDq5mDKzJcddFvJOMzg36YbVHQpwHbbmrbAcVPzkHUSN3JwKN/J5haPr+pzIIB9f+i
kS5myHK2fJ0jZabuPbU3PK7qd6i51P747GoXSDreB2scV0QOBfY+x0kVqGy5l8JnmhM8J45h0SNI
sQkT2nIa+3tlDV6T/kBtrBTk0lW2WNAYPG14RHQt8dilhZ3+DJZe6ak1dMWN115fL+hA9HPbGE1P
kal0ZhRMWcRmM9glXv6xK7iD76mOIkFnS4Aw8P8yxVuDIPWMlrS4E6+uMm/p3M9+MM9qOcuRg88b
c65Qv/kaLVZxdHXvJNKsSR9mZPYiKxUiZcP4uR6BZaR9X0bCMso5j+rCbNCWp1AWnX8hN6VE2OlK
UZXq60gor9iaa5Wowo5tJqwkwJzEYaJyVTmINPfkjbvI4UpYYgfnrbajQURyqLZHWvADPt0Hv6dj
AvRyYEDMJc95EKQH0TERS8dsCB4etmXsfUqqUBS0QcezKeCHu8T/5S/YQgPzZA0fIh6zeka4woxx
tc3xfxurR/ffSLYpCMhowartr/xkuJakk06iy8LjQtQNL6tpeBu6Vop3V/kr6bYCmaIMZIDo9DV7
ExEvCoVzeLIIZnVTM0hfAfqBJM9VU1cN44i8LZQraXoeQC1IVFwDAh0L5uEhc62tstX18pB9xZS3
AbAmF2HEMEr/8M7+HvxaS1m8r643Y2SzQN2cJf2kJRRH5Dmy8YIxUxMPsRvNciWgHCSPuFcDy7vI
hgHhNokNz2eBsq+s/2GI3vfvepBfWt9uN8Oo0UZVimK4P/3ci5oDTOgKG60HAebrHa5DFSzJaUrr
9snUmN1tgFPG3aA/TfdKtps7uM1HPiQg+6zZkpBVJYEwiRfySIeERKHov4RqEaUfIoy9dJ2UHRzb
ZE+uYjiGOVB/D3JXbgD/OIPvn5XEH2RfIfBE2vdZ+XfWG1OKzg0AVa8DD+6Ad5QBd6nTDdBVBHDN
s3EXQeq3kmMVmFqQjj9KQTw7N3zjD87MszJqQ+ws9jLAkIyGQRkYabANMfZNVOr0C9I6DAzcujFy
vg4X4SSfDm8HnXMXonjmoAqfulHSbicWFKICdmCDomaA5zcoB50tgj2DkjaFD/N/2gHMahWBK0l7
yFPKGjHikdNTsZtZ/otRU2PWShUu+HqEJwjWj2QLkCI4KO0aAK0KFCPRJnQ1Zblx53/RR1kIVTME
dl8kq90EAW0bHSMHPC/Z4ikrk+ghdZ7GNO7l8Eb0r3xlv2vlr8jpMMFjFQPXrS2eq5xj6nUqCHBV
s41pmElvtmAaf1iv6MI9KAgckqq3MN8zDHoZht/Wu0kl/ICskPDc5zqCrvLCfmPraTFQE4Ecpxbw
IwTcfPoGWqQ9EAL6CdggOtNatQpUzMz5PY1wHHFNkEcW7BuZltuwNthTQfkFAJb45kPKhmF+w+0O
t7Ykzo6pijTG0rydx9uO0tVuEu2zKkXmnemVoGc8Qw+zXAg8zpmqBDNZCITxY2oaxM4ozPmdeDBv
nMPsrIxIZpae+cSANyayv+geyBMQr3JLewiCqUdehsiHH2yAi4/nhoTnp9qJJ8mKsgCW4Go/gja2
K8EzxB+h7f5R5MTIMuw2YUUqZ2VluMvMSDHZEYf6jzzoXH6xM4JL8qreDCGRSF2msopUU8RmQum5
mdN2l+4zLhj+ma4ut1njj1hC/QDpaxjs9Rex84qgHn1nZzh1tK37JQH36h9gYCAGVaCSgvMP4w0Z
itE+xvG8r88zD+ZfDcmS0mNKp5Pu8ue9PfJtjRQdWfuHw9nxX3vKsMKm9ewENZRzEbk9CZLn0h4y
g7Mg8aPjmgcA0aqxYxpzbUINV+F4muiuspeNSanjw2yFENIQO8Pv9Bdasl2QrgtLadhFyV+Nqd0a
Ju+5aRd+Gzs+33Oy5RWYWa8KkQAg3uhDQXMdbcLim0+RlhPEG+AFMCgGUST2UPwHy7FbEJwwyWgk
SsOfXIemio8O838H7RGUJRKrjG/eVljepsvWEYpW6Zy+RyRSu1yUICNYCuQXRGrku/Ppi//Jnwid
vkSpQhkd/kNMlJHC75aG/uUwMWb2yWt6d7EM2z3WQSvevCGxghPxRPhPf0dRcwH3bxl+9F/12lq4
DI1YVt8BgGiMc40jZnuIdOFxtI9mGozcuFnfP9xj4YR60NEZdQAYcsnnX2Ao7OKrd8EaaWzSwy+7
eyQRHi+14tG6qWRyml68j0cFy/RVakGNDBgekqnDOkj569NG2TRLWjWhQej8dco1o6TSzBW7r+DI
SY2fSWgr1zV7Ly+5W0CiIVeM6lHjN+aspTHbLYxCR+1Ly55u16mWsdOPIC/XjiyYXvsOsDOJSooM
3fZfZ0BMlqWtxNw7TJeQ8xjvaMegFyTlxWXrQdkxeCTsG7mZFZqjEKqE/u9Z5ak9gc++UNJ95v15
6uANMomkfobFZ+2AJhAUI077os+W0iyfTjXU7Oe6+UOptJqHRPKpOLOA271QXGPxbMTn49RT3wFq
kZIwUaAJhv9irz7uABZTCksDLUQ0a9w868LD4tWUPwDDJBYK2wx8iCbHfzJt5eTanYdJIpP8/oxM
eVOYOSiUzpD8GpI5LOLB1SzX6SBGeJeZ8Iuhnd1NhUQMcqk519Hc3DLZlTI1Lw/sGU1Zj3RIAIAd
js4xtKIENpLbEAwik2UV/CsC5gc8L6WSRZklDe8DXQfq9DmM7S+vKen/izQG+pyL98/dTChmUK/+
uR168M2O09tPVfpCB85yISumdE0Ikg1yGTaI87X9tr2Mb0Oaqd8bBh538m8qRbfmaizdqn42c7ft
+K5e+xWhPu1c6xHUhUC0CHRoS0fT+XNl2VhsOVG1EwCpDAK8wRbHfOWFi8pSUraY3UJ5/83Ri101
xLzIeIMEIOrjVwbT96s+K/Sci6BZPKYnumMZ39yaxeeXMMgasd1tJZgPT/rw7PEVJzqYMiIfRueO
rSvWUHIPbWI6SCNlviulo4tK6GNsFJzUlII1lgswHLf6xgLie4wdnFbxqusfZAOlTLZ1mKMS3GeF
EZ4VhraMezBoJ5qFAiFFOG3B7rhePBEZkDvjThuIOUfiHzXRHpjoCi+Eolv5tbYizsJDuEUYcpEe
2piAM2TlhqKFnrnipO60vEkRjtVZNkd1BdSCZ1WAcTnC+vpIAMYHcX143eVaot0R80Rf66sQZXWT
z26MDqRZ4CdJsRN5a/sLqggcJ79dzfr5oJTwI8lpwNAxnjjxxHLumTIyzmYtL2GEgi1Am6t4fOpq
vQjSV1WhGcIfoOAiI/2zMEEaOG+iZqd96aFly0XmugaP82dkBsYEPcpyQDubFJ9C/UaK/+oCtr/P
LSKmHBG4GcC17/AC630O++x+50oxt5dpxrmyGiWj99wYdRLwKkUKj7lliuA25eie0HNEeQEHCXbW
UDd5BZ8U4RiXhEaKOrwG/39NVeouxKWSTvkCSMOlcoWr6aWA5CvSldZ/XAz0DAJ6D4UsMcN3d7Rf
QK8t4ACUEgOachYb+agfR+1QDdmc6WMb+IUaTFbUcbzL5R+NL3U8mMtAYhGh7ZCIMVQYjy47s8uf
3c+HpSkpKkuynGqY5DOx6h4Y3nP6hPhnzcrkZ+eesv2IxYOcBuoXJr5HlCXZkeHpowZMP5XpbRMk
HwYgE3e9r5OjJ4Lx8PgQj7+0mX5yqHWEHiiMHHzFKGp0THoBO9cL0kRb1hlSaNks9M83D8QjPt1o
d8Z2l8MDAYMMfz0+gGwh/EquCkt4E5skXx3nRSm/+tE6/ERCu+IZRoKs2hrOmKjB2MrS16Lsnz/C
D2sqFTj20APZRkdA73PAGD/wYNgbxSSvI5fVXS1G6DmmFn7pOr8KDChTP8neigJtmDrKSvf5nLEa
medfe8d9wEwRLfOFuv6PGQzkuTZw//HljQZ/GQ/igMgn+Z7lgvlqbrT+Hk+L8zCW0NCA9wDx78j1
OQYzlygid40gJk4xQRPl9G7z7gH3wessZLaqY7+v1TRHOmbQI1V7P+ctB3k2eDy4QJyqJG/QsTUR
bGE7HE/cChwpIC/QTnGUYZPbzTBIZOu38ibAWb7abLEnKCC0edmx9bDCnkctuuyzBq6Z+WQzNOB+
qLlksk9ezz5sEhR58Ac6D8F6EcsUvD6MVlM+xh1Y4vxa7ZP7/wiwesJvRV6S737RbOcY7k1vKdww
lgTb3UoihIcoLtdk5KiBM2345KSghfoKJVcqt0pOLpHtOC1P2rLo45Yg9CSjsGzrIhvs/ZbyvQnq
NOxW3jdHQPIrqnm2wdZEAI4Zs0GncQUenHWOVrgKktx84Xmd2hv5JluWEPSq3tKtHs394MBZjT5c
NYP4Iha+cR12um7+2MGSCiZvqpdesou+h5WYbpzlYUVgo3k9QDouEfTGISjyG0eC7Q0UW08gj06g
VyXEyzDBHPkgJsyTv+uO5eoRwLDB2fPQws4WRmnlCnAw3NJn4fayf5nXztQvVnb+iUH+3RkQCLxT
CHqzwYHVAGLWE6TtnqFJChTWRPZv/wpYwJbtlJ89Qs5xOyPBySUu7dzZxOanOCazZoDi6IRK8PYc
yhXwHX8y4RgX8C8X77WMy7ix1fzm8lTuMjWt74H0b2w0E52OTFPVxL7wiARgAwR7ztkOq5m788xd
aeEFquAGxLdXgmW2xjWmFmTHsPH13b1peTZDO8tkNhO6oyEr/rbxpSMlMllVS+0RV4NViCZ2QMgL
uyAdRa5EYw6hlvdiuOgur5BQmrrYlMuFk/5F5jeH1Hpzc/LR6zs2XEgA8JILVG1QzddfTPLrawyK
8md7IhogcuLislW2p0D2wdFxd7YIHzrDC2/pCauUwzoNkwMkjECfXifhEjw2MUC3x+K333QfegmW
CURicnzLeaVPVD8VMiWAxykcWW0R3oQAqHebfyG3XH8HkhMnBDRceVQKHtvtPq/q0nlWhJGvfEox
lo8ydlil6E+H4Ne5yLmiNBrTfWumolScVC8dSuMSbe8YBZJx8UUPzQJF638H0X4EE7M6SRawDs9Z
ZiprqXV4dDM3/DwCGHmuc/zAFKWFOjkaql25G5GzvPP1MfILyGIWEBDcFZJHcXpzInGcBwugBZWk
GYJlJAsA23XC8jsGJHWZqf7SBSUPHUtvCQ9LHOkMgm0YJ777CytSNrbLjb2gBwA5gf08MHUw8dqp
jxXVF3T85xbqnn043Yk9CXbTy55+3zz3cGInqqtyqv9y2zTlfnwID2O9K3EyvW+7K7LEWuXisWoz
gUoqUILHCeQXa5yBTQi76Mj4SMVIkH/ZV5tVpjUHK5dL2BsFNBNHvMUXFIuwAxldcq9FDI31zDd0
GTqTwDe0L7wJ/YC3QdRQ8k73An9kvgZsifTkHxhjkSBfWs7kj5fXcUk5zsbQePLbKMYq4PdDfExp
5bTdiG7kFjbgIEc6PhjEEYrmk3Ca59Ss60j3cQAz7CbsXQ1nNjR7Qxv1ba0YIP+C1tl67FcU7aox
EsJCv/AkV3tWbrStdkxAhIRbeVatbEa3J9GnCISuYjD4pp6+hYpSa4wIsbbNBeN9t2/Y14W/uWwc
ypBwKHHeU+Tai8G0jN/uXSHgRXqU/Ge6PIshmQ9xKTtiOxb3U5uSC+F6oMd1Jjkv6F9OqK+/jDO7
sE5gkix2QDNP6wYGqJBcLxiYzJwzRc6HsAJ505yTIOzxkC3ER8lyNDZ5WgD8/NtmzRR1BmDuA10K
EuNqKzG+3W4CMFtoXqhS7pwrenbDezXcVN4oAjjheVbGd7Jv2x1rzIPGgUuGn7rdc/+TGHNDsQM7
Cr/MeOBfTcKGLSsyjRJkZVSgNGv/oTin0kpoPvrus3uevUleplmGE9QrjEvAT/tnQPOm7NT36jeY
rcKLokOR7au9js0cv6erEGN3hit0Y4Z8DPjmVUD249P3tOKIW9LMTUI89x0c2VfJ/EsSn3qMrrYq
Vq9SaXPpDbnyG034oSYtTszV0PdJRIjOCkMtNuU2lFM06PNgWPt2blGP1sW6gPVts4UQsHQmVRd3
qZCjOS4oDdKdGvUVIlazRezU6ZL2feer/F3qBSMs+tO8G5RePgvPwehj/WUEXddPOC/OeqZR2/sy
tDrdn4fZILMt1Nc0KsdBt09r8/2/9IwOYJgNjd8RuAoUGyIgW3gsNo3jqC6ItQs0FZfVKCVKt7BM
N206Ea8/itfeHf2r1BbVghVswqONsv8tAK6xoSVFF0GItQOFLiWoeLy5izVJSofT1heE1V7ZZPhu
UwE4yBH9pzuLRjgDeRe6lbtfgL1ajP32ON5V+d+MhFo7L7E/nnAtMjsa9P28Tua9Uc2oPAKk19Fj
swXM7ADqSXkDq5iqVKh0KXJmZZtfLgT/8Ub0ohNZssQEn1TQQRo9OPms6N8lLbjiiCw1OkIziepd
qUR3GMy6IR+K+wgIl9aKnFfbwkyYtBpJ4gTcMr7mm9jHi4bI/jVmmavFYj66Xoffj9wbN7LY0/jt
tPqWWoO0+UI0EF/iHUgUwxhBSShPttcdnjlXICdEdhbxfbRwNwHtRD4fdTuEkCdZ6P7Rx4L8spTK
B7BYS8xkmvnrWaPDIK7xjJ4LUFNOTCBYo3/l2vIYmmeckI9RAnlKJTJoiETV4aKng5O9YThP13Y2
+I4XQ5banf8MpsJxoGe47MjoOwPThb7Os27BnvuxR0O2L72Y6ZbqmregWoKW8zBZV7MePeTUKeCH
7+O87OJ9TkkwRyHUNwqzyeN3zNUjCCjFt5ZuQ5JKxyErk1abli04tCDnGxk2kl4DXNUlOxRHwHqB
XyjqHGagIZTzf7GNkXSfNwKEGwbPrmXU8uznmfussWIacwXcavkUpxmrYyidwTpOzPTTXi4JetUe
U385hw2kWlejfHYUK2+3L1VPEl3uMsjJgPbCci0zvCLtZiz82XygmCYnSd4seM+9Mh6CJLFdQGK4
EustbfPnj8bfrmVBiMNYvbGwKzPoz9yD/uTR7zJD4uFD3sn9BzPwpkvd5kzxz02e1ZpHAtqOGUOE
NAXnih5zSpO6KMUY36+THmhUMThhqTjUR1Ej2PimQl4KLtLtGKaXFrMksFDIjDjmj4uIqzskbScZ
4TSscX0BORlHYe+mP9oBRu5Q+ZaflJEZhOgluoxE+muj+7/VFMLIP8acO94ngt4LaIt1i+ebJu+3
Ign0uBNJ9IxZfE98n0Yze6aEDWwltiiLrTdbylbh7qxOGKIDyfnUMlP7qqiDzluQglEXs0x3L3/r
iRwqfrcqfA4Uq8eO3IMY24XmaixsUSgiQA+N9rE9Xcdk5ept2XnFSKF3uAo+oWLQgkA3zLzRPdwm
165pMkIIht/JQJUMES8/DhvOUB3QsKuPHi6+yujR6NtTyBJjGWNAQkbJRRzFaVVE70lXJFrB3ze9
P6mv0WKsrkPGaiKPZi5tRlmgPHlq99YlnVia5m9kBf7FU0oEBHVmtTj5BKMcwh0l4nxlRXOCjEAH
4j2bp/tC0yQdJrtnPoJZLLP95xNqo9WMEPaM+x6hQE6iYbmL7ro4EwdTeiFSXz5vTcqIo/03oZDk
alWCcSADcXlLoFWlKCWs9ZP1o4TUi/LkS80oihVGfZkbZq9DulXdaftYE4gKqYQK38n7WmAc3SP0
/NTr6hluyIBW5HRKrDjOxWuZVSgtdJtGnOzv7FOYj+inXM+AovDt3pdJa0jXehZltb82TMFLOma6
qtgGeYtTISRDiyvz0VdRfUKSgpzrsXH5HH70w0F64JTBrKD0JK6ncS+acBn6s5gbDeHQCDzfjEkk
/h1bjnsBz22sV3O8jqy3g7d/9b0+/iAsPwdFPkd+agD6vZfOdYM40Nom5YSuFJlKg7tjwOeiUYM6
y1LIyia53R1K/XWDyM4t8DHx4jEhg5milCdMHkd498qwwyp2/pT4roMKlkzx2WPnyUt2SSM5SNJv
R0IPsvmwtSjG0AHL8r+Qcw+tatUMjTra6M153LQI7LoL5H5xhkwpUSpofi74wi1WINEIjxTbIjkx
G/MX/CAZ4sGVzGQT4k4dG8+c4qmCowkeBerkkbyEYqoXPFdwbY+x0HO9jekXoR+NzojfCulxsu8g
B23J+L2VJ4w6CDtRVN+vK7xzL4a2BF004ad9QK6KfzU2QXeDWhHEJ+QsrX60YsefS+37kmIzwGCP
sWJQI5i4hP738UGr5HN1Fc1AJ2/IJEmN5rULjnOINRiHbSuQOdnJVppH4qV42Tt3qH7uynlPbrbU
IJYGz+7CMsKzMydHcfGO96lQxooBTZI00xysxPgbtOSViteA/TvRQ9Dn48/N9E/ChQsAG4zb8sWZ
tzatvwVeZtfgzxBroiBUNXHHkhauhj0cXR3azHm8D3BMCJFtbRK5cc6LN8u1a8uVi6xeuKxyI0DX
A2Hmleqw5UIoQ2bqaAwERzuCwquoFfljpUtzozmsCmXLJ9v8rYmzGUfva35z0e0Z0CKMtCtvdYKR
9b4mCYmDaIBCYrTYEE1Qo/3Q8af4dnVdhfGvhtLaE4EHGRCIML2GBY7dq1EmS7ENFCyPdW2t3UHm
oZbK7oaoVLrUkigR4kaFVX1sWHWPAQFFOVXuzm2pF8w4h3bFs6M8eHkqh3K/NU0mrGBqEE6XGD6p
Q1wddNvcDHoLZj8fx6kKMOxlCkWYn18oOuQqwijEb8971YCgZIZ3riay922oUOFryy5oKMitdBjC
/v4+AXNweIsjZ8OX4pEqFwI9NEbPJat1XOluGUsZNteAS04RVgsJ7wh52x0hwjqvVaLyuA0yURB4
L1W/WuxXmI+G1WQ0U8Vu3DgrcamLpSbpXHIGyuHRGrJRO6ENfVZSY6osvGHrHImWJ/9QWUBbN9gq
2LYL4E6Nj4K4BYZslPQCYZVPjR1tKkTBFVnXi9VTpw1F9/Tn+Wb3oLp5oKeG8qhHI5uyjZ5QT1ac
O9wkUzV8M/DjV+KDARrBA/KspnWDfzZ4Pn3P5Bq056sF4VsWW1xvWJ3xoRQlHpPxaXuovofm0KHr
/BqIIAyeKh8pDngpm9+UxQQJHd96Fsa6RA0iW6kLOSjJa3A8mfKATuw0dcv/tzQdMJ0IWChEcTu5
B114cdf1NnNkpvVFqV5oLO+fZuLOeJvo14ux67kVDJEcf3RlJIBa0L+lwIMHNWqBG62Xvqwc4H/q
QLuZw4JGItkEvEoVOPHbjvUY8X2S4ZssmPikGJSsYGXc3krTFtmY3l6igLU22HjuExwI3UyuJ0FP
HqSYFOniSCCuhPXIMbJ311KAWeddrI/R0YIuQIBRlBsVXET20EOPHznFo/wDyPO6BOyAGP6O9bnb
koGYxdfY5xZlWML5ZI4ARJrAgp2E2SfqH4GqoUImjYW307kUDsCyn09RHBqUrJnmkqtxrtOvwPn4
CYlW56EJ9l/LYeIKejgHsAH+Y9EZywEFLcboG9iCa8XGE0h7rzpntfjFJfDHw+SPA3KudDZkcvsg
QUQABEb+lN+Yj9utsbaS4tC6fs6Dg0kRS5QKgMUdkzvspbW8kanFEtKrl4e9eflsvdDw4R6DCU0g
V/3+uoZb4RInbQd86441NMpim6KwXX37Ps+wVgFeNvXbMhzcGns4t7l//zf5MPjh4NKzwob5REZU
kNp8973TbigXdrf3R6Vq2QqvF3FtPjAGHjoYGMEnTHo5PM/ZiwMp2HNlFNcZpUjYMivG0TGgyz2b
wuRRZvn60NTdxKS/EFNztTWat6i4HALBnfVv+1lS2iDr1yiexaKPA/EK4bFoSqFsu5oNY06kMxVf
kSRhh3F0EkHgGvdg7swx9Sh+CJieJZCX+Ku5AF8HuRGIVWTiucWPl0VdqcgdcEXjKrCNsd/wno/d
Alhu0rL6KEDMGUZUVwV00km+PKCH3/8rJv9D5u7VqJisdsyvv/xFhWNOI1FIcdP2OLzUbg4za0Ql
9THxCoxDVqvStSPl8jUEAzb0iyY76TidghLnb47Me0ABqWzcrUW7+c/DghmlRKru6lKfoDs6n7Ga
ibbczXsGefAZ4ICxJ0m1cmLEUUNHBrNwu69R086VkYHT0vh0VljzZGQTztpBAzigNgVeuV2SumK3
N4CMwPqFRfvm/PwftlKgtqOLfyGn2EMTaQQrX/Nps1GpPHTjlhA6znI8H0KQAJhDtr7w4JiZmJB3
pRVYs/1PPcICommGVGIvaD7kg6xL84+5pPJWwVGeIIi7BjPpIJjjuWA10PAbBPn9ro5DaKP1x5Je
90HUnsk3Z9kr1ogrZU1sSrxCu8PpJqqowQNFojrJr6FUhkZm9y4Ilz3rLYihQDGEJyMd2ft/r1eC
uRbnvFjG6m66e/0BARWjkPpQ8bvN+e2eodIOmCT0wvImvj8ehon38PLi+AV2OxNqc1vmr3JtMB2Z
Am7A8/X7IgMsHhwezbMGtggQr3MyzST1+APO6y3TlwiZJjSvFl45EYgxN5Z7mzt60DVIZAIiZEy5
18a8XQqfKLco4uGBBXB6EqaSSvabM1IuC5tnthTkh+zFQRNt0ebCkTjdQJZo/DpPguzapBXPrDdw
/flR5raEFFzdeZe89kILnnHFZr53vw5YStxifAgofNbOL73ipdXn4MTK1I1/oMdp+tk3Zln9skl8
+aJine20GzzK/FhMfSJE6H6mGKalwxnUxFe1ECNZjytzHvD/fEf0XVBFJtiwprcCTxTEfoQZzR98
sqMtCDcAN43pOhlgpPC7qd1eeWNHIvwatl6E4lifnLzxE8BtzjJRXGWBFqlev+MtMVSQeSTbagXm
c5kM3Aa19wkec8VfuEWPaaWgSGyA+QmxF/wB8dz0FeQqDdlSN2Jm1FbQ0ymaPzKJjuk7AAAJ9N/n
1K7GqoLidJbI77h9uuopXS4YwOrIS5jFusWZ3Bzwttl5HkIwkKTTWdBXbQIv9CIyqFZxqboKvrJF
eFCSqmpCnRVXTyjF2qTz4wo4adhYk82QJxgr936RsWMl4ApxJG/rIKX66FNDt/tFItr8IkDlnkUA
nbk5ULlQnqCPFgamWWWSmpjtM7fOYVNd/nPcL7xZyKc30+0Rjgs1eXJQ64JKGQo6irwrndH5rtLc
1DawgoFIqxk3BfCCUAjK5nC0QmSw8AoGv0JjYIWsZCoN+zSuYxj9/B4ZP27JwhOaIM+Oy6WwyJFt
BYlXwmfSMfCkrEHp9A+uaaJDdiftBNNN2lBPjjI3uYy+p5s0KR9ftkT82OhesBD2tzUl+U5ZGTP2
Fz4xqQ4Azn3ZVs3Q7REekJrD2Zr/obGTVXKf2lMCTfnV1/MNY/8oBLSIcD6F0xsYe5FElhUG3b/h
fKMssO+ZhFEN2eKotT714tgzhWrGNIFqCYHbUTUKeg0g9Tx4xKvr0rRh6ZduM2hpzReRE6cZVHKg
/3vLFSrlmSLtphRaZcCShr+Bwmtso9qD9+TUley4USPwz1LLsGs3DHT8ftKuAxrRF6bwB24rzzA5
+MvyqNJ7rq3oU1TpzHzmoU1S0lwchWjnsoWoI3WxkT2wq4sEuAk3BthUqlRUz9uqJgY2gY2xrPTq
zWG9e1tScBS5e3EQ1iszHGTZuZuWhEPuVEo/SO6LBFydAU+11SlzWTZlCuI9+fbfquIdcHtuGiGh
R5bDZYYCnkbQuRuv7j8FErFdPNrI4sb68aYQAl/cUC3Q+OmITTgR5QPd95rbFpazIkEdDcRMvLdt
pe+dhaHhCs1YwhzMCg9nkl4ecERCgcwy5roxHuP0dSGRUmD1n9f7Gt5YfYeZrFCCZpwwhjAq6+i6
mqnVTj/88dKG2IcMg3p1g78BszLreSBZurq+0NGzdSnK763C7lmsNVD/HH557VZ2kKDTkn29GMCx
qj2EBV2mCksGcnOwhQxh0C2lwMX6p4o/utGJL2KMJYVruTgIKbq9D4IlX2p4KB9gy9cW5jjP5vxR
A1yjohrjpUqsqyUbzJdzRttjw+isLt+xPXf8IuG93SkY1NDyJDd/ByPc+k4ww9wewxA+xUIAmi4R
g67KzF/zZtxpO49BUUrAJivpoHcItSDAEjueKUaRw6+MzBVvWv2uFMf3weQaH5m0l/45nBRJdbBP
p/3xp6ru4CGD45ixHKOUhqxXFnw/GLBxTAbPjo504g9AIfJOXimoSIJoDJ/Aj++3AdGS3kOhQxho
EcTSksdVhhhMfAOe8noetvPGUSRxpkbwlrr/9dhU7HRwtb+bUygGirysimnMLthsxwGsx6bWA80n
DmD11nmUuFsIXVQpgXHIepFtYbFMEqn24EAqoD7AVec/+vYf18MmSgsSP9nP/tfiGRXh5TMMQ5Hw
mrVHHCanAZ4t9S7ieicoN4bV1p/2UbUIdshi3I5YiOXzWGesbArO7hXMF1gumyG8g15zX3Xi5+dj
y1cfyAOizS63bWCVGDhutSwegULUEC8vYmCVIlI4Po9Mmu0CQ9qX7sZa5OVk5+man93daL74fkiv
Xhih6oSguxQ6SWb+30yg3yXA/Nuh2W9+YT61o3ue0M7WwX8Kb5xP0EP1WoyoFO2YUOQ9NjWERxvv
L5Qot6iyu3dIrARiFjA58kYc2Mwk7KeCksOwkWD4IQskPI0/3b+Fa2muKE7j4NcGQ+9DVc2pLvDa
RnX5hHKVN7XfvwPZz4O3pFuXaudRSAlTWupKUb5qE5RqAkPI3Y+ZYk6v5elPJ3MwzAJMstbaf1rZ
/RqCZT1ixs5AOdaMRBrRKd2CSYvMkSypyQyE5fUkMaKP+MJOjgOGT6jap5jKdjrVqYznXtCUKryA
+IHlZhqyk1YsezBx5x+GzH+nXuVnXsCBHLSngf013qNndytaV4kg+Av07mn9WomClxuyAZYpdsWJ
Wcwvxgv6eBVr27Cq0z+gR55/JZ08Xz08FzW24oRWhrou8iIVzf04ZqYr6XuZzJozfyuoi/rgrQDQ
k3MAZzEYZAhZZTbxRH4Em95Mg98CoB7R8ZFqKQ5hNRKRqRJCT+Cqw7E+3jDdm1QqOvMgvlCbyHes
2X/VtKUZrhwpJVZ+CEWl0Cz3PTGgr0Zd+/grmlc+XV1mc5XL0JuAKEejYzLrLIvyBxp2IO7EAcdM
4RmDWXUGka6CTu7VN0zihfGMT1qKJ93GL/IMuOaVU1PJ20szFfz+ZhBIwIswb6JfPxtBtyIwtQ2o
TtfBSO6DJrz6BJvcnd76tWaS2ao4TTqHAUbaR4J3GQrjM0/wn+qYW5Di9AR/Ct8o0AOtiM9HTOgv
FE7U6i7an1jJHG8bHHlMN0tqf4ZgM+MezMFpnjiMH+aRHiFy9U891DPpu7ZoUsHoz/9qgzS78hAa
5h3AGY6pDcZfX6fwmXqJ7Y/uQP2/Itknk2uiN4J5wMv+wH0x/n3ctCjc6+buSveJ2LXS1o6s8/hA
Frb8hzp3pJwcAUDF8Jn2ohUWHo2hCRW2MnZdudkNONphSlyMz9Mrb5upDVVo5lkm8G6ot5oRzc+V
ZXr6/03PbeB4PBEyfG3zCFIFYs0Mk+6Wuz+N1IW7kmgmVk1CyEbTqCnRZGYlBARa4xHER3KiTrIJ
nn0TfnjqCGf2/lrsxBGiwX4YhpNJ1+dbgOn2Y0g6oObGzGTQdsx9iZUexHZLRsLi2U7sl3K1jKR6
G+BoCYyq8DJH26TTPE++CnMJruzUwDNefQoNhaCJPnRrwvCnGHkwBPxrALeCKQnx9a5U9uZBgmU7
ff5ptn47ZYI4x9sEBUjyQwIXBznB5jVjOWIC/as/ldeDa4vU/82ihu7q38suJkCMtPrGx5EiVotS
7EefXzn1yqHgklUMjzIU/KqSgPzc11CUHdyjjkqBJpJRx+iLGybM3CU7BIbr9O6+0RcwS0U3WtnK
KWZSbnwf3ZZBMZNmVCna0ZaPgpbGuLwKRFCAdS+zGG7tixvWMbqNPY1YBQ9bLFeAu9CSPVrQYu6z
CVdm0fWuO0cMtsdTA4c7pZIzOoFdEsj8y967xpOErsyaOUzzWlixXK1xMBWfCXQHgmn58dpsF69+
XdcyBIZtuvy2Eh80Urw6lM8o6Jq20v2cKLDWMbTxWSZk9/zhOsSR4RX87eZ/Dq+ElqjsR7pPfbNP
u/JgDSa6NO67KQ6P/Gt6JZpGHva+jNHzFPMw0K9q72fighp2xUu6u+wwPBobt3xaGbqsMypw28B9
VO1wilHjem3OrhJKlX0svgCBHxi3jhTTVmg2E2JQZOkZQr5EW0jhg/+veu0ggH8btBIO40RZTpdO
H6HBo5RCcHboAsrxW54krjGPiGsU1wjC5zaMZdLFv9MgQeMlO6ZROjXWmUwVoWc9JmqEcm3VNXVa
kaBIHYtQIlRgolAQeyF/enb7K2dUOq2BKmshfl7SCb9kGrtXgNUn+ul9oMOweylHFg9ChiCQNGnE
KQqWkpRmqDRowyJWlvt3++z39wYxQCnIFdw69dbclyc563hdRsLODr80hDNBWMIL6tP4c0tnztD9
HoHsqykuvDrW5KMDX+/CNFp5VM95WCikisjVeYr1ei1hLjGtNgEBVfMhrvYEu1W0Nymd+W7/FwKr
36GukLZAF6s1ySQJEYNQ+ee4VO0w9ZVrkaGKpYd3E10CK1pC2lV8VfmV4USZcoR1RFeo7bm+13WX
SFM9ogbngD4MqmKwHtYaZRC375H/kL96ltChj+AckAic775AUT3yNzk7BeR9RUEeetma917qp7zm
KwegZiDdKdX90MMqw6YKHJB8tCGZodQoGKYd1yGxgCa2ektCGzWmCOAh1gzUT+etr5O0z3PjsTOi
jXRU+UpFPcydCCtk3V1wLP6zPhR2bIKjuKMja+A5VkQIBVDWJEOrDTMHtP9WZccQ1BQzIMoYok/l
mvHQZtLsLdBc9f1zDBhyKfs/fsEDrvADdMJZ1RdOkaTliPvP5strVgz2k2nGnzlzJeBh5SLRBdqn
+vuzx7PSBU4hJDrWA7sqRKgzx/MTwXEkiveLaXbNtgXVcIVyQVUbkFSJc2l9mO84Rnq25I0NQcKt
XchIEFufI0wbCjEhhaQJ9hBklet2q4WZHFQCWOtRzkXxBTdB5QJfNHybKQwVoogDECD+iD/LcLwo
Rjb2clY/obclip2Azm+R4HExO8UOlPmM42oqGMOorqnRV6CrbmcweMs3jLnBAF+xAn6HBxM4juKE
gJDyPm6HL+eVCsh9XDvy6243uQMOh8cMboNRVwxiIxj9ToixJ9E/JaDBA12T4FoOGQrvBph/2xNp
0W7QEqWV79ag7bURaRzIV6N6ZQ1TfzWOVa9q45rqzYWb7/ebZMzEOqH0oUG9IvrjE2FOw00rODbP
L6tlQD7eoW1Jb+1a9Gy/hTJR/J96Mze/Jj4e5I6V4xj2U19Tocy6XhUPTAiS2TeycK2g+HD1YTki
bvGkm+FyLloe0dG4CwTAe2SNCI6y0uI/Sv2tAM7CIKFN16gX7uVmZAhmQsI2rpLhvjaUzW3Kx+Cd
8RTcOtU+Ja4GGmnKZk4kFrB1paVjCgT0G3gJviOPgxwzZV8QkO6VFOotWRz+slEknLf0tYPV+6vS
OtYoKxpLh6AAoNMTjq/+q/EBEfujZLnpcvE24SKI3Cfc2rs1WwguW5GWmtYFeO2wHfHRaG7blDzm
fl369ovKDp3qde5vhcylDRIoih4SQdk4+JXGSzfoAS8L79pgiQs6WpAdQqbXeZ+Vh8b9tLWYYWD5
Y05B3CoobdGWAVfvtUNScnkl6vAG0T5X+gjYbkzqawUPF02n9+T04LSCXs+juzeZqYkqX6Y3XcID
P1YeqIw+RYLsOJxXF45rJbbFOVifFPeviRF8XiqNgMeU7m1Uxhm4ATzHAK1CJlhVeXQHrQgMWp0F
1Ho0+a1GfKBqTHluxXWOt+WYhNgyYgZVJJjZhIkZYyd6t2kMfmDZIuopPvvheP/1ghXPljBXi6TD
eFCzIRI7S+/7LL13mqDRb17rgzNP71PhmDXlpxRBWoUa3L5NTsobB+/kO64W9zIVIy6gKfn7cD2N
4H3gJdqYrQUiHu6cGL0lvexYj4UFMpGHv1BPpZX7zOMZWwURoBXGi/PiMraK7G2uonvX+fPmhfbZ
jYjpV/4t/bnUn5A/TGGBChCE6iwSWXwvrQUIa5csWM1rlZDXiBTe9zbFzJZXpa9ivJ2cXVTagQ3F
L2kdfwLeAAitiUg/9mE3jgr9QJzIDpeG3ky3cNsYeyi9aiIR97FAhXK6gkFb49jeDCNcEVZ1wHRL
xyBimryh8izUpWzeFRT8+4gSQgW1pAMtYZhzJzm8hqEyPnHotBhIaSkha2+0KBK1R0Ye02cp3s+J
8Xu6b9zPFGBygpyPtVGCHcjovGDHYBQ0pZNJKLZSH5Ia+oY5Tscze9bWAZLJJQC+ytBUa+03DeUr
QNTp0EXIXiLld8pOpk2m2abXsF86twkslorR4Vj6B1MREB9AwiWBhKfiKugTwCKGp7jJzfNOd1B+
hAB36Q++zVhVVePpV8FurYYpDmqKOTYHthUlMhWwv1jx4nQbdJ0JaCYTrlxm0jUnKQN3roX8NFbf
zGRSZ8DxzsyQTryoS6Pzazf2X4d1qp72sXIDvgFAQ1d45IpKmktObsQHT+v9G4F4oSuBUAkXMFFz
VWtw/1KyU+DEDppXXCXQ0MFuroT4zlohKoEauZKT73CEHrYU54Nrp1QjM+Zom1lzPN2JM+UMNMtg
dto45xCn5stRwVc5n1x8RLqkqZw0Ce9gx47N+xUcT/lVQwYVIdXG/bkEHzxAWT49gEU4CkxsalzJ
z4Sh7DH10B5vP8rxMtq157G2bdkP63+7lLZTbrSU+1jBW+ADAmrCCfeqrmU63zKTnxoF2Cx2LH+G
bejLE3qj7hUqHkR2k/1DjbBjmYXEzXtzYyFx3/ojiIJpBqjGgBOGxwItutAED3UZGCGzYwFcdW7q
OjRlyqPcs7pZzQSbfOHnJEqjW7QiBTtJFwUbllD1JSXk65InSF6bqC9FiRoJd2SvUk18JKolYcJe
cTduSoiTJhbuhFkci1hrsa6Q7uorfp6iVa6PNHdkIzcvlAyWELIbUNwBO1Z/UWIGSo01Bx/AXdg2
EmK1IbbTV2y2PnvdfdsYFo+4IPAja3ssEgkLx1EcX58GhEsFpDcx9NLnJA0RySWUNp+P7NR1ltQ6
Ghn+nfEsgWeBjtA0SFO1VPSpiLH2770Ly3MG2cQNPp77ntOsusKE/80Jb2Uuw7rQpJ7JGjahYzGH
2iwj7MqSu1XLCtaV+Yo2IzrEgbPUsTNG1NDxvwAZqF7aoVmWKN41uqEmWngxvg6zOJDBm0ttHuht
Byo5sdzYtSkpm1tVQ6qC9/kvWU0Q4TWNpv8HQbRHPCDdOWjWfLt7NuJ+jdgLKD1ZgqaQSCvqFhA8
by2ILxj/h7MHKlZnput874feFu6Pg6XxF2E064TW1MLjkvrWD+fossbd3IHmAID4sqMYkxaFpVC4
5kf/dY1LEamr29wpL47vBz8GgltyO7b5EwsnOwIGu5oL9ienwRL0aoZFi19Y+hbWIEwytkURTjir
J+mtjAFSdgRHvbWY1Uv1Z7OFPzYse9jWcf/+LTVQv5oaD9qjLvmEdbhR+qc9DpaQFmAptpq3Tycd
DvG8AZoLWY9BjwXFIv8694UglQLnCDeukzdgaWWVirr96P36hDCAu2gPl3TmQFfLZwWetcPicyq6
eJf/76CLmMfGmlRSPTGnIOn+kDeLO8A0/+zK504cSeWXtIUMZ8aE5nCtmfRPcOpF5FrJbYyvCDea
dO2O5HrbuFlM8+EexgfVzHdXay9O7DMfzxJ1DUQoZjt0UeyNHneTqf0fI3gi+x36X5+2xoCl5CPc
4OvfomlD3kZvljYYNLjCcaVMZmkxwmUAscDV5TpsqOBSsZJECIqm2YhObeP1zKS3fI3CDMi7ghCN
216XApTcuY77ezfHVP/aaaSruU+KNxPJJXM/jBCp8u2JYyAt85Lw4U7IQZa2AydnTsZAccsUFoY8
d5p20TS7MWbGmHWz2hpaTD3IcKDgrhcd6dUL27df7SmjYSy1wvF5wCS6SREQE673LMrtvpxufw+V
K+iZhbuUjspoCk/Kkl1c+P4eaPlnYD75XhROScosL9t987CmTa/Y+NuWYBBXrcUqy8SLxrFxvD+d
z0ql6knvHh0J8V99oi1njfsAYlWpLWbdlj0sssCCc3kXsE49y9arjyyPmGPR4lHz76yVIAMeJOmu
J5CYfXbX3LNechUDp7aYTEAH70YIR8TGcV++DcLwDxWxbsBCRrEKhn9T6vETqS2kvGihT07KbKUS
JNHr3bgbgzo7NBvf+WO0tWicMhKaAn6ZixakkptP1BgufJqQxUqqmT2+VBgKPOulilmj5h3LDuV1
dYBwUK4Du8NAJ/8AQJt8aC4f2H99Imtn+eEIIlwqPfNqNxBj5XGCQjWPPKdPJ8C2Ji//uewZShMq
fLDLnkxv4XpIhOMVgaKnLhHcEGl0PNCACIs7SQB/5Zjl/ZcZYzEss/nXvsCQvd9Zbza92j4h4fQT
TXBvA2NJwWYtJiRDSmRivc2lkcggA0GqIfminxU1gr3pPZV2F1pdpwvbtj4y89xp97Wglom3xrZ9
RYOcq/rgAyBv6dd5DswPi5lZh2ksDIy1+ocd6RDPx7laD93sRQswa/hmwBM/QMlxnHaYe6VXcgIM
YVAZtsP8PZYbp9Asf2jk7z+XbMK1d2sRIB09/6+dOLW/DZi2Yuq0+XUGweeMhSInwCuAGCYO3XKp
o9i4JY3rh7gDgWaH0qCHaeoKlDyA6S/q8TrWxy9tm0o4k97VpGpa0TDXF3cvI/RgsdEgsL75u1u9
DU5XZk5y1ZLrPquhcBqIS17CZ/0obmd5IP06Eja2Z5z5Et7+6trP4XBcFIKCqk1Y7YH/Nar4DwVf
U577go8Weer4Sx824nj0MiapZ58ORtSdLRszy+NP76kTi9goXqJnySde/VxL+mVlrtTrUnGu8MJg
pwPEY72Hkvo8BUnGaP99zjL/eypTHzW18f08RVT1fuPqRzSap8EKkDVeQHzQlXQXOYOabCdCIs+H
iMKDSjDu/qMbySCj7m9ZQXObOgetBryKrPdAOg8+4gXuBUNI9FUFIVxTfj8WoRuhzGyZMEunyxRl
TdoGl230dvBM27pPvZOrimdpk2WqLmkh37G2inS+2CFf6kBffeKYj0IVamPRTF6LMNrxL2QXzH/k
PQpVPSsVOlC3d68f0vmLZWz72T9U36VwzyYqVfEc1ZS+LOa1f69aIatWPyi4AKG39Pn27alSEt25
W6QhxhUM3UvDeOvIxda9PWCQrWcFdN0pDDA8JPMmDnMw54+Ko1O3bh6eOFlq9/MvNdshlzsN5ScM
o2pGpTA4DWtYwSPpWe+2gWn3uafhoi2bux8F5cEAcBjdgLpjNRQNl1x9o5Xx9gV4hFBTFAlKot57
mi2MOTRvMveCzbFBZl7QDEc7LYdzZcOOrCaMCxbe905yu/f24f7+dAT2kS0ozeMQNrXIUhdcJp2w
QVT8gnf1lWWB4yf39PsZkv6do95lplFOHlESf9ltP9Lg+peZLzhgklQxNWcO7GoNZx5fOzM1dgMX
NX4z081CFmcpw7EXTP4ilkK4ushfcblReWSKoRGtSFylMahN40OJM47hNptOE3wsQ6unuNIWqP7/
4Wwv6eEl3mvNrywzdJv4ctG5oiDMroDhsIOC36B5+ah68In0T37JTZqJ0aF0hxCJWrPREBpYP5wa
FyiU/3CMlSqpe4V16kb9cAPBemUPOHAOnRiiiD1/r7GMNkdn2IFBoFBCLI0TbI/Am48n5xaMwskz
qqJzIRg98sx4ZKU8ZP7ZD2uG1Fnfq1D6iVDvwV6PKXE4oVViQKw7dr0hQoyy2zet5cr1qZbA5bkI
My4dXc9D9imc2zNcbnHwrgyjn9Y4PzM7aE2n4RNr+VAnTpCF72wZivkPFYFmCmqtDChOUxUnFHiS
VgFfsGmxa1/Stne/Yi3ElSnFs7bK+p4Gm47tTiBjn1BorTxSPBqnQlWFaappN9AEpU4m6sqyaYau
WNjnFKM9rZa8JS8l6W4nmMNbEjSqIWxtBM76QasxNi0hxWLiAiSlficVkOTyvXu+HOgLoTOfcGpz
Z/Dq4QUxTKc6q8uZoz561ECTvdvNFT4ZqgOVNIDUnv6Yl86kvJvUhhyvxgfYbIeHdPsoWILjXMXv
CTDSoxvRXrUBgkdBCy7o9XO35NJ+a1DLcTTIak540J5KHb8/rC4482is7AJC6YU8h8i/8EXM9QB8
hb3dylVgdycgJ9KiVragvLcu7zxRWv1NgUStXcgJ8O/yrkzbOLJLJarRhGJ+0nHO2oeVWqPMZF8s
1eKle6Jp2oqMQ2Y/rC5Hc+AnLfRjIzWYp/TZnyDu0ZhpWk+aavymwkhg9oEUgWVHDqj+nGVzMB4X
zkEmGCNRDR9Is4zebx9d5QXHRAN4JGhIkPT6kBAooS8H4ZW9qQJpjgj72ld4K4sG6z6KQZvKZAAj
8ruxX08B7UhuNygrOqZYdizQ0GUasU3nv0x1L9iDEE9zFTXeiuFBPC0edIf77NqAdMTcB7SsX4jl
U7Xb48Ranb3j4XVcGymjxKSQQ4SPfWQapGD6WGF2EsGFPiONg1FTsbHbDtbAPjvyHVKj1DHD44bC
QcP/e1tg7p2OU0gWmyqR9xgq9jEHQUmwJCYg/lRrqgMmsmyDPOjac3G66t3bSLnA9PySRQkfex2p
kDgBUlxXV0TBnxHtMVGI1iErSAS0UFxGhazcouuV9qnsIM/79pGvm9q3VCQelI67k0vmTcOzlYfB
pMMFBLWqdrqqT/6UVWSN4YaEfY3YWMWTtHrLYiTtgWrBKhWQ90YFXvIW+I+G9KBv4Op52KfLLWAq
/xeiNMhFHS/c2HmRw/yCi75WQkBmTtv7OTxbobJZAvVYlcNvU3SnR6dTyc84X/avNusv3tATXHyc
tm49DwfE8gnxBAWDnBnkdcQ7/eFZtrrYqO5omr3mD+0gO8eYzaN/cuQqrNgEkuwqQOc2q6UXc/Ga
gI1kulRg+Pj5AFYG/wmPs0K/TLmRSTx4MOH2xC13jQjYmKyVWNFhBzU/FbTck5E1Li49KQQDi6Hs
FA+grznZf5eAlXoDZZAcUhpbP8BLdS4pvj1QTFOPRVmGhc41JgA9RYXAICsgb5UQDMZoFfDwvh2F
j3pZMgu89W/O7tfD9b6tPvNsjifcNz8wMnjxgZMxFtOzP8WikZkxYlq3sGuR2SnD3nfTZs2783Fr
wwDQQbZTSdCCjFn3gOF3VkeQQOxa2m8e0VQPwKP6xaVaY7hx96Wgo00KkIEATNxGH8GcNwQh1KpH
ZqRM8LDNTdw7QYn5IQEiJScCBoahzgOI115ShRj15uVIm1LsC+UI+3ar3EdkwtAahq3tH1OHyjo+
VLZGzwvTYmvOAAyodZ0/cisftg6XMjDqA2W1jDk8czvJuF9XLYnn7k+DZ6mMCMM5skUbUoAGKNLS
lu/ElwRUFlt0FsohHj1gZgwwrgBTibIuSUT4nqZgN33l4yxjmUvv9Tt1UUtXAzE/eQ7gpkNGjuwG
zV28u5MTOJl2CTq4I2hK6kxHD25MU2m2+16PBTTzQgvKEvlRWV1Hx2yssG2uDXyI9DqK2MrgvWty
w6LbUKIhHkw7HDPBj0NlL4hV9cIoydXpP4wCA5InmUgjtf3QmwNPNCRUn2tiFwJjVa7Cgr5mbu7/
nx2gcpJEKE1oRA08nYSxPTOQgP3UNeNV47i49sOj1imLMHwBBA+eF3qqCUnSdSdWcpjeu0aH4rHQ
//Setv2lT54DcltVzKBNbFENSh7s6HiUfRg9f6pVI4wzlPKjeB+s5oAyG6aP9bXg3V1nL++CMk2x
eg98VXoCsTI61fHWuklN2AkU8E+LpN5kYa3CNhj2m8tPYywAN52W4eWVNfGFz2OPqAH4cVlRnEei
gCPb/wfZJZec3NLOmXCf5tQtfsvRI51VuPI7PWRF6bW2ReDcyU9hX0IeloQS6MCUDe0jS+mAeeWY
ZKlbN7OaeFxR3dUVzrC6XNpWtDz1hkXkm+EMpBDcSyvzIqQIbvaSQajzrQzi5nMxMeu2Tnmpz7y2
wroQfMqVyi6OBBC5KzRXzTLvYf26wL8++chi1duJCm6NJP3/Mi9mgt0xS08pBpFbBz4rxYiZiwAr
v+idJCD5ZhAedYYmXfQbrcjoiEMn6Gdn9TcvFPZpIV1k/NoMwEdjXoPVSpu8o/DIJsbl8p/Fu5yU
dK/fuBYJjwLmCccJc58gAFIEMr6Ga0l5ibTBVGYco9ejlG4Fn1E8qt29c7Ji+G+qJZStARt4GzkS
RueNBwJrmNma+XqUt4cauh1dyxGGsINBeUdhjdn7rW2Nb5vEk/Uvp8SGEkAhEneFRat0880GFy3R
DdJAMVfszm7lG10jLSgL/bguu5VjP6naveFIE92zJyk5DA/iTid2/Ps5mD/ypj2W39IpbmAaK3J4
uLlH7ZiT7ydvmu/xBCKRTtjN+Lc+dJFZCC44Nq3aDuRJ1nnA+mDbcW4SZgV9DdIVMCWwcFEga/up
+Jsh9gu+S3kCxm0Bl2uIcoXyf4oweNthPbXeMzRX0XIG8F7OfM5ZYY1xE5otBJRvr8sVEfF8+VBm
6z82sZfy8xoboTDWiIhB0RJWRas/Pgx/dgpfpSupPSaPfaIknNVivo/8cwB9tE5O7dvvKFKAPwHc
RbmSq7sgA/NdJdwqffcddY+ES/+oWXp3TKUAAyxVm0X9TWPqi9h/+UUEdiDLs8pAnys42DCXFIW0
L+5dOBUaoS40gzPH+7HcHh4ZOGwV+RknbfAgbWSr3dutY+tMqJiWWuonCsMg9H9q1M010D05jF4i
UJrFG5Z9hbyYlN7cuq3W0BNqIbpCUsCuHZDf0DkmwZ6y5+HFrFXu2yg2svBS1W+kd2cH4xfdL0on
wAHtMTVhiOmScUsWq4uWoRSoEBFmil00EEuMZrJkUjHtlRPYaSk1BVhFU293jUqYiCmaZpRwETQc
By6zAkH79sA/1Ncusm/4pbpg9U0VhioLUzj5GdF1mpZAkx7RSvHVTa/rRUpQFLKUyUU5BOcoyZSy
S3WuJkjczWKJ8FbJ+8vGAE0te5glMx0m8F1NHNj4y78v5hLou+ArEzmX4S//TQg+Fbq7UHrMzh9X
lxFLBCf7uJBY/bwz0Ji4jdzceRwe4f46iWrUM0kF+b7Xnug2Db0pbQMwInaQ4ux3KOP7WUtulCLf
Hg2JF/KRUFNFpk6aY9qIPQolV5DVx10UApp/A1qgKAFgYE9uibor8u9PS+qst6MPGjpUB48z3Gzq
TBOSnnEzQ1x8igo9t0wMFVLm5ezH80A4RZN2GoGPIa8k7ueZIlkP1hVnk8NndAfTomCX3EluMKKZ
s5hNeKrex4VpEyEwjomg0yo9NK/2kbzl26RAkUjNcEIbCeUzDfsNq2bN6cOrFFekauH0XTTLRuI1
omqLKTVeR3HpTXX36D/D49/d+zP7YfMqahGJelOg0vwwRufP0kP8hPzbECFmUC7HzC7Q3sSuWzxL
R5dB14/66wZsg0qicS2VWxdMCCQnPpmyXy8qLXRTs+BhuK4t3ckxnifU4adov2YgVa3cqYtTyLZa
5yDnynVQuJPboAQNHMM9ak1vpLhR29TCM3+5718P0ovbytpbjbeHEtXEd+L9Dzjt3YaL46MmTWQ4
4YMrkKXvfDp0RWwfrgRugNxLpnlL1hB6JDwieLH+BdBVp69BbRMT6B1Cd7ZatKJ8ohyjZVLHrw0z
j5d0rxrIFX8QWrBkwXOlpSkplA/l7fWK/6fLvqptDGkzLEkFINJhSxcLEuHJBNs1Ulprv6tNhQ7F
r6GPX+/uB54iEYeM39wSzP0ZLAevGD1SV195ieZf7GNtTimORitjPC6Y6mXO+SI12yPpCjF1OCAn
+0QXV3IzFxjOTkInmimW5qRwH1kgbPZL1pgbE5oUxbs7Yf2HNo/brgekzt5HajSyPQTyFnaRvY5e
+5JOZSzTSs+ra5FIWDpu8qWWICzhtQph22NY041O3BHGu7vZ+a9C/ngKyZ6Hhsm9FJj0kMgvSMAz
kxetOskjhLOp4sprw2jKOXWxcnfzgJk6QcXquZARt85p5y7Q2rLqrVuJFoV+Qnoikidkp2e887S/
PHbaiRlvsFyoXV3dQIyxdYbRMtA/91CwVXZxA5BGeGUCle+sWI5020Mtkoay3mSmNq+D6r53bv0a
AeFJ4+yhCqx8P8MKFdSYYj/rWEohzAQQuWd14GgAwP+a99rIz8bfP2nfWkKMzXuopI6TMtgccQ2w
lcamZqHv8WZ7mMweUx0139CUwIG+ydE0ttOQFDnMGl1sa2C4/SJw7FXo2APoSq7miRXVZrEd2qSi
JeXQuE3MNJ9dY54D60OCEK9px47JdJybdT0Wa4K9UbK1DeqyiXTc3v/8N1AeMysnWzUv02zLt0Bv
gLfsKdE5eOX2daA7jK7JwQUDjnjKlkZVDnRCsdUXCK0Ofu0Jbo5i2T2nAXFI1jCjnQ+6DloRDya0
WgrdZ3Om3ztAtCfsVT0lyHDOUxASaietJqLsAH+59sZdkIXQDLXd2epdZfHm/uo4xbuIh7YMI9MF
6VoT6FUS6eJb9jY4unYNu1mWqXj53iNu5X5u498GHq2euqs1dnrxLzNNy9MW3F0YiufjSmSyPTnn
3SWYJlNdbqmtulHmq3dXGNrA16B5ynJQVSPnwPxNCd9YjB2JH3ZBHLY2Q0rwGxUqsfUttrTeyfrh
hQ6DljY1IHCvvxYtNh5GP+aS7/NUNG56oG/9hcO6BtfkiCGs1cXxi2RrRrHp6dWqE9YzFM8e0VpQ
0+EDkHuznqlB7pGVtAa1WHkOV++ibmd0gUsKAm+fvQvSOkdPBbyI4wSbQWKGJJE2nN+1bGB/xCkY
ZQCut/oD7KkBM1jbb9EYJS3dW2ytg7qEWfhLe1lTLxpxDopaBC0soGEatvL0oOvp9CGY99fY4ZLx
CmYclSSWbBRG+LSmbWXTGa967oU8Ud5QXQhkB2crUMhT8mjDZsnfpdOf8pWapMHl6QmOQrseuXbW
DeCgpvy5Sv9BTt/WOBCeQeon3J37e+oSh8hRxTLYrj7/GPHe5qWdVSCFkne/wNoEx1zzHn3a2U+u
H3fS+pGlEEL2KzzZ8fYOMF6fdSI6elXoKM5dicNVFAeU922Rmd8b9g1ehb16iQ1w5Jc9+VkMHilI
UVWibitPaJsdJ5Zaig9Ce4Y/z7B+9aFXztbyLM9QM1ExT+VafCKd+jHlUyPV43b7CSSBtUpgVU/e
i+q2VQAsduv4+PWoLYrwQhNE5rpEg6t9hUM26Drjbfawlf98HPGgcU5XG2YLGy2zuEz+fq+0RBT2
qSDt5Y+Umx8+tHFUONHHoloVspc1LrfIW3Ue55BdZ/vr6PSSUtCisIHKmSIR2p3tlN0RgQpGpXbu
WCCwq5vPwzJkaCiPttBRctnqPQ9ymkcxrdshKZfnjwJLOxDl+Sap9ClCSXyNNbEpYY6fRe/d5L5t
WWwlB5dxht+uFLdL5zJ5H15Yyb8K3HQxAqgr8uFNTi/wHKDLJuSe6wxk5wLZZs755UXCNWhEHaTq
yoz+haa2R0nVXx/zH9JWEwx3BWoBAwsraFeat7j0NKThvVC7VxlMe/SSzecG82Nln04v+IzeVta9
Q4FUk90Li9V45G0S9t+LDt42/0fax+pK36ZkHXKjabPnVTdELEPKLz84V1D9O8ap1XU0WQ39K//p
MS+Xi2plL4G7oT0PjQtloSl+MsTPhmD2BeSdbS8Oxo4Jhquh5gfHb7BJ2J/iLbQ/ulUhTJFQkZpc
jwrbweeZ2tnflTsCEy3WVFCXyHTAVJKeyMs0rf5m3UG9yZkDfjg5am82BsqFMX1BYSh4WWOviDgZ
uY8vqI/+8KuMjKqXj+UuelXjYuK6ZeN7E7Nz5pDxI0zLzMxtUSA0O8fLfNQyXyfQeRflpoPCRtQL
ExRJgE0tB8Lzw8U27oMa9b/ADjRqXl9iK4Ak6qmPXGlJUOlgWHUbPsJlW+dsZ53TtjDD++v516gD
7CPkD6s4PeI8LdIwWJdNMs81PH6L7nfZKs2YtSmaeMR9I02aqTEPgUsN1jaN1eDIJ2hk+3dMQF78
+5c+R4Xiea2CMugn6JJV7MWao4oQB8u5Jsaw7rNHUKfbcEXUMBgBQ1e6D9rzaCUZAG24MzQK1dmh
VxVBJdYYB0jh+yu6X20Z+bNNSjU0zH5V7SAMJOfaU524wSHSLLXpuy4OYwVdjz8PtMf6/GIRx4Tn
EmOLGEzNyGYeRTZdd1WJoKXgzNW0656luGe18Vus8vWYVka3YzWKaXtcPmqVH3NUsNQsL8TCL+vo
LjqLlbXuAHam54dHVnMasflBwmJR4K+J8NCB0O50eUeTGtclrhZgB/XORqSzZFcmyUwDiN5slcI3
0BJNzYgnI+N7mPvKG+FaZiEfg4yh/lvhBY04LCOTO5dKicViRYNP0kSPmW5Ru59OQQJy27xCQmVU
AlO0G9ANKCV+6oGcl7UFp8YNuv2mWiSroO7TeWRdzWJC/VYThH5rQvUI4fPYNd4MttNSrccaFevL
/+XMC4u5e2yl9+RUlwf78Fe3ShHkmmmLHYbxf6gDas/c4mKvxN26j5oxbk4v9wvq2xlu2eKPJgqD
PaCGe3XCucBcNPRG5N/pvBLfUm9HtTzocNvMMET3iNTEOep3AonFCYP4rWHZL5GgizvYFZD32+VS
hkRjF1vIiCy9dGUmZUM0fTgN4tThJvdyziKM0Tos/sds2Rh7HviWUcbFoubCQNNCxeZYFCWOzQzp
bLUEA4p4+4zAIbn5oi7mgrPyxtCXpw16lR8a1NE5x0oMS44tivRyTbR7Jdrp2RH9l6PefpPzf9Tn
hZw97lkRMKFYWHH12cSGZ654POtIPdH/OT3qFs03aNNbdjzkpRlVcWRK7tyh9K0+XTwYl+Kf60hm
WQnwY4iHVGHA6Y11VsrfkBblPFCr82K4A1XKTzqd7rNDgnKKBdYAwqlIj1GBslovNW1/iDpBFJzB
A7KED69iYZqnb6CLvyLYLl5FYZwmqvTjLxDmMoSCpasWh+6P8cMK4gyuyzTpUXxY+GHLEvlVuah2
WkghLbo3YRp7iv735YnDZSgYsJMkh1LP7TJNDjh4b7/2gxABs76LrElOsbzg8vgIidKDC+a16qfn
VOTCLJAzQx4DneVPno5LDsEFOSA0wLetO7LWUEFdmkFMeyeahTvHWJNigq+VpUjz/Bz65iX6BLVY
HAserCyOfj4lTFtZia1JVQmQ3igtTV1IRu2TPD2nfCpspaC23GhOeYGSmovIPwtpGdK1jj08SRRd
HVkWTNN1vDaNXfgaco63L5Y9dxzMhd+CJjLSc7A2mhL92hB1XeXMl3Dds2P/AVnhHvitwQAp7N1i
YolX39ll5VTO6zuj+UUbURSa7najK8ZhSffKzyoIHNFhY+xi2V2VTDosr64cVybUmQzlmkDkDt6X
RMhX32Q9NrAn1C7XAM6UrMNUkxtb2+wmVny1+OmLzgbkk1UGybh47HYdaOjiXMShv+Pdf106qlo6
rcZPZtZRWGnTGZaKYV8U/eFgPGC3a41tLBZ1DVP4NNb3eTl02hqde1ss2o5GRZqOO5w97crU7Z7k
MrLUnecCPPFsmyiH3A5YDgPqONPJLtqc4mYojQPg6qnWe0QnX2mTl1cHvwLBBrCeYbZfjq6pgaoO
LaNL+jBnSE/mY5hcphYuUJfAGcEQ9igBI8rSZDzOx6dzkfQZH8+UdLKRjZSvEFiMBioKizSIW6R/
ZEYMaJrh1ZFTDTcUueA7Qkox4K5ClRyCQQz4bASrJgk1voZY4x8ajWz7xz9y+SyAeDRvB8HcPMUT
9gRTe80ecXH7JOzi6nFKuVdAT8YRzp4FORqeDQUAFDIgxjRTSkhFkUY312hxteuaDUq0+mrwrW/i
QbBnTVRVkAsW8XV4gQOFy5Bq2kHarSS9UUEgyn5d5TgsckjIjHi9KVuQKipo70pdxwt2ii5haZcM
u8FmBny4dGxwWJO13N5Gg04RqQn3ZxhVREHTqP02EXEPgD3VJGdEO5cDluNlOXSW6EM4Z+6Mn8eY
XdyotxmcVpjwa25xd9i0Y6P/PN08hjK1DpfNPS2Ie0lOdKm9hq+CqHvwdPomSeTcZAAFoeLrHEcR
vxXIVJiJCRtPpWvyE3oJ+QiqBrUcXAF6ggRM/FA/XjODOIL5iLfJMvoCooWqBrAJs6Zbz3406w09
4axkj6gXlyV+SVdUF0YEE1mKER9WOz9CX5jsk7a/iaj2lkCEqZci6ZeaYVmXp03QwLjLxcWM0rWY
bV6CDLbPzgmCblPIKqzYWamsV92XTpOwWMryRsSGN/nAdox/jORUj2IPomWhxXtDc5Pj/OvdnQYh
1SheVYD/4eQ7bLVwh+D701/h6jT0cyIBrDbZWRNq8U29pcLPzcuEZj5FRr1/tLlDJyrL6bXO7ci5
FMajz3VK1kAu5iBR5HEfCMY1PAez12lGl6tFjw8cQPsA0CD0STdom+5TmAB0NY8PBwKkzD1mouwR
3+XiMSRTLNOdAKzC7Sxga+h63jVFueSvZurarWmsPr7tGcIzLmtd1oKW+4QW7iHqSZo5Siiounnc
u+CEsSufGXqa+J06URSmZez3W1yPFRVuP8hmspMft5iaRShIigrIJZPr10vHMFigW0+KFrxLNFzc
0J7kQzwStCxS/OQGlZt+YZHgNavYbx0iT16770BgVj8f/Ak+NCipIGSgcfRS31wN6eXGRCaHCy5J
/IFtzDKM64FZkXke/7y6pjvOCNwUgpAYVBCycwqBnnq0fnfrwFXN7UswcWJ6/lSxnPykx+ZCx/s2
C9p39miPbjNYSKlPC53dR2dnW9ZQr3E9pWIggRtBTtvARQURg+GWACxKFWNexbmBZ5ouO1xuEb1R
3FBaxD4ylqHZ8mtOl+GQSJRgGXr34gPBs8z8hMX5pKftjymdB60BrYXW6jBbvDhtE4AukRrdiVU8
Fi5L6jL4E8uZ3VORh4TrzPMoFJ2j+ANRok/buasdEFZZY5iHAwkB/FwYWVTsVJRRcGvKUCPRpX+n
JSGEN/kcVg+0Dj/gxEqUYELPPQ5ZlZwT2vUxYjiAlcDEH5TqrUkjvhiBjOvvtzuHOjAwPwIPUzS3
lrIgvRDjViOhJEZdwDokD8OAC4C6GLeqpAYd4ll0c0vVg209AT+kacaJPs0VRZ8va6wGn5cLyZ9l
xdMxEIXjNKK9eOpZqyjRftUUYpi+hvsrNFMdVq7yV8Ewb7Pu/ORMli6LlJnXP1JwAeY4QFiJQGHw
rYEONRCFSMP/6RDN2hinUAiAXh4h87QUwzJZQdY1mvG3eseHky7p1jSqYyTRynGWhv+jNcVmp655
DrgCrLtV51C2yOBpscteyQPakcZfyro8cEH9MeYHcVfAs5JOkKDfY1Joxb6GjmhJK/9CdEXkMchb
WWKtyIGQf5jD5GCdR2V7Kl6/6UX/oMOtxReyl1Jch4ia89a0ybJSD+KYS+v5TBPNOwMKb+Lf4/UO
WBNvUKsNo4nXN6MJeElc8axZINnq92rFvVpUECNgLiR2QZrk6SclTbuZaZF+lk8IP6ExLq7Jfc4B
tH7KREErePQnfInwkU8wpyMc23MuMHK6whsS8rUS/2v46QitXAhFoFMLDVj51Iuo1GF4g/Moe/T2
y3WzRdpnt9J3Zxe0S9zsP3hi/ObAOEEiAd0ZtwnzC5iyMY/pHFAdUlzfT2YRtKxN/co3eiCWcrPo
/LBjEY9CG3YbnstQ5VORqzJjrkrrnWSTl6ITyE6ZuUyuEAkAwNg85zqBe6mdufgyRiXaR9HPutT8
wFrMdIjoGdpoNGfOE4FXXVbeLbCqICLuR5NtGmt9ejGsO7RZVH3y0XOei8CFoL4PPtr/Wur0nbrJ
bWDiu6tjL3ZG0zfELbj6urg7sl/prKv5SAPsrteDoHd+B97gqbQtceeB11+4OAZKci8rzUeufcUO
fwYdZdPghPvTmH8QbCYu4EDpxekAZi25T7TfHAkl/4PdKhfVBSfc6m89PhqBO7SLmGLoYaO2e2Dp
83gm4GpPT+9asHw9OFoGTtR1mzS/PHNq9BHvtcgjQeROBIX2JL922MiuyW/1XCbIXpGcR2dsEQyX
Fxenr2b20nrIrodI1A3PIyWizKds8zYjLvusviLTawy8V1yi7yZzvgKE+5B/vRS/GOxuu6kX7Bx3
FkKyhU0YTuwS/zr+7cDtA/NNn2GVBDgE/gsADROy7CnMG2ipl7zG+f0D2i+un550xi48RD55aM4F
a/hXqGYPn3MYkZzCW+S1D4yUM2mxn7wmQsF5tZmuWPpDLrJxL6eQGoBXPEupT2HoOqgg4YgJ5UZn
ClA1hvZQuNtiXXWpQmFkDcK5CuCAsVQfDHBb84bEDlvHxnd3DatbG3SMJbGahTVjbxVEpcpm3xFW
Jc9HP9UZZmp/JovULIOShGv9mkS75VYgXK363s0FGoADGeXakXxEF6vyipIash/s9voREc6ABurM
wh9sFtBwro0Q7UjI04cGgaXq7dkqgonXsCkz6OoP1pspPTCav+iB9gPtW3HMQID0g5widLdaH4Rl
780WlkmQzCTHN1EqaU0yZDbp1WCIp4raKS3RPkB32SE7vn4J+HxSJMpi6kH9gRM6mW41Lg8aCT4p
Oa6zkSxSnL4Ft2IP5LZD2hJin0rbtH5U45Cbgt2Y+sn9AbfhKmBXEBud/z+0lenHgUhyN+WNogMT
MglhKUuQSkWalIV3LDxATG1MXU0HxcJWck3UE3JweCfgr12HwiqN6NpTpA3EYEQi8UH1TbAGCP9C
IpCbHBtC/tqxBff2lE7p0rb7rHm9n0MHGK+v3BE/ZXBgMiLzTMnJyGQKoglNg3X/PDw9hzNA1BWU
uaY8OAouyENkpJ1jkMjy049scbseEp5SNQ9aqwfPYLpOeQTiIOoiQ2CaYYU4KBbjU+9pOB4X57BG
Oxgo7NWKj0BjMbHsJ8vkoTcv4MOciLBS5KnVn0h6ejlgytJEzFDX2Vk3+9jAGxxiHBo/2rgwLGV2
YDZH8NI94z79MjgCjH+p0H7TU1YkhycVmPcSwEHio6iqqGghqUtoW0h2j8APmWglO+jLIno/jxIW
4XQl5/NG/5BPCYOaLgLyYAWaI4TVXB7ZczHVazocEwqc8cv7b5nwLwvzsMgGnXCLz8rrQySX6taY
w9jGndM+ck2gIo6At/WJqaNjcv0t6dg3qTt9vAD2YGqB6KfLdwe96YtiklmIKF15PuUCrGRqvvw+
o53FqOR+43mcDDrOjEmoVdbppBT8btwIZLY4T+K8XwuIC6S6goQh3g4+xBmWqMckoGlNedQuwt9x
F1TEDCNErqT+ChDI4eDxtPw+hqh0VIS8YXnBB95ZCCSZpQttHHeqsD1H4qGLmL6WXbm/QNh8gIpt
4nmfnWDSIJVeE0vg3X6dEcB2fM6ZlurwDSHHDAudUX2Ow7q9FUO5IfhpuBaXiuw5ofM7a/+dUzIO
0OzsX+8mmjN1BbKjbnsfSde+qukHAYlhi2f443HxeMmnz/eSZktZhpidPqm3fiqtACGvCv1oj8dD
1YH4RTZJ2nb3ikZlQrBSL2SfTOPqfVV/YYkNDoTcwymZ5qbKOKF2AM4q22WS713hPdnYxTxWCnxP
Cc/PcnyOfvSWQK1c3HoRTmHxBSTS1HCcL+asoCJMcBKSparXzHi61Yt/mgQN/+9A0xIpEgXr3Q0g
eCWdGFM5ww1pAZ+i7wNyPko1aCO84lbncTTOk5S/OZr3QgN5r70pJrR+kuU4SS6yZnPOTqkXMk9R
R0kAIqXwLqqHGIeO+bth7GnyC32MiY5bQrxqojc6PtFYQ95bCXa+nBUMaQG2XjJPKa61WUFXAThB
LNIJ8OqgCJb2re9cWXsdwtFBTrMkximQVWmlufqbmKaBbPXI0m+TRhuNna/Ghrw1IQdBy463aC+6
/xw1Xa6tO2XNTH5zutSjdmBNrYwttSuJzqSNAIQHv35RtPyWAEa7H56LWvsCy6NHhXfW4EiAZ7A6
cjZxMzt2TK/20wPFaIMWX8GQkwKBIiaJBoIaQuyR7w/KeLyyeC9V+8nRMd7zNxAnQZdENhX0cnnZ
3XWaT2pxqTsFFzTlukatrR8dhJpt8IP2+CnFs7FjXLtQ3ogSyjBgThsncrU4ysNlbVpQ++DDBqIV
naCCXAUWJctrSfEBc7BME804optLpA8EDTT5QRkPl5YX6jEIgW9ZPlwnihhBjoCY3XOkf5YN+iy5
Qbxy0RVv2ZSZ1bXJ9CrrgFSLRqGH14+uGmsDZOoSTGT8Bs1zYV8BNG4RhiL1I0l0b9Xu1/P2r3vk
p5+Y7j2saxXwiksgb30+gR0Aw6WsxEWfR2wQlmmNT/u/FiTGtQjzqSFFuIcnQ0wZPad/lCy9E0xo
Zuur0wUzjsehA9WWdjkDxWTxY5i2SEcNXYuFdoaN3S4zktFmKy76oA4Yuy7xyB2gFgfSQ/dL9KT1
qjUnBDxqwLhhlskxRcjvWIsTwLE+rUDvs3hzeekY7eJDd3y/wttWasKm3oy2jrQ4CInnet+ZN0GA
bYqa9mt0s/zXmhu6OMQnjHNCmxnkfbNoqPdvKrRQCAs7dJOM1kDFBQi1BFz5nXOvS8zjua0CPLJ6
ZOEScNH09olimwXzyw/NtoZCK3DOc31f5xwyzD6EBrCYuQG9Q0XeIpQII7eienLH7Cvlj4C7lm63
CVlcBHTiLMmbcUM0sf40ZdwT1CPbTnsvqY/tpgxkPT/Bioe2sFnt9EK1rPSFhpd7mWPfwDR/5+r+
2V0XHq0xB01EMM2sLYpwixTXhu4+uRtj+LWI64XLezpbeMxhekFdU7Sl78oQSGRjojKVnT0Vto3o
LXLzb6CHkx4SuuJkY1AoF5he0qppEksbxWY7hjcO7E7DISMXrkPGgNqg0pxY3D9wq4eP6fJuzh2K
qNeht/7kZS0l9tkthQpqGBATRjXNLKAY09wOZcvJ/33/xl4batJOB66LTzwEEelCazep7thW93yg
HskOgU595TCLGDUIQGLLBhjZmOX9cqoftR4q3RMeVXNJ42Wbc9VWYK5oyz+7k5Jlg7jomyemGMFW
TS1k2jLRw7VXlX/O4X3jXa6KtmiX/5KgZ6XIot0RwdZ62Nhy1cYA4E9a3jcRJz4dKsOD2jCOC/vK
2OgFUxCpEC6jR6hwO5YPNxdA8VNTa7Rlyyzrx50h717+Czu1+d5xLMFWn7mYP7c0/ChF/cQEZnFg
Hdabd1XRWhpzvQfnjDgTGkDf/eizF/DoecZq7qUxNs5C/xH4vn4z4XUhEXGyOoS8/krZSeThtJXb
imvhUJreKbWIPzB0e/bulW6SYzWAHTHSt0WVt1MdSyTLs3vrbB8p2+Y5Xwn06mVucvQmAMncvQQO
qY73ngKn0VroMmgWuC0VPgwWfwxpD9+KnPCgpd/2cvTX1R7G5Vw3Ldf48hB8tx21gOpHGtTqSnSO
C0BZZJxY5FYRXJ24ezGkWFMjN7bzL9dxRzC0qIdCpp+qZXBaGGoooHXZAMSYoK2s5e2JLb3pCrpT
OaV5XBgX/9P5JswiLtuU5a/MSK805424dvHh6N3sVcNYKsgkEHoJyVY1rV7WxBSqhz+6/+QzzQUG
kPjIB2ubUrp5SbqtLl7cP4tzV9rpn91EGVw3eAgt8L61QdYGnxIfO3Qfny/iTTQc1dBgrt4lFSPE
uSv0uNmtQmmHBJxZYBu6BY60ppM+5bZwUOWwwkVX7LJoWgPE9ZqaW4x1FBA5+ooq5js4rIB0tgR0
H167IPN3bX1L4pFWeok6xkqPi2lBCqrZI7g7Pwp0hs8Fx5J2FV+R9QH0o+GavH7sZbfNs99q14Z4
2rUqhichcMlNTGx6iMvi6MZS2jMSHWLMVKZxqFfzEGdihlPYGJAZoIycEqu9FqMUXUbxa5zfkXMP
X86O77D8hkt33rzefrX32wGM1fYfAVVThpBD/BILddsbkwELrA2qIHJn8qD3nObny0MYrs9/EtMF
fsF2yRXZJEyPi0LRl2KGKSNv/63PA2OKnpD62Gcuuuxq5Ev2xU3nuMM0YtEDk43WIZuYWw/qAlQ7
XpcTvv7KnhJ55jyMs1VimVLAF0pObtRasOCkwh7ynNGXN86LA0zQx5urgAOCJnvPduObi1d1wUgF
RvpXfkaJlMHfOXqqMnwYom9dHMLcjwjIWf3B/u10yZhAeEDVc24Bl/kX/1T99UFp3Uwihw20he3N
aNSYJvQug4SRR31Ohg3Pu32lwYs3Ydrw3tvosMskgPZZIZHXBW9MlQg/ybWRLpLTZFkId1PvcEyg
Q0MhFX3DemMVSc67fmokrJktKPuGmxdWZ3nwygagzhzJZNJTWwsOtsQcYTibvP5NHwM5Hz7tFYs+
/ugHdMJFU5ztFzhr5mPm4R4YgqgZ0YCGMZzvftb0H8jg2JXcwMMwij/bNUTxR3VXyMoF/wGhn0AP
GuF4J89dZrijTbonEze1EuKQdnkgQSgPvmJZdV5SqJHWlVVcLwQS59unmUz80ZgiypTPBsqHyjwp
mGdS0p4ttDATDvgFMphB0I/MkiJcmnp2Cd5DXtu3BS20PsMIDrblXHBEmXu/XnMHrtOKlPzF601m
N3w84pMnnHkIzQZwzoni9LV6uqX2ElKFDcqMwbfGz07uXLM7Zo0YiOdCAEKejwFuVFF/IUg5+R8A
U9fcdTyTDp6HLQwhM21Nyr44+IuG10cgUS1YLNzG47zbKEYte8NRiSszMvik1TTy84cuvAMzWwpe
klbK+WsuovD7ZcDqM1s9CiRl73jTEUQraUkPCLLb/D7FZraMCkl2iXAx9MlYG5WBDwNjrcUlfN5U
UoFpnbeFHE2yM73MMBUYCObnP6BdNBtL5Vc771+59JneU7Z0lNBEJUbe4WHUSNIXTWObSehCv643
Qq5OLEhtkG9Qrg2F5COqRwGSErTbX6/6hrWeA3drDHzAUPkvzM9LWD3LKMlWQAGsrW0WoV/zJnfR
rQCgSo82sMp4MirZFX9/jTmp35L87RGPpNhoN0ddXadiHZlcenoWbUhsiXeIfVgUzP+QQhiFMIZh
FllvXDh2pBQBRS2RwMuX7I6JDhaauN+y8gmqOsvAN+nFUeMzyGYPTmr2zpYJfRlpq9puTGkc13gO
rdQJZ1KybJi0bdGe55xmoH1BVYYrR+nizpi/JCXILOynbaZsdBCIByRzdKuWXR2hK+p7+2jB1YT9
BGtmTIUsuZsn6KBLPPO3E20dUB2IiDYn9msarv4cobQWh8+EvSB1DhKy8FR16r2WCZz0To9DspD0
jDgFtWGNy9n1SwDhZUPn6i+Dpcc0TbYiD4toE9pB9GKkMaLt/7AJ7FkS3nOnysbcHN2Gd7WsPoaa
jTcRXYDfzzVkWH5+C+SBxklu4IEY4FTEDDyogxxEhz0cLUvrgq2AoKDhXGy9oFRX/al/JmTQaobh
AIoGnC9fvme950r1z26eUUlkBmMgdEvYWDxNZDbxhByb0PPxkUtgdQv4NyPJink5wlWelhA2N9Pn
RT5aefowE6+HqIPntXLcE0aVcVaC1/wJ5wgjptfw5vhq5VtlpT53/LCUH3TEp0Rv/F63R1OQxtfb
Ehi0t35yR9XuXWPGOAaOe5uIbF4gUgr5DyVCs4ecNaHs3lMq00KBJzv+UuWsSwGBB1f5GrTgbZ+J
7FXYWLQbj4+8y65twk1Uc+g/D0YAco+BMWqTNUW5YVQipAdRSOZzGcqgKvUS1TbftUuH18L1o3xa
etTlTCwdYUmUo7CP2j6wQSOllZDxKdTuKgtdc7PkvR5p5QmYf+D/Oaek60U+9LmdQpi5gQOhmSm5
s4vAyPoR4uFXbtuIyArNaM9lSS2wQD5l3pElIRtrqn/7RjiLYj5TSgJ6Kdc/QST+bLYT8lPWomLs
swcdHwTdF32Q4ST0MxjBRAcjyODbEEKvuGaaRPXroOgXER5GVBhdXytqsh9VywKrHk2VC4xQun3X
nCOWOvp8Dkz2WLz+xzHlKV4H/vd7YD9wjgflD8xrLhte4uImU4uFyRSvefNPEttzMNKPe8R5TX8N
7kwAmWfW+TqD98YIopdwmBhV1YiPzzNJ4r4p5pqglMYFuDw75wI+S8E2Ij6hpV2sAX2Ex7qdRz7o
2h1jNs08afBN1x9DMaffVg9YH4nCFO8rYAtSULFKtwMebJJ9YeJhCByj7qWNMafCO/LDh8r+hAQT
a5Yoq78Yy5DdAqd5Ka5iumTnvLze4Jpm/CUYj0OE6/g2Fyzn2rEUHqAP4df7LuQ/fgT1YV1ISFOD
JyMKseM/tjVAWBfL2oJEh7xqO5GAU/iUC7J9/p1PRWWp36oJjYT9F7onyc/KmHCGng1hf5+UDxHw
DVMPHGl4SRD+AYN76lR7uaAA9cb8HR55lFXjDa6yRqQGLFvX3tySeL2Ss4265CaSii4GIJhwjqMT
YEo0bzTQe9LYJntJ2JKVDetNI8B1qbPtu91Xyc55uKwH66tYmTbRo2h32yq97RtxvWguoBrG+eR3
enczJiJQDzXFekewe2TQJ3htWdXuNC/PbLBIdpU+KYQrLA8Mha2PviP7x362T3DiMTHxPpa3imqL
HFsNkDG/y+oclFkPfD6AckGGltShHTjkRmQAZW/8po5LF5dECk3TJJDFTPnJNgzfPem0U+autLAC
wiSfWc0pXjZwebUknyMj11OR8SjSWV9X0SiiNnifoqA9cZxv4RjZaSgscxYd9uol3BhGFwrIcfC5
WVlmy9wLreiUaLE0mUhkEo63vFyLYU+RPVxDMwYP2FN28vAeWr3rIhhNca3Cgeu1THfTk8DHmbH3
9D4x9S5jRNiTnu377JH64NcpYLO04bSk9MlFV21oTiGaLCv2MRhALaC4XgngmA1YdUQmelyYDBRM
0Z/nEoa1N7DfJdSjuEO3+h1PIUyD66Nb4XRq0L7vYZBj5FyR7FacVA806900wEYEk0UyYCDXaIrA
FHfadKFcnuHC+orcJvhJlTRrZ8MvaYDSzJ+//U2uGRa9FTiv2Vnu3UiPaPS4jnGaQF/ROwsfbs+7
Q7qkwRuJeKbFVn4g8LCk22oD9snYzGw1S4iNPWXSM5ZJnVKiEH5rjjXCt6HvggJsJqdXlO2T2YdO
9Jk8F5j3EYMA3OC8XG0kn1wpbI6+BZcxhIQH9JnZZsiI3XvkKxHBVoRNdU/aW5u2l5Tgaz1iVp2e
IKBt5FwxnqJDMSKjzheZdp2lIt6IWp/NtpMmlwvCmLz8XiHMLo6QUl5ucnVIUuFUecxzzdKemRfA
2I7e3NdXBPs8fRHB2Hjy5JrA/tmM0pTKHMrDxcjhMd6ZdFWfK/btaEfpZ4dv3Hryrp0LvdylyOEu
DV/8DseAk8UjjDnmViSqxJGfN62hY0zZn38zVovFyW2z/Ir6TCfWx2Qx9Sx0+61/Mgnm7Hg0pSy9
3IasK+dYmDuARJS+n+tOFkJOvHKrWbJUrENfJ/QyAOKdvb6KV55Ah+YCppjzXvIcxDdRODWtOuXk
mSqFlpYmLSONTGQnAs9ZBj4CbvR2LEEFp0ljoa9BvPW8YU8Vo4EP3CObtnRHHW+2DAmSIxYcPNh1
4mi/rCemjCDK5Kxq7BvPQa7tYFT4rEbmTfSpbGndfDvnKG2sMasainn+I8n9BEpa3pniet2tbyO3
0Lkx6mCDeLUiCJXTNl26wsTxq5EabdsSn3aMho5VsgNVsNM6stTm8naB4PJLuKPyxipnMAZZJRLh
XqIAEya60/teMZVTP3zrtFx6pZllNazHep0cJPvIbAHqitgO9NQr3Nd78xeSQaxF5SsYREwKiU4o
8Pi3ETAtag7DKyzi5f5UJivN8g+3QNFApKaODubp0936yaiCinVNdnO3XEj7PQXUxGMOfDEhcrj6
ND947e6/zqDzKz+LkeQ3fWqQRyhuuo6WQlFtUu27TjjQcUGA8aPk4QKk+yNfmYjXo/GIFWy4hMs5
xFMiaW++yMLULt7NICxymeoNuL5NLRf2CWbR5hYmFfmCGXdekzGRdiuqrxZ2HVSVvwbgmLeBIMHP
+c8fJr0GAeLFRflU+BCSA717uGXYswgPA+ncPLemnLrIBus8UVMqubcqGxNOCeixMv9RRrOJvWrf
1qy9RH/LoS6Hfp7M61y3GZ4hOvp2ydJw17haYibLhycwk3Jx1efZoika2cgSnYEgHldzqtihAKQn
Vvq0SQII5d7mVnK0VpVPsg2VHdelTAPbf9Ee/kNlOqVcplGAULg5OXSmx5DRV39i55qO4CT2bELS
wJy/uLf4XhrebesL78Y3ApAdiRh1VEk/47BQbDDQkjJGoGyh4ehXNDOT8pA7V8AR0NuzcqwnQart
I9jFdoPjJYWY1BeQifue0PTlV6gQKRI9lMuy7MUsybaiD+wwp0OclvTtTFG4QDQdJv+QV8zhigmx
rGf2ZrHP6fW7dAh6P2DL8600cVGdeqfVhpNqctQcKZRUCn+HyuJERZlG20U1JdkJMKapXekVZJwX
3qMrkEStA26VciwN9EdO7xt05QXi8TjeeLTcgoGY4+9TTxDPt/lN0Drxc6oh0aJRA+AIgxOC78iV
rFQ9x/SDYdhnDl6CUawOmJZJ3Q9mTO+pjcJrjqcDeF+QqHDkWh8eDPpjTm1hvGtksDZAB/M2j5EW
W4YN8Ddath94yGpf6lZU+2p35x07Mb/OEbFBHqfAF0vfNQb7XJr9MJYcVbW8384MiwXUdl6iunDT
hZR9vgngnWN9Q8U05tbRhGoSySib/cu6TZnpI2qdLpRio3jUyohGXnPwgMBJzZBEGVcvedvaDNxF
Yd8bsHqBIVSbXtzaF9C1PQ/gEB0vDE5GsLk57u8yDAamCCcphal7FX29CZ91fmCKtGJFQVupNyQv
0TPkoihXQD5hk4KqdAZYxWF/I1nr6BZwwg+aAwzPDHkZ4I8g8sSerDjfnv3WTVd44TKXVfnfVpSP
kheQ9F+TGDgtP3gMALKiZw4qjzPshYjY2dBwPowHM9xyRZkh2pi3F3MTyn65pLA760+MKnojJ6z6
YpRd20fXARe4FyW0aUpIb6jaJCpW8ozi8eRCe+8eJ6t1FOFvWV453LniQZdZaWPaQ0MIZWDI6G+y
hToaS6f5/MGatprF6WFnIXrbBPWZTXJbRIph0slLph/XRxvcyJfRPOeWNsXmHjBHf/RiqXMX5081
eJT4opLOgbOtVK2hd96SvHmUGFX8wJchHdNoU+5moPQwxahSMQtCRTHsYolsL6s90cBzryEJLOiO
CsQWMnIj/y+8ajanAGi/usRjiag2Vp2fvPXzgEHubs1cNw1a/LTNGlFHxeWVa2N2uoznDPIJHAkg
Xtv6OudHzH+OY7tRFKQeTi+jBCY9qxfysyKhZqSao1uG4WU4rgXOKfubA4hny50qzKSTOfU1sMjy
eGmAGdLhQG1Bz+LqYzW1uy6VgtPtdZSLlX0uKLQcLo/YqgdBRyOXdOC8aUtYQHDibCWGK5u32/RA
10ptOMyGxqm5p6ewq47cM/AOotABoWi8uv/3RAwfqZ3sK/3ncMDMvwUhuZcrLJpDv2yY2Qtg9Iz7
0NVHj5e8wdPjHhmG72dxPdFYc7LH9XbeHi0MM54W/TDCpWzFx9a1kcPUv9JM2J+YBYsz0cR6m+Sm
EUeHH5zifBv6XH8pXoJyxFiWp4M1tCWQ3CXK3ln8RSZ7GT4wq99r+LV5jLsHiBma/snB2WNHvo2K
/mHBv9+USBQRloFoceMS4PhEhtTzBTF/Ufp0bTbfuq7QjcbuQUIQPccM6ITK46TPz+iSfHtrHI1q
u/LQ2kFHrqT5WwDZSZrHf1vCXfI7de8aKjdhKgcETmz9fX0c4ua6UjNXZcYMeXgXbF3S+Iro7oMd
JYHzqUcRrb5ta8NL2wpEReHcUDrne48HfCBlMLBWzwZKiZGzN//VD7612jjvIfRh6tuwdL7dmcE4
qebcCGynZIMcrk3w0MlYwheLB67tRNFMI4iW2PYe3kn7eKzFBgj0WeSSgfu9/m8f6oHbiQivedpa
lfkrsb5o5THPzXVyHL0JBcknpiHrNQ+4FdDbd9QYC8ln4sujpMDL/cFNqvQ0lSswHKN7www4BvPY
uVLASLtLr5X9UnKNH81i7mLyotXKckadwqKzmqEL1l3hjdcra9FIAeRjnqd4tfo7SaMIH3y12GAw
DIpz9CSy97SP/6PenORv16FN3qgo5/87Iiqj6Hncqho+Brc2jPAE9dHY3of1Ga9+s6bTDcQNEOWx
9EL0cnMTGh+Wx33k0/fo+FzQr6zUKNy8AOGcPwLvHBnm9l1g9GrBWeIDiDDJIizbq9iRyX2ht9Du
xUeG5YBeZQOBx2DJW5BXedl1GUw8QMT2/fkUrd6UX+u7sKDsg5B99NxuciYnBmqxmLYFT6XSNax/
bhdLj/fDu8psZsw0Pdi0KuqDCF20cD8CbJQhhUifH4Yii/llSD7s2J32B5vje2ygdUHut5RfLb/L
p1uQqqisXlnKCbiOEc0vUr/dKKlW47JzOnvKwX8klJSGAfMizQsjpwQQ4OWN+JYEf1x8Zk0mFLNo
Y3NEnxO1PpKWbFXnyMutY0Md0Sv6zLWaRxbXCkjrDvx+fcI0uVgxg8WEntH5+bNq77liD9LEkLrh
P64rvl0KfHd8PjLNdBqk7DNqbGXT3w8NZ9Gus4nJVBA6ktBWKDjFz2QU+/UcQeJMtQpHMvfBAUah
GnXSEMgjOnH5prJhXZiXjctVNH0i+WnY+N0acOPHSR8mguyEg7Zwo58J9QGoEV88R4C/XxT5e+14
LicrhVXnfW+MjL1rfgQh2JzWG5HpGxD2+AVATax+39Dn7FGqkKF20omMnKDAKdGu8YUIXwVHIIfD
E58IofuBXG2h+k2Iel64WcahOVCcOllNi/cEXxO7AXIrS8Toku31frWSh4ihlZC1atPmMi6jLOnk
5WqvduXJ5/q8mG3PPFwYiYLNeGRKaSei9+PlokN48aZJisKU8TWNPYyiJZ2mGcsP6cfxqOnfcyf6
h/7BEmqUnjbS2mqBughdPc+o2sgRCPoa8YFlYPzAI2LezvXkCPph84RKzuIj/EMIn2jW+qizrg4f
k+JrlXuz318GDRnf1nr9EA7AFgoHvfzd5PWO1epQ7c53OaO49FaO5rp4qf1/QGJpeJEv13Obnt1N
UcvhOWatJZHoqz2lt44A/qI4FPsuYLZxWn+1rTiOH/VkxbUSIrKWsGnW253FZKpxJmkygUzdrAqk
t3ZoTNCzZEMDouo42xbtFhy9j0gLspOCSCDDzTYhZRk/xkv9DXRRBQa0dUgZvB1Vz7QiTX1a0xku
K3zvCHIXfeuAyV9aOVN1gdAxTpZQp/1zA8I+9mLV1mUHnooeZ5SntHUikZ8AmdLkCZCy8YWwdiWk
gy477ighlxl1NwWL2BOOxmwTS0x4ZGN3NyLgjSRhHUaK3txqimxIgUPXB/Sifwrqa/wXSHBU/iW7
wvUZJm5k0jYE+Etm99g6UlsrNktfJq24j1BL0RFftdK7lv76X5MTotgVrcKAWtP7JKc18N9Wk14z
o+eEmdp4PSDlAIAUYHjARM32f0sqH5ovsSLkmo/Nvr62MxxgrYvfM7Z7orrMoOabvAlbjZ29OCX8
vuxG7WDeEzvh2H5/WyX1+kA+xQbqoxDwyyd5D8a0i+J4B/PPwvbKP/n+19dd/pAH99TR4qHLQzbR
50HpGqBdd/cnsjW+zL4PvY9jPbBMq+mLom46OincW2IEsbsvhCq50rSWWikqZVD9XTb27LgrCiUY
vRtHsbWFiOd37kOnjKlToijllIqm0naLsTEbeOKQWQhMA0SPhJXKlT8yblEJp4Bd3/2Ji1iw01Rl
T3owbbQdrUHd3nR5+UPe6KdwIeTJZGGbC+C/cY+QELlVakTH0nRwFXOkTvQEp+Uuk/aiOhM+HBK0
sU6jP4InshglwBnBO7fCvXvmKk+PTn9q5qrvVQQjD8U5RLtLWXuchrS/s1nAui9YhM//42CziWmN
6hTkSk4v2YqK8mJXENE2Q2Ms8zEmSqHzX3PWLVU8+rpHwQxSrj411gwxP59hzrDwosgSswqGEjn4
feHtb4VpvD9+GtVhun8AXrXNDCYWL5FXSU+RD+0fr9QzR5b3KAPypDky/nzcFpr/hd1iNPEG2btZ
Fq9fpo7jeuRlTTEDzlWSUzYuEy6dT5Vr2AtgNnom2qsaOiINXtvAxNCvafWcu6LgckD0ZrZrnNlt
ezOpZbLbW86lVYK3MgcpDYDuw+WrUi7gqndq7rWgRt+jwU9TTX5ISUjD4MYq7OWgY1Er45VUWQkW
eRCT0rjY0rgoDWDUt+APGqTmTor9NgxmHa08xA4LugdwnI87ckBGMxBguTF7+GTmbQti6u6EjQB3
7dNOqjwniMW1TPCxBS0cpVD4rCDGJkmv+h+htXSRA2KU3nufuuVWJ9JbsURN0/HzVyaM4pvHValO
Hxho9MEvL0lZFF2g7EF+L+Jr8YnhMo0NbTGGeDt65UipY2sC1tE7iJ7ngJT1AP/vCB94dEQWvScK
/+PkGUjArwQC6uWMZlAKgiGDH367iOhjXOxW8VbtT/4mRZ0AA6xHcLBgEVdPE9TUJTUuBVTvinya
315aX6PrMYBvEPY7xR2bVqkVQyXALrkfYSJyzoOhGNsTfwAWSOVBoWB4IlZiyymV+B6/2eA47BzG
0JXHZ07mhRmY+Y+dpRl+yw3IxKNXr0B2+raK7CHzeI4M5UgYQYUnJjzGNGY+aPAI4uQ8ZQurBwQ1
hHynf0NsTmp5Aue7x4rRAGMWGZfJiPnfOOEBQi3o6WM0KVdVJmZN7BMwlPT/EcFC/XGrFwRSYWzK
5mzmABopdr1Y/E4f3ssWczrkMnbBQ817rCq3QxqRMhTZ6uz2Btjv4wazzntAcYY2RaRwtqKRiAb6
xiFVj6T1ZMdM+UDUALnA5xQrrcBd0HO7nI80rOrtaWqWBdfljkCupImAqPZ9Fxz9HJEVh+ELR4da
OBmqNWNUvrza8SLOjLr26QvjWk2Yf65AtESYSmbEtWZ6mAKjEKRsUP/TKQNnoZFzJW/UJ5xCFBf0
wLTnfHdEpYO8sXv57rRWW7kU//5FHTnKQx9H+i+aEFBOcY8Pu/iNRwYAwDsr7hfHsm5ee4vPH9ma
drUoj8YayjwhEcUeRJi0uqMnzzb1Sdd6FR2GofEBPaqFBPfS/aNSvWceG5kvg820QLCdZRRh9v5x
Xw4S+JQjZBw+XC07sWM85F59jD5rfiY8P8FzHv5J0pPr+Q1n80gqi5YfJX+OPw3qQUofx+CMefWc
EHaMSHwASmBhCJrXAJK1dba0lrUcgkSkvNeCgGJHE7EvyfCuHoTcyzgmZviofKw7ZaRq8B7CWCXr
dtHXupfifImTPUlrR+7+cJ9RG4sWSD2L82gkhQrbaVT9N/yJx8rIitC63q1LSs8x3bKt38vBVmea
U8BQu2G2kL8/yJy7GI+SC+lyg18K246p88mmPXx30EH9GJpJvb9U3rI4HwGwulkJPUlVn70Guftk
d1HQdswZkWTzTp8rGAN+OwXprAJTfX6MEL7M5LE7ocbefIftNLls8w/x/optuPm47P6bfCCw32C8
kLzYC5dHiJ9RugAv4TTIqPk82wnznfOjzl0XuWKDgk58dfixsFXGAmh+ooLLwSkCz02SvteHKlLk
T0uFiOMdzB93R8w+FVFFHzLM46HnLaxuaV6A58L2SsoAIgMFzPbojlyoAp5IxYtgJt9UfPjcdrMX
sX3DskODRdmx7JFN++t4jkqHY9nDPOzTOW8tJqcx4EoZnNNmxqj7i64fbnihKS4lAXUV+kn7WEg4
xymmuhyt0CIYW1i3z7scbinoRYEIrdFqxr7UglnmWNxRuu8xZ/Ruokp4y0abzk82VtFZhiQKFo3G
C5W4m0ms4gZgMVjn82T+mP5CZrsIo/AqWicxpjHgfzyOBeRFQPwgVyIC+4Grqfcym+QSW7zUmwc2
m9dnlduwYFCQU+QbXaYFEbDBxKvXDs4dj8v8qa4pdlbRQ5vnwB/rmqXNWhaN4wLWg130wOoftri5
HrFBV+KLBV0cXSzFiuZF+o0bZFORU6sZQdyhJANQgM8T3T7hJkv1dfY75ANn0l1QadyKltjSbKx1
KYJpqjdycuBzprazNLmEJU0C8Vi6CI5T83Ytgl/H2xrwkRNbMe/mZUIDBqbZpNZJVFYI9Ba3D+aw
neiX/Rba6cpC1pO1uHN9yj+9tZk6P0yIvN1jxdw+KPRUZm5bjljjVU3uOoH/Pbe0vVYQCDoZIVNS
E/Qp+h2/t2hfU6ubywlY1vuFboH5d2jr1t0qS3IdSJJGzCMZH27GanFRJldNzEpYtNYSbmoS7NaX
9TUNMFDhVavugIHzCNEoYTEBIiddcxjfBmXPrf+teSA3W7b0LiQh4Cz4OHxWX4mRougVskx3z5GV
3ahdhfDMnQ+AUmbR7N7HrTPMRKDpvbRjPD4m1Qhp2XRRkB0GdJrIAem8mbjhWun9FAhBcsugZvB2
2bDY1lo6K8UNwQWlA90Y1iYW28oUHGBNNggnYjjdvPsSFnWlV++CQkdefQoYk6NlKw+r4/hJ3hvZ
SPNQcC0SQ8ajov1ogil9Nma3kttIicllLzmqcD+rDE2D3D7C2eSdj5CVHIQ7Ikm3uJ79ZIx6Wwt2
+n/cXZt2EfQEve2B1HKJZuJi6KN2TGMGxAwe8zt+r3rOt8AX5tNgOErJvUqW9n6wWkLvGtw0xe3g
JD/qNp9DtgTSx+a1dxEqPp7ewj1MuR4+5TxODtYdW13y1WzFd81R2pnxfgg4J/Qf2NZPA9Gmr/wD
Venh3JH0WJJ9djaMSKHc3CkpiFTaHwsnf7hCnkWlQeVlTfe3LKar4lSBnZ6Uf/S1Hr3Mqpu3/6Vs
/Lc2PYg/eAnKi13zH+QCKA/IxvS8LHkM7JEIlfge8ay9Ma01OPTVMXIKxfjqEbc+OxFNve74G9Uw
txIPqywaDpUqao5Sc7xYMwb5WUJGptPLa9SkMdRA5EkP2KyLMBUWpi19IKzZioWde2/VH9pRBJZ/
xfo3LF2zSOv+PErxC6CQuVWgPfKv5ASn2rz1uXxTxojYUZ+7Y9X2zbCR/6AqjP3QNH/ixH4Yq1Wm
PadgXTmKiByUq+7/HfDQyIxCEG1scdoyhad7P0l0+dd8CIu4gWnWsbY910H1VsZ44+c0SgCi4HLs
1mkBteSwL4lVla8Mr78exo+AeTHYAjRO7t6zMtnNMJou6FDmDjwL8LFGhIrnVCWEQSJtXckbrw5n
S0ca1u2ddpddPjphWDx/9q8Zn9NOpz7vc4vOyx2hoiCb1thaGn7SgWuDpQPRu8FkDvgMS/HkItmG
xFMmF2FsE1/UFX5tFGTUB3/3hLjxSgtMf63ev2g6m/w5ykyU+Ar6PR3tPNWT06KyGY6kxf5uXmN/
waM45v6lE4YYinmyxyozBXSjKG2P2cYtpn0H1MFZfTr0rtpneaW0pog5hy+8rHtBoKmgNVBUQnuv
f0mRcAhUzKBitJegy9RbjoeVvXXUSogPmRcnmJvHMQoPFjEvb0wI1QEYTeaSXaJKe7e4nF2i8WDd
nzgQW1oDnynJpWLPxRGlKC1QRlaRR4hR0SVdWhpfC1tGKR4nDS7BhwCwSKzcMDjHZHN1uM1lfki2
kiDMbwGKp6QzRU5/V2qHHBg+clp6i1ae1UdgP3EpTtgxG0YMZuuFLXnX0lpAS1WIkdNPjw1Dne42
VwBKkzCCbrpAJFoNa0IkkNFZCtWpAI/AQVmH6M3vAopW18uiho+54ivUED4mzgpGwbPLtUNibb1P
uJtvyHELWLmYAcq+8LVBZNqM29SF6ycVLCpeWYV0vQGSBXjbnT3yfllUaL7z/nGan0dfDJe7HVzP
+3Pmq2It1zJV91CHocCgcI+orcm1rkldT5BFYGPTg5rP/a5+0/I2Bx9Fg0JIB70GjepTf9dvXwPE
GcfeWC3V5rAMcK2ca5HP88Z8C1V8nifVAmOjQQ1tQujLyPwtohBYQu408UTxlE1bu25ZwlCfApIq
ZozIg0Q4tiE/hkgGZaLMthV5+JSDD971vOazwW3tcN7IY0IAMieBvLEm+sawBQwc2982xjM4eHED
iVuzHqCsKuZi6um4b0ZUAuEqqkweMmpdk7ah5Wa25hRvrudgI9DnQU/6hP6Ef9O6fTUnJBmER0Lq
Xk+hSOvtuXEjMNFBchRaMpQKEOEzzrstpOEoIAa50hGS3/fk7OES1+OY1n0VIwIZndUBY8vv7zOx
9Wi/gPSsUZG4M+ohHhSN7Bb1+3XeUMVMWD3+bW4iG2+fOPoGFPgvLZJMDVTwe7KvOYHd5jr9r4SC
0+t+Ltk2sAw3cfU85qNA2yVuB92yzpXsrkRhLtgN2c+txzrSyviyDBjy/XkQoicICX1mvac7az31
5j7V2ZbsOuYkwy/PbyGFk0I8x32sbywXEqV4BskvJY7yUrQIonvxrsDViOW8dskWdL9zbKm+CLO+
U9gAK3rfY6zHFFDXR81o4apma9rZwP+NJb/NoiqItcGzT0VZ30vHmh3XNkwYeTAZRulJ3ddSVc2b
iO7na14yeeKp/W8ck+661d+/Qjh90ZmgzJTgYtPgAJplXSQjyh0OT38uRcDRFDMqaaFOGH8KD4P8
5xbM/Kliq/9yy75c5sLbt257Zsmoh8OSLvgLtuv03jdvR4CnfXp5Ecqs5Kk673AHxnD16cp0hokj
MAnVZkiuyzyBsOv0gigDu9veocI0BnkO7epObshaBIp7rfqLGgt3xU4CE8HHW0IYBrlaZWI6eCny
mlU9yCgVfpIhHBebjC+fOqIGYvOvAYuIjlKm5KeIsrD1BeP4FuIF2YKpO2HVj4RTPP+Pfj2njQDz
ELETPOxy+ZjpIf8l3gDr52qgSDhP6kb1ImjKTgOE2owfTf6yub9Kq1bmFL/cNwQQILZP8HIqgICO
V38NeYFfL9Z+c+N30H+pB9dWZOhDIJgqHPDUQPlqXBmTwlzyw3TAnTEDYrBnFd2bUKjQMCq28flX
wl/OpEsiaa1v0w2Wg+REQFJ+NwOcBea0eMd86WZDo7ydEnB+5RrMgDsgdlUF1MWNXoUEt7+HPHQC
ITZt7NoHMgFdljuMuBZB4NuS9kvXstPMY478BAItnU5c2VoMXmOodd9GqSEjdG1stIEjirxMsAbv
D9LPNtCX7vPARWCvCsEXRTsdEJJGhFt9g6oAAN/ycT1CeGUzzOHMCo18FxeOfPiG6Txqi3B/8Q92
USXa3T3+1YqzgzBxyFPJQjEuMxMThAMssHn/NFTHHeARZmoajkM3gxPxvJG5PjhE1uZy+uVrZwkb
svNbvU6rq3vZ7Hur43jzz63jKGKwuTWH1EtThO7Ch+t+RL6toAttj2bl0eMDSO6QFpdhKueBhAHL
z1eKaelR2ZiVg2TWa2MD8oPTLR/NYtRp6kkRggYoyiy6V8oAxwveATWK6ktnJJgpakGghfPjuPuq
dV8hW618l4NgKXTbG4cUPsJeDdoEl8myhGmRLpFG5xdcunNYu156L+R9Cg8qlY+fhXGa91A52opP
ruii56h+y7Ekfj6Y67rAAYmJDRfcBBXdq7wOecyYI/D/0yBcYxvAqquIuHItR6VlrTGH88rsnLRb
V8sPt+l3oXHWLFh+5Z3Igq3QedhnqASx1qwQ5E5d2iZfCUbQ9gZOuhDvJy+tZS663nK8Tm266SeL
3rOZ7VJ1IH9cxgvv6hqhr+iq8zxYWY+OgKe+lYkMtPiOK4ngkJR2dQSbMJ0sMmx2rpVIAJtlgWcH
YyKLW9khMXoWDAzpM9veRAgRkfXTbCZxDIkhSQHLka7Phw+oOhEHxEwFZ6KTx/ljLXB7FV/KNaGp
ZLzryoGnmO1Z66M/xzkZpgqq/iLq/mphlIEK7GAAeg3mjq+jhoEbmlLzGRClsh4sQjcW1GZMYfBH
2O2aU2oWv8jAgk6i2oDF2MrCc3Jwstlx0jwoI4p5nrtrEDjEA3Z/0JrgjDSGOP4mpVw6GJZ23o1K
+bl8DwnkE/KSX+OGh4eo7jWTsIqf7Nzmu4OGe6fb2AJYSDAhcTL8NLE0RSqxYUC8cpt9USX7emAo
56KUmJKR04qpb4WynMD5Ulp+LR5JRKiVdoXk7MapGjQ8uTMCOvueuv1fSHMYGxDnv4VtkpyNStgh
GiNasKEOa4BasRjld02BVaaVrgowJuwKr5+Hfh66CCmJd7t0SvBvWNWGaDf2pxJkvjezjX2D4Poh
ztHXpFSx/NC0xBHh4hHXjZPwbBcwrePzrDaR4nv5jdNGJznwHPM3B+0BruGysFuuw1I9yx8K78NU
CQW0e9pGRy+DQizeL+jT0/u814bsOiCJlLfqMH0WlzWkjuS1AaWl37d3PKwRN15Uabhqrifjdtol
BRn6z+8PixPRY9uC6Tuc/PyPUACPkej/whNZYOQYeAvyv2kTY/nxcLshQaj3lCqnz7hlshblUhDW
Ql94RTt2sfIvEFCuNCC7KaPYe9AvGj2AX3sOblDjnxQgcGOxdz/pHN168K97NgwcE8y1weqtpncw
CgT3NP6QerY5RyMd1rLHYlUjZfqaW0ICwJmaUGcsgHuyzni10nTNVyA4pYaK5eOPPpP3QLhCbAc+
3Y5oLiWo0y8mg95eZ18vzN+lOWdciJIotA4aDYQrtbAlcYVzKSFEYYMa4V+v/QIPPNs3shD7TIiL
HY0PC6ausEv0BFnKoqLEfutjtHQUH6nRbX+xgyyxmgW7Vtpe3pgrkPsjr7/N6TF/RTxrVxxe78iK
mj50LubaoDhm8AtVKG7Ksky9lxQfz0NEazbLL4caIO+ANAfLDoAyy8WRijqHyR9y2nDVolnqxUs+
GUSHU7Q346vWt615d7D8FTRTu97+fce0flrFq4pw5GqHFDnFbHTqPXDuo1Kxowg3Xc1pY65fgMiD
FcErohb4kD2uEVDaieV5Mc0JPtWUA0emgL8l/sIlBvDEPh97GluNAOfkbFG2p7XxyyWk4dHV42Ii
tR1gYimJLnuVb4xl6loJXvnXELnnsmCgfZKcnvQQUa0GZFHx85fdT1ewXPL603FAfMK2G/QRhc14
yHD1ldgWuAI/o7KvP0q+NBRfxKvZ1myT0zVlxSlMDEQnlTLJv3hRewCzxywDfoJk7ApdO0BGy++d
iCctXhROOSi/BMWLoQeERe+EYasTKDnvkTg6McdGuz2hC2OG48Wjrxlq1Wmdf5v29fa+MRQt6p9A
ICQTr7AVxyoMke26FYPUuomaLgxGmNc3MLRi/+96STs5JrENsqwZFBXFnYd/+E+Emb8MF6mXX3eo
FVkbaUJtSxtNDch0XWSE9JTvi/4AqOgAh1shWlE5IfpS5UHxDKdti2wiLVXtin0Tjtf0AyNAuGA2
Ktxle/xzFPKFJanhWfDhoUl2eJ67dnxDVS/NSeM2j3oHO93LbAzpQiQJok3N332T/1wf1m3N2rbi
dUukRfmwYoczo2cy+HOO1NoJS4+CfJGZIuB/CahtQAaEXf2rHHuCtZRTQK3gxy63lgx4smEleVc3
B0EKE8k2PDfj1rSCnu5/wI/wKrqfJKG2QjaU7x7aE8Fcibbe5mDUz1EZDnZYmlU3p1etqFLHr737
sHjSTJb4wYbEAmWn5Yf7b6edO4SEABghzK/S7CLs6ci3m6LlES1Ot831L18Bmam9JAEUbxTQ31rz
ZRlycubJ7fMOkzDqW0Ivg5g8Pm4DF3jERytAhF1DETUz66bY1CRUv5ToWNW+8GltarcelsbgTTyB
xQ4KOsJodqSdRuKr+2gTL0e8Y7ddi+rTX2GuP0Fi08wfbQ72DZsx7u4YGJiQDQDdqFU6pzTGRLNN
SPuv/XUm1IlXAhYNBHIpLZWghshiWbPsYpwnZkvgF1U3CwV4kRsWWF0x/jAk0qXfVOe0cb7iALyO
mRKLrYgCSp3LYcP8NegwyszPiIKjs9T+ryrlkRNuQ0zorc9fAZ4MB3sa1uOLYrBTGOxQvv/qU/Sd
0ZT2oGBEksh4NyD+z1T29NxDUDCPqrhYSg2JnOvW+RC62Er2xEb+3ahkRTobIPEsMvkdjlLyKP5z
WvnZtv4oXcWDdHEGuSZ5snQOXZ/L2y/dzSJJCN8c4d5dWdoh62hkb8/dohoUP5IbZpcTUtC/Pv2T
0B6YNOMQdw49I9LCbau2DVJQup+s1RYPgwjfAfNvV3hJn2tKwJ5cbn/GZnxwUDvOKd/DnCgNx3d7
5H3whcoXj4da4VcudRg0VxooqWCbXBD3pOZ5aneSAOe+1hKeFxH/xOWyZVWAOmEiURWQEwRD8eD1
cm3imkoOKubTOPW/58reOSVtBdBZy83zA7wzjKN2aH0Io6tTI3ILyJIQoLd2/WYCz107Jwux9p4F
M+tmBlyardnGqlpKprzMz5c0MEakX4XCYIlx5ERtXo9PzcO5dkW2Og/B4TH0uGlT9gtn/MQ97axP
+wAdYURgsRrTvMaaGmRz+EBbs6F6c6rpjlswc1Yf+RGEuDaEZVfTm1c+iPmhV5JW0hgEQBw46Ygt
wHNekbQtUuf1/VNlnuwT+suOhfkhq+A600huWADyaOp2Rxgv6ttu/yg7xABZKvYSmWMM53yRKf7E
OZPKy6+wYkg0zYFhSAdKEFOLvL9pn6c2MGECU8drsHnI9tnsXPw+wi2guTdAP0NbraoZVwGaTd1j
EJXxfyKAizGKpz3lxVUgoGpggzbsDyR5/a98sMZgExgKJ1lr5vZFIuBXmM1X0HfBFB7MBVVfiYnl
bS1hB0YCvQfY+W9kwPk6RhSdP9/3xBHWKi8cf36sdFL89r7a0nj+snCOlCTR/+eBKluxBej2YMsU
HZjOX90Am0kqOrgBdV2DawqcoDfiA15kT9PJyYvc8aArdZ8nsuSP2BtpYSqiwOO17Gj4nBDphKUH
+xg6RP61x25MkzHyqex4PJgS8//zp2z6hwd7Yq8RSeusDyWpKr/z1Nx0eMPFLuHkB+wIVD1EFCCf
8/JG02xa8VY6IYu4ndK3kfs2cNVcRnj+H+zXqIqXNy4GnreIv5urNU7DNaiUXaXiFVeY6/N2GdZD
LIl33dYTVzcwddUlVKfOZqoBJDOlYLiii4xq1ZgON7wpgPYJpyiAOOqjXDmaybOhdoN8GK7FHkgT
HvfRCcrQa5uqODDkJnG+vEzejoE73is7nnD6Aee3la7Tuey2oMcnXqDNdqHFoWgKZkfpdj9KahqD
P2NRM2x+IrMrdtRCXU5Y+YQmS2r7boAXy+s+lb3VHWOnizZBP9DOHCq5eIZnGYxw2WgXSEsKU7Xc
8W6QXFsc8BXGEXAilEcFUnT0pgrtHHZHRL7Z2nJZCk/VGKxP+fsabY/poRlQ0zeGZCxGHTTJnXZ3
M8ZeGEr4lnXtPVtr0L2LOXYgPP1fJAZzNtUnlBkJ2R25ZQFaAeLMx/GUO/3U7Izj14vzp+eN5/Gk
ZIcoAU1qJFt0Mfe7a8APo4tmx3lp+oPnva+gbjf2tx44Ve+sD6uyx8EBUDsjlxnUaeVpKubkfkpb
bpDhmPp6V6zIU10ZkelO9cOiEu1c6a6vh7UYJ4Hoem9oLv/Df5CoKc0WORKLpRxkfsBE6d/BuZda
U55jIykjAdkyFzilhuTb2izUBMolPBzpeNj1me+3qOLoMFSDi1faC3BwUlhFuTDS8ZtB1MsxUnFx
wZCc8Z8KVcTT3ZaOWUCtlQsuunleSblh755OevmvaO3RcEkzjEB2iQD3TXXe+0T6l9C1/RM0+9Mn
kbZtvKD0EaH6R0kIt//+ebwrZhQ6h5ZbFbTy5K/X8V/EHF8Xm+DdGuQ1GlCzi1SKUr/k5yrxgp3z
vNLNDYAq96lGMPyXheLkaoVeZs65xYHYNGSrrbv2tsunE2LR7i36wJ3klRZnks8c1cBhw4Df7WLj
qeU/Y7oy+xUmnkUj1pYcz+3xmGFeer8Ujns63sm3xri80BfbufOc43QoH7nVXkD6AmzAAR9G1o6V
msuzrYf/jyNNPafl5naENludshTAVVqAVu0k9SJ7VNxeNL6LBtGDG1LAZZGazCJ8MPJYlgQ6mKA9
xkdhJVydLL56sVsqsSf3A8VOezjQGXQNtsnQiIkx732oYGCMrr0nMLhOmzbyrkDa5WH7lX9AEXPT
r4fu45MTrDb++CYhTDYJWM4RK4rPyurkpEyFCQhobYm36fqXv1Ju7dFGxURkCGmHQB+bLm4hy4HO
w0xdeqxBps58zY9Cp35BEapsx82ef5WwRqUt0gwo2jMdQFWhFpOAkE/XpUCIppBmsSCj3HUMAc9u
JeRVeEsAhIow8LZbxYPHAAH9HJQ7GZc/dLTxKCM2OcltbA57YAasUTV6zCTBYlwvXFiqVCDPQJJo
k/zamrz61R/9l3OFOehQ+J1ULJxH9bsuC0pM+PoiI2N/hqyQ+cL2rOFrHkSiB+YRD2vU/P3+GqL8
gEUXEFdFFcpSUxJcIgQC85ntA81PuRoH3nVWTxNHGupJN7IpHg1ybfU2W5qQlr5e4AsFpaAWLNt7
BNui9mCeORjrTRC4jV5iI3l7+F1nIhzXc+SCfATV2MypGVDYuoV8+F9OjbIkxDqIFeDgDylzlPuX
3jG25o3SULxkMpmtz/0oTEAWm9LkucEhXSjRRMrINRCCL47KIpdZwxGu8lLeL53ytxxqpny9ePG9
C4aWaGmuskkjxoLjFOiBSRBzkRJmyNB1Lx0dlza3x8ae6iPeMwRO+2Y/U8SeBAHEv2Edg6qzAq1h
SwE05hnNjyHLnJBZmHsZsMJqktoVGRvmTlbCGGeRAWODP/HNaCE5uha3T6mcC48OERdm+0fbMK6P
mhktRL3fhgdI3jFEGOSulE+LL9ZLA0pQM5m/+cbdnzKV1VCx+3FV6h3l3h2c4AU8nqO/gYOYcxMH
3Ay+KYbd97pjlVK4jDGs0PjueJzFOu0lZo9cMJW+mSc5FDJw5NcbPTdxFi6vi9ajDav30MxS+p+Z
VmJ9d+Ym0CddJdG/u62A6sMBK1MaR+2zTOgvvZhSxODXXdfVayClizsyPRGK7snYRgLdzM5xiVLm
rctKAtrJ7/1+yVlSwNBu4u2vEDe6b8b8V5E8CXtk3vu1601v0m3W90sG7h00TAfTUVMZuQ1iqjvR
K2t931aiJ+EGhaUdqHvzO0KH2xVYR9uVOfG16Sjn3l6SvRo5jsEgrVblhHjs6gycz1Seb3begXJ2
1NBs7LMGGRpbkFjfkeBN2xrHjzrv8rsOBDHAs7+CLbCdJVuFiP4E2o9N14We9tlY0MsTBaOxcjyd
eJ5YltX+XYKBy6pWtYznfG/7XLPYAwlBq+iuPG1WWzIs2c8W4Wbe5OHkVxKzJ2bqc/nx++heCHXX
x1NTq96feUktSWxEcVFR2gTbsg2S/8SxDt9P0fO+MW70IT8KgN8k8kijISgs+rgbt+EL7AlAveyY
RzdaC9DoScTrDZsJMIIQIgcskc2UpLFAEIBAAFAVkVoF2c/XDzH4LPRX/SmWy7gIuG5KrD+fKktg
kO/1WjvuCHCONqucXLYojGHU+uYv1RqEWshXGj4OuQDmlWvpTuxaXMh/XOcjDrxREa3GkPpw5qaq
lTdsBbLLRC1Y5NyfW7ITmVvMtLsETllcwQl8eCpMAC27RUceRA6k3764qw2NKAn/lua7OiXEuQvS
c1EHoqo9R/JwC7q3FjJMmvHf7UK/N7MGiP/2LQ70gLF/3gePByMY7hwg4Oi/Fc+32K/Q0+j2z7S7
vtnOy1hFEiH2yIc2KZp4rOWMUzyxa+jb8jYmXAmNfc83bAzhABCQvkrObvS21Ef81/TPtJbGCbOa
y5y0/XA3QbF6Lmd65KaFu8jTm57KnZ0vjRfqtYMa5CCBa6O8tCUkA9afkR8UbBVH+DYPbX+baYzj
U56+b5E5VoSnXK0WO0dTZlVj7k5cIwl/bgeKz9dakd8JzZ4mTp8/mawH2JqLfgPMOuFl5ZDKT5hH
zKTVihjrYFuIoIsBNwqrM298vImltpQL7zFLszk7DW+AQaJyxxSp5zhKZ1IyWYYOpMR6p3vpQc4m
XzwoqTHXr3ArJxyof23sCgD9//lqehZE0CtppR8k1kXh6ajUN8E5sEvvx0nWcmUvMbo4b3c5U16s
GPZaOrvFYGFZN0fZWkqSDCz53LfZpQvVz7V0OYF3H5j1vKHfb8vqtGdvFPByfPtrhY+pqvWNC+9I
eNvOTfV8y3Uv7cItQNEFeB/3i/MdKFP3KFvGuWESOdiRIIsKnTmzi1psWgYUVVB7h4IkawyL9pn2
aVT/Ve/kjVGVARiAfxqmypI4pj1pOI/hzLXQC1AbWm5nZjpkP1lJCskU9nZ+mj1BnNDgXpZkn59z
a0ZUksvKysDeh+IuOijdpNULWmb8UGDij8IiJg5GKBPDsNwhDRckPSGNp50XSrCVPRrVgiDRuQ2b
KLxTWRj1tfs3aYYp+qyFpS1moyCCTBs0TRkUrNpN3FgPZ77R6F48RnmoFPwUqtxdgL5dpqtxtvvX
ChJtLIiU75uGkmvpV0Do3Y2u9RYB2oWklr60cIrJQvXbuTu48zPMFwkOluW/vggyTPa+Q0I+VcIE
2IIp1MjX9+y/uHya1ZI8UFbUotYWBqO2klwznSR2Km4ag+/3fANnCU022NXo4o0dlTuXkWj71FxM
eS5NyCzNzXgQNsnzn+x5A+9BRW8DGx3q388BdyhqO1S9h4qq9cXYIgr9uUXWb+HAlgrrifNGc14K
komuFA1ykK4Z6tGimBHOOLy1DVwz3hZXLtb8VC4hPq1+BLlK3S+ZCwzHdodmWy9DkOTY7lbxP1GC
s/lAmA2HZqwgVBQ8R8zhgVHAPleQLeOebB69FfzdsSMVJz5BC2MJe2eUbIeNCZt/d2uWFSutVSfL
UA8obcDDRZNmz3UeJPpgFjNnS4t9NOxqE04kDv6Ie4zkN5Ewf2YefVnXDGI6zO7hE9Zn6Xz1JwS3
YaIVzyj5Cn7FroPjgRnmDsMv9z9FrxE+0z/V/Q3LjmJaMkriAL9Ew8MXo22jmrXoMjp+2jBGfVMo
EONoIB/LEqcuReqtlBuRuk+Zf71rYPdzMt9QCYunT5DagtvcbpdYDKbD0G6PnhhGeQTJLLHbZTda
8HEYFWV5Vzld6jM+JSvEOgsY6B6dNPVRaQVZDBZSU1YKBwZ50lLA3Ii8BSd9CiMZ/jFpzI62NnyL
/Iw2unEfDATU3ikK7TpGT4IxaZd7PzVTHtid/bJQ6fhunKNNrP2dhdF/pkcm3U1wIGVcJG2OwuZJ
cz5Z41VDLLT/v32nib8XLzBsoPyfeKwcuMHnryFJzTH4tPTXGryvG5ZYziwGJIlHlrAZgSWvqVYX
HHFvyDui8jSWF8FtfADvxS4bTm5nCdIodkCOm/B56wBFxyoSG7fePY2WlBgom/WP8dW2T/FQjcmO
bUDcZdAcYlDlaQU1whQBKjbeYrv96dPvOq0GJ6Z8d4K4GVZqMpRJinAiPWoI57NZPmmQgeUaqK40
O9PeyLp+/O1P5ZxQunDi31UWNUsLvze2CsBX/2DHew8u8arzA6Mnrx2KcC6nx/dNlnd6CseIXWPs
uGWWRE15VuhAoq4XHxEDKX8/4N3VBDRLVVgGL+7bQm1yQAK555UWw546k4ZvyclPakh/tXBT8R5/
fYMFO0M0aJeEdcq0vigF7TO6drIOBlOvtxPw1rQWxs6y5cde51e4r4VVuErX3gORK1brV7bZZTSU
90VkqYmjFFD+5Bgrgrc8YY2UoMCDKPpEdbN81zxQv7hNJF8XvvOV+dXAKXYbt1EuYXWlWCUVIgwZ
3AxHl1lX6BvIdoxQCoRkOksWHlbkQNQux5BRFCSIlLR9oYGdqbLi3Mg1bANai0VHM0JiHOvxR6EC
KyOja6mjpG3RQ2r545SmNuQ09SZGqpeMyN8eCSpN4jpThZQYkWbNrx2CNLpxvoKKpYo6yGc9yZ+7
kzxVR6ZcW+39ALcKPeyjFY5hEMNWgy/Fn5KzqarqO3HcEgV+YDyyS8T6SbK++sjxa9JO8Oinhxw3
p+F+2pAmTdSFtw/8W55rV7K/H6PWbSqWbZd1A4AHJDoCDgw3oz63w/KFEYcVdsqq+amhcPUASuS7
Fu54fB0I1yERAKfa4TyChlCUM+d5SD3vn94Zz4KisLPkfgEuIIiylaB2n/VZs8otpQKPpKnwKl5H
6H0zz09G1vls/UG3HubvsWkNx2pNEwuriT9YOtRlTkw19deuCtBp6nLbwKdn4eTGNubCA7gnhqcV
kOzFeW8WC80Sb5lw3zjCYoMjcABzuXjv3vziOpx0YKT0VRXJALsJEbVIyyWn6J9BUAOcKmor9YUo
bSrZ0Y185Bo+UUZLGrzpZcuFGFbKh6qZ6lMi2iUQmxtzsszX6G3s4qJO4m8E+JZu/Fg0gcrk4Jkq
16+lJumM1ulWRwXAiiXh+Mix0c6RNuadwhG92K9wa25EoH9bo/qlX50eowLy1Ff9Fk4gQXCZTsWB
Mp5/17BVJhyZv8v8DNxbmbw8qzve4uM4dq/4cxjLiO0bbdjo2qwWdbGPIP/NEE3rG2rjUFilt3GK
LTt2xdAF01qOdip2j7yvy3Y3RMeHXnelr9g/L3gP+Nd1kvqnt7KY98zCorQl32AfwMFB0rUTIKMm
Gv/K6lGOCOQjQAC0gG6ez+FOnhJzoTJMhEDWWBwbVvsEAYMfhU+mLSr68A+11UppRv7qvkdY7Dl+
maemwnvYC9CFCxH42MBCzbzuXlRbq6tLtkTtSGeR8VhtYMMgC6NlJ8VUW6yAdGJ3rP+lVYC3GPpH
m7hgtgReJQaz7DfrBplJM+TymbiG4TdVKejEPHCzOLnGREKa3NSyIWckPjflQNGLLZVpvgxqLY8i
QdE2QK8mIu1Te3cnGp9wzfMakWFqRpcV+DxqECaqhn/4YdnPdxt8cyev/vmUlr1WvYfs9xeBaLKL
GvTW11XAjelOmHVvif1vlDcbFWQNyXnfa0p15l8EVq5GIydZazAxggH/RdU9c28tjyeWIHwAePV+
jD15lhKL5KXWoEpUM4whVGg0h2fqxMfMTLFddgS+bd6YleO6sP8jdy9hN36ZOg4NI5CzSsESwbm0
kmKdObEq1cuwlcC0cZs7WGM8bwMvsxyDjiospI5+2VNyInnCbqyIMJsIRRkqCmOwN1FvflO0l4Z2
5rIom67q9NrVq8XlybF2u0IlpEIb+MBLXonsPdomc5F05yl856OdwL6n5SOjqcKP7kgYkKwyAIcU
ZP/v7rjICt+k9j535LKBDZnz2+3Bramm88KLodN5k9E1JWuDE2yGYTvdJB1mBFQk/bCOKpQDw57L
11aQ7KFBmokUeLaZPiiUzdQoGB3DgwdUd9raz4FQhj2Wkrd4dcuP/fHZT0uy+zV76QDTkWW9mDSE
8l/2LGpOwjtIgK3WwHrARdmx9Ma/a8lpnTt/jpcPJKJfayYaPkcFxeH6SzAw7wrK5xh+81tGWfsC
JeesuDTADy/UP7F7fuC6WqDErA4N0T56BP3DKov4J0CnFJUy3RWo67UusTzBlKTun2rinAiY53lQ
kQj2xnhaVxs7fC8+ISe0jBioLmPPOFt3+cBXCIpZa24RNZ76nvzlPwpdrpXisZTgTMfJUrCGqU0e
7mJB9Lq59LxF0Rq8gcdd7V9P19ngHc3Qg+ynBSY29jf0Lwh6Y2w4sGwOncFIsNbjmlhzsyCXCOvL
kIKFsb9o7I+HuB3HgqMI6sJa1ofvuO2IALeUgR4l7oTHqGGV8hdX+xg7RB7WH/Meydxcp0Xd51u5
pJhKcXsAVAdutAukOsdvCtWJpPzrTRltEWVV6t9zNao1IgA6sxioH/q16gh5LDr/Z3u/xwjnrD3W
x9n2/SQiTR4PvB3gEtlbOPBVJYOSMcg5dxf/KsgAm1gedL73gSjaF2lMhGVE34mxvZinqbhEM4K3
UMKmLHoIWFB9NoG32qbs530l49t7IXOoiT4NVAcjR6xZhymKl8o0bVCsTFXAbyvvxFPpRXNc7jtg
VkSSKJkboZmiCQsNvT7//yUO/RLvT7uMnnv6XNBcHpzm7GrG4D0mk7QAb6DJHnen86kJaATahgB2
nHtKIyG0xGNc5dmnjoJcTccp0mhGx8d46jqFgfpgjdDn5rokI5jYg/JQSlx4eCyKxDMFGOcwMM38
tAr3agc3bPdNrF+756LOlQgGXA/JRGGqi3WpjYxv3PKVRHI/vn4TAE7oEaRNMLf3xj4Z7Hn0M506
TLYB0fevpi+ZVrDXTL7t+jXOB7Y+HjM48uSs0F2eyUlee8amnP9U4AZIyAyoL3AAan1JvXpqftlR
LNqRnfAW3syC9yI4UPAgvQvTKfuSbmKh4AeGh9HU0LDmiHZXUSSDzjt1tPgNCJg/f64Gzhs5hFMl
H9iNjnA236OGZ2MsLLTqjD0FBdUOxkmkOic91/dK7qsU0VxJX0H2wMJM/hJ3kSYDf1jJjU+J3p84
KqoMhAaJQgwvQO3fSJNbDg14ZJ5IsYVTFRC1EXS9qcUfhriEPglRBMRa5y68B3O4ZNNhKcxbV4dT
7q/JICFjrlxgECpjdThieaQUIo8E4lwCOx9KXWxCF01tVTh6Gf/3dnK7GlUq0Qa5W396qPIWYsQD
eFFJMao8PLQlx/95t/W5k8m5PZMejzWkqSTyiD0PUu3uFQgJfZQ55RC5M3S9qTeKQQfTabVy52/B
kpu/ECEV5X8b2oipqtdxDB1GodfvW+5HOgkvm3OMOvsUFdPeRqEUYFdRGOqY8AZ9sx1bWPXx0TFW
oXPIdjiL0XzOZ/ayr461kK6fa/H6N23IlyZA8RThvw+eeVpelpW+GjrF9v4S702CpN7zqpc94tTU
0R1+rKwZHVnFtDU+RHqOcSnaTiOSUOtqnN5MWy/RTXG9XJ1xITcb2r/M5/DbBfAH+TexxoPF5Ims
lA5hHwPdpJkwVpOrrUQIJJjaiTwjdBK67dMm6E43uZ5nu1ZLiSR8pfYUV20WIJA+ujAEMBEw0sFc
6APCcYyUQMSpu7YDmN6lKQKN6dWQDexcCuamQvC75WM3RQg/RZB8ufrl4r65V6jgAtEd80tBSV6/
INuWji9qhmE2y33c9Uo/3xOd125KjYU5/n1uz8dNuovW66t7L3Ne0FETwuQZgUWB8bhK0Ntd/nPQ
RIt+nZaqYIluVvFKuj2BqOGfo4Keu6mG8K41k5xunVks8rMZyGUfHa9O6O+okGTaRx+Sbh9S06W3
iHdhQq1o1R50pvUsVMxS0R6OBF0j92my5ZbAlTeURj0usDw1snANTzLC/umtQwWLQblZned3XSgI
3W8oRBlgXeVDCEo9B3xXR5SNuNSHCpQqX1ir5bHzfMgBErCN3AVxhYzt/Tae8Co6wpWwCfrPF5Ov
0J6R1sdeA/yyN5rvRYPJEJhIAYDcvzEeMxJbNFsEi1uZgLvsGWrWZX8UMgd3U6alDWBA7G5W8B59
PBYV4BjkVkAYaWXroHp15v9tVOcJue2uD2nVOGEjI1Gm7KLvXXpL6Lj0gdNe8e8wnrmZ0zb6iitB
/baWSu/KY54ynrr4Pvi1Pi9oJ7HA6BFEqPHlL/UD9Qr0gXc1qhd0XEdq/nJCjZz3QR2Unv9tU/ps
a/FfphB+2rIqc4pWtmLB/WHL/jpuVhp23MKRPyEtpCmDgQrXXTUWbeli6tFeoC3d3hZ66G+nm1lM
88JSO2wpLmTXIrxtojR2FYmPR2YZlWlwLegP3BLYA077aDwlwMkOw1tTAYdJUhhOhJ9KQrsZM3uF
wKroiNeFpZujO3q2ItMJmLkDK1B3ZMOL/ppDcVLqPKxUwkioMNNTtPV0cF74AHQ/269EHuo7DRuF
pFRvl2HqQgRJpt6hrOvWwEpUILQFr62cnxHAxSthH+TLFo6xMlN3pRHPxoTOvZi2yMGVdSOiR33C
n2mhXHHla/q0SJZGlARDpEodKQFPajrP6Y8WnkBJzYx+vjmGC0U6dVhDbUhRAfviekcJJYCa9+wa
+egENgjSrylgYI7VfVPsCAQWQ6QLbA87fSyOmQ+FkkyeXKff1BSeOwrheD5h5jAc4QeyZ+EDjhv9
Bp8WOt4quZE8nwaVTXxBoJ0PzKd5rCJHAOZOxiJdAb9PqADR/Jyw+vCn+uKtCJuKd9UHmPFW+i/w
8k8h9njiqjcD2iFhA0lXKPwg1rpk1ze57ZN1dI4GZ+rlej+o8bTLTY8EHlp7VxqOegpMN9DL8o96
VY9BUNlKD4TypxKSi7BsvSD52SGNuam81W62RD2vOBQ/2NDCJlAQeumaVTmDEu7f8TtNf24vffKJ
x1TmEWlx8nAlIa5XxjdX8tvbB8paw0SsEdVWoSF746PSsNriSYuL3togdLWYlTMutbRJSCBo2GVF
TEE4QoIMYUl0PvQPuy5T8Xk/Ycugol3w6Y2jOPZZrSl4ymlAL6Zbia2Whgj2cLLzTzPeXjzr9eXm
t3Lki8GrK93+vYe2o27BEC4UYtYssfapJ7F6ERkLEvR5m6jyRCQLULYdi6yFPb9aTMqFtsxFO01b
oN1uvNf2nA0wHU3U817ba2474yPvZbp7yeNCPfB26JsG5cA7xFnJgWcVYjB9u2CjI55/IMOnGFcT
VsVW3QVufnUNMDoacQZHNOSCO9bgBVPvP0O2v5EhoYxi82PIdOnBQP+F3JqN2ZkdMWr1FBSSAdfM
GjPBuAbHDjisgXdtGFy9iYYLYiBM8cKOy5JiHtcyyZh6+wmei+ozZ2RRMNmkEpDGhMADtuS+KSGG
fLz7TLapHkk3eoAW77N/6jacT4joL0bNmoqpWNWhGxGg5O/WjBDst13LUKyEV8FJFgZOluVrzEo9
qqtP60KNsMftOo6Aava9JLxIfVOgVX+6lWgpGQ/H0O7386DEV7D5FhROsH6u35U6LGjc3V/eNjpC
1WSFD0IRNgbqC5NgwD36jACLrvUM8sDeBsWFktu+drcaSnKI14X0IxS6yMiMuE/o7n9T8Y97zNXa
28NCkViTeR/ic1t/w0FTjRn6fA6ENlSyBZnHgf+YAAGHPubvtpOzMmRsmeGXZEDPE18fuWRZZRaN
36O6HSPBK7mFpIqbal3MV2K7PAslrRivDXjOseGiZCjO0udQSAD0qqfPk6+tN8AaMQAzwAs82CT8
vQZs2pbYScSMWCtNpe6Pvzgwr6DNquOtzOvB8l7n2WoobtJwRUxqOEDOTQ5qQYR0xzlMFUFP/Qxe
8iqOioCJYu3m+Yg02i3J5xzF+g/uzZaCwz1VCvReOonMQYqWCehKCZPGFfDgWYgs2tH1cdJezxZA
xZhtSlFqovtavvhDWQCIKe+ctgttMnXZCgjSnsg9i75YzlW/1dJZmnVpWo2ITtHJMwPy64BHN5u8
qApe4sdJNKwzBKun4GwT3WoV7q3oJmZ+B1gPY+fn8vwcnwc5hcP1+rIpNLD+c2d23ppnMUGvtjtO
TaN/h516QyBLru8lXGwW2e7gaozkQQ9aup5xzD66jqyXtUdfEJ7G9eVG6s6JV3+zNTIcppmFe+T0
RftpnbS42GvKTNry5J2VNtCo33EwCsx2Fgyut8resfCB3q5S1wgcI7DyNNY0MjiwdzuUwmxKxppG
ni9gnAokWoLoPDJVn2idCBRd1iLH9KhYVoQMzXAZxh8WOk3CipVA+XrjYd03zNlVKaEZOoP43tMC
zhclr3yExYvtE/RCV0BYka4H7iDFRaA1rn1q6VAiNHVjTslUk3L+NN6mgP4fkW9Ka91PJkmTDtSg
yBXrKzdXf8IzMzaujdSEkvVvXuIxwjdQGC/jHHZN5ViAnTMBmTUrsY7j4HsuP0ueqGE5JAAeS+sw
j9KMVAfQC3L6VMdt9osKwcS6YB53qO3C2yhOo8G7QMN2fxukl3ow9IkyseHPAPfef5xqxLTL/5VT
SrZ9ZY57NhqC7uXE200iwn2GvpfqUduADX9jMtKwcEank/IHvdfDwPiAA+ythNvCkFqksurceMCJ
1pN2R1P7pRt40iDlEwbCehTcmmMH0Cnck0Znt33RgUHOGFFd1k0JFD+mL+vyraQy4XxRjqy5RTvf
UAEFT5e80zrzjqbXmGpuWmHVRoccmbB1OKXrILp+LGMN8mDP4Stbp7o8qlTuuKQFiao+oGW3wVB4
fP2bJLeH9R6x6QuzyuzFOwDBEUM0Ae7kBTdZWO+X3+PxuniEweZczDmxqjp5/X2c59Kqc3JSyj94
X6TCvDGHsv+8IrPmoiOiWBIa1WYya4rxojRfi/UfdwQWMdHbApKj8q9sXj6JT7bihU4+UTuCgSJ1
EbdRD1wNuC26mHeHm8wQWCZyb7/dP1jOu3WUSmJlyrmHd1HByizxISRtk130jJEXf9uSH/v+0BU8
LnaioDdOhPLxGb3DaO1Cenr32uTN5rg3UBSWqGPCWPEtc53mqnS9zcg/Ub9PaZrNbXbegwm7Z3Jk
P88mORWbg/MzNOMK+rmf7ug9YQMgu/jwT7LwkdBqrt4afXeve0/7Kt3UHUZCtzp3RZ/pHsr3wk7L
L3N89l+PFNMJ2S/+03C5eO18XVVotscs11LdGdjYtySnZnzgSMoryuR12nvg/Er3Sy93cVPYm08K
teovHAU9aJN8PYM3k8fEObfrjSd0Cf7pZQBG0ZvDZ4tqyHuQVwMsK8LcHNx0TgBhKDHZckqQ7q4W
xe25FAcK7eq3qJJXOYUDLY49j6dWEh2byfi7stGg/6gyYTevmTJwIePg8SlQKvbh+XMv7TKdiVDn
mls2y6DL7lK+SI1Ult6HTZe9rE/ppgf/nHydabZ8eGNwie0p+8bxgWjYzl+zPRxhHIJOt0RwqFUr
LyMyaTUICzQJWlQ8uXTOrVd+bgjSOAz1Qu/7gy8DAINE8+U3KG+w+U3JFu3+Gku3rfa2O4sQ+knf
8byJFpPIscPHMsDmOjjXwL+axo6BrGBwdKihxV+ghozGb4n5mA/sW/oG4IxW8P4UA7Aa9BNqOccv
IF/M9EANvUMhkK67dU45wlDNw3uHadFteVwmYD9RwDrs/MHUw93dggTGuvljndu3miEieCvy2dhf
84J5/YY4XuxR9bt20AfaaSiFh1tWalsXlAOgKRsZx9EuAB+pq6BtLUGH4uoFwCXQ6o20l9N26x1d
vnNBSO+JIHhpa+Xx0DEuDA9EUzEbNfX1IpKtq/FbgYlNnr9DY8RD50o0rebHFCmomM1WGTUxmqaf
cWi+fmTAsEPgvfM5Koo7+r8H489pHDCmsD7iNykwnluhF9GHQTSGYq6HquXINgd1N27Ck6rGG4JZ
h0wW2kRderGNzAyJDSqoRcyp8hzbYhLaS+VXJDFLDU8wEZbxk1jiXpSMqapgpe4Qcx0OltkxSqgr
MRBW48cpIaXb4sbsFtNapMqv92w1t01tmRNQcASLxd8TW74wamngPkhDjJBB89jWxJiMHv/puHDW
DA0eGwlFEB51uLQhVs93Lso7YGLx4HCZU90qiuvceqzD5Fs/az3J9lMLHqI8LK0kcoC7XQTnSSzY
1oRhiIi+AuGHsoN3x6/e0tkKogJb+afn2jEXPBmE4LQTwQKBMRIMNH3QgzHPPhAllER1qgoADUIF
4B1CV3FJyS/cf/tGCxWOuJW2KCodxAOj0DRUdFYiAjSdKoAG0bDxFdg7CALp8O9dllK+LwUSeDnL
A7eJkzrVauTvEBtdzJwns2+J7k6MVbzTjjP2P2OGc4utgCTDyluLGVqCOB0Q5u4Umbo5Oy8kFI2e
eogJuGBwzrdc5x/z0KzInPwgjuW5hmvZtZinLxZvQxd6ajN47zSExhtiHnwkN9tQ80R07BAD8Yxp
ONhoS3ePCfUlbgz27WrIM/RAROTXzfEZcs7b/v68rcpULNENAKOanK8zUVnVgfFLscWf/VlmgavG
1/96qC7d3x9OZ251riQoaJIefnXFYyU2zQSYtjTygTlN2tQX3oF3+/YMIjFfvz1BpyIZGEVUh6ZH
cb6MkCNfJeKResJ7X7UpETA6n8TuzdsOTdD/jG49GsHmTUPcjkYwyGnE+rFoaPBPKNJ7ARdmun5K
1goN8pykx6fftV7utyKBsqx9dgnOdulnHngcBY7QRXdwFp1Jr8lSGaUkvvHygnQksZ5OfPJiwvBD
X/bs+a1x1teqj69WgqKmeqpaJ5+rrymDU28WXQ6JiEu+CKvZVAFNYmiQ2PoV9F4FWPREMBwUzBQ+
jtqXXqL0vafoVAJ/R5U4MUAbVHYVUIQD2uRAlNsSLwpirv2QNn+AjcVeBKDjpFrp1XAusRH3O+Ty
qWL51B8oybwddBvLBRBo7+fmVxLglkIjx23BQOYbQ9m47WC5pAtQIUHykLzmAwn/Pnu+tPAtcFrI
7Pv3U/7T+vI3yXWZRAxRaA50ZpCaNf1MOIDQZUMLbQqHSegBwGA7eYRDLDux23GQh4biiHEmL65c
ul64P+1OVkB6FMu5pT6C0wDh6qYOA6gNLdmgXP8+QY20nrn7znngvPP87/KBa/h5dzP5GAKpNZg5
wXWKo4N+erCExV96vjSvbpRRpe2382bkz0EuShXKxhApRPAIgeR/N21fEdJQQr0GCknH0gHFMuaF
VStBFUCoL8/nVKYHq8j/St2Z//nOaEGyP08aF01moft1j28iN0lXGb/2H1HvEiwgP3fGdzuUfUnp
aPAtP7T8bfQDOm9UQbiIouQARamq3VE9roRjW8niwkfboJGLZzA3jWAUAV/uQrreWWMiytBdPJts
Venx5w1EGzQm7fZYWUom55HiJzUBetuLvRq/Kiojqr1atvHevboTM4+k4Nus7jh9LD4ze6NXnJGP
MYbbgPrC4/AOssSW9+qjEiDIaVDd7bSK/3dbpS657Ecc2S4qkDcMtoS8SmxqwraQ8K9XlHo7s9+7
yumE5JFd5lfiUmTtWT+1rskKFM3e+eJUNmfESYXLzb5xqP2/tD54Z4zMtdhq4O4TCDNJYsjXL0Hl
UxEee8x22/Jazcb6CSChCuRqp7ypJ/e14xKr31igF5fc5STKDyqwoGvIp/CBjmkHQIXBG2/eQsIh
zASBaYiPZrrOhm/FpHfAoY46Oc//7GFWg+1IVobSUvZbBaUuv0T6VCF17+WXC+mtcxVNYT1x99xN
XvDiiRqJ622SDZZaOhzVGAcudFHMnD5/gxdRTm0jXLbtLQnyAaGEicbMMbbPsC5lwthBbsroCiO9
VjazMQkf4utpZcRNI7Dx+e6r0NkWCYyDa/rOml+Jsax7eHD/9U6hY0+bHjuJ6EukcactxWzh/Fml
gG6YsB6lnT+kLTLy+oJmSJWkTotoYox7POSMZMjMII3hBJAe9dnyjmFsQKv06U0REwm3fBXxVpo8
ujE2w8YsF+PwiDttakfPAOCJqG0kGnn1y7JAg1D6e9lLeukRfkwghZPi4HxISnBlTSgx+Brgx8Bb
PnHPIuRlEZeUxNpeh+vznKySxFUDDQg2wPHw1rh8qldNrVcuc1qILl25D/GpJJ68n/u/y6C2c5L8
dc3OizJxY0pmq2VO136dJN7NKrzB4r0tasuZd/nb4TWlGk8EqYJJ05WwANC8YfDq/0vaPQXR4Joi
agCSL+5lXC8+xQqY8BrbmD+ln9j1etnWFGVN7InKLdEj5PYbZhyxjUqEARqrMPS4vBo9fxbJhKL9
nkH3QpHvJx3UzhaWZw4nTbAuxA8hoNQLEWR3FLP2qcFSHQllsh8HvFxXgtKqFO3roMZAaErvDjNr
nf4E+tPKkTuo7InaTtzrlEfGa2HPEVzb0WR8ddUSUJBfRkkfLFOL2f3/uW06fWcqp2iJPIqQzhnA
X+7GXuvXhsaVF5BJAIXNxAuYU0Ix/JcHatrLMHqDNIgdHurKr6jSs22XmAAJhNd8oYcchQ8pyQ8h
hAYuMYaidgAhhHcM2DBU0M7hBrFy8+FfZUfRQVWBFrZbLfLLjL4Y/Za6Cu//4PSxcfnoJwWhjPY+
zryDD/26W3O5rNNntmG7Xtpo5bm4UyNCStqEhddfadFzPuzCej/gig5VwZ80fVqVw0vKaGR/d78u
yB/o7067J+Cn7ksDG+GjiFPfQSNhQgEBGmJixbt/K42/CqkRMckWDtj7G8qH3MKuS6j+inLGrszk
+KL+fFrL5/D+cTuyQjpwWm9LBSmlRKTc9S5bDAaYH4VpsZpXy2hZ7B/Lsb5ZGHOraK4K+ERW+qsB
WJZPCom/KArPwNl/ozTcqE1E2FGQippRa7BzOKiuN40Q41oAXkekf78TIB5nfWNuaw8aNBq/7FQ/
YoGLtvZ5SbnBO5mJZJaGs0emc0dV1lrkUfu+aV25Nf9lvO4GBBsqa/dSuNdPJG4B7lwLWYt/kclq
iEnwSPbsDRjuyT2GhjHBAw24w2tLCIvFFs2g44U4TJfDtI3ARK4rJwQ/P7I+pZna6X65fdjj2kyd
7wiHP+G4aTY0c1eYEcGv6nx/4hJaa1/j2rkq0GjGj+I4dqgEMSbELBHQiR0AKNWvkjP+tuGJ9cZx
0KNnPM10KsY19TRJdjFtAkjOO5ia+HDY5HW4tIgCQ5o6KGN0gAUM4UCg9y/nhquh18St59eKlp7x
fOd5dElZEyGnCF70Zrv0x/RCyjEiuqV4VCp8gYXuf+grlDwI1j14+wVRG6AFLiqkuT1UfW/CH2D1
rInkIiqpkEZxTCOBKPICEbaYA1AJ1Uwq/5j3EQ5Zx6DbQ3oV8TRDQVgS5nZlbTqUa3dsbEbWuSWz
wp+a+Nd3knDjgwW14N+K+EDihYe7C7n7i7iWkN+vYXXfni2BcvIM7yZVO5SzJqOciFx3O5XDZ1Qp
8O3khOBdObUKVhl196qEuCDw6yX/EHTwYn28+cfHqCaGbiNLO3lB8e2bXhEGruKFq11ohzSkNWYj
IMfPyiiQKzIAV722MAgO2U5r/MvtT4YtFXdft9VDqrrKFwmW8NA5knz5A2vFZPJqnNa80aSXapX+
1KE75Tco2inOq7yiDPhIsnD9gLCmFGqFMSVXnweomtc2FaFS4y4wfXWzrR7VnXrclg0BO5hroWJn
FQh92toTUfhNyjfMMxqDlr6cjukuGOeE9zoBmcrUYeKegnO9XTkuXPxEyPVIQvZq3U7dT2yAnu3Z
ZJyfYT1v3lB8b69GKJ6iIfQNWnN3ZElS7J1XExZGu5k/aoAcEAyF9Wkl+u904STMZGrKup/hEVfm
8nxxAmZTdaRZvsf/CxtL495NXnMVNEC1xdfzYZKCPicB27lnpmVjm8OMmv1fCuHS77ED2S89xtw/
cEfbIq8LJ8dXgn95iZSJdvMmrxI9JKePVRS0/12tAgzX54LbCPHCcKXItdcsCUDkmxEIxhDTct3p
VM2skgKKVuT70Y2dh/vV6k1evxhBsPS8SLzyCFzk9sls48pJdtxl5n/9gGD7ZdvV2UlAEwa8bdZr
GcLpzjc93OziFGA02OOJPU8pg1t/rLDpFwBMuyjrenVVIteWkcbGXy/80klQGBO6oHwiN7ebYkfm
/SUTSeEiS7LgGI8Pw4l9yFvKAM9hOcv7EK8p4nrL8o2atgm5RoxxviWacnBSnGfLFS0YlV+aRKLc
48pnB6IWog3iNtQl0JJoGe7ZnBOnr6aidOj+1fPivXVC0EaKyyW4+sT0GcINuts7kH6H0hV33m5m
aYETEM5A21+aoHsGClhEURo6MDYGtGBOhDQfQPNonvB+13bmF479F1HIG+4eZjh+7ZqSE4zdyaCY
uFr5pcC6DiKg1fs+kYlNfEzIuYcxrSRVMSDiLsRoxpRe9tSyc43YHlcqB6xeMLoJ/p+fBz5GNsvR
X4TYwecSRV3ex6b2uzXNHAWaXnLwSaUmIkk9aIhZgab2ux1LxlfpIJMLI2YmMoirzyOXdruRfUL/
C+aj8QGKvsPhsgajaqjGoJbPFgIbQhG/v/60iDDXzka1uSUIc9nsOVKqkuu6jCGeFSfF8uVRC2QA
k+Qdl6HST1UZvYuV1p9jWhXbEyso/FSuziCR4U+m42eccP5C9uOY1+rpqCLtN0DuzpLOCrVRFN9j
fIE0FFvo4g3A/Ie2/fw+5knkhAVmFhBNpNRmltC/VSd2etDLHRozvPLlio7mywY96Sfj2KZHAW6A
y9h1rXjlHeKM7My7CSCSbwSGX37VnovUlaA2Npc4rYssF+UCsqtgEe4LVIznXbG42L+S+6KFUGh6
dntTh1egISbetcbLlOkdmVQyBa59C/DoLCSKCswB78d6kj0p0MrGRrTPnmZyKWvcnGTGjeBWu6/D
sohcb3CB1I5B5cX1IoQz+XpvN9WWPoezgo4DuHKsIjpGrjP6ulFB7ozFs8N8PZPyyRXj53r5bcyX
6X4TnMpCRHQ2cMXxlT4w5jKpDVxS28+/gCZMM00nRRGYJMUV952fIWXEm3XLtMefQ9/fK/Rt0AnA
Ek2y0MOSOK/F2CZgJ3uJtvqTvYHTbfpnEpODLoNP3ofpr9BKQS8JXvtCWte4LhHLj1QJOAgxjFXN
a9vr5t5dKJcmmbpcs+AEHm2PwavRHM/e+lZMdvDmWl4PP9MhMXrcUIC7hI8HsEQq/c+NK9wCJ77x
85zL+YhTsfJBMMz0rLo7IGL1xCFhvA9RxKQ5+c25iCCVlyb2wk6rdohB2Qc0lpMF7kzxwFDlrkBK
Ob3Vky6Kyf8RADA+Ng2e8aejU20jWuQDQcz4SfobHYPSv+xulAHQaM+D/sqcqKX7ZnPT0AMYQ1OW
tOAzFpVZkln4kzc5nQ5MImt51SjxHLweJmV0DbUkGlhEopPPV8Q1K1MzdxblL3bQ7vd2lbxRUPYN
CTImoe4LkVQSHbgj2OSRvBLpiyS67WqZWWvsTuFdfY1dZt8ZEzcsaahqoGRXWmxBU3BrcA7KyKyp
6zPUe0xVQlVkuzMagUQ767CVE/rodQ6y/HCMIBK3SHxZHR0GsmR0maZMIERWRZ0ysVWn0k3dbs8x
ZCatGhzoosuxEA3rGwQ9Eqb1pvOOAIBZ7aBoxC6LQzw88HZgU7JvCRVIQOKGvE/k2tGJlgxRZVXb
Hz5M99LPz5kxzJ9v/KGW3J4Mdyl68PFH7lUglPuHsZYWwpTnaNYTIMgA9jK3jiTH8MDtxn7dEAod
2TVCplA0hr7yaYEmPNkRj2vGIsKdteaVdBncu9Jh9IENDpPj/Pm4KbVEBed36hz0IiSpzl9Wddsl
Czd8vt4K4YOzeK5odIB86omr6qgER8TWWtA21JVYLPi5Ng6NDcsFxoGci7qgR3BQYn+EBe6ASlAy
od1Mh3kF7jG+l9o1s3fxmoDkQn93m/p8t108/kOJjvnbO/9yysTLz3PSnalQwLvaoBzJfaTiKFol
qm7CR3LRr9ZC4ZY1OBxDafUndVys7IgoTcQ3rwCsRdrV3zoFuk3vNa5euNqXrOertbvOaRxHDIRs
TRGjkesTZOwFvJJg1f7HOSafuLPTPcJjfFr52+6foepPeM16zirzNHHPTvEXHSTE3IH30XwB3yMi
CnBRVeVptWTLygMvnGXyrqI4Xcm+XZ/+gY5gzy8ydlL3aFq57urtD+EDxMNWY7dFze1RlRccGc1h
s/zAOeO4DzI4igezGcxDRclES1wCg6pevPq2TzK+yAUPaMF8J5kPgmSe7KfXsdmhAn+Q35mXOfjQ
xF87laytab+KmGsoWRZjyS8gOyYzLOvKVvQhsFg8Fi0h1RJaTMji3TaThx/51c06X8b7nwdlaann
6CPx2tf2CVVsWD23ABeaaKWeGAk4FebD83B2oL/1jv3/OnUimDgRA1DnWrKWLUcnUM52uqXdZUQA
d4M9DKCxTmL1dRbRuJEAG4T81kpCFgRvIP2wNTC1bNVqGpOwIybQZCgUHvs5ixZZHO/y8CYrBwu8
5IMAS0Xeu0BA/K+iOcnAoa3Vx3jnV4yIybF/lqpl1bqlHjnO0t7QQyBMGVdYLdD4aSBdBd3LaA7P
ltMZi94zZ96WAj0gn4czBhR4l6pxiWGfwm34PQzUcgnNVeHRb3C9yD9BLUvH9/7mBQo5U/3FfXbf
oQDHZigXq6JxY5n0QjMxYUGQlM1V/cYD0uYuRK+VrLfqC02BAfjyKW9x3kgN2HYg/aV+NvyaSo0D
tKcyWPwh5So5Isr6GTWyZvc20zlyHAzwlyLUBpZqOXMxVgry/HrC85JDLEG1XgqnbMKbWyajMV5/
1lnJJO0rab+I2kmaXZNVGpSGkoCHWUyN/1CJXsT+NGVi9w8FDgtF3IFaMRDfh4AgdAfdrhc3fk5A
WcykiMX5jsTiyITJuERn7r0vPKvDEkwAEzgBLU35YjO/2jtEs51JooRa3Cb3TM0X6ve0GacClclT
z89dGjGEi2dtz7HhZpHNiGOkI49Pm+62C6DLa9vI1rvzQYtV41s7K50Sbx3Im+xncXrMwdAAXN9y
zfftmgAtzIoi4gkGYHnza05IkcDhGNZJ53W+fJ/SjnGz9JWAEBXbfi4AARM0DMEOUDfMTUCb1u0n
Owg1yfSAJTbodhRT1OsbUTPeWbivoXydvfYcpgvPN3tN6x8VxfxWjlZ0zBiYeSe+1ZAkOTkiNZ8C
LO3rJm2PKJRdTkOT2YG8+qB+y80xqJPncFWr2eGOkLejyoJGxf5T/ThIgQICdj2gVngmC20RfPwx
i9ytkz2S5AZfzDUzatU+2Od5zFeQFDau/8/Q0DY1yFfPtxoUOtoDZjGRPQgEf18TxoRpVo2lMw7M
vli4iJvdlBR6DiIgzTcMDYRb1FMi0WtJqXWs/0NRlwNK2zO2pDaSZtHmC743vn6o+PQ3wwPyHwZ1
sUDLtzKQZn5/kk7ERf3/Jhje2g5WAItQ0t2nM9F5kf7rvg6xQfdiM7TdNqoKUDqfiB1uUCWUou5Z
Z9KiGE+H94v8faDg7KZvtFg4EuW7Y+V1k8PX4vQ1m6Zp+WUcAjjxkxkiQ0fAAheEmuvxFd7AVfwy
FcwSPB9m6olO8xZY03UZGWhNknvOW+yYKfT9lM2sN/eqwnP+3qu4hadpGM4O5q3dk1Kn95uBPDyH
fivyQi+LlzaUjOpMDJC3apjetGscAKdso3teLAa39uEsWDBaug/4WbmZiIV4KdgsS6YlaUWX2r4s
9nKSher7mL5tmilp+iq2now8A0cY8ZGx8zoaRcYiyJpsBjmWckZkQIFMUCgtaN8iDdaytE1U88d2
2hQJiJjJdn/N7C+HMMTqqN5NxtI0TCbXNz6SHC9VZNuuiaiNd8I+KiwPByQlUpTMjDTvAglg7lk3
ARvsTYqJxFYROimG4r+PMpYPG0BYZR1PPan6bEGa08Dp39BB9KGsDrzELG00FJ+XFSu3xcb+g4TG
1vE1VB8ysSFkkZNmtHaMxU9+2jdv1HumkzoTpnu0q4JrYb9lKQL9KeGPr1H+5tgOrZ/L5sQzeOkW
w891pUg7x86eagfEOnXxKiFJU/pghc5Rb7vBhce8ILVkUC1Vf6LoCYYhmhlJ1jmiShj7ouzxicZr
pT5hqP0grMR7FHlDkuZqZFiOxHAR1pSJCh284r1Xoe3bNLrSjqa9+4E9RzYkStHm6Fmod3Ne+uhl
6asOqvTpGy/e409HjZ3v2s9oBy3N/j+fyygqJilKTMl6JuZx8PtLRfI2PdvnuSJS+HXlFrm2Y3P9
KIPjyZzvLvcUpZ0jhlol+7eZxTe8WXEXyL0+Us+NxG6KUmvPNSMotqufhlpbDu/s3pIC9qO6+gXq
p9p1sYUJOLFKaKUymdLZJ88peJ3N469lfU9rzlR1x6Gr5Mk7V+dk7U6ABUa08YDRc0XXgoDzsO3b
D+JQyqAVQoZ/wkgCweeIGIiHPW8FwFxjpGv62CSmZEiyUxvk9FfN6JU4P61TlQMZWcADe6YvtLve
y63imrwFXNyHb99xkMIKJ8pvloiOkFvKmMz1cY90dMMnZDSjhhNNTwHw1jbtdajXVe3l+ALDUf+R
QONw8QdNusDJwsNy5klfMougei9uS+zRmTPPZxmRS2WA5wd9piRAw9JlkFdDrhY7+cu7siNDZhfP
sR0CzDN1cLA0ZVoTU/A70FueiW54A2A5B1uzLGFsmS78p+AzHCjyy1maTnPRnbRw6OGkSeS1zbe9
KMJk3H71vgku2SeCLzq2wv4uJhHGSr/xQvYtzuDGxYbuu8HTkP6P7Xu516GsF0G1qiZc+VgolZ9z
zn35bY0ggMyePhhQCzbgycGFO616PD05lFP+3a+K0S4F9ZHCDuqTrsp62rRfy2tq8ms+i5vefIU0
GEnqzpQbP62qKjxn24pzxEcp0XpPzCPSg90EQ/UeE/BD9eXW1yb3wWQVcMcqmOm7JIljdq0YSKdB
k2T0dOsp+X+cgPNgC6G5H3TGEqR+j9FcIKPnTur6nL4XrJ3iWGngyb73GgbXjyipJJzQTZQZhGgA
iS49kN25OK1iu29mMTwhCRMMzbSrcjs5Fd8WTaM2eW9rZ/H0ySiPSZsA7D8slA6HxN56sH6deB95
5dM4yskgGZLjx1tddmXn6ipWHSqzp17W2SZmuCYzUvWAHVvJE2FTb8C64XZECkFKBUpqksPFd+mc
ce3qu59l6s4nVjqJuOUBecPtX3amCsPyBh2umj+x9knnZ1bMS2tJLSNWX6iu/29KcHps9haw8Tfv
7TWMY/g17EilOAMXBhPC56k0YobaL5pi7uF4nUXEUUr2YlfwzguXWBhFtntzOUG4aqeb7Dw6kPkv
rFs9gavdLbu4/JgITpulPz7zA66aENwxy78k35zM+V83vgEe2QvnSwBgrqc4Kk2b6JG/M6mH0hfc
P2Mb5/h7nBJEhV5kXRLdIapCaMJdEf7Q6CkN4QQ6vni5opSePNp0umDhBV4bzVD4sHTZArIT5kpZ
i1WeLcHGWMKk7qWR+AIcpXwalFBbNIdHRUoqwL8nuwZ/R97KPeE2+ylQep5zV8j1KTf+g1ppJXLk
Ui6MDIOln/BfzVqlcpHAOCYKkXbtN2hV06h+kaNFMKFDBxw4F4dTRhCPdKTi97jXTXb/3UxCQ3Af
QS8YRN+2kUd/5iICTN4KGR9M9dbiPZt7hsqcc/8GetKQKh9GTprcyRgQO2vcMBkRR+Lou2s4t7s4
uK2JDvH8dXJjO+a3l8KdiB/MkwWfDuewqoqm+9h4FjJWGzWqKlEfJ1QG531VhAEBPpBJJKpj9iRF
4CsreWp9LsxG4mgzyRWXsnX3Ys57TkbMMUNhVsOtz3UHTgPYcVwuwoE3DlZJ4rbQdYYLeyUDF3eM
28F2m6513G018uosoveuVGHvZ91/oxvlu1mhacamzApLGkKHs5GyPbdlqFm4wLIyhVat9X1QU5Em
nMncV9hGpv4YCq82G4/1W1LGQMkYjhSb1Ny8g9n6XnuiDjzaw6XAm+M2r6sKSjYt3zI/hnt0ragG
p0dbREfwUEY3lyTcObqPAlIt/hy3FEgoEbVE56yVGiwtgBtCqueJ9/CBBMEki2iamSE8Pb67rtzU
IqMF0ezKjFZ6coqNh9C+kvL+qUGnUidT+x4dCNqbT3jPBl2/qRYVp6zqZKl7CIQRSNhu+qHgXQBT
KTpGrkCm6pA9NfUR8SfJJu0izDwXdgx4tsFp8+B3+zK3ZgO4uHEtHSBB+QMb9QQePKu+jQr8hMgw
Rx8dk7tPCes75rdcIK9bq8hsmvZQN0XYLcr+2rqHsMNuvAxxxC7MnXG77mW3VUCj/k4rjX6z9HTk
VD0KLDn0creAgOtPJbKhZs4OYL/DSFTyexH8SZwTiZPBDgvuxYKPT6bAXmCJVVKYGIg6ufDPTIqs
E0RtL+HKdhviZ7/edSoPDKEAH71yslzNFmqKXRt11CN1fwczR24S2p+HN7q9qRgB0s4LzTEoEGf8
8kdoNf0HCGFOrwe88lfYWvleuI7JCUP5ESGC5V8Tl0vYStwhNaFo6LpPqEc3pEOeHRdWik2rvYNA
IF3OvJ2Soqf1UC0DtOTiKUK5ZwW2cd024+kuKKbbhOXXn7HD874vHO/hSC0vL6W99VHiZf3EloQg
msZrx1GJCC8HjGI6Wna174AYQRElMxG2D0D0k3vpUSspRn5AOWgGWIm3WQEgIsU6QJ1wT7YkcfyA
GDq7pPvnhILB3AVX2g7xC1JNigQfv+uOV1oLtDIq+sQyENzkBFmPN+X1eGy+HUad7beiHQykhhBK
RCnLoZ0GnUea4bRd4VURgcAWzHiczll0Zrs/8R6pOpWa7HKKfkXQwAwkUCFYNngFvIrbBHmD7kae
3rSYtjsscQx1aB0qBDl4nThdWNOULKE+zvLRCnALAKFr35yUczsz2XdgiSaG/dPE9HWANz/MDGwN
+OyuHmT9UaM0eIhUlIyg3ODcv6+3VXnykOpdu3bViG9GXcOM8ZVSVXgK1GgM8IFmq5zFRH4rxMJ5
F5c5ac5Tk8aU49aBu6NJR1eKRxz4u1MkAGgWDd6T3xaSBQQgY3/soxKjQcFiKV7Daph2W0RsbP7g
JmQSBF3j8VB+gzIuR98uqayYy39qqohEClBo1dCQcYqQ7Bo3DWJbRGtFBIcBWx6JpwI2/iZrsfWW
wyQuI4D1bAGkG6+4TZIEzCBGZzxqZlIJ9kaEx9dSN7u0bnRUs6FagIjBzOSGkP6X3aiC3oZeUd5V
84qsMiYmqyniP6e/7CxNgyESxhfAWNaTzDBnStWFPxYwMlPcq8Hqxx/O7ki3rrOxfZ+0CJuI7f/W
TROM3f2dMzm1lyzIwODFIwBwDHSTAm4CkqFr+MMZ7/C06PPQbqtzjCwf61xNW9YmD7hRfpy4wY4w
w/CuUORER21khIhBT9PlVtDyFKu34ibVRQHBvcQlrHag5RDInuoBNkSaC7EkypKI1OSiqW46Nzb1
Ddw89X6rE7q/ArdXFrMret+Az+py8FvLR8QmHKJrCuqH0k7Za0gcHmCsVDLXOO7CeHlZ3wWJm7Ij
RbWUQ44Zyl2TFE7kGnoDAKPTC4I1rYsJoz3jCwnVLj3lYQ4JNTcAXSzpjO9uCKfhRIvp+5OO2Aia
r6SPEa//Q5FUuKVzbGmOGEv+gHZHBP7+WK5FQacgj9FQ6tUTIpvZ0xJ+OnNcpZgou834TiwWyjxf
9HP5BiKRvD2Dg4F4SrPGy+N0yACfXYF8Aun0WAVQ+NY0+Klp55Fb8y/VPRwWaav0y414bAfc9Z6M
ccTYAlW+oSz68QXaUIUgt+TwIy943uCihYnDUOwgNVyJhaKrd0Ao5Ie5tZp47ZRJqHj+zBdCxvyO
L0Ve026lQfUCDoYyOsjtY36K1Kp83IowWI0+s1i+aAVkWJoimLbGwlaUtah6UKAl81hk7yMiQFB5
lJpJd+/ccQt+FbkVOo7FziJ+9lnqi8+1O4+cni6XQrmqO3xPO8YA/rQ6oAH+ydZ44jht0p8Coa9H
MeLNV03uQzN92iBURSoX8jUmRHhLU9WMCXG650VQNKgVe9e8vz4NI1bWp7rA6CgXGuNtuseb5NUo
bNTIGY239T1MoVw8xk1Yr+3blSKJNbsvDPWZVesKKpPo47sdqyv/aUWRi0FLzfzSvavtTxRD6Qep
Yp5UniEeK0tTAgNBkWFoJQmxvXFR92V+T+X+oEe2v5BJFAN2cYiUWTfsC26Ievd153YRcyO2If+V
KFXYGuDMOVKYNb0mY3YdFqiOJGwZt7ngszUhmJQBxAjzF9ieFL9NqdlLZ7cJ/s2J9tl+oheSqojc
m0dk80GX92pO72pzFdLD0/RGZ6g/mAURmxU0jgQibtxSpq1w8tV0ThxJEkzX6ctQPm+443/uwGDd
MwnezJNzEF4CR/fVqwBKOq07vBfTAqF6282bh5tCJomcgfBM8g3fKzYOemEvI//Z6nGe1lg/URGV
NY7djpzfeOWChMOx6ooyfaauJQxAV0xDvOL8HabZ16AgKpz6KlXBt47pVFq5vDD/bXhoK/cJyGOG
zj8NMImY7F/+DdVH/VLIfuHrggnop//UJ/274wBpwoBYmyFpWXZ17L6AoXJh+rXnHFvSXGFDskui
kwBhoeqKdo+m9+pDaXvdG8Ckj1YHhejGL3RqMFDj+kXm4Tgmgjw+TPQ3mN6S2luj5nLm69ibvc6p
lC8KkpmP+WxNMQi7T3sLj1rizPLN/VJVeGRSRQrSGBJuBgTd6xFzOBMDdC5sQ1xTzne9zKMvrrvC
U1416z1U23C4ZoeFEvHP/a72JTa5Uu/SoHxzuQw7aZ60SUECblRKo/qiSemMmigXF5/cVwJ5/d1p
fYyhYwBWnUwpxB6WXyD9W0K1I/OojEcQ5SxvSsod4nYCM9DRKpjAZft9iqjfwITS3f3NojK3zYLp
L9eo0PIryBe8z3yU/kGdvyULLcbwPHA2rEDJs/ZbxT3N5/wBg29sZddbrxxdb4ezuL4hBcVipgTe
hG5SGjiNK9x04BYVShgrZYmDA9YT22WYmsbopOtekCGgQDJtKpaGBBmHOItmjYjSNz7x5ibUIq2U
OvgfljFLBACde/Bx4REw7v6JhICsvgUn8ZtivSKZxe+G07k+M+FxrI+pYL6aElvfmv44EKGo6VvU
+gwth04vrUR32Pz1ss0df+wqAD85UdxDjPZzyRSO7nUWdfiRNxu4wpIE+XzXuOMD2xktvDJ5b6ho
u6QGZsF4FDmx/wsN/UYUbgsdRYt96oEAtvtSvb3jf6+48+Z5BhNvS5UoZot1luQDMn1hKLvOe0Nr
7hDj3vQhwvycAWJgEU7tjH+5rxSppNTTyUzUPnUjlf7YnHbEijpBpgqS4fd9st5uDGWY/KvDv/8n
TH0KFCcyCZojssE1uKbUcLtfGvRVd5Gcx0vuQOBey487EX0Ip1Nc33wX89xiP4gfY3IMzDGex2q4
i8zWbg4sZ1dGEmZv8L1DZBTqQcdy1VrGl0KQjvGgHDfKhM5aocV4Vc16Hgw2EUyfNnRY//hKPH1Y
Q0ftDX/wc0jRM/OS/Kh7SRiqNoJhyMBzxrnHNjG7u5HAhq9rtlU7hDkB/q2SLq/NR+baS1bhv/Zk
In5MgLis09DiDqv6pB0DOd5xl0HuztswhLE18ujvqj/W99V8uSM8VOfcbyBaAh1lHf0Txv8x6XXQ
OfqDPNpZ0zHKpMNkG0MDQHP+77ilAUUVIVESmnLCm0BIgrOms+B44lTGR9K4uwJ5YHNh+9W//Fvz
QwgJvYkpr0MfHHuTl2aYLd78IHhJzm/8o0H9pNvwn8yI/e0w7ez0wK8FIBbpT30ZmgdfkQPjmbzi
1kk3G8EeGxyE1pTFf88IVkPviUXRic3ORk3awqxVGvfrpSHkzL/4XyrYOAs5g9F0dqX5HRG2kNeo
esi02L0yUM2va8Q2vfCta49lhafhp930oolIqcxP48puNCHH+YGAxTkLyNc2pqSrf0da8KlOpbEi
EaejBg2lMWBv6QEy8io9JWpxjon1/bNIdasbZn4cEj2Cvu1dAIHPYDIynbxY9ItBljCiE2CSV6Az
OSYXAn8cYTjRFTQ+WnaT5eLEESQJe2LBX0WoWQWy31uypFHMD2TniXVFx23878U/OOtQvYNeR8wx
gJiApI7F4BJYQy7EucOKU5sOq9PG94ARd7oWH+HYLpDujbXnU7rkBhSz+WeF1RNEHwY84xC1mvqF
qGikmDTGqv6Op2wkWvwZkR55HWC7QomtxCMrYUM/SSrjnKZey04hiZ9StowfmYysMRBW81b6+iXN
CVEGije9AurUG5KLvzhp4bRTxNsDL+Q50L7iF0ye3nJc89tIj69YyVlPUc/m3jl+GVBBsv/A2khm
2o3s4nnVQyU1F/8PWP63M6W4We4Nq1Eygu2jmJu0Eh+SHXPOWMKTqI6UPZMOuARLORoxoeOw3vFS
BBppM8etos/C1v03BZZx23bv07GgNarI/NViYYt3C+La9WGeXboOFrh6E8PL7/MNF58v7adHdwyw
ZgGBehzEM7ByrLP+Argg73KW4RlfiVGC8/+0+wpaCuc1FRn3jn+/Veg3oUIsUVcu7J4L9fN+h9tY
DCpOFnN0cc6uj8WLgcyU1f1UluQjG9tqZfnB8Iiiqh7cDWJ6/xKtJtoNKCu3HvVEFTjb3zMDQ/6h
+UCSiaso+/u93DTcP499dVoshAC72PtR9BYYURCoD6/EcwBfxdQnaGW4TwV6KPws68st8uDQjgVz
N2OqY170qvAyUR4W8bcicB+GIlUka1+ynBOyUl9vFROQ0QMOsVays855qJSPR8VwWwZYJKlaCAjA
az8whOqyuBcoFr+HGgEIYxPIzHmG/DPJI6kDFt4JJXemYzDAOUKxfSf9hlnWLyoar6QEr+e9QIlq
DTEGdZp8qIJMc5mifPHumNlLPyitSFfF7PtcE3o+GMUHEflZpLb0KsQ2bhCTnSV5oM6Us49Dwpb8
Vr6fw/rRi1TnXkIDj8kcCdwk9R5Vga3dTt98aeY/TvZqzOEexYR3lBKdFirNPRIKeM9hHQvqT4bM
5MSQ2gAZIYMZ4nnoAALkdMiFnMJyKNy0DEIghYZBsl8hdzCv1nGkkDevi0q+qECh1fi+1PK1Nsfz
NAXM/G6uaS1Er9CPNczPdOET9/MnABMjJ55h+Gj9RFaLDfjP9uPxRo3OeKRc7Jn3P47/aYk9Ax6P
jdDoeBPuNc2SmPtUB2eM3vSZ/iIdtDSYELlLI+f/w5VMv2lSXJFOCYtKaNsbOj4LwtW2YOU+87GR
PngIgXL5msRrbty3QynYovQIsWL5OnYyOe4TE4Yx4irr7+YjKsgVbUPd2IuZ+O00Wt3Rsr8zKz82
+IUgaLo1iucW4vuBRjD5utIdAWYstZCmRIiT7I9gl69VsnwHWK16gTPgi6wy99QgT1Phx7IxSdLN
nURQNDMGdrlVDSbrVY8G1vHLtzckeH6BoLBYfaAmSQLayxIMA4lcg4VYyx6mvEy1nos8a7yY+1j1
Q6p5mmVRzOlFRYLPnC0Ddjd3oGUtcNH98oHDwjrpgFWzGFicboV9wo9wEUrBYntDZuLygFB+s9JQ
VPckwXkUvkCrkc13vLoi3If31BK6zFvxsFi1uJ6UMuhH+qT6fiL3Oxc7GGeZmJOLyqtGP89umZTy
N3+ciTBR6tYwIJiOh0TzpTVjeQFlkg1g64tiJ6KaYFdgbTpYn2v3TdYxyq9Nh4ZKL8GvVnhHtOGz
YyU9HwtbVzdQJRkLGthvJpERSx9uVf7VM4zUbw0CNwIBjc5t4PLIpEePswXRqiz7GYn2sQovH04q
Rncmi9bG/MqdIjxHuu3AG/TUUnB/Cy2wNicatWu2vq+eWsiPgqgAI/cJF+PHnaCQwPhz7OVt+UaS
RY6yX1qOctIBY3VFOOY3yUeP8aVORliFp6ZzHZcQqV9XpHgH09MBiiSkQV/fgZUi2ZDURpcFm6h2
fIn3NzefTKO35wHFpQfrMpSRLipanIxKEm+1LaUobwVcq6T9N4S/NipSDpnM60g8FtHyD8wZHLz8
KTuGqBXb/bbSZ8FG4pYgqNp2BysW7TTOaEw6Aq7M7BZLh+C8jyPnybauYY63djDTjA4UCXhhZep2
5HQtDI62gZPzkFmZ9ca289oXeSeR/LIjZuUDehAiNVGRGUBQoCHM6vFBJWsUEUOe4gSb2mfXO/OZ
flPLPJdxEJAXkCW4hd3kP/wcyJumY/Xu1Pxzwv2m/DM/D8FrsM9YJXRyElUPc2Ls+AHhuM1Yld+m
IDXOWIjtZ07rdrSzzqkxG+ASS85WZTLoMvUk1FJ3zAdN+7kszUbn0RaxaGzUxbnnajaihg88t5TZ
+ao6OZvS1QFWhxcs/iNo/cyarQNL+4cIG9Bw3123K++FA/FcRhKvNE98WvforAags0qqkEIgsltK
kaQ//VjK9PJEJ7WtJsdWqA8Xy12RtsFjEVkpv1rUImfPbcy5l3wNEkCHnlSWw7LUE6jj1ZtwLZX6
iRwpD8XlkQEJS97tvSNbojVKUbbxXWKljY2Kw1/83K0dw19gSdvuyC8+O4NIDk4oE2aOEZlU0R0h
aJ+rq7QSo7WmFjFIKe0D1X3Yo/GBAjviUdvQOtAwOKzBjrtRxW+UAhvL6qajduGksdgI/tTOGH0W
lnjonZj5MPfXlsD4dmIG2oXpavI3L2jzFFrG2V+keEpSzDOZrcsrfj8a68sWfH7OPJhxvM1kjxgu
B2YXpC+irCf56T1+/7VwonDjI8iZG1TImeSMHoVqpqFldJQjVxaYZjaWAXgGQdHRrz2zGTV69utg
8o8qDWd1UOmOfLHgVkaeo8EMyKOn4piHLagISe2g/9zxODj/kDnMPKDfq28YAb/B6BJUKSSo0QEe
eaDLIlwJ5UvouDhyQWvlJI7LIdamqwQWNVRHY+bD7ZrQkA60KPm4NIS/oHHywgBeUMAZ3MyWrs2I
CnjUTIfXM8IJnk6e9pS0qeiP1ftZIRfR2Ovp92hVK9ekvw/pePzd+FcOPtjHbbspmEExUiI/ztxQ
mWp+r76DrpD6PGli723Hwpq946SxcGA36VMDtaKb/FZrfaWxByZHrBpqJZlaOfb2nB1dvXXc1f2i
8N7+gH5IMQqvKTTgEQzdqdZSCtGsSwWfXeKnchPYpu1iRJyhGYjjm3nmXaGb9Ss7z1vNe3LX1nDK
g67GEcdQlOzrjTUD0xkrOo1Uw1P6OeYM4UdUCWqzQ9DApLm7+1livGmcOIDAkKdgrcyHDRumyW43
GJs/azrd8NBPBMivdVCQ+lN69Oi6wR0KgDYqg2gQQJBSmOn/S9vPSVCQbXJ3+c34wErgd/sSLVeQ
p+F6Cxz+LhuM3FQYisYeO00MFccRuRC2dOtyvRkaNC9itVd3LLF8tMhtJfotdfPUJIOan1fjApxL
xW5btXA4ADdycciJmCqTgzTtwPj/WUljD9z8qGzv3l+f0II7ftJzO6qDKntefQkp6j4aLX8uqhr9
qP9X9Pey3/ugoFw4yDbGCPRW1lVWXVciItj00XwVXJquR7FHjpNaoeI273x02XGUAp8stEc5g4th
qRjU9P/+UftvZJwqHMhnKu/HLV5BB6YjTD45YK/XKsMq0Y3Sra0swk6LJ3bJ5N0sdGZdhCWCFuL9
3qDYYAbrUefMM5dhv1NprIMZqiwarQJbSQUgX5KFrX0qIIlXcuc7VIJBLoK94hqvnWaJyQktihbh
EbMCroux+YT3uYR3BZhsB2P5dVPfBDmDNwclaM8s5abHVNYakNR+sFMhEi/qXSwMVtmUN3y0KPI5
zKD9dnFbYFvCQ3lI2uFLWV1yO1sxGTLqthEDIzib9X8BLqalWwf5NI6l1WB+IksKUaKzbxJc7lrN
1vATqqzHMRxemBccTKTKMVgb2xyyNfJ5aLY+uq2yE8qBSD1zihVpDh2rS/yDZb40W8Uq2HKeFq/7
8/oyDfIaJ703qPvcb3hjupWqjeWnE7uUelG9pQJlgsjqErWHXz+CENogZpP+44pmY6cfk4qmBWW/
+RU4jLgRhLaO2Po33d5NYaFdbSMZZdClbY8iTzw4gut7RChjek4+eelncs2X5rT5UpQhsLl9f4SR
QTFchMC7WY3qvMvSNfmq35UhvfOG8idg71NRImosdZ7t9WVKx5BARjOvBCSzeROhns2degdZOv80
i2ZEk74bdwK5M2rBqe/RNSIEdYEcXhYPGOjdxaW37jYLRSxgsZce9UUEy41Oht1fJ572zfkiKiRK
8c8Ji3yWhKYXCzGZpIC0s+UR8Eqt92nIsd0rsRhnlMJQWB2H9xxnaO9OUDNv1yINsTxKOUrY4fqV
l9kstH099a++0hWkVmfCeXSM6+8t8gIeHaRFiSB1TgjT/6fKRSKmocu7wIYjaFU7yaj5fsCU5f76
o3GKxZnxm62pgHV86TEUjN7Gf60/hGNUDy/hR+QzRU+OEPnLB5KCzFREc4OkrhpDKC/dIvBgQAue
8i+CY/9OA+SsXJ9/QgIXXcXFIIWTTJqwKxVUle3roEBURDkHWqBxy2ByzeKIDPbS535MJMgY3FZL
xY+1/CB4JykZbiUqaoixzj0akkui8gOxtTerP+QqnUUDi6jWUxAc0G7ayWA3mW7D2ddlLs8Bf5WM
OKMeZQLAXAWYncSjO/jgdmLfUaL8SgxU/bdH4FzK3hcApk1APAhamNqwUVQGZ95VZgRHkfpuEkUb
UbOi8VRlOPJyR9sbj6bKL4JFF3tIEnXsRP5qbJTHBFj6oVA0P6QGdePD05sngaf6m19XDmFoJsNY
8Vwvl1pXbKSeniUI49PfvY/gCucqW4yv4P2YG6Q/BvJdcesstjnz0e/3Z7I3Wzgr3vfT6FLOfh+o
BE5F/yOKO/mA+g4xyu8lWUjA19STgiXVMKH7Zk77SFs0CME1Dx9pd65bM+IBagRumAlIOkhFgq9/
IP6dGFDM8cdLFAQHBZlJmhxYrYtatpfWQ70hTp50Vjf5VX2zizhUs8GzJWNW8zUkbCk2utAdk2eL
NoicSCjyeE7f5jmcLRHcg+aEELY2YLEc26d9/qx/Ecx8Nv78VNuBpkpkFve5sgVxuQXP4M5i21Lm
YUHCLtKbxI96El3Mk2VFTvlWjbzSmWxIiqBynZZ9vawnOydpF2YZ9aUUjcmUfZF+UUrPIPE2Q+vu
DvSnN+W/DmD9nLJhCU3KsQ/CCEMtWkRK7Pmi3s/Z537GB7h4a3AhxzQbGstxNBF/JIZq+de53+yh
IUvBnVVjyNx8z9pVcwuNx8tUciPY384/9AVnpPcHCaoA78NLs1qH0jZaxANhslTN3rhYVCQQ/qox
k9FY6O4tC35peA8KxZ1MRSnUS92CO6HZRyFa5RJYV+nyf3E4oUcHxZRepC/vcizRmQJI57D3qyPw
5KfUDhDAGeGhEoWnjsqsPf7/lOxofLyC0av4YacSWT69o+GUybpzeDIjhUOCIi/GZcpV1z7OGbqa
40BXyY7RGK577PwO08f7Y5DGAAzGtbDnZxcfRsTz4SmCSPu+Vz/TcQ7Og56tUV4/jqMtstVC0w/h
QGwYLw5q0Jg7UydddglQZMoF18eQIYaP6yiyADZAkjfhua5j8X4JQBrAYg5B1k1BNcttmSD5h+xs
o9EURThXdC9Uc/yN3QMks+7t2P1UdwyXR8Ss8OJFpreWNLqL5GhhYxi9xkKjbcBK+cAqzYVR05ao
KY4IX73JEzP87vKaUCK8OaWyPOdNLfSZRe7svy1/Trsmwnl/k684qSrw4WiVXtEdgYgkT+iswztz
txE7W44lmUJ9rUdl5w99holY0F8RTGHiEQRYDFzp/1vDeL/Al/xSRVXKdu0Y2YghhEb/4UAojMX1
zjNaoC+GT+rpH1Iw2qafptrTMe+R0dCZ0x6tiLL3t3MKGUybRN0yQcHvfy2boi8Vvv+78I0sm35o
9jMc+zFsShmdcZJS8wqCx5Oe+zxGk4KOc5g7Nn8Sem4bxvOHHkWqPkI5PYCI22wMCMPRfigjZpmn
cJQPOHYCvlGJyvHKOSG92q2oLR6OMV2XDDbAYeqCfdnG2za0tmeZUz3r+khJycjjCMNRt1iEO+Jr
Qo7OJIGhK/YYXBRdHPctnfSUQ62AOWKeEqIj6tkgQd+vubXlNsfoi6k7jcmL2n4G5Pwrvc2JodH/
QuEqc3atVcCHrAE35wrvsOkLbwBEN8yX9WaM3yxkgsvpvyZCeG1sp0XnVUZP7YkBoNVZOacJaKh3
Qg/fRak0p461bZJHGrAndhmorVc7C5Puz33SdWd39Sd4QBIsS51HqlyS7TJwfAq86TZlzJ5GAOlT
j2TnmNMbhu7it9ZITyD8E2rkJEJqA0D/2nVVzgJ+KEowGtLyw9DU7sohgiflB/O3GNaLXZtGIu9w
Rodc2/y55O+qXuJ9HA9EFnf14cUGwlrcb7VFAkji1mJDILyvjl562aoiVs78An6WiW+qO9xtUaTd
AG2m9YnFTLxtyLpWZCKi2ywrk6BhWDkgc2f24n2Ku5DUAezLLA/egtuuzoejLiy6PWVBmlSk2s2Y
o+FhXbCCNa+tlH+JCNxknpwo2W3eRUs5cUWeNImAHSBptV5CDQyHCGvfEtwVZK4tLj8maopPnXAE
uFdRblEHJXd0y9SaNHOnqv5olhF99yPUSb4BILCEPgYuDX6ifkxB0NM6KBJgb+aZdrQlXE6EK5v6
yQDjYErMCLDEFmhhheqC/uhrhyOStYeLvHQVgndYsNVEx4QDfQ5szPohFec7UefXd3VdipQ+EL2O
VPaKUPYsarRO2LKA25N0D7zeHa6fwCdVtuvgILc0EB7DuMfGT+m/khX7OryRHtj/oXarl15VSp7l
cRSa67fZMfbuU6V0m/9XUxnk+AmXTBigIlc4MXNAtq6xWKARzBb5QBkuUj0DwTCoyEtqEoVQLseW
/I9tX7aLuhCamEwLaulK3QKyeJ+ygeghVAMQCwsF7LazF20aMzg9p9RGGeX37wYWZbjV9QZ+Z8gz
VXeQpancW2zwRZDtX5+dpzUY7bncpW7/E0n3x7/9GGVDmfJE34EfMGMd4pHdm2Jwj8/5KJNTKovj
/BDHOt+XHzvul/nDBO2jiM49zCEmVh6sv5Uoz9L7ZjAjIr/utzdjdpxpsbWZmIco26Sc807ubkMX
6EVbpo7kgR0cVCc0w4jbDQeNM5h0Cbow2uvYeLqiA8mCqzBG+ry8d5nQhC5s1W2gIe9F6GU89+9Q
pjuU+C/IjXXEUTJjgc43gUxufWjV4Nc1869Zp76iJ0dt71epgs9bxB1vw4aGnUufmCEGO1yb4iLC
rzzw7RFgjq2ivxCPO16R+99RX2SIfk6jz2IrmQR5aENPl2lbXQwzpXy3is6bWlyzSf9/yYX2dJWD
CaFrB7WMuo+oSduIlju4zazPDnppjVoodlqGPChqGLGx3dB56q9JJhIgSvwGHkBX0cUs61Sw3RZG
mp1hEvqFepobgb/F6CqFwif9EscEOpQewGBycSm5ixyacrSBW5C03ehb8K2ygbzEgSfHb8MWuO4d
rIHKKNTLhZNtwA4QUGsoHEVKzbeEuWiqG6HD7pTbc2n0GfpQ3+GXL0XtSSzm2i3OXzWGKxTlF1kh
vodnl+KvAZwKr+2K6+P/5Ox/lm5yRFD8MjtGSvNN32iRwT2IQl7JHzzaRNeQktsfArb+oMX5Tmi3
J7edv3tPT7o4dx4IaNYBBw69VltGdPmaHCX3tNgdz5LHviXmm/kgcaHvbFOqseqzXTQtDMsLKR4r
Ob7euWoG7/+WJsNt4gAvhCkIEHSC0WmN16k2aHgxj+NM/clWcMvtj14XbYRryqX+o4AvFkuxpvDE
fhHNlrZYpaCWtAZD0t3RXcWj0tEU66hcS3A9rgAx7oYVPCgK/J4q7ti/8enGjFMXHhmMb/pKykSo
OVrlp4LJomgM6HuLiDbHMDTj5D0tK1Cmw2mQxLKprY0xJPU+40sUsKxjkYs6WYfPT5RCihvxzjmb
h9DAJB3Z//oQ/yVtUoHPDStpf081RNy7Pi/mGDaVRs/fPbZmc/HaJWe9xe+ZofuE+RQvbe4QXc1N
h9K4yM8gE1IY+jt8Ikpqfn3+KX1tspkm71bbJNltXTR99lyhtOj3g/fPt/U8U4WlgJILhih+qIZG
C8TQJriOZ7uiOO/iLYffPyPs0HtVO8C2g7m+Yh4l0bu12KzfaVHHhG/pK6x5hW2AOuk8UixTx75y
4E0G8x6sZeZqu5nK+4ykxWwBjoHdQlkmgv6ChkJ3rjqsjAa73uJdmXHinFN4nHZ9Tjob0HpGX11b
fpG9usE8mKHdmS1wSQwFGQEvRLtxE4t8hO3WCnIKMIZWlzN/N0PGEdC+8cAG79zzVyudjV78xlbF
0RK7KyWw/ARc+asoSbJkreGeS2jLpoZR3gtPHDv3FGDpRxS7C5z5f5pNGqOk0eMkqUB4LSgY4cbA
LCjhIjbGycVO5izDknwy0u/D9ODcf4ViGazbg1DG1xvfFjlG0F9RhpwxpU36ioG/ZwMTrOQI8qOd
iOxkTauWpFE5Jo6uWlllkETCYrs3TMC5tkfNZQ29f2FWeH8yHOnmyEVdd4/LN0lyK5Uo6NL3OZs5
zohClSEv/rkoK7QRiBdSrrS2iKbc4YZQOnbHUpT0Ct4EDQpchuygcuCCvQtcNZUa+DEQQ8W822aJ
LPqbheDWdis9Rvn0vqBa9mWHVrMDJwAyU0qhosQV7OcQBt578I+7j90zsyYQZztebRzRlfr5BYV+
FNI0gM0sV3lrExd+eL3QJErXv0c0prkt8mqiAONX9wvhHWI/fnjzu5gqLRAg5XSpdkrCrg9gMoUJ
jf9Bw2+FAYNEVSdFW8cLOr3/NnubV2vqSAaqj1+2xdKmgogFuM+VJ6L2bfPrc9H/Xj6nD28VCr+5
Hrih5jaLmXJUVm6w5kB0sVL4UjbAfWvc/UTi9pMDWyhvZ5OaDvUzE+huAaaQBRI2SfsGecv7Cv1M
kgSFKYAVj9jjbb/4ghlG++x36r8mT5Pg9gah+stG4EjbCNR6DTIuB8QBiG2vrV2ocj12OhholPKs
B/aDLmbPkvWafeg1uqrpWAKHM/k6r3DN1kSHTIjC9qek4UhymXA9TiDkp2Y/OXpDEOWClgS7Sm1u
rNpVkgAMNNncRowBYVP/LkrAmyY5HgYZRH0Z8oSgWEY/Yhcf3NC9n827kcLFA2Crvsu8sF3tc4a9
aQ6cckPGlGOjzk2i/gMqxF+SLNT4tKjQ4PlqzUqmemRstsHhHdVlcoLHzsZKP8VvAX0Qo+zqaNjC
dn6x2lW27oZAlqmxn622paWUygq4DKbtP82tdZQma//Ep4Ddt/WIdmnFBg5HYh+dqJI3bj4fT9MW
n5b/T634vripH2p9dI8mWvnASxZ9DNuTXJyMKaXzsvdhWTiC3FKUd1g0QSH8wpvpcFGyEwlR7Lod
FlX5sa06TfbNFFIYBslOM2H8sdZ31usyfEMenLEZEzt3FdPSGiFb3bu2jZojX/ZWI7/D5lwj5mri
4uWsTmAaExKZyP4BlApMC4cNuvkg4VZsTIvwD6LTMRrZhfE1MjH2CwBRN+S0UmQJQp0w7tHMEKPV
UUw49tPj7pZrdDPTaAE65sF5b3q2/5XvRbYFcDUgXEObMRYEtFwjCLf82lS2jKlGUpwJ/IBw4b0g
FuwqbBa5xKOR2yUyD8AaNHP5t26cniDuQ98iM0Sj+0mxnxaUzhRYd1XSDo2wtIXe8racqAmTfOtt
z6CTaKAlurXg7gVB27KBjr+WPjDfO6vakRzdyDRbNGIJW+aoYW+6PdKVuZqJoRusQVyTT9jF1wlW
xAhU/dlY5Y28w5wDmsrXTsPRI85HQE0cz8Z5CP7aajocz5Gcz8HRxmpEXRhHDLqhvZAWpAzLnt/B
GIlqSyEuhI1qlD7kVF63NikSy6Bn76bCnLrX1W5XCvv+w3Rb9Lpa17Zdq78mgROb1tEjrRPZnpp6
U0YWtm7AeQzxZgW/s/+dgo2myP1FnmNghwYw6s/pJodpJmoSCv+G3pj994mWBcvvXrv65Xz2mFjn
GNaH7qVtpOHMwJnU6d6+EP4w997ASqGsHXt4QZ/6A4hkIGevsxa6UWjLOzlh3Zo1SrcoZK0bgM1z
tEPm7upIjPuGfX+d9/aY+EjP0dtfwbFmtuK2pVZNbjMrkpV/XA9pyVe8kbZGBzW2ayLG5MgscN6v
cyfkRQ9wAfufwpqslcTzqNYsNuiUrxj7JyXc9aVRjsohWqVi4TqAI8EyfMvk+qS8cuVfLZZPVWep
2Ke0KSIcE0jiPJRxz/pLtuE71B8pnVM5qH8lNkEwDxbaVZ1Xjl1CAvM1ASaGMUN+fDLDw/QSRjmM
AfoR1F0Kbry6J4GGkqNuzsYXtOE74dVyshBiJhIRjeKJN92V9nbSWI3dzRTRqnn5tFOIB+n1dEAu
bYsAlo/Nn6GeEpIOlt0k8WPSUkWizux+QRjtb4+1jY9zkbggs/1++jG11poAPcSzI4GbsReyE16i
xxECVI1d2bkX4QIcFoqghpvPCIjy5rdyRtZ7OGHSccNxy4UsbTsoCCkEAQ6pQ8U02+1RLDvly3iq
OSyeLAfbo+yykctM9XcE0y83dPEb7rd2/vZzGpbunz05GApRxZvFokuPk89o/U9U369CWzIig5VA
21IF59h0UzdOrujBC8JdqH4XqKsiLBm5q805rSALLAxDjofjtbQzLgaQucE/+dWUw6n5fAboBUOZ
ENm/YfSQ8foKH+Z2Vlh3sjLr8mezWDEq0Dds5IVnhIMunIuRXrixplrUhB7j6cdnBHiltWlIXVt7
3m/ZLyS31l9Dj53hDiaDujFkFF5pFB+zYLANzHPymREWaMLW8njbulG8MU2VPA5/pNeQz/EGtVKA
Kfs8dpm9basbV0ONA4j4WBLRJftciqJzhEWRvPL35hSKX78IenkmCu4hdeGpPBx09+x52R0fVPPF
BwRWInhbLuxPKeHtczOYL6jsIZFf4NKILE2wBPFOjdX7AsyQz9DpEncNqhbd9XBBKI0fzDwQwptG
Egkr3s4DDwHFEzlcSlwCkLRafk/3RDyp1MxlqVvymPdwqlDOYmyfK8c7QXkRpvdPH00hHZ/9OnMG
gN3Ac3nw8iawkwKbXEQphBgAVjmJ53hmqzNDWr30usb+NFC4hWBdomBr+z4BNsqHJuOcpERnaaiu
dWElLiThbSBOKhO10FNftFxSWMADaktfLNYBkXMyso+pHvGb5jCLp7n5u1Oqz9r2EPp12azoqUFS
O30+w14gli00bpW/iVP5IcP3BdSGvsNEQB9M2mpK+nXaK70nxsAxvRXtSGkHYEIaJcuk0KrAdSts
lTcx6qA8OrmgvSW9UK+uF8G50uLJZpYL7x3fcV2I0HO4EvenMNTcEnhuWNKwHHalGxxFFIWlVefc
bhBXw+7hmrUPOZNbtk3sO3ygnkADI6hZKmTzTSMTIKysXrSlXZlLx3CYcarVpoElPaZ3XAalossK
gt/V082L1tY+LTIX0uQt/GgeEsn/BEO5YYOKnoFVpqsVW0hH4k/06Go5j4IpK+JkQ3v3rPtQfOch
RjdX3EGJpQ/QfZ4KakpbyrylmK3GIOrU/Cmx/mEIPRFiKA7b0T5p8n46IqZaoRLoSWib7UnBNowQ
5v2yNpmsPkj4flRvTGObAjr/vrenz+FwuGFjJhdwxqKkrcCBntj9eVHUwtJN6VZjV8Tw08Zt3NR/
VhAVBPM5qGNYNfv1uIIhgZIThhOXLMPXW2s6ppU351i3bwIZxa2SdOwtW0/zk39KYp2pv4i11tg0
LGlk4K3gcarnynXQixTMmATaeEjOxLWaHS47O94rE8G1bD0H3C0WSui8J2hl8vQYYRRdhdZUIJJl
SOx4aDYdMbSghovWxDWU6m4DZrQCyuDgyMCI6iJsD6+fgFY9YgBcGomdmRGU/LabT9Gu+MrgNCPL
/wP46A/Sa0uEg52raY6ibwKXL8PAKXk64WWMR7HgYKA+pU3dwU46iTls0k6L9YMWBkiloO16xFFc
+SixVmNHPwok8nD7fZ21JqzQn60G7l1pQ+Ufv1pS7p4t1MZxUA11Ds1xVvTiHHctM82C/pQhaYhA
0PBQhtkLInoMYO32bf3F/xxuYLYfcd0hNXuF+pyarJgUGFb0l6FsvAiuUdC5FbKiMwf2liwbKmkH
EciVt/vxQOgDiYlcLdUrszBDC3EdJaFv+W5qfiVlb8ZzhRskaDeCHNRK8LiDyvqCuYPMOs8LnwOv
Evvk771w/VXdYYUiqwdQEAJ5GJ/6q725hdKBHPTy81kWSDUXOUHDo2QpLX6RT1KVLRhyQMQ6uJTt
dHImsbiBMwZUg/cOSHd7Blop0UQSI80fQlzldz7sAZoMhdWOtw19HrAAf1Eb+8EmQN8Ajd5J3hSJ
g+vr7O6fHQCXbNGRcU24H1ptn5FMWjI2QazRnBel2nfBZ2xKBP0ECsEg2IRoE9LWek61ZfttXCrT
bQsSzPwlWStAK6DeW7BVfIie0Pd1aBXpYttKRr9a6nrj/D0Q1SwtW1jQrWwB5X3dMCNWg7KGbtkm
J14rZcRGpHDLkmuP3NNKedevcneOX0KTvylLjgIc+Z8Jf5KOcbFuIcGQx7KVWDawGzOTgWejB+Gb
HTRZi4XeemWiPaeOBvlDm9pM0hl8oJzauD8DIkPjpf3Q21aV12PT2G5ulcwK4AupiEeisQI5++06
Mrn2E261mwqoL7m4UCC3C489OY2/4Mw7WXs10k5eWKi+PpcJqNYqcoVn4g/wxu/FatcqTUnO22jI
uqkJjgQCcJIkNP+E/ZD0IlOXa4Ylv9RHxLXtXSE/8HAdxVT5Mz9/jM+s1JkeWbc4oKyx6ulKUS62
mYKamBN97IvQQgl7qiqHYQIPDmvqzuiQP/ISzYwgWT54CnyVoVdYHRMwYxXZg+bTizo4LJNqyIJ2
H/cbafdsKA3/3IduD2LvaTg5lI0nN/D6hHHie6u/myWaGfCK5vj4KcwXJ7YiqAq3T6QdHDdjAKOA
yJxekoQ3jVocM0vkffH67XRjDgrHw8peg44kMMROOaOtlCHEJIZ1g6qZmB94e+volGQa+tVpLmDs
NPB4wkpsNwHROR9vlncY7tNtfrkNY6WH/rS/gsUGYN8RgbMHTBtjfT1BA1xjNDtHoGn7tep1WFqY
4u39K3Kdp2JE/msyQBCSAruyRGDrLNIzoJiwohqrh2+963EUwgRHuZB+fxqFP8MO14hEZz1o0PFe
Ud7M8A7yASyzWolaoCCQaQUk4eUEScIfXsByYYBxfPHvIZakmYsEJGuXnjvil1lrtrkFvyP6vf3j
0ltabdS+9WijgZej4Q0FCLBV3iX1uW9bq4kFMOzsiBjVX+SHssKgEGBJnK1vHy9kYV3ZDgf1wi/X
vPQTcCgC7oMAP75BtA3az24AX3xDniLyybtspzxO1r+/3At6h02iQOlkpGP3NRfvXbbv2cn7IVYa
FG5+RPtY/S7L27tIzVkqkIZB8TdLsticT/vTQ97q2g6EIK8jkfD/a8yLfN+6W4EeXxBVflzGEs1N
9RZkgFqZT3Bs171efuJVUOkoM8dCyowweiDoZWtnyUNPc9MXorxWTtpv0A0Utc0Ph0CQvzrYadxF
+ztqaMDCMMKcOZHDYzDdfUKPY6HMDLabeo3LFPJvVLmTqAEfLY3PKnAGwCJK6UBjoUQCmxJdBOiu
Wzbh7FPC7PH4c35Z/n0y+4aXUSH6DhECXrH3piW39dvzw758mpM8e5zcT7Pt0C6IH1MaKfauxv1X
BbagwqQ+3H9CoCq5Xh7po7ZLvaBuDG6nre6ehU7l27TtsKXDXfwcaDy058ICEOurt/k/yGpkNCHo
aWjNdLup0Xi98nbl9ulU60srXldPdCBA6gYQLDpS6E4RxujwSdXeMnrML8GVIL68xklBuXsG2GiQ
tJwCnej2EVlvq9Rm/Ve9WldwrBkmxMv8qTF9OpJwmymmE/XhewzMUEx6lPy31CChtDlSIhQ73Adp
NvguqtPjBX+il0XePyg40CyGS4t7c98iSKTIVTa1tYziDg1ng+pjrmYpHULDdVppuAL3CEDmZ6Gs
LpOP5MS2e/tXTib1ddc4lch98y4zx9lvPpt7nfoXv6LWunLONTkf+Ixc7arKWvEDOBvAghitzp5A
ke1lKk2UyUUpm+wmvP8aIyQthl9dF/9rOtgJBHaGoRJjBSRWar0vv/Gl//wEl7pwuqfBoXRLza1i
KRQ3AbNycFmvZCYutKPPBj8NLlY5c4nO7IbV8WI9qMgnhbnss5a2fHL1qKVJSNqDgXAIJJULWX8g
AjPjXyH4+93DcATalQ2QQw4IYUiDnryMhJP+/tcTBNZ/4bur1WJyiYIQvyoQ/y4gH8wXAi//F8Gx
5ofJn18BI5+akq242PJYkFYws2asxdjMZb2L0iq3i/JY/hu5v8sra6fCYqKunFZc5WMEEYImVSfF
1xOSQd3RXRvSO3/0UMhgKIU1wmPdPmNEIEwt0Tu3IHXMs8RdgVEh5LxIPZS5qiBmYXQ6+ujOYXJ4
/iLB7tbwr+lbRZDkD8jWEBLCU5AhEri6n8XYXnOpzHlAi5sIUanO4wVNSWZJN7XXQIlAYgd1EXPp
K2l8WDTUcQuot7RVnC69C8JwPVsRqeqHoV5OBG91+5ucqci7GzfHmmINiQSNdkca50pUSNtXCCSr
Ojw3hGSYOo4SxPN0Cz3MTuzdsVeq9fejVKdAAhDg3Fr6cfT1pm0nsvOw4JnO+lUZYXMLPmUl6cvk
ZFryeKnXir04m6cgYvymukY1Do14Rb8sYMJ2PN/Yl6OfkNSDdTLJ6JG4DZkveLvt/+sNy9V4V++I
HCEm9ivIoDilWU8KceCPeTp2qrWKIVloGeXBO9der1JWkhFHel0CjpElbX0+u/ZnDWbINlePBSvL
oO7MOi8bShRXwpo8KshcgFFD3nxyHN6s5+HNnTbXVbB/T7OCUaO6zYE3fJYoN8y/RrGwvWps0AyQ
P4Cwc1tA51yMK2u5OhFLcrA10HT9Ra0l4Chf1rITYxsvtVGDLh6uaaTiWV28bNA5dpO/ATjlJINB
PHhr28uY/5sqp3gtvj2N9l7Xrk5trwtxoyiN+JcrAWiOlrDunVODgOCCaY8Uq4ZA/zAWiW7eV4ot
R7TCokx8PDpbCHYnh946VF3hA2X4ETvS7kq2R7vrT7NwywuXy/oVGA5Yegq7yF/KVrA4w+iI6xWy
FZ9+v3sr7F21DGf1t1FpZKLqcyo1qNU5rsqMr47NvPrKjwQ+oUBrhIN+0y1rbDgwR1/JHCrK4KJs
EXv9Pnh7pfOwMsi9Tkl81xmzZUVYkv58mQ+7ZDGS6uiu8eHWUQDAfcpCJ0kl85PAUjnrHhHextae
udnbCj88uTi+Xp0qaiVvusl4n52PJBr2lxWph4Z/AMeE+fPMctshz9jLpmQt3zYKhIj8wS91MyPq
WtGp95b8pL+RLSooINPxQ2QeKLw2KATM8wHKhVmcJ0QmM2zMrVygiyvI2CI9rzDD5so8yiUV9meB
KP5gqNN9qdEGl/VkJzMNDx+6TRebX9sHAQPbq6osHXN/zHBqAKqh92ss/q0srlB1sVMNwoqgFQNc
ndxWczJy912qKzX3eslhnQAXldWJLII2wtS/5C/L7cAdsK2oq8myhPznzhedj54wD498HcoQG1S1
YnpMClnNlllKFbuFV4FR6e0vRTPlKNHIrma+TCaLNSnyaZIWlqhCSbWw9jdVWt3L/BHTc+CRe8JX
xtB4nyESTSo1Ba0E0lUXflA7BxmvHf9KTy/q73AaS0SBDJwSWPaiTLMd6FFSl/1Ef+uUapocikGq
6Qp7ePC5+LBr/qrP9CCZFI3y3q7mf89X1q/Hjqbkqv1NzmYgJctLfqBC/I63xfL3tMkGR0DCva60
ymd1FwAb5EkxuGr7QQDH5WFtMKGhrVpao2M21YLh+N0KsXcy0foB8DwucVaEY9Je+ItWz4BklZD6
Y1o/37YKAOPYVPuGw+O+zxxqInDtib7tczDFin2EgLHwahjz+A8yMc+CZ2oNYvaDECUZWwPP/Dwk
C0A7IHZunp1POIJuQDVFRg7RpK0ZkwqFwSoijAJybMxGw2exB6oBnCvE79wYEKh4RANAtD2+V8GP
k+5HCZA/H6X5uBRKsUZPmv6atH461SVEvzHqFLzucUuNO+BwcCPehz7ozlSBzkGiro7BPMt4tCbb
IYcW78n4wNn90KNTZEIFPT34Wc7bQCHuHC/QfbJixQQyNxqkLYL+3mtWocdeLchbZLaYNHSzws7j
5A/lbqNcfQ1SGFpYHU6ec7icbWUBXstYR2si+pMoxXdsx+rf9MpiRZ+T4G6uchYQS6DOWfequbrG
ubycsAR2dGzHrnuzCf2EiVG/SkzDPYNbvgfiMWlW3Xf1nPZBWU4r6gkWxDDlQWsQgzE66ZCLw1Ab
dayar+fKc98i7fA3TTnYt27zMa4kCkoIpfN8UKeRPp+Z1I+hq3d6Xh9bwxYO3l9nruVapWJ3io/V
jkrlnL6xd8we9NpW4rr4sW9u+vdpOLX3D8Mjf5uUD3RIeE5B5863xijEFxxd0gslymeqpBG1mcaW
wVm0gBwGjqGp0dsIP/zwZT6DB0wdESG8LcSsnHxckkVK6JAXlsLGD3Gm+iOGOSuCNJ8+XfH824W1
mGLRh4kHn7iVsIBzZai+kEzmVvaRLhZKH2WGqPRBL5GWD3whFRsAN6jko1cTtXhj/rjwsvwDKaRY
el8ruW6GD1ztX51cloSw3ky//1PykNn6OBMEALSkFVLFqSK7gXp/iq/5h6Yj6DbI2NY9TxUTfigF
Jrf4Zf1TR5YxzrGXClbGt8UrZJvZ3cqjmbhsF4MUswiCV78LjuVSw6HWlyguF5N4s/qdB/8u7HE1
NIX+POh5KcKUHYAGnl/bGaAglDkIfr/7KfHYhkrvIqsP1Od9sYD8cl2ek8OrtnsqqB99KO/guVIr
VkKyyaSB+nFaOk1gVuSh576BiyeMSCfU+5wLzoRgQjH7ME71rFuHQLO2+P25fYWr7aqvfvZMpXay
Wm9N3bvonnJd84bgMatL1ND8Vj0EBWBHub4YvGvMYj7NWrm/ir2s5KF7HKzQXc2HanKhx1YcVdrB
6wo63pxNQfdC89An8860He1Dj7JMNl+O7GDyOUgYQZG4D2IF4u6/n+ZGnLgdS0w7Y2Y0Q2F5TiiW
tGJWoXMiE3vnbQlgWYaxFlPluq4tiOnmcLAFTA81P/wq73D6PVIzWGim+2buctwb9dyEddE2KVJ9
rHgcynI4kvZMYKmvGokxl4A0dt+4hHOOagRhAHE1UrnEPTdHBpQ6DUtlpMm31R90umdEYb8Zjrgg
Z81HE11osBXJv/fnOft9fGHc7LlZA6Tp6nzKxhRzkbHUXxQQPzW6DmrJl/DJWLTeayCy7N4nw6b4
6Yb9FM7dXcp0glMhrNMZQ9bO8VDJBqzdeDSABsGsF/TP1TSdFlbQIJ63nj8zGSCRA/aTwR1M6rCj
yeP62Wb7ve/s/mk1VvmsJul555dx3zrhf8Gl4dk8cqV+sjygvrlFCDD+MUEBZIFHjsqm8wiai4sh
fR5HVv77RLPZTNc45iKcuLH0drEjw4x4E/NgOAcVDjwCTr32jxl7B9Gsx+uhQ1fv/+8OBIykbENJ
pQ4mMzUbyxcLyeTmXJJdhucx81+QhxjFAgh4i9SYT6BglbuXODZ/vkeVJ1AJu4njMgV9y2po26JY
hYAWlc4k21LJnqRctdZFhoF2cUFvQQGi+gtElmx1MH/28fGR8G9QTtK9keE72LwglLT9FDJ4+6H8
/Ei8MlJ5KAnV7OUnwnp6mFN2CszyR2E5ih+4gGaI/dierULv65oqKdrUvxuhm+W3ssh3yIG8dGBG
AZJy85lnj74DyQu8XCbQ8t12gn6sfOCkWJKybTExdkSTF4jDwGN72N+joREcYLyvzzw6wqd+ctP5
lhObdSsLg2gxayJm+/SngL7WuJqRiMo5T+HOvJQucZkwCFnWj0MIa7tz2dM36LVXzRNHxJoXcLnK
BzsekzbYDmV3XycomTeeCQAzmkHzoYuDXlaEVDOeUsaVafLpkoO3V3i2yjKVL5sHerc0Pti+K4pH
5nDvMpeEwHIvkyI46dQZPBq4rRWsZaVEOBBWPtw5NfpaZN9mmY32g2jfakQkjd1PBh1EJ5pzxub4
wOpMnltyqZa2RyS28AptCuZUqaE0FZG9PA0/tpKTW/DqzK9Vrxi+N8CnpFkEYFVNJRJE6dzXD1Ax
luwwU6mE6bWjIUzzNe+X//KUYzYvO9q9+mBbOFvBk0htOk1cpwttUlC1uE5+XKfmAPnZ6GEPXLwq
7/qBSt6+W4IZ4Qzzs4lf+Xdv0w0jo78aqEk5Ut0Es4Oe5v3VbffPdT48TtXw9zZj9zo9vhnDff97
ZqvCieZQn+SlZEtbD0lvrDygC9ma13yMOTQe+DCntOvXPJlYwPmeKS6i195L2YFTObSt2BvUd/g5
fFeczeCImIIE+2cOqTfpM0HsWbpxJVJ2fTNnHxP7UK7ZMN7GGtgirPRt/IPVqEZ/gnim7olxx+9I
uQbXSN8Cr03Ik2r/ysoYO1HKdBz90SNOpWbD1bYYFH1pI3Mq7B1SEvk3OChk50PWlaCAIxuBPr5K
0sZKGYqNnsbuwc2lpY+SfB88GJdsGToDK9o5dXXGJ35JJNpy7aBEZBelW6iTLW/4KpiFXdnVNcvJ
a5Q4fEk3c52UHrFHvQ3qC65fy9oWKMcTvcYC+pUggAumWjUWzvRuK6RST2wQZp2O0VegLzlB0v+B
LdAlQI+9mqRjhgfPCMa48bnn3jxbi+b9xBv1FS4l3jDdZPHza+YHrO5L1OWVX5dH886wEDfPRkVh
BkoKYzFyxpZDbA5wQIrR3+EIf998RczhNQTVKfCv/WulqrTwZE9dqp2KsK5p6gaT1deS6mTo4hM7
ext4T5t5gTuvZAwQAFg7TV078hlLzyOmuybw88B5ZBl56GSpxWlbUx0YG6B96zwTzfO8aGzPpVJf
E1p22BPWsPVmkR+0hqcPWfb2wQRRka0GfWyP/FG4i5aLJxVZsrhgAnsRyUVzIfRl7qD6Qdy+2SAc
g0eCaqWNUjSEBoylTypAtm9lv+HDFikyua0NTlrpDGMxA2N98McJ2MiwzaQNpb73TzLsISlG+J8X
hj3EP0Q9wFzaHcC36IoMcsrC2vD2EQ5sDyX0E1sLVoVrluNCQtSXfIKUdTpBBfJt1zoe18KkVlo4
/Ean3gE8dfyr94HnbcWnCytFLM3SfZHyHo4/+UJvDrfuyAD3kn7Paf7i7VsHTADCgJIav5XmRVtb
B49DLSvzppMOCsM6ipPeGw9UAfthg6uNviZwfRXrOxcZAkZwNAxzR1Ug4QfF4/5UHQfWZPDFpibq
2YprUcnzBCa3Me3c4bhYKQor91L6FKfVgR0DBn5kXZTbUSGUtUQKXt4qdh/TV+/QlAwEuVpdNz9Z
aBLUmEqN1y3XUkLQLfjBHfmRkIh5u0uJ5NFfLL0OCdJUzt6XI2cbopiP5LpZSd696ocnGrXgV8rr
I4kQ6waYSwPFoT85UawRFZx9F1Gy3vTaerJT6dVLcDjIaTUy4O5kCGmg5ZH9Jml9M2HD2lrOQOnW
SHuCbQHN9CDXMlTMr7x+dKCkaZTTteKMH8GlAzBmHJNpVzTtdFwlYNr/WEPjpL/C1Vn7QvfGvNUW
rrQq8/UJg3LXy/RMi5iE8NdIxFhgQ0wCAMp+InqEGj7n8zPsQOpqoT6H/y1lAIiNE7vw87wnYQCZ
l38cGRUsirN/xl7Au99aVzJsXmvdAGO7KVhvU0y03A6G9qeufP89/5eEcHi+wIol/ms2HQ+54vyb
w+RbXi7PaU8RNAhfbj5Pia+se09eQfcrGkYa/VSdTirVjVS6p0ujYoQ+8Pq4ao/KWdZ5204Xz5eP
kz9UGnqB7wBA248lor740PbSUbL4DvI2hKylnIhaWBEHtGW/ls5AfFrsd927Ptz2t8SzWVZ0w1VG
zagD/R0wdzEN6pB/rePNgaq4Fo93LakJoYnRqp8UMu8XHGao/bSoBkjv+FzuKNFzIX9/NnRPv5jB
Q2dTy1SKtOJqjOrzN9FxiAv2uhLqVUOl/0E2naZwutbRuT6eouystmN6XtRlBXs07rhiqzDkDO6n
fIW9FBwyU9PxBXXH5fJ+t1XCzSL/VJnN72yAXe00g6SoNWW3DHX37rjZ+s3/Hkhroh1H2teeYyvy
Eg5DMBspqiLP1SWlR5LK+ba54tgPeNnNGkOHcaedSpltSp1FOxZNxfNwDrnHSqUjmvLRRJ/3dWYn
3BPDVeuoOUuC5eSBJ2vV/q9nJW/g/aNPwCj54aursUagyBNKMmFTLFBf2eCdZw5xKn4po30rXpgO
GiMirBBLhiRQjz5VuJBFbO5p2KPWmllUwZDjm4qeQLIGnafwwuhUj9hx6Z2X5VZnkBoCm/FVmcTL
Qwa9E8EmNLy2pwxjceAhrmaL5WdAcQyBvSIz110gU7rMExHi1Nar7fcmTpms4dbZbvQm4eDnYP7K
3qudvMU6NriYaBwy6LYM4s2UAV7wo8TeYMYZDUiXyYHWjM5n1XIS+afDqcznGAUoBuNv5XCva539
BVVpbMnhYxnl8Hztxb9YZDfsdcrF+M6gzbn0CvaHN5AIJvlP6mey4rw6plVEyhDnkN41c7Q1HvOn
HHJP8CbeC645sW60KX66YrhxIPdMj8y6iPC3P6/pzlK0zhhXGdDIfMy5K8+ZYhvkthu98W7GdSAk
c8FrQlEY4LH2i1ztz9sxwLgMf+qkmJy8yxwnvRppiUXpJ6AbYXuKpfrMYYktijjG/RkDKEYSZQeA
oyOxNpIPaXOgxkqMOPmkGFEuhAEfTADp0JvvKkVpsDFKwdpoOv8uFLzySeHkAUmFC+b3jblL6x1/
Nq8oZCOpLUuyqepsVvnvsuBLCB7/hLm8y/NI3SUsqaC4B8rzcB489BxijZkVHdZBkyYHpQ1H6TFS
hbg6fkvITE52gCSEiq28Ftj0FOsZFjIdWyVYxy70d+tsdieo59VLI8L2KB+90Rk7YS0lkX2yGMSn
0XiCq0SuAV3dhT8od5i5iP4aSyvYo4tA8rdt1Vdcp2aR9THtkJ3YVmmzLSnTQdfTqIbc6TD+maCq
LzOESMwyhLZeNkPhkEN1kebn21IMoKV0N8n65MuQsmmVaLyNcZaPadRz2kV2mptd4AE7n+FZqoF2
fCJUfleZeV7AFJZ/55XtI2lbpqen/422fNu6fo6Kvv9vCP/YBhG7qIpkk3SwTfXtFxHu3lyNP4pE
15jcim/jSQ0AfM9fT8sy/v9ZWejam11fnWALgi0cX1cVZbbcd8F7lrXLvS/qPZbq231sIbpeIbKI
JuY7lpbA0BCpUafYmPzRVa4tjmoCGkiE2lhU+craCQMFc8xnf7l17rqRz9XR+tQrxW/NNoRDzS4J
3qdsCvCWScv1MZ2vhGdApdkrDYTMFbEHKeG7ASsWgpjIxOgisjik6wVmSYzlla3HkQTYfceWyr2L
eI9JsRSCNTu+GFnCj9l7qrwO/AsUcrJkJsLwD6B6m+xgTCTaV4q61xw5bL+l4JQxgDNzW0c1FqLL
8rDLWaCeaYjB2/o2jxpXNBSDWudRo6IG2JO2mvwkDck1sI81mqjqvWKC9bZn1G73GPn8LIarEDy7
qe8pCmlIafnBqXeqN8JWjkMEmPUY2kYTNULWk9O9FK+4lSyR7DIQuvxXeoXlIbxQrFA27zLmf8gl
CRFWw3hGtmE97sENJVmxZ/ZDvY29X/KdseU9SPhFLIYY1o5ZjqqbinIjhI3FVsJz0/eEDKvJBnIC
+5EQHEkKxpUk0oaGkXViSFKDUKeJlfFw6KASc8NzENm9QhxBFeUjAGb2itT+ZiQfiF6VX58OItG6
GYmYF9WHebgarC9K5o9D2hKV8bupKAkDJ2ETQAXmkhqkCGx/iON/71m79pSLDDr1jHKI2a1mYa+T
0ie6jDTZXvz24iWPNIB+8Rml0F2T8EdNoFgYntXWBpc/p6PNX6KRf6Adfc4SCiPxWwVVo+CiEHd2
eyX01Q2iq9TsdGp7wHmqKXN+kW25j/fOu4QbeASCZB1mxmt6NNpGRHpizD/+7GLt54UogEkgeU8q
ljwT8QONXnvNBwHuvvlaSNn6mBDAyEKQN+FlYILC5HrPEd+rM3FMx3/kF61gqeCL9Xust7oUkeku
H91b+TsBj5F2kuMSPAR69R0wgtiia46eSu1Ou9qxbdp4c4WNaIAIQfUnnIkth9fQfy8zsTI8yl41
7R8vKJQot2gO0xp4WyFbb6tWkn1IHM7W09cCwjQcYMDcfT4tTSLfK7SWv5aSA5sX9FPa+/xfVoxk
r3zX5EK1ZAPEI8I4TxCGlChU+4IXBCWdRebNynJiOEp+0F62RoYM4vaK/DAPEqda6vqY5Nowf7Hi
XkeDZqfFwrscQPV1DFWJZjcBW2xVlI4XXTqCWiBYeb0M6iRiTbltXLj+Q9SSRzCDeeGS6cJqsant
Xs/hegDgDwxcu8djKDj+VYlexrmhpis9ho0fWnMGeFCTitYe9SeeFNXQWGFkdSke+R9aKxmtOdkd
FqJetsHzYCXMTkXWbplyONLOmUSsM4EhuKPvQdnS7CvE+NQybytQRtC1SKPF8hRifKJ1UzY2dWkr
3GSwSu40FOjVtqvpEqNym3MonujjoskDDozAGPSBAJoA+wzvQ4x828lkma+T8FVhQGi6STvOcNTw
rTTYMShVHOrOwl+u0hDExmh4oMYecvAqjLUGlhljJN6rR96xMsKTjLfUqNgL4hlsJcoYnLIG7Vft
Xm5okzMJEN42ezPXYnG/8ig43lMXKgT+a3kGvdseR0Um01pCsmUszQlq50lb8F83EbKQ9EwMkE3r
GI/iHninU5sbZv12dBr/5ZDpfQooz+YnMiwt2+cZit1bw1g9XjKM7WjSmQFLf2TA4pkp9dJXFB0d
lHLaHvfbyovQDQzivjxSVWdKP4DbFavXB1CZd8kyR+L/LO3ppq+D2/cRGtoYkUmcgKPY5GaXKV7i
dGB1X5iiVw1MpvPZlxChUL2xYtBpItcgUfFgu4wQ3jHReNAhDvM0sT/y0r+30Mkf70ponBSQL9uX
ZW7qtrSUdpHgWZZC8pUneZAssxoHpDKSvvVsfE+/2xrQI7WzlJyWuVnyKBJ1F7pCVU3Vd3geqwby
8JlTu/dAaH8+IEWzu20pctVNq0TRuA1zJh4iCmJ5mgBrLiSW7fAVjg+v7nFhh0yhRzRlK3zYN3O9
NVKbSl3JC4PiIxjbD6fVfPCzZ728t5nrsr/YD62+BmcHZzU2lkwKyInEdaRiEblHuLcoI6iu8Nw5
N83KQECOO4fkpuXEUYR8U/CsAFyBEzyvO+UJxeuG7rQLJ73Ckbb0OtW81QaIn8VbHDeR529RvkXI
uAdL5QNHODyPTtiS+yU2BGThRTkk05IfK/3gdRyPg8QF1cKElQ4p+rg+kpZKeu1nrgf1NYIt+ZBh
CT2p3JGIRZMxIgB2ii3XY17pGcY8LW+j0IOUVp6h11WoKXlvrABHlmzK/AWSrHu8cC9Unz06yG9T
J5oAbWzXWfGbAF87eGoxDq9N3dgXtwZrpxhXRtzLmMviaIQIVIzr+pFMumkD6clbLIILSuNRCi5L
VbIAVHBoxAzr+XpMcWafq3rdDXLbS4PeXWE9f81o4PWLwmYH8zZ+MxztVC9lvHvx+KInTC0tyFex
FZO1WX7nA2xr9dODMXDqQjy2tAPZK9BB7WwrrZB9dBJLdOXd/jsYJNpXLaJv/4fvbCPgF2vv+yAs
iSdewdiz/Tq9B2cOCFe2kZ3d/dPI1vEwX05yXGUX054QUIuW32W26+fdrVSi04BwIfqqUCEdFO47
QvtNHihM1ckZSO3waMkCkGzHpGaXmpfcRGIJqHSfN23em/KD8Qimqv9DUVcECqXCZOAof0NZDtnw
9u/71mB5+d0N0qQ2aYqeQyQrdVnmi4AVlFQW31ygmHfgY5R/tu7AkkJVOdy4xawfmxRGbdMqRE0r
8UisKR3aEUwOiW1u3Zb3/QdwDD6XBFaSn039WUqi4pZyBjnFeSNYsn0FYUDD65PDUfZDmcPWfAPG
Z6TZYDQnktDL+8nhQMV3RvxyR4vP6aOvoT0+NaKe78klVJOVegfm2rAwTlCMIjAs1FXBsHbvQgXf
VIgQ3yiYm+5ZUHfDfWdlnBdyNTty2sODduOxMxywS1buxHULahkL9GhRDz0MivjdEC9AAyPFVbsC
at1y9sbihzchGWFG+2KJfOlE6fOBCG9+7DPSZ34uNjHi22fTxKVuPZWFyVPKupJ0QKFteQPgCpg0
tSiS9OZc2Uk23AdwGVzeeMJsBXiWMM4MD48RyJWEGJy55+y5JARqkaecXhJrocc5PatllZleM0BA
mW6vQ3Tk4WvhCzraU4iK3SL7f2Y8/Ym9/iqSj7N7+5FP7xfPFsoAoZeEWgnspZCdhNiQNKlGl7y8
czxLZKuaAm7ePwLYORIwT6mxtAYdiFeeNOZ3eRUX8gwYSjUgle8YvFgeD+7p34uzWQhV1fscoQz1
faUVhbCswFGe1/n0kT/ILeThFVG2KvfziErX2MyKlRY4c9PVC2tmbE2dRxCi2ulPnKR1ZXSZg5uS
tb21J10kmDhVkMVzaxRxhJdQgnm8iT52Hhk4B9nzycB7q9gSzaSc4NOEajuRX5vfUKE+6zJv+pgB
YClgQZRtbWcRXxothfK8c4vN4obbe2uXLG/EEZTkLfoLptYkfmvM+Avm+KG2KfqRohJ9I4abp81l
YiwwUbhVvlM+TnhOzwi8+muL+wkVrG9tRYLwvNWtE+bm6mhy2YeIaF7ZMoHRHYaDQptt3rwW2hPf
/y6C0d6YCQcLJU+njlzJLX/11DRJWY0exBCnhA+vVGOEnZau5RCuTwW9UL1zaX5NybnQ4H0OKHN5
HNuPgHwkaUKsa6QKPNOUUqXuCuSrCQzcGe9RJLxTin58Gq4FztHb/zgf0vqMa9ETlehRhbs/6GsP
5H5hWKFob/B4/EQsk2mADW0CEik+onHFhl4XRO8VyeJUgfWaW596gEYW23jdMKdhcwZH2aUO3wgv
/JgjD2J5HJadqYselGYqOF1dm4evsRnkGS7WPnifGIVcsLf0U/H3k9Zg0vkUI/7GbE4IRlv2ZkWf
i0yK080tXkpNHaX2RZSggRQDoFA7SzGKbTZRwz5m6fLBG7EF+P9XiSQFvIVyF67e9ekHkSNu98o7
L7M+LccSsohmU7k7M5fNd/gFfcCoa6sA6fUpEwMB2yxp7zVODzEzskabpVSnE6NaXIXofkrJrUMe
KVVurOM4Jn8JTdGSS4InTU7hc+mbUGKgcDIaj39iDyacf28JPZC+0ElUsQgI6pRPAnkFfX4BKK+2
CCk9GWh6Oy2FhrifkNjZDvBvchboNAMbMqUYG6rRNxpMfX0whj4mrmu27SFA1l/QRs3pA2k0/xvH
KNJ8ljpvoyZ2wt23V0AdhCs4tH/8OusLSDfdg7g4JxM1O/ec7xKePov0SsLWydM3mJlj0P+kQdVV
aZCpC6VRjJ57NnETTWYPb9hOo6R328AbPdpkSH7uSlJt7cKS+nM3+syqbMzMNPN7KF2ONwVUFJOV
uVXTq01aigFSkxquyz7v8JkvBRQjyXTSSjlgeU+1qRJC5GOb+0npVN5ArIejbLK+Ym8NriBoff+a
exmmh8FTj21PmIQnXT5dmt+2Z7fySuxqfWiTGIxEX1TW9QEwv6w42kM1kod1jItjiLR2vSwyvgi3
laOl7pOOqqQg6me8i9MA8+w75RafnntEvHju5PX3k5zaTsf+Vp0Ovt7Z6F9CwLUVDqTwrLDgT+y9
M+V9fcqszddlsMQiyOo1sUh4LaPQUhAlBJqKHX262oEuxtVf7vVEKuAOZVy3MTxSnSTgpQ7OU9jz
TApDWDh8kbRRtsHxrgMebIfbik47QrXiXAjxt7+KtY/kVVK/x8RwrzTyd0RtwGWMWcv49fh+8WEN
9unYl0g1vITF+lwAhu5ksSSgj3JBy8dWx8F4twRaFO7aODfSVSDw6uJDTdvNjBdXg3JLUsEdAGUj
Tq+zRK8DtcaawyaFlmu905Zxp7LTTrofdlPXDt0ENgOhtskygcLrHhglI0OjfVc08PvTG81AZP2N
eWAF6NDA+Cs971aP6IxaejIcdoYAQuPveRGCDU3XNOX8pr24kEFaGFTxipRgSm8jAhJPsz8Bk5CW
eGe7M0qYaW+K6pacsc80QmXV5+MiZ2mIwO5OeTxz3nBGsihCNMFWtJ5s7JYVg7278MAf6F8l/8NI
HBaxGk5lI6NegF24kfssm8JrEIVC264FQjKj8bujgyI9CZZbPzihxUtTCCBWYcPSLAlcgN7PSeoB
y/8Se6BEBGHIbnSBYpNHH2uzCsLpRFsWL47kRNSzWTpUn6uyAjvymJNt0a9SOOCW0ZgP7EnzKDuJ
H/21aSAmztZKX1SmuOppojNHKjeLM25Rnb+nBBY2VmE1cdQ6laXhl9xGays5EbJlGOXKmSSC44Sv
G3GuzLXYV5qzJBMZwoew7vkrvaSw7tnpVJi1hna9JBvFLyKfpWcUf1WrKaaveqTtKYyI3CmRkUFK
tbBt9Z/vFaYfCQbqvU0ZYtzeWTm+AFOJGZTXKpGhtkNDvK0QPYf1tt3RhnYa8GcChQUO/BTcj2Kq
dqrXG1R0ytL87dBdL8jlgrv2HRbfyuE0V5WILLxxGyImmnwiy/dbe1T3hdSvff8IeZasQYiFz+rC
x0JlvPa5uIf2FjbfCnHOZTiPyvQwU5f/EAkiHe8nhWKaQeYZHgb0iYfn+atmm7a2RWnhDKMVzcMB
hp9GUGs9PJ7EVrwQ8sXJ90h/MafCVObzzRzkyh6j7/HUsyc/qvUv4eL0McURRSA35tITtbG/mH4z
4RrOBaBb1a8ljCUod8ARW1jF6jNzCb8wzC1xr78++Zpja3X3EQSTQEAlAAy4V6QYn/fE/ukLJe+4
29FVVuFbOz0m6Ges18KOgv++kXpew9XDL64zCVtPMO5rX0IXDOgN3gXYQ6+2h+aFpbPd2DJbAGDo
FFb+bBXKyoI6mBM5d7/E4Cm7MvUQ89SLsnj7vriQmS1VN0Rk5mF1UUfEYYtPrZq4unQLUoTsJ2mW
1SwFYp15bPh/vijL7MdWH0baUrfMBVvfr7O9OnqUV7SacLqEXY7RxpPJCrPO5g6UA7nb7KGryi0j
0Ut7Ul+7M0wGBXyD1K4+kUPQpDbLVmjcJ+T2iS5G1vS5o5MV9Hr6Bw1CUw9wjw3tlIptKecuVlcM
DUWD0W6iBtRF1Ael13RYytBZ+DbeSlL0qUcwLnR+1+j0s/CoClrQUFABRcrQY+MMpnQMvOGhAMI2
Xlga7vj/+/wn2oZSsGgwquDcfnUQ+crmsrtZUKqalrvOY/HbfxA6FUpLz8ZqEAzVYh6gJyKUGzAy
yUKQlJoLfMw3HSQ48AlaEDxkiEn9CPgpZOcuSLQ8n5HS3pkkbvu/R3qxLoD3LhdJPLnNpwXpDBmi
VnAvLT3wT1jaSO6i0QMMYjYyNRyzq7xuLzMDAQqCK8iKXEF1yuCFEHYnnAl9SUaxDlfY37SYMaV8
ibwqqaj4VTMapc9NfPPwea5r3WOxrDdaV0KarwZ4KmTr/Y8BMm/rryEl3Tmy4zEi9o8hK9opiOOC
8OedQbkzckNRoH1ecS75K9Mfc9Z05LgMmdhb1cMP6BYXfgKWnwQgknrK+7hyw+DejbVzj4zCfqr2
7Pm8/o0hnX6J+Lkw2MQG3S+jbrikeRv36jf3JXuqAybSKRyVWwXeGYYegzXddEi2sOobi/938++X
ocXT/MmAY7a/tJhYBKJxHJ6MoPmb+sOTN3vBNevIutCWQlC86KAGY53h0TF9tThQ9DVM8wRaKjSf
HnjGfP5FQkOosHIca1bji5rZCmlU5on3gpvSUJSDMHtavCfn+TxlS8AewNewxwpXrTiCw56H/N5D
xLI60vG2kpfcW5i27N04QFNe7YWxE+qLMj5GhFlWnWXrJ5n9+d5jzSY8eeWU5x1SgCs1HZGcd2EF
wrVVzWGVcSRkFMF3zc6AANH4+QVkE40fmxZQJTfgILMZAj913ikKE4iahn6+C0wyhF1ichZP5NIt
Qn8vZMX0lWbxqRKZ2HcAUW8nkZ+nk78nKkJXL3CHceOtJxm5jCIwCEroYoAc0v9eAECaQR2PnzDg
Q/ssO/MR3lSNdLPpSCFiFtIOL1xUgmIAdfsY2fxeF6ldszvW/G0a06tdrNrj8sFp3c2KYnOD0jv/
p+NLgW3ekGja/mPFmcwJ17GkoqTH/jE9w6LYBJbIO/6/MT2UR4bRz2F5JfVB++KpQhGp4uSdzh2M
0mxxx/S5m8INNybLqxx+i+LSGmFj4Ne+RvQcMm/N1Ix1xKT2jrewR9KEZN+B2fe1qZFuz9tJxsdp
T0Hrp/AMmc7y1ecI85UK7aub0NCeki+BuElGH0agUGnGKmpDc9CcxuLq36WDVLqnPtGRLwXFjesn
MhdZ2OUpYMdNYeK89iwOWmZX6AMQuO7JeE3lEssVqp8C2ulkGXhnmuTuFW/uwybcp+yWomuztDT+
1fZiT7E6n8qcdY8xoC3zerl9OuX+Ba7/Df1Tl4mwkwdmiaCXcdxtIHpkzFkQcObNmL19kX2Gb0jP
7HYFacohAjoeexzxFmv0SYgalvP6l1WZDi3ncFS1jLIHs6Wu4Bnr4yLzHTnTPOfybPsOxSzniC8U
NA9lpySnh96bgRZFFVcQQp6+4tenyauubx9hzg/RuYp6Q4EH4ZBVZ9R+8h8UOfTPGK+0nOWHMfZB
gEHINaW8Ff36wP55e9q1ewrASg8T9cHK8Hx6eMHEOEfHm6mS1LBJez2k9t0Q/HQ9ejfUdrZRfs58
DD63aH/wvlbHKzRrkmvw1MrBKAKFbTHjnolENtYS+IFT2Thv09FEADscOt5aBIsAtsw3Vwxf7W4P
v3Zaa1p7FK0ZcOE/CXIiZ0rietFp2w5qQUUpLmU1TfucmCmoILsCwp7lXo/UNpIuAmzQoFwl2zwt
++AN2MDfLRr5R+nxreoAuq5ni86sUHLPj1ZjIz7q6ANMSBuK7wuXOfk8+GExcH/7WOi4LOwcLDNl
ZnSn4oZbTuASuZhDmFC5U3tloWEvPQwPEiqflFg1DaRny6UY9LtQmNTy4AN3DXsVgF0SrA6lp8/f
LaifuOgYuwcjHcPUOiaYCbzR6PQl6nZ65RF+tFnjBtlEfdQNFLQUK+nFKm9o4Jhna/zJI4NaMcsm
sD6Hpl3ygX7cDpLaZCqNVp4rP/V4nAEac0y0u0jQEPuDP+ovozOPyfAhg1wNEKxlorpeHGi/WEIw
RuXo6v/nLaCJwAtA2M21+RvuAfK6qHyYP9TiscdhLxlS9eE5H4oCWtGh28BBEUPdsde/1Ho7Grwa
9+MWQlUuF0H9T1t/WuaVXu+jVCSwqQ6TJdqW9h9I2cc3rEyvqQg4FXYaBCwh7iIp90/2kdcskd0K
XNjiQ6Id4p2MKVh24anHSsej1aWHm2WXDlqw6qJ9b2a6N4khBnsP9YhamemUhjnUU0K3BYgrxlDl
7OjhwDUQhhUWFkKgMCyWWJTyEibyJkz18ublhBXzRh7YBTRXSECZ2HNqWP6KVLdi5LnmfDZiIquF
1bgESA140+O7pClon4FGDmEhZQq4bYAIS8e9XAYUNI+ibLY8nT+8WN/Ou3Re/o76+0zsGd5hlLTT
nMbsPAAuG53GWv5vhxljsmBQLS+yJlyAZbgMLHmjnE+tqbalQfokbv60mKyREa1HAo8nom0RSs2b
1yRvItd9B1qcNuDHEDwtinY9TCq43JpBPCN3X4juqk1mW18qmfuxYLuq0dfPSt0XHlu6D7zm9SP0
5xTu9XLFoQCRetXNv8+qFun58TIsh5+CCMggJxI6Xvs6Gmd12qHsEGvRdtPOvr7KTYpIeDoIidrM
4FtxtuVKabn0l+bJLXSrfLPBL2N22XlyRotGX7bnm9AOrbryXeJRJ1A7M8V/8RqP7a9a0k6N5SnW
T83MkZ9rCZio9zfJ4/ekLWyuspati+bM6Ogjn1ilZSQBbf2f2kjJSCpkWkdJt7NHuONTEWrftT0h
3x4m4ufN48+EDMpAZ79MIZRaKvOPrcCSbNOp1TRIyetC7SkhZeRoNo0uayd3L4vhLa46S2MRROlf
EZAb7N0BaCoMeasxCh8oJte9JtfEQQ5E62E/qMle3AN9R6Di9JY+9/g0MNFjrqrV0huH43d7Sesr
qOO77Fdl0VH3dDr+rl52Dqpuw8GE5CA3rYo4kOb5te0ptC9sOWVapbrriyVzhdJfylYSr0CNxgNx
MQuHMXiCDWPYU7qa87cNMfYq+OS9k1NeTgz4PInrbOODTAHVMWWh2nmQJUWhbA8x3RbjxR+xyhxb
Pra1EVz3EYa60RPLjcfUqIQPf8VrhVKMhPuBK7uw6gr7B0O2QMzbcXv5W6HiXLdApM30BRV6Ef+e
C81T8YRrfz8GnN38a1EFvkihA2rilIyZsKRAbSiIbTlPKe8T4HANUqHOj9m4Hl8k/CI+a2TJUwqg
c+1nDb8CdqhoFlBSkioJfuv+2lqAUehUIG6YjGL3boQg+fKSeV4Y29F4fiJG8DvamZOuDRd98AE4
+8QAKwN4XdKIghXJF775wucLW//3IbtqlPUaVVZKg8w+Wru4SvSV2k/m5A6A4t5V9Z0iHAUELxSv
3wd0ipFGxTrEPrQKpz0E2AS50qatUj8tmuAve0SoFcEZ2u9VSRbFlBnb7dlIHibLawN0cP99Jlrx
7j3v2z6qWTu0GLlShXbQC7J2MWhqg6Prq6mk/DjUq1liWlTtCJ546GMhyp141aIzWjINteIX1WNK
9dZ9pvrUpZbnFzkTrV239Ge5EA4PjW31clTSFkSMwnT6z7otZ9HKwXvKE5S/OR6QVYHWitKxdcme
XxlDGp6jkCjBlRztFWPLqQl3QZvW+ftb0zTzT2WY65ixaDvIIbOTfGNMHUvC9zdrUN2gciIWvDty
aQvZcs/MRP4xvVIb0l8lsWDqHOEoXb3f/vvXP6mqtV/NZn2p+BC78qNrsQjWcZZqDCeGiYxXFBbD
6pG7eZfbfquHLKzy+7TvKFeBH4wSTI99nQrllG/k+8WLTxF39EHQkdUB7rpBCct2udGT68nC3CZg
fojdorVOeg2nTWhdftNHh1mJj9ad/BAckJR0x3Zcl0ckOb3Q/mEO8Q1e3lckrQ05uvnBzbjkpgPC
ZQWa0YNNAPi64X3Rx6/E03tzRsLZEcDfOMP9HuCnxO8Ho2bxjc4eSTIbTJWs/y1AiCRcyQOop+9o
pmLS3CKcyDmfce6A1mg8Mvg7Ro68tTCoz5cWKGrdAmMK4DAo1SGGG8q14sraw1yyNbToqBW9lRq1
O5lTfNDhUyzW2yfJJl7Mi4tEdpYgNwcXA4pyw1W6pBiwms7PQNg0MkRbFWv1xnOzapeN/SmxqIQW
dns0fxqoA3IN/xQX/gRaKuIKcugVKDoexj8PeRePZkWF4cSTWnBYu+Ssl4kncUw1qcUeTcW5eT3H
xfX9hIfOd7f/+aMDTgTILaF32+2Z7wZhWDHW+XuM/+vHiRhV3svQHbcOJg12DIfrydbw4xbTc36V
7JMhqO4qXaj/zJOrXDsjIOFiB/m2jIyNf3AQCpnwnydL3lNZqoOVM4ZxZufEdePrRu/ZW7mVN12i
Q6T0QFqCx1MLlr2h4WRN9Ju2om7t4/nwM2mUP2ChWvrI7q6vkHguzR+Y3eWzME2VmIG9OzXzPnpJ
DgUMxggmQflxUzY+lCR7hz2zRLVNaQCpX0v4QQrHwlH+Dhlm40nEwCKsvdUQY2ntNtVrmGPBQ9HE
dJ6zpx7yDGddE64yJ5q0tezhcygp8bv0Ib9rcBZoqSikuZWoQpD8SrubxBgr/dX+Zsx1pnVDX20z
LvIj93SUp/Q8pcsvmgvA0S0alS1tJM2g/mMMfHeC7BLEXMcmvdp5HS7pY+NRbU09P1tnqjkYD5TV
UBYSyWFBJKW9OYYz6lOJblME5LXCP0XMqYnu+oC8WEaw16gcMEmYQUgymWkHuqO9XtYf1K8TGknz
rmBWrVaoyl9EUmWnwmMhRZi4iQu+k/q7EUF5Hy3fCNhLjt3hy5RxwglcuNMSZo84a5L6R9WVe1u3
OhGhMHOfXdwW5rn8th43wnLZ40YzROUqF9gR900IbHAJKCAYXVNmq1q17Tzn3Sg5e7dp8wN6kBEc
3v+z1R1n4AHe/8APeRyzQdnfA/40KkapZ2fWwtzp7OkuDhezeytJ2wJ/fEVjiGlXN7as/supNTS6
43de2omt/PatOKV157mK4V4PAZY0JBvB5MJtA2DBJAT2zg3Z5cUymSarJ+KlEOOGEdT+zU5FlyST
A7GhTNnsti3yLgzvjSh0A5CQD27VhNQ18w+yCqr8yyIDH2vvOdSMOCPfRTi1uM5KXAtnNgwG/wCK
qDolbNsabMqaeT/C6Z8v/Eww5Iino9+RAh6S+buql4YC5gCGwj8eqviVJDUuQnlS4RSohzH5opc/
GbqgS+PFRkgw/WzclBbVKG/c+OJj6VwvFAvJvsmyH6CGnTJicruTJDL/GgWSpDw5DLKSbOQ4erw0
zhLmqWf0DwSfj2JFtAiD7rMfdAqX8Qp65H8voWNfSKb0jbuOFPvCyFmM0ZD1wPXM/2LsokCbl2NR
jUM7hy+A3DH0jWa6BhejY8H/adMuHA7ZaPjwveX2eAx5rojAop0ahpLnWmsb2uWnFio08a38FO0v
uA6Q0L/4Gnt2p7sooOhCYFz83YUVFzEp1lfc1pkgLfJwL2J3Cd1VOsBXPXX1WIBShKnkPHXYOFZG
plXsri82sunM680cninkYWGDORv2DxUFwZ97gC8oYsDjLKgei2EE4Negzjl9FSATNbwv5jrsswiW
2siGAEte2iEYJRJQrO7CVYV1kOYaHYuMkMNXmfRyhW6RI4FybCM8A6MohdIsCDpofZAuC4MJPdZz
wBZV+sq8tEcBq6GkWLzXjJjSnefZywfLuBqYCHWfNwh0+T9bC2NORKEWpywq1SLJhxB7gDBRqhF0
Vwsu9vp0u/eEFVD8AzcqkWDs2XFUx0OAoZR7m/5qW3AUqQ5QHuHDRDc2U4BCABIcsl5NAABZx7o1
diSeN669jHO23ps3jm1NHjeshqKPRV3XU0hipCQlLwGz/wCKoS/B4YMqsXxW0y6qh+YrS/sb9MPz
jARZQqCtS21jtMKpEvHTIp0AYjkgKV+DEHEhCxii6KR3vYBmzvakGWCUg3kfm4rVPvhiZPcO/5D6
Cytr7/ZMVtK5HI73gRcxUrOllvH7h+6tZtu7ySYY4Tyzd9YyucRYLtY/wx1szBUO3Ju1JDyN/3Jm
JhKdy0AYh3+G+vWLSjBlGZwWJULSTEBiGwBy4JUjTNoJQnpoTWd9cJvEczFb01+vMS7KjvFBMiSR
nXnR3tMEbz8pleGm6V5u+PPvhNSvyETbBIheDNSB0xvzwJiLoC6kAJoi/dntMrnQqYSA0LCpzm40
0w9MVbGiXK3yg3maBGqC8mMvAENae7tR0fbi51o1tG0MoOT4iiHAIebnQwsf1uPxpLEaaV3zlywS
9iSqsmnyqXOU8terszvvutp1oroxxiZDo4qmMfdWkzctRH3ahfYSmuvRrdqEhDOUSh9ncbxxDxP7
CvZt+LWn+kIa/bTtN+vcp6uygb/xRLO+MQmfp/8Y+g4BRMADQfDlgKi/73KEYSkQ7dn7oS5HPpzM
IjWTZ2WLTiwccp8X6Q1BZsSjFGZvKXPElTw+iQkQZm3FN6YmYDu9ZZfXr1doMcEHOO7lplH1bhRI
D2DEo9iZF4j2kZgI50YKnijGKK5QOemnKFoWaGDgobettzDBY2DKrNlQOZirrxo8EPUcYNcWF1Lr
ziy1gduX5z+21kf9icW4Br10xWOlDb+RibbpfQF4Pd1rCSE6HOXHquEB7rmiwQBbsDFLTOfY86q0
iF/wvNLvHlOwSqDpEsiSBWOZGf9LI3ec9k63i+iTBFyfI70/2cLPKJeunl/hV8/rgZ62ZwqzJoRY
RtQnonreGfiDMy83icV0MWQcNp9I3qgCSPgO82Ve9TJj6z1LMoWHoJX9LImwSB+eTgTy2b2jVnbN
pfZhTqYdLgTt+LggtbO6uM0o8IVDvCx4FwUAT0nTs/v+8D4x8vZRx67yxS9mgTx8OthSj0QrPdCK
bmsnuGZbXho2aoL5UuFR/QN/d9SOjxWEqtV4u4mzlokxpG1kDswwm+K+z97lF8YKJfNmk6vujrO3
yEWAuL4NQjzAhG/A2ChekUiTwtZrHyn30wf67dDj7AHxpsvDdF3uNgbUII8UhV6L4SWTPv3s5ke3
ujc4cIVXXiGbyt5AZLkc7CDmaj/HI/hKuY44ODU5J43gA4c1VRIKlXI6rDKmUVWsIiCsq0OXC1lQ
Lwj8+DpT/KZUntK20evzk9OlZse5mvml7CbDbg7Mss7mYSNlG2uDowxuNAg1y5Wl86KCzLwwWtQg
fLUHygSlF+mnxv108SLMQRuatUtxeXre+a2SOxgG2BKdgHqQzmCdLATEXUxp0lxZ+Yuj6xkOQ4fL
dE3aEYYPKgOp8N5eK8DtsZ/eNixf4GI/u50Bfa1HW5UjDOumZi5xUQuRX8YzSA4O4MyR1ocMHDrK
V3YBlMkzdLsQVRlM79b4TyZIeokNhlCVTDN80xlM0zSll2cIdJxLpgGnaogObS4LU32+32sNlTxu
8xmxJlCTnqUFKDzglS7yY/LZbCyzQmv447FdzHRXWOfzn7xKTJ/kNQ5TVpthwqavPDOuLN3H5Go0
B+w853eD9kpUG+Ti5BIKsT3U6XrMwwvZScdtF9Kmd4DihEEsgu7bQuITf4RvwrWq9ur1uVOjxTDG
X7CxejAGNpr2Bh7/mkPQaJeTLz8Cn+NhS7/9CSdyOqqeGExuzxSFXWcQViz6IrIZcs6REvQdF5vi
wBNyOxw4lM4AheftNq+aIPpH0uW0fhq4UeDeSkjI2kQQh4oaMnrY3GX+Oe+Z3Hpb45jzchkWVQZ5
P7wQnn6D0ZydVksGh2a1L5jxQFsj4f3Kv6zDjza/ligrho6353IuLYJGbx5nV14sXy/2MR/3hDK2
zeNUhttUCU1HZD1n1uVlBFvaDev7C9HJNJFytTnDiQw9gaRdKercg0XVnKI7SitRhB4h1qs3SIXD
022JWjyehLG/jHxrqdDYnsGxCW9qjLsxl/Axv0J3r5eMvamuIW4sMLFqhq1vvwA8IMFjZMDfgd/o
et6fEc69UBT4yFidr/V1yxgR2Zvr/G4LOVkDkFrsP8PZ1kMwWRSbM5WwwjD2Wjeni+EaNQy43hSR
jlu2YhwlZ0z+ZEntLatJMfK4JAJLF+JnGbBAyS/I5+KfBO4boQNh2CsslDTuWlisNuOXx9hGr1cU
xRyycdAwpbu1jTXnHx2kBUp67LFtrNLh/ScXpbWxrAc7X+2iR9K3ML9xSL6C+4NFyQNBLlM2J1OQ
FdPkncynnMsXb8nSAcIKyrTZpeqiZcR1ux8DWidU7GmQ2qIY/BisUJWh0zRUkaZJSyxiq90rE6Mi
13sBrp8PnhlPPOiTD1SM0NVjfk4MmrRg42JzVZdK/1ZEt4X7GuV2yMEs2bGTopftzkXRmH9SjB3P
zvNGhu1fDBrQ95h3C02Rdyzcrz7yzhpLyckIaL/lNg/DEL3KdKx88REemLuqAm9bt+8jGjxpfAsk
2tVSAHMz5ESQNhU5w6rqF5qN7+m35dZnC8eOLK3u1BiJKLdrrVL4ElW+NJ8TRpZzZ8B30zVnl7Jx
T6AVCX/uV2Bz8RF6v9x75evm6RsAiQQzicqqZTFdr3DieWZ/dkSWntkt/aZ9BRjMF9XJEqAOu4/P
7tb57T4T8X/JFRhZNEio8UATGj82JwIRzSzDSX5xM+U/s7Xfh/b64XDje/1ZzKyKNcTT/sQ7WwAy
E0BZ+fGsbUlLwTX2hucmT6Jg5QGizlWtT2ygl5O9XyVHvFHpztgLhFDH28ygQ5Gsiz3JY7ppjYtt
THJIVGOE85oQPFuUT9R6R5xomlp90a598qsfUo+s5EuwclIyq7r7KFxWXKBxwXumUwTqk7ffPoa9
vByb4eZMaEeisDXlaeZAMPWUupSELYdsTBowCnUFNCaw3UrnWZmUv6VhzypG0kalqnJ4AsGF1T4q
pUOnPrKTZZQrxhsXWL3xzt85m4qJpD/hVcMzgd9Vn/IMwPmymd9qMCfGJ0xhVf1UrZOu1KUqTwwm
WI3JBGkq1QxyQ66FLGVuqnrv0sVR0aneBfrLT1JT6GebTy0EDzPKxl7fpYKLsR4L4dpjeARKjmu2
GAPtmULCYz542W03H/RctuGPIrD2H19J4p6vRq/FjbnYysuXJ8aKXbQ/2r6y3zhGz65NJPEKv2WA
MMvVLlGF6M+8skwzoSi66Ad0zfQpGyxTXmD8/on4gy2EEohdzrGZ+LISwUhTVWgD5s21CjAZbW5P
Cza6CIVbBcrCD25JvQr1g5qRWAPxs6RU4K0uLRZ0dvEf0+dgcUkJyCRfftfKhEdcG6w0Fp1NJUbL
QkKiLv5wx8G7KvBeQwOj3XmgYL8eusJWYg9inTjAEJaFgoSKR1uwKHnNqwnAitcfsBAaDNeO/z+Q
v6BJHhbWheoB60GssXIJSt5ncktpViuZLDH4XdhD7DvIkuyH/sHWR8mCSsYue9+73BZxarlLaLcC
r+vale/rg7X2aiqXC+a1y6tbYQE4GAkDPshOBGz9PIsuMKWk2R9Y1ejGFSvf4nNQq8Dx2BmABE+C
QlwkTtzkVQ/v+FS0xxcbAUeBGUHu6BdS2ChyPjeT7rvweBjK09Se49s4xt3AJFS3rufjkgiups6w
6yqIydx3Xufzg/7qZRfs5moDxAtg8+Kvi06SvOVBpxFMAR/Vt0Y+JFIwipB7qMKS8AsOGis4tcF9
vOQ4v9sDoP0J6pwSDEiS3U+O66WWqhlipZ866IscCdOAuatyEcUW7aKnSTZeWwlThnyV2P1DWMx+
nIOOzvfKurTzXx7z+F4xj6QRHTD41sSsqkMEi5j95ZS4ndTpDiIRXC0UdqgGPbCNf02XGSHS0aZm
ytpAMGVyJ4XbZwH6NW1rmDa854ZC+J1DhUNgifl/+CwCAAmVkvFqhnFZ2kCJ2e8oNgLyDVYthB5u
L9rUeA+OkDTLJW12R944WVVI2gyUWfykH1LixL7u2CWZzGILbGzIXMxPPJ4ZR8yPlpdMN30urBKd
NwuJEzMok1J5jyCjwD0hNdk1n2AIKnd2POQ76F3LAslEvjOtcQRQtIjoDhNCydnJsNQQc9KBYmlp
aXmuhC3rx68XlLzRGmSh0D6M/vCdVrugp0+qcGhV3ANkviuVhfKpREi/zGEBEPuXTRi8BvnVTeGM
W9gPN2jgo7bHApmXc56JRmgTx63VQyNkPVrXI6Pb81y71y/Hrv/MZciQ/Pogsk33RJE6m0/W3Rt1
Kl62z/ZQj8xVdaa14qw1i28rcgjkR9P/n1XioP3u7UgRKg9XDHut/EIm0vYAOG5+U+ylNJQtyNYs
2sK17pQsg1nn8C+RNYaoLMxWWnsy0yH+Gn03K+Yd/NUcJd8GCb2tj6HZERdUQ1CuSM+OXTLPMwBy
a8FSxMwtxPQ8OKRSktle5QehC00H2oH6OoeAKaS3V+Wtc9uqXDr2viXHVrZPdJsg5sf7KqlbJC3F
9HUxiG6/XUnX2PSuZ2N7Ey1mB4hReeFDA4963qYX3AN2WxFDGKvQ1r91OIl4vvfAT+F/ubUA7BRh
RQ6UaXX8+eTVOHZ0oo2mmxtV3modQKH0+OIoGwTk20LlOh+Uedw/TRp5xp8X5Lv96lC7HxAwzYVC
EIx1lq5LoVP0dtzql/ZAg/okANUNNak+BKOn/XvZXkgN/Mj9zCrvUF2NYF4fJqYUXSRN9Xpwlz6W
oY7sclCorvnuhXa7vMWsQ83zyMHTGlCyDTA/Aj7BvKXKWdQTU96vgPT4+SI5LT0orEVRb872P9oQ
VT7iiKEZo23tXkKO7m18uhjhjaHoFaJImD0G52xAbKQDjbrtOdJxi2Klbr2OlsKSqGpopECShKva
bqYV3t49MEKCkKfncdibDBPSWnhsFOpKcRt3P/QgxgeVoMaPRT6U5GXCFmaNfR57SqBpP6HFYdIq
X5WZgfW3uuWhZuDzjF1mVMQl9T5+WmTNNqkuFRu9vk035anfvKyyXZGj9guZNT4cwrZ/kNWWIzVY
arY+ZvBwbaKtlQDau1Iu62xmYraP5jiiBuLsBOxYsRP63CPsS3bqQbG3w0/BA1RKsw44H44IwANO
T+u5qcmw89WRpctD+oF0p2pEGoX8eBSf/LvaXjdwUdQGkWbN3Ckq5WRZaX1NIFb8iWFkgJ+bSRGo
10Opsjn2V/XG/nvPkc9/w9Wt2EbFQta5QYWHJN95EEAbtoq2xoCm0xmJuWec4tjC/rHmEAk8WPcu
onWoTehj9m+w9XOKV9TOXwo3SxD/xlsN1j31Y0WLjdlKMDvhlH5y9Zv81mqW/5xrtyUq1F6WlEVP
jixiFRz6Lxc2GlqMHWq2B/1ovFAlKtDbKOhgQawrcTCQG0O6KmhQzQYta5woXAAhQXZeM4cBJyGu
Q+eUyyYjWgjAD6chc8X1pyDf9PZ4d0J11D9+M1In+6UwyNzZudncJxh6LPCrNt1W4Bv8X2CeFrnB
ZIXfoLR9fKMFjl3dD1uNaTHDKsqku5OU1TGUPnfldrqOluWyQGYEeSF86+ELsFcZ+JaZ1P6Yun7f
8fAnomaCiAjHhCBvXhdqwpUUTl/cw7/HMTQtb4bOAONPtr/gcn61fxWah6i7zUoE9LVeKDoB4zbF
aLR/Huz9m0SWtF5GXWuMgZt7/UL+p1NcVjwmosNmgYpsbsM4LJ3vzEJxDKnmmQ99d2OMbEW+/5eL
Ag9kB82mWQ/qZwZs8NqkVf5VB/JFiELttT30/y1cTS44hFvrZ/QGeJnoKjOZ3nFvJVdrseWAatu3
EJv/p9OEDRc5Cr020pPd3dH/jF/43MbaLXzpuZcfqBVcQexgjLMSVAsyuvuKyglp3VkUIHwsVoDz
/IlhV36D8p1vC+TY1gdTPZfG57iWeutHKicrVly8I9PFd10Og6ldPoMF0Iv7C3p2UyTp7qYqDJ28
Rkz1weeeLSihPQ/87oRzyTprdKjuSykpNJrxboybGHW/tHxotgo8QUW9ai4BN7yt8vNoMc8icQEV
FlRvaKEtHqrCxyXq0FEoNywJeJTHrpBqUQ1FS4H1J2Zq5jxeTWMmIXnJViU6GH+NF5M8o2AX4thk
0p8BrdEMYshNCpdISg9CLAjnq1li+FE6r6Xa0YUezB5Nl5YrIkylMWCE4e9rbWBSTialShIdM/yQ
QwzEn5kitFZMJ+kAyLdvdlqkbT1qJAXHjDRGQekZpQpnQeiDqG3Rjikem00cEjiayjX3OPdNV7+x
QrQlD1xrH+9GN2EcJC51vBg94H4ze3xArQo+gAAuf13dJi7NLarsocZKf+uaX4LLqxj+Y5EPERpx
PGXWwsBevEteWM5HfhKV8te7SGgAS9fDU3q+BfqZjQTwJKaNW+Yp9OCY05LtUZ+zTmsL/EnT/ASy
0OQTeh4gmAUPyYuU5XmNz4WrlWcccDQ6DKxga3Yx7OFr/bOkByL4TVWWX5IfTQEvBXSoqOzZOQLR
FDYAmSA8rZNThQliw5nkn/GVq+87pJQYfv5esYwSv7dF4yT7C9/pEZmkZKIdlXNLDouIe9KATGtp
mmoCCzrSUjcxLbFA8gCT1U98+xfaxAzi4So8OYlX1yxPY36NQrqfl9jC1SDJ+8i1dT5HCg2eHXgl
7FsHl43dlg5fJ4MGtZZMujgNTAJx20tLZrLNALHF+UVcKHEE7UeE40jPK3ZWVndhoV4nlEUN9P0x
T4PlOr47c1bnHT/kIpVwBjQYoY5+FHMiEHUxTWFXTVkIOdY2tu6hpcxclVNMRtP2XSDdSrLb42HW
eG+MVu13EYCLZvJ5xG24Z869OrwB7hmesaVVJRhKYrcWmi2/zS/LmZGDccSWJ6E9w1QNLc3Yf8FS
Vtf8dikTb+9X0OqgivBG8nq/jKwMsgLIt0Se59K+eEDPKp10193K1dph7jVMQwUKKQQqb79yCG2/
ahXItbYvAx3cpVP509cMiU5zYcq+6elwXrpR0NWOsM6WHKXNf53In7BMpNPuDUU8yaLYjWEzJRPr
H34MPzQqBHEP7RchQLHGvt1PWhb8bYcw2SrvHLIwEcLAfKjd/gw9HhMvlH694lUyzDwPgBKeD2mn
Bc3/n2+fAH1eL8qEXNVLuCOWo3pOiLZEKxwcBmh0mEuozzzAPP8tTifJpf6OL28CPC063wFJAsGd
xWz1rmoU+6GBuUCHjBpTNc4v6om4auDu5mx7uNIN9Uv5K1cyBOJsqugr89jyiv4ZiPoTKRDbaStU
H13sPipsYFQz/ClYm2qYrrak4o5u4+ACoSQjPXZ/qcUK5uby07z3fHMwntkFI+RKMZjcLbRw+kGM
xlqrtc9NsqvQiVR1HqOzftDnRs/zJ4z2schsF4vv4MQHOEQ4pNt5fKpzevaA1J3DNVzwaKsr9d5X
o5fFiymcHNclR6zV1RJH0LqxeJqrtsWlVkKmm6CO78MRPF9Z6rxStOMkQTPfQxHen/+VEGfJpBsC
yBOoTgrOXaYkASxbdy9hbAlXBKIqRBnpIYiTSfui9DGQc6e2+Fauw4aSntDMb8zhYRhIji+fPO69
1ogk/xWqkq7jSH7VV3D9d9nhY0q7ShEuY7W554wseeGwLdvGf/IbqE+vBYd/zx6UU0G3N019g0Mw
Rx+a56zDjpxSrsZ2pJzcfLhkEiB/iCxCLqeL16DnhqNCLipzjWzb0hsR0o+WMB3alkURdnUjdT6Z
LLIc6dcYQ8RQrNGtPvalPCyzhR4ysC7hwB5QHkTVpnLhLk8HVBSEL1XJEtGg/UCMWRfrUUdlaHaa
wxokA1rvBPm8h/7L/37THuxoU0yOAORG4t78cZz5AqYIEbxOSkv7fSYDsZeap8OTUYFo5b7Ok9GH
Tu/rm9odqkjroRUmF8QuVsHCKjMYbT2UEX/ApqC/WxRqT+/d9UXXvm6enPJKs8YiUvHNKuJol7Zm
q8t9pDyYh3kNhjCDm/d64bH5COork2cCx3KpQNG1nwxAepdtuB4w6m4b6wpfr2cU8Gu+A2UWSY1M
M06bcivSXOZr9kHohE2hEVnPMcKHZfNlAk9WDvP6gZpj4MJOvExIWKBy5ZdUDAsRy3oC93Ji0BMX
eXqPJHKI4g98SuPJwYPndxO31VhTe1MHMvaxYNymeqY/6R+mZ9FBXL36QjbG3D+m2hCMt7LhATe/
zak3CpHWHBnfeeOKxRYG5P5j2rmQYEpm4BSu1NAXvdvuiFhy1RedGgRC+HVdSQ54vU2N/QzK6nrv
DqH/o281XxNroGAYkhqTYh4rXcSQ7vOdjfu9b0bm+0/C7Bxjl0+pD7sAZe4W2p/UaD1yYxKS0xzu
+L9UazGtldV0eHci0TxcUkNxm+M68o6OrVZhCcXHipzdnqC5Yn6PFhtfV5ZBzIKck5hYrhYHdytN
ojVIwMIP0lruhd7IAOKdgYVsB6da/zENAV/09ycLrA9wk8/J+cYLyMbKOApjhwi1m4wMJ6p6VHhZ
e7eT0GN+jgRE1kwdJmayqZ/2Ee0ADX8rv/l93/EVD0GkJIBitU1mkFm/hjlVmme5Mf+0DmvF2byy
2OtRMAHYsDAfnyfUXWp+YMqGPo1YWBcRh8OlC2EUERX4uV+aFj4cPHi/94+djDzxZmeLchk5z8p/
bSCxDeUuQNQuq6QFqBTpyLO5djI/koSszOJhdBFfPGttnbDJuZZg1/IwuRUrokka91DwI/7MiLhw
yuL1x5w7+Qqyq8XtpcCxy/rXzU4nbxWw/IS9cFmfpVq12CxBej91ytH2QI8kDhT5epZPU3nC64Rh
QcFFXq184ejQYPRYYGoaVwL1NeQcNdoypHp7Yknxb/y1k+wALStnvvb/yKl1RkNScFSbOiMTyAsc
PE5wqaRv9ttzPmhvyJ1lrhFzQujdYQa8X2unodS9DB3qCDTB8ElhgKFXfPm8x8c0m0QX3gEj69W7
uyO55MJacAI3nM9HyBLWWFSKiwbokX6lTSAER19FK7TQAb29NyNZZFHLcS9e+VTgELRyTeXgPfHb
m1Z5+XDX+TMmCoGgySr0EHET38VxZiWjQGs4h4+JlNyXN301sSb1bo5MYtScMZhmAd0bj4tBnvb5
NJ8hjkXzDlufClsf1MYInRvdlo0YwqAa4WK3adf2yw4qn3KBRkfD+4szBWv4hi2oFi53I20tYb+6
HPhZgWZVynd0lGY2sS0a00Uag0HlBPlzkYUS8fM+lVLAZWHri6ajSiyN2DCQjLMzuJ7OsujSl/7q
ll8N0obWdbKc1QLaeOsvJowpfZeFeqeo7bj8v6EokT+8TLnupFiatsqroemk1QElFeXoaw503TkH
U8ApuFu7J1aPBw6ezMftQWfncTjZg4KpRq1H4a83TO1Y9QLmdwz+LRUU7OIb+8US7YOV9oJMAUsY
RH2KpxclLE1PXiRcBmbwhf31cg9t2Q/lVTenip6wEnKNeIaHYY1oZGg+eZlGwlBEIm6pN8wGMeRX
ynuvSB6UUZJhAI1X1deySMWLa+0yFCU+gQ7D4FX1MA6Zuvq65A//fjssj5XV1xg4J5qRGTZEkI4z
xtRKi/HOU3v4I87Feq3KSrsOumH6oXqSkOjt8y5m19HZe9wwfKnSykUx/eoSq+Mb/nWbFTZp5HXQ
vGxfPnqHXif405OUXQUil2uozQIwiYQMj3An2rKgucAZ0shL38EMzUfxh27oUrvaDSSaDPe42xFO
UadYINa293IzpeyGM2TZER8x82OM6juZFc6q3VqD7OUozrd2VPxmKcM2MlZ5T8ML/XxToaxkQewv
euAAxr4FXmEc5fEmtdFSliQ/dXbhEpBPSl239L/xs4aDIfKc55YCF945rbptLCev/hdN0OnPD061
k6GRMnxa6n54gJe433UbRm2VV00jKxKqQqsCr5HDnwglVWehh+vr6i1D+ejcAByxOae9nEwzyo5o
96gsztVi1FxEmoDal+C8TgIY9xMoPZw1ZCx6HNqpMEtnuxSExsOWXZPjMqPRIgeGP/TTPSzA0i0V
eVKabyASBgdrgMugOWzpZxTlXjfqKm5BlbrnBfy7/N4cf82ps0788nAkYkWh/GsltROR1eO3Oevz
lwqC8lmPocHRE93Xm/sBk1YSyK4hkYXJaJLoggcUCr6Xj9vVcWScfkQriSIdoHvwp+HTldojzDUP
Ki5Cfv2O8hVTxpcVwwpT95a5JuOsVtSoclapSUnw8wW5AHmelWeahg3K7Wv4VE107Xj2zu3X4c0E
gpqHBoxS050cTc+ffPoQXmrd7VKFno8nB37D0thw+/UyBpmVMjdZ2mcwTv+IHDzBeDHi918qbm3c
IG/uEp/KR2PaZW90Bru6JXmzvs2Bm6HXxBIEiQ4DP6sZUsXnBgKcW8mYZTddQZPb48bI6bs0QIR/
8ydJDLHZTHCcLsOAqEa29DrQYGr6tEWVver3Z0hSHCfYy23GSwFZBkxMP7W3CauJuneXj7JFzH6U
xCAqulO01UAhtkOPyO8P7UAAQvjvCXHj9dwGGbkoMkzVNtat0W7K2AJpcaP3nupZKjfUSWS/5/fZ
uFOjSqTgnhZs+BctQ2JDDR2Wa4OX+AMtSq/QQq+ntn2OrrEW7BS374taMh7XdGf1twqdkD/hYzbu
Unlalb3SwSKLBDWjjyzkMxNKX3MJaxb18y+LOv5CsToGQ88tpoASU+Vtde78FYfuHUsFhGf8sg59
cgeMqkqBlY26xbrA3kYLiiEsbDgCdt0NW/rriuPbGt4rQuAhV7WAlJN11w3nOyVPhKlIAVCxCYV7
3nVMW2QxXbz0HOSgUMUS91BJ2nTPEO4x1AFe5RF4hngWLO4DR0WXfj0JDvw0v/0CBe0e3wBkO0Wq
GYgbyURoevoMRiacuvmAi8/tcTwtMkKAdCkdARaD5vRw/uhL6Pal441dP02fE9Im9dQ4/FVzOfCu
Gd7zsLf5i3l02fqFOCKYIbLFUyxNTo07F3Fk28EelOWYQ0mpLRA3U6y3WQi6wl4uvtufOjWKEbkr
skINI+FCttI4M/Apqw5a63kJscxeFgfIQpJtelgR8llyy19mcuFP2fGrT1BmSHwuYtobysAlmc7/
ibrRpLtrNOLA2sDMxD64pzc0EuMWJ01V21t7v9vUKHCROsiJEKR8+OH8uOebm+C1f+p/UlRyYd2e
kGWPnCKtiilrSsHfbzBi0DXPORVfso7nW2zE5xabqg9hcdIMKSFSguKbQVNHe0sQNKvRR+vtBhFp
cjjSgc0Ls5Hi1+PdjAhRyOFDo4Cn5qrKqX+cYiYIDiqmMbA7ObRh5QUjNE0sGgFSL1Zhyb3RrB3N
LPVglW1n8GbvFDVQtxn6rvBq97oIYdzJfA+3J9/loKXeudde22bVSIK7MUzTjGJaKmG4oxQBtHjz
tTDiapUc6teNTG6TujijxqW+4HnNSzBAeSLD0iFU2loHSmsZv93QeU4DmARJgLDurbfgCL3Pv0uI
dqCFiPV3qqaixBpEYX+Wgf3qhWOcZMWtHCDH9buYCB1CsafpKF4fMNTGDviaGA2wV3JY6tYwrJmd
clX4PToKIcS4Kdzx/E/qHU+Yd9QVufAgA0G2My9Xy2RNgloRKUGxuhvxbAHgLKPXCw89dme+ddB8
kJURpq0ZJilhHtjPh8BQJmQSckmP4SIBAXt3Jv5+AcVTWYJby3ZYR3OLM9gc9wMtC7LEWjyadiZx
ibYYy1gpIihVhiqIrtXcxBt459X8bZQzDQiIjwdPtgpIYmnzwG1yq40WeaN+T+SVa/jLzEvgukp7
j6d5rQbbqt4HMIAVe9NBW71hKjMcTUB2xImzHcaU8wzhV71dmZLEOw2hJITJYJW9KE8nm+k//n0V
VgtM69eR+BQ7FpLR19oMZ0l1c/NdWsfLVGJkUsXFKuDiKpPybw8tP0VEW5wXFiZ69B+qJD+ClY9Z
js9MUfevQf2aUoM3/rO7CaugtZI6hotcacQAjQ25+NcPMc41MKtiQ03zcQKev62F9ZznEpdkEoiV
NJPmFQxUg2lhxNA+cGByUNpO4aJWcn96J4auLZCuOUL+u/WFP9kP6pSAIqATEaV4oXJMByEPfEdv
RkTz2YLpe0z8YaGdLt6SWpa0OYrC3xqdNwoFYGU2bgykuyqOi7CxET3YwZKSK608LQCVyWSokK4q
ghyMgSF1e7X46rDUt8zyor02EB89kbKPSvfUvpl9NkjwwkH576PbfR1hm/tCTyLmx9UZpo6s9wLH
fe8E/pD9r9JX4B9h6LOPjAwgRsahCx1sb3MxpUtRxnhRwpH3PbRZq7l54R1zwbJOvtvLyDYXXZUg
RnBuZpsDJQVPCDtW3Lxdz+5qSEoN6ZO2gCufZZZlWnNkCLylKiNeGVT37Z+MVDOqVWG1VplZh2hd
EFTdH5LJ0ZCz0lJB4a5BdEN7UkgGUrDJV7hNifrHmAmt7kECs4mG41cUZkEo4iWWM41WpZPpNkn8
+d9Kuwy3D6soiA6k9/zMkKQVlGPqm+lQcEK81H8HHluIP0S5hMnfUIQ2gN180tnMl8+bU1SY+HRR
Yu7e+ER0GZ2m6xmwIEcnJ0NlztVunCsuPaNa2w8DagjUdOdbxQxMdJ9KyYFknMz3Dhf969OHuM3M
i2s3AFCOUBWWtEBrQrZIo/44nWgJfEY81SKM/zJR/alMjuY80C5JKqwztZexqqIFiCZ3o3hxwSdY
2uU3FD+uybIYW5uVdO/DGfeEZGu4m1zhWilbPJre11qosjSeBvjjvOS9/zMnpUOIGeVRPGGW/1M8
1fptrxNSwaImFfvSCfLNzG+Rb3+Gm6tSIzbbkhKU+71l5MyWNS8Eyc9+LWaFB5mqfvWDn2SfyHH8
5LohCoBfNZCIWuu6jmYXKGEt0d0Mbrm7M6XwQYc5yiWAhHOxDqIsuSzT9hIEp5sG/+bztW+7eex9
3uBiTEC1FKPo4QZ/DTyiBjzX9AVdFnU/IYKVfMnp0/fhBYoUsYbu+9G3WM9bLXQHmY0YteAULtLI
th5XIM6tEUwD0yZUE4k/TfmCE8kHsGyMoQrmq2/9gUGdq06tZ9P02GHK4bSW13zyOgOKcBZPTj5l
dhjjzJBBxW5b4CtSMb4KIgVH98An/Bq3Pi1v0i4kIPuyzvJKVhVjEfBEUJ7abbgdS620MTcW1SFy
l0iB7VVitxOEzdGgmFzYUSFWvm6AN+prxst+nXrqrx7aUIVZ/BpKYVJ9B0CnuMV9lQNOFeO6iBdy
sAd82Ek86NEnN6TQAk7dGqF+L5SG0ijGE4QqHUGpVME3vqEzf4nMmBVzFkf7PQ4otVTIBs1syCgC
DKr8UWs6TPiMiYT0ln1ofruuN8kzjopt3NLrBQdrUaFa2MhBLSw9L60cjVWLa8+XHM2944rQFcnb
KgfbyGxOnVArwx5mgcc5R33MXFGo/lnjMcn91uEi8DXmy1ibgxw/C6TdgVKu8iKGmeDmC0xnMp6/
VeK5lOSBSclmZg03jjINRaFXT8/ValvhOqk3pFsVwqx/H7O8PlZBcmy3iq6yOXg0gqeIB1aT8CbF
Qy/QN6/WG4yazaIe3E/Nf74cVOOf57BYnXa3Lr84tb2KnHVDPUB2xW9nUpRDVNX2ksBgrcRw/nSO
j1zL1I0O2/kn/DE4PitrtNqKdCrzHOw0jJOex74oOlx7WEcTDV9nrlEbTo049gIKFaTkJEKAUuUh
e2E+m3F07E/viPXmSM06Ilr0Cq3UPxcfI28G7uU2/FJSLz+Zai7ge8tI0BquQ8H4o5n0i84VZa4e
XOuS2Fywi0RV5iASfiN8zdUTGDi+f2y74jGZftRjGWzRdHEA8m6EGKX7SSs+JJQB1cd/9DjY1xR5
9uO1cFo43yckZYNugSDxXk2CJxDKzvPy3pjk109PI0kauTmMYWdEngWo8XvHXXPDFzKl1Dan9zso
GnfwmLWHYd91VmkyBMpYUOJ3Qr5kcK3ZbaZ+DDaG8ie56bm3sbDBnNLaQ5zwmGgxsDy0x1xLveg1
C9gC3VdrA6JlS7kVg8wBCJJcJjxRxD6pRZUWBRMX9D2qN53SJKpviTXIMPuQkXvMXYX1+EUXnWGT
LrCGrVw6HZg8vCreJYYKOAtkcSXElgChNTfq9hyEvKW5AmDqmYHuLXrxxM9pzWRCF27fUkYagtW7
QhZZKOwjzjJzazUpfFxlqJH5ut6FEKXA6D89zAEKLwRdYY6zx6r89uWNsoEY4ufel9oI+AS/NYoS
uakqdtlfhHtNk7r8kokbKQAwKLZGYmEXUPOVXlCh+TV79zQ25dBIO+DNOMzFH/HRlCaemrFC6HUQ
MQCx30hLwxGMFcekc1M1Oj3Mcx22v2YZMvtdl+GSFdpRNxg8ftEqaU7SA6ATrPNAZXA8oSa+Yedj
+kMOQFdGY61Tbb+Q4WHSnRNQrl0UeOSN4CF9wTfklkJx21CJ2bsnAps4ghS4vZmaB32FZCklJNz5
tbP+qrpHKBsNP+xV/AztEymhINGVFx8nprSWmWyp3YS8edS9Cli1Ixes3VysAXn0QfMvJVYjecZx
wqRDdh1AULaLxusZdFhOlCyV9rLDhKL2lxe5T177Z2eixr00H5CGvAgJyMr2WIt7KSXLDxvrCNIW
naTgGai7463+OBY3sbkEoIYuZAOgoAlkiGg5bf906xTV4SyfksAW5j1BiY0aaenn42xh+PwrFBJh
Chy9anV4KAG8VY2SIPl+7q2hqejoDopwhSw/j105SNYId4V4LdiMmXQDLlcC7Fi+hb/PXlcq5gRn
tULaFSp1dOzJse/9bQWiu9JIreFu67WnRcwXszM8Aj6EZbA9JVdOo8ega+SOWpHw8GYUVlwiWaCJ
SiVlxKGtW/n/NTH78ihLzpnFNmMkNQA4xK0/fNlFjFrk+oSXQJUKC5q6IOpEcb0sIildz0qPsS2E
+B6tUL6TJ6jDgdkfJrqGOXSDqPWsUmEN0BwM+vd6k52YitfO3epcM57ZO6xZ5XQXokyk8uggO/Ed
MwpoeWfrLABLhN42hy0BVe3uAFERQ4FlJHlVSUmkE/fgE9Awg8DHbQRlFSloC9QxsmDthpnTH6X5
/IQgj3lEC95pks5b3P/WGRD7OaSltd/w1WX/Cd/TIlkj8cGCpPxcV8KKSeRlcNA2LzWb7IHzKSAg
rSqw74O3ugIKDnYn9r7fQ12GxhYhXPNGUgPxKUQNWxNy/gZ3Wc+kcvk9hs/VcJAPSnBCjO/I+ZVl
1z2LALzgl1wUS2VFD0DCXRzJX9xJkhv504vQk/mIMdzNUf5EAPlgOgyvk6KT1rGNzkD6d6th2uYe
0J7ZMo1WXpub7uNSiepC6aWNYOEsJvftVMfeptx/4qM1Rvms+R8MqwKt0+phut8vksLhBQDFpt98
v4X3E8d6zLc1DeZChqFCvt54w8FOADbbml6ys+lLV2lJFcOXCcCtNcsryKwZjJpr6kkhj3qDYf0X
UqxxybU+itHRsbuZGItqq/yrKRlXYIIx1EJiDJjePDspP7D/Mper5i1YVmU+/9b1ZAW2CUT0Fzvm
dew3V30gN5gskVW+3YprD4BPFXGAhqPM+PZjkLg0AHknx3Gw04IwBEr5X/K/S0J6h0ZbtSHSL9i9
i0pPsJyYE+SB0svrqT6Sur2OengsneEc9q7STJZSK41YhxYzbn25Jj6FJOKpkyyJwaVLv2iPtkGk
ZhcnvHqJ4g6RhSHuT146epvqtZw8ssFvykPm9iVV0x1JLYgBXapMU956gRDLFyUtRH4sy7rStuUq
SqmVEARhzBwOXauiHfXfZeRe2giLf1Pfs9puy5+QoRFJftXQGmp/RwK+8WGDOaRua16VvpbQ6r/D
q8Kcjd9Wvt0V6oENudjsajBJYnLuFtGI4+6dsKZXWWkGPgsvZvo4OVPj+fh6xj55dZtiCl0Htlr3
9A2r46U1lnmOiRnI/De7EWvkB4U9HUPCRkGw3L1Hxay5oUJB3V09WsoMDTVf+EXpIN8J/J03DDg4
m0/smeNw+ktjOCmnK3QApamG7AgbG0js6TdI8CLunyFd2Ef6Sg44nHT99JrlovFwnG4815io4Eoh
W/zjfKAiPGZ5CC7E7GUba0KLQpeVrPlwL0HXNThz9Ibhvy/OHLFOQimzoi1oT4it2St1n041KNp9
/90n7vkwC8SBzyEXdz1kDBGufNFN5yV1MfBGBaS+n5iEGpvalbQaKtuvd4LBD82XCigCPAnl9S4V
sDRx+lzb/cX6ircKrQCroCNpO7uisVqslOEsN4yDPUvJtENCktxa9ub9/cB6Gg5sL7IiADq+oifV
LXuRzp4sGBK+ZbhLFd62wFdjKY0ZzSMb2ZbTccN9hd/kMOIXaYiKRKciygsqn0o1iWrOOHLt8stp
pQimbjW65PryZy23FWgC1GzWAFWuTG/jXIMALI3cug9RUNUVl5L7ZsT0OBbXweR2m+KiV8tC5/GK
UglR04+k+m8rsE/2vjEGqYDF8KEi4AXDp1OPLV8VB022+gbHdUcQsI8H60ZsZfV4o34fgC4C+RyD
E6oGZEnUvNMsNWe6t89BMiFjzeXYEanmum02hkXbtaBuuVL6nYcbtRSityEYz6LZNy4J5yr14+gz
0qD0VpW7P0tXQVlGOdlh3Q6SxF3x6Xob/FrzIqkr8RYUHwN7LfXCtJILJygWJ4HtA8XYdaGNbZB4
fPd0aaEswsZCO2nJ5vf0Cmg93CcH9QoeX0zDvDNZG1hgi4SnVE6smrVzoLeaTA4iz9VkrtRa6Jc9
eC+f+YXDNw4cLlOn8AwV7q/mj4xrxFMTMVOlAcozq2l3gudlnWVOTKcWxPp80dTacxvpmLHlbocK
Y4/95cc1uJ4tZscsEp+Tb0XPASuHSDEQNyYNvzUOrYQGLuEf/ylDXwiqU9mVsKd9HuSlE1mIkBfW
NpBM/2d+roPgto9VKmWTyADaovj1n3Z9mWwDKUttzcp9+UaBcMa82M71jPKviIwpKphRc18Osz3S
pIwL6pz/5jrHYN5zgLN2dZ6b8IiAaMueidn92IhvznaGVvKWdJPZcCX3+eCnp4jEtrSOzeSh3esd
5qrcmGJelAPmpG068Z0Ppr+k8QXv9NNw+hIBj6SVIEk6wLoeIM9q2YiIT1rmFkZk7O7j1lxEm1gA
GUlN5u3B3tq04ZTEKm13Z8/E+izya/ZWoyJ2ZOnpvwnmI84RrQ5oLFHUJfww0gG+mH5uuvZooCmQ
I1XWx9H/9v4Rux+3jElxYbeni/A6GZcLXI0mi1ROWjO/mri+osdCpfo50tAU00/b7lsogckoTg4S
brLkV+jLhd2YVPMNFLNMGlZ6rY+K4m6y+903eSi2sFrLt+PaFFdJCXkyJavtfl9cVUYa6Mfa27ny
sW6KBsWqXIGWWgM72f+QQ/AZelpb/8MOf/yDJJgEptKkJ9oUhN9haoMoXKgg1UjcNBH4tVUdiNwW
Qc5TSGebudGslzv7IWIgnEWCbQRmCtoAIFFXuA61ON1kcbfyofmH3+YfxxL6dTVlpDt/7onVlTBM
bT2HASLQWHIb5iVP7K0weMkqBnrDeMSAighELkGf3RB3V2mm0+xg9WMvN2CV1KMJ6ttkRxVA5v+e
nrcvSlNALr1HH1tm9KAIqlMxb5BtnPbOFAkzAoAQ12n+50sFtuRAOowN46Gw6Q62LzmQgyrTS+x4
mGBvNr3ZDkTw5GzxAhw3TTvjGm++IkvUjcc/UJr+sOwgimF0bFSohkjfVt5C/5D54uAZ2Y+Ue31d
AQ4EISybr5w+iKdflAeAmbCWTYHSgQw0hML/jVpW1CLAZxAWJwTWuRKT3Du4EmN6hHaJ52dx3tVk
LO/Kxi6znIn4m33BR+wYxOvPoEHhe6iefPaGJ9Fs1EKV0rvvv2mHip5bf3X7rkM7V9whhUDsiti6
GakPAM6WP3Fuj+foC5M0ijg3s74ZWR7ZoENxnRrxde9xRZziHLqHCRoowYaXihaq7I3t1aJvXPY6
vZn5ZlsyRchwADCPfI6CVzuH+tIlDT+44ZndoJet0vyGIC5bysd4z8GvNhG44ph2sLYQXwuIrWGv
Z4bVAoL9SPYngwchYzq+AzztgwPqOqyZbHfXjtr+WpVwykRsswfVZrtfjKloMqJt0riByvvcxZ2m
mAu0K+Do7xuw8pVaTeHaQY6pNgcIeQOOTaju7q3+YEKTYvE/h3AnkFqUlO9jA81zlMyQhcarGYNt
2t0yj88KxuFOHIkzeZ+RHfvUHk4w+NYtM9Ut2ELJuEeAxXIbOunvkEMvrcv2U501hgsHH9j0uLOY
PRLf87M6X+EE6zpavFETiA8v+t0a97ukMkp2rT6DmHF5ed0g/uDyVXSO+St/JdvKmySXGtxBKoV2
SmrbGsxVZ1rIrNlzRmRg+VeTwZ6O41f4y8RgQNpE4whWvmE2vSdNIUe4BCXTFCps48wyg/Um6zzQ
gqt8qyGk5MlYP51IN48Uil4GlpRPtBjsUbYmYBA/OA0hdDrYnVfTYwoMqMZY+YbBr84A6FUjlcEi
QxZP8drL9B6nP/WmVLACLSj2TVkdqOcy982w7YitRlsfeTYbLhXnTqGHvZOpWcuTtALo53sgQUTf
d5igxqR580GPeY3zdRyAIfoWgip0a/hwVdMIWt2Hb6SKS3IZtsKu/+1xxnT6vNRWEJIsNvBu/rwq
lWJQY9wBHRf3g719MvsYZd4K+Sknpb9rDGRxr1l1M5L9IAlI+JEZuohy1Cb3qOydBXpVyLIfXc3s
zxl8Jo+TeW+1fsVNfZ/tyzD47/SL0EM8nUU1+eFX+KG0DhMMuQ3goMd2L49yJOplg9ORKexLyO6Z
U8qiS85mGvigGSTjul6leW0Uygxjb0xyExLdhEehmNWmBBxCwqHqNPCpnO0ahg8tiPNZZFiYROY4
yyNnsVhOzG3E38mLzlPUn6aR8Dr2eI1M8CP30n+shkD9dZML7+CX2ML+uOrS4uV2nkiELffFC4uF
VadK4ZmYkyQmfocvCLmJaf65TpeNMMd0zfFquuzhrYUq7qCkIem3nHPfG+E8YO5m/g1pw+Dy310y
eGRGGSM1HXkFlIYoAhGvS9lQw8J9ir38MEkMVlN4x3teF8o7ey0UdBI1mclR3JvRI5jk6rkMNEt3
k4T1eaySSEExsZAFzse3tlJF6Svtby96NI7nlHJ4QYVek+wEwQSamXxQCYz2ITkONIJdnZXJ3AYe
auGoWbXp4ZUdTGy6vHBps5syfaSC8a5HqHG9ZXY1JFclb1oK5BrjCBGgeWvbjMPXsiLKX94qgm0F
5X6N5DehDt+Xtwu/nQUzocYgAAZGfRiy4o0z/ykmMrJVlM/Ku7uD9xn+9NjVr41QOzTWcPMqzFHB
J0HliBxi8DxTgyfPxGAeDucvNXDdPfNlF3hK1VdL4qmQSfFjX4GPZKqCIwVIcmJ7VKrBRQZWFEXe
ezYPmww+iv9wvkRZwbEG4aQ1FHQy2Hsa32Q+/DeBVyOp7LJ0qBZVl9sgL8hFRxiqnobaDvDeb7Dc
0+vXGcqfcM//jwHVy6F+htU2wO7LmiLDfjhynZpF9NYggbk9CLTqfwnsNnGQW/CWHFwOLohawi/R
2Mi3jUjYFgudBAjDWhTawnDbMsedhvySO/yZ57HlVKWyUux1gyboySu48T1FEo8O3iOilkKj6Zi/
mcMfBP7+PWXKFMMkhYy0+epptAvDxBx7v2XmLJr0TkAP29B7SESX/f56aUf8M3YLbvlESZvUIWn4
39o4Li1cY1SNK+FUzHhlTg7gNMNLMvnJpd2K0G3/WoAHj9WflsflAnQWGMgx9KT9yz16foSW6twR
CGJfv5GyNJrRr4hQpTS8fF7O3rpHDG+StCpkJxST1WvMtcFEOiEnV3S6JhYGMuhGUWbDEWwXXM3o
IVEGnjYhqRjyCOSKimI6JWSY+Bn+JHRBPsTbaEFsFY5wydwQlhx4JJW1Qzy358782beFKqQqrVR9
3YGwT9sxhncAB0MT2TPyeR9yExnuIAA8kiThLK7pBIW2rcbaRgLrU4yV2/mZ8LfquDRz12HKFGpB
rhtpzoJNbbCpYxdu/xnEonX4aELbox3lrWMmPo83PoRmNGoWdhI7o0lQA965DGGxDAb+BlVpKVre
xNcFgbt8o2IiTgGsMBATo4l/GOPm4VG/6vkVnTQjXg0bseAubjqzHwl6V767L+ivgt3v0IktdJzw
9dR2Pai/r/tOl8IJXhoszUi5uLbx+pffiLdsZhKInoklCA4mANJXbfy69zkR42n2gRd1ZfoJcpTL
EfpTROz/SZN1EX7dC0rZXhQKa7f22j8J2V/S1+qxg9VsE7PV9uTg2YpWgYem5/KYbxGnwJb3a3I+
8FruTMlmRZdPDIwNLyYiINcp2jlusSMKjkqKkEiTPVjHPyCsxBIFCedUlUFJ8FLfh8i9p3L5D5an
8OpTPzlmS0g2rdDQD0qC2QJzi1CyDfxmHG1rxwK1hZc1ts8u0BfZjru+Sm7m0qmJG0aA7VjZ19f+
kiLYDePiAGu+nVQGAUpQ0KqdhyH+Vo7/OwJzDRAg32XAHJESztji6TKru0MYRwx8gbitP1jodqTx
OuZbopi28KaVHDCttNAk7sForYE03Qrj/iqP69FpB20RJe+m+tb/3qCQRc2g/z/PdQFSNLKgvzhb
Y9ej+e6KXKGk4iUD8swRVGDRpTBSLomWvscPe53QNcaWdBaMIfbkTs/n1C1PuddINhaflM+Ez623
PiWgfOIPIsdE2/DgdMLb8gv29CVXUp7zn2OlKxLwr2o+mSdfiPqHLi5GI7yxMTjlOHt7nk0cj5wv
/yp5yv2CI0++B/kZIM1tjx4dmL8eLLQO4Jz902Z0fjGe4HnVVD/ZCvKBtIZNOfd/Vyu6Fj/sj8kl
CqoMiqFQtEIroAvr/ZkTGOn4MwotlZy7izlHJiGzJyQFF50JxFKpqdQTASX6+CVXmS6Ze19gNcPl
uKe0+QdngjqzcKniF48rptGTM3dqK6yS00e6WjRbs8HbIBioJ+GRXgk6sUXssgJvAGPilzjTCQ8P
F5f872dOdm5AansS4i5j+EQt2YcfMPm9HV95IjX2YxeRhyNd0GV7tRk92/owEw5FBVSYiF/FwLjK
pSiouK103ZPUqOyRKiiqXzg84rVpTkwQGqPwPnrGccrpMweAw99z7JcIC8mv/qzB0eo+WYK8fYXZ
nQFVYceqI/hdLSWenGJ6qoTYjDX1wwt142j3o9znPxnPz+i3kBLF6ORn3mni7OTGmddyOC1WvIF0
VA0rUiRZiWAoxTyd9mSKRfYL249Izrkud4bzbDFCohQQImSCu6LyrO7byG368ani7BufZrif2FRR
k1j2jeNazhvygWkdSs2/FYb3d4fBp1MSBM7CRXZZgFtR8B8NeSeZYkaq+KvXziqvr0CKm/O/EkcA
5NhC8o/f5iS4MdR0WLA0xUqR9uQpHrMSFvDII/vsykjb9pDdVWt6hjFPgtHTbdnXBFdRvLS3JnP4
sq6uJIVCdqFJdyFwYiqfcC3kCyCavHcliqsf7GEc+B78gOLWB9ZHWpWZpw3G6eh6M+w1p76D/7tt
CpKdd5rieHo/+P2nS/mtFUEisUsUG2I5OZpt1jTUiAiCBkZcuIA/m5ls0SYyOEu28xJ1aOJVYfvk
8bfUhR4x9yy8vAj/2h9XDf9/lXnHscXKZsp2mLKU//QQA5YpkXHidmcZjQT3AaYwjvL9Q36wWA0e
4tdvlcZ0CBo+AAgyrvT9iZEmx3t/SPm48N6rEwdUTYd1GurKCEkiKRDytFaeyFxyke0TzpcleuWA
uJeP29qOcyzqpVc36e0q6OcAqMsDCpHrxhkXPYJGdPoAnRo9FPnR75RKKpDpW0qiDOXecVFVZg6F
d2p/TGG2Lp7w8C9FahJ/2E/kicYNSY5axjG+GifIYqtcN4BHbmFoOkwofUObwcAqyhiM4wnjC21W
3BycysW92K2iKCRqrLDMhp0VOEqFL7G5QkjVRLXVUk2j5uXgOZcfCLFAOmlfwCr2OftX1OkJyWkt
P/622kjJ0wDO9K209ucIgZygmmoAdsXQfNWxHVTqyUeMhuirmcMFYi2Oas1RdTwLFPihjVQbl3qN
yV4zn2JdgSYsel2lFEGfZHskKSIqTzUy177Vn5Ojb/vZLvD6klsgyA8k+Kd1bOZzFfw0XtFSP7Zv
D6NG5UJTa4NWQbyPkh3VQmXKTKYmczstikRsgasl8NpU3KtfLJZBImIVkZDC9qnp2L++j1ycUJ4B
eV2gaPvIV8R8GPiFgESO0wLUMrdrM18Xs8lX6r+z43nE8xDslVjz+ofCN9sBHMVrT1czVqKcqLSj
Krf8YuCIxAJVcIWAfmz3fsERfjEAMj9z4fMXsEa8+/89vGkItYUWV5hy0b7QsuQfBT5uKHr+zM6C
2wfllopZpUy8u/mqbzJg9w7IAFe3TX34lXAoweFc3CZQzDZ9kGDwZ1JnEBMK43Hro1C5C424qAse
l+uSFG0ev47lc2/koJXEl7rW+9puOuawrn6bCX5SidBQA4VAAsknEEOVTwkPDXut7For9NXQ9Unw
HfnuTPhKl6FlyjLG6KVXjhWrDwsgEUheT7cwSzCizTdbOWHby6Q9b7W1zz/RQnYBqyBlgdkgLQw8
he5YFnNzBFUn9bqB+9IR/gb7ghMsf61gQaiTbrTvTYDikwLKyOHTuXH/feRonAWJigtUcJ6QKHpv
YCfNCjfKZ2dn+EgTHcbcAFFOC2xTMLxAYfG2vsxpHJ5emin7R1kEXqhWA+Fu1BHYP9DUqzMDw3Tl
o0IWo+Vwxza8wpvnnq6276lFskPNcQCfc9MOnE/90cVGUAEHVy/sFNekAYIevo/msLIhtuSD7SoA
6sK/iXQp0tfNaXozrhpMdwBQsNNvfB6ztcsp5yNX7cndtZYIegdy/55iWZc2xFGV+ecuTgXx6nuz
RqL4sk7nt/oVFXhkjX8QSQk6Si/r9RK/Mdc08+w2fKQgxmMReFTaeqzfFfp4/DGaPwMY14Top0eK
AVh88QlnaozCHeCyY8lIwUyrl9NMqASkKGPvT0I36v7pg8OAm+VQQzwI1pVpPVEc4o0TpqOioO1J
FI4MjFtC2Ing5LeJ4DRn56/wUszuJRSYSGlMWuc6Gy8nDk4h+z2vtFtGm/4WUMx5gFx/Oj7sT5+g
cqCoLUExVpChVagy2AmqhgQ1rgVLh7d0gEtv/8RotzXrqxcBIk91xB8xk3xmw/qiB+tZ25JoL+uk
f6QipaYgHhwjXe/DixhdEe7KPFTJRb2T0FPPuu+LmRnsgeUI0Mdvx4goes2cHrDlGwssu8jC7PnD
ITFhC7QCC2aXChnAih4v+GNym5wzWmklyf7f+iU9E+4Qewt5d0UqjJs/WVhW925JDsK9GeylbaSy
HYMp4o9ai/+49Ebcg9GHP7stVoL6nbpmfXjwID3jckX8SODPSgPUnV69MZRfR5LmtlIbO5Vcz+bC
PXIZF7O7E3GWWSz9I12bp2vv7q5s0gb2WzEt0rqH8qVHF4i0dWdPebW4Nu3sPMYPbduG+zam6guF
ri5qEegYS+TET0rY20auDCdvnSHx7OMtmm4LbuwpMmeuRIURXd53oA01gdso5jpqOEsihikQp1kJ
chKPhml4bcjIp9eY2fSaow0Zx5VOkyoTP3R5XrOLOtLKx5ZdQcFBkuT0XiXH9yR4Wn9GfZMDrqdc
41DpLpp8IBwo9fOS++0dCO0rLWcn5f1ZtUb+uADqurufRflWpfzBrPqUk/y1/9hVZa+8630BVbkH
5UhVcFGzcuyTh0lcI049TIEBb2dCDNihXIukGnUawgbX/YyquScNfbzipSUmE1tY5lP5jFf5F/rG
tJG3HWZ1dVkizdufCQWfU4d3ap93EAXjZjBWoIQi8QmUaGDSyOyw9o5MDSXZP440jBZZptSpW7g8
GwY/GbGJpJF2nwqh9md8hhPRypxUn2ER2a5ypyshKKOyzkF7sQQPce6eeZmEGm7OtyyG8zA4bslv
6MN7I7HtRbVU9CGPvPflm2neAGiBRQQ2h4FcTZyD8lXSDlt+u8GkDFsjoN5tq5HZYbfe4czucL9a
UEXlNJ3VJNbyFU6XzNCija0+28uQUYRTh9C6lwuBg1OoAtmQXAaoHg0RnovZoF+RRGFFjhOi/vRw
vQ+CcXxoDVFSkonOMfGtxirS+bu9m5JwQbmzlqmZBd2agln+tQxqrJJz9Atu+D4zm9w4GMfxMwFW
y6lHmQb3Hyq3PELMdClkCyEUy+5RgCGUmm9k2Smg0/vRoXZt6VW+5yeqj9X5sgG8i46qE3bkDKNv
IMd4NaG4JnwrBDo1e3vMxZ2qUoiDDuLY631zqpbjpAPUVpGhDytLo95tKUN3SmJCIq44D1hSSzlq
SfrVmei23LoNIV/f8fMVNynlVplvljvxXNKji0DlhR2ngMnnn/EN1EdQlR72f3x3ui8RKp6NgUu1
BUqCihSX9GidnpUlcBg5/hEs55PJqqRLVWHHIPnul8C5KWBqkEumgu5Ck6vTKMX8QRZVIbZ50A7h
b0VILcOminABYm3ze3q0K2fvkQETLH7AsHQubFFyGAna3Y6/VxeQ9fp8f+E3eyryvVw6xvyQYLvc
8YOtsgY4Wbk3cPbGO0fVAlau8ux949Kxq8KWecPyg1Rr9wOffBXTBfNURDwDxePTXJM/idLSvI4D
krUUPFFwqos9Axtp5oOd1IZue2YWWs728aNxqWQTDOHEUWealZ3uhYz+1416Wsnk3n1XgXqRb2Uo
+FtbgfImes3+YtLfJgwr5QM73DmEwT6AEaQKPXFlZU0k+NVeIW0wXwFV7TJg077zqYpxy0zcY5Y5
c22J1q9Ib3axJKAjtZdptYcVO6L51igcCyTTtBHY/BQw961oLZGDwAsvY74BQpvpYVx7RWtyH4xl
tStNxHAEroNU0L3Q8b54p6JpccRSNc0T5eUZBmqpPEei22fKOR/fjamcHZjHm3T+t0l4vr190tdN
2HckVQMzsmpjT+YkyoMysDtU+BDJIeicMFfCi9WM3zP8LzAASWESKfZFoIQOSTuonsCV/PYWZ4Rz
WtNMJZh0Va9VZMLxWKYFxdjzPW2nUJGa96rW57UNcFRQ74s08Mgou5jOkPMdm7AwyCUUJPOcA92E
DOfzdpcXmVXhNG7R0VJtbLCHe5qTzs2SDmyyK+c0zyMc/PaYBJ3q9P0b7hLLEmi+tCtfZ17/lu7V
r8uhp4KblSSQdsjsmO4hCOKvVSE28xaVFHkzh7KQO922PHqYkKpWvoxLgsmIuh2tSgoLbVf/hml8
Hm9u1GSYCPIBOIIQaIY9gBp8HbvTNmVgPyjrRlxOBx2ZhuNCpj/cjJXYPe4z8VqNbbuOZ14hFRSv
glzOYOP5YKDEGBhewIdwAeojn1+ECSH126UXA1qlAn2L7PQZIkAFIbDKL6asO+p4+psAgGFrl9VP
Ie+KFlX+scUe2v84OSA8H/6qGPmDdVoySPiaM7G8Uqmk9Rbo3dxVE0A/TM1S0KiIf5SetQLl4w7k
vFuTwTlB9jmFr0fgzYx6xnsSFePN1FmisF0Jk7lcRfalutnGd+y9/V0Vz1JrUei0FYR0rDqMVTSg
zPs/lIJ/O7Zz4OaMYQ3tCWqCfUd211ka3JgYEw+EL4a8bEWi9YeUhQeZo3LBEZKEVoG2NrsyL1pf
gR8P0nvnSrJl7pjnt1TXFS29HyU6a0ttM8vOPLeiKtsXI69L8SSqDFftap/cP8QBr37SDXdxdhcp
2MzfAn/LTFNmS5BuuP8BbuL3v0Hx0SeD0ztsOtYecG619U+XQHDYDsXN+xq3jh5BTDSeRqpIu/4Q
9aoGt088MWBzKg2Y5GLvvw8v4Kvwlrpb4GtoUqSGjJ885k7Mvc2LRFjdRc++RgG0+RD81glYqvsx
gF5m9chcJBw4rLw44oL0tkHodZ1dMaFZXPS0ekAsR/absm4g/sYtg11EfTvgpg4cjaH3iiz7Rv5e
vjoox4cqV0SPghddBDAhyhhtBolDcrmN3CYSn0uVfMPNNFB5ic/gaei203Q+Nncixis1qosAGTgm
n70UNAuKSxuWSHxQ7yjwz1S1S9lAk4NVHe32ecEh8XGcIqjCwTBKk99S+o5zERIwRmm0itRL6MYv
6f6/KsLvRQ8CLY84/Hz72ot0egh+D/jBRTT9T3uO/lFAGZarYN3+0D2xDKKJg35ZOgX5ZTqhpElg
LHp/ru+vaRjl+4UimXy8hnyb5Zseo7C3sOCN5bsZXL55Dt9zLVC4tX2+TW8Senex2kjgn23VMEGI
ZgeSZcNiGHMfqx9AnXboDUp7BVC4R15E6guVDGybpUwFGvF1Q6ByxO0t+mVu5L/stGoWfcq0kYxB
ie2Yg4kJsoeSdE7s5ESutEAH/NVyC7Pqplr0aS7d1IvVSpBmcpDhiIsDkfRafW+YAuqjViA4Q/2L
n/hwQwuOH/J/gKuNBwa4e/DhVB/5HZ82ua4NNupc80AHxQ3Ki9nQnE62Mh3zN0wD4JEbGyKYx1cX
Tm3U3Rn7kLlmtPjz0FX77eDiaXjBnz3d42wJTVtcVeEbVQgzevMIoZ8uU2maUR12XN1RDQP56rDG
Zq7utvTb0dP1mwKlwMYijXdHHNw0t821NuZHx0wHMpZIUa7j1Nx2a08sRWaYdZC9QUCDGpCgwB3P
9lqxU3h6hicCNj1Cl73boxj/rePE2PYDjdKHOtE2ahKAByuIRHOpVt/EB0sM9PjWXJbpYjZoyECG
mB8Z+AR/sWUjFvwpssMpcWKmb6Z8ZFtwQiy/zc4C/FPlBYrEiLPUdPHF2lLtTwvgzZNRCirMynDB
MKd6K+dHl4CGr5tNXqpS8CsQiQ+vEZOvB61IGVMsaHtujW7qtwWpIXE5US6Eax5jNN9jlxbtEpqj
HfABFjwAjGryFn8ujsMqFk3tNN25BWuV51cul9DrAbcdAfYyWGh3L/N0bhrCjZBHPFCJ6c0WBHfn
gJyVmZ2mxb6y22i4gC6fqv1CLVL8rlIlHSYwT/qTonOGZ1EOczor8NQMD4Dds5MK8mq/H8hqfGvq
HcYuYbVxLoAsxswmp2xNJ7S2AhOQW/qR5ax25lDOM34JI1X6Bq1yW6g9mOxNrnsTn9guEnwPVwXm
F24rLG81uoQpUaS5UEcCe9SMBR4Nq9mAhu/tXgjC0X6cFtmKcPrldL23NCTvSgVh2nziBj9QXQLa
Zd/4phibJpDL9H8rP1o91v/zdCx9s9KfOG0V6YIwIP32w0zaqrjDqLV3pNQd+cF/ECRM1XhHkf5Q
31wfhDDnN5y7oNlfrCrZ6Cffj/If6hYGkIYi+7YCCrEGNCLWynPO3TvKmmCFKelX8NmQr/b8abeN
Ugs412doLCoS0t/DFWLtALfunmkjNjTfmgt7wMpW2IvWBTiiiEdWFkm2ogRDCqiCXMmeSmfolVnw
UW7J02al8o2mC91bl7VXHPLF6tGBmni1cqeyTyI6VsZBPlwq49VC/eMWOMjE6BNp1duJdNE6HSRC
DMKMHeOSbikvb8gY2uNH6ZYtgiPp73TcVnVthc/2c2xDoh63ProLksPYT2WUCFty9fXPvx57aOPm
1UZ4lnQxpC0dCvan7bCaNKcgVWksAVyNjqz8qazqNqdcEtATetTNkF/Z7tx1DcNwvoSHgFscZiqt
Zy5psK/Ndjqr0ae7/rMiFCZ3J7ya9qjZOyJqyfd1a/1/VgDw1jX1o6uBusDS5Fp1xXM4bygoYEVX
QINZ45cNkxESCOKULpSE+9UtZE+WG6EzortS/1eWRjRLC8ouXflmB9fgC0sCALQx1h1dfESkAhQM
u1J/XRslj5bPB4IZaAsW4SobJHVGEzJ5jhCyrbzY6DFTZmiWByiRKoU9yINb2Vfza9tX1CPI3jyx
PlG74X6PobI8a+V4n9maeF0iZcHgp5O4qMmdu+8Bl2fDnSyH9acitOQjeQsQ/5ZomHUewRIK1nKa
5PtVKCx2vpwHObsonDak8mR0sEe/gDpvPbGrlh2m1WHLYrEbQfQOIWg/0WAW+t6Pq3iNYQ7Wty36
q57j4Oe+sS9UM/wmVUsFCo4vqRBmHXnZ4GBm8vc34Nxn9JaxQ82+Ec9dyuEUTaRJd4AZtgXLMcsJ
r43l34baz9W1uVGhirrgrLG5Y2PlQ0WAgMKfHKFZ0sVV8WkjWOJrU+2Jad45cv418ZJx57Kmq9iV
KOmHA1GZbFOaB6CxUdDwDC4K1ASIKAmd4DE3EpMDOEHd84BjciuR1jcSzPaz59sn/3WgSbdnA5B5
7LSNniKUkeAcZn7utNrQ+FCrGh+d7mlaSZ5juzMmQ9H98sI4RzTtcW1g1y2axopKQmAmqFWExZ9Q
l2fqNlv+p/GPVoT62DfZqzqIe3bJa0y4RsE3seUlOj5sbl0e1Tip1TYyy80WCm+gyem5an8h+yRG
4tvrBVz+2Y3ARzrnSf8F5+FWd27+utYIFfASDBt7FMT0eyP3RM7Lgsewns9GEJ0QUE+4RmsDZVn0
v4S43Q0XpkmlM29pz0JYTiHkmqAqvnw99T09l5626dl1oN0PMTluKsOOa2u1hKKSm0TqhbrzhReD
SyZvYAYqblEhkhSQN+azHddHjr4qz91l7Rs1gmYJRJinQokbLyvTtb8zxe0FP0aeCESSZVGnB3mC
LYxrpYIedt869LjMW9/S7okSRFmPBOIOQXwjRPXBzzYeceAsh1TkeIqcBPKew5WEES72ss/lzJ2b
OTTkb2i1nOc5B8yrzOy6Ie5GgYwa+5gScmpsxpRvhmGs0I931XsWPkCtlIPWMSWkIlWgU4kvfHWs
i7roI4gSATa0SVsNfJWXX/5asib+OKPtGrI1T4AT7eqIVnR6q8Rw8LXEmu3Sy2JlbjvFII/bmSqN
LGHvA4LjDiTJnJuuPsoJpyx0DgMzymN0E6FzFNv/VCt4SGypcBUqxT03PT4LROvnKPvGqpUmBS7k
DJ/nSnf2hOxNe0ww5+O4UTtPPL8UZis6os+xuqUQmcqh3PfM2mpkxjMOKPbj5+EG9mhp9Tuqr7KY
fYlBOpArB1LV/3tSA47f6v9CsN+fbmxv1sd6awOQUvRSxYY03pC4O52u+72EqYCOd6YYJQr5dPcE
bMAUAekFmel8tV5V5M990oCdMZP8dfSi2AKilb7C0Vl/zHzZ8at1EJs+V3PPmeyYWtHHNQiEeHNA
pE5NWF+TkG8ASUMz+5mp3vbhn0/Kbx2VIBsUUzlKgru69CCtEznG1oZxJKpaMI/QismBTbJDYkS2
ggGcGX6gdlIjf2RL8EiPuZ35f9UwRkxYE4gjQgON0el/g1o9mrKLsIP8t5mPEwySxBO1GeQDazfm
GLlZCnS/LI8cg6WUVeptFfidrYIXlwuWScBnkbSzb9fP8bDlw/s9/TJ0YnZ3WlPhsjTZoNAxNb8b
6aYrVlaQYyw4P0zeaSLy4YQp7A7Xi9hKpjtH7VZfAWKQYf7xpxKvH5jmnMeDlNpDmVtKOuc0H2wf
KUyn6sHtmgUuky/rKwqcGcFe4SDTaF84A9MpthpHuqxv+wd2MlwKZAAWaYAXMzZTwNUhHlw9C5Lc
G0TS1UwqcDka7aMyWPBovSamLlcWk0BOLFz2VK1R/mBJk+unT3ZImlDfgRntpWt7lzORDb8d3B4n
QHY8L3ZM4KfuFNGUe/jC8e3hsUu3t6SfrHb7i+VowoSUEoR60e4N/CDJKUsvqgsZ99onbHmp1aMG
YYQTVbZcL0ii0y1O2xrrjD/KasS7Y0g1+je7feo+czF6UN5Q+V8f91RElakwC8gaRXFp5mZZ6RjH
XQHkownXAbp0sgvIh2ZfK9gJwPI7s6B6sA/I9mosS3PO9gyuVBWnD30VnNMt5cSM11F1sK49Bjy+
IVezhMQxNAqNXavoKZIQJrgfvlTnqbxaABiXejYr1uLR5XaF0hI92DSU/M+40REAI7IoeYVB/9C8
53eAtRTzOPSNEOVmNGMjzqI19XPXTj1LaK0WT1565+gwrjQzRkQzMUV8ZSlCNA/1NZlSzLJskhE7
bWdyBrZHQwlIeC9PmoNJUDz4Wm8N8brqGzVMjahUJgkX5puqwdi0diNwCFnDMYK9PnFEWeg2ZMHO
HhpQbrC/eUhoUKYJi2DOlFdWQZgDTdfwX2xR8W/cPZZUnvrGE1YKsM+vSiytFYjtduvoKU5eAeLn
R+a5vxrqog4ATlkCS9QBSYjt9FAA/2dA5panSMvMkWDV0hkwudYHtEvqAhB3hetQ2dsLi6z3eyZl
KeDVj4A9L71C2/aAUZAPHNagxu5bSNoVv0yd09gZ6j/VUWC9KbwXHL9nXzkei1ukwpkwqkc+nJ8T
TO5GCqvoWFqDyPZZCcTSrTsCJEiLs4BUre6q21jeSTpmYd6xA1wRwG9GIM5GYznPvfJF8WBOBOKW
s9EzBZ0it6WRV9N4fZlwjMcb7hFATo6OoH06qe1TE48VuNaki5n25QvOCU/N8MNf6TmfHAuSxEny
lzUfBj5Sm9BQ6tcEReoQgu1UUtMXyzomsjCXUMmNPgtUqzAH9FaFjGx/LihksP1NXvnHCCkpWuEO
SDXVTFTUHfzlLRxovsWhkWQ73eLH8/subl7sj5aerkyoF8ol/8owTMwO+eIRMetJ7QaZb1MTNcDB
sYNLjQU1hNeEqZGP6UTU6aew9gGerRIQFjeR3vzT99++PXVUb5HJ4yb7oMkK87o5JDpxA+ypG3MJ
tPUTkOzyXtIH9fUPurd31OdLI3x4V5yKF6bFMRa1zGsUnsjpFMTOmYZhIT32H/tyCcVzl0bfb64B
A7JUANe2YNLypJ/WkaT9gLJQElu0NkCx4MOB0IWud0pBJ1CZaK53jpZfsRmMWDVRMirlssD9Kcuh
OCwujSJUB9Sc1Z406annvts5ITRFE70cYZBlHX7JpB+VTOVg6a19DfMOgNQVEEjxLto1ohdBrBX3
jWo7l09O2z6PD2ZtqEJf/7mxi492ki1nQGof8fUHJJF5FSvkoSsRgYWYBhkeGvpdGb/3SdA7BzOx
bPhT15gyb5AIzWjajM14KnaCMkmW3LIVgRo10kKT4pqiDCE2Zkxj/uuTERRO+n/P/g7z/awyRRZh
bfkzcjAiOEaWq8x2pJ3cV1JcYskRz77xqw1MfzsBqzhyuLZcbRoqSjlOR7ng8BXdkLpGyzgC4HTK
FhF7ljtz6r2y8qLM2jlT0dBDbC7+ErqaI6sWD8Wx6f02rYBMhqhoIDzYKKN80TzoIN+IAgx99Ii4
b1XfJpfdmyvWUPnEBuzyV2ASqU9CHyx2Kf/fyr71l+YNMfGwQJwuEMOzLQZI2EvdbScKti/zNPQM
p6zJs0NKuIpXvyeqFIN6L81YTOQJB2fgIsf8LXVYctDN3Zm1OsNzEr7Q24vw6b1dqZMkTwFznKYn
NvE7pebWITwHto4CxmPzmt8JpqXe/yA+ePfwr1XwNXjTAI5IiAW986b4IwfcFUbYuc576z8ezeHQ
OU2C5Z7IrR9ob6oL3bYc9Xo21CP0Dexxb9/nvw+m86MfOxGD+2FBFf0W7LJOs3PBMl3rWDW4m4ut
KesvTKYOPFDfdnJSomAgSuss3DfaXo72DAyse4VZt5FmsXyBKs3prgHz5D1BlS2FGrewxekJJ36O
03PU6LP2579tRCe1lEd/tVm+xeTlt14GbUmXx1g9ZcTQ/Zq8ttOyo4bDJtAmyRuqCOYEDi3dfxpf
8TjplMB7xPmbHLyPlp2sTEsbY+7uzrxIm72xqCUqWg3zkCBV0if1W8bgjIoRkjNohG2liruBR4MX
74QE3+W7sqHKgchU8Q+kCzziU9Mu1o5ESHnG7EMlfQFtawFvPBorI02Rbh1TrZ+yX5cDSkezuJ80
3mryY0RpZudXPlC6ARvAmj5bh1aGiFMZgoqz3u9bq5AO2sO5roKovF3YrmkRQForO2+T+HW44HiM
lfXVYN+PYmrBEKLBmIUNL9cNdX+efioc7aHrTVlJ6rlB4u7iIEqLS81UhEFYmreWYwuEZmeGcpgr
kcCwTwh8Kkb0jmqqMulbBqWlC/mP03kXaQBP1kn20yTsa5mi/TlXsTW5VuS78VXlqXJQp4o8Eo9d
ZwY5+TQmOkwYjprBnP2rF4cuW+UBgYf7Vlp9EN6dFnAiPoraqeH5TT/gFZMZ0LGwGVBgqieZipTu
cIlZJYvn4HGlrtfRqfkvRUetFRPiDFPbDYYFyuRG2DDLXWIAGJSEAID6tSXDSwOLmPpSBN15sCCw
tCwIaKsb9jQZQhwgHDwvS0Tyz4EnOwxrra94pOJ60g7ly/ReOERmfX9CbgqXss9/PJev7Mb5sSm8
3PTuipHiWvAUS2cladx6KT6klTdMNeo8ulYqNxNDiydRuPmq8UlGlQEG/17fvmVreclaef7Ln3DE
IA1lDfRP0tGXk5wkjBNGBWRRjzu8bp9NHFJgnMotGrGijL2WDQrTVPQnwiw52wqFcpeQbdkTyimZ
7NZ0ESWD/dlvL5Va28lWZxap89J6G6SXBGMn1H7/cfE1ejUeHotMaRyupdz1gF9230Y4rtnHi6DT
Gvf7Qf76Lg+n1BMJFRgBvqbpaZrSVoo95ZEUf8WavJ7Mb+xJOeC3IO7Bbk034Au1RebdgLsRQzjn
M9lvi0Rf3YJ2aPGr0grU/nwJoEUWWP3BhElDb5+EzhATXngFeit1tNi5teRaW3BE87VS7F2HVJw7
/F24OJZ4jEx7WO30lkyRfkgxdVytAbiZKgwVjZSg9rYPGOyzJtAeSQavZW3ZRISjid3AriDfGGF2
5Vr0Xmo8ELLuywM7GMkAKLTTX2MNbaS574FPR8D6Y0CZ9yPuQeuGZ0HoAM4Da3YcKmEeGV7+kfHv
wzKngbKcMnzMqfLS4YZY/8cG9+cTG4VKuJhsdCZS56X5Nbb8HEJd67ZDt03R9SoEPVxo8c2BbEyQ
zACCoduTdkyuq7lDglj7Hp3MwjgGFOWOiQen1YTBsbNINU1ARY5zksFEV6SG3lVWg1rXDImO9eDO
YSM6P/lHCXkvLwNgrLUm5DSBDaRYhhYOIYkhuXQ/n3Cp8kM2DDwFkx50TjrxkIgDFkDf8CukulMH
xG8LtDutOAfruxQq9wEudU78zZJuBsDBmykKj/HEP1C8KxbD0lixcSoXAjdEkLfneO9KuSwLTfT3
k59wfvL4FQe1LCfP83/CF34bbOHaWNlACogABF7gifq0GeqYQ5lwRmAAOEZI2vo8n4kPcokN97YQ
8gAltqIkK30xn185sgG7VsmczgYf3Pk9UUgJMYmp+4w4orWrwJPCAZQ/AKXAzV5K0Gqs2w/JjsWP
pijT6tFj9Uhr56Wzb+W+Bw8/0unQ20xHi1IxkCXTltVIEqMw6Cp8UIRKlrsE26jmvCtQvT6MAMg+
PHefqMAmmm/5W6EAKfE6M0RnWJutlt740lFWPpzs9VtFjl1Iib46Kaca93RW3O9WD1lOLd7O3kV+
lUMMJ7MQnpUADBVNkTqx17oJ0xGhlETuvh+LeN0WZactfvbeAWL3YtmHpyzBEXLncixlCdiAWICk
1Ca4FXgXXFRluP057lp6GTYWRyjkz1UQ++6Enlv81d1WGjfn7Bebgv0/JbeTw1R3AIaVgJK/4ee2
8lYroJAx8BvzyqMSPHy6tZkK/7SSDDNtdbaBtL9WS5CIJb1KAZ42hSn/0a0qH/PdW0XN8SJQ96Bm
rZBJzcBhm9Ye/98eCCuni8DAzFj5zFGSPdiu83fhNaqcmz2RbOm75x7sHsDue11J/RsEjuAwHovM
0SdTr5P7IX0uZ8v0b0HUmiJIJjhyhc5+ny6BGX+6twsGi9HW3XdSM35bbBb6i2Djlm18PgC8qU3g
X4LplIiFtGIx1l+JNTP7HydaKcImlvxr6xVttMlv66XiGKaq369CbSh/wvhRh8BcUDQ6Nc7nTB08
m/DCuSBNZguu3a+0n5EmQLe5KStyzG2H9Jtz59OphOLnirUsuJsETqrSmz/QAcIME5iokNKN4WCV
KM0+App92ek2rVY0u3wnF1FV99hSNI4yfJnGiPPwKEKpSfsLWA0IC0ilAXagDCwSw+rqGodzV1SH
hpPDasoS0zGRsFqOtME/QB7yE2Fe2BW1uMg+ZfgB/nrk2TCOY/PWDFsFuiWeFX+n8X6yOIq8dDo+
+TDILi58V1m9js++3gTauaxG0PxrQOXBMo1u8BOSMt8Kr+AoYxy19fkpBe29EEQrnJRdeOHP3cka
xkvgrfKYF9ZLnP+IURujGWwVOmK5LqVbgs1dpYZE2OYuNRfQIF/OgdmNuCiTdvNuJfKcxjEAFxqk
n8w5TdzhiT1eGu8Z8t4XPm+RMb8uGeP4w7pv4EuVzesl9jpCBJoo73MvqL9uYV37MR/TXwVV8Mzr
nq1xo/8h9hqUXmPoaViOI4z1eNYgId1XcC9EfZIo4/+4Wm6wC2w0fEJEKgP6LPXcN7Al9E4ceSXW
ZNuoS0MD4WxOIFSsvFvKEkq3vKTcWipGiyhD8iWoycLJVvd6Jquz4mCdVBLM0FK/hRkOborz7DB1
f1g9RtVFKiZFcaycbmUqckFmBzlRVs0llR7uk5zqopx82ZDibyeHLUMnH/WbGobYnmo5+4VL2caO
gr5rI3m7HLTkUGap9Ft8k5ELxJDDw36kwv9LBfbmzS5UQVv6uwPZczs09lOd9n6aUJBfgwRZVHFJ
CGtGvZ4YY8wuIWPACVggsFrssPrpbCGjtWDnxokirFcafdmO1aPcrfJm60ueoM5MIIGfIPNG+UE2
/IVy+CQjbn2BW2aK2O52zQTY3hMo3Whoj8sOdatrXfDXmj8ZJoYjE54QwNWerSCDv/GVBHHksaMz
6bcvqBPRpvYXScMvLrWGr7PUOwSg4EMDehfmGrB1Q1fi0GLLvvGh92F0AxiSnZiB4yJt9Rs6wzG4
tADcvYLleKcMIp8QOSv0G+bN69YbNABKQ1HQuozm/QQwnhXbm8JKtoBaK6HdeFWOD4O3OH7FnvqD
wLXlXqYCkYNGSBPGmRKUyFgfSOSEyBc7LEm+nOBQhFZ7ftGToBpiOm3ole+fRR+GmgWdAODWa4r8
EDDarUoHjAcTj2eicPRLZDK1eTkqMrgUrFomDI8w0n71D/eF7JAktxZY7S641VZM5VyL0icBgsWd
L4m0IevW4QRoGWp0LyTCdOBKfnUGKD9pqSYBp5lpLjsFY+nUDgVPpv2XmvCUaO3hPZWX5LDyvRwc
s6k+fDhsi8bSYVuA+/d9fZL3NZSkJDgZkC+XG8nagkeKdINy8QzlVbnkL3cS+s0FrLQHywZ5fwjV
VVQ3qsUqqsWQWcMbwu+qP7ZqnfxRjovXf+UrJG50fBzjz6qsSJsrTp4YYtr4cUkJRrMMd9+Ot8Oc
SrPnL9x1Y6DIoxm8Nfp+mBjMdR1YD1X69gUbpU5f5SKYnNQIyOXn5pmTHZ3SwLCgE7bL/tuTNdCl
q+u4J4WUfkuuY6X0n54KEicZpjYqSmyMbQUUFAEKTjEVUaHT6voE+1kL+DZG0muV1HNDKIiN7g45
ZKF6OLsAhMHgTK5PyIeUy0RQ8qwnNi+ziY6YMzLD2wJtUHJuIoTjPcV22Ad+SCXu0vOvCcJ7YiE4
UfmoyhmgmYFfdFR7LNmziwfAoAKJuT+OA7T0XS7rI1xmSPSQTMjn49GL93qO8TCAlZaSYo6oIrBd
t+65D9mvSx7yRLpufvy8zV9arobdzZPYesv3agW4sAEi6l0X889AsT+VNzAx/6539jmVyxR0dZmd
UOiG1pqY1pYShDbX0Uh6AiAUgPMUVws3b547xx2+oWQ9/n9pe/j4p9pi9xrlra8hvksbsoCLLpHy
q1pih3X3IpfhAkeWsVGJ5TeI6VH/nVClXIO0eJmUaJzWdo2kiqc8rxnE/5Og0IMx14iE+HU8ETn5
+XVf+fbHsT/BEdNZlB1PmwLYX+uJ3WKAejNvXpcCWKbIHF36DJXGFPyFbRQ4eMBmmykONMt+9zO8
pSObNSB3U8EA8Vj5W5O+rxO1faj+EZWqd4c/d7VdgDKLccwar/LJqL55iy9pDkeZBoRrYKksGKKK
V8PIRmdyA9BkvbdTJndY0O1DdOMncj6i4J+cRpUS91DWGXAr0wnJ3oA5t6yX6ZjZFLrKiwryewlh
kEip2CP3jf3LaZc7KkYUbuHcvATXr0G14xs6zmtSQM0OZOmDQdBKn3OFvQwqWTy/kTccedb4+upm
1krPGUMbZcm+Hux/2N1i1X8oAHeI4o2qWngfjKsh8wL9vT8g+pw9NP1UNazegtZAedZGG9QScnpK
jgAVRQ2od/yNQu19JlbzEnNMajqCrpWkgWf739A5PsK3RuRfVi5C1kA+n/5Uj9jsMr213Bd/yMPe
Goz7EDSfKdcuX1wLsRrCLytnxpfuMkYJ7+ijtpV00/kviJecmluIgu9SdJhq+nnOK6/SZaCnpZxJ
jC2y/jArzHVXgouzeqN4QTaa1nLvUf+/dlmF5y883PgpmUkfuvnhmL8P/Wqu40QwyD5Lc1WfZUWO
rs9EOi3CJ6+osP+Ei37VNhPu4EGiKc2Mnm0suPfviptg8TR+ms9VM9qdfbslsEUEH/y9pIwpYuS8
RnOgTb41sTlAPuJKCwWY/WZYNqryW98uABD7Ztz6BfjJht+lbOHr/sRJTX5dhucLDMhmAN5XBWFT
8QOVc7nkRMv5BiY32uEgMOuO0OISU1xTt+ZOfco5GMTj/1QgPwHxhFzMW4BP/AbvIfWYWssiOHeb
vBGmTA/as6FzbuDNoM2BC7NMaeP9Wc0h/NnY5GMVgHZIr2vo/anwKXGs9Q06vdmaY0xffN4bPPDl
308lsGfZURTPLgfERFDFnZ37GtG7WR+BWJvf/1cCfBQe/0EsFRfiMpmja4tS81iehxAwZbzTITEV
Faeuk04eBBaUyD+Wmw9qCJKHwyQhEvqy1wzVdwrKr5ybee3amMxnG34+FTQ4GqAkx4BWRmF3jYH1
OUW7yH7L8MjZX/cgryzXo3WH3shFQMD0Hn2EZ75ahK9THuIuml6tp3bLONBzg+PIxZACkIwsC70z
c8H4nu8SKrh5OIf4tR6i/v8IghhPB1tUWAE6ERumnHlkySv2BHtLjXjUy532mcSml1Tz9u6DCAbV
SSByLiDYLZqSu4af0BLeAB3U0bHo/4GQv1EGg0q+yEWpAO0kGROVmTZjT3p6/QFnt6/uSn1alKU2
UskVbgyK/haDqr6aAiLXxyKKgUGiiIB+rswI2HRrRV2vOvJcgpEZ16s7we3whEwnuYelRRGrzQeE
CKYL6TToafko6tdRGAut3VYq+8GPEyp4sO/m1RfPqps8zhcRqtXnrea8G5C+b7yLciv0QrMwVM/M
qERSHTO0tM/MaBRWmNFIy+XiJTbd6SaCTg4h2K9RhNU/IKyV3VSD1u+4c9YMz5DhJjhXw2x+g24/
YZ/NlvyXZfB689GzDmDmBfG0TQ3mz1XfI1uhU4p/wmGd1GXQFzcHOGu+yysKuX3R8mjQV5c10PMO
57EReTIR9j39aFmInLf+kEcv1flPOBVet11XGF6Ec+bioQzQnI9gicX1tRoeaz6Ojc/01Czo/Vgq
k7khqmtzP1EIIqZR8A8kPskAuZ8fw5QjG6mE0iXj7GkO1rU/+34QcCLfsb55rqDJzDgDd1vVaiLF
E9V5jhgqRHIi8eXnR+L2SZYu4ubw7y9QIkqbszIdCtKjxyYAVwIejeJ7z00xR6Wle2NRZZc95uoq
8xNuAy7AFQxWlKEekUHGH4jz0GA8EpDgMfDawPTraKJm5QQAUm5gd4UBSQ1XRDPtrmWpHcQhofV0
TGS+xVhXjXyIeU0ZndbEMvCRq4l27MUgiAJ50gDY6wbTI1bNH1SyRq37Qd19Uu3UTIipvHMK7klq
1uBqaJjnMhZE/htuMpj0NFQEP5uhc9llZ+KlR6VGy1TJSvQl4g5Kc/fdluAVJfqo9hftuh8n3LdY
4awG+xz82RRa3LrKA8Q5TAC/AFVCD4ygFqVrB6EmIlATW2CZwTAhepMALguS1ith0rwbZ2x78OZX
9pch2gtHqRX1dbA6kwC4XHy43bzEh26w5kIhjNxv5Ad+sr8sVOWnC2s1cW0zqBbrqf2TsBGXOPa8
o1O+p/0hOOK9KKg3kRKbNZnZlY3acdyZXunwVNwqhWme9xyj94FJ16+lOfEIPZWg6f2HGEl4aTNt
BwhxbA+aFxVjSThI86UHy+M+5BGUNhE+iwIPOgpkjR77JIAmPpzRifL78J5OuGvDZF28wtMTlDJd
Tz9jHCbKsmap2LoDnC+yN2fd/SSsTz2fSkpGwq5M4JNU/02UE7kqugALc6B8ouVZWKV47AmKFlFg
p3sQpD5X4wSCNritJu0533B/rafq5gxmBN2H5IzmkN6V99zOsSkrPmVIroPY7z5OR8+bFocpB6t9
T0lNw9dK+3z3RLiWSe9X6hnDQ45MZGURMeQyc5xgBeuB9RupuAS/cc9i0i+OtQjcgwMVl768gLo3
o34bDtFf8LUU/3Q6s6A7Cs4wQkDDuEMIoAWTScrdaaXqEdVica2VgaUez+t5cVZ1DMn01kwWN6cL
Z/k6Zk4aENpIA/KsGX3MwHubmqNmn0kL3v2v3lMDNJ/5lHHt6RPzIRDMoUKum3Izc0LExsmyP99E
CWBkhoHkeRF3VhGALPgDjS51fSEfuIO9ooe2qeSRsvHBE4Ply63qDhqkY8pKEe3V9/zY4qViNJuK
so0LpE7eObmDkxcFJu5duW69lognalwbukLbDyAKT3RoPUFffGXeHUCyTG0lvPfcSV42cgDBqSWa
Sja9tIcP1AahBH34tcl5fCNtU5UqTVSrrLY8zrEHoVj+INrw6L82zZi4AfYlg0aVUECfjxj2vfVW
KGF+d+VrDYmz8ZYu1yEfJPUWCdP06cGfkFFu02XYCQXfPAFJRqXTWkMn+EGNjz8rDj+B6vJfF2Ub
TJ1EaBQpT4eGO2oZxEVesz+DKDHOs72PmDOhzEHLIRkpn99iWWYwlbNF6rPCkxPFs1+rbNcAfd+H
8dAnoLG1UZ8gS+wgyYD6rJaBWap5165DtJOXWIBZZ96Q/FRaEfGb39jXpxeNTcNWmOFncQrclLHK
kaVoK18EKQOxQkB5awdGTRSmbzF6Af4WhGJU/dpSPIG4kn7V2xV7cUjeXLdgl5jW72jiEU2XQMFA
hnnPYUOh/fwAhgILLNgPNWz8PJUOgMdXrpXcySFroDwl2291ylsQ76IkZGNQKwN01Yn0g24iOj66
FvmInzunivO1MTs897gsUzxJ5vTFruB73A9+QXIlVMfR3HWBWZxz0pOzWPVNl9FzA5L/lTipP0rc
4o00LFm8W3JxxkNElQg6O6UFyu3inA9QB3zZTjrNjA8+mFTiYu4G4+djjuQ13VU5LZYnT0PsBvfU
THrDYrRJBHRB/KcdF5242lg06FDpWLG41ngHfdA7xvXNAig6TkCIrQaoFcHILkcf2RPnNARGUavo
U3fAU+XNmX8Irvkl5RqIC084fHFz6+Ku7KwiAzdCDO0J9x5Q9tW/hFTYrkrgoAjIpY+gOQQOzUhs
ziFIs1uXbI1gyrN1L1eM9+xQJ7cGIQOcZJvUKcOTQdY/WoErnQjoLnluF03tSckSghp7BtQ2ywCp
NTbfzKwX55ibiURqY16iyM7s+jXEGjJBm+aEnz3tATHMau1kWrA74arTwzjyXPxXhdX6IqLgZpyv
hhHiEIf1T/O4e9KS37QZ9WY0T4fZwBFhK3vx7szp9kGDmjk1LmCbVZ5uVnheLoqRGw76IgQ5BlH4
xQCR0k6im/v6cy1USPYCz8h6T4lh7FLkCI+Z82SQpmkMqw27VVU5BO0cd2SCNYhAfblJyJ6lwSwM
l1iyu++ydAJaEM+Kn7gd+O8tp/2/lRwg82JHcKvw3JqIyUc6rkV6GMf+dPUktYJmKto5YyXpUkhV
UFfyQI2Rs4wVOLsq28qpfAbbmrGwJL0HLIjTYXZWdGGTx53FfdzM37Fk+QWK2K4c2zFRKWYKM8UO
ea7YKCMHHdWsOZm3ymJ3OzOPzcNFMkQbRuTzmQHAopQ7ll4bD8tz4+GFoq3+xmRaAw8bgMJnNYLw
09Q+/TiDgdPdgpnjagE7YO3Cb1/FwLaCOqNtEmKleqBGAC6iJQlxNn1g3ZW91AM17D69FUUjmPBi
o6EQymaEL42lpOkUbOntdRWfTcvAzT9IN0wO8RlLZWpwtSkLzeM9NZrQv7VaW3BwzdacWxUIvqSy
l11mdJ/xjXLZx3OAem69Y89BmSH+6cEpDW/5lmsgu51BbFRnW0cbV5kfKZOyIEtvxdtTEfsd3WMJ
t+oB5RsdKoGNAY8mfvAJ8vi0u4Jc6DsgB/mRPZvnMEbZSwRv38ZiKxcs93a7JUM7jTiUGTPN5sr2
sJZZ6EB66mk97oHlytaQbmYovn3aa4iCtakY+kTBGcWfbjzsES2I+fGHNTpWkmPhAGRsLglha+X/
lav3VQyCb4FptdSL1P/OdgPEh88LrIYeUpiyRAfV/xm0QKv6RKF0TXCDtd/xHE1faZuoQHxq0nME
hluYTUAjy4LLvZRfZJaZJEt4nHsvkkoeYzEGyCQI3raXCct1AQH4T9FcO1lNQg0mS7sEeiK33ahr
TVespbcM1Rb1ddiJnJOQ8+J+JhNO9nZOhIwCKTn5h5EJDirGoN7JLfzR8OvhxyS6ZL0PsKSZy5Qj
LQIKniL8sfJ0R6PPhm6e0qewai6Q6fAJXag6kR9JRZvJCjj2J4AokaDfEnzR1zIPHna3pcPT/DvE
KEm5jQtluuSiA9K9aLQ5hfC2uRyYu1L+O5cZTJG2wHd1M2P5jLVWqtxcYD3RmzHb3s8wI4WA1Lbl
0geC6KDeE9PZf1LBIatqk+B5GDHigWSurytZYmgUMZtK+vZmZo2WfvKBMojE8XTNNVTCaKyLtNJ1
r68wTPkqcOhLhB9IBkpUhDsSYsLKsN3zr19MPaGlXEBjwdpew1UZvmkRN8D8eFHfOXcjMeEdF086
MuKmNWyoQ0hTuGgEeEvIU1l1JreK9wt4cqzM8bTgM+VD9ZU9Ce3VbKgAq9fp8S7UD0/JxO5astlr
+COeJ1VQgbhMteD9+VXA7QBr6wr3xu1iUl12thpOVn+AOzTfLaHxDFuoMDHaMwnIWA71OhUNdE2V
9bzIn+I9wyDKoUyH7RbNYPHaJyLFwdHQ4y3YtUHvfrBR3BjEkzK63njcJ2V+updFP98PkcsHXGwr
PMDOwkMG5gZdg2eqYQpR2xuXzu+u9/qliOS1lTfp4IATpd1Skl1tEaewTRiEMKPbqqBpG79sBp3i
R8YibqqAZEkJYp9cvWnVQ5NQnV8NVPEex4SQApfgMrLVBcZ6fjIPfb02InwdpPcIHEuqsjCxrTu3
mNkzUcuXkkuj8jFsl3MolvS5Jm6/I1YtqvtZvDODM+y9B6xuk+47VQ608GxaZY5U1a7RWtHX6vnc
3tX2gFnsz2ERjdzP4Gla9A39RDBY24NBrF/lMgsRfuqbV1ecN3Tj79RXuzGyYADZ1M7MSdUCTtTI
K5bh/W/AaQ2v7AninRKEaQUfproqmq8u2G+T/vtpZLek0eJef0HcHL6JxeZM9792dT5cgJBRTgg6
K4WBHIUwuJ8psjeXkMa5XJXECwyVcroqa7THHByr7XBoBEeeD7nWIAY/j+TOv0OwFaqIQZMUactu
NgnrCsTlgHskJHuNxiKMyR9teRJLKrjL25NwuEZRhZO9wV87hxxUZK44sqMT5CYbovM7THonQKkF
65N8iGRGwGOz5hwETMOiQxA54ZR1Lx7mGYeNsWa8wTtqwKYXtVrllSC0aoVRc2P4QYs7r+vhb1M2
9Wf8IK9+kB8XVAsMquT1k3r0ssqaNkdNXOvTP9ASKf7lCkJ5JVrmXCs7Z5HKCiZmsoWY3irAkl42
xiDZ0PdXx8WAMIWigk01DVvk8Cn7PHMVvRcGcbkUCJqo2Xlskstrr1sN+fFeeUaAhAreyq8KRGD3
1JyYVBjS5S18sLTmjHN/Qh6GbjBbBG0ed0oayHVpjPBD23XtOOKX2T66orSJFlIRRAZNsDtNLIMy
QmXgsS0i2pwvdTxl94am9MxdMrOwbCawpM77ZItxR1OceXzMT2ItR9pbyzzNlNKpyevDCrTBOsHS
ZtrP1Pdx74RDc0S/tvQ+v+jwb1g4Y7qASeeRNWYKK9KFFHNW1IU9c5lSiVAGioPLhBHxrfVzbJev
M7S8yK31XfQGOiZlZuItBjvOV70TOXbe3N7cGHX2xNLnqKYl9nVgH7bUVKipeZjjkG62zeSfDV6P
9RR4CgODv9u49720lTqfYX5gPOxUWL3+MXN5ZCd8IV7owAz/RUUV2EtByn1RybYqeKA9xzDZCOzh
AA6Al/msUa2WEwTULsVkHI6O6BisqgWlVTPsQ/aPW6n9H5D5/QY+n1SjPNu73vq46EhC88iue/Dz
txJSdSnOMrgOyF1bGWDCTr+kRsxGcSSic1W2AxSn4FlaYCKe9Ug9NfTDCDuTMf8XlsTGMqsdpbvU
XRaFatHX1EvaYGE0FVjdqvVZCyFfP08mCK2eMqZfWR2QCtwCvKZ1zUPGm6GIZFCiu+4Mff0pGmZi
1Md6RDPViZz+M+eDo5HGDa4Eh9A6J9avY3NYOFPEFlJ9HVmzHLFaag8UBsNgC9qdFWMh0FEE8qMW
ZHlnU/1wDp0yZzkkxJso/YxVI6HAm1AKvvaxFG5Rr0+YUiuSsli60kmhGJNNAlt5rHqfQwPu5hGN
jNcJdZKiEUzicSp4qIvQfeF0tfo0Im/OE8asfu8ltclXc7/Pzi2vIuMK2uP2LuPw200N045Zw0jV
scJ1+jTMtJRqu7D8jwrGMgPW5WQWSNMPa55to5FCoFQjyLEgnqxupf9thvbWAAVZ0RoYPpthbctV
qqazaY+IxgpvY9fBCke4Qr3hmGm2HM9hlt6DR0b5dnEHFzI9qZMWM1OSZaLcPqqc9O9QYBIdztEy
rgr1SETAsy0FVrRZ/RCcHBuiU5X+oPnBnjL3XiuOMD2RHUWDLdNbvpWqAPRjtiUQUVJSRIXv0lgF
DhS7yzuDMwNZPmaQmB4S44jG6GpzgA1bxgb3r1uw8e1DdyjnhL1fSgnTQvs/XC1nN+MPGER6TKaY
kGl6aHmvUyl8Wp6uvKpKCocN+0nJ4f+i6OLWfE1+yWG42F1rmI/XdFxygDgeKEGopmsjZONBgGjC
CEDa4aNiW1nNhYfEejBI8YElhOrTnjS9h1CZMv6QAHY+jHI8bpHu/2Rcrl51RFfw9pxeHN5nCF9w
Q+tU0XKiJ9+uvJsloEsXmq3ZcOUZYhgP8HFAg244LtNwJUrEOLykikksdmbeHqcm2oh+1Urb97e9
VRIh97m4LAVAyZI287RC2HIfEYsbQpD4YGFgkE4Yy7LsZXSJaqj0+aXrg92oEcN1rROdHyLHbojd
3DAAZk22C8JyTCQl7HIoYcInMrRN7JNCeiBuqU2/EqaA/cwFzCRGoCqUGl81Sw6DqG+kHfIKMvH1
HH91cL55/OxdPLqsOIe2WP4np9WL0qF+s0au2pXhz9DCL130AY0bu3oGujUCK5lFEJC+hbomVogJ
9m8An0ai6bMgJi4Q/KPsgh5a+jXE8e3wmwXy7nA5t4Sqj2TWqt6mTldBlgW57lRue/Isg2gnJuwE
zvphG78HztzhoNQ0RKU1Az1lQ+Wtdkt51UO4XhCP2yNuBV4xZ4zYMw0bMhGUgcZBXBHIyP6S+xW+
nCSCMeE1vks2YW7O20hFby1OBAAY3Ax/a6mV1PXgfEShCKPIIo+rHRB7f4d2FKI62Ujj1J8RJPps
3E/8KkgGLWXgShSm87sVe/o7tzQJqgtrQ8yxuc3X3ThiE9TGmWSfA84xD5OmtenZPEeRk8QmRz+m
aEVeFtqDpJk/3xA1vsbSznsbSZsB+54aytHEfa1EDtXArfjHaHnWHeGfkyxxh6/oX6qzLBXgR/D5
ywUsiYI/o/5tRoRAAj9FQvyZjbdnfnmhHY+vTfsoBDNtzkkWeY0cSIE5k/19KU2b0XDeBwBgspCb
s/q/1OVedlZSdYhA9kt35ZLDvZBDkE8WEtd5LtKx5HY37Y4ljmPg9EhsFaqsrWMF7SsVeM15Qzyq
rolTGp54jN0ys0+xVbJENe2aCYBpk1tIG7WGGeL94xTsCIShAH0d8X4zzsmqRYzuZh8HL/2S0SrK
YOpfWRDBU2DEFV5hkErm2iZ8lMhEm3UkxrC2EIXOFGTZoVmv7jphAsTe5c/3Oudv7qk+8ZI1rR+n
p4v8Ytd7QSKQ4KYhjbCPrUIc/B2pnHO5WP9r6tZobRJz+hCCB7WQM+Uril5shEH562FWWEjUgKw/
2zD5uIJYTbzAptSs+8iJtmInZc3T7sYycwJTbeoXc+u8PEOZVjyIGQQaFPX1oBp2NdrRy+lM7tH1
yoMpagnbDPoBxcpn91c7ADjrLP1LZ9NVMe4FnyxTgnyT/lGDhF+WEDqh9wq3aJdlkNUsWBb7x9JL
VuETdb/Oojg/Qurt8m4lQEfjebNQtPkv2lb4Q/ylTRH+C7EurwOc4ldbjAjztrAJwhedBkh/51WN
Hyar5x+5xM/BevU/qUBQWhFWAGgTjR2H7v4S2bzjMVDlvgEz22GTyEVB+3RzrVQj/KWzy37OHWZc
7UVf3QhNPzXcFaTmebPy4tHA/S2SPoZ+fhocLEPxhBHZbyYppFE8J46m+dt4moGjoOSQntFJEBL/
ZFO3vxOgnfSFkY+Fd9P8a4UajdvThO4UnUFhhmPMX/XEpEcFLXbXy+V4Bx0rgZPrCA+rmlplzF5L
MnC6X4ZvIN9YLXuPODDagZnWSXr61mvZ6Gc4iRvC1mSyg3I1hw3ZQHBW7NEliy/dOLa4VyrUv8xQ
ruL5VfsT8LvQxNBsz+wwCwvp5f5z6lct/Cw3VZkpTspgnNgbWinL3mvefYbWNve41H8/FgxlJvr9
de1iD5KAXhgrqjRzlZbIePR1SM9y3eWhPn2V/hwmkyy99HmhntXHrHizPXruydn7bdeovsABmjYU
SlYyxGFkz+Q9q6fPorAIDieM77ufFDdW6OV5Gx7ZSeQjf53iUL0zREtOzwsZvaZxOrBohZdLYZcm
UwpNdfIdd2l7+Khwb5p/7/NqjaY+x2PFRgiIvuVrWZM+SavIVnusVmNtWkWMxZEG4L9x5+nnaYRH
gCRviZBmOO3qetKGhrErPFm/cGe+TBMiq7S0kVOKHHrtMB9soY4RT9JqTUUsL4uf2NM+Sslw28Aw
taObv6/XnOqx9qJYZ9BJZ52zF58qmRxjNBVg4lPh2Iwe9VNQyorEAoEtyLw4Ye/M9jztaRAoRbc3
jxC7/xycohPSK4BErKAORumhfDu20tALoMrLf2GWY2ZJbE0xYWuujFCTYhKrPwPOKYX0NdOpWzx6
xYwAPloqMvGRQp5txgE19gkns6jvY+sXCkfmvjbZT2ODwNpLWdhtYP/Ood5z+SXjCGaZLzlQ0Xo4
aoinZIIqc9WCmgC5k0WBsV5FlXKy//fQ9D8atO75/2+aKfIQxPp3hg2Jnbpb6YoBlW5cWtiMO2Xa
4fbjxj2olBbcNkI/p0DCgzhZbak2Kssxq5ks4FyNp+y+DdPEC/7hkF8twwbdYgWwEmjin2yzyewo
rqxb60WyGO7PQrJ4HLFV0T68eGOwcWw6HF6w589IHPL1RBZzjwnHzvCXOJoZzUjShvBzCWe2U/33
/zEGMLIfQdcJ8pkct7xCNyiZL8uNB9Go3DwkkuOqrK/bYzkiGnY2Ny0nU2OCJoHz5JBs/ihTkjVa
oP3FI6QNzR1ibMBkejEQe6OqHxcY+3h9L0EZ0ov161YU4/Tu0SWLD1LYlrHTWw52uOZ5USqnfVxK
vRGO+kKuITudJNVBC4DSkzGk9KxikPybF/CftOP3Gau2wH12nQW+JxnaGx0Q19BWaWzMEJ8PUK+j
oScMd8K9/Q4t/NTZVwnTJt+FkaulX3xDGhinrjI8pHErIqbN5PJaGCve9CLxyIEcaLEUGSFifH0C
iTKWZWIGt2N9za1G26C6U3RZVeoYDYfEg8NUS1yyL5TImNwABnOpr8syyKqx9Eci5Y0sH4hlbybX
Z4g3IRkexwEP1tq3EqL1fDaChI3euszlaRKrv5KZ4MX07ivFNu378g2ktVydTFtoHtle1sEYuq6Z
vNAu1CxFfMp6Bt6CCgbG2snvS4hB5io0AOfeS3x8v3iiImjU+MgFZZUnwS+OW7HojQhlrZKhHk7I
Z4iJMOuAfxCf+APWeLZpfZRvX8Hl00PsvGeEcAjYa5jPqxWPsMr8amTSO86/nwp/OMMnE+LSOVhZ
RYYS5MimPQfcsCefdJDE6OUblp23dzyUbS/wAtOLU+RY+NehGKrGJLij0Fcdf48D3nMtfnds8ccH
itgApVDOiUqKC/8+OwxDKjELz2BKJ4UDCnmnO1j5FYkAxOMj+sintWgyqv7dBSBskfoZnnrXQk+b
gSc/ic6/tN8TP35oiIF3ByappPbGCYWSBO1JpoySyrhTn7UiGqBrCcLyJ/++XS9WYnbbyIysmV2I
lK9/tbuosKo0Krn/LfsW9SjDEfSGmg7WobpfS2eVb85POTcPYw2vz0GpRMqKSfOyrJkF1BTjWpc5
i7boudT9NFDjvrUL8Dg/onGfZMmYNnhOGkqVDfDUOPmkwK+QnUCmJx8jvO2ONBmN7dAZZxbWo/En
V8Ptc9irYLGOVLaGn4T+MRukRzyr5VUiqkl37zEjJ999i07+DHS4/Cq8g86j2/Aq2+umOkGuXsd2
8e6Was2GVxGLHB9tg6PbmemB+ilNQrOGII2I4gIc7852Hm0AQIXHvcIA7j0VJYTxROzkVZ0BxmGO
ZzR/oQCMOzDVPhDmF4JFcPfJ9kR1OCEOOcVqhznNsYETh05DCfriB8LF1m0Z+jdAr6RZXuy7Uyg1
zrpSwlMUZS933fWf1JJflYTEUWTQQypG2j0vWaYP+PyIk0/Wl2NNl/j+icvvgMA67XL0p4soCngB
u+NXTc00GM3osOr5H039aR6W6ojFut6pa0kIAljztTxehjYyDoN8Kc0TT0HoWCLA5WTe3mNpCMEy
iEl5D9sHWpnLvginIA11nMMolIFHNI2/Ctsu1UAUPTaYL6kXuO32P79smYZSe9ZRZ+tEFqkDdX0A
e7HEMKeHkCV6YBwikQuTCWG0UhjK1khg3LtA3jkOgR/10bxkShNYLBrNdkfxM6ge5Xrhn9nH+Myk
AiyZAtAInKNRmycmlgT6e8417bDiVoN44iCLFimwkF5Erhib1FhmTXLtLKtyjTVrwRHMwM6bsQw2
33CtJVfxHoUHP0nQPfr5i2ncDQKozOZOzUmcM4XKObJbaWRZQiGOH4x4pEQkPKl83boKPTacDubK
v/zEPNwcN/gb5MGt8etIbm++jwQdPyONyUbDDwfBd8UIIgucqJvrjCqWCUgU3ZzlGpH5poljoYeu
J6K+qFpcNuJH04EM+ys+kvrTS/6JvVNsZrra3id3d3qnr0jireWMWNu7eY6asNyurHbUVvN+MXKn
Sx4WUY/yWazm301GrB0pez2k0HAR3PBfzlyPI5VP/MHmdrQg9e7dTJlJlJws9Ur1qlIkN721FfS9
uEVNFEtMZQt0QEyy5Py6IjLLra9Cg6vYTBALfvyZo4DRuWBQf6yWOk7yOqcP2lGFSARUWdRSl3Io
3Zab+A8Kf7KAD7RfSKTCO7yT4+P9CP+pLQyNDb0glU+W6XpjEwfW/g40AZ9Yg5FUncJF97Njh2mf
BtByJYTi7dzJe3+WIDAQtid2ZS529HIZ1nqtXC2lUSn0I6f7zLxqOCtYgumCjC6uU3pufkdtjYR1
c6tkLPWw60me3nu3Pd4XnSioaE09amG1ISoez01abdezt8lBZjmfKHLJzkzhFfvWnMjvDzHLR/gT
VlStbjTNO+mzXLIhE94IDpkVmTq8zZYKPhTeaTPBEGpkcHI45FnFt8lBvOp2sW2jAgnPGBVPOa2k
i3k5QS3ohY9/hTdpSp7R6pxMSmvnOJ1Fe7j+ZAMyVhAMzcY7wlIbIvhKi8UzOTk4LCvVRxGSFTIq
w0rqDR0jgzhhiF4lSlwPqquixqexYN7my8gRfas0bzqZ6blbfMcgIYlYHzY00deKBvK/6saqr9Yj
hzZjMQmRfQLqTa1QKZNF9DanK0Jf3Y/db4YhtucSVTUveJkVOLjQ3M845dxgUJ1KbdXfgBho9bYq
Y7PI+Qpt9bRoqO4wgXLmaoeGSBC+tM6UVN3ULtlZqhgKWKAJZ3AAV4oEXs+fjd6t87J7wwLMxg3e
Dlrigkhj8Dy6tH/odG3JiuqZzLE+EpImmiHvPuU1wFDYB11kDWjSmfd8M8FbOZmaT9NhQicbWos4
ji+z4JExdh5y/kYWNIfpwbC0Qh6C4pja1fWGxMijtAiVX8PZW1zraoBixornls8dBIc6Ax5+9gt4
9LOKJ+X5EnE1J9WQlL+igAOH3euAISo9FSqmP+kh4fZ3YuVeIipWB3o3bXVxdcyfCv1ZBC48NGN3
P/GHCoefwMtYX1boUGPEHTzaMeroe0rPt+rMr3bjItaN7YiiXeUlLnJulSRsB7AW2DK+BB0wNfId
0JeZEHBKOJmj8NQyqgU6YBVndVGa5HrRUIpHCm2A+PSagCkQVoY1qtgcKmSsVNWXPM5yV6sf2WrV
rRLDV8FLq/tM+q1N393QzUaN3NzNrTdfXyiAzK1PV07zxit68AvBrEBhb1tBCaJYnGYRtz6048ll
qyjMenGKCHhMhB9LV1ygQcozudJBaRQA0HoDTpht2pcfQNbWfkE6JCDD1ZbUz4hVHCyt4o/PA5UV
tliCF8EFYoK9bl3uDiDBLgF0rJczv6i27U4U0L9hnhfspQlSx0Rv1FQiAfJt2ptwO29cO16EsdLg
5sbHIR9k67tFDTslUUtysMlFByhRTVxn9p+ppDCKUGiZlri89l9BHgLKxz4cJMHWEI3WhJsyxv6m
LzZMLeZOQZXaPT/ejh7Ul2NPLQS+L7IgacIqOa8d52s94orijFlPDliiaJupY+/sZ0axO1jezYFV
7tuY5xG4FuLm8XeRFA1HtYvmixztVMAi4TQQ07YBUrAaTJiaLWOUVR7kJNFBBvqgfFn+o+BGS8nR
yy/Bkbj0Man/D8VNlNw2/fBxRM5JRQvjQT8VaAb3DstNPORueS4cO1S8fzgov0BUn5FDyjiK/urL
rNFq8BSbirCWLR7XE5P6EiUcugHKVQKw87v5EszPbl5k/ibhEmqqua06ZwZXlZifsNny1rFljSE9
KXr9oR7HMZucXxQ1+qr8WQ74RB/loLK2fvfSfAgp71NoS84++ZcEBjDi28lsijM3rLgaf8EgtrgY
UzlrtWbD0uzyx3uW0vJxSW1BXMEi58R6ZnzcWRXg7BAuqg16cZAElDyvXp85k+2xaqdFQFj5adoT
+OVL4ubHqZjjaDRnq2jHyYYrZsn6VRVioLatUNLSx2yopyO08xubF40v1Cz0K9qUUcCaVXcg9PG9
wp0mpxH6I+qO4AJHyAdreWxV7u9L4KB5KHTsBOydtH/YgEXOH8mffpY5/lDm2mDNY0xLtYGb91PL
vm4U1dF30klP+9RngYOXthGiXNd/eLRDFLG8pLBtDnmsVNDj4HAQlVIAtWE9UYapCERH/nx/PoRE
T9lxehKLCswkuh15SyoP49Ni4IGxUJvDBNxN65CBXZL56GYPtp/u9l6A8s3yFat/ecFi8zbri44d
X8Ou6hnzrTIvD/4x5do/KsJOSA2+znet/MIA8SKRK6NoW79uHIlr0RNK8uzT7AnDwloYvw1Pjjau
euWM8H0aDk6srYu8eCW8HkSM/KOxNcrSO6mKGJHiW1ZlO+B68hcxUi2R5HD1yPnM6HOKiGv51IT+
aFKqUDjZrDRL3d6DILBP7FP/x3+QjDYsDAXGoxZiHUAJnI+fxiNAY5+EHDeli9vzJmLXT3amJeoP
LM2OlesE3hH3EhzRoFzAIZ9vIQZ1LTRZrOj8XHaTyhd2CRhN0L/cFn4570SukmUm8AN50W/SstgL
ljy5iiP7VzCia0S9dJmitz2otEZupi97Nx3eN/lCH2eUNa8/yxcZQEnRXXoJPjr29/j5nH7FXvc0
b5FVmnUrL2Df5+wavUDvg4DGrdQ26rlXdA44hBQAIqKSXEahX1bglbSX29Z3UGuXgwNA7M4MWBr+
oY0yWmCMYE/R0QWo19qYj8GGowEFwqeY7gi4WOUgQZ2Dht+P/5/LM0g8E/FRgouR+RfoQtq5JKLH
sfkwrEXIjLZL5XZQvGYaxj80BezmXj9EqZcndMAXnGk9p5EeiWTWGqGFzanumxxnfNf5Ammt1fYK
7f7E182mfUtXHpW15xVzGOEvDa/hRQoI1TvZ60N2pQBis1BIXFIDLMRaCMTeRHMn7S1Fdj1U27Xa
evaMtsaSsGWxraqStNe1mByv51bA3heqr8i4w6gDk9iZsg+3N13QcwcLHhFwctSYrBYFsU1UEWyh
b9cFJyF4NF6jsfzQ+Y4pM+6jy0dqtZiFtBWEvWXQ3UZ1xWOVVs0UOefyRCpgwEJVTtOhMXFGtJCe
tmHe1EqutV/pX+vhTKVzD9veZNB7iQildvevp1yJBbyr4RJaKhwcTnhwm763b3zRVLLSrrMTUq/f
V57s93OPIQKUVLcNCGN0BryrDsMwnomX+CTuUKvxSdjV6trD4vOAE2Pmo8ahyGgjCXs2ltKDY3/e
F+dOqSlx1qNRbLcUWqLGBkOB6+uaxQf1CBqxqq7UIWtQRkrWahZsjLRYMmuS4ba7iIarZ9+Z7KpT
keV0TZADinX2Xmp0Uq7iK2K1/8M60Jv9WskrGWdq4hTnbjeeYk2jFafejYFIKVipBZ8WIBGMaZt1
X2cvQc211JlCeyodIyr2+5RGSnPSGC3YdqG5d8yTIAz5MBllmURP7my9XtVY5TDXIn19+Wd1SyeH
cWvIWdH5JRn5STflwddpcq5HqiX4DHn5eawPnY3S9PcnLrUXj+7HjbGDBqbk7Or+5RdF+uuXxNGC
trbrrLIhHTyQgus9BVoxhVVW9uX4meYEbQN4BwSVKRIsKQsse/0EDVFMgzMX2yqRN180ObCbwNbD
m5clJaCA7rwnBfRppNO+RgzVkBBaX6EOjipF5t1FVmieKVp5vTLM0ATI1yCZRiddNZPKq86hTnum
vgKd9SkVCkI186PwdGmJRnxQbPaYw3dW3R0CF68TL+RQZZtI6HA5adR/h32jRh3YJExb9R0r1siu
ipeezGYk0NjOwdSxRXRPBgoMV/1vNog/J0eKXV9ReVqgRollX5jBrgZ487OTkt3gaGRoFBNo5jvc
23k691p//XdElhmvfFX1AptIr5Cw4H2n+EMyUxlQnI2cpDcjz/R97XrSu+eQUuR7xLFKCfGRblKA
IVbnSVzQdaSg930PdAFXW6yD4mFWsGnihAE4qApMwsJ3VABSqgWeKc+xgd8uIVMa/XdQGp1xOJA6
jt1ootA4CoOmz8VwuL6C4LQd3tb6n/M9QounV1qpY56FFRl3njr7OBngPh7/2N2iPACkIndRQMPq
YCTKJxIraR9RrnqHj4R9j4zi1xBiX6CPMdJtyc7TVPRt4iz+S8qU4DxOfdn9Zk1uHr7ISBiDSXTU
mWGrjuE6JxNIwZSzhYyC0OBo5y/uvV7wp4D8OXj/GaPqXyjapBQVr/RMnLb+1oXeLL5yQiq7xQDm
2myv5fc8tu8mFpNNtw56fq0F/FqExZmmlgkJCSn7tau5oWr0U1XKlwI6UkcyaqAExKZ6vp+w/7dN
bx7uq2uMTAWmr6YzqLatWnM8VJMo1Fc+1S+O/mTwdflh2mx1duFrLShsyTSk8mEhdnhj6Eh1dmuX
kWE6p/yMUvsA0kEWDsgClRjvSyIUw+/6rXane+f1alnb5wUO3T+CoPaRdRhoFh3ISb3wzdK5Ge9s
55CSB+4rKnt1i57Lobw/LeKzBBILSwkMoaDv6kggl2IQAuO1/GKDgmKiLNjkUP4hxobUz0e8SRhq
kNtfP16W9F3MBLJdGq/ItP+2XrO30engiA2ZB3/6JX39IKkSytuYeZ1waELMvdhrQWMkuRx3uvI6
/xjs8ojrRZwNgD+tYCfzgX8GpfKa7eMA20yzw9BEmg8T2rnWCGQNxajedRqY3XfnNp54Bzc7r7+r
cSFvqbwIEWyRv5NSBBDPL3jrGRxyiJUkX+c59ghANiMMhHeFPvg/K+30MeSZl8h0yCP9/W8G77lS
4P0uKO6aSm4bmL5fRcHjb+s8vi8tDnA0BHN30RuipRs7qxvmtmgRVWidkKoWtLJuSH6+D5hHWAgX
Ndyx5SujR/Qvfca3iupIt/JEUqr79oyg7Dvtx8GG/8d2P/ynpjUOWu83hFRQvyonWPm0f8H+jWMH
CUMkLsQbNgI6VHtnmdD5O44MiDrerjpgBiXcjhLz0adu7uemcdpoZuO7qRExnz2zGivN8lpTG6Jj
MGd23yHymrv7HP5LQ4JXpBAcp5XBR6MRKVBL5mLhA6zcTfhgSSwfifoKbrbYOWRjgpTvp4wuS6YB
LYJukdF9eVleFD3PwLkNaRbXUie5Z4sJ0Ce3S7F/L47PclXO9xjv50R6jzfrSKSHZ52f4F8FZpNU
c1GVbCQA41/XtLCtQYw+deium4k2Tuy5wcIBC4cqwg3yaxIzuNEOgaXI1NWZj574ArSHnsA1BqD8
u5cj39wPR/xm8RswyzFdYyrMpPPbRCJWINoIkKoamfAqEW0rV3Dv1R7CSiIYjTjUVBtktf1srhj7
MEvIt2XG9CfsHH+a/nr5qGza3v38E/LYB8GwM5uFBDnUCelFXi9xkWMNv+WUPxxphJ3UwBY7zX5T
weBdhLj/GxwvFgIfAO1gvaCNTPnrLxJoWQCOh5ivRKa5VuUKdPzLNwDtIoQpPdKo9qzkr6l+FF86
EHTw/I7tf/T9vQXX8DSB+YicH8xQTIWR8OFXSM9hAme5gAmsU7YqBxS2HeEy8T0R9ivSIB8LVPv9
mEGb6ATfzmBi5QrxalVjLOgzujm7t+4vaE3wYM38ohRSQ8wIqEaj7RbGfCcgrIXPl09q4jIL9q+p
ijn9K0NKCyRuZKjS5V2nYmzENBj+q3zT7GDT7MnByLu7qBS3KjFDy2NflBOj93U/k7jVYReuiV6/
lH6eQIy1BUY47PrwLgBleJigPG214sGT32FO2y0/ab8afSPd1RZfhvB10JDbJj2HMSkXrMusj2JW
tQvqTsl7ed6nrbIZfpvslA5SeDqkH8I5FfR6WmDdyq+OmZn4DETp+y5UHT8U1kIR5xK26Nnq+r0/
hqPbSsb72FQ66HJHHCYrmfAATtrGA/TNKq4eVLcHN2B3xqX+Ucd6U1ZRsA9iu8SOxc5+Sre9PahM
vsEFDVpdLDbx9Y/nb2kM9i5AELTvPfCA6iuvxJrdt9FLP9BSJ7Kz8pirC65xzai/tMcoPnRfJ0Ro
UVqUTJj3nHvs9ozlrBGNXxGu3tELR5ciC2TJconT1toN2TDg/5VDFH3MuJKx5JuAQd6/GX0ZvmC0
6JUFGfiyehFMS7oDmHdluAtCFjugQmCfQwqATlSAGOVV8fPVqpaKu/DYZl0orG6J1AIwJ7Bl77ZF
4ADD4LVtbdTSBPp+jlboiO0wo1XntQ1c51wikdoO1QyW0dcsDi3ZHHtVkk57K0Qdy6gm/rV6rhh7
2vgT5SovE12rOjFmJCcrmqpEf/xaaihQwFiAF2UoZK+Kmi495Bw693DWPc2ceFEVjYe2ksx1Of92
wjCuGlnTh9ua2HHEfIBsvTJo4rVVqEdFSqaeefsj+STvLgLsf3J7M5PVHhe43VBwXwkq8zGV9ibY
jgwJxicD+eNc5hpmYosC27qgzdAZAr61OwSXOxZpPj/lwBpmbbzhTMuckVOLxvK2afgC4jj5m2dp
KAlqhfw+vLwQWUsCLPF+/u0cN02sNOHXAY9REEiGe7z5LkfnpbOFdTKlEFaXt5HSO0rGN3JWIlmi
OlJuP9rBxo2sUvJmLtLG/a5gfycDDhfru6XDosG2L5WxHk4ujdwT90q5qG2+98MQDAcoQb3jE7tA
DmccYpruzVRTAogHWI3i55xu3I8iNexeWz4fVfSPc6n9v+gndUMMMBMGsyeSiAL3brF9yTY8cY7z
2QMywCvWMDjMCg0kec7p88YOrmMWnMc135Bxom9921+Fdj1Di4NEyLDl8y/eAVkHl5cXQg1oLjf6
a6/sF7jqxdSOvJP9Vih/oS10k0/60NUdRY7aKgqVWgJz1LRJLYEMGGCmmswGiUI3gMinlKKhOvec
gN1gYOTlEE/DHcLblJnSHs+hqWSY84f8cGQq1LwnMOcWqVeM/GE323Ah+aRKds4rdTRD0Ne8+NK6
64R24TbGjcRNvZiZW2Lq49MGiyFWXl+KUhh9etIcFTq6HYWNH+mfUbvL7eaSOKNzXJvOyW89paN0
iVaOssBbIz3ZnHkKOZ/CoSjkFLmioqb4TW3+ne3W9vzW5KTXSCErdw/CDtGdJoFpPrqgMMSWxrpL
lmkoOLIgyYnj3ndOHp/hMfGqKSAiZRvc9mdbGGOWSArsHNH63q3nD4FyWB2KSxAka7sOhErvupBH
ybt2mK6/vJ8AmQN7833jSU4yihI3R65jW63q6Aq6TPA7HAPaDHJSOXQ0OX6z46+2k5h45RTuQiKK
GOgNByPohkwpI/pdZ58Z8rIFfTLuS6+PllOIu88KlCYFX/njI+XRPEKHpZL67us2YJ9DE6wnepTY
VejpodmrVxoQi2KkvMfuhgJaQm8Azn8jR3+3t7/wy0N+rhY8EarNOLOVtOVBvhW5lyPsodXmjtBx
edVAU0/zoXpmQu5Kv5LPZoNx5Dy+VsCvDE74X0eSctieLyaxXRSjqyzyv2nBQl0XD52NxCOIgnu1
Qo/PZWY/pegP2zOnbUpGuRnPp+iY18nfwbU3UiFBnx0jdG0uVcOjgsbBbSwGMEZQISOLRiJ7PGpl
ubW1Qqmr21n4kbiGtvWC3MgNEZsBPhWPEgNYToU51g5g5TASLc2ZbySmatEckndYc/hiaS1tZSlT
JLgcT6heZ8cZpcv3A29UA+tE+/5JM9quYUhMDUvirxu8nN4TQjmJz0MsZta36xrBMww4MRwmpp75
kFqSf+YoV6Ov1jtbTVwqbbqrnRcRCLB6CeMe8iAKdMM7vCyqq1S2lBVd3JFhAuEPtvOABcgic3Be
LKD67M0VUCSozLNShT0Qu4M1/BdLsqTY/HMCqZvnBXw6ijJPSx3rzCKPMAxvfqV1xOq/C0GfiuBQ
WEmLkDuQ4aH4jbjWTmUUdtny+ZsfHwuVSGsi6rcqRGMG65eIneDgogECJkwaT7ZB0IGNgcemZe0c
aKu0jyEs8sLR9/0Py7b00q1hbUeAEM7f9vKzYPQ6jnsNX1M/w13wFPhB5GQ96aV3D7LsgnGKBWSq
Hv8XAhmuAct78AAOwqQnwpMn+UfVcIrUxkGzVj9BCXN9stcLGiwNG8NHkn7q6Q8x4Zu0Y3YxoB36
JeW94n1FgfbyogF5ArPVx8gEHwoB7yIY3yf5mnHjuJCXVQeHm7qyEUMki7MtENZu9zkcdHxlqUlh
iGjDLoRWIldsjZHrj66fNLlVWY73/eF3PeJH9k71ekytoNNGBSdYRMLEKPu2LT4IAPPnc/+FrKew
mlJ9+lWdmTrUb1LpYw5cDZ+i15mWgRdmsoNMqOcndoqTJU1p0uS7XrpTOw9kbJWRYVUxozc31tFz
0+NMEXxxRl9etI9TxFC8OvM1stuOmVClzyD2zRf4FKn6KM9MzSuSne7t3V0mePpb5+v7lCyGmb4t
LfOk7lw1E9UiuUNwID3xbu71Kq8qODwKGUR9uC0PNB8UChUwRUCT7p0cLS685QhxAes7ZmqXcDx7
W8cjL4LGWajhJr+hVWSTlDWwBNPk1Rms1jGWmW/MfT+7vfrTKgjA8/NW7HX+ihX+USccplKibalR
GC8T1XmyVpsAeR1577FdmKG3qvTIHptGxDltO0E2aQbCYYsAr20jwmVkG0pMSenwt/znb42l76Ky
j2ZnQENp/IIQKzU1O83AaS43+5kuKAJPEUp5kPxcXw3TfJpUjgbWijl6c2jkaYLuDTl5s40Te3qn
9bj2hlb7DPHr0fCnsxa845torPIQ50qpMF7pFXM4OIcDjfAM+YkmFuKM8KsMEZWReScdU0fYEFTq
HZmnrS3Pq/yEp08S0KQxCdHsfcbbzcS4xJ9er5TvIMxmXR+AyuLvQw4vloz6y9XtEp6wHpesHy9H
QZvlXqQQC/3ztF0eGppdQ6yoXv7qwwWo48FspY/M0P2VDFmfc1B19mS/N8eEboDCW2lZbWLqIdg2
m7iGVLO3EcguQgwjMj7A4FANmxXfM1SLpjy1VcPd6IGTSjaRWhuE7Oike9jvQf3EYtKn3O0ZXbUo
m/jNcGiYDPc/4jnJ/444N0gX+fpeTn1g8FaOmvIScUILBlvq+sre1jZCp2pcx8/4FojOLAyxa7pl
Oz9ygsDHr2vu9T7irX6dIoov2fcZGt3ZsTsakZofstkwbq0IcwEdqpjqe0BN38M5MMUkbrxiRIMa
kJvAndGy3bcmIvwl0d4Ya2TyfGDgyrVdWluPQce6UQRk0B6a2KPH0o3k+a4RaKVloX7SY5LMkAj7
J5i2opnTJxXpiMgME0X3XfS921JhCBP5ZELoCWPN4aKHiLF7CZZX3G6UNh/SxAYSB18IFMDdmL0T
onCjRHqSzgubVMB0QM7usL8Uy7NInd9jfjVphM+mql6IPIoBykiq8ymgRJMMczQV2t+YWLXtGLWY
muvn0hRFjgNIbfrjeeCUNKbp35O6U6Iv23QNB6dcHQTa5fgP38F025PZoNsed6sjT9fjAbDrcmHG
kSgqbZ6OiQ1ujXyBIdM4gwuP9pJg4Hf+Th0z1Ijbr4r5yYYDmyp7BEQQ5wvRiCnDSB6Br5BncbSo
gDgAcGrFNhNoyFFNkeBY6SRyUCyZeCh9WlZluy168N6hAB2xDKhuyWEXfdPAFw1P2SI9sQC12Gcj
LEjVu3SMjyrnXfXeOIio6Wa3ZHJQANiJ0jGqTyIaJiTRo+L3Mv2yaEAkhZ2Gqc4JyqyImEcQL6PL
eVYbo0E+FQSko3fINPwPhpZIod0wTC2xvWUmi3gIK2DHdABnbTq4K4bL8LXx/EvEHqZg4AI2/kgz
k1Mn4gvcbo2Ywr/jstzMFym29CMI0ThZQisS71wW1nlKeIuast7ZhMkErCKghSJcPYUlWTIJbJeQ
Baii/JMXy+vz5Znh66p/EcCihu74y0Hl5mYxjVivSNH+jwrLjUZADzpIb9DIV6qskEL6jXrV+dd+
1JYMoXAbT8AGWWTHgEZPqaxv6IJ4PTVCZ9k9nJD+ih0282HVZrXsRNd2rmh1LUhcfiwTKaxi+oFn
phJEgg5Pw6ttgSfAsJjWOnD8OQ4qow6cVM24ukCrBYT/Y3gec0qSXNns6qghQ7OfKCpbNgwjarlT
88I8WGsH1LTwBUneu82yLDv9YhPtEDUYwZwemzQU1Zk7I2XsiZ3WESFj4gIsSKMGR/wyVEbiliX8
L9kjTeK6b9DMEeQir+UEcF28465ImDST6gtMGb2aSBJtoP2/MvCMDqu/TsvY1nIzUNpIENr8pf+7
+DSMXiqBhek11rdwiY/tMO0a6NSsqoawx9/sjr1RaEKh4BvfR2dW6RLglVmr+doMoYHrHw6SgSKf
1sHczXUwObizhsl4rRnDdPSwv+yJzPRzZFWYfycQqZrOIMGl2I9LYE51ItVjHNHcwTuWFDKsZSHA
XSw8iXN7clV1gn+ipGljvbFKx/wVd5xpHGKOFGDM3/QjO1H1wwR5v4XulOML+sZFARSf1Ps1s/XX
3Q9uJqtrM1YAmnqkWlnz+oNnRVy/2jJFNSt6X62fNAPebzGXVy/vFeV9OcckaBLCnO5p4x4DLoP3
3gJecVls/9FKyVCW7pZX270xngfi7I5aycXwd9FC2uOSb9qyqfHAdQeT/y4yzD6E9JYm+lodTV7X
TnU+CZsahz4Ycnl/EIf/7SYPyz6U+cAq77kxzm4GNJ7xmQOENt+42NiFDZf5ZGbfVCsdRmn9tReW
qY9hLcC6XWqgm4zJD86WrKaYMiVgri6n9R/5+f7eQOVw1L6IPc59F6cfZ/3okJ/Ch+WKSO8gOtxe
xCDQfrQUgIr8Kg40S41M6bwk+/kl+/+NZEg/WKBO7e1Nu66d5gH9AOsvt+HVpJkwNfZs3mKCGO4c
Lci3suhRaC60DKaZfwe1ZEbCnCK86q2y+EXTx+iWo0hDLIQ7STbo0A9FKKR63UCapuIbhcp8RMJH
Nh3FCxFlbNse8a6/wHakScW2kwMGj4ceJc7HMlUk3wIeXWXjjs9uVeYBaQg8AJqHsXnsK2mUtg9f
DgeL7GjF4aP/gam5xnVoQ51UTjRdQwU6nQGUTcHFMuEV/o8YjMO4T3zuTTqjOkbQigK3oXmX3h7E
EReet9dQjOyamJO+wqHO3memoHCsahSRQr3nEmQssnnqlD0wbzddXX+/b0FbAjejne7COdifhRGh
Qf5Y9rFnN0qL+/x4e7NIxra7PKkw6r8VAMj8QlsKQLItvpu0BiR5XwXFELOAtHBkosnDdqlQN4uf
rXEq43HTRbR04Za4UKdqRNjRXeWCEW7jB8CnR/bJU3LtSPpHeHxEkh6qvXVZ32SskOrj25tpuCf5
N7lCZDOMFX1DP3FpzVkOku3HoXThGqUZjM6FL0YAh/zE+gu0z4opJwe5Qz2miIK1Gz9f9w2A7ics
vkR2Rb/zCK6daMNIt5xPEWeuvyVCvXMrUhleC3DzNIGaLXzZj7VYpBgQrsXA0axajgDhTZvt4V2C
oXAyCOAIYi8m9CeSigKHEApEyW5h9gDPKwKBu/7SGTpDnSNhZGBLzE5NPpby78bOusSol7S0sNQa
XVpS7jrJAq79GFbulNpd72wtUywTl+IMyHFpdnr8phnOO1zTaw5ZjafFAqRQvuznvZBIhnL15S9j
4JAbefBRMJY7DfbMXV7szCM9Ast3kahj33hvuheVzNnd4Jj1PSbg01JH4qL0o8OMtaKS8z+xKDVG
x0XA9mfyQLHUfO1hMB+8nOn5ZFVNFN7hBnu1PT4mXYpQQpXYlsxNAA7Joswk0lTmUt8mHSKi6EN+
N5sjPE+7Bek1AcHd9EGcO3bFQzQ3AVub0KAtUFafRaaM4BBCDfVS76CI8bu66ycozE/Qxwr7/rXp
mqWXV+gkdGoWWSiW9EfK5AyFuWz5uA/TBpcmNO4fqGu7lhjtx4QE45CMpri8aYTY1VMqEW4jV79p
z80I2YYzsqRnMMl6PlW1YW3hTwmWjF5MmMTGxuXwPHa9eeMODF2NbwH77FqQTTS7oVc0YKY/Eef6
sLHcqDvTzdq/gH9crXG+/h7lzVSFcn1YTuJSa2XPHEBvblMzCwdzwzALXnNj7fHmvECJTJ06i36P
rxu3oXduSHmZch+5ozGSAqu57/ZRAs4Vj3wOni5sY+dPySbLfagHLGcXnYpFOXAP0tlNaAXebB0d
V7sF0wBNIbzC9Udwmp03fvUnmQCfPlfgjF1tMIE12kCtMTygsDltWByFjdCRKa48681RsjUypBlc
SE5GnFy0cc1Dcr1B7xJf0rsxGaZgYx7ATBmjh7HGpZn25NT534xEMoArFgp3Mz7zHM8Vjvyo2isE
6g/35ftleBRBq3KY9XWczHZ7VTN/VMLqqWHIjSXcyWtwV/bGeWCOppmEFNxQOLnafdLefV1Ly/Ei
1P0grjnEmNmRA/krunStyBNPrt0cjj68srn2+OA63wAsSC2N3hvh/rJIirY3S8oKfohbsOmVOO9U
7EjyZNNpFwRb7BFvIvK52BYkubc7D6Wvj0BvYU+qUhQeuA54T7Q3h+sFUz1/i9VTMITL/etrXPrT
rFLcSTrDiMm8Ivxbc4WJtcvlbEwJM0goDzETvTd6NwIm9vjLPtGhMtMOxod/2MMJ+fUwP/tzYh16
6fNt/c357xCs6JHmGqd1o+/11EMnfYfa+9eFIsmEa6IBicrnRVaQHB5IaU+fYOTkmnIaiakg2v38
fRvHesRabNncilL9OqCg42tEAJOBjwCTfRaCQ8+Z9TD6HutSKokc631ZXEV4Vegll4GUwozo1sCs
G6Bpq/9EYSYC5t2B0O4CC5vZxwUAXfO2UgBnn3hYY86fOvUvHthHYLd61vxn0PV6Sid/ssS7Gr2N
VdvDQcD0uppzvzCr6PPlHKTU1JEpD6iL62u8hezHvGq1YAdMWIWIdcdhyQbgXzEGFxTxbGcipE7C
dNCZ0r9NyIgQxPgHPBKBY4o21Bo4FHRG2bC2f9d3LEqYbAQWrG0da1BnvJnRfsEiHYAX+nyQIBoX
gwAzPxgTIdyFnRRQ7FFNdQMBt8/74E5DvyhHVaNnVzjHaL1pkTZF+t+NDsEPH0dt7T8Zwa8du81L
nhi+P5QbMoTeIppgfR4GBr6zbJX1tc7w4ISxdTHXvBdLcg/O8IypFyacdF+EcXZyJkuXO00OpOpH
CSStNO5oG4p2Y/W8GhJ9GhaTVyqbnj2ZoWZXH0P7tn4CUS0Ea2Qi2rkqaaut5/0EGKGqt7czg34a
PpUcVILc8LgdMr8VoSLRo2Joa1j3Qkm/IcchaGrmghdawSEIgny8oe+EzSqbJT4m8liRJqkt1oDj
vf6JKlJGN1Uz0QUIDET6n7x7xj4vQZEFNAcS0Z9GSa0U5yqdVDssOMEBI0Om0+1uTzmcJ3MYbIaq
MdVws1TB1L2oYn5rKo3UaQNN7lshk1m7KawSLh8lj8nQIUuWkm5gQLY+J97uWfz1xIRiff4eTzcq
r/VG/md5fJUQycSOJOmr55xreQ2WlcQyeJXkv5VQ9Kxf3gW/TojMdqREiOWMzUHlT8ND8cS8VbiQ
/MtlLsNavdbE9fTR3jzhZ4IGanvlUUfmB75F23Im7VfNu+hTYfrtGq+uGUQ4QWSYYKNctuIFksZV
mmMHW8K44qWLEx31TnPn30Sb9RxfkfqiT7e9Dv64rERIry2YVAousod6gwikJVXWr1LwoYonA3Cd
z653gVOZtaMeQOHWg7iHo2pTprdublkaffBj9WQWmM+PNZwsTzn7wCas7QVrIoFL2q1egAD1mX78
vr7zZtldrm+XKQn9NzjJyzQaEXaulvthds0Xm1Bs68ZoSpC5el/dinrpkQcSuFx5QRnz59MVzNtU
Fwm3lxTc+hAwP3zYaC8ORGcpftOIIJvWfgUgkqN2avrD8YoEDiqgBP/cS4tsQmm0i0dNy6yXqu/K
Bz4q385OIp3ESqbB6M608zJ7cbyEyWALZCvd2Ns2njHYH577ykIkpOB+MCplDXOe3HgrEMRcFGBy
5wIDT3k2ktKKsfvmlizy2kPC0gOuJQW95PxIgggBDyQF40jtOI3bUrJ0p14EyR7f06nzziNOhQkQ
fnD8foCM9pHW1RobDpbyqqhhjURICxJYoQzN4advSr82xh8F8xLd9jacxIlNPm+3rhCYUSanEJrb
G6UpAHtpUipXcHz7C0vYojSzWK6kKeKjf6w3q7MSSo+GZhOssWLn5fJk9n5dKjW/vDAxm7VTftSo
BzCYbT8+x60wtVkSzBoZy8ZT4fKfzft0gjqRixTRN9tNuwWprQfQ6i2pOGn2aDbzSe6ICwHeMt4e
5W05MLPXyIhBS6y28mLsTyl4kjYag8eF4arDIwLpaV9tLm7lP+qIr3keD6hC8Z5fBfgqfebOxEhv
bn4ThKVYk2bGg2quUAyQn1LMe7JZCSTf7cSGjX3lzv6doKhnso2wqOzpyVp3vv8hSgPa5Snb4dGw
b/Pk/mZ9QYKyBjtrbnS/RFF6IahceaMYC7S2Q0CPSajBhNDrhP3lCODdfKFLcyBSHCKcl0ZrjUoA
X9w+O/DlkkFrV/LJq3eEhEis7CXFVEkBBqT+JiLGFPRq1rUzSSlMJy0Of72+Xj/C6oYpXdTcufrC
4RJBiTnk6JNlnw49jAWWmUjGgo4v+BL518GMBMN0aTT2uZRnKtgbFL3xQmUQPRI4+dWWxBvO6VLA
6/XEyoidh9s6Cz5le5hwtFQdoZ3TTWO5LpDtHiTxTa8r8HBbzJVSy6QWIa5d+FutFjVawubanFLz
xMry2vGewtCx1ry7wbLaey5jXnBp+XJorgZ5ghtlDdgDIA/2WcsPpAcMDlIjBcnG9qpixDRiJ5L7
93p5Y/thcb+qL1FY39NyQBKZPmgC9rnYRb/TUGrYnSxnwmleGtkCUSRGZ8pMB/xCR3QeFghvM8B7
s7aEcxno626vy+SX7Q7tFZk0hbyeOq/qx33ow6A3rQPp/DVNlzqBANxBx43hLMxJ72jBS8kpAmln
CZQnXTS5+GxX0KSLhd0ts+Y5ynyDwcSL7IOZz5dFDID0GixiLtomawGs2Lfwp7sGWSVoVEQjig2J
qFke3I3Bmj7ubr9qr6aUlpLRKBaELJdNxS0zZI8NUM5gyMfLLrAoCodqs3bbYqPcmW0DN1/q1eC8
OJ1JH422BncLBtRHda+wXSYHh39wNsiUoxrcxUounHciF6HFsgaQqY1tAVycP41ySua4mlisxNDP
gisRkADPibjaGsOyVBsZD+urz3G2grMYmF2Dt6aUw0wQGbUGjvCUk9Fja10OW/yHzQ0jt28PVsF+
bqWp57g8KuT6KPimOfUuQ2WpgX7ls1rgs5XRDyrsZSXsQV+a3msbi40sOBG62pVvTr/OPTmMk4+O
ra0B2NFfsDRiFgdN2huqgycVundFr05hlX36CgQn5BfO1Ev3pDPKlxaSQ9fKWse+BEbkcdxRnf3s
4QlRdLhpvSepuPCm627tgAmtS8jhOaye1OYvBn1o1ddSzfpnA8RkEko0Z0B3gKriFuhqc2ifOkd2
2kRPcDYRgXc/GD4Em+z3TerxUTxq/ikRkC7tGAF1s60ChzVyxNv2pqv1sUtLJwfvLywLAc4M5jDR
f7fNo5Qg3wSx10dOlZIuL1dcSdYCZOXCi4K5LcmCzzsNHE90f7/rWOfhmPLv0dLIFhSWwCPe72qT
fmcXN5e83pOV4ykOG08oUsftY3qLMsfPSNR4d7cH5mMeaIrH5I+K83MHZtWVjV+DQK76PD9Ai+f5
51hFyEDq72Uyj1yb0iqCTWDuXLsIo5+LFUpSppLySGHF9XDCGNXgMg7HZc/S44+88VG6t6A9L9if
+SfGHIQyj1NtQxb9OKAjEhFxXQVAHh/scx5XZmHJkTe0R4Bw0DBV0PJFWZDh43BGA6mGXA2I7WZq
bDICaGwOotBx7cCnz3lpRiOZ55b0R8QsmyJdpgz4ZzND7p1KoF1SxwYhugXQ9MNA+OKHcelnRlxQ
hR9w0HXYMYSapMuFaYx1hDu3elkNW0Ysmo+2z6UgJniM9939SP78sUw/9yIEK3XfNHqTeGZ9uLto
Ds2BMChbf4Gm5khvPCAkBFg3TMorpmXS8m+ipydauXEr7mNuF2VYhAREcmyZf/mjwwp/svhAFC6R
6xhMekPfQZz2k7KNl4yKJb+lK8tCubRgfTLIMpEVqB62DBgIeosoksk0bKm4zgNLdFETVX10Rru7
xwd9G46iFNcQrORnjztsDJrMpk3DeNssLkeTJNKuFyYF/x+E0bgIakImxYMwsBL47FTfakVL0kDS
jrk0si5qbVbk7MANVhE6xltlLGkvD4drVJqwbILLsQKSWcTTn/p1iMvRCvX9sZ6r6Bp5ia7g/Ngb
PBFMT2pEsMDnX3/anW1HGPi+hVmGP/7H4U7U7wmjjSA8q7QP9n7hv7KsnpVN/Z74YRk3681nJIn2
1dL3tFm0kO4BPQQhoUOvkbJKKL9VFktgkJLzhHRKtR5DETfn2cfiBJGN8+fyVFRKCdzczQm+QePa
FulgvaTu1j4+fJ1Mnz38d4iIhLqh1dpzK+0019SoINk+M37wDbADh8cw26v9jeotds4lnNZcCAl/
596UBem//wWJQqybzKNvlo5wEEpWHAzZW/VGDUgScLKc/GZYWJdMVc3G0vVLe485tPDVQOJaG/cz
RwgnDd8yV92CLHFLZE5LjH21m43O1+hhBrO860tKDOfXxKtqyO99d0aYEl/smEW/qWfPKRWau+sf
dYDKIkgjPlBFnIoe333Xbq+hga8gvxdeIeOwQjXNPX6wuPMlSZ55DQLy8jev3VldI3gTqteyS3Uz
L5rmutOXUAwtgt5vStoImFD0sZgl2CnrFr64vI0RouDZa/Jkh68SlCOOLJzDa2bnQ/bPd/LNE2IR
hReCP1RStUTqYSnkkYDjOmVddHn9eGZLh/H9nYx46IWhlPXv6F3Htz4poQCA7k5WhJ6TQMEVaKRY
72YI15tRpLZ77C3+7kRY3fsEckNgHEKF66J175XJewjyZZ6Xizy+nGoEoL0jIawmDAnPinfWNUoL
kCISyjMTEPNTwmAVtfWPgHXVV4GqrC8P/l9UR3f6T4KnIrclX/wjvoipcLu64jzjY8ZqDM7MuxdL
U8xDA+B1FflI/OVPTAYFwk805DZYXwyw4mp/mAfWk8CU+Gz8msMVfYztU4UlK7cxta+ZBn7sSUbp
2GOB9ZgyInjx670rSMatI/bLRi6x2PTg2FR6C4uTX8a8f3Xztv5LoL3pjYrh2IGy/FqTtviMbe1H
IHEErACnuBTPRQShOfzEuueGOVxrDSIo8kMDw71VTWu5iKtPDzojJNqj5gak05yQjXwBVDJe2++G
6yDoXkW1uDtehGyIvL8xpYSRXAKy2mRSk+2raF9rTLya7vLiT3ZXGtXiNn620bxCV3iaSrOZ+Xkn
yt2tZwnfEH2X8HokSfh1rTbmvJw8LPg1zNlIKx10NFmEZYrrwQ/aws2tS9K68jryMpU367UhtzMZ
DcaADXdTbuZXPR27EqPQPlg0mS3D0iyD3QCNopaVoBtFb1Vsxw5yoIhK4nxyS4lAJTkVyh/lbe4/
KGKa0nxX4BcJ7DWZfCCRwpqbWmstFosV3jmtdKRWtR1bI7Ub43WMDD2btqttDSyxPdpvv5AVyngV
EaGyJoAu2N0dhnx7E6BcBp+dLUEFZvDNDYJlEnCRwDlQFHxeBM0YOKCtc81NtkoL4XtZstYbOVn+
oklqXuVOTaKCsnzOgxGjOK0gfjVfh/tVAzWAsMo7+l9kQVHyj/R37MN76SUeXq2c80cJpKMCSTQO
RTmghxSV5oc/fT2GCo+us8Jp5l4l2uGRHM0Jgux3aWkJ/8ASgbp/A+MakAgCCRAHZ6UcBN604+Iw
DWIoztXGuZVqMgj2C3pTTSDygJji5E1zAlB3NSyY4joXjaEWJhmgIvCsENPhJ7a/4yQ1geOBvZV1
7EOxQFWshCk52RmgF2dVmvvAowDrTVmVBVAkpEeHe+z7J5Tjtk7Hk8k8UTZuCmB5dp4q8le8RBOc
Kom9Dlyz1vCsT1YECZFNR087NYtKxVVeqNuCM93giINOySHgDUP/W7GS3v/R3gK6Ha7NnzFmmgr+
C1D+AZ9lSfbmPqsun/s9hpfW7+LIGuL8dZJxpa1o7ADq53OJVSGm908hVGjZcj1Yruk5rZfY6mCa
eM/h5wQbAVLPsXPxi7MkgjAkjkEZTHtPnnJSdXGz1oabRLExzydWfeE2eJUF/1/EljAl6Xm6P+Py
ew+Udy3qeu9lQM4FUZvWZjVJgyJBuj6mByfbIYqGHNgzWS3MpfcSUtaaD1OUlVdvrz0TrIRlZ4vw
XVkorrH6SPTZJ9W1vxdaKRM0GRy1DQZA4qDILPRzMMABXz1XHpUDCGzqTRG8DRnE+taU4LXnLzGB
uAMsqjsB2fSJl60w8jwzskyByxK/wY4Emoho+cBi1XbiURk7EOnzZhj4FTAP4MAvoXsHGVhlHdfw
nFDy1o/8YaU1H1VXfsncLSqR4lXOw4rvblu2YkG7rleNLsHZ3SQdN4awiUTFeREHlGtRFOyJISjl
O0RXFQkhfFhMMKQssKeLs0BQg4sJyW+lUkkCJXXysGVBD/gMNE8UTKy4WKCQmHQmfrEq2iMmfwQP
aE1UEbr5hE3HzWMlhOTvwvk+g/rtmByqkpBAmH0pPH6yvS+Vs2M6JLXJ7YZW8axUIn7YvrmCVWbz
59GuPBE5K1s+f0+ri0y7DjQUWFJ1S1W9qLI4BPKdNMzGvqukyNViWRtnBruwU4vDGHXo7PPQgdvO
oPpIkbqkAgtdtgNIkDnGfapA9VbLDOnD9WFJ4/8YGyDaS8nVzjJkJe3KSihDm1a9Rbf7e8d00g7/
HiRz651waUmCYOjSz9ctdIT4ZUnAueiK/fisfHsgL8xBzIGus6PLyxDmFy94QewKywfWTnU1nucx
cL+9ss4lDuBjClRw20gp69tMKZhaJcp54l1+WMt1hZxewN6kSwK4NGzTw6xJvNp+XpbynajVE0lT
r0Pin68PNKiy0t+ep9fUzOaGQoOlR3bXmg4ae1LiTAHveSxU/khFUzCc95pl5xb+7ziy2yf+zjNt
vOIlnREBTvAWz9SKt6fboVDkh8hZcl9nd+4c0I2eFfJvl1tCsXzYXhk4kxW1ySLHNsdZ+UHjn9Le
70VrZiJyixeWCVfsWMq+JeIz9IxDc4Nj6fWwHDdxwN+PnYsPpwzUkYrksAErqWYY8LI5e6CSdTAS
io7iuJmqG7IYFmzx4zRRaUjsER8dcMfg09baJga5UCcO8I6HJHvcsLNxcle8+cH6n5Mtt8wUxKYO
sO4ieal0CESM4pvl8CO4lDFNzy2rKIi6qZAvaH2CRAx4qVtiqir7sX0ppIr3kqEFVAsbT6IAf7z3
Kp+/Cj0ZNh5fD5El2jKUoFCqGxd/CSqm+0n3LO0JEYvmluD7WHw1naOYejuVCo5ylNMxqMMGZsU4
l8XNcB7B8SSwlohUkM/2i2f/Opsjyov9kSN9ZUwSeBCMqbgK6ZrjJvQvL3Jj9U5IqV0FyB2bWWYQ
5JBSSncesypfH2vMc7qrGXoJMzFspRMXx1wZOW+vwxdncDCC8jDBL9FhCCcwEysIfbpQcms5ZBuZ
celD541x3UkkjEBOPaCszLLblqphEmjG59apCBqDdHZZyx0kQtfzizNXX9I7i7smUS6UXzXagpDC
YW7QykAZPiYvEJLjUVtip8UU7FL/kcwO+dCS3WkK7ZHSNlw001LvYp3vzuiYYlePxuAnjPHc6Sp4
nupXrr5p2//7Oq/6H+qVL+z+poz3Odhnf4kx6N8ueaQ1H3YOc6O6tb5yhTnXPvxw4UFV4PQq58Zu
2TC18SahuGGijPwHkXUrveVr71CHGzRfa4DyqHLh6a2v3rh6ZF8DNRv9im2L22Gf39TCgtq+JLJA
IGURrC4JMbor1BS8Y49cGqG2byLKoP4BS64E2plOPhD+weij++OTyLE9Gk5ycUbpXo8iPYCEa+nJ
G9mdAKDDw6aV2EOPcsWqKVXlb5qGa7u7F0VD/9jFguj2q6o0u03HYbhttdLL64sQuIwIiAysdAl8
1GZIfdOa6L46AtipUTVy2HKHMnJY07c1CYk50zqzmW2/yKIVgbhzvD+4990SJczB3fXVE+gvIUqT
gTcJogMtVXQkdcY7PhzJuYHiSDR4rSWncVcD3hZStLOY9mVN8wcvEKD8+tegpVuehgXNQ5V+T+Ze
52mz9XXbBifwy574dagPaLyhq+WIswdplC8UbJ2G5I6Lfw9LTrKbgBP+fIcOR/4NmC/7zRHps9Tr
tWiCjFPhVRPHrYOiGqJVbExR+713+uGyM1bI63USQHANR/c2+6aiezXS773oJQooKYNCuEpjzIzn
/x8sOgTdxeZGnKds8yc2+SizAK8nXMk49aVlyvuVVNEp44rbnidmNjeW/ICOPpPQuzj01CXbyfsZ
WT6hdfY1fGuNGX4+Y6nVrqMBCt9MqSzyHtjkok4iZAWH0vKtdqs5HettYiW2IcnRnochbmRxqPKt
NugkLCk0uGZNq7LHY3dqHoMd235kAoKHPJvMk5S8mmKqy/1v+F6HT4Yv2VUVP3rLxQs8NpjNA9of
ckeykWNwp3P+AMX8mxnz7tLv0hjld7iC5ySVmPCzul6+8L1rN5T5O7Xh33bee48yGzoCsbplAzvp
MK39QaEVEg6fr/JmhBzLuwsT/lHt8kwzjmmU2QHREOWpo4oEjE1k7/Adx5H6jcUWoeH7nJrG3eE2
mUlODoXWMRInlWtChzTCKxtuzCwEleZr2rTkkkshQDDt1MIs63cWtcucS5X5Ph3Rb3PXJk4T+wfX
8623VzbWYrz4vTXEONTifxAZzFCrfM6EI7wnANY4mXTdAR4CQK+moH+30j8wtNw1qJ7tZIyyRzQp
TTfRWRXHEMC1Q/Immkhm3VohnAUYAt9yeaR32tNtp4KUu+W2wGNukzPFETGLELXf8pjYEUc85zXU
3AU4Y5GOI+V/0/UOBqOMxrTT4NjAJ39DURt6NiWNqTUO5naE3M8jErJmweGiqChOSeMjAOjdzOpj
ExNmu3gMU39iWPiZGDml90+EQ6mq1EogdNhexd/PTZQRY6ZBuk5fbYnaoJP9U50ErcBI6nx4JB3e
Jjfg98+qyYkJN4UB7AmuAFale4mWSV9ckAe5E6exXeNlbzj7ifj/cVUKHaGCeiGFcUsOcD2XD/oz
FHALuMZVgCkg4Dkt+P9fjBTxFnUM/7CNJQNUNcjkWBq2wL20Jj2MLUB9LN7oeGkz0qK7Ic+3W7Nr
JvBz7o1tg9L4QF9KKp71Gxu5f+WRsnuUMkIC71BfXr/FkzT7Ur32RDaFukJS2bwsi8htyhB1fzQ8
kPAWGfpnGzoabA6ufh/B++4l6A2OHsMWGPLU4QV6YeJKVpoE3nGeQ0kOk5s2RRvY9/rX/EPHAHZq
ZofJ5bbY5wYUvUAWsHgh2cP1DI8mQG+RCK0YhsJjRQ3g4f04yHZ0oF0oZKI3RMYkdEeRlgl4vDiT
HIt/zFkFdVRhrcyMrz43q5/q/INUxZtosCfOrtHv+/PfIrlkGvmRYkNBPMknt0BvnJX4VD0EqRcV
/6fohiScdg+dHRapokPoCTBvPbLFlCxOfR3kGulzIwWk3lyLALf0B8lM7Na5hFmafSnd9mQpDyKN
yTuNjYLH8rwK9pXYG0y+JJHpAcP/3M2WOMoJhmmC2BaAxZgtv2/D/xge/nCINrBuuWk+XbSUhOeD
0G6ac8+iXrpVmhA13gwumev8R7Z6DMjYAxWYrc3W5jSxh2WfDwc+936HUcfZAUlmcj9zj6MbGFbP
9PILsK4aAJa4NJoe2L/w1Agqd8dxcntVDuKS5sMkoa8ynpHFnoUcEmmyiy3ossLAPKu5BAAWWzu1
gGu5bwwoMW2u2KtwOvMWJlaEairv7f2tVR33Nd0NT8jtcVn24qkLjUeYuiNxWQq+C5NsV5eT7fwj
j49Anzu60m+5pZnp2mj67NbfjGuWDeze95d2F/41CpqZPR8I3VSUJSTizW4eMQFgEHThh4Hur0kq
rAAXKjPzdNqZq/JVbyp/6jMtBzktB8f/koq7q5/PuuG2iAlo2h3vyYTqx1UrU2ym17dXrPrBW6xZ
pdix+tJJPjYH25FCu+D19ASsNTAZIBqk4WssrssZ3fnNQIkoE1qqPABdKIH0o9bAzaZ1i/m6E2qL
ELprIkKJAQ2cc1tDZ0lC2H5+ToYR2dHEIFazt1V632NLtCdy5hteem4j75js5QQAGPX2JrxAfVu1
fhmV6mX6djXrDmRKMHMJwLwF84Prnd6O9As4SSHjAuofFeiu5oPZyNo+m8mtwU2bs8WxfcuKEbWQ
vzIhvqOe9LD0KP7nnz/mxnRYJcHSLVSAyzMg4HJunGq3C3As2lhXiN/PtpUjstPi6ka6sjn/e3kM
jns00ZLJnWIHhDfu2+MpeQFlM5anCosTwsZZQ0QynBS98AWvedsUOQIn5+mhdnGKoQlr1DNLVB7d
XcXj7Q+rnx3E/rWO2dIRAFZKNGVDLBYVHDHa4NiCkd/jah/A1MRa44gk19ic7WabBio/yMpS/Y5A
DxuxpRFdo55WDUDa2dKG8EIeCi778Krnvi6PlTPAZfbQoODKKVIvfadcKRwCOnVHGz8r/bf+ftTR
Z+OulsqmyX19oH0GTUEfnk6Z0Ie4y9z5abSJUvlAPPcOmBGHbJojFY1tqF4cfvlPgvcOMZqGLiZ9
qwJBxbCm8qjPUkmQNTDFULzCxtvdyr5Vg43HMYV9gDmBfNBOmdKhHpDSwa3xlLyTDPJBAy00atFe
k7lehxU0AQZd1fLB6N0kVUppPG+dnL7Aoc9IhX1YWWn+QTxvgRBmJzyEUPyw4AvxKx/6H+mCW8+c
O+PnNQ1nERD3P+1oheu2EhzhtH+k39fAgU2wCqcocAUYOnqJYOHoFrDnO5YBKpGXmvuX2MIWWZGV
ZfuOM6P+7KCdP5RoPhG19OKnRa4MY27mkcD4mmPI94dCSYxbmQzrGfh802GPN9YIipIBe0Z76ruH
kMtxEXuiUgcAjB0CLFByps3t8JRMA8gE7U70H6I81xejo13+ir1yoIpJ4W+LLv51XLQ+Y48ofx9T
PPe/tBhnh8WI2aruBxTeOZqDUt6+YwoIpuz6IsOTP/ZsBdki9DlRJlxpc0ZP21rMEDVtWxZA72pI
89Sx/nXlX70ulNgpRRZuDlcdHOE7car4yCDanDeWoEPDvhSsPycaDZ1AnBQPvEj/Qg+7hOIb7k6+
sqEdVT/o3Ha5w4ifns0RarFgX9CWVvnoWmPIych3Ldk6cabTrV5dpj+1tyjhu5xoBP9v0UuZR66o
wUmp6qkXO1uynkSZRBFaspkFFfbxmmqU2W9Y7ZB01U2Ty8/R6lmu7XfcD/tj7zuHlOrPa5jgq+uo
pjm9ctQbL7nBMFnobh6h/YKcmArz2Tk0gPSwWM3Jr0iw2d58CBVYpBpeRsZ07dWmeLvypv5lCxM4
ETlpKSewEZQxutq6a1e0GkH2ATNXr8re5/37+FQq3U6xFB5SJG1+qyQGxGsO/gsXnj0TDsjxnBEO
J6n4ZN1KAK+M5rU10PghnL/Ht6/5v3ZKEUDGfYk2yIhIn3HaUcR06sxzWyM0VlfMju5WAM2i7LMH
5CpWR181CypyWCrz9TvtlNnPmqoPbq7H54WA2xnlqDDvTvsKsDF1QaP9EpqUdpaCP2+c8VOSWLfl
RTxlD89PfDmCFpRGHCV/ZYAREXXB0hSYNsq0lak4KvVWdX5UlaMUh2vyU+zkO9r3UFF0rz4WBuvp
WdgJCiZZ0gsXFuRKXAoiObrvu72DWI1dWXRE3pL22PYHlFxlAI43NZkA0gPhgcr3P9T0oIdFHTBX
iGxK+H7u+asvVNnLmyULi7rXWpSMadNvQ43A8WLfT5Rrs3MTKHBJSfhBTwBCkuEmwitZbxkMR7dl
VwQiPK7nPC6C8rfgNNUBpvB4NIScr0iFwj7IXDxsrr+LpSMWJXNLJHOFqm7HEhOTrKc2kkWxHGGp
eHH8MWVafuJb1S3H5PsrbBbL+xKzbiAwoyU/nsn2Xvyi957bEA/Gws8iEb9oIFrCC0UTI8VBrH0l
QTh8WLBpCT5pE22aLbMULIWSVpLyeLhTxYBWehQkKjMqpr21gWZrYPSnyprwW394NRnGbA//6I6u
ATzkSiINRfWQPdTV2QafEzb6ZbA1KY/kZJ0kIv/7MaGamWnVHVoAxz8TgvXMdFiVWdJlq4q/gXhc
H3FnKG0GEkJ643Hv5hPZ7Bsu8+rDZKrwtoO3WIm6fIm206iHoonmE+fMv8HsscjF507egsKRPBBc
v2LxDCoem4oMX2cICMZYrGn+mDLXhCr+ugDiIX27viqze6/ryiZCexCcpOJBN4gic36xh4+ewjqg
jWS7FPAJalK3wKZYLMj+6GAfc7/eZ+0uKwy/SVJP1HTtyK4/Obyl148JC7jtiZyGbdubU/ToyL1f
vq1i/FW14vQK7tpnmGOL2Mixc/ItQ5ctXz1JTRqHoY/ofSy2TR06GDBPM+Y2ejrMxP2aKMOt7Eb1
3kKrnikYfDh50Q24f9n8mNSWJ8On5HcBEYgCSgRjf8XZpEM/9suo7BVfOP+z10ceztE5An52o1sz
3/285ANcJ4FZRpFhR/b4wUYya2DzcJ2TcRMqWjH7aPtsDoPrEqlifib10m6P+yzbbnQi3Lt54sGo
lfeXPIHUvmTtlUz8nyrH60MA24adi6nDv4Qb039X8np+efX5bIz6LJfRR72pdnG3Z9QtiFFh7nGl
aGa/b2HznkFTb3l1JVsEVZrGVcbKxu5+mdDWodE2PBU+LoYAgLJBjUASyDfSKLhrTZ/6oAEbXqog
wdPWoqsQEgAAafY49Hg+St/d/wPqnk5yRsYxgyUXZeHN10bXDktcU4gC6pr0S/yNnYL5S4YXGnpe
hdBsB7EuxgJgOxlpinr6wvkog6eJk2OS9uwHu4cp3WblDq8sIi9kFROusrppMBTEe6tDHaGWMLDM
NlWr5m/RYWnNaWBl04oobbjh+gI3KL06iDk81KIxhwS4f5vZJc70J/3qajZ7Hm3CORGjL9ICMGfr
TUGxxNBLZ4XihXbsd7UjJd1LJjXtgLtqHy4qeTTlDBTtlL/4dgqskLJKJKY/31CXwKg1Hsp3DqYs
ZwMv6YZrXWaEjn+FArSUNI/BspPTC7G22xxFa7eK/dcw+ZcISAJmTKs663XDR1D0OFXZV9qvpIzi
kJit6ERGdUthBR+Zjdqzv4OJxZ6GR+lrAqCGX4uA7ex5fIIEXwGOYx06sWTkMiGdJ/lt2gP/iCZ7
GAsV9IsBvXOWWoxbdzgpXX2b9zSrQNWF1YWnk3DdD5ezj5Z2Kj1usWQPKx+0BzVktkm6hCsTt+J0
MPOVNBogX7IBC/ztcyzrKM+tQvNhwbs7tB7HINhexp2Os4G1TinurI8iGp/bWUNoqf/Bp5Rp1AOo
3UpRVglEU21QWwWUsMy6QlboO8mgFhm8ZIsExX8noqQTeqRHlvnm/UANvQDA99fuxfJapV05IY8d
CaLlPAuG42F7RkSdHgmKQys79lTDwKDk9kbQtHtwm12y8xeExi0y3eV6OrlI7RVA6i0mjRx2rrXQ
Bp6FqDjnfwsPdiws8dI9cEnctGDvOj+Ck+BpFAquXxPSY1qybBLvD3JraUkuoAdGB1QytBZKTszj
gkkRUjHHtjqhPfYZfun1h8Wnuq+chhsfnEYUmg8VjgtWRDHwQEY6brnBJgr+Gyjbc/VJ/zsxgtCx
srysBLYjXR/9FkEWag2X41zU2oCJi64q7NQIJZel+f5fo95MvZzS3P/lVsXAy7C2AFoDTTxETJxl
/Cr1OhVPaO+oEehO8MHYG5iXAEaFKNRTE51KBDVpaf9VFI8Hu8nB6HWUjTABxqqxEhFTo55GEKpm
8L2o5CSVwVVdCS3tvNbCowbm4tOWbiqL9gkONBEJTBsOwqGtYoc+Qkt/86OtYM6bR/0uEcIBABdw
Du4OieaHvG7YCcQ3TFRSNW+E0/TZBjYxMv7jdIbuhG9MleJJdSzRzeyGn8OAaI7tXoA5FODf6fEE
KhJWLmSonAxPwQNGqjgQ6ODxWDGFL3AAtuuTWFd223xaRalli7L6p1KKATxEP7rZ4wp6CZ96Y+NT
S6J0GnjT7NNUDbp8jqFnGTj5hbl1I7Ba3ytQcrJfdFlNwHrTHoOQnw9HwBwIrqfHd9J7KfgQmHEx
Mt01IL2Go1s1s6nxtVmvoyzZWW4kd+F4n2b6GOqf3p3LEsET32PCFxQVPv0Z8X2mMrWwU3mNLJSH
Cv4R/RtusGe+QElmtihL62GOMyMZLvcxFWuY2y5F+y2o4WAuuj1Fq89zFShsDUeDnqqatF0CKVtj
3TcawAdbQvaOI2YzY4EDG5OaLzrLLxxBiJPHCaUpNX8k7YQtmBm1VwlVF8R/3VaMeuA2oA/+oF22
pLIxtMDD7C9AJedS4MMJYp2gok0pBebaVbKA1xKfyyfnzkCY1vnxg8aVV6J1e0vGQq+5bR8ngc4Q
BbEHsuAGhdud28/3oPLgKFymaOymVbDqZUbQYlqZ20d99O9mfpSV3ftchn1kb+ADZgPEq1VerNdi
PHpNnHmwYTpQGCTz4bTiN+20jwj2fCuRvbubeCl30av7bITg6KbNd16CEEQnsjx7nMs9N/hrt8VF
+ZyiEh7Ie51gupCUd6fhLTZzBDehqHl6Q2i6hexJ1GcKmvNnsCAbW8KuB3EBe/bVHnLGACRKSmC3
X90BF3IXM1RYtju22B14AlYv6ApE7ENpZf347bS3HavAkvd2F0tpW+wIXkaIBWvb/TnyUkR+Uzbs
w3Lj285iVMX4jU89SFWIrP2EYT7YO6ODUc/7yXqfejrU5tdP7d4F3gmO0vKqJ57Rzq0CJPQHiYX+
Jdg4cCgVACt84KQIroWdiNxsXuaaKMwC5it3tQQRtxklPe85+D5kSWsM1JYD1C1LXeHwMtFKLQjX
QA1xoChMzT0sRqN62EvWI1Wi7sKQJZOUpcUYHFRnB0XTBMPxZkUjgJ7Dq4nVzxn4wvnYWwTyJXZQ
/orDWQFlK9czNWzZJkkSYO8g+j4nOjsAR7GIjlx0R5wbbE95jsiP794KYGTlHjkwRqPpLq85KcZz
S7gDHTfwLQWX9mw71C053pS76LZ55yyvwhL2quK0EowWWRuhTcEpltVi5DxChBhteCq71TmXXo1d
ITMN0m6H7O9LNo+U6XFtUvO733q378yGALKV5ZPCLwsyFqgc8qs6LYVk6PKkihfHixHZolvs4/b1
9bzeNTrgfOCiCm0orE9Oxp329ggbA9SouiNhxIJS0n+jn8YoR0GF+4jZLtvNvsBGXhyV7ZXfbMmL
MfG6t1lq858uFO0Imz+hX8LpAV+HXf+gYIUPv6Knt4LjZgXxJNm/ayZIm66opx3tNpA4xVEoprbx
m7KlYGsHLt40QFDXIIABOhgDWdXCgUUIxxr+6BP80V3Wsyb7umdkoAv9+Gcr+zny1V5H2k4MZOIe
Tv4VTy0qQXBb9D8F7maJePFNjjZndEVNCtm5LbcX40mEkzcRSR528EKUoeWA8nTso+cT/mLgA6mn
4e2I/NfDj6U9Tizpf3o10jJVa2LWEO9HttYto4kogJ6DxvG4BTfox3Cl6VyUCtZCW9FgBlr/EUlz
RGUN6eWZRbh119V1e18U2QGwcpHs2nWCqkmq/OqKMUlOyuMRFXS7KNum4TUXVUoetCyaHNAuXex5
DFBxV5ENQHlK7yV65BrA4wTdUrpQdcW9/lj8AKcvxOaqsLeOaGIz/xYc0cIOjM6EMcmT5Pv7x+Eu
jcwHQBakxky19EpPfh4upSvhvXSaW1VeCNtUPiqoDv8w11nNwhbI9AzqeXXVi9f4AMIl/w2j9Pv4
Gj+L2sTQ646MXztMCCzqntIgS/sqXW9dx1eEqNEwjJchAsc7W+JCywLVSycho1f8bONz5I3IBirS
Yhvfh9TgjyJFliwfykNbSD7qQ3Kus8nyl1SyfUG0IV8kjWMv45Dj3sK7v1vwr8ASvqn06wqb5m9s
pC4zmGIvjHpsDUUkeD+KZl7f4wc7oxGQspMFT1Qbclw3G+jEMazelae7rW+T2eXW6CQ6em/+nGFd
S5apytz07bdVvN3rmnmagyLgVQqOn0AFoCGpAUH5199MH07QjwcPGMLiqxyEzMNyfVPaocMIpHwM
gl1PsTMRFBujjFNFetSr1rYYZX8hCLMLHeOMSNlfuH1s1WN6LcDcZkAGrqo0JQp6QAElM9x0lJPh
H8zSBKPbstKx94iuQp1I6R8vH6M57IRn0BRTjbuJoKfOuzQGQ2+9JWvqJuRMN9yMn2g/KcLHIcEM
fBPmFF/f3wM8Iy7ZvrcHB8yqOQg5H3Fq6XYR92TER7/iawTwBJL/8sarrzsvHfYTcdn/TQLsdjD6
ssHUW3Ze6ZMdC3Zcadi+Ql4GUkARpFT4oFjTQR7q5Bmtk458Oq7cM+dEJDBC00DMHjU/abgWdgSJ
yi62RV/O/k0dLN0MnxGo8IfvnLV2KAQmAgtkMxNFahrRsYFEhp4CdmuG3KeW66al0MY7lIWaFqWA
Mp0jYCbyWcCy9axOcUFIpPUTuhZIdvWNs0sCCZF3ftObT97avmTcjokcEPspAGzVJJ5jC6rR+rSb
XAlqv0eiie4aa9iQ2t3tVDuyVe5mZsdRNYoquhV+5q+Qx1xg6PoMhWFnOoLm3fv0XBpDZaxszxsi
CTuGLSAfZWNzd0ufDCM38OQ3K5qi+pc6ZvCQpqQkxK4CokNlfkW4TB6ig9VLL/Rtcf8stB4Y1Zg7
lcY/JSHJzJzXu2V+Gq4kt5n6rWvBNQPEVJ5YxMDhLl03l5KeNl3dhEshDY5qSEPk6hrgI9mZGJ8l
jc6Jfq6mojnCBrm050VSWy7Q9OdKhtJbEsBBsR3hdmmPz7pXLbwn6loWZ6OA3mWg968//WLGTghM
MlwfRkqqR5vMrG4fjlcASK4ffS985Ec2KKuCwlhVk5vYR2gFeS96YGM02iR0Rn49+PgsBIyISxy6
7ZuQN81ENbsvKb7iUKBTxixMn43o+E6pT5mZ8s3ubxnwFqhD7ddGren+QUQCLYexn+5Kcz8wyfy5
DB6PRes6CVcSrfFC+DQbfqn1DfRU8qsBpcLwbUL5DAfn7Lw8UxqR7cLVCAt23RiyCXKCBpxpnK+b
Z99+5xYaebRD/SDnBPTkJ7aLeBCjxSTD+m+pCGwCHAHPYaIUyAF4yhBbXLE640bmC3mG/rFhPVQo
NE1sFsg6/0gTLYwf9JJ+qJ8PESNYanY0Cytz5nK3L/FewslRE9pVw/zYuDo9uVzDuL7BOQzOQOrg
c1dTxRLBLBOyT7fuwQU/wQY4sgRP+FADyqQTL7gcQNiHNGQ/n03V52F4mFiCbrYw/3quVjpJP4xF
wSJeQZ5nQKeRZ8KCxClZjUfmIXSB9ASjkzkSbUBg+lHPD8cbJ6cdWfRi7LPeyU0FOouEL+sgZAiu
AyYAyqkcSKWB5wDJU5ddDcwshLTjVlwCdrXjzALJzahV3TEXpEOfZIP6Q/lJjjL88bDyb25cwyk4
5Y4Au8FBVKq8T7lPA8Os1wuLfxo9zGeKscX5qewUFZXiux+ByEnR1dKuNmEwWDZa3S6Z0VxOtZGf
isVn2uTsvJl8TnUW/JAtlI39OdlLawiw+OrtgnrfQ3PluxwN2Gk53A+WfvQI4MwJbJc9GwDWZizp
2xOLwOdK90lx0ngt3Qex7ZDfc3A7HPdsYQ3A0tH8hEr5gTEtZwohtmqoRojZEvoKbZiZ/aqFseD/
VaFwZGmru/vZ4y5Xgy2/s7+JVVSBKXyAywEpBNbIFifsFF9i1ENCvMUEmvsX3W5HzqU1vjuezoSm
HoUlxkqo+dGja7psYQxPR9v/0jiteGFguKYdL5wzwIa2yGinmyljjZevh+eDt5VCxh9k5YGb5BZO
E7WqOujNFwn9pWK7iv9MKcFWPhsFfaWzMNpIl5GZ0YbNsL8JuIuwZX0DUO4nBdPszRSKEBrwGyYa
7sgzx6JWrseQv1YJExFaWDHVV2oIwOGWSvHU/4MrwDRtVCop9SU5pZoQNR8pHweptXxdMMknAyAy
1DGBfNQWVuDVovGGlIszMHlCqcnwmsEMqPvzibrwopg0cQKEZKMruqUduMmdnsJEhFJg3Y3praA0
UodLtYOBz1HA+el/8KnSO07OxDvrQQ+67NI1fcJB8JGsIzwMd3evVzdSgjEfZbF2ozco+s3NdGXr
D6iEPaholoYkDgOelITW9V8taHaytpP4Dm55i0FUEOoI9nPSV8yejdiv33D0C5IpnaX4JsSVtJLV
f+E/xobWhbcUThbHTQCanlPb8fjDdVaIBhFBJyi4XfQy0L92aIFZ6lj9O+AeTJfEWaMYPok11BWx
XRmfOCZ9RZPAoolLwrGZkJionwgHVTK2KnrkGzt+4AwPwKTx1tzlKeXwcY+u4PvS199WK4Bf51r7
VVPM87cR8DYAzV+7sXrgvUBMpTSl1Yuxf/ebF8W7G/xDTdxQh+DvH2pRYd55CKU3KKyTDhGdJZhV
y5jSk4qKMcSqajAQqNxZMSdgSR/TnxfDC3ymeER5hPfOBDs8Eeb1bcM16k2IHt5ochGH+RRwTRoY
fM73+0IDGdwtiFdhJypkM+9wcNWZOBJMj7dddn06xklAgMRyVYLiW5TDWfDw91z4fgId/Lsx7imT
sb05Gc86CFo6r6KeZjIqLgWkKcV6HM5i2NH3q30crMYwiSkSyMIJgg6NxVJio0/4xTbzN8Npy3nm
7j6joIcAXEnZEB3THIaEoVjhW5kov0ovEVWUeLMRcfdjEvXDpmXJvSCFXW6TOgHdplr4/SEbhSdB
UVG4NQNLIFVXziIcv71YlD/BDXmHxA2lOa8RZpga7eo0TKh6fEcQSJDwhW2kCvJfU0TjwecjEhTr
KveXFEIhxBw+hxuacE791WcwAm/0m+PcuHnjdkjhZz/Gyl9HoTK7K43FgryIwcHpRSOe5gFj38dx
rvVEqvNlfAOQNh9QquV6eM2TqBPygARR1Id9c0zwxWAPv7VCzjABAa+huh50ggY9MOs3sjSeZX8L
HssRnBy5EKFZxCdSlUsDV4whxBkSJfcoZdMSrGqMLTBl6lvcr5RydloiH4qn4zsVfYO4iRXeXlMO
mhjXrGgqDPZF2Tuu829qngBJTShvCpkkvlwZ8mvDTZrFllN/2zfBxNIpF3GaitzV5gidIsfFNvmp
1ojNdjc0Fbxb9CzSW9a8UETwGK1gyFf7pG+SYbgWi2lgVpSArOwPal1BlYbr2TRuQ8Wkjtk42BhU
7yPE483czX0+j+1W4iliIrWXRlXX9SHFbof8xrmsyjU39OC9E33vJn7qQW/Y8XdsR1fxQxyjX7F7
DXm9TO+F2Rapa4UfCriHbrnSlJRFpw8X7/SJGZJ1vcBTWwVH6kqvFJ/O5WzZIrasW9VF5NMRKjaw
uwYWfCC8QM/9B3S/M9Ri6f9V6uK39+ncOwQNM1hQl5SuOp+xE+2CJ7xJVRuNQTifSqTgb6P/XTbS
mDpb9dFyqaYixTkZUm2gAR+eBvGAKdrPvuuXOr7GKTA5ndt8agrweXAtOanbH+1bMj7MmTENNoeu
AvPrt/KvUxMYHdEAxp+RBskyTGeeDaX+kimwOKd8ZtfantzQB319xdThPq6LhgKxM7eVQGz7PURg
EB2RKFFFss2epT/zlL/FKZmzfmaSJz8+FDgV2g+2Kxp2bPkLlvceiPr8skeICrpxVJ94l0ojG/2m
iUy+v6muAPanQQdAJr8PoXqD2L7dBuvO3K4qqRGMZV58zHozk/fJe6gGrg2loCbK67Q5Zd5nI6ja
cfsbRNxtgR7qbRPOlRWWGoIPROhz7KeET2djeCbjUsBYc9exwqYK8BZUnoDtKi2Tap44u/c/6cbE
b/S4VGVTWPxnGZjt9MNI4/Sm/w+WgpbTNc1vrClCHjNvGm8n/duqamMVVRpyUDNC0/l43k1YWPh9
mHsP9q6c1OEZCnhztrMeP6hEd5mqMiYoeRWJy/h3D70jMbV+5Tp1frs2/A6Wfr4o6lcyN5rqC5bm
C1x1EI3j8dQ+YnigMnZ9G6G2hTLYvUcv4B/Tmn6IqcN92rxuI14f9tM02hiu6iAzPV+3XCbglwHO
j/7GiNmU338TN4hAr2aj4/q7NW/mijFq06B4N8SJIfRTV2kIak5hKYVlrgVzhhdfL77lkXt/6fSd
UKCSwco5gUkkM2Btd9FRmr85MMa48UAImVlE2Dv+HNZhu2Y5fhkPoviiZeeYisJq7PvbDYQcCevU
z+crZIh61xfs2hzREdfavadgAv5Lf8pxZ1rUTdlrJRH3DcTh/xuUvLXbzCc7mrPqdEndJDGkETbE
O0Vfwe0jETNg3OVns7yJpN7DMU8QTM8eASvLqAXWYyiOjcXFI+QNcYvwTIMWZkmWdXavs2nsSiYU
Wsz76H6e+1y6quJTwq6gWE3EaS5QgpMa7l2Rv4TQ1TQCnZxTdAipuIxHlXcZZa7bMHM4YLN3KdRw
stZnvjkAd4I3VMeTuGwfQ3qY/xGKnfcXFOe7UODMqPAR4WAA2hkVt1OkTjWO8sVPNSirBk0S/lBN
a0QaojJrDxULhUqpR9/aO8owwst1i55QRC97B+CYbQfEUNz1/4ovBuZFYYaKCTGRm3FyaJnxy8B0
BoPZuoDC2qnUkTPNYUb+GmkAW2/2NqoRpG3snSpqXlGlVlVRO0lGN1aDYIolZux17jpMCNO7cVZL
WaWFc7EXABprCZRoek2Ugh0ZPvsXABo0orjhGhgWhBgKFBLCk3k6pL9aHA9Xm1YqACJNr+JO6GXU
ax7beZVCqBQ9WNkPNI15BkD+/aQyP8PNTGUq2WXeaFY1GXPkvnniwhhgncr275KmZa1Q+TvB4yc4
Mp6UpNI+0eAZ+V/yekpAY43vpgl+ESnDrMIXYLVLsyMyMbmu4en4X00SUzAz/gFZxsz7CFX29z7V
twVSFUUUkj/oWHNwHVwW5yIzuJxzf1Xg8//e/hfu6MHkVZ2P0QjiU3t5xPKYOB2DHe3AmoR12+XF
r6Kbo4gmy0SALusx9v6Zfb1//xk6PEETVyCNgY//6073/iHhMijw4HfJwErMCI9IuGD6Zft2VGiz
im3bK2X32XftXjEM3LgoCt8Cd9ECgfcHpEuI5tH4pCvR41xPgNcFFvm6+i2ECOiiRp/gIsgSM1Bu
JHdRbKS8xZC1Fixyoln8CIuq4AhUPwtE3MES16C/ZNKHiHrac/5PFnFelJ0Y1mPxhBpEkLP3/XhB
vouRjgGFk+jM8meEnSD4wYlx+FCIdtedJMiiuA0NdPPFrz98yxrU4HBsjRPAZJLKUv7hXt8tcOkb
c7jvMrXrydbebL2k56X7d3sPiKY6qqgIihCafx2KWpQS1NUbH/DdKdYbNhVVa7zFBqw1vcUFoDPX
wvjQJBSszB+iSWxwcnp8bC8xTEnx8+0IYcDVvTlgD61Sl9aaeonmYtq2I8oDRuJHQfhVc/4U1FOD
adRIrUS6Y/EZhZcwtWzcgo17WxHC+oLBR//gphX7DfFfV+lNVEVCDpGfgiA5AHcKQg6J6x8QzuiD
rEBb8ZKmcGJqjtCjE71kAI7+ZIKQtAraY56ia5uV9rDwqW6QOkkJnyKPfJkHaeWYjfrWcf0wFpk5
Z5H4FdhX/u9TtDI4hmaTRuESDi4eeV8BDXbaOFRnsc04gw4PCP9GxyaDE4rddPsvIFq0Du5qd5o7
j6UMvGgg80XULQeXk1aYz3k4HI+IJ/kP19ZKbM9Quz+PHmdw61l3kXpgQUw0qHLBwi9FDlXYLsMd
RW91pk97o0gScyok/L9fIbcKN/R0R0TNGSbtxzoqAyI7QHjAnit8616V/UFEu/zj/Fdz45DUVCoq
13VIR08KxjEmHfbJD9z0XhwdA+LbR44KxKFx4oZAeaEujW7uB3+DMqEoSxNs+iwKvqY2MnvQ6nHW
Gvryb0RkSd+NHBf7EGMjTrh5xgaOXqriV66z/+/ZJbuYUwyUKE33GuKLY1U81iJ7E6wH2pFSNeaV
UmGfB8baBwSB2cAH4ObCD63uCv8zdpGf8OdkQxglhb0e/cWAMfgv5508gh5UQoEB89h/1fPgaf1g
NgN25IHTkhirRTRy9+r142huVw0AmFPEHzYTP85tsCSyooDHTPdImly25TI2dmDBU8BGBmfRP7fz
onqM8WfEOZ3N9n3LJwfhO+Pw4ojH+2MHmEbkLgcYpaWv1gbu/NyU8Y/SjoGHs04RCE+sw+SYno64
vdUMqIJTUkv7yuxSzicUmgPrTLohYxD5wp8LcLxpHogpuFs0nU3gSHS+T9+TwDDo6xlOzolbbNdh
+JNyExBpqxOPphNi1gYypMqFp2LjyIkOrZMdONwDt0Ct31P+Fs76I/Nw2R/Z6zMY7hnZAEFzam11
jQOWizzHW5Rrybvbirka979bmvL7YcboPuHYBJ+cfrQYHS2CM0YxDbroWpuHF+1TjVoaKhNwyJmG
lrvwwNAQdJmq88MEqvJwp6M9tZ7lcaoCI2Z2AUHHQ9by0LT5wxJUAEr2uCHA7qONli6cPe9Fuivh
hWcYWXYyQhuB4NGIyLjX1+XrGuU3WUdwSYcMvetBjdLJyfAFl+MtFVnzCxomcdcoKfB7kTLXd/ay
XtHUo5xycEuin9hkbXuukKkIGfKTlgWlMjWyNFANuy+JkkR5ShJXVGd62r8zTLoEZ/uXQ0W0vICG
dXCOiVl0Q/+Orv3aEKSWiw79aS0NJFjdAOxff/wsbkuDOkCYqGX+N+IbjopU25uPhoEnNTMoAG+k
KzkyWQTLqiXefBFLZprn//AikEq8C7mcm9dIsouQpU5KPc2avNuf5lDHsF2zZl6AjLeq3s/JhPYW
NobhbOYN+Qu2wLhx+rD08BoJS6wMEt9KOzy65KaH8k8B204qQzaf3uyVmmCLNuupGNHwP2nfJm+b
w8zH7m4QtC6inC1XoeettAjV5ai00kfin7VQ8QXPx+T9EL+0LalG2MQ9aLAZ6qL1kuhZEpQKwItu
XruP7yuX7f9Sc3SHLk65+uzH7QuzElSDMk229bTg224sxeXZSFjB5gPMUXgEMaXs/sUCtrOZLeRa
Wo4kSMdrWfUBYMzyq5srGnL1eafYHXT2TPNMz4YYS6dJT6KnJZtGD8dP93Zchkjc1+HcxxTJHuWT
y7LlXd4zH9qY3eLQ8YJsW2PcSXF4fVQEyMLrL9V9vXROKJap0PAnDCAtYNgpEa68iRaIFvRxR4UZ
nSappXgKAv2kxB3RZZbRs1dDwJ2gc/YvlBX8hlCgjPI6AQfnIJUFMk4Itsvy+eczFYGqFCwvu7+g
ZkV7J+2+1OlHYsic5zphc5GarJLlDdWRJrxbxhg+H71ZGQxHFAwMvQHKqNRGWOLulQJEjHmyvZ63
9MbzGVvOy5G08gQTiHDOEJ7b9Tbbfl33/WNm/dN94F41F6gBp0geIpZ03xCurMRsM0TUgW5bFuXG
gdU3JL+QtjT/8TeOpRluMevMSJxtYFXx+gdq/UuGPefx6f7CW9ZF1pm8sZoMr8Jy9KfNSPsnf4O8
1jks9pXVxX33wrFIp5D7VUzsevY7o7smI9w/P9Cxh4OhcG/bxp2jNTdO5CWm5Q5jXFawKpR+asCE
TIpB63M6UA9hqqpupZcWbhuXVN/Ma2Mr/gJdp+vBRx7pqWxp0aMr0upyLqPutfqogssaZSgabjeX
AlCzb1dNTJA/gT0tK9sxUWu5OgclPL5LJxPVOLCeMEYzqUvJ/W/Mp9kLrRW1n7H02/i/R+gnfnc3
bxC3IuUgpJbVGyXkqMw7DYGQv5EHDBEc5HaTbOyteBcoQmNflDkRPTY+AH3qxUHLhMqSKiOzo88i
woO+hEXLeTmvvia7hiErSWQ0YeV+j9xX9pd64FbOdcFstnqAxPe+2g+HCEH0SraozfGNypeBCQxf
DbfLYafF1z9xWQtaAN0bBXc5fphxvQvo9NW+VmiAWgEAgnwqpzcTbgTIqItb+D7UJDNEA2c4bsT/
5mllRDsmTS6nv0dfm7ptshYqn4e3qN74hRKTvZkojkaaNaPaJ3gyqrF0+M8/iqEufBCtpRtYhKeJ
ywWHy6aqSGnfYNn9+XqQS4oPiG4aQhGCwq51MS9RCtWXA/nF9MocRQlPRmKlTJDhkG9x5V5kCeZi
c1B7h8OD2fMDU9dO4aVReJiWCNUe54FumoOcyshyiFOluybSmwAte95MzwbO47m3NUCK1rFOXdYM
cWJ/WEqUh8zb4IetlsIIsatqfp1hu6rHijvAvu7pBZUCbheEPN9L+SDx5ADOk9wrZvXWuvkbiUwb
z4OG818xf6pqGLi1jLC7WjURe3JUmNM+q8BExA2sUAkOfWsVNtm8uYq6aXwv5mh7cvW3tnKYviG3
chl6gWcnZcKKQe24P88zJkLbEcNjKn3YDn3i9uEaXxJtNQUdX/TcHbvlCfzZWyblhUsMd40nc1R1
5T5FCwnkKiyfg+tInO3n1NZ1ROibVVUn54LJ4puPzymhDKnp0sdof46A+j1Rm3Z2ySq5CkLb0EbX
Lb6RIbYfevs7ZO9kH1Fdh+qAt/1squpOE88Iihy6xP9IHSnVF9CXoQ6my/y5sLvhSysRmN+X13R/
BqjD1f/b09UJyoSK26X2EvBIStvkZnZg5UYXx9GXsQWyspcxgjyqC65q+cZ9zLlO8h+58b9GrypR
+ScVMfCVinExYqAo9SaHHMRhccPUjDSVtdD80KCt0KR5UAbzl0gIu6Gx2UXuFxJfJyC28+22RZzK
beK+hGOwGOMFiSSb4YY8SnLT7c45ZH9RQTP+07G6Ijs8mMSJOjmAItRBo4Tt1GCw+ErVudj0fEYK
mD0iXmCJW+XMkUAj+zfh1i8Ra2GNVRR5sVAorKXZBt8EgcKus9Fe9UI9H9wk3Kvih7qMYeHLvFjb
SqkMl/vctjfnB/szyKSUmhXT0BczMfYHII/YtdT0Y4iRx7H2WIJJM3Aklutx9MlChyNXdXGfy+Wu
joQuRL5Q5UeMzbDwu4HdGLYe3bsRNHAFzC94mfE7c34AzBI/c8WIp9a29D1LHiByp1Pht3CBHa1r
CrvIqgV9Fk2kjaF8yvg+DdboqmQaHVsDQdRjbuM2cq8urbhvU9NphZTKrSaisdQo6Q2w04iWDhhN
nfVPH4yY0VTSxweODqfXJcFatfENpwdyBlDhm04I5VaOHGyRagZjxs/8dx6akIILK5GlEFygHbrg
qqrpTgxE+0alnjeTKvrx2iASnx26ylAaOI2nax0xrmeA8mRR+KQQi/4y3Uc4JtopbffC5VLHIoOA
4PciD3PrKuT0NsIVNyOMgQpaODiIgTtJ8jgElp3xM7LNJJoqRYChEU1LoQTZ2Meecamw1KRlTg86
xzjDbUzVSEuZrNoR2+u26pMC7pHkwdH+rh0bl+TeDquohF2N4HsfVzrGDx/3U9JqLOf5bMKTOf/V
P6RjYa2oq5hHHjwjlU2ORQtYWx651WvZOVSeZbZnybOP8QcganLhQU1WdEw1pTjpD85WZPevyUGN
I8mbfE4n14ZkfRMvSLxQIx1ErP7i2jMKrErhriZXXyaLGXhxkYiyoRFsBxg9Aa7Cj8NoKCNFsIMh
EfaTIU/yctlknxgcPUHFqpVuVWmacf1y1Xui9gGS+tdysIr05h9pHMQGtQwoLS7Rbn8IQt7pUIVs
BjnrF+QIQ/9jyGCXVxHHE9WixVz10IxEf4/uZWxaBymWSRzfSpi2xWXLj8mDcfVJgzvQ00iy1lgA
wAYu7XKW7SMNkD0LK8oUOjJGEXljmvchvYwcg+dCjaTgTcEwLVpZm/7i2sO7FO3vPHjROmcNjT8m
mzKeP3IFFcSqAK5Z3vPUClvqp2gKQcGTLBAXs09++/vAuLrRv/vXwU2EWq2c9/dIRtflz13lfntL
gIJUn/MR+tfOkHwC5kV016nGlc0tM7YAnp8EYjFc5TVXTNFfpLzCglmG6uRaUl/ZY5+u79eiR11O
heZuLb7EW9QC66m5i6yPCtNRBINErq9c34VXXJTHLw+YKl8PAKgzLpNnJJSo+b+zCtetNScycPr8
j1uTTRKgm7agT3Z0URYqCSzuRzl0uZbqUtM1OsRyEdYho3bPgkZASfcBUENIztfyVOf1NloNExWZ
WTZRvPAX/DiA1a9I3diRQCaJvFXcEjdUpi60lwWS11S02Q+RC0B5MDElOaeERHg9Mr9sgGoIPD05
fmm+J6kBc9LR6EYZvOUwqOJrW6noZFoagXb97JbLXnzG+KoqZH5R/jfYgqO1Y1jD749Kvz5nwVF9
807Y2Ypbip9FJaTXfFkbG3WPO7Ksa/l+OFLtTfUYvRZwxhrZ72jahFXQm5fCfCISmXIUyB7i2kWq
5nbEdooC0A45zeV+8yDSfhRIifvYPwLIwVttzeoSkPoHgZ/xL/9zqHgrHnek+HGptiHordkPFAZb
+dnnF9tP2np2wnpipT7izRibnIQCr0q8xy/c4Xlnq49Lxm2u6WY+1BtmA0SsmJ2oaY9Uo5nNz8hC
cEOuTAuq0Rvtwx0f8CrgzVJfAYvcXlYOTlDEb+LC2rinzqvyNigjD4eug5Z8f8lAagqnPB06M9zM
vRNDYfH6m/P1bj8M8tQO8L5J0BH+ZEWttsH2gsEGBR4qUBd4LYjh4zdUxjftV4Gt4w0v9QjUIE28
Y0qDI404wHSkaRvqGttK+QpNOxhI8Qa55i4gJiwkdROik1G6VKGgikQv/hOn0CnxPwugAhBOi16g
GHZLRmJr7P2/5CQCnC44wX2PdAe7qCWs67Izz8rYmnNK1PS97XzcGeDiHiGXIT26JxHPkws2TON2
9CemwntXuTZkhvE/U2uCqZwLD+TLn2fsgiBHKBats954g3eIprN0XeP2ntY54M9TWkh59vmqMivs
TUqQSa0bTrih7kjkBHaHXMuBY8uTIHLCaEUPEvlhq8qsMQaBnIVeaT34yaSM2Cbww5bih29szUoZ
YcshYRWkjw0CXPSDygzRB5F9Kgw2I596joxJ3I+SGv6VAvVD/3k1hqxm4fEm9GForYkHt0q0dTH2
6hxV9Olz9jmJZWI7RtZ78I33PBmL8Zyd5P55dOBV6akyzxPVP72sNXI2ZXsThb/oG8PYYTahXHsp
M03LO759+DgCySJ7Q1rZUmKpMQpbdpuO8r+/aGYggOLyUSYevWjnWCMvS34zdYGxkqkzn62mYG1t
1Og3i91pJOZ/VSmIx/fqpZm+4tSGAI/Z+Qq9OpXq18G1weFn0pdu7w1xDZ7kvC1yJHpQSUk0sNyQ
1iwYkqHERdbNB5cnYiP/uJ6cox7gD9lhFj7MqlrbwxQmxRlPnhL5LJ5Dwq2FNigmC25DekdYNNVa
5CBbU1mfwjaGH5QyNVTjqQt3o4lrhwGCM/Q/OmyEN3KSSLvaGPMdgltDfseOWhrMNPLs/rYYgfqF
ZN772v4UyCDLs7L9B/8JUsrelUKbxVJn8D4kyO6wH6vX0/SI3/n+I6jcpSzbGaVHDQSMv9KnrPgm
KLvq876sXuB3FIDGfDAoZ+8WUpM7/WIs36KkQ2DFz5tGj+UBmgDTEaIA8IHlTeAIUyHiM4sX/nNy
/kiMPzvWfqDgkPx9HjF3UnBhibVUcXxoXREjTXgHRTk7a124O9Lybl1RzwILto5nX3W3rsTa45vM
2Jj+tCbbCnDpxUHngPbJIfGNM1D9W78TzGu/k73w0X8LAQJEvwb8DvH5okkF5zcAZ0f8+KkVczfq
YQjCZsYJMS7NWYNc54sETQ3oAWp5eB2svGskrnlm/mTAi4jehF3c5z9QuqrU1VGYBUggjWgg6Yky
UrkTUF66AakQItilQ7OjBAYVlvxP5FD0uPpr+UUqbJ9SBeE1iIYbHhVWJYJthseHHJ5n6kmVXhyd
gS30kIZ+ajhjoit/+kMVAhtPh4+SbmUhd98G0AybERdxMi21LyafKRwJim3sTvBZ2CP58XjIfe0N
5hbojUa+5boF0/i69x7Z+uDoV8SivEsh5LR6bylFMzGknC4dHjdp0kmdmcj3VpixcssLJB4Cpc9g
hlFW6n7976rtIsVNLkA9ePUOdvQSbyVkmscw1vPaqoXqO0t02Wj5p6QE8c42opQ7qeDHM4bxIZ4K
hUtJXOwwf/+NYOi/nR2dSBcUpciXBBkdsHbWn6NGuus/72Q62I+5U/m3YO6wxm5RoxlyOerNApYP
lnFANO0RO3evaOF9uIRkUv7tBHAMw6BKF/gu659XoJr+te5j8wkrrEGZEE6C31V+PBBMnonqgSjR
1zG8G64e7Nxkja6Ie9LJCNDRPDbqjJZugYnGNzqqVwQxiY1pbMDIZOFUr6l/Yv3/1IsLIUa1cJ46
9YufpRAYGPLXiSybIbA6TbQ+T1YhcvWr+acEZvdhlxpEF/lQ3YkH9H8pGosZs55uOBRoe7ZrwXjn
3KZImQLbEMCl5F3uDQ8zMU/zvAsrTacXc8HVtj7h4PmfpJ2SAH+sdfSLZe2j8OVs2LbX+NpzvjbK
S1Wm9YPFm1U0K/p8ASCU5t7Fi4UJusirbtSeoMAXr2DUIF4Evw1ROA/n4tOqRvT6rqWdnk/mX3jd
dfbOUCL7UYtYZ1BUH5VmHMq5BQNh5XlMjZgs1towb1IngXcTs1CkYqnkNiv9Cd2Vg7iCkFhktAhS
ETfNTqYZgYCTsI591J6zmwdTBWAJS8M+EzRSrXiaf5fSz+DZDfhAhs9vd1KqDFHbisLp1gjjwsG/
AeBYzFfNKwV3HCj6cA3c0SnRp/a7D4v1HTCCdG80hjY2p6ZN+V7s72+/wcHdrCKprgD5DUTmd5dO
JVBA+tANqKj5TZY6oN8PWqF0+PuKL1p3kCYXFDfla58j5RS+8N1oPQOj5xQZgtb7PNoGmEpQRgP+
uft5EVAMg/xWtl4KJwiIbt8JXP7U/lCNxLYOGJviNyga6DPfeGzsfV2Mu8fzfi25spLxc5K2hMTE
QHQpF19yR4QHcvDjLDRa7UVh5Mb0Ps8ynMaC05avvx8vXXCOZxohegh9uT0ZLuSzelLFfL2cpzXe
H+xHPb1gietLLChPgPSv4pdO2ydF9HaLTLqGzYoY+0/YEu/Q3qGVB8gJI26JC9zw8p2/wrYSV9Re
XxcdPJSuBuIr7Y5AkYazAarjURTlQdJoiBKZzdNsH8bSJ9pcZVbPT54aIqdgoCgqRxCwTPWAVAFy
xwv2jB1Ek1PzHBc6LPE2xtIbftF0SF7Xoc5IatmWGCQ2W+oDbdgldZ6zKtCDn3xQDMUcOXT7BXwj
gwgeGYbb7nAV+MVm5kpq9BUqw9lGd1H0ACEXIc4iz+jNkZYrDE3h/QuXzDV7krDVRDAoLB5RI7Bo
HymmnXBsKd49fY6mSlWvGZ32dIq3vYaWNoRLQbguh3NPdVREpG9Umx11t19pD4/UzAVtC/TAcwMZ
73KiAbLZXIkrH3jPqEGedavGGQI+vPFFIYEafK6fStzcsvVyQk/Q6ZTq31DLKnRkd5vawO1ksBQs
5Z7qq9jTFp6cPT/FNEifBS2rZJXdcnuAA8M1y5M5VUOQdOUokLFqiEzA0Sf8WTXlxnCBUfLbNOj4
FAK8qS8cNbCYtwPMDNpjCICE/FZPcaq2fckWT81U1SQ8upRJd+Eree4CLLJ0CNSGRsuXa3efiTDU
U11tdApyf70pvDc0EGcX+E57q4RPRVo7UuJwnEgIseNeDJQwERZWWYFJEWvO/53j+VB1OMlL/OyG
99piyVKjl/k2DSQEp+pe5Chq5Sa+gOr+55MQBlm2DUXzxTHpbtfsDPVuQ4n/SRbPf26p8Xhl9LSj
ywqK0QTPaQiyQjaAYJV0NA/aVqNwizKk3rinlVD5WSk5rz0s+qCc1JPgF5oTJYD00etzovD7YBZ5
MXoUumVGw8l3Dm222h4Rgcn6gTiX6xw4GphQ5SeplFXodj9dOHbFRM1xKHn+M0z3ieUJll15doXo
u0Icd3xEvXWDdoilWdyb1QYeRv1TZ89iwDyU42Xyh1zVi04fL2EQfrUCo4N596SAbhueWxVLc4Mw
XGIabpudZZzd7SP4zT57IAMwtXGaJ30u+euRHIkKoPC4fP+9Z7DFmKoT6B9rCR7Z2SVTPy41KOa0
eAJ9AdXJH2Df8h8dw29z6Ml7cB8Sb5THhooGOYmqK8R3mbpYKu7s+UwdksAv0GV6UDaJ/aYWWXBu
xweF+8g6nMHwcBAOmSDkKgapsj2qG8nrhlzHA9Al2YAdE6TJnQBdJYUjawsJnNdhaTYRiRjGiPiK
pqzqBLm/x1ZnVNPpj5s4DP/uCRuuEwqZL1JYFlZLNXv+qq2UNXgdxAVMIEHs5zE7UUs9V3I+Mlfv
nCIkBmZ0JtRrAbUckZi0c+YQ0/nC1tbBa7hE0qFJZVIjFGix3kOzqDwRL7PNObi75Fs9pdIpwro1
B5PA8Xlg7xKfS/870rIyMWgsyreWVKhPJuqwZjZy7REW6Pd9QdDOHaYufAvvShK3YznExoQincRY
1x5cJwIe4pH9Gs3zk+mS6kg65eJbmTvrtsK0N7jra50UBAhKIfbohKMrwZrvuaTdWPkEBmE1f2OE
YxKB6jPBagulJ9oK3dohMZxd/jFnU7bDLqiNQuJEEv7x8thfOWSX7pffPOeJyZZPNrGs4Bqvl0YR
nxK84ELMXuMY7a6yc7ZHsWIDfh5VLM1YnX85pToo8nfKrLZ2qqE7fopIWg9FXTakVNI/nHS7D2aU
V5GYwIAMMsoau7tlEnNZ8s248k/U7AXn4tj65GSxyNHg5qFD8ehdPb6eAPRSPSq1XOAdCOM91/er
qtfbTraFbI8sXdPJq60f0VpYmCbIqWhI+AGXwGZ6MYKiNjMlerD/ZYSsWE0ya8Vip6MNFaDPoDCu
XHaOIheib9nvP+DZXdc7voYMlvzK3GiavLmben/OUo2GTcn48ktqyc4xy4/NJHuKT8bmsjpihSJM
9zEIybWemAnKInweBj+LdbKok0IyWTA0vB+TuNRcrgBnSxAtQa/ExxZny1dq+mqS7fQfYR9pQtwC
JP772sG2FvNzimw25LG9oqkhbT8dm3lEpzKHD8bbuM92wAJ3+sSCclncXbRHEaIYjB7O4xsn7BE/
AdLiQHoNOK3rVMQ4uhGpTEThdnW1p8zVFlq6C9+i31wP7wdk8sQd4pgfLlE7phmlbh8z7kOA/w/e
HjiMgAJA0ZhQJIP2GiN2jjxH7rTO/hmv36Dv+nofsZw7WshiMPnBv4iHSrNqIBTHmiDAQnEQ7wid
JJXQwgPWl4g5xEhDnBwAF6Q5qwe9MjaKJ56aQ7UE0Uix5fldYm5xxR+DNDqEP2R6lO8AY9rUm+uc
ydw4n+ZzAzD55atYdINu8g45eBSh8yCvxWrDBz/bCCzITLaQb02s44MyVMdxfMPenxZDxWftO89R
37M9SRF3ZTbP7zumgjzE5NnmhSadtE7kAjetliiy7KBwBsVxz1QN3CRPLJRR/YNb8P1MwTafyQy7
dsd622vWu3wkluJN+FcYqpCOHJ5fIP8MoZSIcOKXyZ6i+/cRfirshKOae/6uvrs3UyusJtJyF0kk
LETcsd4jDTsYArQvlvyMeBrY9DGcbnceLA7f/3swk974cSpswRCQmndfxKkiNdGMlb58c9BSM5OH
kExa1G14Sira9ToIYAk2uGZeNk6xGZwmHwA64vDtIrm5wbwUroJaXK9nFD1DFn+U69/v38TsVock
WJ+fm3l5ZqLigFNgIimRO3/gUW5HtXaxqk3IE7qOXzPUkFcQ1Rdt6YfCXsMKiOpf2iHTvkRjRjt3
kRic6uSbbfBV2WcdWRWBz5Y3fXCoLJCVUuIk1ycrf12vdkWq5ZaYohqq3de2Z2sp6h0KZzNnAKMD
13AmsJZXT9lNd55kSXGsPAXxo6GMLOznCUEGU+LfJjbKZpWwCI27s7+0q2l2vdPxnmGDftdA02N/
Ki+JVb6G0CUl9NOen8nqr0azGY3YnePbNUB8SUfSKf8Jsc+8RpXfPelaQlw8U9NBbCu8R3y2NPMD
/NuDS0e3+rlBTuWZ69AwJo0ALnrmEY16QT10+T1L6wRz+5lI7gOSjWLln+tP68Xdb4bap0Nzjhu7
u91UPsu4UlkMEEtg16jK+hs5ybRaB7vhxw9YB5CDfm9GrxOgLLsCkrQQPFlMlQlYRJ6B0exLiQ7K
sNt7VjygwmEI+iGxvCK4AVF3hHveIPSDPY4Ly5WdhD6y8K3opt7dpua/bgDIzmggv8m+QgBOLK2l
U+4si5s6+fK8pK5JLrk1VAB32VLzQ42xVpm1aCct/v38E31jtgeLaKd5qpMoau5/VhXpjxLdlXq5
N3DiF0X8XfwXW8m9h9Z7sKQCmFZeWug9bLggZuBKrM0MaStHuD0qsYmZ2ElS/FUS3v23LOwcbTXx
rC7Yhn7spM/aOtILO201v15gbMwrcjCQRwRz+4I8ll3hN7vAk7Flij1aI3GqFaOQL9kjbCAxI8le
/D7RLi/T6AbvW5FoyYj4XE9zx6ZgaCIU9UHEPnzoLDB658n7Cf1KvLdUUYbgQl9ufBbVHLSYdIhG
Z9S3qvYpmUPUYEK7BKuNYFKQGX8/v6Gy81w/NjOkf9ztD91YH9JTbMN1I81ipvn3OoIqmvweG//i
i21JCjfnjuKxFyFmV4h82r5kj25HB81RuyUg3RdlPi1oXxc4UHm+H5DiLI8hUtMLD+pufLwCzcPC
KWaWG8uOEKk8+Gwrez+R82YK1TQOwDEwwFtdqky58O2XVEcLHa8S0mih5lO3KujweRqExy5hgB/4
m0JC57GtH8RybFvShCjXP8or6QA95Qg+o9HDH9rOPF+RdyMcFwKJmMWdOOQ0rjDdIg4NEwleWrzw
AESa2lYeipiiepgdpHgTOH8WfuA6JzBRCFyDlxy7C4Rr8TelBVcWu0NE65LuBdcdR8TmC84KJ1c4
PMudzzIZFJPgGC4J4B3GI4CA16b5tVer8I4l8aYPHUx0FxiDQigXMEY+fdkx5nFOdxiEqQfQfqjr
gsZ5pLSBKvzZp8ERvEnh9++OcVgi0jeB+km8KDlTxwbEvDLDmmzbFsbN5bog0to7W09EqLWQeROv
HvevVC4eMtsuHzPLJWjssN3r335HYutHrrYhkR0KAfD3nNqvqp3ZPGPcucCwivii1EIiBE0bgcjA
sXj/74jY7HTQ8Pi7FtqAjimq2L7ji9FJQvQhGLzkW6uwa8apqRQgL0PQ8dLMDEbMOAekGjVqbebD
v4Xr6F1T7ngY8p1Hv0+BZRqJBQB+7c70hSFoylCmDV0hy+TMKSc55hlqmygd+AlyhNMRRyXe7mX8
+URbMyphlu3qNY2ltPIkBMNbxFoYAX24iV6+PeFdM1snLLLrLD5mNfNsmPS2kyJsPBFpovFI0e29
w67X67znL9zlkKcORLXzPiWnZSXeUkFQKMxeMhJTMDHUsAqLkHNSyjL4tYjymw8DlsmS17O2+Yor
ycbS0275OTnBwfDjgSP7UVRCIGoYkk/I3xc46Etx72Hh7tMIvkE0+5kuwOhKWkvlFLaAhFaxQ0pl
tKw0oYWwOgKND1COxS5+XDzAkHI9zIPINUE0gTgQDHVN25PT+GD7CSH4xafg+N7g9y7JGnJg0ilw
BLyDhNYgBe7I57q3hvbk8J0uV8l3dCVOLD6ZH4/qjHqQ7qDOZtqZq9NI8OboZWr5sc4+o2Frpt2m
Vc/p+6ECKkLKmsisos/6PTAX0DJSdKjjksnI1dbY1SNF0gaVnjSR9GRLjTGg/eLozsfn9vNb623q
lnHGYuopU5WvCc5ew6bG/wEHaVtApkRe6rllBeTJpCQXrk9ePpxQM4uzxhP5CnkuC+OKJoTc1hAu
GNSrBNlYYh8MJAZgt9t+GjDGzfYicDt4ErjPL4kH66iumcFh3RNTu9U921K6JT5k435GUIxdbCww
wYrGDLdfwrt6NJ8SN7N6CSvM0oYTmZWn2rQFQ7pBfZLt6pZpG4zNGZm0vVhLoNcdq4lvpoFWUWES
wlt6QgLICualSCmNqDBPKhhG3l/u/s9IRns09EAEdfZTX27khGHVoUZ4CGAl+loWbFNqiohFOt4i
qQaENZIpP20CzRp58TCKKS5MVxJWzswPeyq++MYBji6jrMa7129bD+ZVXEiiOlH3RTKUcm90qpx9
yabKMn+4oevu1XpOmvBfrkXNvU+9FXUzfmGoPQlrL+7i7LKEJttNeAMT7OEj+fHldf7yW+FDCUTt
pBsE93vFBQrHqUOmKhHEWMgEMpY6oHKRGCX88dDcLZ0qvObLBGJWVZFnP71Z9Zz1o+Xfb/9uaIgb
PuAN1GdH3CG20LQnmxym/ZRyBj+b7jYGlGqITTUL0152Sqyem2tl9Vu6xQHyiDyWBJmHHehB0z8M
QEC4nKY8uL/CiiNJLJSnvO6I4QUu/zw1tTnWVeJYxBF0VvMomPPr1ErOpnM7fAc67hf9jMKzJbIR
QqEGVJpJcb/7C6Q+Ppr4sSuB/lxqyKZ1S4/uJDW3Nk3H7qxiLx04PkSg9Cs5h7OuSvsPnYsn23Ki
C/gZw8rC/rVSXELPYf7hym6lDc2tnFCqHMdOembHblyhKFoPsL9BwGFpSk0qSQgK/TlJUtuz4x6V
ioBiMZOSV9cM3q7TXRYAZOzfHWnJ3SLd76gYFIx+PKa3YzMw7u+vcGG8//zsTKvNqgZMQOc4afsl
anO0bI8AeUETpNhb922Lwa+VEscjsaOLrTlXL/0OC+RKoVyk9qoZdzt/C0PzFuZhFhl3GRGGIqW4
MpNSl7zrx93oRns1E2ztQLfJ2/1MCbuCyKmQvFZsiACKOzivZviGN+4AvJ4GtGdXEtQezm+JRMMm
czWSMWJm2BjNSeKXclNJ70DBSh76pqDpTrkrZmY+N8F/Pnt6hc795o8ZYF96LAy8HpoTahrKYppk
IqNRGRWAtYmSPN87k6AoCv11O9yLlIdtlSutYMuWTEWqR90q55nwRW5yJGD9a776xWhHKWzUPJvg
IOZQYYe/pmKZwSool1aemUWSX2b5LKAXvyuyNJ2Xlin6BzzdiCM4uCJdZEuR1w+78JmVTWx1HD4f
i2rR9aACXM8e22N0QNQbqvTLkE6dofIp6eA3/SMCDtO/K0kr/taR9rvXE3y4S/ezN9GHaumeRs8o
t+mQon6EtuY9HQGTlofqj9BntgxiHYtvLIsuLBSqBCjTsgVnzbfRYYzfIZFssfZqpPr4TervIb7Q
qhTTXuWORitjreoutPZpCiAA0S1Vt2XDLqjBWUF1E3DUSK2fRgJOiB8Jqa6mELTXZ96RUDjFFTEU
wGCSmIBXOmbqHhpCIQSqjNE4gx+1I9bNJZjQNuDwAbDEM1ZjbHtIz+aQdrLUrGtS8g5Lo+SdoiO+
rJO2KQNlcNBnPZRcW8+RTEGixJQbAceEd+l4itfRm8Pd4Jz9hL3grzMoqotZ90f716qfdUNf0aVF
vrGzBnsBXxC+GbJhLcjW6EMgUUEyBE+VaBXU1SwurNH9VLYWK+ZAJ2lDZqKWi5jPFfO6godcJvVS
Ltu+ooo3k39M7Y2HafufduHYUWWNhYNGXPeDI5ajlpVZ0oScgkD4QwAppm/ZFq5TW2wxOW0EfrBB
e+rWGG70EKm57+yK2JshuiJ57OMZIcNVFI8/4xDaks0gl+cEZ3C7PoA23v7KJ+wkqHx3i9meKUIb
Kgo1/Zhmi4LDsXpJyKeiaALfJRseaFOhLuRkJzrVHLrAnDyR2ujB2AgJvxM823tzVVEBI2xvQo7P
gwyc51Ijnuw5F/xaTw6+7YaOLy2OhVzQln3uL37AheJrARHzwqFVXyqhns2nKMN2Y4ktLWMPUyj1
DPc+3qwc1w5wyfXmfbHnJAEcRKt3HHvcz9apYFoIn+NB9Y3+SNcc+kBFFONgjbVN8/Gm/8rIGofs
J67t5XBVblf07y/W2AHAu0/OLZjI52lv14EXr8zDYGkVMJSekZyTnJ//VN76zHzS79dBNlcqgYtf
3Xo+0RNlVVuPFFWSiSgsayD/WdpejgcqtriDBQHfWMaSqwKSZY5RYABJa5tL6JU612ES/S9KbUX8
rPjQo58EMqhS9w6HSvhLwPL98+//V9JL8rHMWAcqoL/ifAwdeyV6dNxAuqzGeazikltXHapKQlI3
WOUKlyw3xXrtQ476ULURMlolgcWAWBmdc0E8x/rmPdVuglyrxnEir+JXP5J9yb6VjgnN9HxC4q0Z
8GMa8PeYl+7pjCc4hrVsyw0guX9zXuLStoG7JkWR+faDN+W6+89/7qhUlqcaGfDAuTnCvfgOLVyG
Mn2tYxH+FhvfcuURJBTMaZ9ZCliU4HgvUVvI5pwVfls05aXN4zrBJ6TLnfisES9YeRO9jaJQoSF9
hVBNnpzodx5EbYmlkQeE1B9rz6I6+gFPzLl+G7o17suJ9H1wSd1uRbvi6ZBmRTUiVGNnJ/dgQgWn
UHOYgpwY8UUFg1S9I53Om2aFjE41F5+PBnYSWLdho0fRuHdEKY8wxA6j37MMZMqfBzEdY4itTbtU
lm/9/zosv44XtoXBELNOUSeQPyGuPE0dLKrMg3nIpgJEGZGbWi+kC7u08myNwxecpa0HHibSUYma
j9eRnkQoALqLfg1PbuUc/RgOviWna8k1fSy45CdylRzLO7+YTrX4aIjrg6U+fvypJuexuSL8I1Bo
HAzqU0VEzgW9giz0/6Cb5+uRGNV2KHsAhzrZN33zZ5W5dpe3DItCWCdfTvs+EmxuGkIa0k80IC9F
mVARem8siWg5uNwYET89vZyn89Z82AeftOMSEwws7X8dt5wJ9s2IMZlQjR6YQ0JyZXS0oPkqKJ1/
294eGGLdBy8rCsTc/pvjobAezRyAjPM0lCFI3moJHiFklSsDyIImTSqqCdxDXCO3d4NBciYp89P4
xXhFbcmo0rKWNaIxjEYuIZIRS6PMf1wQjnSLAr0l8wGkzc/FnYkD4KJn0Pwl1oapZSt57FSdDinc
CPR08a3EIzi7DY9wGCWyu4hoixSL/qNwpTtHcSXKnx7D7cOiF996LorlPZnNIDbfrEBUPcx4Hzm1
dWNn3qQTNxiHEZWLjoP4o4hhu5fZ2crVjL18O80VoVEf51Wc/aBiz7FJxnw/8AmGbgu9PpbhkXcC
NVGNb2P3tMJ8wQ+jg2Jk2yECQB3zK/0i0xvWpnaBf87De6FSJGpOtJ/KEH22Y6M3RNjePYld43Lx
GHx1Fs+485k7HnTEy2qpT43WMLIzT7VNs8tO43JkPMREuTJ/gxqPwGQgPSWHvUf216rgLDP6LdXl
SxwCoyy3S0qlDA2m73kNrOswTep42B8e3EueaMc/bWZXGZiSjpMIGfa++69V76877QOFjxaAnkeV
X0oMv4pGSwBtm3IVzrRMRzoPs0d6mBtuJJlGgAyVWY1QR8AkPyWT4ny++m+K3hDTUb8HFumJWh7r
dnUfL0cs65tu0J5TN4BAJTpVl8heyQkQ4oNKu9eKRZYI/v746qohPmu36OMpyuNvDtFR041HtcJ5
PT3iQKDljn8B9YfCnte7W4MKL0cjWR8rJjZ5ECajZqjiSRU2W45pOTLbqZdVTMk/+nqRcktPjNoS
YUt9HZCbD8K9q3QhQ1fH+ee0g0kmrIDjmwNcWKA/cti7zrDkSsMLG6xYg+hXigpaPa41SD1cYOQx
DMrQR7NUgSwsb0Ys1idXjwgEcVYlXSlpbnbHV/H2es0WeqWL1pUCSW1utSYg4uwNDlnqOkj4ZjMc
CQtYmn9VGsP6XmCR541wZ2iEWU6R2tzlgke3qIMDtTh3rZsnTk7TQnUyZlZXUmut8CJ/ojjNjObL
2iBVV04mjTnLbhkLGnb3S/7/ulq5saQ6PQTkfgSDtVVtkLXQ0jnOBGX/ZP3FGo4dsZUe46f/VKai
3r5DXadp1qX+vKm3e1J4Wyzvgam1ay7HuDM1ytLsL/4kNBTk9rA3srMJdxSFmkuuWdKfCgBAmri2
ihv/dKfHjWTVn/I3Hrpn4i1+pnir48yyPUgJ8PwXvZYarfxl/tcAWwr6BXOdYh+QL+6qXG6WljQT
RpLLYhurQRzBOJPOkpvkOQu6pcBwK6Kq6pl04c8kOE0yv5oPa+zRNC1o/zn6Iig6lJ+e+2dtZVrT
yU2oOc9UPB6+y64xULv5crbWKwUTyTSAYKc1qnbHef/MsoXLfpbfWm6wF7oicCP74Px+4Z6bSMnt
iNPV7pzlQiE8RBBR+QUirHoeI/7OY0+KyoJL6p0YEbvLV4HP7eRXfw6EQxwSxSF8uTAcwl2a6q5V
chbgu+qAz6xP0wTzor2ZsTLrVEwD+HR6YIRdYxRAneKWuEC/0/+DQV63K8AHFQk6PlhAzlQmWIDk
fMx7FNfqxAeFiFiFbVBNiV7tG7gLFcOAjOvqLwnx68XdAl3y+vztjUoXXu8kysW9uBCh4Vq21J1n
/BOqQrSY2YLYOAm76Igsl9yn/VJ0R+3VejXCzp9e8UYOwHDwqQbKKhi8ie06orav8waK2/jCZKyd
ehrMa9V01XVm4PyXORzTrmJgq5L82oBeHpKeT8NSp0qNnyfU2MQsd4Glw0GRxrnygQoHbvR9tr8v
oHUxIc82wWtLr6jBNA7R4pUk85UxdS/GOV3SgegcPR5fybGUbrph8xzaVJfTtkjfrJqAsYB/pA9O
CmImeEjed33ZdEWLlBHjlt0CeUGZ32UXJJwQUKtSXpc9gDgACZRtkrqtbI6yO61NOWb+4X+QUI7r
M8QtIl0V9Fu9LbGvkk8xuVrwAOXojcrQ9WXNOHa4HN4PtPlpFWt/nZibDru2bsGmyaZ2WPCa8ZaQ
TJGlUWfH/iiwbIanCvpvOKnqDD5GRlLex7YyHBtO/VXiwEyf4LysJXu1Ogpz/BhEAfEMTaMVbZVU
a/c/75dz5+j/31YCuSYAlWXdLHktDEogMr7GrVeL/ytDUWdUOTJF3LUGNAk/v8zv98uteSFwzhDi
MhLERIHtgHHLHjyAykBEWadphcsrmj5GiBmatcKMv9AibeGkohu/ML6vJXz8LNj2MNQbcIHQwCcI
jsGfeRf9/1zRn8eFchd6vTxRhhFAFav77OJSWqWRFcXzr1quTofxWbIyhJ1BnO+PPQ7MSWzy+6Yo
gG7sbmJwEOQdP3INbV0QbP61CZnhFk1tLcBe+RO6/G4zZuuvzSkKHnY9uZW2mzH5NYakj2aiWJei
Sq0CIrwIS15mxNFtmz0n43SsRLqXkEgovLi4upxVQ6LAQlXFnrO/fxS8ULbNYkGTrNNLsH7A6x6j
SUQYqFNTbfhUkMZf27oKgAMIS7RwrE1ZCqnBVHwH1njjXMN2ew74WeTzo7cBx/otHXO98bqMTUp8
iezq5Y+CFNcrrjAgY0rcLP/a+pDAAknzru0EMgCCLdEJjAXbMu0CalFEY3cMD292uRqdxg17ojCV
ClrxYFfSbvSPewAQkb/XjKkmKfQKM2et0a9mlQo9OrPHGohvT5/t4qwcMlAvMrxrqA+QJh4Z+AxT
kMJ3XT4CsdA+kfCszHEXMwzUgFXkTgDMtF2affR4GW7blcEnWH1qHGnS8slwVlCsKrDN43RujH05
qtF1NdtZff+dcVQ0PH049VXJlMO2202qAaFE+FsKGHGEN/z1PnktQ2qGydWj8lIp7sfBwtnx7lpP
a2sGKk9ynJaqxiWyEyXNz+Wu6GF7qPZPe0UDNW7wjDwBxykmHkOJl3DXym8o5m/BD6JGK/tsJ4Y/
BjGQ6i9tk4LcW0imE6nI33u/o4vQr1LBKob+d1vt8o1poBV1dC67Fg1OOCTQUM/3wLLcy3j8cjBX
6hUtJwOhqnPXFpbXADrN/xU5G7c7bkihkFCyAA5yXXIGJXJ9WvxZNfFpwJIupY9XZ2QkTYj1qf7V
cBnfKcOYrsHXtRkTiBpdTPLi579EPf7WGyrHpvpB8ZE80/f9+Eh87LbsQLMgZjeLRUGmvMlScxjv
b/eLhiDft3g/C8tVtZB7Y9EiNlAXqgYpzQrAx0kZuC2lZFFPdMyxmCfBq2Tz2WOIjdp3+zfPC1u5
ugpvpOMGCvyunsA0WHr6nmoUSCjVMOB34D3zbsJouzAWTSWfo2XzaI28A0Wym7K0PCto7qJL0jCc
EuNy2xRgczxJ0TL1y9GrtCjSpG/UehC9yb89kjOqDCBpFPain+gHoFEkIikivDcrwFG94wm6HW28
pxEDUdo65GaJz9zKD2ziLsYe20zMeNlBMYOp7sf6aio+IOBugIXs7lwryc2YPoaknGTHvaa6ny/9
vGXGhOGluUEz18jX7HcTxtLpRU93smBYsVeS9Fjvz3570/GUg8PHsWB+KzBJXWBodaIkvx3+Xj9Q
Ki+BqDWqJz78q8f1YdWh52NxLNDDAPy1E594oAH5ht3cbfajV5ymvX0BMidRWRbrxWI9aSUVrO+4
fSBtSRsBl0XYtLDtgXQgMDE1cqKP2njA+waho1v6XugkfTjxxESbTb/WMJ4/luXAxhpyhjaR2ByY
ty8KEAtpUaic7BQHqpxc63aVCzEsCJuQDk6L4FdQfmnlV4jJynV8MjsNPbyU9Jria2JdJqpEFS6p
2Bi/mfKZ6k6gXTOudllBEZsfl6t0178zakCOaUtLVce+Mvhof1PVww0tgc6hfO4Fpj1aUK59tg2X
B9PvCQUSJslTJa52x30IEka/ZOcNJn/Vt3G41ou017nmWN9RoCuZHEcR+Q6y+AHSGFfbqTdllwFZ
rxeU5WaW8Q07WaNHhKfrbJkVXwY2Cbs/uml5p+gtt9Bh7e/4gsbzG3gA1gT8tbx3UYRk5ey9SFuo
pdfH9SlUweyGAqnbzZ1ZRgU2vlI6EKQpUSkqiLKbYx9iw3dXgvsxZafNJMEb/UgtjXlhGkagG8Mo
/tOAOdVL4VpHowF5X3KpyzqB7TaOdWu8J49OTpAnFRtE5usITPgGaZxHWtPl287A9OZKJOfHxbOO
m0r2kLLzgSkorl61wRcvDv/zPncfQyx53PQZ/1BhVZG1bnccjeI9QJgFPXo7WK5oq9D1no1uKWo8
bKWnwDA31BBAffxzBzBmKPai8jNvi+wY1fEZcVH29cAUcV3tvjKiROQAQKSYrMvv8uikGxxUKJEU
/RrcgLtjCBa8dgV/j9vnzOH0bSCZoDqchC7RG8g669uGcv2EnUF5k1b/XTZ+GmNRVBAtzEOCfh1y
J/A0lG8nEkvgwTbHpxZ+vwm1HAzPfchX9fRVaDyaoPt5EEZG4dJN5rqTBpAc48YGqoWW2gSSe7GW
FS6nekwsLVo+rD/SdOtHJwWEOsA8vSbVYUHw6/5h9goM8gbLMRJr5E1qhLKWV4YK5Jum58Yora5l
k6xtRuA272spiNwuw9xaxg/WmzW+hH+tGLGeD/KlWKfzGYpwqIXOe3n+/wEleLGcWbUbQwHsv9GW
3u6OcPHOPjAqy/cgnPS2W+qdHmc+jvk6qoYMgYjhH+HtzPG+4XiafMyGlZhipinT9iWxaNTCBnHn
A5siwd4vTmXQrsqGm69S6mnCb88mPDwtG1dXRHOTTyZa9QwsthYg50Y1dQ+UmOW4p0+xFkRFbMfg
BOLrs1tiMVWAXuXqnlQtrI8s5GpLrgi/ZEacGCnzS74Hkn2sQDV08Kw8KnRwa2pMI71QBxt/efBY
zq8JV1dUpcf4nlFxJU1+DX/QqLk8i+KRNU1T9HoLPZN7Cd37a1up4zLnPQFlSWb9YMkTo+Cxody/
AmTF289H+qszlfXDgrxqxpkDrzzCmGd7MqOPgbymwh/DOdywIurTH1S90E5FfHn4RMKB7Bk7Zoh5
6kBXYhhRTxX1ueo0Y/altH1PTYd61hpc0/17eXeIwxUyUpZz7MZ0KlnBZQBE6oVX3a+ZWT9g/FUd
Ie9LlJmO86lL9EmB+vWs/WocOgD6OKsvSiaSvOB6w06qeWTxs/U9qUxHXYBuTMX/vcB3gjKJ7k9A
ETOIJJtD5ti8CPbjE383eWyf9skPJJD6W8vALZWzCMo1cp0nc6QE4+drOhwP/e8YDE4vOkkVnN/a
rFHB42vKorubUMnTXBpYtLmWgpaM6zyZ1JxA3zESZAAwBLymvy4TwxZdjy2ACfgFwD9JPW6W9WgD
ZLa9en23RSGSe2P6ldZsbPJA0KiLKlslmYcX0ZqM92/5kgHfXewMwqMCTEqMqG5Yo2sgX5B0avNt
IH2JyiZ4IvvtzzuKDpmbySWG308ztewEubV7fQwT61B4vI+mmzyd+EFnxC2aXfEn34f9yj/hxqtv
/eksn8EuiG1qlW4MGw88jfPcRHlvhCWMo+ONrOrw/+xipDaBz1gzTgwwNnxb1+c4OkrnVPPUETrt
c4QgGF+NeudOjL30w1U8/FMy2J7Qe2XKUZcQHxTt8Fk020ar+EjGJDCikkb46KK7SZuxi74Wsl/V
bR1ZwQepPh1Q0rgMTpLBTdHHl2X+DDPH92CZonUYVWCAyrdImI6k/km0NeJrVeusm09u3/ghCuA3
h+HlHONSJzn2m28brIzIfojJohZtbOtlxkZ+0vMBq4AZcwPQ1sZAdNRuVNyPmfO7ZtuuG+Zvk9pa
BgTiFe4fSDiZPuskyXE/AzMh8gJ9P3ShiKadqkLKtwp50WCBCOZd30uI/lsr4AOKkJVUHE0WkcED
FM0ptKMUi9q4OGMFyEfrOkZk8KZ/d5yhcTWkom8neAteP2FNdDQc/kTNABJ0YSJ89mkJjwkJStvy
IFuMsiguA5Hn7q0yhrGvgEgFRjoXv6tbZ7eoCA1jZu6+AcukcV0LTerpdWYjwDvE6Lz8kPETHNtH
dFn2tOp4uZYT73wGR372cY5CjZLk84AognQCG20Pwn0/kXtQoO5zJc5bYdvAX6hqgRtpnfc3q97N
eWJW3Z/5c392ihyIBVo4PvzxoAuv5IV4jocKlEICNS6DizVvdX/3+VGVm4+gxIEdH+WZ4GgEIrA1
s2QcydOmHFSoG2Up9483YwHOWMFEPrCnwC1fkzcn/Pb7MU7oQpSkOE7ce173Spmcxznp3QceUKGB
9XuFODGbpn+EDkyCjLW8JBE2vgpG9OKhbSv3BM2RE17Vu3ROHUcBT0p36GCmjk+MRWXxAFFmb6ol
oCLc9OYWjd9k+55kZEk5AdeaG6WZ7oNRNLlGeqwSn+OgcAMiqZpctueSep+M/vtRGdByBWHTad4V
iin7DkEIy+CiGbCSYSToJuZlb2dx/T97bslOJW83QxZJA1gweTUxx9n4KZiOXyGblIAofxw9LLZw
DcNY6mak6r2WAEzl7j/pTYwPrc3hQy3ItC3lxEgvVuvCVyOxH7CLKXCK8q/rp3ImQe8zwNfchFBi
O8L8DJp4AEf38afzOr5zrnnnOjnd+x4iRVftDylzyNsMYz2q36FTlYZFPVR3Ms/fQpAsFLzBhYdE
eNUtt+4ycqu0kSUno9CHgln3w9eaqurYqsUMCPbLZ8P6T6l4kRbkyg0UksgluGz8rXgwBEfZt2Lr
XvruH4DPmdIkwUp3fToGvOcM9z9VcWZPoE1d5AwECzlOXxFSG+rBkWRRZCKfVuK3gbUM8F6Nwo0J
LJyfd5S0Q1Q/jBNPV/iCLdUW857Al1lmQexPFzzeewskWiYfqcI4v31L23xoAsmMiP7hGti28zQ5
YQVUUInFJOPPippKHPcLtctXAKRmfYhCA4dx8fcLb6fFOWA+ngYmpPNN2ahBXbww13zH02aLqyrF
iGqwbKKMkSI9WhI3ZeYd11s4wlI0kIUF6J/Z+vBzec2yFkvdvD56q7NrhbCgoyIXuGcfFAgPVhN+
rZ+Sx9OHo5gydjISn+YtMNcEPay4R8sCrYHTcwo8Jq3zANwohETt2Yjb5j83smSuF1sBnDC6LkQK
SlBpor1+B8DHr9p960AlO4WZTd+ZAojTQ5q9+MtL5fLToSPY58PtjoitmGUEBJpAbiVrsXpbwKR2
tCYUO+7Jzq0phOdAgyHRdvWHxVR/kEykOTIErxDXtQ/NEwKkPaSxMO4DH5iRQH1EH6UW43heY9mK
+XAsD1IjryGG0iAKGnd4tPEb3YKfqxKcsSowraKJzFqo48NQ1iDjLpupT0gAPW3orbTKbcvsa32C
wgiUsDMZP4MwPzvYZMyx4dxj4dHMGODT4TlJH65AhPQpus295V1/6fsCHPh6t5q/P4ubi9GHW5ig
pOK1Ek8bkUKsDvfywdyg2VV5Ia1woVI+wozhBvb5bxFtFzz6QDUpp8rLv1FBEehq4x4DtZELaV3G
HdVgUUok4MSuXV7KCrJ+EoH9S7HqE48An9kPPCyRYHn2c5kOmSUDy05dT3NIcduNnuSJdk0rqg9I
viIm5JFE4Oup44bdS9Qk472GN8yt7OePgkfFSb9jQLIzDDvuUJgRqlrOIz4HuocpH6knVgsHYl67
RazVLVk+yFpPDgA6Mf2f3T/JFDYz9qfDMl56z4fn6Koc6bZLU0nCr28CSXe8knw/S8tkeNtCPAAR
SCV4O5yzmlADNVYT9pHfWhdyFOrdn+zWbQ+JFxUfIy/8jnsa+tXBw7DspTwcPE5jw+QxV5HOiQXB
5bZ7r0cUhz7bbylX6S3NXKq5fzd7OFL1q92Hw6j8yXY3Gi8Pq/e8eZzpWB20JAMKUDIbFa5y75yk
ntIsANWBx2vi33ivR+N4sLyPyXha9uWZx8bL2FSrtLkpweQ/SjCX0dJA6IlZE3BYEkCXwyxhhODS
gvDJ1ZuGr/bAUZBe139UZIU3GdVC1RXdZ0WDMY7Tne/a5kYGkoTQmuGV7T8Ek4Iy2wvN5nbm5Jll
BK/8405tUyi/ieKU+lflkR4Nvlw6zXCvKVrUUmQ+9wpLJ23j3wHvnB918yeuT5lSJ3jpp0VlgSxJ
rx24a44zsKMqll3nOPPmkHwwYfncjoctJWnCJjpdZ5wKmXNA9P6l0egY1y85r5jjzqiznxBQUa3i
eHzVtl/HfftLviV0N/ZPB8ABjRFJsFuxaOKF+ZvzTQPeDNS6FqB/7dufX2jEyLvr5JWU/RLMyoWq
CIaM7meJ5tYy0ukTVMdCAylAQPtlofUICCcf8CIeQI8wmFD8osvd+/lLxv58OiT4M8SvwEUEGDSj
ML2HpyDV278odoa8KcfA8tVJzGDS5eyJryy7TsOa8VpxXFQsTxqcfrbTgvNnWjSk4eSEXoRExGzJ
Ad67cEVgJRlB7OoHI2DFiLCWv8ry0v6hyA11yoqzOtykFxagU4gW4gAysKc8Io3xQj5Y9xq9X1CP
DDnRNjwhTD0mPz8z+NykMMqCv1RgRCRKev873b3pWZOSc2CTIrCrI6OJcN/FpWgZ6saXhaZeM5Lx
F7hzI6HeUJWya6yrUjJnH3d6LkT0CFLzbYpDntskNaoUwM8vxYDtWsMMeNlZT5O5jm/TBUwpnEcS
jlTYgjF3/3ABoY4MD8+2pvycEiSjUAffM+lIvKIH6HVuuEttJdV7SvcKqSeMy4jH5mNjfztOEnYd
hIbdzvRxMSi4sZlMfHMtqCVLC5P3GysNVdZTyljgDXDXcRj6gMstdod1IVX43vJ2zKoUeBEoZJDO
Wrkre56byA9TM8K88h0jORDJluEFzCDzXAiDXPzKw5IwGb3LvZ/Y+BFruzYzV9Efgnl0E6Qk05cH
lEohJbbhOFMF0vs8H1cuHWalIn9l05uagh1X/7MIUJ7AqNUhcBqbFjZUUhii9YfxCTy4J+7kUlrv
tZrRRyJ05fcUUMl/tJpgyxI4iCMyUzkGrga3bbz4Gb2B+V2gssCzy/q7FxkalNPt1hFT8yl8YsfT
+Iv+GLcSnIEpVbZWi31Ckp/pdkaI+rHQkQMl1uzCvDVce8mB3A4J+K7wZfQWTOgvO6D5Tmr6vvQG
SVeZURCa0+rw4nbQtpF90VbMt0DBxFCXcWb3x05cVm1Ew+Wwo1ascjsOSRrVUJ3YwaPoz8ev8POr
efYeaJgMt8IenjmbEaDZ+KSmeeQeFw8gkGJHhEqYIRZtg/q1KihDK8CuCqbsluAEkx06pVjK6Oos
wz593CGyWgNJuQAIZHUBdnUXNWvbUqZfQHJSjAGOZJgGkPqHBNceEH9pqLByUMcRmsFGLUyI+LR8
zEGy8gezD3bax0OWXY9tRE2N5gRl+YqGijjin1LFIl8VLWw3vRYbhKoc4fGDXegQWf+o5Y+3dE52
2KU/BfBCc37pFnEt9VxRW4ohmxZnyfMtGBl46zJEckMDlI2O7ArGiRKxnnUXb4Y3pOTDmMmhIevR
uByWAOSCG/T58cqX6IwiX+etkbaJok/LH1JDUtYkMJ7BRbTkjSfbfUWhbZGpQJXs8rU48Cd5n1yU
p0e3XuF0oe3vYclJ3YfCu7N7IihsT2odOaDhBfQ/3fRGKfR8JJ6o4Zcb0LKS1Y+YznI3i0PoIMbB
t0Jzj8GMU5s6XInSPXN4qOyLchwcBXCcIKeAvpHeGttCNK1y+Mtt6jOHN5xyIp2vRpa10BhVgMcp
tsL0pyBI5lkGhWP7pxa5iAVhFfMsjxQaTEDrlYiHMcQskiq0dNhyOGLpR4pp++yKAKjFexGu8SVK
0Mf1G+0Y3q8n9+GOaFX+0gFh7EVk21aO6qEyiSmwDgf0BofKqnPE7rjfLa0fDd6lYIeylUrJuKQb
DtZ5XOfgd6xX0270S1FR3TPJ7ExS+rkD/M9/UljsR/awT4/ZuUrTIJLatnw08DS76+BHoXIeR2ax
V1XlCQ2bwRECgUdgkfjw2Lf+LGW2G5710Y85CbRj8G/tvvbacywVQW5/mrrH2LB+9CnxZYeKymT5
mJ+0enmt3HFwpd89mijWZ3t3KJCvT/bLO17j/6XzNJ85AQUuEHssj27yxge2Ohq3hsZO3Xx3Cq05
05PFzvLpu7QeaowTd/JGjqndaLOzStWP7BFbN4krTHxjZNGC8rG7hyZ20hvv0wKoUChkOURAhpGC
Rldx+0oHagABdBw2L0Z+I1OsPVwjBUVb+sBpKSRsoY4HyIMXKX1lLCuE6KlLe3l53HLXMPlCb4uP
EjZb7fq1sRIIKvQSmpgypn4U0EMjyo2pgyspwTCQhyAmssZKewaSGmgjrSsv106mJDuhO+xtmaCv
BnnlaRSSTcF346V+gb0gP9BdUjOr0FkfDbBYXY6hMCSGY1SWxXH0yLELSG4Eyy3x6f9Z5XNrgO8n
d50a2TbNV29q2fW1Uzxlv43Dw73wU/kxL+VqZCyCv4IKu05MNsE1xd7mz2NGHKpJ3Wwml83mmhMs
QWY7GKP80K5Q8srHurLL/boLAoRH1Kq6Y9acjfgVWG681ocee2hfaomEM2JQdRXBDqm0zoLdCk9T
zgs5rLfctLDYSaFUYFKIHHsuA0reSSMkfMhWamnqinUlpjzfBPLRlpqOLnjfYiSxs6vr0Hg6HFpP
JZmG1AuomJeEM6Bsd0VbK1QUORAEfGVmUSp43xMTyHv77xoiAxP6lqwbe9u7LqWqFC8PSwMRsGaI
+2lvubGFckr9siR+5MNDL/T18pWvGrgv4Uhf1mWRoO9bzEkb2eGyyVXiOGaDRKYdJOpsy2TRFzyr
ff4nzl91AIzpQCpIwyog+sF0Gp2ihrAuVRla+UtSrMIUxN/HGgo6exTbmiTiVMaIUP8Bl1BurQmV
Eu/59Tv/fz/skXwOJYCn+6/rZxPS7znWu7su0rPNkVSqlojmSmNV+IS9sZUTTyRvZGZn8xmfBu5u
1mOVl4N1SG8DqSQeXBxBWvg0EURhMgo7mmxt9FbMl+JYb0eC2Po8AHLgvN98Yx5UaGw6Y8WWjxi7
rhyo959AWpYePbWUFmZJIE/KhndenVoodtFyuqEuMj6+STlRHVr1KVc9fMGyGaZwgDgXc4L+PE9x
TXyD+eJaO8hJht2PtCXlYdLJQ0PL8SHnQJFw1uiHWsFfCaQDmc92+ozVpwaZgcy1UfDr5vRKDCfu
VFSwlew9O6/+g16eJTRPKiKzyg6FVw1mPg9N2ApWbSA/mNEax/eaQFy/jwE1+bQJSV5xPe07edHs
F0RfK97R+tigrCOQfGIRF0uA7GAEqA5su7DNse6kst4HrXpiRcnSsKbzOSMWdl+LYwnUwLnlSJNa
6dqct9jkCypGrUMhuX4JMTikizmTRYm/mANX8RBf+ZoOlcXhVqPP65CerI08r7BU3il2YA2TetII
ud76heNmTW0jZDGFsyzoeQTOgPM9MVzJzENEcplUcu65IKEWrRjL9Iy5H+QOR8wERUJlHQ9MfDBz
PUD9BEaBBKWYNOkuTNRcQUzQQmIsUyydn/p1ykokWS/k1zmQQtlMjGbttTe4SuDCV91G6CCDUaWo
BjIR2sBL96HFVxi2iZLafXHVLJVKkMEpAjEx2lV/4+kiSys+F6AfC41SiVHXKqjG9RQG7bUa8AU9
32HY2K8oqq+DbhJtzs6PdyknmoOTwoXLWHtY61jx39MHv4FNuRNee4eMcNg3DvVzWNQYQPg8kuxn
QVkNX2f9Bxj/Awa77p3+EgQbUWn6CWoQ2oC3eMoh+UXIlstuVffkzyUb9QEUoEaXyUz+Jj7GYLui
4Lqtx3u3kk2/RQ8Bl6/ICQBNKGo7zPUkxQiFJ6it9dMGwOhvhUoUroDnh7L9MFcF0/nk1T88N7Wj
208Jr4dNeqsYN4hG82gjfddCWO3GIZHIPdSG7ra/g53eluIuQ2xpN+40kXqLcyRl5CgPOtKcqSGn
CgdUbcKVN2suLIS05Z/q9Slpm614l2lPR7V7/t+E0Rzt4JVoF7O4U3JPXwofDy1auRsAXUVONheq
0nNJqh4AtRd8d1ALqVJ28YdEmBJxqO0gh8yaPKDEJp6Tri42kHyTNH0+6gSfYsXFCDRDhtz+CtV/
Kv3L9av1axSLBa+PjP0vHIJrxzw2BuzCqKiPPUrKvBUV6S71ud+1A00UntASAaL9XV5f2IWDHbDV
XgvZlnrZOoLb9aiNzTEmLHcetriCjjIHQPpk1HDf5tcMqzPZlAVzTfvKrdWAqMDXQZQPJw9NLkpZ
279gTla5qrjiUgqbz+Ba0axuVkCF21H/QxVaqS4kgGiTD3EqoA83TjL55RSlTI0fZSIp3VCmbxcv
V0qT8P98PvSa52hzSv+h9KQE4vEK8Tl1R9+HR0R+IKi96r7vXP5FbW+z99gj93VIjXEMxqohnnWu
lGfFOejdbhaI2QD/q96vcp3wLblIW63y+CN+LCBm7FEwX3LNK48jVXu8qs5tF/8MtmLlTAOBYZYC
sEiYiw/zNCCG46iR6aefShd3y5ICrsaX6jQtBFJsQ8jg2VZKYcUs+DPmB25oS8fzqRqmQUXPwCuK
YnwovJlVk8mIiEO186tUeFtkvU/aQm4LnX57TVW0opy9HGF7tvkqZHl60kfVN758VAU3xmen6qMT
Vg9dh5Nlz9JxZxLa8dGj5M59V93UD1TkURwGV4C5ETvA0qWfIQWOXVQ2MfFolgIsEzHX6pvfVzIo
w+a4OCh8kC3zUd08xPQ4lznFxNzAQ9eYYBJrwxHPlSdOnu3EQJ2olZ4y4PzpYML63k29cVvU4vhg
/BGEEa6TQLdpSqO3+kYQ9P+PLR9y+1XdlrL1e8GpMISqDIPWMBEMWngP15JKTDo1lDWTtarD+fRO
TUqE88UjXieL9y6tMfvzxPw2bI/hIm1C1jsSNsaGeP7gIYb9FbE+5ezfZRmZOaTRILTHwt7UUlBy
5rUle2t3Zt8j/AgDvUVn/R5yOAcwlp0UerDnduiBOP2YYn2dyRSqvWCldsvKiC7dQ7Sd4NH0/sV5
59wrwCxf8bPOONW2IR595wQwKCuh5vs2xScSbid1LIr4Xkap4QZ1vUTXAfTPvTy/KTjiyZPtPFEG
NWiXZOBrxL6JIQo+3zoHIgPROHg6v1INTvTCjAVer3ohsq14wsaXXdxA1B0yZksQYLLTVAs9ZrjB
D2ieoR5Mtbc4ek7mXQrANGr2mQJb5LfMq8dST+BUvej2Fh1mSnZxc94B0IVBCXmGZCqkVZzXsvOj
BCJKo1sFRmHlPTTWEj7MJp7uP2Ia5JlbKwuuknU6egPj140tOYPjQwVDSboEoutx+QtnPNeayJr5
7EVkHZhdV6RsPv2AVQeKu53PJT1jYG2SCalqJXvn18s0Ko9tusHgQsuYjm/dx7nGKmSEI5S7mUlG
ReUnt35wrEt5Qv1bnTMfc98MIyfZrJZN7NaiVQ+4nKotaxEpKU9g4X+Vly8IDRPnyBcUZ9RFa2cs
fMRDfflyh308D78M2QO5LYSc6uwlto3gtGsTPQaWmhHSByGoiTr9jBWR54uRquHNgL6NVkblJLYu
IU3Wl+bqDy1ByDxe6GjcZroFvt/SCxquaC117rcK/eZbXBfoPVLVbHRtC8L93tdP71lHXskJbJR8
PjPq8WhF1T1wXCJtIOhDY/zxW+LKABznZsAx9/xMHhhzFK+eTN4VYgwIxcJ5XSELl51sPl4up/mH
Le4S4dYcbYwiHABflzPZSL6fEq+eK5HFTg+8FUGqQKOwtGl78gIbII+zdz3TvoNF74A3rFpJdnqs
1wrFt+8j+2u3s0HQ5hlcG31W4MtRmKj3YCsM2KWB0CMriS5SUMnrN6IuOJI8d3J1dCZKmdBRw/8/
yKCBw7vFuIDNhzNJohXNYMVJY7MGPfdoLrf38QFtd+iBa/uhUqE/0bH6BmDy7fxXupzl7dlVmNiw
JXTKFzCEEaoSAQWiKKVMXbruEyMTzsSa7FyCVVVzNWRMF4misF/smVhViASVHuSJcyzpJtLm1eiz
CCjGatTh1Zw0ZZY0E6IyxGnwmCcl6NS5DNUe0HcQTkwm1+QU/gzM+Pex7DmiU1mblfGfZqsHUml1
N9Aij+Xan8TsdS/t7prXAaJynPWhHXbvYY10JHAxJjX5JAn/ByZNaPTvDOTgnXZUp4Q3+Zq6IbDk
zyIoDOMqO8aZBkavC3Q/nBh34UQ18n9WtlzXFsBiqQUOMNx2fNNvVwLpB1ye37Is/8ku1AcZl/W6
pj1GAjOLuagur4YujpTh1wfyQuSI3a2acNHJdVs8PABk+NuK0NmuLH7McfZ7+N3HuvWQPu4Uaa+/
hxnJOxkniGRytCfszvbz16iG/hOWoqHh8z+WaY7S1U4XQWjCrw5Q5PDWuu4rSUgE9PzGbHWJiJOm
f+OOt9awuBIclEIeintI/X3e5zOKx3AuIqgN/3ojWKxkyxpKbfzXYptgdwqVWFlPOoFVv+0MKdB8
spNytCqnxVeT6g5+Ev5+/gzksOSS68gRlo4Arm6ls+LuFp4btkJBLO0SDXXDU4V2CldxWCDu1HK7
OrVLtBPUPjVgcoFi1fn311Q2LWkqAmPEGLEVBBkkmJ77mwneQKnrewEDgfMNzF4kmRDTE3KOrswc
f3ky3wwI7qNmYXBjDrf0KBELdcKSPQ7DViaRWjEoGXPagQvIPJ6g+8l3wNELBPU7h4R5icxHuq/y
p8SwXSrzHVGUPPqHdsXzTRVOdadyxAisyXJsk2/W+PEdrySZ3ogJNi4EmHdQkv46P8uvlxcerZTL
6rYB4/cDcrKLzT33fDISm03ViJDpTFk/62hYjixAu1pGRUiS5BViIyv2k1QFiNbC6UQiWpTwYrL9
x8KAM6fGa8RbRkmHzAhV+VFYEF3Zx6FYySaPpMPFdEexDEAbC2WGwrnN4tVpw/F1nDj/Q/haRqKe
8PnvtheoqTW3YUoDBncvgS74jHfkPM5ccADFLQty3QnzNjzbTKKzrWzjx/EaHeZeCiUr4/panVSs
7JptlqxjUFKgoWZKVqh5f49atDW7+czE++PYrT/iFCOVt6PTJXATXjLl9wLgwqP0PkLRICXUsVSg
T/lu7TpRRboG24tDrZEoowlYUwreqg1QfL7qkMyOLgQ1C2g2RMIu4fiaJKto1sMkCtvEiI+Yh/0v
f4TkfsF2GSYSgqT+pgIK2cSug3T/rcTLXaGcVt28qTAJG3vQsTZ9bo/md59nOUebNblKuLidcOYV
DAXTalHlXGQvwuPh2gE2RjNE7Vpe+lEgXyXtV9JjhdhNgCutJoyWE/PTzJmg2yX0Utv+02QRgVuF
qqfruvDSXWc9Mg0T+iN03n7cTLXHqUdyx4ehiv75s6KI4jsZNkgQBLOy6rbKqjftpSAD0dyKwmWF
KmCiDavbmSktPLrNhYwvqmbvmrC1/TuPsVpQACNxRaiSB4UUMKeTfVbVlECvtkISWeWanM0SNs/9
MFBZfDXqC2JGfpEQ/8rgZ7/GH4HfE2GTUZh+hd3fQGiOuVlVuZxcFZnJ7n+75epye73Yk6njpE13
OrXP1FDBCYfAnhVZRXc6SGKCb5wRdAs4oue0x0x3EKn1ZzBQOqYcU40obE5yB1a0ELtRM54Lw/XZ
ygikAo7iLoTzyikzqopSBPcQx5K16b/y6LFW9aFOM4TxDYOb7bNgBZkwxS5PgnZ68DOqAWoLZB2z
X926HZyZqz1gXarjUfDy4L6LrpbPff5fZHebUTJlTn2G1ueNa7KvHlvoctArGDEIwkZig33uEFVL
AhLjChBi6BlcRWQ4YGJsk8HW1T5KSMEJOfwu+gybBwMk//16NzNt2vB+usHeapsSihXceqDrrW5v
EUgQUiqgYG0CYyaAjjip5HriFeVvIXsTSYaWKcCOE0GbudJb4J+APbKY3utCrxxcrNChQbQlbxyL
uByCPpO7xAuvvmLt4qh0lv7Zw9jRLhTs+PQjwelwwhf2ceD77pMwzmG63k9NVjTn7YyIQ8cmMoS4
KH73HyLk/Xy5JI79IVTClgeW73EIZpz9LY3pjjOuP9qpNXRjtgBz91y64IjVxpKbFIuk/nD6A02/
vka1q1t8hPISP+/8Lm69jotn6gwAaJ/lpIbc64hzfYWv1TTWTgFNP1bzNehtIsFViTtY4m7mLzgA
2DlgL15IMvdvRMRWxf/X4iclik3XHoHcROcEmD2p+wWlb6NRvmaivYgmG0CYG6/+kH7m2978KWnE
MbIyoxF+01n9ygJypEkwSBsGeJm1DnAoyM9cJk/aRg8bW5VGKJXfDaniapw941QmlyEnBUsEJfCk
W0PdN+Fmj5l91X5wSqcUQIR+mYrwNhlulHQ6vAxn56K7RbAJUtHqvyYIlEmpalsOZPVt8cGYJzsK
xfF+qf6IhHozT++rDeKfCv/8wrSkdehFkMZBbLNLQ57Ze5pfHtcv9vsp2KfJA1yRyk35fy/Hd9EU
O+5TKk+KXGNA8WWVLFMPe8IBUkuErXxYGieWkxg2P2xVHlASNclzgE0Z3STpG7Z4xBtjB0Hys6Jt
TjhNiKz01+5kt/rQ5KLhpQ2jBjT7Pcfch5fGQ/l2B+Mp5lFHXvdbC1UfxJteIK9YD91/+dBDjDa1
+iL/G9Ccu/DMw/r9rrHAuptNT77mtkZ6L93QJE0R5l/3WD4Cet/TcxyqtG5uChxGaDmVNcZp0XUu
00o/8ionbUlyxrO732PsACGo52FJzONq+0vlrng2FTBwmGJbzS6n0ZABChnI323zIcCvA1ao7h6w
gXduta7IN1d6Dt/7ibZDnE69j6efm6HJR0o8nb/zLtdejN2YkNheVf51ymztH/SIxui87NI+2JyU
rk7dRblANAw0tmqXchMj02k9apTM67Db98UqZ8JepFr3EABC6GOaZOJ7s5sWf9XeErSL6KMuJJxx
g2gxpgnaR1H9briUkLuhd2b8RLRsLInK9mtZA5c4KqyKznLgXq3PXjWM3GIA8IP0+qBpFAF+f1Ou
nMhhQ8xZLzd4XKvi54DJ9RpoU2GGHKfSZRxLB8NsPn7kifB4yy8cVskKbxlTu3PVWRlBbIQtTmtE
mcUHOGD8qthsa/IRSxXsuclsrEFspave9yX7wbQbCfQt3R5vrIPj6OB+nMclxPcSCFZwfI/IPiY2
Ni70mUoz7xHUxka9Pd9Mnx19deXhWOH3GCWNUzOklXOjib4YvKFgFbgAXZGmkiVS8t0rhujDFm8S
99bYp3gscp5Mgfegmf7bzRoAxqF1kAA7hKXCflQEZ68VQeiRJtJ+KServDq7Z3PWjoSACqx35TzO
8VtqBrPSbi9ROIn3ixftOd5IHF27yBAi5PtWg5T6bzVVIiCsYDOKdyAbxI7Dc9m2w/EmTM25Ph+K
b1GJrl/LdPouS2tmuT+i0ik83dC+vNypniDUXfqTYcjUVa1PpDW4WHKSG5JPRc3jAvFmBdX9cb05
MYl4VO6Lr2ZtiKSlvg6fDQg7x6SvRXPZ/o8VaQ7/1U4J2Mc2U4ENKjiA0t9qwE38Ljpo2SeAIlQh
lbzY6L18+Al5yfOuTDmPiy45z/OdrwkI4EYpeUJu3rSByyFydGpx63gKhzXRjeLXR04yUSTDtvYs
Uc2I+9TswWPT9H6DVS+TTD1NXQoi557UryMMm25L07aOkWNNTx4JeA1UirjQXPc0+kQS0kb6H4js
5IVycquFBquOnJgw4fjeLhi5/dSLdxmGxIgRqDjCF3q+SibemtPlNeuyuSZNGlie6jeN0HXmd0a5
SXioUQfyr9UyRjag0hNvWN89slxccygxo3d/d4B6eSR+HtIUGZpXHOfV3uSMlXlRYxYb9Vx/EoBI
s9HvNi0mWXBd2o4zKIcOmxfwYSSC2oBZYNIkJdGQeYPMJEN0/8FLmlODiG1xljnTLm1LUAMzJA8k
lVYoRNxuRe+90mPZLEx40kx22qb4PUso9/jRz0+9RVztwgW5UyyWiXSYdfwf/UZdSPey3z4jwKcN
C4f+fp26++uCo45nZh7RiA7E2sWPLdjLi+jGw1kLfM0U/EC2IhMdALvGnVXrGgXAOzUkxzSUW01R
mD4pMt8ZP8/ykwgeTJJ3cqBNcrWMgMoRp3qc62bIZoIzPpyon829FZlCq2zu/d03NW3nWp/Yan0I
0HuAv1MBMmGEhnxMjRZJPP12XDoLxOBrX9F/WnuLQuuGX+aLNs1dmoQuVKhkXPIZb62KkY++l+cq
hy8diybuKriGI7wyDPAdVsx8omJ8SlR+na+J8gobhfGFNLuzx48CoxBiSDz2x05+Bg3yNOz3k4G9
0qxIFu27SkV5akuhGWjSLnTeRDE5Rr0gdShDctvo/btZn5ObyzLaHsTUItjHWKyno2uvrbf+56wc
djCBSA8Eljdlf+tresMJjK8Fm28caiDdKoHgb3faRv+hx8M426pBMsGpkW2zAta7oPRJZjsmCIU+
m0FESJoSlPj537GK4YXI899VtM0++NYRSjEIhQO0wl9EHlejURujpepwehss1L53L4nNqdaOVXa7
HzbOtYwt/4UsvyevJjjuVwpwdbLt1aTa7GoC0SqzmjlU9onW39g1ic4kL+CxFelZDo+w5dFVfw7i
AL0BIcsiJv2nGlWokwH7/9PZnC6SQihC2I9eZzhgywg2LjE6+dYKUokxxrsVVvOg8VhnPxdvDjdO
OvCmZAzoHMGPLl835N+Vipsl42z+PxcJnjwDCn9+zpw9BHEkrmUxIcevuS85RG7Ut/9G+GTswk7c
kjGn2/pTlTYK6LP0iACwbssACG+KNUA47MdpyCdIJ+TW7J5HU94cdWlZkDsUsR7RiqcOz4mkmnaW
Jc/MSE1Ly6lvwyNCBv/JchpXi6uL/kN5jY5zcN6pIrVH5wtqNfnu2UnMpxFzokibnAiQ+IPzTQHh
7wm7Kypg9QeOOwaRtAx6B0SbmY/4fQudbx5+Q1W8MjSKVPs0KD2sbzj2Se+Z+EM2CwiBO5fSiDxo
qrhY4F8EKDmiUwhz59g0/VD0XZZjyXk2ndlJS5juRu1KLkmciZcPQqi3spi5DoXZiWioQYixCcSE
j/tGv9HWK9veX5OqCZzgMUo+MctWBg4rOhTiXR7STlKdzlTYUCcRaR+qQGBHwuJeWcJ1mXTbsCl0
62DBVL3POaC2ym5ofUSNNwP42+4dkv3NavblMD/JiNerGqJ4fyP3u+fLUte50Pt5NDNdOjH/T7Lt
z15dWDE9Fs3Eem1rbAKmbdFybdUtabU8JIdgwasPEJ8iH7ZBYLNEzDb8WSHbiUmr+MPry9BBcKz5
0viMNcDpl6pWRec7IRy5PPwx7B8KdNPto/Q6JiUxYWWkkhl8QqejkG404TCXtqLAMGm4M073VS8N
o4PZyKPxd0NvfBciYruyyvXMYTw9xvyaMMeKGQzjuzSMHdfllyoJYEWg5lACZ/mtwa8m2zaIv2pz
PUCtFvfVIq6WKgyq/WJ+csr0/MP/tB9Dalcy78e8KonG6nB0hdjo4BTZIEVDU3+sWgwsNZH2MG7V
OGOB6wEZqrr/X7+VhsV8/Cmj83JUP1ySw4/VjIbZjx1Z1dJns5hLYpDLy+wsXY21Uunpro+B6qru
kdvIH7e6upAL70bEzNrOEuHjHZMUKP/UchJKNgHqSmLZXqiDoiMm2tLFSfM04NRZw4gBLC2wnRdr
nmgdIBQHpkJpBTQApS19zpDlLakvy9kBPOPAd+UwS3m3M/aOV0z9k+2fTSbF4txPMDPbFgObZCfs
LI0/fgPE7Pd+e+6vsLbqKvZX49ViyC4ze1ocqoGCRRPfdupA4gD/bL1PS5BYOdO1OqmjMW+9slUx
dOnZmFAk4DJXBFuMURA/XbGk7KuHCZXPCPDY+DUD5lmSKpqqq4cT5zLfWTJzitgKGj1/b4Iy86K/
gxE3G26BVKLCa4rVwNPEjfkfV1w760bWDingLldSCB+K4PNe8EhLz/kT0Nzx/3EP6s10cMQZLSuv
n2J8l9UKpryexYJSLSY249qMaiE0h2AQrydRe3gK05kWa1+cRtZZwIDti1sK2fBPHWf5E93u5f3T
eQzDWNcamEcHEZOyQcLnu+tFLZVKypQucYe3yxNBQiUaC9yf4akAqUo0eiczDweztrk6FgY0nMcx
6hf1jt8ewQVoN24MfIwfbxkkIuWSCM3WuyMfzUC+mj4SosOSFL3K6LNkFi+l/NoffE8c6qWijhP7
0A1NJZ9528p1WPc4fYBCOw4R0WeDRuKJWYPeJUGpTpWAHbxp7Li/1CTIz3ndbFgBTZSmO/4EUmky
4tsOZxfuYWQAkAe0JWmRffPtfqi47aoYJP3nl55eurTWXtM2gm81K9OBZv4CBwkoFaYxoLTL9P7H
HB6HunOuZ/eLFH0NQq51YIFk8BhI4FAI9m/KTeHaBiIfN3kceu5mRqkXS8dXpOmh8K2MzHO3pyiT
iT3ThefH49DbruTv1FYQiEtFLoqcUclJ/gwmuyeJrsoOb7zyg9uqzJPq1XfvOvEOT67sb3IulLRA
0c7KLX4UXbrlBeEdrIzV7cNTReL8P5JA8vbmns5va8OjrOSHvRVZBMwwhzv++2qCMdsDorxoFLpH
se54BWMEIHXA5HiqQMyAQ61Q/FKHxRc1Be0C01ViOVRzY/nyU5ElZnuNGKifCFctScpjYjyfPzN8
EnNlpF/h8H2UeQSRZHhYpsWrzNrjAxgRwTafKoxFTWkDliQodP0fK1hsC6Mg8cQPz6P4/Hz1xmkq
kzBfYP0mLtwrEpIO8TTZl4zYjxnUSGqgX7XRjX8ZAOmeqREVClu6c2DECh4GPVZ4Wwg+8vMilUNc
Vs3YLt8AhNRGMTaI2ay6Sl6Hmv4iNdriB5Py054AE9sfwLKSOJ2IkO2H2pvhtO18M/YG9eo0KIe4
UY0uH3FPkmv1h9XIgm7fPKNL2ezlGcuH35icgc1DGGwcJ/Jda9dDEE7axkbKD0a8XujlqHC1+KO8
b3G+g/EryypAPnVnc5282LtKO9XrLhk8Hmn6w/c5JLXa7651WEot81RzSBqjiFAQ2OxxwNzCnokR
hc8/vE+HNcjioM09fL/WLB7KbYRZYodTtvN8ssFMXpFyrK7MvzZYNFv5AW/LI1cCkFAiFOOaemsQ
fzsFc4ayLA2T9hQDfWIItQl4CJkWlF1xk2vo9SDWseszu5X6CRPsOqNaD8fD0233wBrIF/BOhGKi
DX9bnO32MLWe05m41M/k4RRfAkm/AkdTgmwj/hNxnq/QhUTJaxORhH7UqKkAf8olh181Ul2Bn3BK
y7JQBQYe3IQ0eFNerEhkquproJ8oAEQQvtEfHOYMQVGnUuHQVX1Xn2TQZefqVl85zeGm1+qKLO6e
iGDzk1Pd7bHFyE1iDvMpiuWr0yL7CWk+g6x8AlDx/uEP5gef5BkzxHef0q0xPifuSyozZHk39hUw
RPsmewpxgxFTfX8ClHWN5lpdsw5WdpYr7d3GWfxO2BbsxXSYI5Tco7W7VsO3EvkcMKUNyCXAqKWC
t1XcE7CQZbd1OQGuvskI4UbpRfrcFaQPisfWiXnlfwKnADYuFF1TWnK9cEhRrbYsM1fArH6wc7zi
vkwEpW945Gpoi+sdNEEO0o8hhJKVHKzE9Kj8o7wyAuTdpDH2eFs1fQiJY0zaGB6RLMIJ4b0nw5pq
PjdOCkA3opT30SCfIu9QpGO4hW1L6IocmlhfJIGRN9ESepS5f4hKLNc5N0LICVKG9n794nEKZgDb
RwuNNLFhSrSNUwQ4LSa8hj2FlrKP1OHBH2egGTdlH5k1qYJJ0M0jtOQi3+a93ONgskxKEY63qvjb
VM1NdXsO7ZetD8K1dbGOXK4A8rJ0D066VObUgoJhZlUxnvudiOf1FMcGMSyzfilVoPsIkii4kb1l
Rc2/bt9UTdvpyQkSiQY5Kc53i/Tw9KscYVtM+Sz2gyIhqXT+V35/Nc2Z+/FCPomoht0eycKBIITm
2xF6B4OL+MoZS+oRh9GZu3yrIWfP2cce3VGYY0tT/KO0ciSPyz5JrX3QPhvBCz+9YlMspBvWORdC
vBowciNy4d4+OwB71zZYiVqhXaxGOxcjSRGQAwEsFmh6ddXEPOu3hTeX0fruSA4mDAps0Qm23rCs
P4EouVGg3Jrn7hnDjUOia9c1npGG41OkRElGQK1nALJ5zUOlPQoNUKkwCk7LC18Gg39SzXz0mpvZ
sOs//b9VdnS/HJP8RQY7iSwYz0PC5fJx0pO9QeHGMhBuK+Mbbf5PKfYbNQGZW8YnxIGK8jVEaBup
Q5tBKnI00+83sAn0YIjosjWRTSiE5L2MFsyP8jucTVJ5sn9vHVMxVvUlLUm9HKseRxlUcldirv9/
WaMcwp43lwF7GuQi44D5BDO2z06oDeel3GmaZ5Du6+4nOlJDyiCz3nXmqnP24CCpHdJ+8sRthDFF
ZbsQ/QUK4hcjuA9+rv7+L6Zon1vSBRssZt22+muQCKai7aCvWxMprLocwZ8gKeR2WW9ozebL+aND
oTGhh2GN+cEHeEwUcPwIlVcne++Ngso4QElHi3G3XDt70ExsxJ2vancJhOAu32K4R7RQLngRr2fR
MlBEls/+cO3xOJqihEi9xE9+W1JiX7/WeAjVFJK9tcu4M8QBkCvb9MJ27sH+SuXqszWvpz4ITOdP
vsKRsm5MTnsr3ACh9qyicVZALVtSNQGyILDus0qNpCfNHVPZfnSxzgXCeKgc9i1jBrANefU2fq+M
nIZr2e+RtLxzUzzDcMxcPhxtxhHuyG4a+yOZ1OABJ1bOY233gY9rUcvRUxYqh8lYZ87BTUGbT83m
Q5ce6/WuSwwGeSJP5eaWPYxmKH1g1C5XsVc3rag5E4iTpdqjgFk2TkBuZXc/8ZCyNaZRJaRHQBWI
v/Q6L7L8WpQhY24dvKRLwarnx23+mO1iP5G1+3TSP28GQ1ubdRwqlei5RwB4imWYtPOfJ2VqJh1o
1YCFs2Pu0Izyi5a7DAH77gnF7ifMQ1MGzktHDH2Unut+24XEvHXoLZamh9LYItH80x7aMS1xUxkj
fDR7n7vxHv32RrUd0jdEcvQycqmVIqlgEbxDq6O1y+ttm/vNAf2MbjqFolne+omvmQsHy2/rsi+/
bomVzu6G9mm0uQMOQIP7pZz8b5EKscZ7Y6qk6sq79szWGO9htGAmAMECGcW0+sGN3g4W58E85KHU
yFenYoUY+c/GpArxji5t1LYUJcx0VeTMDAwHdHbbXECHPAwst6VzUd3nRp8YfuBuGvfqtZzvvcTX
qk2I2O54WN4KvwMcZLsfY670z91NU/aTaUtthbqNLk10y/CGpqchwWRdzzA5pTsaZu997dXtRvQY
Z3+ZrABT9MWETZK2Lvz0DxIQKvULIQuMWCQPZTyCrXvC5lPeVIz1PPuwhYt/INMpSWJrx6AnSNV4
PDwlXg4WfbcbS3l2m78FeQpy6vqIlmSsgG7ImYsIsKE4CW9IGa2jlQfACKI3oY3gvX1h4oJLJKoG
QTOH8Dd/89J+2CXCCDBF5r8iix+czBWXefYrLrc650uupgUwu4EjyJ4gsBhJ1T/f+/HWUldC5IwZ
QSHWECSR/MQHOSaKo6ABqYB+Yvxiu07nIpYk7FmwMhfjGSlIsyL/HXwdhe9K8mI5DVDx/UOrvgLw
pEN5b33xjYm7frAO5kOnjmCkA+Es5nHIpAXk/LeSG5SrhL1j5BVObFcHsbXdZSu6aCWAp8UFyYsv
pFAswdM4y5V5vlkVetQ36bVmH8MrwQjO1LbGTryd+GdVvXHs/WcdxH8SEZG53GgO1L7AYoljQ8/x
rtF8D5LuETDea5ZvjPUcvPdNbuy0l/ibQMJYsY8KnyORnV0jMYctQfLc6GU0fArRID8XRC7TNvC+
OHIz4itLM2HNhCS1sST1X2jMV8C643PzQsvsuhW81ozR/xEb6/4hLAHlVhjc6PNMk8XrgPk89qxl
ImWcJ3TbUw0FjwN4Unj0DTX7SxXxbsedENjyBC3SvvhyjUzqPS1OpZACdtUiYS3lYmjoQ5cYfzPj
H+zEobwDGTgDu8WBNFWk4WAK7+SSsdMNiOhB1baY4R550Ssp0S4M5yc2yw0kCF1G3I+9njLfjm1/
1N4HN0bZTqSPWhLjC1o90e21h9ZbJh1Qj7a1qL3hIt5L8ca3NMPJbdYM67ncCYButru71bb/CsDJ
QmVoW5UmV48cLMgMb+/mHHk7IY+aWloviebugXhwEL8U/80SU9AYtW+5UGLaPBlbWIntQOKWJKC8
MaiPKGX2M+V3R6QI4D8LEN+aeCsHhwfr8JYsoWXlOtRoxVSDhReAff4KuuXzge+Zs0Xsnt7Ap6Jd
t+nS6a18c3ndCtm4DmXhA6WDcO5Q8WaNV5jAT39GfK5CY63scOpcph83yjdOKqIPSHqcDqGr+9B5
JGGQE30eQ5j3+n4kS8XfGbT1R0f+sUHi1tzLeTKH0swqgCtMbdLW97ihcqRkBo2IrhMiPXA6MKmX
jhahU1lK2D6rP5ltk2iVmLGy0u5LzzI+63mGCeOIMOVmoRAc5bOfg5V2DrW0g2UzbFkjiH9qONnd
fYEfHREwfYySuLZvqdUOs5UkLAhSV5f6AoIjuHyBzI5UqspY/en52QprvAFfcw8dALtZ13HazyxT
90LL8cTwxVvsSZRTcj3uULDnzbzEHt9fw5NFcEjcwc/BsZas7+K/2EyZZqUCYnjETfN0nFUF+DKS
8VNAK7KluPjv0DcAUwfVP9/E36F4X0x7WfbXrWFTjHPNSd0NsNcpUsdcdKSAB5Jl4dmrxyTm6lPU
ozrHKbF2A3arxYh+gWJBQuh4QTtb3c3qWFBztbEpaYCMUSh/TUi7wlZndlzsa+Nb5/tBASxXp5dQ
gvaiuGvNoM30nxdkEHPn987ulycNlKY8K+/t1xwEJIjw1N7jtWAhrtK8WF4wPtlw3lXOvnPZi9Eu
viZhPvfhQSTYXIMmRmxXpvGViyqOxt/2t9i/xvRNrFRruvF+lzwc6WeF6sP/PGdeQ0WOmGjG5fi1
ieam73dGSONFFQ00FBtb6WqbRopmyvpT2Id3xtdjwsOTQfsarNIAiA9nHuJuuL0hHUcAfcka3xsB
yEl0AUTz4oyWJP/f7v8BjzyKvMOFXgtX5x3HCAfxk+fv3tfy0d8T377xwUMuATfPphzOtgXtXSmW
r5RiSzO9m0CN4LlLi71nT6RJvimw9xyO4Kj5ENQHjotUEkbNdyC3H0jtWPWZDda7NY8dWoLojJAT
nIZUoyNvSKbJN9CwB8l2DhAb3AufXNfAGkQJpUhKOwEMyTT4aEiqZKz9V56pzE714ucxaaar9mzx
PFLFlRZBLCLrxaWmagxlbzB9eNzEHPyEvxWQuW8pdAprSKzaBlrrwq2PPWqwSEel2r5w6T+4d9jv
yRVVM6nlz4aPIdOUaLugPCcHBOppTh4nAVZ31Y4cTDvKNX9Ois9AVjC5YqCf7vm0PNqli0Oyo/yY
o8s5PuTDszDYTgS1l2+5/O8vXHfSqPhRlN6/fK0KwqbeGaeh8KpGK17Rs2bn/QIzuTqcqxyCFn4I
dscQ+7n8mDNIXbkk4IyR+1xwV0mfRvSWU6o1VQ8dTHFvMHob8wIto/ame4X+SpGRXH4oJZIvk3X4
tnJWTsDnUppJO+eL2idLX2z9h4+muI2L63NrEHFrfEONdZSh3QVJEpgLlJaAlEV6TzUyabHYh41/
6akWeAHkXZIBZEmpdXEwMuaGLHUE/3xjFQbkjYxbZMA71EPWZOdYDuaeKWkGINVpQPVpV80FKPdI
fozkCqI1M85Y7dUBJvI+Rw4JuCIkmqZ9DW4aBy8xZjXbmciZqRP2jLJI9MxcoVaqlkpaFovTDayL
aLrpT26JINFepEJduZXk/+Rat1Dn+w7xg0k8kvwq4Z6Y5a5BRYxV1ewX3TVTdGKIW3PLsBtDrA4q
Y2jTbwq5ERltTeDkVuQgKsIp9zZPNnNMx/qdiqf9Ux2m6ZQEbozC/ZnNOdJ4YQpwWJ2HHCSYkpWu
NV+UJP5Jb3IgOEClk6pBamtOKZQan7yF5I8gnmN5Y8kyLh2WKEnT+ZeMG5O+cunN/DXx9Y7xFB9/
BypWo3h/JRSHmIpmSE6o0m9CNCJQpecSlbm8TB9z9OSGcFyx/uZcKj/5VGDqrcMcxUp8lyIMrSck
JCFMPPJhN0T+bug9HIVGEI6+bOdD1suwe6HqROzIV/Ai0LFhjnSDAcM0X9uMNvfge/vmlWtJuICx
StxANURQg2RSZKzn32EPbDz+jfqsE6OaRcMalOYPvPSDN/xV70zAXqcqhRIYpQ3sVovtv4JyNyiR
Bxs+REH42yx/6vuJRJZ/VF1XA9ABBIA/eyWiOI7bHsHlyvV5MIXX0AdKK+K0a3NYv+hUHwKwsB+r
EBs02m5Uk+QTzLJ/EsYBHK4PFwNX1aL8ZhsvGVgoraxIPS4xfMZp2rBGBse8Eyaf2nczY7Snji6j
k6+xcI9oN1QX+p285KVr2yXiAN5cXHkkKWhBjy6tI5jnQaU/zmvRtrM+0Frfi01nLG+DxXU8eVvp
f1V3yxNqZXlsxlMnLjdX4U/OEAmfQCdY2KUZeFs9JqXkZKlCNqz446SMg9/mPcyMSROH1iVdD55Y
cZt7fF8/8m5igP2drZgsKgXFqlwBj5Fxnskg/8vPb3E3LEUUZhvaCuYmEs/CHT/JoeFzMHfZvtjX
qbm33GzOwiarwZa5sViL5kxlWC/ltBoO9tCtWyF4FB4o+bhr5vBnTX7H2Kt+TPjV8l/ZiUSCWtMf
pQQ1tVtZej9PbELxYwtJ6eVF5is9f6cy1AbgVb9m07aydrOeYG/kjy7cq04YDXVAbeucZQY4qKo9
lIcEhqZAq4f+uyg3Oej2IM7f2QzncYxkJ5SYTI1p36O/iAPqcFzVqSyOsXkKP/FGCWGnN7mxlUae
zxV6XEtVqSiFteP7Mcd8+KWP1KEHbMdM1FfWwMXEufZGHtcXu4zLpM1euKKBS9nYXHEqz7eOHXa1
7cA6z4gfmZOwjOfhBLYyHTavEdh0EykZPiDm2n+ctZrj+jbvVRM6t/ijN4HQg4hMWqeuIa6itAD6
cO4Hi4GdGW/aURwRNZRwKfyb9cyNlu+P8jbswC5qTsIKH/kddT4o7qDL4ocaR+PijYdVrWc/Nr+V
/cyGlVTyqaU6pkeTKg/yn9BUag7zyF5JF9n8jkMEN4rF2UOSl5l+zFEHrqbLFacfDH4q2ZjC/f9/
jRD667inZzyowRGkDGr9UJcN+OlnYObwcy0EbNCz1+wQEy9yAL1Inqe3w69lyD18A4gdG2HkuR6Q
cok35l+0iK/73Ev6kMJ/31tUxnoTOCGQuiUU+gXyFDrmlPEjLU69OCs5NABgm/m3igwr3iMCsCXr
U+EPTkM2XAfaNXIX46kyQ8akFeHRNCoSl24y/qL5GPVkIkhi34JOp2p25sALZr9zIvD6ciE/ESKd
v1jrV6ElRmpWHqYvQGDebMUyefuw3zF3SiNxjc8BI/mRjVQsgkvoct27by/EP4QsUbAwdhURt7v/
C2wM02SIbVr/bRG+Gc7S2OPHfGBvELyw5vw0MpwVsEAWgtpe6BWGsYB2PSEogyLs+pT9+4ZZh4X9
qUyrdwioGSPIGIDEd59Ms1jSaTZb16sFO5tlZp3JGpyLzlwjDB26b15qK6CLOk6NYeyUT9ptPv6u
/z3U9l1hZKwCBAd1d2VuAlWvz2vEeTe2Nin4Fn0Dt/84CP4Bn6ZqFb/sbbbSahUoc9/mrlRWYjqG
8fPgIfqDdDwliLky9UIHSr+FUuVhiZEIeuu3UmOqpgX84WkPjmSwvhcSoeF0KDhcF3aZGOzT9l7Z
XmYjA1aTQHBgt/aJ9bZtYFq4OJjHhNG3/BnJ3Mcwqqdu74VtmktSq9CfmEwTxm637vxeWRErcbsa
zc04q7SM+I2d4VAv+zqi/Svsth3uWxmAFigyfQpyoyO467N3T1ZdSGhk7QW/RhAjpiL9LTR/Tymw
o4rLtXjH0G0MgkfZlzsmygy7AyfQoMSInoK2uqEXLJ+atMXZ/66C3g6IS49KV5KBAMVDHB+bJ3+G
rnyGVLqLUg57TqYcHGDBltchvn5sXvIAxM12oCxzVd42sPa1fjkFWLY6wQ5lXXg6mx28hnBp46WT
PsEuj9ri+kFS3omAp3UFyCoX+tdDO7ljN5DCYc6/CXTTd3izee1bAIDcz/IA46P0Mgi0e2tEokWW
LIETZdmhgOHS/DyfO5OzuBZdJgwMnkPNR+504ij7LopGb5wbI5f8i8I6MgpwdtRlfzTaPgFTjYZa
+HFnBk8ow+dENhPnhi61KRmpXjOD1RI3Mpu/jlgFTA5YPpzXwAsIKUKofnRM2y8L7vRgycKq+KMo
AVDwGL9O6WCqHd9IxXqM8W9DE8jerJd8oNE/T4JXQ1m2waROGiezkLK2JwUYFVZw4Ch/rJmhUU5Z
+/tXKv23TMkVZN7JHzD94kopJqAMKVjaMyIG3ZBYFsBBC2g2Pas0E/FdfXkImJca/sb0h/S1MB+K
7dCt+XbpSzArsz+R4beKJji840xC6euFzFdx2AjWHJIlcAq/jNVEaO6GradwmDbKFmJOtrZuQirl
tCc9cQP7R3DjxLZww39d6nnv/i3gKL8U9afXF+NYXdonTxjoU7yPZrJBCf7GDFc+sOyBPh+Dpy3w
aiYu5mJ06rCGVIIZrYMZvPjCil2u/YpriaD28dGoVrQDNlJEAo7BiyZ4y0SkFtk+U/woxIDmzc2F
HhgskShooPWraZEZ5/7iitsBDM8XPpZJdJExijOjnukRJlsot+3MnLDyIRcvyqBQKScqFy1jJ2gp
FjLeVd3rJ1WEkCZnnXx6/AKGIgR560ypvbEHGBVxR/Pxi5AKt3dxmyESYfUWndQVxlTVjSzTKe9J
A5kxC1GZQ3u63hGO5Qtpc6TzbKAZQYaWyY9JMH3pax3WD/3RxxVEvAbienY64A+ej9wZAYxIA6H/
Tw5u1JnzvyvuTITrmWU1va6maxABudtRz7ANGB01nhmA1gxwZ+FgVJyhFgOZb0lthmjVQ7aIT4jb
v1uo18xcHAz/VLWGu4/Pk0t8DCfIjFiBza+NIDYrtsWwZDcCwAzIR+C/IpJBXYiOAIlU0XiQzIPN
hDfRON5nPSHqCnp5GxYQvgAnxID8A1h0vS/Ud4t3laJA/nZXDUaV1Aoph4uogt70HMQ2usw7mPvo
5+cd6giJeOzisbJn5jG/akX9ygQikgsCd6kSESpMrsZMu+uNTs6OF2eP4kpVD975eiBQUpkY0KEE
40K27ypthOYymkMdSq+k9WDpQ0m3ajWpkFj+vVtZ/R7YcAQ1IkYeOluivI221UyqZEZvFXNsqY0T
z7dFaHaI27YCorlfwAoBuLO+p3C17qPYeWNepTyf/qsH0FOymg8KJSs3H3pA1oqPapwlis93XFCM
aH8O6j7eaDPe6TualJkQawA1CZPfr0V99U5SQilqMJ/fnLPrH1LSz+t+s/f27YMi7BXa5J7DBkaJ
C8ZoXl6McG4N7CRpdeB/fBxhRkOyxsa7xaytKmkXe3vDVOxmjHnoEc+O7ts1SD8r1I90KAhZ6ihE
r+YVN/lnfSAl9VYTfbbvl02MfHNZMLFCLBM5sy2lQU/Pi5xdnx95mQdeNeXqA2hY/stCNFB2dy/g
y8RCRRSR6BfwcfL+VzrMImS9konYvlIRSbV66HtkxriEzztAB4tWLVac+CFPY3dgmY0AfZvmvpS9
t/tKvv1tCPfotHh4Gx7SVT9why6hEca3g6evNcEYRMaOldjXWlJqD24Pb7LqdJKs8KRnUA1P/Z+x
r8L0LbWcSq2pVvT8sQSM3A5ld+200Rc+owteCZd3cczqae0UGGQVFaEkjcYYHIc61yXdLu7sExsq
xYlZIRWqIpiZJHAUJt8pXf/xI8wM1JSE4ZOYj2PoFvVBQQIBDkrlaPHF1ldV7VxcjQNAvxNZUNqH
pi3dJz1Sn74ySV0ypil52YzfJOJIHcnL31dyCW0UDIaGwKDHdWpovPdZVLBoQT7qZQb4gWCZBA5X
0hPXKZ0ChAvtryQIUnYhL+JEju5irNHhecK/mz8TwGhTMk9pyxXNqJDuQY1Tc2TrUS7UHwH34Rzk
jxBCd4/nKKpkNn7RDIXI82UhHoSHjTB0w9GzmdWoPiAb0EG1M2DNDVQ+c0TDssTsRdq6aYt5nu9J
yxz4WIn+T65K9cPUOm0n9xKfgav/3psi+FJoycwk8D1x7oEgtyUpmCpzqXsUPfbkFf72b2WP4VUF
Oe4weRt+nfjLe/nP1wnmEa4PsK+EQ+vdMYKZt4y5oxaqICsHbDcCz1dNu6HLY1i9l+VpB7Aem3qO
aQQNp+GcTpSApclQ/fGSAkG3+IVUcTImLpaNkKr+JasAdYvvXsim0QIJYq5Rn9K0cr4wv+PND3UF
JgymRNiEUKPEtZKoMKw171P9qxwKj6DYSO6xcJiaUCFH8qtTv7qeRSK74rkPWu7fMWY86RmASXt/
9T4U24FiRBlldU/wz5C9/pIshd+4IYZfref2RaOrYqp5wspTt6h96cX2MQAQhUbnih6nXywnb9BV
QXqJql+H9CA7cY+wu+bYdbBKgg5lzu9IqjkFGIoWAANhcukuRg1qNpmdpvAuZEasAkVRbEuOSiZu
sgqCLnnMDwdCnKXI9m9OMGoZC7bUoa2Ppdf6aHHGVxEplSVT3NAyNONMO0UZb3hy7yAY5WHhWV3M
aPl/GeIeNh+mQYLn6OmT2vhUbggg/sjgS43RhiQ6Avzi8Ft30s7h10WR9zddPRbH/wJ3jdSKAO1u
3VAQbV9JIKTsCV68ri+xttGyebdU19mI9d7GxO6vlkZSgRAFk/S+i//yL21xuQJjxJsIPpaISzDs
wKQunN0Pm29kKHqNuLKEs5b0mWPH+l3L/gLUwCQbZ46pka/ZtAQieiyE5sgdoxGom5Xk70sfRTof
DFGUHoouUBDUvyp+yN0WtGouoLBmQuVT+QQyI9rZeKfg2D8NKPp8OlAS8TGknlhgH4/XG1bdz+Bi
T4BUAwfPOyx+1oYnT9ployEt0GNPqlutLrgGJgBPyYa/YstzJJWqkbGTjasj9xyXlJVwo+69LsDl
SoJkUBz1jEhGjlcv/QJ8zW0bk98HygP6z5WOotrPJk45n4BCkKEfPB0PfXFp47V1V/G6mHSvfPLT
515o3dARd4oAzo9U/JupAfdlZF+JCEB3nzKer+HymUHd5BHag17LKmvrlZIKMHY4ObESzQzyvJBU
/wuHOYKuFciJXn4Jw1UdX+phWeXeaNcnLiNUP5HnfM1Xa5C251Ie1gEQnpgHM7s5gG8aMY2Mavck
C1EAKLSRvbeN9fYsg0ki7SQQA8m165qvEE1YmHMnDLiHN46QxOVMDNWEOX54SAi3Qi/NrRIYn/KO
NGOus8CFRFzWHSFVUGkMDQDSlMpg9nQG0CDMZga2SIkEeb0MkYzvyEg8QLlEXgiEJdg72iUI/pq1
KI/hnOZ7T0zNqnjQNkXTHYJX1VAjP/cO+NaPLH4u0yOtX9DW+NykSUBVQVq6NLUGeySlL5mtZv7n
E/6lO0Vos6HdUwtgaDt/JaMQfXS58vbgkd0oYpMke8f+eSefJR7MLLejlRaBj7MMuliQhKEAAkbf
rUq+VYWVU45ij1p84OLj7avp7sU/CundRdz8Pi8IYjC6A9wCFICGbUke4a2G+oCF+vVW9C2jVdyi
6ApOUxYSSO5xXeSq2OYhwWr0OHcKU40VeRn4CSQTTWnKNOP7/uzHEbzXJ5CACDGIp47iYluyhVSa
NsA08LpTm++7HG0E8Fyk0+2j/SuT4uqW9aAb8s7hS/q0yacL1Iv2PKRKROQeWm2/9RuhsMR51da1
zxLsiDtvzMdWuRbwc4gJKu+y8dDX/fgYssfMsPfiDn9oeGm7ZJHA0OyDrjcVBlxspmiAZmLuREi/
PndYZN70hYv5x13H2fWqJ9eOgY76c3M65+acgVPPBDBX+d7Rj7K7nBJMIzSLBJdRzP8QTUTPO86p
3SF3yHLSuJsiDt9A+cVbSEAlGNskAXvbcUwoftPXrsuMiRl+djO45HYEebdhdgKb2GQbRUe22ieL
K+R2mnKBiCxCrkYrhw5DqTul9ZeHzvxn5Dob95xq3tY9MZaNgHZ7i+LFekZDmRVTzFxVOAhbflij
GwWXXWSOLiFTHD15tuOLkHyX6vNfShJpwPttJNQv6F+R9EXSttSG8TtUkgvOonF1jvwl4alIQhrW
qyoEnsfzJeF6b78n3xRCpvqekoD/fJReGgN6lnbewltfUhUYtXAHSrosSFdOWJVfhAq5qXjlLk26
54OvL7hnyQ4g1tXO+ZGj3B2PW8FZoBuEroxqS/ZJ3SO83FNVvxTLfAGi+eoQSpsr60y7JmLblPRP
HSxLSXK+p6E0JVGJAxNEJHGXwWW8OTO8ArMp/kJCmmBj4gRa6PZFwLEdaLCEYoBO54Lfn0sJ25ch
T6XVPMo0BtPKVh8APzgCh+gRgSOkcqcIU9ciY70JrLCSRb5BeYe2q1UrN9zNNPIxEdPRy8b5dgd4
n0lWhoCCgDvSq6V9d6ivQc7r25RbMXrjaiaq3fXlAVXHVLkFBUnXYPo4i3xKIzXtjoNy/5IKhy45
7JzBBCcE+6T2MVwPecVmbxu9oi2ZKVzl5anDkFZT8SES/OondC9VX3+CsbUOjXHvreou40SPA7Vr
2uFwRhwCdBc5kVqzjx7NhKY+J3cWQJlsQqRqHqOMqlD/nEwDB0g2/0Ak0RGrqKCr7bGJcwcLdzDA
JxmBt/qA3RFx/3kY6TKRar6Ov2mOaueVcBwTbMALnMtvk+5+JCqNWqgV+fn5XF7HCO+RKxtVK2aw
intd3FFgb2DJDn7rWM5t8E6iiIOXsMqH3PwTAlLNoAU8u5fskGYYjB5dVzuuoLzRyLD+oQy3BnFm
EArSWo/YNNF1v0sdV61VKrrQb3b2J/WQJLHz9c/Hzky8JO0kw0NGukcIqDV83BfUs00FguuGrcDL
G92+XX5oTzpvZLDr48gxcYr74rO7Gfm9D0sA7XI/IVYtSyefPulRnu7PGqOlGe46+P+3JaJMBx/8
cactFXVwDJtaUNiA6ieUVba8P6oyMvjjByjm+I7fqQU+0BIN1mRiaE9e2hUgqd7xGEGtveEfxs5R
/hNwwes0Y8ftqfWwKHhjBei6Y2PA/BGTfMT6aQajP5eT9jysk76FDfiieNZgMCwsP/Hix8WCXKXg
08GHGbzLc0zGQIPrdbEdNVyVLF/xgjqw9gnTgmdkRSZ17Imnt9w3NJZmrt4k1JCzUwodG50onufn
3wlFIN21v3q/EF3CtFu7SS8KhRHQE8UsmW0oaT5OKx8Jdto97ChiQCsb7n8MLLhnhFo8zlzEmgwn
mBPM8fwOFW8JDPLsL8GHd9n4R3GFihG632fP1SruCD+haIDPIblALnIa6ZsdBxT2wEg+zoSnMVjH
KdXJk3VUa1LRklbQb16qIXp05mT46ZWAI/+uL5Tc6vXMUIJvb71+QfOqeRFH1sZJgJcF3J9rpMOS
RocmA/RHTvl/pQCkLUA7t7ruAvjJXdJ8fW6Y2TkrO5qW9TsU7sRbUhHBxVOecD0Sy5Peo12jLLzp
8/UYClrG9VXFiLQ/Fzy9n56Wpi4PyuBJn0NFKGPSJeEZTNimtqcBu1nhFFr/uGUL/csifMXgg9BI
YrHwXlshOGL/HZHjGTUvPXHGZfAE0c+3vHV4KJzG6Pnr22AF51eCHCLTWE9EU6i/BKTE3YqCxID1
4awkNq0l/KhYNeCd+mEmvrITr7JqonCFZNVsqjRMeWxvsCsC3YnJh+0b4T0JsxpbR8TVhGvJ5C3F
Ssux0+gfSOtM0Hj2bQTfNEHi3tEqDA9rI4CtRkZnUIAOs+dCRCEuQk+1ZSzE6qGaDWoohO3b2g5/
tjpJkKiIHH3xXUi9tcIGZea7FGTnrPDZhb2foFTgMD01wBv9Udu7GzGRoQAUjAdGGQLvVToXDRro
xXM9lYCYRE9WVGNxkCCXvGPNv/M3/Ulu520fTtN4GxNK/J5CyoRHwONtKmVyncZyOgoupDq9wJzi
XhNPeZKFBjXD+z7ud8sHttEGwD4eYq8IxAP2eHIspoYAKZUtdMMcTyRob3x/iSVWfGMV9aRYxjHH
u15bEy5JR9AMZ0g1xy3IqEB89d0UvkNUOFWB9cbd3jszBrv1YD8hiMxp23fJMsJhxdUQBD44/OkP
hJad4iF9YtgG97n0qrNF+VtF9Th/uMiWflRFGo8hTjFav3ai/E6QM2BF0qmaeb/52kSdrPfv8FUW
vke0AaerDniO2V43ScQajRkhrycSTnG254oW9WdpQqktUwDrWoa3u/65Pd7Gt3hhPgQGNIeyfVqm
q2C8G/eTi1F88I6Wzrj2TkERh7ArU85s/o/xOISE14K0HvpaBqovKnwXSoBQPQxGUqn2tmChvQLq
ZykADmzudMbZrvRxl2evqnak1WMm66Cc+l5T4BBuCQrqwp2GBikrRoWAhlkJrCAK+9N/xEw7m+lZ
336u7exlRMysGQ7aQiygJxQrsZ6KCBmsU4tvUlQI/9N5wdxSGqiuj/nsiN6P6udoWZryGsEScUIz
65HC6EfkiP1J+uCmPI6hL6A7ZVEpdtuNPtt5DWI/7cDR4glUFZNO0D7blrJBwt3jiN5WPItEvhjP
28wPx0uJR69vZhsvo/jA9MtfswZfa9gyK3rFnh4rZbHBG99aVm8aBUjes6yOU2PC2rfTa6yJ9Jld
MnAhrpc6tKkj6p08Y1FBCwNhGwYO7fAMdjk26na+6XXkzmWrPHGrZFSVq3ugpg7SAY0pj7Broenw
QRUfj/dBtTGj17rarDdKq3xXnQV5tUaneJt3OtoFyLQc8rdeqeJbegb9Ej7y6aOtCBpmx2z9gUoN
40qreWwHv2p1+QLp2btpcs+WmPvoam16xrWeSfk7GUIjtHGgo+ocFBfi3u6CKWDN4czxKvpKmEG4
mbaM+PhDYEF3qyFL3vSOqvXrR5VZcp1HMg2Vxld2Ch0UBpd/9u7lBDRLpz7mAmpw0Uo3ariMKAz0
xoxttp8I/mnVJKfJ4UmUWaZO+O/eAkMKSHXieumWchRmIeRca8QN0RrC2bVGFkr7pmub5Pg9GPCh
vO4+PNMLpVk4AzkpWFUKUzmjifklpLYQa/nDtbedDiOw5CLCnF2yW20T7MekW1WcRHGHjYOha572
1o3J1+ij1BGZEeg7I0dO30jbxEbNp0W/x69J0tFkVM+jnJ7JgjuQEW57tlJJV/nlQ+wHlxy9DEiY
OmpzocuBIhzDpdJiYHcECx6ZLQAxNsk5h7jXokXkuy4mlCDEa4Y4ReiPYj7vCkujSfzWmC9Fkjy5
HKAcKgS7CLYYMu4Tk7UQWUgXai1mK79n8FXjvGGSYCkmCFIUZdcNhwj8nbdkxOIGpc7T+837XrMs
sBNlF8iSfEpu/WT5WIPwgXWqt8TzZvTAxnUf9exTnPpsTWsqU/mfLmD91diYj6QilZQEygTIQrZi
6wT3rocBzweUiWsU+fxPbRV4lvBcJqHZv4Sqvo6pc567cvcv1FGWFxYB3pvY4AmG9bbf2JoIB1I2
Xh/v0ZPMPeIu3oWQky6cAAYt++16VXprg01ZareSL5M9nUf3X18oJkrp3MczY9uSN1rLs7Ke3xYe
kdZdB18pgzIr6Jbre42E2fFKZ2t2DBRgsa8dmm2fTgNeBlPwCzCwK2eGOKJ6B9U2wJyfND18PWZ4
BVvgkRR5Ee8DFocMeyKQPOhGhcBChq3P3SFgNlFLOzlUlQqzv5ufdSpq+DNfWFLfVnRTuwyvmOVf
mus1+Hx6kIY8IHvohy94W8nZX3Dryenkr1H4AY38/G2Vsnb5EzVjkfsC5XNvrMMjT4CETiGZh12j
yQo2hesJsGKXiMkmcUcWwsSvetSI2XJmlSHGYG+rcKd1iWFdCkNnL98kb95mAMKb/lKdg/KD1Akq
JWNwvTYajPs8IDXkQm5WB2K7IV3n6pkTXbYmyhJUaPj9FZXdAW8aXyYWD0aC/iRfE8i6XoimNkSv
WeMTwkhtFxrLVIghaHtLdu/mdQd4S+gA+IIhZhSfZ+5r9D0XLJ6LpWLYAnBEWUIhYDaz3e3CIaKV
R297RW29AZRugzCqAx5rHIL1MwfWZlokIrp7SW0Me1vlFUELv0iHP937w99JdF9dKBxQ/dHjjZAv
M0vqMH9PnI8qzcnx6ZE9+pcH9qRlHuXAABdhtlGSVyM9zzndg2agbAVFN4T/4+eeWdab62wQCO1k
XNLklP1RwOFNiNdvU+vCnO0vjbxFNNMg9xx23YLrTbRuPR25RmJmE2c/JHQiQ+2hwENLB0MmF1RJ
fPGvu2LVRlE3X4XvJVwTnQy9BCuuqN2D7wbOaYFYmGW3hCdFGsL0UFsH1nBq9ZxkZ1IE0l9rq6ME
5qwo+AlH4MvHUJK5W1bXJdwL5uOUX6wiyHjumcV+Jj5G5M3S3kfoeGtcjaUztIU43oJlzeB5LHjt
lHw0VChv/R9BfxGcMbgewXSSgLOTqpsK6FofDQLsMhWH1dlTMR2UNgdKG/Oz1PuK4JnJCNSXJK7J
XS5Aj9x9AMnudxPCb4icyApM1I331fjEMRvyeXO7odhJPXYTt6QkBwGJAP9Edqv4KPEW3ndDumJn
MT8T1vfOiDX26AwQJgfbG/hwmR2eDQLvMd2BZHIbyFo7H8IoURsHA+5A26raemAxzFHXcojcQMLE
aLkfJQT/bNXrfpL9WI+sXCePP4h+FzVwCzsU8b0VFUwjNu3ZPIvPPdLUNeH+a5XlP1iIlpn5BlXE
ge8zz/gNvhhoSaQbG/zLWBtjQUjd2Ox+h133pEc50H4YngcGdkIYtQodGWudt8W/wPSN5kiZ3QmI
8W11NGaQVndlzFKy5Ezgoac7YL/NpipXuriApeg4fdrkbXeM+Yy5pmYO1Nrxjx5Rz/U4gNhboM51
sH0DWyopFoEFa+yt6N34WdRn4l4l8ZwaNk4CbquQRaL86Bpmt6x5hsBFWtP/o+VuzgkbO+edFe6O
JWm8vxY3VHN83e1MabR1vks54svZvLIhHgXQ5gPaqA7aHZvjsxLdepuibSNuoqKBoDg/jEjEqM6K
slja5EKxf2zaw7JvwYUf8B1kcLMQar3/ieHq18NlcH8j7/VLn+b79uLSl81zRmdvy0hSs4g5sTih
3GWMTRgUTmBLMi5/CagiJ9zPDcw/xSgzoaVZ2U3AsiifMZrzuKYCQgybDiJLD386yJHZKSe46+KF
tYk0lEgR5OLi8D6RdnkupRUXNEHoGeAbiBttAxach9VSlwPfM0SeHJ1jjHyU6wfSnDr1ibVxDHDi
0GWmMTnvB6QyX/F5f6zv3Nw81Aka3kb1VrHFYVCf1GXXBo7v6sZ7rPsukM+BhYBVSx28SenX4fKG
PTr78r/KtQSeJg9W28Tn4XY1h5AmgefKb9YIsxxoTGCLWJgicD+vWkne6JYuDV8kg8/KJ3zs1VyU
qhmrvShf04+t2KsX4sU3+KVXwnaMU2mHXfOLPpprvLxH8oqe6bMSivNPjulELhLS6iBLbHlDe2+S
lzfCdm3ekr7Bj0IIYo/cSBUVwLApzLcGURe+catLc8OgAesMx+TsquFiCGb82FG/+LEtd4lINgQ5
A1gHSTw1P9t8pT2PoowVbiE1mO4f3osbDla31mDluL4WE+LolH0/nugz1M95y3gJr575DI7UtkyM
0X6TBEdtbfc2SFW5W2/EInwQNyWf4+DdiJskBNrcZfODdOBoP18o2dk47BS+tYlGYXC0pwEzAT/9
OOwp2KKQ4yaYwM03zBztjq5ZZLv5LfLnSrXG+P2hC2b7Rz3nWH7xLLIL102WqAvHVRb+GJzxBnd8
jxlDgLlM2FLwv9ZF97Zf7Y2Z1RHfdG6rJ/ex7xUUub2RKfa6yEcQ+WV+iduzXkyT2tEdfuN2mZDY
vWUKpfMsM7iCNc00d5GlG5WfnRsN4+quFDKPh8yLb0wUsmB9p7Uz2xxpmtSrbcA2I7iahiimccNB
Htpi0slYY7qSwBVt+KaS0YtlJFlrDpJSt961hEXXZP7DF8kB0v+nPnEfWAN4jRcWjk5zn9fwscMd
tfOfksLxYFQxgvAS4+b/Nq0AUh0IUvqGc2RUHrVbJALYD52MMF4Y2+jfur3nfDYAutKKilrVgACq
ur5XYqOglRFtPsgJkGvsr0LW/Is6AmxjqJQrisBKE01aBX5XGEt4Vw+mDPZXVKQ1lVqW2mZptBVT
68PMZzECPkDabEgRZfEkrePQ8KJGiv+ofWVe/U4hw1qvGAaGinpobZUoiFvjJJomgoynCNEW4moQ
fJdAVcICqJoabBR0Z2wUR9ZnrQl/2rDD9lfy3/XGyO0COb8gxg6wxu4leuiWqhsMjJGX8gsZXFVW
B8FWHlSPvcx/PKTtfcDEd2k7dBGdUDIkDQdAA8AX1QhTOfwehIaUOvy14z60uXXTYZVKWM+WIz6R
LTLNJxJQv+XO9I8U34rpqqimwIfaRlxDHcT16ts/dvU3LbCPbqztPuxVGm55dkCW37WZawB9oWJd
Twx5ptQhQ2eXYDRRoKH4h1ssgkh7TTyVX3Wm7YCbilOxk61Sm+GVIyhAzCkoU8VArIfubWVwmBcB
A9oYQxsNdvwc4hCrtR6SckDilOO2R9XXXbTMQUeeGFOVNN+GHGqC3vy1/eqDhWECIS3XYUtyqPlR
z6lo58sWeeE+1g2F7KDICN+Q5V1SJj59LTC4jXHBCE1FYoEI5wS5LZBOgJpTf6hyoFwGV2NXnZuF
4Z36P3UfGV1Sk0rUffieX/XTHVJo5bpqAw1wUeuVx3BiB2MKN24rejJPOh+eRiAB11ktCcHhDUhj
QJ7pmPq1qydCZ69WNlPpy2kb1J5svhFmcNDUPEy8D/cvn7I2fakl/sTCGadmveWskYSYmpt4o19p
c3qkski6IGDnopiA5VTRWn8FsNDz5hPMlyd9F6Tq5m5Egq+kIhgZIN3pHciDucMMhjgf4SHL4iCs
TCUQI/ripS1t0Y7vz/gvZ12uUSJY2vD1DGG4NiPFw/qsaswEThs0F7QsXt/Vwhqj8POB6u+38F/+
LpJOTnRE1K+RN8+FzJPWT0BDgRbWSEoXf9zEh65fdwNyrQrNRWUetvyn90sdUrexxlZt9Ov+oKa7
hd3M2fELcY9KpvboQgCfPLsITy6ZsfDUypE1MfzoL1/cO+3aWVYALqO6QkS4tXhy/oU6YjTMttXP
XpXNKm5IQ2LCRwtccv0kOEsgY20Hm+AzvoybzCPjGuOWGiUpSza9Ld6QfQODpO5by0Qi1iAmIXc/
3Du6mVdQaL14D22hOcybIGMwRbWSPkKxPpYw1/HZ/jzz1V47Ax+hBC16GU6fWY3a70MBMaVtYWJk
UYxAWqKuShinu8Mkw1taMmUfmqKz/mtVUWKh1NBT2/QlJF8HTrjCaTY2epCgJM766DgQ4GEG1SUc
8kk9/hcYSOvLHNnnjztgkaV2oLwV+7HsCbhAuor8W3CS9nfk9pQe7nM4p33BEgFKm80T3qq9uhaX
HPVwbqzsqCRdYJbbVeWPMZKDzKv46UMHTMHnGOdFdKcaGtYekB4jwq39cUEWg0784B6ma5QXlspU
837SGi8dhxJHmt3Z1mRbIMwvwdgMSeeII/5AvtwW8/SPBEAooybvCr4NVdcepkR7cTcwX0AHdAPk
bU/S8nQN3qaPZXn2Om6bBlldWW5nLbdniPr/OdlSdMeN1mQ65LPnBTLASIne3QfH7s68HaXRS/th
NIHpNMLZm4o6Z8GU94ikBhGOs6kEZjKbcJhdnFXhrth3uN5whPkVgRQrSDMnR5Kc6U7klw5BVPlj
ewgaj8fhVcF3TaXfdj+wm0HUe6/SUzM2QZ8ynTzhWSjdlkz9a1LdUqPE6kCdsauorbHxpD6VnSvY
uIzFkCZJ5pushChnVcylyznPJHT+aybgC9ZlE/J/bLkYj4FuZGEv5uacMPE8kMRswBmlN2X/0zxN
sJkhFxcS2Vv26BmejJ/HdcEbYsXgWR7UDkdExxEooLOWF/FTxn/JvbawX5UJKcVVPb6GitEslQkD
04aXrnRGxHlICWW4A8ah1cOb3BApRAVZ040aabS3VZb5m9KXSvNdE0yw7HHbtCZGCdMv55YSXfFt
qTGaACXRRJGhv8+InlZ+7FokiCPLg/XIHMz3toVK9i6+BPqGKeRvw5TbZ36XJieSlVgPjCY1q5v9
SDCviOLBHJFieioXilBCj2HQ8eYQ/tqfGVMhH+5WVR+oj+PiFHhC1+EBDs6l6YnV9pTNc7v5NGJu
8kpb14Ff5IuFgaYPc/HLtcbgsB4Xfp+vEVOYLNtnQpqWO9C49gqAXlnfHOCOM3kwgbMIResACJi3
eqykOWewEFGAifPdwbhScuadqQKd/op+KQdP22qEUy5/859TthxRJflV3oDNkI35qOaF4xrdrFch
nJmLQCfJrRcrraNMadHKvW2VZ7VeYqM7iuDFCRYLtMLOc4q8ElZ487U7IFtlCmnkjSQs0yPILupV
tlK5LxZ5JNbTSvWWMVxhGxhbnExdYwN33ayVwCLgK97DGUl1zAQBTn0jSzVlHQKm7k/ahnsmry4r
xTk0nwUjhN2UQlaP9LogZ7m4huwKes284m3SYCCqfK0OK/gu987Sig4XOZWucwgR42DSx5RY2i1A
TuNv/QK5BbsJcIRz87EwHaK9Ilb/f1outnDbPnN+tpBuSjKO3lT7iUVFXDZNL2Akeb2dP+/OVgJ0
U6uaFWuIeh1mN0e5oBM+qaqNt4iCH36Vp3LfhLF3ixraS9WyII7usmPr04A0V+yxI12rkGnOChPT
XDk9zYihBrrcbvjDjlFQ7kPU1w/LY1llz3r8l7kCqmteq+KQN+ctBVpLPlIt9qKyff3Fc5I6DTK1
kQFPb45u9HmsmgeNqyCWuZ6bQUviC/2BX3Rt1CtJfJAyox8V89RV1mHZH+GkPEvN35u7tzLwUYDO
qJfwqjIQNxjhq/uSKB4xy+SYoOk4CVA1HaV8YP50kRUzLInJa2qWI3+pOePLsz9Tfofh0cRIX4Ul
yi5G9QaxGNf8eeDoGWAg5FJQSEYR7ncd9b6q74CBB6FKWZZPXwSjamd2gVwMx2ft4CQsumI0B37r
Jw0nZe//e/nUvwW6z/7EhdJ69abJvUFNXEQWZTckUh36UM+OybHF3ZMDOFplGwH06ywQbopdfscI
e3LGXAL52nB0lUfcVabId9v9vN3QIo8nrbtrVCJQbK+2uKeYNbkgrmumYSSNToqDyyyU4lkTj7rf
9YCKwa27PO7nNOyQF+DnOdtnpbdOOFDbZVd41EGyVISobTAC+vDUKZnZSeJfc45gVIr1QkVvjyhX
JiYVVyx6Izp+cbIs+nXpeYVtoQ6T2ggzv1W1m+XIghGYPXTbY0l8x+NwUwRXl4SAPiV+HFeSyerQ
5fzzUxMK9xgXIM2q9pFrWBXezPrz+q/7ZDkELXXxTi/I6S8YV1JWzXuSKSbPs9NjiBLM+0pSUWl4
SsOdy4hg+CnMfM5nUFYH04f297+BTTqLdRo7OFYrm3KvAWmJy7jz9JyOX2FBL9VgaPvtmLNjCe5f
jgeFLKRMpv3xp+M8FhkNpJN7/X7wL2o7gz4XJWp5KMtDgWtwHJRb4TN5NlPQsDMp4O/3OAMKky/+
x5+ln+lXZBuGqbRSwEJ0OoJ5zrt3lN4VTSQj+SwWfl+gE380rRLOcS6O3XfMuS547HfFiQcR9EXv
1sptmgLN/sH7mAEyKQqMpY8BdnF7KNMmiPPw9Gcb2boZX73tX7OrOhuJmcYD3yY0pV/CpwRpjw0u
SIsVQT0lLNXRWUesQP4UlLVJdx0SdFF0acHb0z+T0gdwrvsdUi6TovsxO8mLZKkAGIBC4eu6xkU4
8QTRHNNhi/cF8cEhWktWS0XNPu82w1x2mN9UvGgpuOg57ELPTWmZFlbzUFFZTiEf8fQE7JE1fT28
46TT+PtRrRJ1EFS3QoF7j7m2eUc78e7QPoy4sjngTwRPSmqpWlWXnM2vf5qF9R6GKmx62qEH4R0A
/wETVzs6JrOvYdAMyUwcudZNF9+wJ34XtkWXK3GjojPGHxfcucQmTPH6y50r+IkImqQNhO8RMdUO
rmYigNtv3sfpL+iAnIABGU0P1S0c9qrye2TBH807vPwUvzBPIUGP+onPHRDVG10DwYAzF6NtFsgq
6EEuV5vDWWUZ1AOa221P9s6lRdyTlO+k/thaSL4yOymOP8/BUsJRuF1iVjUThZmTqey2r1FHH2B1
g76g4m5AvQ5rw+HgSBlzPpD7dW3fwsI2fnzZD1quEbUUF4Ds9tBnH0DskEfopG3kvRBZX+Y4qcMY
+h6r2V8b3368tCEXbqvrLvLVCShhNeshkygajgG3t32YsdIdRqeUjfsWJuOKE8A02bgHItC3yd8b
lgozSxYs62w2J9yVgZtdwQt/ZcPMnRX9WnlVXbBzpBPc1cgnRz5Hjmln1Q5+hqbNzUA9IPKNxjUv
YfsGYx5E2HOFm9IkgHMh7PzuKP6c0tLZhxpXucRNqPv8xxf6YcfngIRPEjtmoPA9MPFOwyc++V5Z
owxw18VuEYwkwTsCQUsYv3ySpYTu4sF9uRzjUKfHaesVVTyi5w2yEf8oOKN1zIYadt3wNf2tsH+r
xGxs+3T8QJbZhAcrylc/4hj5LWqDqBwK9eJR8sQrJvZ52z8n1qQfApfM5g4+2DGJmFVHnCZqzX8b
PGOsJzCpifjkp2b6MwfWJ864Xuvoqp11uwPD+NrCW/i3VblAOYyMcnlVDfoZFPQQvZjnliUOOCvn
f3RyWnoGNxL32kMiJV8wHuDaoClAYtu0KBsKLZ5ZkI9VZ9iFrE70Dbn08ac2nwmFbZmz5HzJDhQM
jY5jLT32yHmG72xsVsfxNcDR12hlifoxiahOyYS2zuJ49QPZ8xLyKlkqxr64cgzHRdkHfh0BbLFx
qBvy/CFItFtpOiBzsI+4bkio0TK315iUO6xFtkBmMcpAaql2Tl2J8tOhCg7Y7geXmai2jy/qOI5F
+EOva8SLT7A1mSOXao0VrvzDgjKzVj7OP/4EccJ2XwUrHGny3VXrG6kOh9iVPE4fKpuJ46z7QrLf
dLYRtjCsmNusVys6lMfVdU4U9mOFUx2/zECLKnzQk9kzDtYZkoM4FeN/ocNFxUZyRbb3GPhYwUbh
woueyZ3yHAnf0PZ5d4X3/7GMQ++70/S77B0o238LbGbyxJOV9ILI3Mk0kAEiIT0rWzNdpNNnCoKY
lpGdILsTb/ev+J7q8vKHlQtmNeQ7yLVaUIoszOvPTqlqBJoTy85tsgKsid2JOtyT8sg4VpYJkFp2
tP7bdsFwQBy6clDF4vz8A3Kp/RfcNybywWY7Xi65kwKYg97UA2asKjzZPzp4e1uk9BuEvo2tavg6
9LUhX8JpRA1AJtnW337gy9lnCETl99r62NFOuFBKCCfqIIFaDDKgnK5tY5jsatJE/JRVF1bVmLn2
UzLVPK77ICRkVXIpHAWHwACpSHL//FO3WNCj9JxtJx35kSK04eGl1FWOaY/HBOMoYIG37kgYx+L3
Rtu80NmB+fqPVghEGiS6qYEhkoFymo3RrhtAageDBbIvJjqxOT3lAnAEPqQzaVyW4y0iIO4GAVDz
WgSDD4OMZR4wD3UZWS96LHz/8RoHhNSMDUcQGdBCRotGFNJSjoRNHp4UKtraqUbX1T8WKR3T7SZn
UydokPOnKd/tiklxazrIVyUI3oYQMny8o9ogxUSD3Ps1mYGy8RjneJHNhsKWZLS1A7NjTdJuVNTC
NQzkgWydmZUYC3i+uODPfQo8OVaZH0Zi9Tx7AksS3y/72xwotvZLfWSXBSi4nMjNfk+9z5k5KIJV
7qYtBd+uvzu/ogUa188jKn057diW7oLma1oT0ydUwWQn9sSFM92Fv7CoCWzMKWQs8wACdkjXmdjj
nqZxfxP/bxjFiNOvf1unOadVGMDr3Tb+Je1MK6vTQ+615E/c7TNFZzPSQFad8M68rNCgyKU5tusZ
epfnlls8ud5KzO2JXZjUT4dhMLBtZ/SpcT5SzRe3IgsOHkf5HcIJHb1j7hYBIBRdKu2jQAjM7IgW
DhRe+M19RJkTDywC1OzqX2tJYKXMImPXZ+5769gn0bNDSOXeIONE900ubyKjAZ3IAGjGfsqZjTig
tRlE9doc4YW/D0NJs93gCw1HT5PJI/fV74CtR4JOxq4lO1X6XTwsPH+IWK7g3e44rAIWlOK14RXS
U23tMBPIdqF0nZYcMrAp/6vU8FNDFzSSaX7zyJ22EXNyfb1X9fxgo+ou/XrZhh/gGj3VhMEkRjba
m76668ywsDpkiF3ghRIcuVgUPB0DW4Waa4XUiyoq4Ivxb57TCmgWBIRNt2a93Yw2Z31rFrENZQk/
6SiXQwVS03GSb843OyE8DVj6Lx/BUDTQl1RW+GeUKbbAe50v+MaaKVQq7UJ5P//udUjFdX3IikYa
/IYMBu+oOwmmoQidRII89Px203s7lyMi/8pSyodVZdoHQMsqbOMI1mLOZxrMaFvyqjrDcFU/adAY
kC/U7/eSoQX0WHgonClGpkLhgstOTfzKtZOriFrO+aPEbk0vzkmWQDDBnWH4vvfYo3TDDWW816UL
bmCg8jsolyY6Q4OnIjUYbXJHt13byuDIVxRMXPngo7XAIinIIFrrfx2wTfSBfLBhQcOsR19q9kJl
8VTxndJjLjUgK6luT5MR+oHDYM8gep24dARRPKlKDg36GI+VQ23P5RlxgEWw31usOY8L93RbgMPQ
S3/lLcxJxpr2cAA3eGp/VZ0xJHyfBulNxCnBtZLNCHXkb+20j/C+rjYkUfvTmivJzkhIHxHo8fZy
wr8V2ZifRvX5e+5isSkmcJdWgbdFDyM557wb1+5K4dxapkkc1UfjXe6sPEEtvSRX7MsXKpB8Zn0c
IQWvaYfnz8kj+87dhLwA7f6oUrvIAvXFvwHIKetXaRePGeOg+jmXGAIHoVZmd05ElrY3c3pAQTDw
JqUZH19NAyQAVtdVPvaZdsMALfRmio+ns9YYJzhvY1vs25v337lBYUdcWZVlYtieBj63jb+UrcX6
2RERcdalCqsJq7tdfSZ14+zacvOHR2sW6wncFBNxNFKIsilB/w3BTRB8xXCOLbBvIsYuWPgL7pyv
r3utSuXUj9uuoJCYpFhCBS+te4M6htwFyLZErwUbefPDR5w7Pc+CRvoI2O2zLCWPUmYTYB/PYUVh
m63UGtVwjVDx67j7RHpT67w/7Pbv6bAUxM7b+a7LKdKCGzKXdFFcyF0Qb5LPxHWWS2sZIYZHtBWB
fbfmzCUtTOrSV4N4cRGuhkApucq0GM1MnRjUp83Eq9icbcFAkIvZHmtaJtaDFFf1AqSrr7LyHtt1
xmI6BvA+Bo2YOh//31NCy012SdIlYpD5je7PPXIzfQBpBw0I7s0w6R/heqpVOMEsDu39z+uT8Pei
kT/7VsY/B7ot6p+vqbF7QMx6SXN59zGPemvJBjqkUV92wg8l8QB/l9bwORR0u0RsqmA5omNX+EwQ
KoUET2GdRx14zv34Q/rcfRc0maoZPFaAgKSvtehReVWknaHXaJWEB+DeA7TyEDN1BgK9WHWGHPdk
D5YyzfAO7/z7TTr7LNaujtXtAX3G23rw8mcvCco3sFhgkDB7emBVxpngC99lLVNXi7yE08UCmOXo
G4/HwTEUqNNIouH9kgJSNut6/kxbvjrBAKff5GZ2FeIXtysBgEuKe2X5HVLNT5bBST52F9/+gvxg
TVI7nCExkxIWKd6ziFcKlrkyn6r/CYVtdgXPUEoWP/tYPeAcjkG5spDexIcZIPqg2f7zJR8MX885
VPfSUQpGZ317pDfSuDlL1aWMyCprLiOMGqp7szL1Ty5pSS0HmE29iLAt+o+JYgL3RtDcDqVbVd6j
IgApKRzjSWlq8+6eGAd3KGYDWVEMc8FUIlvyFMZ15a51tc+hPR7BpmyWAHPUyka8i8skOFSyCNyh
3kaEWiWz2sMFL4iCUCv84OFu/LtXiwxMu6XbURwpIrHvEzW0Tn1+M0uEU/bIZKJGpY/zudrzkRXK
7sEc1yW+VNq0Fii7QdnRQ29LkG/wPtlahlLBIJLVB1d63uBm99t3YgBnCy5/9UOV4lOZ4Q2vZv/Y
YPOqbvmqZJmetdELpyLzLMyh06BmlBIh/WKg2VzfzOo5Rie4Am2gJTzaR4GIFWc5lHkRoWXUxmwx
5RpeSZ8PtLMXcEJ+xyUE95tBIWrXusbRjEhFtM8VCb5dO9PAohngVz3b43ZnRKytgbgKf+cFwo5B
Tiq+nEoUg8ejwjRZbjAF0SICSjvBp+ioMEpxvjngVefDz9Uf0QryouPriHdudvJbm24wFnyACZCw
rskvpZpUjrJ7sip8fmbtfziJDHrcaGqvUYVcqy+wXPILHDpdS9psQcrDCMkIZB5UhrGqqlwlHD/2
wAv6+jsenfIC20WDFnBrIptvMXdeXSeP4owSnyVyQ4KW6oxL2oTXolT2/GmPidbXWjTIEmsmNKEz
Q79WoKPbyhIO3tU5aDGThUJhjBeRMvGybOabAO6DJNtCWfq2HmCzhMSccoRXmPjTAmHad9rK65zZ
5VWrk2iVP1Zs2rQyK72pJAt8OQvqS71RAAEf3nkIXX3MvicSG4oRLMh+MII8/xqDe6pLhuj0QW+v
6Osqm9f/ZJFgxUZGasFf7pmliv+lEP/YcRk7ZD5NykMK71euV6gFnFwbn44Zyxq1ELKg+Y6EjUzN
bGQ9ajCwpxTwGJMehflfP7q4w2z/+JoVg0IOQYCfiteHNlLOuuVD/xa0vsYDFTHCKDPIj2TxJDXM
/Kaas8+zsvnCnvTFMi4GDoji55NGMMpalbP6+gG+EtK2bfyWm6leYq13TQ5cvOvgbaa6DpqOnVKt
OBdstTjoCpgi0qsm9aEfviP7dZlEWvurkh50M/aNE/zfeFcN+rO2J972T3H1oywYxTDgj87yYKaK
TSPYGqnYL53cnkc2TuAYXKHoyT/lz6p8RXmh+KdNjfCdNHc7yw9jqCIFPgpQnwzSz4mKZJbJnF70
cnSUab/NR84hrz48spDzR7MUvbpzygYaM3pG/8shTmkNSeBapATb6nxsx/wtVDWILt35SgjQ/uSl
v+D0KxrxqG/ysqAu9SQZZlHrryx1mBejO6N2plr0Jlcmmgai5Vn4cRAUZ6aNWzhseh2h8hFMzns9
xdNor/W2hZAKP2aYbT1n7Up0EmHQqtylM81/RoDEokAdMlgiyZloULuTH95GPkUHss7HZ7HmBn//
JOsaPQ7aYz1XMAVRJ3HcZ3oepjNIX15s3wg2FEIEVN7plivy6IY+2mMcPrvZxM5T3sVJmiwicuhv
ooP6h+k4PIq3afwFtO6Bjay5+5jPgKLxnKpetXP+BXTQfK8Z48PbIHpiSSahnhqM8hc3rQWBLRbe
37Pljn8lGMmHJuxYUutkH8oi+dNg2lGxXLxuNmWENVmALVYLf1mLzph40y1pWH2dfaO5XNkchSlY
Fxid0yMBxg3i7DLaurXNakUsZN667q9C99MoacURWRNlYWx6G3a532vutxAF0Eee8r16GCAV5er3
K+Gy9F9q4qgnROCqZDppWvboL6NpqwmX6B2RKdqTuyyizamrkejftHsgS6TXvdYNVgdkPEShlImz
PTzeUYqszVlEN6+XjEFMpWhbFNjo8v5KfXbDrAe+VxhFTjLWseiG/tbrvLpn3zLy/I7MB223iFYH
XCw5NNeS54GXFC1cX+wrn0msmgoxz/nt7DHE9wDOsPWRW3d7M8oTogAFAwZNO3GF0zPgYfRLqBzR
Lq61Roy2lNnpd/FzYW00zTqD4iEvYf9mMWd8pXtWqnOLP7bdU9dLiB4XnHk1wKYKhWyEAI9ZkudX
Ugp0P5Fd2Ne6XmPwXQtU6Vif2kxXort4N3QpWkskYG3r5TUYmwgn/B5lHqj0P8qMSS6+h165ikVr
O5v4toBC8JZyFgTGtxfsecdWIoO0cRVdbABzmRKulLulUwyUBglfInY2nx0btCQaYW9812JpZ+tH
e3AKQYqloFHu/2FHzeb0QiM/BWpbXLgV6Ta/h6ZNjCPJgfF4BEvkhE14cF2GmmV2XEvZSHY74zeu
ime2txloG4Uyyp0m3Gvw7/yybvVxbdHjUKWTmmxtTdkwYw5gNsQ7VmnkbeCm44YkomJJvZw1MxVp
fhM8EL8/6Z4fdeV3Ln3tk7vyted31j3leZrcffII1AxXvk0uNAwrK6HX9s53L+9Z8/4NeGPc61xa
YT3+w20TpQPA6Mpke1ko3WwWo0RyBCGDY4CbQb5lfPNiFUzJDdNwGVO9hEYrmsJKX7QY0dyFIWmU
oU8lM4AJ9DhC2OIrBNsXXc1foLaIyJ3q0sqUnvZEXfXtdzQ9n1/Cf7E1sT4T/SZ3Q2qtY1pbF6ls
Q4APpizzDipAsHxzBs2DJvzpjUudCOMO8l0ySvzu1EJBqvPMpcb3GP2qTNGIGBzVixorwb6uIvKf
qfle3wOycxz0AcsBHJjPB6VUn0nKNLk/1GIQXQ26FqCdZH2u0rQHdHsNb6OWvG2mVNK7zZcVW8PO
mtVKIXVdd9hSaI6Xui93UdowonFiOdROvUkEgpl8os6H20OMZj9xoXt4jApSM2sMaM1bAGJFY/ru
+mQ/hn44/mCyRQ41wOPdxHFNZR5KVmB/pVfXMGdE/XZv9lNzvHUyeMdAoaXMcRqIUwRdLtA8J+uP
A6mZ1iKOkpubgAsiSvNilctofnVCBOwrXiBOvtIkG+qHs+eL9mi9PzxZG5jChL2bqIBVckzjMFEo
CfDYaTEXcd/YEzAdAH2wPnFQwfGc7yjIk7jqPUppTZm5lRLWs9gik6REkF3I061F4jQLiSwl8nfe
CM0ysIQVJ8ISY6FycG3ukkhDVEJ95dVSD/NvmYTt8Rntx50IJr4CcmJCXhpj56N7TcIONR5RVXIK
CyJBkr+DNYNtYZXswPJaC7HyhycWYReduyaaPhVQmwYdsbEiNRyYFlQIDd4+ROmDpdOZrn6+lSCp
FAeQMfABMQSdddC5o72ogdWSGLu4LA7xEeRq/JC2BfoJMzHuHJBBfyLwxDf9hHQh9x84lf5jpreJ
xlm6fe8V1asWdiA7tKpg2+CmiDyrOwoh9O8yNXjf1JANnV1NfRpmsn1vXmEeu72dKD3cG3Y3AwTK
1tkZsfRz79AZVJuGzE0m70CaFbPzvB9i9h7LZIs4I74Og66W+2o4itYVqX3PCvD2TtKegOoMQQfx
1ppons5i7VXl7bFfbqNjBnBWW3x9UK/RK/8zVez7oozV2hfiQbY3wMQzPE1XC3OWzbec+PUtxnkR
1XOMfcwqFno5nsIYm69YO+lgXAqV4gNBCL8wjLmSjFImBQF0Yyhjd8SlO/x2NICor/65DjUf8vAN
WP/3m48FeZKSFUFGB04+6Dw5rSujFE4EfOxPtpOsZBGxjyRhb+ETBtoMQCKw1/dfR/H831C3mGDn
qYYEzlroMinNP5tmtCodIDDKlBiOOiR8vh3PhxJJ5Dj1ydyuULxSwvl2ONOv6gq0T9+D2Lb+Vq5p
3xfVxKA9ArpeXR2EwP7haGLSVac9cWr1hBgXntHjmFV4B8ne/puv41JNWcPiussWGKk4N4Sp5R/q
D1VKwf4zR+Z0NVlEYvsYCpx/uSI3KeCq19Y+uTMM8vA7kLY4GuEfzCD2Z9jHF8Fov/3j8Q22Oq1D
xOFFDh9U0JZktuvl2vdz8Nj7F+S2XgkN4RX3kN3t3U/anOx2eHtOIOFUaToipXFSnFK8hB/Kge53
MmKo8oTtuNvkaRRN3ZTxQ73qi5Rx4UfojsF7PyY96OCesw7wjitAzz+Iw+3O8OPhtHyMBALMK810
ogESBwpldyPSs0B4fbES3qZZrCeRvBMRsxwkRGeToBkoP6BgMX9yxRnsBCzNORLNfvbu4r+fehFQ
LHL1uw69K4J9/eU80neHpliolN5TASyV83Kwt1iKb8D07LdhHSKc8styL//hmmjGPZb8vw7EtoOB
TWk+BfCkkpS+fXvWIaQtiT+ojm72JSZUbUHpw5gT3dEeprcdTEUW+LhWqQ1eyjGcc0+0bs0XjmMW
A3VThAwlEkYNhg2Dyk9CRC9L4xp6sA5pFJHXfNsuZ/b9meuxVTYwdhhytJILrD6M1Ur6D6cQ0GtB
9GziXUnt8eJVUHnW5dPoF8Aca2qf/BU5xfQ1cRar8YaQ7v0uKRm1wAcKdZqH9/Xx9DlYW/ZexxQV
RT24mU2Iuostc7lQ/R9Aip6S5sbNkOkErU1hlIXIpQebs8eKdko+f1riZZVSkL1zSYr0wRZQLupz
p0MySvmM7Jbft/0REgj6gHp6oTfWW/Z9q+yhD+hSpmXnF7/mnBerT9pxsj5SyrNISrFcoOs0T+ij
2lnVZRUpxY8EnGD5/IuW7O4Yc5F/1km38avdaYyxlen6lJTvL5oqWQ/0pboQ7C9IjGl8O1Dv5IiG
TY26SviemLkZqRIlCWGjk6ib4RTRmnOcwCVqcu/7P1wkzeAnaLpfNkYohV90f4L++9uMs6GjL++z
PCjn6KW5W90xqVMoN+BY7ZKf8aV63nBJwEWNKQ6BvMnlaCZbzcP6QTFLJND1rOgKz8JmD2S65zXG
A2IIeQyAILEiV8ryplP0QjebCLP2+lW97KjZBS7ajMySyG804H3Woo33HhG4LPn25I+pgl7dbObm
MrXZ1w2Cm9vm5VQhbCs7ZEnvYGlQCFMiTAejIVtxupjuYJruHx9PFT0LpV0T8CjWWxj91pTsDDMh
fT5pX0ShqMoBpT9Bh2fK6ea6a8Uo51Ve/6RykYnLoQqa4nQ9PgaeDum2YpTBdxd05XVul8aeEq67
g89pc8tBwmTY0zLpk1GqwVjj2ASYgYN1CBDu5yZSM7vr57g9WIJD/eq5QdYG1WjbRI4VOb2xemK9
k9N8hVQ/zWq184xBbuc4QEDdNCttUyJpgkvKPxh2k+Z8T80Ef+7/3uGLvGOHw+J5aD7NPLUECqv4
Tk0Ybt4j3R+4lUDg6dte/IZBGoVPcXVf7aVVkS8K7yMGawi16qlimBrAi6x4PiinxrWVxMSi0gTQ
5bsgsYHDzMe11XWqX584RGUnRG4XwIFHuyV5aQ1i3ogWx6e4B2jldtW0dcXJyADwGe5sHc96HeNp
7qzzTiNNPIdX5B+joGoEECaK+VD6p2esgvwJhJTDkvBrZGtCM4hA9RLKkSK21WmaWCsIl0yHjfya
BcbEOQylPaWEvfA2LLkZPdwu6vyi+8X40dxrVcm5Dl6FNQAPeh/yOipZmCiqv/JG6QQVdoFn1n3A
ldh2iZ8NIodQJeq10ZF97JQM2W477FMVoSlBuMdPKoRW3mmEePl8qk5K4uWMuY9tU5KEMK0udnma
v1Fj/fmz2Aymx2gTsZiTlSyvdRX82sjdXpJbhXzd5/gvljSwRkM4SgvkswwEJXjzz5HryoMcUOYK
C9Ht9lJqyzurJrhImcYuR62bhMJaFuLcn9GmLtLUz2n8ET7EpgoGLod84dQeobn63XzSblt+R7Sm
vm+/wtEH0S8aJLZyp4p0EDkr8VZHzc5P6CZCYGFfpwfQ7tC3qaRx0s0SSBDAkKCErAIbHCFioHIN
FHQoFzrovNv9n9Ps5UNIBbYbh6UtrDz/q/EdmcHOOWrrlVjRw+QTf5S/otFgkyCgY/wUToF2sUQc
RZA/2vNV9JSTzUIGHlvEEp4K1Q01/1Jj+o+FnrsLti6QRKS5vghaVJvJSi/pIKAUB7SpVTE5U+br
3Jdjr3ZNiOgbfoDVUzkRXslYgFldalWuYm/bp/7fEOJbt4vCTEkAsokHsFy7fz0yJ+tJ3tufZ6rw
2tqkwJo04Unu1STG/394V062e7du4YJuR5JffNLLJ4+YpqPDeXRDZ0eTR48oOk7uXsCPaQ5456zg
yUe4Zn84EIJDHDhndacFpxrLtRHPM1fcJGHkC0buXkVUO52wPN+vOcwY0XVoe/FCF7NO8ufWUs3l
9SU8QHPUnMDvovT62ec2HcV+N8YMkFOidWbl+Pad0hdAouspRIKTjr6IxBkNpKuD/nHNETuTLOjB
D5GcWS89DKJMKLHYUuP1xtkR+1+7O6UZ24zok3m6aq1ki+Z0BOeJqebVx8KSaj/7iPL14Qy3Th5S
VqnGdtulKm8lPdTBtf6PvuhKybQM8NryM3xGcqdEOXS7HPhSa+e26tYcmOS9pmJOe8p7zXisapWi
rctU6qxMFP0ZNgOO6f+jDRWdfZM2q8XM2kAXLnvwttZ4av0Q1VzkZjVz5ni6PmkEvQAZo99t17cF
YeH9B9pBwKql+Hzud8hEtBRIMmBGM0l3lY2ymTnXwXVi6h1ZkMHGI1b798Gg7UL5BYnitCdgKVG8
SFcpliTtF+0PNgWe7EQ7xTtL3x3+BRU5qkzaaXW+LsPFYxAE06hDe5/bgb9yiiARMHuVZ/t/Ni7a
NVPdHgWyNXzkzALoJ4syDSc2I6K6qkUPR067Rtvm2EPWsmkfuCh8kkcLO4rPYXl5hmS4+PRc0VxI
u5BDYzuKBscK3K/waVYPNhawAv/zS7UvFEw3WBLK3ncBubOoyJt4qDhz0xPGdYq+VtBz2UUXWP4k
GXeveVakKY+HSjlbP9UB6+WPGQjx/D7ccN3rJe9uGmmKyKIkOsmzpbXfr1j7J+RPldC13p3EOZIU
oilmPdJWqy3+pXTe9/h/746aP0wMU/sySHPhj7wUvxQRqtV9kuRwPtbsV+ApeUUhMWwMhkZtu95N
TjxQpE/5wFupa1snhQVgVWJieCrFYW+r5NENEBTWeGQfV6rwCTTGboarrKoDP5zxEkTMEPjMNaAj
wYk7nNhUbIuuXao7XE7BeVCTKmxPROIFpqn6Ft7yD/MEBV/HFBzYjil4jWq21TwY0VEjLhiyhgnG
wNU5Q0H7zggq98sqvxkHH4IUUJx+fndapZQ7mQr4uWMENi0/efEQ5v3traj3cX/JYBEt0oaZFHjg
1kjBoP93bYfDN1Wjs5vnBAXF5SbuZOmmdjtNm+Cfms07C1dMMq5f0ofs2Zi50UeuT+n8VQwuJPgp
2qPMXQn/fxnNejVrdAxZUQ8ufhn35bWg745cJ2AbLI67Ple2lzMl2r1lk7T1tqw0x2d7yGwtnTeZ
rIWV4T14Ca3fK0AnUQtwDAEfKnMAy+TQk4vgiSF685CpOYoxGFZs78iCFBGrXSHOCSOiidpXfm1X
es0bcZA2W12VlSOWyYpwl+pNWBLpnCIpjxQ4mgiozm8m+AzSmBgfOAneFwQSsBlQr88sDKbraRqn
1jBj9X/MWJtF2KZyGmJ37SqIkqIZdQHFDZYqq5a0rfunLciQ2G/W4j/tCK+2NV8Z34VglQ5CfGuk
Zot6PvNMQ9puN9LNCCO3FtTpoT3iyy++IeTn/sYiNthlPqmIfXNat+NkvCPYPbZ5edIovlZGuURY
I33aHPUinsqHUm0jdslxrpbGFhiZ9luUlznscFGBYkWMr8Wj0f6cx+NIwmDm94KIR4Y9bkw4/XyJ
ksp/lFsj7GECC1Sw/cUG6tyRHoB2Auem88AkuEE4tmKcRGloKbE0eHf4UuPxRfUEwGaOwOSmNpVa
xrR1io11bHuKcUxmV9BGPmYjYgbO6v+n2Z9wa41Pv3D3DZkcmH6FdMLVVTej+evCqF2aGhfHtEMz
7zVev84lpVXGMoQ9DBBzCeg6x38wwdHMLTgB70YhPR6aavYQ9tjmRNL4al1Px6WTC9X3Pm0X5omn
FbYMSrcXZyC5blDsJKxXva51LOoqGJ1Pl2haX4hSoh+FOlcArEv1HiOZb4djPu/Ata650KQkRGj/
i3nRhNMq66rWW02E4kml+YnGcu7bNOi4OdGU8zRbnpW5oZnM6iYmOF3ajgInBMiYkdCX0OYWX6LW
leOQMHl1BNuQIk19XwMlfeWqblCLgm14zBGLu5JwHQkIZ7Ek7ktrsCo4TWgO3E9CWQgOyPvQqPPL
4KL/IsPxvyKt71GLB9sOrqQz7Z20TlNxN3GN6BDGNxhHnWJVCM6BS6oTNPNepd9SMvYlY2eJd871
tPXN2m5bi5fLGBnkS0UHHBtiWr6pHUykHB58oO+IxCiZgv9qeWjytupvC6mlbMGMSMxI2R+YDsZQ
qz+/QWk3vxNHDf1I/0nEIb55bm+1XeJYH+N8AEx9tpeounVesEidB6QqvdpOwUfihByGO+4Bzh43
FLzZP5duORGVel86UcvAg8j1QEgprsj+Nwm4fnBF9oWQPIqX50vC41jR3WUdf6+YUftovG2EhIQJ
7DpeBIDXvGoUueP9Ka5NjomoA0hmPL31iABCyNAAELcI8JI0dGlHZiiftwZh6A1ZDXb2n0LkrUt3
s4gbK+wydAjaHUZtqRiKY4P3BN/sYC4w7V+zBRGbeaG2Aou5rH7cBFe+dft3mww+8IDYd2RIohBf
x2/Sa6nh4XG5zWPdXIfPAX+G3cnmijedcS15AJ5IaBDsrzFqCkqIGIdkvg8uJ70o44DS7KpAkt7a
i/GhVyf9siiy0KuSTIVkNngv6lpv7DrtREVn2gxzuVbgebgQ6568nhXo1NX1DJh+7Nh80SloivLm
ZEmqeeHLCaMjc0GZF5r4fNHznI8ovQx8VVB9ZdBAWgIi57Z5aZQWudosKYFidPd9vTkBm47RV1Te
vT+rWi7bcOmtXFF4Uv3boiNdyBNLy2uOsPdRVbDEAphK8ToRKq45ZjXyoIBM30IqVTq0+mYWpHSx
yIPfw1/pDu1hR42GeSR7pHI4n4I6huX4T9YIUpwZY8NmHVk3qAy+PqlJ4l3y+2PzaOxFLC9YGWIP
Xfpj78BISsM5F1FbBl0g7yBLFxgcG3ZiDtyxcvZSuy8Ais1SEk3vRmDzppuanzOh3pJmsqFhMc0l
s2vTzjLvPjPcDiOnUnsEPJG+Owe/f33d/NCMA5BJz4rObbiCYeMEtKosKs4k8vMH+PXwJxiC6gHj
nsVQ8U0ixw1cRD6zhMg6lhdqBQ0lsdDmTMveRh7DRegCldqVcccQnrsdYLvN9pScFelBIz1O6rEj
+dB0EqiGGSNSkaTbN8gXNuQUlsTbEMsPuPDo22Psyw4DW6BytAcyUJtvpgcHAM0xoYAjijLQs072
3uoYbcgsPhgk2td60v3sXgiy8QhsUiK6Xj6x215oycTk6k1vV+gPhMtMsJoZYPITeCeblhVArBiK
sdBZz50qf4EYzb3T61qcne3xK5NPFr1Ow8IhzZQSXaibFaRbRkSqoQhvrFE4uABnJuiOWr+OvKNL
iEdK1U99aT7YSzkTxaX/lLw/EtvLb7hKsXBDeegdODH3YT4Lb3WFpX4I7dAzLm5EscrMfRkOsjcS
jDFrA81tKvPaTqrDhdP6nm20cl96h7p440qJaLGzrmhEJXEtdPi0G2C1N/VemSuzAgAdScBbr2np
ZtFZfYVCdspVcqRSr7mSnrP4eyf2mOPu+N31PeKJe/S6VDSwu6duEvtX6FlzzHrP61GGlBFGKC8U
TmmbCYcEtqq0B2sXitIUSIGwj8wN5j+dvhcsFxPgeqaQH10EzbI0jACvGvcA5FxlSjwj8opITYAj
OaM+cDZ4t3mSHZgU991eFxC6NTlwcH5PuydlH9GOhpfcy0naEpeVWO3RfaqqrdRiJnR6jTndeMgO
AGx1OfF9VC0qeXP73C+b8uEUI4NryVmgvExUm5SzJlzSfH/aeH01txtrCii+tPRL9R1PUtuYhWwV
hIXR24rff3wgMNWe2Bfrp7YRwj8NalR8h2WRcoXzTHsM+BG/pTIebN1HRVw2kK7BiCq9YQfXLxx4
vL/lJAITHDHfh2znzl8vkjEmBozVnwugT5NtMe8RtErAxdrqoz73O/wGV1jsXBhaPDm8UFnW8Oz3
mfe8P74aOwkFqlp6qZF98+Lt7aaS2u35peVEdtz9quVN96xNXhwKE9pOJ6Ia7ZBaEay+yDS/8ebO
F1ooWvXEsna4LhW/OWsAvEVjGqEhnGi+W23uyGT4HzQ9n9tVEKgq/V4AFiT7vKPWzHTgp1kcX5Vb
cy0cy3zkFXyT+EiDYjy63Ds4Bbm4jZ17I8UVqUUj1AKs/pJD+/ZYRku+qf+4tBZmeWn6L3PuSeGa
2tNPLmmxoPOk+BeFB+UdMwLCbxF095TG5P1X6XQp83R3t2wOo6rV14/RBnW7BuLvuLa5BG5AKumr
VZkfcU7M1fXp5Y1hFGWQDtEQK/p3VTvcaE054GKtFAPMkw0abJFr1nMXHGRV2bMuxa3RumLKAA/V
9Lsa/eJToumVuFpd+0T9v4EMsaf5PSqsXAJFZ7MlBZ1kT6TQYMYV1xEU5P2bL3alqdnf4zdVSnWB
0/SGz5cCQbgzsUCrQWLor2H2fZBrPTdk7YLu0hPcdY4kjplj+8QU6oGRP7NnvOKjRYW6frPA+FWw
EWgfiMhBk7pNR+horV2JB+WdHKjALoMi+6CzbW+ORkfLpIjGniVagoZQWb6bIF/NyfJ+X7NkaCN6
Zm+/7oUNyIgb6HKQre9PwKBklhw7thAN0D8WQ9vmLzGv4pXhM3D2xWen6KU5GK/WmPc//A8Ev44J
XwGvMBYZH0+VJDNilbahfocSx5Qj35NBbAWMWtYghYtwzPXici1eVOvll0F8Sppldm5CjV1srq89
n4qtCG6mouxm5lh7sxhURnNupOfYzJphQOBHxUwSaJbAb1DfK4EIZlAxICOmIiDuhszPSQ3EunHw
+jpoAv5vfDxltqUbrJ6FD45TrfMOHpjsvMsGnGDnBKOVVBQj2rXQLR09zc4wWVChovbRj+Bq89M4
XEZ878iyej1ZJ5QesBIyiSz4I+Fu4h+ZC0/pgrNWqTXzOiJ3IgMjsgISdY7nOkZixkLwycgz525Y
o7IcSvp4Y9HvDWB84nPpOPFwDCiOuW6PhVTuf602ZOJsJLYt5MNFRpsMq15F8bOiTxtEadaWxCbN
Zdh4sS2TUoxV31RQjOGQBazaK7IXsogvs5ZBXqUqh1+WEMBrSd/50t0hR395VuxHAtF/YEANGAW8
atReSZ0qOTH2V4jSjs7luu37g1eEEVgr8Ete8LEl0ocsGCeFXJkLh9zHqvLjDH2dtLYEwnP4+xKy
d74Q2tfLx/o4Of39R7vjogb/n6Ccgf8y9j79KeCLpAaNVP4MAeROEUYXt+o4eAp2mGkHJEOYv6d9
9jgNRY7HqHpNSH/pwJN/gBXwpYTY1uCOxxM1QwLUUDjbkWhkusSJAeK827HnuecnH4xXxzyp93Tn
8rPT+BM1aa2cqrNc8OYy0EVLGMCytA5EZBj3yFnBoIspdoeTBZyvlQn9gJS4fOAPMlz1TY0pDP77
ds+mNDoIjuDA3p2w0PlS+3TvF2Zdj9ER7zx00lwlIHYEABJWFrkorCxJ8W9xJ/u98EI8dHSo5Ntb
S5wQ4WdGjE1wRDtKjIbtiUxmv2foVusGCbikHaKlmuVAP1fy66RLWfY5UkwYMe4IF8TudseIEYTU
FM/w8wwOapjmTXYFZV/sC2bkyg+YFRW6wK/OLyn37EFYYT+/jYxAtslj+5OnGccNK+H+9aJWy3Be
2cSrDtcWLhDHf4UdpD032HKfNLg25QgR0yrbKidb8CF3gQHtPzI0CC08IOAOCqFWneY8aiKXO6yi
jrh/7CGIOLHj+rPG5IsAlXd1X425SmhKL8nHy1VFGDgB9UlFrWxKPWK5jhDD5iTglmZH8j/5Wyc1
VV+H8+wsslAxLoiw8TsUl386T2U3Go/c6KzTdFt3CqgV6euAvn52PcZY8n73f7mkPHUqBCZ32lRl
LGS6uf19P6yXqKWkh7whvkC4kk3n45WJ32/ZOZbnau4TKOoiYjrFdYqRHAmQ1hExrC6FCyBZyaE0
dkqnYUEnhNsdWvHuN47wNjHTnnXNvOy5lpWZWLT1+prRUuwOfy4eEQEiSV8FvbDDazUfG5/o7Wjo
HGNiAmYkgGRFyVl+prykCnIO5qn0frJR7RZB4HsvwVGq2ZUFtTVGTkMnPll4hNT5HOLTd9lMp/0S
mIrBjPV1npJh2UKBaOBCCmmHDJBFm4pPtJbmKbHJiQqPzWp0ALo4aOmb50yh41R5+OxR1XtK4Qne
2/QIUJ0MfWNoovdCsYVHm8wWuQs2EP7Thpza1vmc/PRF6EC7F/JgM5SOmz4C9AjYaFclF8m6UGRO
+Co2g5UEEO2vBR33lpNPe5VOCmQ2VS49grvtyxzPkccY1U9o4ZA+0V63eQuHYE79YkLfFheFGFdW
7xVuKUVEL2vCy6XQY+ViI+vDunn3tz9hI03zQ1gyyizHYLQ/R+IqOl1rsoEJqJYrA6X88H2caieK
w5vJwVw4ZNECiltxyAtwtYONqcZeDvt05uTMT6sx+jXkrajAYPKt722qKwTw9JmcvKXG1/O9B6Nq
DF+93an6iKV1PGrjWdInzXNLe5xfbzxWpmgB6cp7CzfP/FSJ995+402xB0dix3y8PsX+tkaXX28F
W6I8v4hzuarE30CGKAu30o6xdU5IlINlE0M8399Qb30bdASUFXangWDSVuZ43g8cODlWuab3nY/t
Wbwq+RcN43SMnhJ86ahTAtoAPqkyey0A7MeP9OMQPcfl8X04NHqVgcRTevmArXRQTc65g21FtOIL
23I3xxOKwZIudgE3nWOIxvVWCT8JOrrvWMRZxBxyzUk/44W1l0dTmoAI+o95BKmys4C5KuMbDtcU
IrNbt5SUsNe5N+zaVVlwtJSbVF1syYbrW1JYJMSgVJI7WNUTAoEZCu/e1A9LRYB8L2ed3j9imBAj
fMOYmw/spemRr1wVjvc2kcYNqjgfzFLEucVFlZvrWIeMC2k0tWHI0W8SD1Y3LW2Bvd+9qzBDGVd9
bUZBx/zlzSRsuFGhW2rOmN07Lib7dCtIDQ1HBpx3dWKDhZavVGQS1QzgfQz0hydGJsONOY0UNPwK
w+kU1ME9w64vyV6tdAlhP8+LHBYVRryO3K1ixei3jR5n04Codq572XrVbs7l4oU0H/Qi8aki2OR0
/VQ31foKHqCod9cXfFAU/Bwu5UVfPRLZ3oUhIFCfPrZ9lV6qtprA6K7npONS2UCwuutrXoyRbFmx
E55mQU5a4naP8ADp9Q67ibo/A88NAUWWx+8x1QW9iu9pMHoooseh9XhPXb0BItCcAM0A8LOZY1fV
gQh/15n0sxsx06+FFfxnAsGDduPzV57D2yELiHh0HqmvzNKrCpvCupToibGCUa2z/DrNUpGI8mrk
XCJirno9nfNe+7vsH9iwmwJdO3SMG6awMV17kpenwHNOILat8F/xzhFY8V1dioTAD9QAf5TKU8S3
LviQYrZxn/E+xRYLlBuRpDrYa5slW92yIxSBQdid7yEomlDMAho6ZTOGzyE/al9TVAIEkKKWl3xF
0MhG29Ec7s6sBcakUVSNYWM6d+Q8cU4ZDfpO2xFo/DrfkURTWon6i65HV+aObzCCVoElQPf8hbXX
qD/CCZTPlLpHx0+ebttZnrLnCU3ZLkHpE+zBpg/JaBd1m0zRQLpWJSQWil+tqKaB6yYUHYL04ncn
RmPqVgbnBCBcYDuAj0H18ICUoRJ4maLEXNA4ubO5xNGwV6x9xcmOY8XDlWvjKvDWMLg6+ct36wr2
SrIsjRdzJe2CkfU5nHHxP+WNN17Y2ZzTuC7CZlipibgCqjVqSWbgw+yfs+Agld9hr+4ujAj+fHnY
O+EFLVjPWMwkDKcyzSk6ca6QQts02QKETAvVuhuOQQ2Y4PEiCumk47qR22aj/3MUBQWKzh6HI6ZQ
PCd1uQcZNRvHzjQnPG3+oTOrHuZb6Gt2yAQHuGf7LZHxO19TeDvpC6508kPbVszHqid2KMOs0M7w
jItWSDbTL5YWINc2EvVjo7H2v02CuRnlU1reHJBqixPf8YnikVwvWZHZ+Zt4cJHpVpobXVb65NG4
ptfG/PdLuS3LifbBwaYByME1vZsyP/8cUReyXqP7aDN1nbV0CvcutlH4weW1Tc8d6Wldw5zg+SfZ
m3cOg8f+mbD3973+Zz9BJVfNra15JHIesrvk8BPBqve3vsvP8vRtqt+if7bq6Sv5WcxjdXuVgBZt
fb/ZmnmCPmCZpPE4seGAli38jWSpL/adC0NLQ+jH3dZrvYP0prMqtqxGxE2ga3yqFTgoVKKji4im
0EcrTIVxUBwXCXn/HsZtnafcO/hSMgTyJHnjZlqisRu09WfZZCz7ovgcOQ364Q5Om7t8hWa7A/pa
GSA8mej0/KMviQtjWUtrRII8kOYzgBPmJF+VTju/D4ZCO/l7t7hcQIxo2Ud46WBbR/apAkdwcctu
3J/uSz81mSkPI5HkgjpycFR3kf2VW5kNW4cZisxpAZ8d03UTWc/pEN8NeSCzMV09b5FKBsp8RaEe
qQSY06J85gg/0FS8XlBg9KyywWsCnjUMH7R4KZXYnWltJ+16zIU1nXO4OuzJI9gmiUg+xgunQC6x
p7PI7LUgX9N/RyJNyS+MimATZHzGosDyaU1rdAZKW84GDDLzRw8VNhX0hIXuVVu9WH+lOT9xVXHz
3l7zgfpxhcpvUOFGJuMbWhcUY3CJ/oLrihmd0mMM6FYM3TBJJejZP7sq07AUMhXvy4J3V0BWUt1Q
hMGkLrolqmKLZJYzJywmYDLBD0pXQVRRTHCBzEw3weR+yRXHuhliOmAL53CoudxUQQKr70pCv8Gb
HIOKI2ioknI+vmBYSdOccqDOQ3KRSdg9szccOIOWiRDBr/6bH5gjXGZhojglOjyXGRzNEv9HfeB3
k4Ivz/9ca+kQcT6xRjGHL2Hl0XzgqpxbDvkafd9+GSi7Qczpm5HDH8gW0WQR+rCOmsdTbIbW0/zu
R/q0h+rXg0BiEnFd14WXOuhQmIt+sjuJ3ZOfxL4hlil3lbCTW0Y4BoEB5wuRT0Tr9elM3dy8S8zg
xRFoKMhbz9bDpjCM1BPxk+b18YhgBXIJf8p2UcAXuvXHDXzTC0aAjFstII8owlEq30eUpP6CF9FA
vodP58U5Oj9hxqldFOzr+K9V8Yd2QS9A/SQpPMOiZ7BpDA+rmO6PsxSvtYNOWCT6QWl9uXGFiL6Q
j1fRhQnKdFd1k+ULZzGtPMW/TUCWgpoMk58a00jSWXz9TOyxJ3oyl3CHDvPPN8sBz2ZS3kmjR3MA
wO5YiXRyAU/cTR96J+uaQvDcNNy42LR8+aadPsnSKfK4G0ZYzncRlLQ0dJW7HeoTVg9kOYYNo+Ym
8bEj981QS/M0fSpXBOgMzk+/9Ozq5id4SCJQMUk3UKS3fGU83SMMOmlBNXd+Fml41qOZfrEZnzkf
s6sifik4DBW62v5V1u68c9/fOeGuWPeyKO9r4HmN84qGzg4R6pDech1JvN6Abl81U/z8p/BcSmGT
aR2WOHF3N8eJLNn8UKXZR5PPElWQTYGPn8Qv11JRTT3hf6uK/s+W+Fe+pTcey3mYwS6yDKKdH6id
jIv0CYYjSYbsO/ujFP6vtCwGjVxO+BnNHkfsHq28ttNzgvw7mJbI4GpK2yN0VDLM4DlgYrc/r/nh
nFLTJYMzBbd9WVGzPYLSodZBZNtuQlCIln32yOLZHfCMRI++2LHjTY5AEnHGjuXHb74gzstxjvAq
pxBe3KWm6CcnHzUHx/g0pSQ5Qu3eSyfdPdcLz5dI51sQpPo9OIngltHKK39Z8YSnONKUiCQnqCzj
pemWhb+mnTflRIfRaQ6CkGTs5C9PouXqaa+ePKwNRBlelf3aIQvjzgSLWdSzWa/+dqDbPb43/VUZ
AEUp7WGjO174cqxbnTb9SBP+v4tBhSJTca5RBKN/6p7pBvUbR5+qXSQU+QiodfRwreQorBJP5v+E
75AhIxuw7kB5fgAsQ1MemYBd8845hq5equ4G6ACvbX+ilMqo1RF5C8esRVdUf1Y0AooejycMAoPC
URPH/R36emGOLNdItL/MxzdO8U9wcRDaifOgTWFizgn0sPDadRcJrdG+IfOb27HgHUvM9ZfkvUsT
tKpZLgQBcOPVwbk/9uFpCyUp1yeX4STOgMk/Mxc3f27zVohV+uTc6eWL8BHAUiT5ZzXwNIkKE4mO
0LCiLWJGJF1M31+LbcT4II+o9fhW3mdHV86OA7+GUnZH0AzQzoyI8KsI2y8fJZIm1v4N+NgIH2bc
1oZ7OVis3UHpM14walr/E6Qanxm34uWujFaNYXKewGZSloIgtbwcCFx2semC6yZW6R7bt9KHeNXy
SJuYZYNouDBjw40hwlx/DEjLsOg/KbCopf3vDRy//nVTUI1ArUmvjJJh8wnDwt0gm7rTDsa6x3q7
4n6wh4IPEWNSWdOPsbc4u8CkRsSawhNWRRfGIpUVYKAr9Ol04zwC73z8d5jECVP32kBP4k+Jj8KV
5wDe+1Q7vfCGU2fx1SZEpFvBo95ncZ/TlrPDE7SMlIqEBlH1cOlkPS+c2kkS6vubIWPqEnf2H/GW
s2OSwdniPVSleOxMWAjfFmIATeM9+cmih7fUV894fkfbfURL7FKMxK+L2TigD2Ra5nZP+W2fAH9M
VYr5qhd5MgorTWT/FrajBJ6MqXtmIBTSWDJm9E+nvZ0E8T1IaDwdlz23rYlOg6kuS0DJ/4cCcb/i
bEIPqSHDSa3mJZ73lls67M+VFVtgi2MH6Er76FBBG5eh13VsMkeVd4t/HF66dXPujelp8a0T0HgS
qJW0L56VsL8Eq62UVqEKKHiFvUC3jGXP8MM3Q1QVbhwCDQVR3OoiwkR4npQF4UZBvPeFj50pcToG
Y1g4B7B47PEmqHzol8rXCoXO62oA43zoNhXf6b0sOdtUtv17/zncSnjbuI04QV4BjAuskvmLpGpN
tvRyX4Fgqsr7gs3RLq5qhKP5ynx351pD3+5eG8scX4PKxydQ06M40S6gwPEbCddTqME/nSzTFQ98
KQVwIgatpaq9FCZNjluRrX0AoCjEUWFPadi46WjLNsz5LsgnMk4pGq90PiF/dSJYJNqKhSjw9OaZ
JZJ9/oBgrBG3z0Xrtsud6lpp5kIRDTBd7OqOAlzQypn2GGj2DisQFbzZCdUAVgi3FGyhqjFMSiVL
kraPUPebRK4JzaELPNJpWJ5OabgQ9K56f5btii2Td9eVJ4RcvEA+A1FUEiPJxsH/Y0lqD1SJt9Z4
7bWiK/qirWaD9QZK8fKPwgyWPPT+wjXMEhAmRqC4sE2DdieSkn0dcVbgDF/K9dFOix/z+q2DQqPU
uBjZ1wyGLwweOaKW+2BAw7bysfKU+oyMWyz/TNCR+LYP+q+UXIq4P6G/q70ukrHo5CONaFzUCXVN
Bt9CahjbJstSehpHUeFk11u8delaBukgTnPQq8/Zh5huHmRb46ju5520OCajppmlXPXLv4A4mWef
h0P2Q1RSYYEYnkOq2kmqXyfcg7VP5N7ArkpZyug8ShKCLfle53hJANlrVXUOOJulHRdN2eAn2+4M
vHhUwHNaUGaSLqUqf16GcWMJpM8ON4ar1NzTxPO3deZ2kvZw4mn0loIIR6sbBODh+BIBbwZoNn2r
XwYrjNpCjmww+saTPzQ611waIXdnLHNC1KUcnS904PCYyW6nPcZlPkitV9Zhh6onWZlW9Qy5272Q
xl9sPN6WF3wjZaUCYJLtuyS2WGVG3emdKItNYqVxdAOJcMBFnembrhidT6gOpR7z4EglDqozBaj5
wgKINJ2LMx/3WpeY8CS1G6RDAMh4oVNFEo/qEo32wnbU0vKQ5eb99eYdguojOOPC68ExDMen1Kgn
37xwcnQQHhTlpy/Nn4Y+1MnavVc3E0W4ZAoSBSEkGjWjeaoV7gVdwBH82jBkuKf9k6jI56tiUJZ5
2xNFJ20+iLLsNYDIGFFpaMCw+wT+oHv8JHU2KXKpyMhvFYWwf8DAcsKvRj2xrkGdvlnoA6xQQZ63
0soCYQx/MxHKKg+ONxedBTbZ55NOaOAipvUFG99kI1x0vavLoL+6bgX5rBi19g1ekK0me/X5Fd7K
8VyzLFQTKPY04QMSU8CiCOCPw+6BdabFv/W9MOjF0C4jHl1cId3mO7nFK+Mv3anQGFaSrxvKv2Ww
kM83kdLrKyzdfQib9mpMmhzWnzsHboVRjjrtzJ5lKxAPt8kDR3sK9yNqH8eHMccLhEHVacQOViAe
wm+RlfmC0qkqMn4I2XGb8/Yrm1wnajS9FhFHuNVMH8Mbb+4o7Y7TWPs5Ohynm0IRW0NZTbDpnuaf
mIpKWBFlgj58/OgEL51hm8Pw0OyI+yBC+NoiIz1nlwyXCn6qlv90OV+uuCQ4Fc0FPzDwjbBjnwH0
ScRHy94L1IKVTZBDHBf1n83mk6ENLlCTpETs4CZXytLzUbXBg5xKYSeo1FIw0VxDx1nCxfzZPN0v
RqI25blKeM/+839n3oMHqEGufIEJOiLbZs/3Vbly4+lC5+6biLyE8HzhtuphsieZGDE2sLzKhw4k
x4/DzvTla6S1xQlZFRodykb+cIos0bW79lGSAeNv8cooeqNxlspV+an+zZeeTCrthwAbr9kU0jFb
BkGf//K0eL+ukineUMGcBNSHwZNg3vonx+HtaA8kPTu5RtsrplBkW8KUqzuIeB6Y3Uu9zKMMg4F1
b7Se/QhSr047bmUH1rdbqvwUEY4tVnR/rkLP86TC5mcVnLWN/2E9T7X3Fij5jO+RHpJF6pl6rkRa
O5+n87u6ksE3+9vkzcqfiE61cVAANrcTnM5qCJMRtoUXAkisXIpIfy87aoQSuHIajvQvTYpxd5fC
nF2H/+qWun/lC1whyYUaVtslIf7++aD7HnKtaXOKZY0IgjJKISZPOiIIoGG3Q6+PCLWSomal+uEU
oePmbwAga0Zm090UlrLJMSLoHD7e3T3XN20q/FAYUIsGbAxvxGKLfqBGzV7yw2qvqQPL1imFRWYZ
FK6XjeVvOJZn4MSZSFrHxvaxsDnaldeTwd72L3xcrP1Nlrpu3NOYVssky7dWuW7ins456yHn93AO
t57eyNyyIDSrpCoDNpMxCH4yKsQpoFJQ4KcP+r17VH9bbo/46OC2pQx2tCqmmk9aNloaCg2qU9bR
QLkZhnGdXOjiGCihpLhXdUuszzyfC0wbBDtnXcQw4afwPSW6o5MIwFmjWxpXJYNGpl0rFS4oJw+b
Octvs7tj8SnprbpTMfs7QpZAHlm11Hx4M9Vt4XWE1zJmIKdd44AZqFu3MfbZ08ZaOMP1RauhfW1w
ePOIt7iM9T5uyRbD6fFS1f9k6vvjesQi731vp93rVe3k4zuaJOXDYEVapvsefqqoA0s3HviDD/Ce
xzjRLNR1P0tpAMfDIWyix2NkjD+z/d/a2t9I9PE1MJvWj01cRjIDfH2HZ6Q8OEtgE+6Y8ztv83E8
sw8d27YPeUFNtaT+wf8AQTySt3hia1T0egMOAxgXE43xwxbitkw/zymw8ELrVyah1Ela/4iwDLTT
66m2mWMhMAZJL3XQtOdwghKv3xjabB9iSr6tucPyfdXe9jsbvHuMsh7qvUTJWIPEDEhen0A5GyUb
LgvjQz8Suc5EPs6Zf9oVJmwmKdmnqxcWT74t+0OZw4y8ETy03Ppmt+NDBpbCEFoARd65HzoHygb5
UaeCoDKNe5kDlzZhMaPnv0GqccY7273q7lNveFl5uPEy4VIBaDZGTqAfspLXqNZaeg8tqzVAVK8R
3ofmALx9e1gpFSSUdGqRjedHpgJ1WmuHXSuC1aXHqDHzcaAkTzqEzSJxU/Ed+clvJFhnCbqXOgW8
aSpCJozx+2Vh409szIpGl4pkVYaTEt4LLU+Ljj+rTwFGf+M51HDRjF3bGIbytAi9mXF4L5np6nej
uc1F2S38v6ALvG7yXvWKlVHP2G3LYlbR7glQYumrOYNmSDFvKOmZ8mvWWdjf9ZarKwdzXyhNIBmz
voc8MGcev46FncJgApLOwqcpbb1rPLMXmDRX1ZGg65AdFKGTV1G6tzOpULM88HBxgLamY6lEKg3H
EkIzESZYts8PGlFJzs3pbe5vc49h1/hCgxcmLHwXd8o90LrYL3U8DgMNMqGgM7xlq6HL5F47FOaE
3PtFyTnCUCR30iqKy7cezWWLoMxVwJFHGwOTaX8pgTQTE+1xO4jaJg2PqQcOJRDuHBwP9tQH7Tm0
srya9ncFdZ3Atoye75GL0dRpDH+/qhlOktJtlFiXP/mDs7vGEaZWXzt/jTWp+rwe4tx5f88XkQGC
b6unF/NTsi649F0LYb18rPxjclNRkBubx8vqxZTNSfkV9g1WiTzCzeELlVrETJEqnXPIY58pmLoK
YugY27qnJKJZYLfOKnY6zC6rPuJgL8o1fMmGA4OSvTISXnL0wnnM6uqh2H66z8asEeyyTrL5nP/V
p/SweIYVWzEOmTXK2SvaxflrLfxnS1/aa+XYhdDDMixBWB5Dn+pyuKd1gzXorM4uVP+nmEPQ6PGN
yo8eFcWRgxHkKcfmZ6JcUZ81vBasMlKGduLpwJIEtgePajqysRq9IUAkVaAxQv8AVHxESH/nGE49
IWZzPwpBhqpgDhvuGj/kAuVcJX1/iB+DlxryMi4mP6zkrvdnKBjp4MFwyfnuFH9ocmfDrMpv59v6
JSZ0pR04Bw8Yi8orwswexatcMPbPam9Xja/1S3zF+tFePx5AevgCbD/bqprAfjJicNMYB2UgW9VQ
QpIT4p9V3VRbdvEdaYkYUpaiXzdoL5UV9gN1smCn9t11+EOLhhd46dmxHj0ubHczFFYjHXgoSQoA
Qc+DnFBaSZgaMIVUVthmhWiC7eDadel1AWzoqJ6WTmNJF7epWAN/1La1WAoEtDNyWjATNFt2DR4T
y36oGGFfLj+7Il4SUvbRO5JOl9jGAe2YjRZMjUpvnDba398v3b7Rk7KbgR0+OFaCLJh0mJvIuWbI
HlDhkXYnwwxrphZo0tvRGLZdEKCQLcHFH9gLz5lNC3+LYPqOhyJcH2PIp46yqFC22B1aPvRADc/g
Vb1qKgQhmeptqs4N0vFh1X0dW1PQsyiCWEcfaFhDxCTtOg/W1Y+yjCrP2jb2knlalWZA91PaYXQ/
ba4DACl1mn2XORV0cFb3GJGTAKySzSZ7DqH5OOqoaPKr/QjL+m2rTM3PTGUml/Om0d2VDrhjC2SK
VVADDHRbrMpyd4DLTtpzUfaZwdAgc2Un372cIsZWNfYzNYwdj7m9LBuyhbbLfCOTr1nv7Z7QbqBX
h0VYKpl5ZouBE55RzGGRVMFSFRSWLY7d4v9ka2HLITkthtXQc1Z91alEqrGfaWdLIebgbg8CS+B9
x6lw/yYGn1KkhCj83Awdn1onTPVHoEkvy2TCB7R+j8rLMkREpdGIau8vx/47xjRpm3sHj838cQCw
nO9SZ8gR2k/wqY8/lumaIbM+dRPPAF7g28ggocWDURmdPpnAfdds+/7hwDRad2Ghg98JUTrqZKj4
3qwZVc4LLnG3ebdRH+IRx1oPoScRjpEdxecCV78a3rOcGff47o94d73F2W2MvrVEzbpoIYnsfFwh
SDwZ0wTT8EJMsmnlMXZ9DyExRXLEMT2D2WP5y8rzdvHMmLsNNjKWf93WdOW4WldGIctPPadJlLXb
s2uha/aRjqcsaK4ZlW7y+oNfqJ3jvaL6QeStBh/Q+7HhLQRpRTU+7ULH7oCfu1PRX4nWdntlwkM8
sx3EJm7W7wEn0RKQrZwVQT43Z9ZFVqB+XHA+OEaifaIyOaDzq96r6fnfoYKOD++dRsKEq1Fm+pPb
y/3SB8pPrI/fTVHoFIn9BPeJImXIvlD4FU2GFkONxet3PaMYp5DsSEGeVkTXFM7/PeydiJmOxZUl
BDMX60G4UXyCXwwC6BhXduC+FsSwXM9umo6aGIc73xrwW2MB3WZOTj0lyybYJZ/ZiKTKNkuXh1N6
r90ocdd+ItnQyaLFd/gz6P9u+xIR5oU0zl6XB2XHsmfK+40WEvRvSWXdjCS5b8zscG8ijAx/Rkn7
JUlpG8Fn1XTNADtn6sjqldCF+Z48xaWxpBLwKBgEnXGFrIO7PKRdoR76e4NmSSodQYMKcLm1SN5C
VIRMb40q1UwHcG6QiNWWFA0ijbl9XljZzThR/aLxs7UA0i4+hMjefueORywIunstUx0P5N3SoBtf
Z3WMehuyZw9BpOgB1P2fYb2UtObNp4gC8QW02CUvjm6xE3VTnYjr1EmcmwEHn+Q/7s2Wp5YOBaoM
LCKprxqsbaVZ2YFhxTdFhNz1T/OfkxJ7ltNZNC95PZGlEVAaMu/W0eDxBQGUv3lY6FA4gsn94YgO
34p9t7DPlOXfheqWjrKI7PpFQRxOzv2M6azP6IJCgip9t8nrCivGxm/xeE6IWzVFlzglf/EJ5pMX
xi2f/NsfVfWCLkCBREleG6nzwEDFrTAmI3Hn/0/wmX39xZjHfkim1mG0Gw9G4apzBb/2yaErScCE
l2DrSsLYHqBalDGOYZn10UEYCw9hnqvz+8RRcjCVFRoDyhKFu2jjHllivbnrsK8IkeMe1Il6g5p4
zrTuDFfd5xSuWvdj982K199rpxxUDV/hpP/D/hF4FTDtG5qun1gaU5Jb+uE5GBVXSukqmF19I7g8
/NpApsVbIjZSWP4N8N+0IyVZS/W18CEgvsFWzvnODtqI2mVwngAM4+W+oCKsvw33bx+r+ez14/dm
0ABWnzFqKl/77RzC79r9E6MimN9Uhjl7NK/ep9qcqu6h9qH3+Ab7ib4pqM2Fs4jf0iA/1pP5abyG
WV/idwOMqecOjxD2fYRXyfQhscnNDBAABpJde7Gj94q/98gJSIp2MWCtkjWoXqmtyo76xNbVpOQa
qqLcaxjz/V97NsaKI0FS9EeFHh0ji0cWW77V2LmR/dl2RTLu1ca8VEC8CQy/RxSyafE1WoUPR7no
pJqt4zuO/8H2L772EAvd33mmxOyPFUdbwymeHnfFpdt8Z7pTOpAEmE82qh2lL07oanNaAyoxko24
1dq9ruDDMKy/vlzWl8e1VAmmkMuNdm3YxODtoQGVs8mfm57N55iCLuFed9UvGTwiGyvAgctksiio
fWdEJEp3hBtcX982Fd3DIZwex8e3UYKeMhHJNrGk3gh7Tha1u1zXSyuOY8eCiu+fulJ3xoJYtWNm
sZ9QGFUb3FNJAEiCM5HRlzbd34PBXP090fi2zLWyobImgt2Md7G/2k0sHlvL1wYidny8s8+lg5KZ
Eq6Fw3yV3jz9beqL7olHU6D109RZDHUwHtpfvzk+esFhOD5d5kiJdZ5rGpdMoALZs2jpwCQgbKIf
FgLJS3rwi1VgbQgqD1xTn6d3YxvU7kXRxfh12BHKFuZramQLnO/dVZ3Bwuh1RheBEa+VNI5jrgE/
Rs94Rs382kLMNUYawtjV+zP1khpzIkA01h4k2j74wKx29fM5gbZGuN3v0C7t6Hw87gz16qYEhdsm
K/p5FiW01x9nkAIfXOWSNiJq3y0Bpknj3iUoOON8kADhSvIDMGkTaisyblwlrQFXdLYZHrTeme1Q
fxFhDCRUpPrnm1NjBodgvSKtL7TprJStJ+ZmVRyqCqfADvV4MkJRMEdz3VfpQVm7Ub25ySi53AnF
AZj9mxHkR2rjKgMPlIxt9JrVLAQJmVKYoBNPsksw5sgqI59zYqDjhDACAUz7CCvpPIYUbb6ClT3Q
ghv8A8d4D3xm8dkyUxESbktJanbP4RLkIC1a2t560UZ6N8TlKacWGg8zX4OEBimn78ZEYU+ENKil
WbX9Db3qqgKgIQRj21tGK8woDBWPuYlq9RMihQlCKuMAtUyDQgpMe35dWSzupuHYhLRSYbzb2ACB
2X0fpZ7kMEOMoBugwDPCMIERdhDpTWtuNnij9x17DOX46PAKvd64Mc8pHFr+ZyrNriDgnqr0hdbD
gWOzgSNFuCPoS4dedib1FdUf6Cp9bulmsSi0q4C1pVXesrPkCkj40qqoLK8tUcIbS7ueA7lVc+xt
w00ba+dzb0DNjT1jBKjYtoHw64UlTo/p663ehQZIoXI1SSJcyZRhz3sbQ0Re/jyka1VERNUpMfIk
LhkxkxMZ8kL3/AlZ1zAu2rHOC+/WkFLtJUJUO0ss8OIZIyehtfj9iIk3KfgvfjXDjxIgV6Nf3YaS
rkKsaRkVIWcWI99JEOKqFoZ/wXrn7a3Sz9j3VxMv/nwLthk1LaoiYbQoPVAD/Yb1TiXA1bWtjKBd
oa403mknubrO/4mdFB9vhzUTIuSHHy+LBCcoE/JzCsIFanTlXhdF+J9CjHG9cucN8GU0SD4r5Q4P
RhUKYcR6bhI3BLNVT8CYSJLX4AitqJvuVhb3MPI1OkhMtcSIyIbgNRfjSdINXbiQAXHgEpLcZhwB
T4wi5I3a13j2SmEKQrihJ247ZA0hSbMJGCwyP/+pD9aOMKS1BSrGNv+WdO/wngwcD0pgoBPH1Ij0
GgQUdrjZtiGuJn81vgPkMxcoAS5p/+oUrDOtTttFl2XwQBiJu4hIlxtCt7CIDwOTox5CqOC0J8b5
eLhtGdWUcVh8wb95LPDXwW3QtrjbczPkKXFOxE8KTgedQelaHJRxdkV1Vp9nKsdVoyffazwMo1gZ
w9S2iaZ3v/VwEuocISjcZKcsqrEyT147+JRvWdz0CSdW4FCMVIqx6eTCbu26kZNj28flgYRusaDb
xflA33as/TK1uerdBN8KzlcgaK6VBvkgMu/oZ5RiUsU6K86/2tADj85QjnRVWuOGRVxIt7a6LgJp
E7m9qxGEtacNqeZlnSAdSOlGAwcdpP67c26bDRbyiZkWtfzrCu0p7Qz+WXnsVPpH7Wrbr2d+fzG3
slzpfvZindoCji8vG/EfoLA6YiCLeI+Z5mRPp+tRc9gqXAVvOCokYYwI0GNHOWZ1+9Lmlzxu0yL+
Ax+p7FL1UFSvCpJuC0mlqF9AZyRUoKvuYlWOyo4xKI300VqLAe7mneXWhEj8Z3qeDKipDvTIUoa/
+m4e+X5dJ+zZFj+9oV2hCkAKeHDGXUv+AwfUp5mYI/n3J5w0tuplQDjsPvze3wvwRT1pJahSZOPv
49n24YuP9PffD10lwl6NS7IKZAfUoGIxM7M8B8OAhBcbOQk4iwAu5AZhkUQj5VNpC8L47MFt342M
bDX+YbcKFFg6z8zjtjN5YhvstcLNqBTbX6duaGawqjI4KfvTfO6XXsbB2RStoh4FJZcbLWuzTzkS
e934JFtPFZSzXdMJcf0W1UKl2Srw74hHkbxANXE9uBbfaI6iXAEQJED1sVmSazf/jK3PlXHqPoK1
yFe5MChIt8BF8RuSDXgaCglSk3dn6s/6Q6SrnHrom7tXFOiW/YT13fhODfCJ27xeFc0bHvdBFwUU
1X0SfwJKXGA9dRHPOnCnMlQhiqSrPCLG+7LnrNeYQvLdQ0V3pOC5eqeLLowY/7vTOr2g7aA6aFnO
khdwMLLmbTX+Tz39/oL3RvcVjgWRFErk7FDTrqKCirNftSEng2sbPv18AG9JhWiJfeuW2ktW1wDj
ahSo95ULDyTNDz16+09rgXfcfMU3qR9lChHeIGUCRyzGLWD7eP4uPDDTKPf0rIV5xNHt6z5GcA+H
O/HcIIfSSEnlULXTbhmqz7EcrY3LLTLHPiR9FP7pxAjLEeFLQatWmlMnI3vM/GmsSdL2NNwTETGH
vSq0j8/tqzGPBtT7vgotS0gFejVnU2uxK0NB6vAk52UnczHrCraNQrI0jY2Di/qI3Dy98vbhwBM6
HtopvG33o4lg/4Huj28TAoF8xfaj2KeITr4+E3RcLTXFWLxUndam6cL4S/R9UK/FkoQySJJI5HMa
w1CN8NF3S10QPk5FJQZCFMgLeqNcQvmzDwyl7hOep25bd6PLncc2ye4cCm6ZoFXkj0fCxoQGLxxU
MY2mIFe/Vg1hWJr444dTtE6v4uizo5mb/VoFLr8PM+wnyJAbb/1Qiiz72aUAKf1H94ksuL4oHnCl
WJ8H6RvBUe9k72yva/jV2kfffqcRxAWw9WxMotfJBbr1B0CngQDWSU3vFuFXyyWWAgWpTG7WtfDg
ufw7aeKXkTCDwiDezmUgudVQNlEHrwV/qEkRhL5+7XAAV4fkkDdMkZtGZ4z0SRXQaUhqI3viKomK
PmTFSOMNtq7WoXnDhbvSsqVUXCDuwVsa4jAjHJ6PU//rZlmAMI5fRXBt1oDp1nLzUPnbGObwExYz
Jfcc+Fd5MmSdWU3wXFT7HLdQp2VG9M9MIrZ1ZvUWP4TRPWHHhu+lIEnzFk6jIiob/TBVUCVa+EeH
t1kk/QFDjOcwz8enHG2BzcXv+B87ByiUohQg8sLHMXFEweEJoVSO4xMwDxKXwb3DP5hdfstTz8/w
P0aCHnjuD+fpIlgFxpdLozjXkkKAPyMt4PLEKzERMfDIeUHx1BtDuWc8bQIol+b4Zge90JkuMG+r
gefO6h2DyX0iJjZ7IzohLa4jSzFsRJI38V17Fk8Jd8rPtPuZNNhiqr7icGayaIH2aaPTdXZXtrXQ
JLWZ03QTzh4h9t6c6YRQ1P1JurR/kJq/2CdoGP0cuhRFs7OM0eHsfb9qHelNtiF2IVHex9PcQ95P
5TkwEJGjkLpSezRwwdaNCBD9gV5dGT9LMKsfokuyr45CCVOOZrRwEJpBVIzi3LWJ9gpHIn02OduW
2HReWm2u0uq6adVV60a3CGKrvR/h77QR0dBIE+D0FyyLoY+7ifJvOhSoHPzun2oD3KaJ/8EjQVnH
tYT7kwI+P0P9dVfAfhV6hqIYKFmQ6v80oPIq6BadNm+8fPa+hY8I4y6ubN7jZNDdxZT767lAmC+y
piS1PMMRileSM7dpjQnzj9PIV7Nn6ec2icG7TwSgHOvtnL0KSMzCUsXlZgc7YKaaoqva20AUgjTW
BbHAsxQZZtlJWaHN/foGHPiOr0R2kdQE90zvWH3sbFEFLV+KqjmdiNU0L2/z6t0oiwp1Vfz11/gB
ax/HGOI8EmXEm/2wzy/LP944UWVT0pIWbSmfB4P/jpwORMWJZXbF3OPY13v5YWoYaQ1L9d2xSkHw
UeXPfaUXw7DP+kqj1RpIDHs4R7porQpPRiWdfdSwil1VYToBnWGZDnpV5UcHF0SWGZLqJ7nHSE6q
LX7a5Gk4ur/nf4fJVL+Z5w7GSuChbsLBHP8zwU8wP/jb09dPvB6NHyfruIMcWgmL1EbQ6Lc5kne9
X4sNBUueLVvejGVmLQqzh4FnMHnvFqyVaJGPm13MGqPnUEOTB+5VVn2HbbjVDnAwpv7E4FP9m08I
6OZJKsI2Y2fZFZ/jBLOPJhpulZ+MhO0vbRtK/JwfprWW95MCDjJRRlO/WKghnrz4ZosgfQtPCOG3
nhHeRphsrQwXUcT/ow4zPJKNHDOESFoK4dghFzOff/uIkT81QAy+xXzvo8C3p585aF2Hbef8Z94x
8DXTK7vcjEvvvlWdGZVcGIdYwIOjygSW6aScI3vYXU4MEXPWI03MbLMXwOqLeJA030js86XMdXin
bZwgZX1n8EvSynVl5xY31lgGOozr61V6lMmxM+/Du0Ite55HHe2dwMvANu5X/6KB46PIcyWOrZwM
rEezHX19Olq/kWomWhxzV0pn6IJN1fU4i/TZKOBwIgvjulC2PN/fyKHp4WO2b4EzjUI8XNGJ+FeM
6dxKr7PmT/pBy8Zv6zNa9WNRjbzdoxhnE1CUILz/y26j+MbREPqpFcc9c97jnmKAZW6u+1EcCmwH
GerTv+3jT3su8gDoRE5lg2RrdoO88O1RjTjcaBToa/c2yM4VJc2qXUE9PiB1sdnpg7WNZl3kjDMo
37qLkR3z7tWBkh/oXwd07n3eDfIbxLEppqXGF7OcLqtf5QdOpJ3kYb+dV94mYfskBkThaSzU+5d6
FoEeLJ3Um3DAN0R6TqYG0wYFMLsPvKL9IDjAa7SH/H8nB5skwWjxo5J+qE0ODTqWvL90NOx7VLXg
HMqetN3/qe4jktZpWXdqZpboxnNSdEpxtYHk+1Y7QchtrU9IfJzdKJs2qpe8pcJQZ/D8IqTIdbeh
yOa/TkWggrCtYmFPU5LmMPTw2+ANk+qTYjmF+dYFEs/akrFfKPZ57QqGR5x1jLpZdskzc3kSR/9m
ctedT7dMKvwBV35ViQyYDCOh+LcV8wFBr+IiEeUPvjARU/hc86zxPbNAhmCP7eyCme+xAhWL9l41
tOIgd2vqc1H4L7VP0YYszFQZYbO4I1BXrPA+xF5M+ohC/DZRd7XAMYY3nYkbHgWXpMeuZIKtcBHh
NbO5SxR2Dc9Wuet44PXH3Qu6Udo6v9SvY1EZfJvndfkSLJ6pdwTbgdNXsAdhG1nbUpI9T68HND6I
VCbQDrv1bueVqqyVcyWNfo4aa8L4zEcXt76jxO0l8cpov4D353eCiLYdsmdRO9ppNVFUX6B2Pt/c
0Vo7qKNP/ZmbyQ6MMCrwZ9E//ENngQXZXlvq7wkzP0+udU3Wq5V2Pw0th9aYrcPb+0QR2l0hFooI
j7UB7YJllR24LCv1vO7Ips536QvKnBrTUJtIrcIFolG1/tPrAcwZG4JURucA/eHq/9TwkAxLDRJl
FXsUC68pMdOHAgsvXiZxAasyTgBCFjqMuH3u0yGz0AO9SKo0k09NyVfJHSD7A9vDOV/QL7qWi20J
7vRJEBMo3ssfbMjlbEm4yoKlDgguFxj+DGrB3KrJaXYt9lOgKNJtUviaJP7sdnUOXKvtDm+WCy2O
U0UF+a2xSFWt14HbAujOjFTjHQB+9w7ShTkWp4bGiWyHPZ7OEJ5GF87EF3CJvEMZwcL7CDumZbYX
0OZ0w2/TOvTxZpAiNGw+dRtDjiXFX7kLj9dBI0jl0TKcRDuxk95t/pdtG1zL/soRyG+VoLfh4K06
aWLLEjcxbTBHa7AcIwu4ekXny057huRDcA1c42e+r8U2w/fcLWl0K7GuhBLIGossfx11xqyj1FHU
HP05Ohu1kSstJ2dfMrDDsGzIzgZI/uwT5x3r0Y/ooZo+FUID373ThZVi1a15fJmtIPClhIIVSIkn
u0HL9T0Wa39vxtbGxd/j0m0sVElQ9sPKEGm4YjleCVEFjxI2X/bg4903B8uKt36pX4lYKy1B/Rux
Aiowugj0WdIn2eDR0HwBIS2gLH2WEcrwMTRd4I4tu59KSBYxxBW10S8bPqaYPaARM8ZBh1HBtHGH
IMEV56W0BN3XHKiSq+PXItn6TI9QlsPAiqoGwwuTWQtd/9mA8qKUhoiIWWU3di7N5e5V6gtI/MaB
jhJOyo37ScWfIegLQeq4thnISeD7yIH4u0HN3pCKkYj+/QS47W3V26EhCvR9OkHp9IyoAwb9XYzs
nvbnZvY1ewzZoQy3OF+LYzp1rWsEeazOt5PQCJjWHJLCLTq2s1Bw9JjFhIrJH6BGyphkrE4zrIlc
biTc/F4owE7Mw3mTmYu9qBDr/FsfZFPHj37/P0FJZ8ZLOa2j2QJr8xG0OqcGzS06WfhSF8q0o83k
ZTU/vgzV70iZKeU7w397+tTXNBHWpurlHw6MOnDLcxg5lq15aMN40SqFuczPNZtif14TzuASacdI
XQIJzhccBwXDFXwmFXJGdbS/nzC+3nkJjCqRMymObKjwgdmfkMA+jkD2kMglAIXb+/KglwhUd6q+
qN2onGJ0WhhTsA9odPTw86UaU1hyM3XjGno0xFn7hu3i/ZIhOjzD/cc4s3OhfKB/9AyCQcuNtoBL
0K6E0vogPFq5OKQsLcg6monkNEIO7mo6Tu0srCC866xwioi2D0uET19B8tJD9iVmUJp6/lICEDGu
Tn0u2Ny709pNN9a3ZRJN8etDiV7r8bGT88HRPE8rMG4h656TT7hz/e/mmqce9cRip0z/HC2Kaczh
fO5aO5hGM8NyLKIQYEkU2+/rzuPiZU2GTGZMSSEeQqQm/3JngZM8Y2tDdX8oHYkE5dQf1QIX7iVW
ENMOjsITpxeHBAmTlQkBNt8LIeWnmXAcrStayGCzGjrfbEYXDy1d2gtLBnw4bSeJpL5rk4EtRH6t
mqob3ZU5E45NEgrXYHrSdBfthd44vkW0JyqHhmn10JQg6wfbH/uxY1apgBjeRm3fbVp5ES5j0wbi
yVjR6+AMAtzegIPweWtzbVgIboz0/e/uTUiI8uWZMUIeuiMyDATsTMKSMcJGjJvWdkXFlF8JU1/7
7dt2PtQ6W28USx6jlhsucSClxCYE4DD4lBx8ZX+YBYx9xVICrTKlzC6cvzgI6utCEcmrxLEhemnu
l5iirFSbYuTCq90LHdcrsVct7hQpImhNMYYnEtkRvT5PSE/uHXBnXof/e0ZYJZYAA3xJDwBIzs8I
XFcNGEtWKej9cEIDaIjeDRH9qloiA8euKoqo8zk8FW02Tg1hiWQdPoS7fa4Dmeb1eycUnesAMdlI
P6UqGXfxXrvoayq2IReOWqon7DlEmed+bla1wfQErMT6m6Aip8YGpLZDZGd3do+Asi+fgw1iJs04
JKw2saPO6muTmwVSrPZzi53HShuRGrEnQov3VMlX/5LXxkcvHrRuOJNZ9y5OR+D9vWFnBlinGZgG
I3lDhI8nt6aBbLk15fHBXEG+JMAYh30A9GKXh6UgUsyD5YaA6WujZrRJEbobvLOWDBXBykLLbnfT
/IUYVSpwew/mmZ/r0xjbh2eig7xAyol7el9V94xX4ADUj1l3Lck9Z61UvtET/benYf0CNVfsk3TY
whvGhwuGfY+YmX/fys92uQWLBlrNo7p615X2VnkbTLXjKpYzwmtS1+6omuRNtg42riWKPhQ/o+CJ
Ro/mSMpON0YKz2Y6pu9PrO9NQpZIG0bWD48vuk/lEOViBPvWqNR83O6nfEoFqi4An4VF0C1Gon3f
RYAq0YDSbvpuHs6wvbeARj3yCmO2SmqmgzxJybilD/BYSookUGyvFt/cI1Ye7JO2KVF//FCjkRBF
R04xGH19iciC/eD+X/8ISwEd+pfIfQ4Z75hbMOl2ydfRhuDz2uhRW6v/vD6Bie1MKfLburGzx8zI
Dvw7ueOGJywqs40ujcwU4QdTc75LVoD+jePyo51BRqNTSVn4sz+HI1Lx80ITYvn+U1IWORG7jasR
fLh5aaDtldOEe1lxq89K9bSoxLn+qgjKiqy5J+A8HGvdWnFf0npvBsNdJQ5n9fX2NL7PEm1ZvYhf
fy+YKb1OvAk1xSAFOOMhZ5wFZhlnDhwPpWk35wri0QrVgVmMBMotG5z5hlqTBr13YC2pS4TbPnzH
GOotsdRbgykyJDP9UaIjjfdfyGPELbBFEE+8Fb/jgFZOTX00PMrgWux+GkKYO1N46M20mAbv81i2
4U9D0E4pAF9NjoTkNvQuyekEWNxxiO7UOOS9pgoi62Urdk/CaTLTIDnmweAV9Z3nCNqzmfnHlu5g
0b44duXpv47/9XPu4RzmphIq/g+jBXf/SN79dbmy48Ud76fIDU7M59782IZpwOz/8BfLw/rr1/GC
XvwiiszkCqQsH5CCIkIEoBlbnDYqlgH/BkAbK6O4M0ipJJTiIxrFi8CAHLy0wNsrftDKgcHPCjdW
ea+29crjkRSAt4SZrZIGeXdPFQOdH+NOibRownbX1//h+7gzKpcrT+MGkvzCnaABBJbknHI90T2G
eR65vwQHUR2hRelq7tzXpXjcUD8uZk7l65P6rAh/XHuiwUmQeGVeWmPdsJ/vX6BsWxQR3P8dQqNm
9d9eqnFRItUuXOkE69B0E7DlMsBD4l2SiIaLv1YeuZBXjGg6bV7/18ZlXkkBDqLhzwlrfAlMYTKk
NRWYyF7F723rLpv18q1G6aOM3OGL+9gv2D+YR6n9jMZ0CkiA4UEHU1SENJqUQ9woL9rNxHQtdjxA
20Zz4L71KixAKyF2eSuwdWVk6EcMoZgkfLva8Jrs1Abhn2UyolmexKItw8ozwrCAbTPlbWCZJC5W
tPuqMq+SQjwTZPCWnHLVkGufe9pwOZzANqw0sYSgFCeaPOTO/pqX3jbw8Pan7YKHYSlsvevftf1s
150gUrpVEShmlX1eV2/NRdE/PbZe/OuOBcyD3vHlqCAkAqBmVS41dHj8VLNB99GAPAOM9moRAV8E
SWyvp/NHMWawiP1K2OlUzYxqDjeT37Aru7shoSxpClB6SgibOyo9nT2LORu6Tkm3194H8GDi7dXc
0a+I0L3BX/u8homTutCEkT/0dIrBIepPdOF7uIuR7cq7RI7VQMxhAT+JQW/734v0AhOPSDB4CHUN
UaPdSfOzzEcOJX+fbTrLCdKQkr8MHwbkQWcQeCpHH7Bvpi9agm3SnzfOTSpIWIX2IQlMh9B20QLu
RFBiur2JWd8uPdNX20rPvgSMJunCL8XRSapucCRib/brIOix93d/z08uojjiMmO9AJpHTN23vuko
KHHco+yQiRi8qMm5XFloMDytgSBhwPTSpLh3D77hX+pGb/+ZM5QqnBXWuh+Op+S8AHb0aTKr9mPi
xxhAaTknwQ8iG9KlltYBuqLKl/iu3EOpmoHu5C4oZ9n5bywzZNhnUsMdhBtFOBLEwzeEarGDlXi1
gUYP6OJj3YEw4ITk/HufjyVf9Bs6exA05CMn9I3q9pV4o0p8ayIDd7qg8/uJeAqggsCDxronP4kE
R2vUcXM6xKTgkSV6IQ2N78qvSGvRMjbbWQfWBBMND3mA4j+Xqlfzae/+Up0hRaQCA3VyiRk59A2T
gHBanxX/n86OtdfZuE48RPCT/8KWpLEiuvxC2t5q3zUDqUhKiK9pmwpV8jDRYzraYaWp9UeI/t2u
fPr1tWYe6L1n9Ec3yj3Ci3d8WHoo9pZ7pWb7Nd9qQaxGJB5PuRlYjWD4pG+lcBpADjvwVJYP7lT4
0OUueXTqG/pRpX1pz4zWrdLgzSe0mcHy3GiNC9+k8TDq/AV97jslqhoRv16N5rOBQ98Q66aDsZYh
5P4HH8qro6bFKcPfMyU8J9EkGxQgGKI974WkIcqkwabzC06UhghqWkc0sSkuzMLuusUXw6Hak6U4
5PQTrlCLTys2J32DVQGWnAT+Z7x9eTpmYUPAX/W+NaCExHE8+V+elnSdUI4QD/cnwXe2IZt70LYb
PmsGUB40heovvj2U+aK1tFVKJ/ORNqhLRD2+kYu38qwYUWwezU2YbYOKx3Bno9TRXyZorBopMZtD
dMWKhN+ojXaTvydIBwxOOA9BCtz39+j+OouaiG8H2Z9hdXcmpChEGJRvjd6RxfG+uusPtbcGgDmy
jyLGIVDUZQ1dp3Zvm57ADzWueso3QrjOezltuBDdnz2FERV1R4rBJFoAYfR1ZsEVYngn1Zj898v5
LzqkRkN0kLzKLeY25GitPU1ePSR+jsPyFDlLlHXnp4ThcU7XOmIJdYSyfllEXZmsfqHV4hlcuags
32XeGtHNkx7V246dizYKIW72wq74I4UK8HN6MV+EGCXfv17zY/DQXLyRMs4RcDr6WnOJfP5XP5jS
x80SQ0Sfek2nCZMqhBOqbeTLnzEuvA24jAsMNzmE6rfWzw/psCP9lefWe8JpYRbZe1c9qf0cQTOy
1hfmb8xcBrZZiMjeJL5H9xrD//gMjLwsKDjTMJ3x8diUnJx7swqX17ShNhEgIRlcD242YKFrEBke
8fCXqaE6X7NziPVXhhSPx6fsVjUZ8xYi5EhztIqMUswW5SYunIw9yBPOlzuaNfCPQtZTaZdpj0UR
1ztltyQh0NfacQ/BGrz02AP9TUm+knmyvrn4bprH0ZX1x5SjsajEzzejf7lPeF3KsH+0y0CH2Seg
/+ofEgj/jAAkjlU7jHm9pMbTdRcFAqLab5Urpkk+e+EgCHxxEWp0rt1Cm1PafprjJS985lDkyil3
+ZmAsmX1bA47Frg5JL2ATBbVTvUYqRXnASeUsYpdsDSbm5dik5s84Ebewu5V1H71pKqxeL7lInQI
o6Cu4ioGD5YKIkiJ/eymPWwoba4XXBolr+Jst1aUsNa9/g6qfgfMG0K6anv83yhek5z5JPW0on2Q
PdlQ203i7PaRbgjkZP8VCyTmEkRtbcWSS6fYpGYl7IyJ0KBPKD+Caj/qCfBpsHOeYviJ9rAbLdOL
f1OHXUS4vyNkL5bvv1SFzEIm/MZWRWv6HET3KW5yo73rNfabvLOuNoE8zpesJS5BmydXJLEbHrZ+
0KEJUlAi9Fl4wjrvnJ3cmXBi7kdkbBrklbfGjtE3BbRDlxeWIYxympy8cC0MxE4InXV74xotj/PA
8pwPtg3Yk059pzh+j9VUZ48rix+u9PX5hJNxVqkd3WMMM4GuEHhEdMCqFCtk3u62RdXBf6+kLfAs
JZULWaoZ68UsUNLDQLQGQ0JMLy3XPrQolAZD22Dda5fBlxv0TKJO/SXWiFhu2dG0JK5FzqwW2q2n
gKzfce4Iu01hHEkDcqwLuokPsGx0BFoU17cyhvPHNbkQUsmFRPXGuhAjkVdbgdLX0Us2HnZsoROH
MDfkpLaz8Ux1rUaQHDNjYrYZdwgk+OgOHxGlGAZt41EQLYVeOBIS7Y9PZUe2lL4oIZmf1KiDZiS8
H4uBU33kRY43tK+bYaOhijp/8yet3mT+AFUL/TQG6zz5nOkJp3FNnDOZbd7fEiqyGllpytEOMyie
JCLnkB3yQ/j2K3i1Y75hInuMuY4IiRO7b5tUt6Lx8wPZIwZHawrbJZy+x/22VZJzd0aoQL1lFG+j
1fJTXSA2fVJDuwmQQPkh49xA+XMgBIYG5q+t/whxqXITibgeZ3igw3E73wYW4aa4KWfyvgZ9jAap
j79ABozWcp+PXZFWWCYAAbsEOjJb0Hdfcz7+qzRGnffWL8QReP49rB8qhaov58UUeDHq20xAqege
3CkEnvJS7QyokWPoJgOHtZJMFhztlvxBn+1rZdceK8auz0Pb3lG0uqiKajp2DZKei1Ta7WZtsWIJ
7a08oJAph0SXVzzGdCIo45To+etw6beh80So+H20kxsnf8J++FU66aQABYnhQxdItgVHOXe58/0Y
ZwtZkfNat1EbLrW2I1eA4epR65mm5pcndXiEWMxu/Spf5VJ1x8DjP7eMxIqNOem9BmA27rGAcNoz
K/H5+Miqt2b92m4Wo7zSdOAIudh85lbod62/fee5CtMvrkCHcKpoTICtzeFVnNO7JCh6kWxhBx/7
w958xMOu11MmAcjiGHyauWhQ2Tu0PUzKnoRsexj6rlQQ33+NZ+QXuzUjgoVE7fVDNXGk8+vKzXAH
7RtPU1Ti8A0m0p4C9c6xt1VC2B7fzjjuKAVpyk1mfAMBs6YkTNLp+XBJF5BIoz9kMkCMXcA8IF7w
Aev1xqFyAO6Frfi87KIv/UMY3t3LmEAIWDSL7TfzLzCNOsMGc5H4Bn72PcmUZUvITdNNoxA4tnsF
l0fe75kkw54gcdXI4XgdCUipWpoO8A0qbwY/XgxuUS+IrGa5BuhbRA2pnHpHeUQOx6asROowVBtM
zZ994C3anqFnPYA2PkuKkPX6kTRrP+MIGLAYg2bSbIs85pIDnf3d6R7v7LWIo16/2Gd8MJetRbm9
EfjO0E0EJ6fCe5CFWh2S9pg5I0Nzfpm9LNItLPUaJfaW6Wod2vZeUMolCdppkgWSCAq/vHgUZuVp
1r+wWF48Vux9AlPPCrisYmwlUa9s05Et2ZTUkUTpOyXy6gBE0VsLCqs6HJHkZ42A9OIp8RoR/kmE
3j/OLA08XwAgFjO6iBCI5DRXlepWrm24XEdBC8lFDXWZg9qZKU1BFZuCKkOZU9NSwXRZxc4Ibid1
XZZx8V9NTC24Y4FpVxtSYqFGpmlF7URDwqEr8ZzSxjveXWFJEebJZ/lwa8a002TWZMvrOD/dBugB
2daP+wSI/KS5MaApFOW/C5jWl4/D7YNhCk1LmrC48Q3tkaucQPVaxe8cYiJUupA9U/2uUIttuMGL
MrN5KO0LkbRNs55Oz2uPJbqrrZzSY9dTXnSqyqEiAs1Imid/mzOEUlMQsSrwRXHlbUFz3TCV+Ph6
tp4bcCrxLbxQlnbvqKaWY5RjxmktOEK9n1dlXBz6gO4laIM/HRqUWZkxsyi7AprG+DJ5U3HCdtNN
2sakzG5JDN1xryd/xrCrvF20EQGiHYDpc4SolH98GmFxdSrkCqFhAdqoAKsJvGWLtQzuMMUe2uO/
BbMBAY+b4UfWbwQhKo69psAtBDiqBpQGDOeflDW3QQ5gxhKGREkV4dOU89UXUMcHmGPeRHoXUjNn
W5zKdkehXDZ+4zWyaRkT8AQEpPzNrtSBuV8bKZTkK4QyzCRKnUEuk9MmRxh1ZvQ9DqiHmI4RFN2L
ctKgfRvPeSlwFtjFkh5A4llPyOT/YWYj3LJ4lDsHwCvvP+fw1+RjMIq0JH62azKo7ZIhC8xxe+BT
6/ppKe9u74+1Mg5z/ScHwTfdVmEQdECcRTFVXsQTz8YMltwYJ9t3FImktVXuB+2+h/Oof1N2HjiQ
y69VUgMBijsiRM37203ikiwIa1Y49xCRc+asS3lk9rR/fJ5sAHZViOYEhxxoYmLclEsQVQWgv0Hw
Vw+2nJJCDo8SZYtP7wc2pa6kspeUpyZBWLq50vyGDRblkohgBkTkX3L5fCKyoKK4jkAjCx28RLIr
G5iaBdCTRNc2/CHnvSbQOx/3mD5y07Lt7nxdvZMFS8cewan/XZc2K0TRMNQ4Uomr5huw5Gzj2ZTf
fbCPO4S10hfd81tXaPXLe7l/GfEe1TTKjHZl+kuuu1zOTA0MK2pIB/mU6+gdtNPLPgyc08rEzUr9
q3/iM46mBMhwnAywNB992OtrytEDtNVhGmWgFJKrwW0vNMNGbad12CDhMSjBXeeRr4d5/oD8+JHB
d/cVgZsnJK9U8oED6rwlbD5aicqiUaj04LxfrwFKYK8maOW81wZpGmPzn5ItmcJirMoAZ6wvqmQ8
U3mrNwhiLNkr8D76D/veBl7GLbzj/yCQzxTGm/TvZqv6+VLtPCkTOw9GVJoiFwGSAT0BddZZCp2s
adNRozOsApbEIj3v+6MrTz/95CtGVU9BM/YIpBZf2aIXDkQ07zuxOmVkR8D8uN6i1xRMFY4F9FkP
cpm4MyWdbZR9fUndaVW6dcl7XoDkiC6gCcACI+3GXI2zVHaaDZH7LOX4p6Xk1Z9nV83jf6UD+Vvp
x5tt5TFaqizEzsTk3RtprsqveLyHHmVgNIoJ7K/eRfqc1fy2wMdPMemweZJ765F1R7vnjwZBeiUC
6w6LxUR+YWXA837MnVESOuzKfbZGmM1yOov1UOdlKh+kYebNWSDjBRAZwD5YuupObeqXqD48GqA8
siuHXBHBQVWQxVkaL2813MZD5B8MIrYjS6I+xyoeA8mtwYlqEmGBWPc7ks13RfbVZih70FgwtdOx
d9TCqGTcCTuI/RAUhITN3ED0AC3iLJEy4ONPgZo3xl+JsC7U9o3a+Zd5JtVrevrBMISQB7fhiIvH
h6OZVXlgX1NS9cvXNMCuGqJLlkKxkxYqH6CfcdIDxoL9CkWYmtXQwjMM+idR1UPtTyHXheNa5Ssf
/kN12+CckAkDEJcqmyMzsCULgRs4P/kuFYJHp1xAUXDH4Hgqpx4jnAjornm0hCz44cKU4YoU1yRE
dxjH9Q5BSTy7RRtbX41kpm/lvRm4hpG2riqobUVMkDS4VhK24sQ+t8Jslr21+WRwLFpqwStN2OUd
UmdcvWPEqaawfRMQl9OOOwx8iwN76pOlwEm/KlxZPCuzd0tN1txOHbNUi+BKlot08c4Klv5VXiBH
hkRIrD2xBWsvqnfjiD5YTaNPwffmdv6eB6fqB4sUGl0F0jb9ZFkDflchjf7FdBo5EDwqZMFTKNjR
OfXO1bXHZojwrlQE5HjxZBli1hlrlGoeKw3aMkZo4tzQgEKU4qaFgT8Wy9Zo16JFQOKxVVFf7POV
CfJUz3DNDE5JFODA638uFnsGeJkjSfNkUFKY3JVeiSfalIofchGuzSSdBCf2tN2p3//aC45JqOP0
PWkgX5/oNRAE3zjpnBcR6QTwfQ0/fuq3iJR68vtkJTnSTu2Ah6tgYd1U6oPWY+cylGhyibcv4NqI
UZjFDNZa1Vp2fsAatQyVb4ExDxgp6yqJxCWvqAP5fODwpdnpDkFyc+nUArJfokp0CXJiZjMfsSgO
dUrvYM4PJVti30B8lMTKqNDQUk4JAqJY8lgR93xAGnm5d4R6ewO3UF18rU10kKfutw6NOpBrFsS8
lPbiZaQTh/mD/rFBRNT9AgjWTilQriUL90ltRtsU4nRUC7pQj+majpyYMfBjzWrRoP9W+VzROR7B
H/Ue34NaYf3rdk7wsAIaBP5luDk2+EjyMun6Xr1uIOMmjpXYrDlG3Kb8oodQVP5Vn2EgqXHAxeQ/
e35YhapaETcUO7PBpIjcLz96EJ1rfeATShGgwJd9W0QYJBVop4w0C0aByGwpeEYLwYgQca9vMWRE
0rHwrshySjaSpQF2iXgMxsVPFcimRVa0rG0trNrNOX2VITmaGwcir6x+02ibLsJIA1YSORhWIVNb
a02J2pwyNAjJSqwgAMrzCJyJCv8+wRVHTnFBesRFxQGB1tvPRDOAxUeFjab4fhiKtnRrHN8WJTII
1FoB6v+FDvM0n2Ktfz6yxJQpfJ40521nud+AXTo5QFELuKZ6xN///uPnHknd/hpVODHK0uGVQdhy
bvJ0RgE3auODJ1116uQ8VaKqdX8czmmTcjnmTiGbrST2cdshjiEIaONTvINWdrxUCoqbKOoqdwLX
nHQc8ahf8cNQWmTFoof0Oscuf5TLibRfb8C3wM8p9iQuAtSndb/V7K/ACBfczFkKEQvzFyQ0avLi
IbxcsowrJ6QuAFNW6yXF++TkLCiMXUiX/L53JitrmjOZKs0b8/UaBUJmZ4UosNA/8sgYsVDWdL9G
7/MStSSwcaVHcM3DFxNCWtAaYK2zBQ3bDy+TCHptdc88HkI25HmMtXgEKMLhzJtnk9RffoiyNRgS
PbFW+pnztAsf5K2/adQXu5Bl8DGvc+dZEIksAzN02uK/HzBbRQAkjGjDBLTnyzkPY0h9yrpy+Vry
aQnfgMiYXfmpsYgGn8oqjOpLe+jszsbiw397bMnVuXwqff17gt3bpZ+6P3nypMZ8FcORFY9svseT
/ZmMoE3b4H7MD765heLQ6AuP4dge7kTaD+Y0+0fSDXUQme5t7IYt6R/RWj/Zz9MJ0EFHYfR0DWmg
BKvXXVi0EYrlmgUbG0N+xhtSNEp3YnykEPdEgYq7orrlnlbO4ZOJRnQB8hV9BTAre4Ie9xaUN72z
kVKpgy8wEnYt2CIauoGB9GJL6iw5JLBWnBHWkcI72SoFotJ+1HIGbN++FvIY7JatTqlohLqj2axU
PxxZUwrLi3w4qiE8/PR+WsjMqDDhtQ6em5jEyVu9eLT0Fez/OQfMTG8NvwcGM0jOlXSwsMJK5AV2
inripfTFhnkJceBIHGMCFADB74Wslrdo4OdQpJZFNEBrtAyJMjOOEHk0Q4pm5lupzcdXDi0NAeC6
wI0k3SGCn3oIx8MWewnnZom6NSWelbpIiI874lLrhMydxyEjxt+AkASd9OViIU7FQQVRKr1KKK7B
wW6XGGbEiDbpSfthwhvStojEKBtVFnp0mIrdsi8R/WdHPqrSK+mAnxOidM5DOa4J9Z60njvj8HJJ
sag0dGyMcGn4eD/D/W+3xgFn9XoWWBvD1c3LlWUIdPzvZesG2HEEDH0T/HyP5a3GBqdYOAqgKjd1
84jKNrez/PIBB9ZnLiWiufpOk2AutevcxqzPviZGqpAQzVTqinbV3oogpiHvzOLSZnM5iJjzA9Zi
LzgU2nLqop4L+9I2UKCCtzgeNeyHAGbzPfQafeYL6keX1alv8uGJcaQXRIw/OTU40EZYE/6e5/l1
AsRNUyPrYq5OOZnUpjTdy4JNX9E5HpivNR6o86qb7Ha9xVFvyIGPgMymLk/p9XJLetT0i2dFanCz
7zKni+GtR4daImqvMZU/G7OWehC5y1iVmyfpKg0gWnwL+PCHNxXDkr9iU6ufdId7yzuwYBxgm7tu
518z1W/yyJ3NaFg73g1q9syhHnPDB6Ye2X7O2dPbMIFzZO3TP9bZql8iUGdx/oatml5hqTYrmdux
M6qhlpl9ZRaiTr3Bb3S1mTOLE0s05BGfiKLdLGSbxngfYx3EaQXGcfNcbc39TR9iJV2gLdP63Qau
zOiiHrjWoZVZ0h0qKd9Bh4xtJVRM1eV2bCZ7FcMJvzhsWqvW9+XDwPuEIgNHrSZePW69ykT+JlTS
jbGdZ2/N9Y6kyQfWPk8imMBcsgjS1pAW+bASjudK12Qg9Ay5rNdYr3OXufRXwHYX1zHbb80zfD0F
G2qg1OYDh5XmVJCQL49OAVorkIUHw+z3CRnxEYntQVc4ddI/IG9vQ4yHX06kmy/A71WCVippsSww
KMXlWmmImCPUiwjMZHweI3eVTey5fvlmMmykhuQyXHkUJAiy1iuUNI0gK3sZxPDR/zcHxvb8TrEA
aO7YyJmfMGUQPEv4r8fTPPruEuAHOnZ1teqA5xcvuHLMHXLKKe9DdJc5S12jLjFYdZ+cmuM/hMGJ
yCLTm90lrcB5ua+pRX1Xcz9HZA3+uRVSRHFemD3E8C3hqQz3SE+VjDCwrgmvuwTlF0FVSP0umrCl
c9yTXKIZ1ZKIJ6FxNxpZA+VXuEIAD/GwYjh2ezX1UCvqs4qWTQFvjAaVzreDLePkaxVkLCFibN3H
Zp60wPS4o20C4GQPVdf5Y69aPoidn0WRZeoY68hLL2kHPfP3dyXRyspgxErczHRkowXmLU5YzLfF
uGrB9qVX2MRPDrpOGzTHtJblExllDeiqTAy2vo4Drl4a4mX5H00DiKOVgDeNnNz5TZijgqPvHXG0
oG5S6c0gk+TUeiDBuXcf5mt8QsBdrTri1xn0t0IvZc1cOUeMWRlHrtJbuHofTKU7DgU+qQMxyKSo
xRMTfmu0zkGQMcMLnovxELpBbp7IzdaNnYYON+Teb4M9+6/F67JYHr8Z8FjUcDFOcOGgEC1k42nn
BDS8HPMfsfSodFFlaxTo/wqG+f/sAnb20bR1zwI1A6LGiqIbnnzrNgAxfTYL9fveMPG9dmQGGTE0
wUIzaDs4fIMJkzrr6xClfMJ473l2JPsEeiJKnX1+GpkYYpwVpYJ8ksMYK89K+84ZuduMF9Vtw0VW
KUmj54Q2hPqQUu/dzCrivVlocUFrt1ym9Or/Awia04hAB6W1Wz23LyTk7tBGOGyVih5gqvoOwis2
T886OTtEtwfST6S5Q64gKOm7DnpeIIeFqbMak05noCLBWcprQvHyblBcyYy8n13DCRyZmqZHwEXt
NHtjdWlGGXvxzca8yCxZyVs/frI/aXiRk4VdZxNxScfcq4KUpZSfWFz+xUzFJPaKqitswy4msPkE
HUdGvreO1h08NUPlrj/ht1TxN48vLo0GaYm7HF3DRoRg6Gkq5kMJRYFNQsmYb3yNQqosQSinjnu+
2LlmMVmzlj6hwK1RWCY/mATMtLN/+1PHD5wS9rqGjOXWgk9qBf74PAClagAeL8aMXrRxDyk6Qn6B
abHKomUZcoa5nv2JTS1ZKqsovq9nlK/Q9SC3HS91UDc/XVG6htf0CQg7OfBdBQoGQrjS/RY5+SaV
80kSkdky0IYvAzaqlJpNXr50XyfKVZ83Lb4Np27l1ieThlbiSnS3YMZKAuTkAmrmlF3MdBWbtY3M
2iRiP2Kp3ELx7yV9WOenDAUlL2MwFtf7Dy9/r5jT2A7Mq0Vc9oenhBUcB+c3DKsu7TgIZXLCQ5qa
golHRSFl9VSZP9A+vE8NAn7kNc/lTVe6r3F0GOH0BizBMmiBwwkp+teZaEDdwWNnj1LDbElqZKao
I1FCituZ22P0FzjSIuMmGwVRxhnv9IbOHWxKFfJtZwyD2o10Yfyfo3ha9iS+t4fQKkS0CbNnQp6K
iFSKPq+cTb4h21BuMRC/P+KhF3gI7uDqEz0iBQszFUJjqewfzIP0eWyRrkir+g6xCMfLa5KimDBK
YYjB4IPpCY/yqdrNAKnZDbiCiuFsgN+0bMuWll0DC8W8NIwAb/8ZGG3y28FWaEYrM7IADmqt2h/z
uOWYNl8XyALBmEJmXXqROz5sMJOvTgy04bOe4YIUsQutx8h58Oz6By1Fm0G2OIrpysfjpLP4RFY3
5Yq0Wyh7MQs+pVUSamNX7BAkGlyaRocOTICAjCvKolF0ntlKAELb95IjTfpBTbYwNAz7KpJffrqJ
fp1HCKjCtL9PctWzpvsiJAeKZ5Cybh7Eh9qfRiKgXuc2vvahkXFYNskO+wxtI4h02X0aj25MW14i
onSlnOGposzAUSBo1vOMbhedrBvmGIIjLYFhGSQrHlAy73fZC4wcw72j0bUbLjmJbA76GSdTYL+5
BZDAgI8gbBIuEU0efPg7ngyc9fa2g+cyFRdTPnvIcJwov4GINHJjOOndxXhg1AhKBadzWX1fHXF6
2yYdXpPMt2FtmMOExAkMvueBuk7eP9rA23bAfDwJg/FxFrVM6tlDQfJEt/p3zP+D3WQwZMpuO5NK
rXFWn/Gu/fnn15iZFtNVLWwfRxFICXXlxFOEcuZ2cLZhI4W6VfOCRXnfifjO8TbaoWI9WjBGR1bK
dOarAtLo0czMMKJBPxwWWVwlKiL1BHJP0CGgiwWF8j8MGy9xifFw1LO+yUOmAJsvfdAPMokKd3FM
eQ2egfCdoG1KkmYlubgDSaGyFliawF3oCMLwIA8uw49cmYHRHJV2FcH6XTtL0zV4hJfMutERPjVM
gPv2D+yJ/F5OF811tv4ykidHd3zHtF4Tbnr+jinlkClxCDTybxqNSdVoSgbgb0UMDQ5SpC12+Nml
3uG5kutwP2owxpjmAa7J5G7uzSHxXDR3DMT1qN6mTkMyklb9wjlVxVNVmJD5FsR94TlSIPREvC7t
8ONk4QgymoxcompCxkF+FnHNwHmn4SbOV/Hixc2z0TE9EyrEYIIL/Fq2h1s8Ie+FJMcD5zkSUG1x
PZLxtQmIiEMiWme/D6GeX8K8OU7+C+A/nSZwU3pvGcLZHkmpODGY+FwFz359qFueYZKD4Lp3sQ5U
ULcyJd3znl7HWX32IZcweYKthuMH2zxTwVW//CsrOlhS/RB0MdQoqUuUNmYxxoXhpe/jedmpG6e8
Wh2R88FQBBCi13C5X8l87q6jIeHKH6BgRFQqPFhP7aTrKHpClOFBG6NTYJ3066vInx8tPZC0k8P4
+DuxFe48BOggGPBtobOVwt7yf+dzerN1QmDlMbBGrBPLjJEfB70o84DEdOOXGvRCRI5qJuoxs6AB
J3Zw1IO7MhHr/+MXHsb/xPPQG/9DVe/A24/HeoJuCSpOrsde57GBwZjCEccOYKHcUwWYK/eEHKPe
hOy3NrqpXwe1GiKmWfICPSJ1p9a82cGZVHHnqZrrYT4SDkfjjECmu0X3sxGmDN95Rv6Pfbew7hKp
VAsQGsIMevcfLJnRRYa0pgCppRFUzzmAi0YOue0paP2j3eLTljp/5W+Hs5B2uH/a2uf9gr1ZsHFo
Sm532fFha22iHVtLKYbZqFqEB0Fy64IKSboLbGrVm77DaE569ONrY9ycKI+F8ts8N2nbB5xyTw/b
d6XHQdF/rh/ugDtfJJX5gr8pO+FgIvKICl18Ldz0+frnM/R1sVKTPipKHbWrlebM27hnujmSALFQ
jQmKNpnza2CJA35rY2/Jccd/62xKOWHzMVCL3LC0PPod3oDY40+ofWjy8lHUeSHiBwgjfrGRd/A1
VEcNeBRy9H5nmMbgw1jcCcMufEKrFpPpY/43kIztZtjro2MEu9MOa6wT76t8Y0ZvgDPN2LTUcAsk
O24gHb6QDh/TIZyiknmzhAsc+ANn9UcQxfGQJaPh5XiiKVmAl9tPoxQ8GuzOBtwszl/lP7Rilj46
VSWGpt90ZgXuddnd39QEyutg6x5ntgKezdQfy4Gk+PT/Q1eVLTR8OPOKsaPJbM4yIsIj3F+FK8Sn
XCZBcPioARDePjjAnDBx9AaABmczli6hzzvtYlJvR7iOo6om1wxtnM87symi0s+Qr2Hqxo+SWnt1
dGT4wVe1YZmhu9leF/kbWEzDa/mxdn2AsJdmRUuFXiJ14gicQYq4pLP7CZ/IA8AMq7fVdVZ/G0+I
zK7d2D+YAMLIfPNwI/gRLozJ9gCx1WMd31F0CbtMtsUUJN8IZ3sGfiawpYXbAWv0t6elr55fgWS+
VaB3mTv1gKdBQZn/nqBDBefJd7RgCgi6q2RZrPTUvHZJzbFN1aam896kS8z72xx2Rw2+k4L/T3mY
Ucdhk+OtmCHdu1Z9GBveiEdNZWgEJ/uu3BgGLgdwcfOfV2EpFnpiwiR2tp40xAXvxxRatR8PfbJA
WxJUlyIzQDt4/MGEsY2bP/qagv8mk9DOUYku1q8QPyBfkrv7VM4IxeBESZXvq5P2faj1YGx3iapV
JPyhOLd6xt8xorLhVZdxoB6Ztr4OAmxylW2PMz4nMileU9sFNNdU28f7+d1+xwDoLYeSi5R2L70R
O1NLXwJXFjG3fH4n0qOD8RhB/IGwdIcmMzECfYSPwn3tCWrylyqtF6VmaWOCkaeIlW/zdWxksiq9
RJoecNPkhRaPSGvWhZS6xZZNoyIhulS/DIW9cclLk1kUYQTbT8UZhAWBfbq/J4PtH3v902+4hPix
95JV3dOowLodaHkfr2Ox9slHUvzN3E/IDuhR6NrheSxsJRXQviKf0SZ1QFQu4fnwrlBBAhDoHz7Z
S7xEeW4ETly7Y8Y95R9l+WvlQ5OvHb3TamkVhLsYsRzkStFthw7tL4AoGYCzeZyUKgDCbM09S8XQ
dtHxjOCe22EJ/OJ5fOSRXVZpR3cpRui+5iMwfj+VSjkpCu8Zgi1LYrjbFtUpZZQYsF8t38rKwFlN
7xfD4oR3DsGZA1zI9QzBIZp4GyXQ2xmNRRbjPk4cHZhDmVuMahRq4AEVOot75wc9nuXRGqScaMxW
TodXVJYtmDKgOjBFy97rbUGFQHgZgyjg4GMiIXl3x3qMgINMaTOxyAXbWXF9CVdbU2aKQ48II5PE
cZ85yjUQr92q2I7ih4H0DgDJeaD1oSkqdFPu8K6xYESUB9l7KhMXFiMVybnl8Ab/sEptiMP8L4ii
kRBIBJl8iazZnh0lDQtfH8/8wg5ZEs8d28sELa5RarHMsjaeOeIQiCcDBzKSm1ZuHgzJgHuG2tqL
xrJ+7mO708Vt2K3mmHacaeSGSjz1qzDouUw8jTz0f4En3ugyY0aD4papBKHV/2bqhQ8TLIkkj/tI
HAgWzDYzqh8U/pK1CyHzkpIK1k2Ln6kcRXZtsdpVn34FlfKNa7N1LWnwbToD2M4Nd7Vya2fT5cw0
72J3xcFyQdGIni0oj8aL1tS2OeFx3FRqLRkeJoqeNBz960t3nmX2x1e3o4HT1Y30nlOOIrBkvt7R
HM3VTTb4s0GiLFpwIaSLHXgo9QdRUgIROmyIVfhofuOaujY47Yvaeh9wTNXfwEiSMFTcke6SMIjJ
e0LqNgv8p1GDBwemeHYq1b+Dt7TVovmzfmV+SPj8/kr3FMG42Ct5p54hhBfGXuHCgIyX1W5qPNl2
vzreNuAdJkjraIhl+U+JXFa2VZuWCQwvnrUV3Lr/8dMgdm8eJ5ITAUhed+ZKNZcH1rw2tWffgGb8
i1nvEbhSeMZ5ZDUHNvzm5KySVpO2HKNziIXJmV/UwovSLW5R29VWGLlW+fwz8JFECAmRYZlSXIpB
WAwib/DxOyBXsQyghnh5tbvYs0ZUq+ox5keDvW+PM/WqKHep8DXKvXHAHk2UoThzumaEwV6dbjAr
nmt45EoIZm175zY48iHDHfrRncsB6KBKmdjMojzlOMA3b2DxwC7B82qqHuOdeu8+QEeqRBIRGzOo
3h5bzU+YsUrPzAgDawvwSo3BuWROcHBGKmqy/ACI5mB+Aq/826ajsY2dU0LGT56huR/5yGeXM0+R
Z6fw06JIZZJ91u3yKFPbIVZln9NBcwG1NeOy3KPqP4b9Vm8N/mUHDltTnmgDyu6fT/3Jh91nub0G
1kzHYvVH8QslB9OFoyMGVb/nLTgYeLLyaGEg17xDZ6o62892zBXtoeUUQg0os1hq9vbtQF2+k20L
blSkrzwOGi9cDN8GM2Nj21wfBdnlTE0aJmUWMie53Xee+D1pzCBb0wiPmJRBTSZIklmG7sCt0Ucf
O2rWN+jDmjR2eORhZ+818VG5udtIVDNwSJabq4vTFwec8RPqat356UhR3PFaWinAMh4OEbl48dTy
lk8440p3fBU93o7MmMlwttsLlThuZd9auNFJjCJJyS911/GgTktVnXuSDjRdOgc5EXaylf9uvv+R
pslZcPHsdgoWGrqxgBq9YigiH7Fa/d4IU8cSOzlJ7IrtOVEPzJbrL69/lRECmE5bZPmCTrdM08Am
q+FPSd/mE2xgvIsKZzg4xjRUYGK4jiDPU6/ae0gIHKOoeGi+6LUn4XYNugaY+xzW9nW+LSRa2Bxv
ov3heIWUFa2IHUgKZDHy57KpAtdYqehHu6nz64i5dUErA7WCseM5sIi1cy26HaDb2jRe0Tvb78fH
R/7NVv20QQ5Yy1wcQNxFCgFD0xV7pNsRDiCjF1i7I0SUSYaHP/F2i7ilqR2/4RpPoxl1kcjEp8PV
/dkyhstw/hM3KX2ozvZQqD+jo6ES8F+E5FMQew2rEheF9Rr0xAnL1IBuUL56gNN0sZa3T2Luaf9M
mt3Tjg2/V7IVQ/89xITyH7X9ja/t5/mnt1EcAxtn+gjp5VHYm1QM06ZG1On5MnrGKPYOnU5VUCKo
8++HMV34uwLjk0uyAe74eGhgqpAYNN/sBCTjw9TrA3L1BiVE0hn5G1KRe8Of6PmN36eJF+u6amzY
5FaMRuw4Olvjd4MSzwlTTYXAITsYlzrwQdF/468WmpxAwj6M579v+4v8MkHt4B5zyt4ZFCjJcqWa
6jKYOlYN6ru7fm2U3jFRwdyFCYwNOCdTfPy2nIvvIyPBrphl/8pEQdp23iBujf3zZIDvqJ4M+LHX
hmrEXLfVRokZKTPbuDfQ9vMYHjkdzjthV5sT7q5zt/bAuxPN8CvM2v0OvceeWVgeNd2KZEu3Wp+p
ftn3kAAzEZpvvUulXsXNtcBw1kFMYV6saHURhAa+xGw9lpFeYVBhIEcB0jaC7AFIwWq27pvHkoux
0op7+cPrHnz9sjsyimHu0P3KX/yLpnTA1ZgoqlwLyBBxZvydvwF1VRyFGU1poNcQ+SWXy76vCAL7
csE3TiMR8TDnry9eeHEuR3ncvWiJ6D3qJ/nog6p2+4cfsW/cQAna3Cmvk3Lo7vlT2oZIzs7yJb2y
x7uyM6D6CgVJopVqLeV9YLM3lNz9+n0Ovg40ukzMJWAS5bpjZzk8m0xqQa7RTRqgD8keFmrobHwf
04Sk9JqcY9Gp2M2pdQz85R97AXCMSC76Etsqa9AyredRnHHIyXZyq8Uf4rKR+BVAKzba4pF/JKTb
wGXKqrd/DLEviN+cJjDbW6kbzNATe4GqvShfon+RJuKuKdFdN6pOhqDIJ2wYvoDdmeMcx+PIevbY
Tu7TKIL7QiztqoHywvuNZGxg4lA4fph39Ki20FoVixHWIhOvennE41yjmvRhzT6CSAmqRLSkfZyu
YNmg7Dqw3xUcFXLuMfkwVvRrpSIsa3Qv9q9KSlcDZdYYvX3TU8YlwmfADUyy5I4HzLoDzGYLTbxL
uLGx19EOA5ZsWZ6yaJh3pyQED3xlnt4/KQvEIa1E4338s8SVvv6+yXfV5PR0rcrsxP6xP+j6wTyZ
I8TNTjU7kSJZ0bKBdnIy9645Z+OWUi5ySaycggdAaw/ql1eLnKn2SQBeoikX7u5iV3bOyMGB8Khr
9MvZICoLP/d716zeFl16AE/nIngBPvnR8ejjm0WcbsH7sXWpDxZgP3hgcnJbQ7RUgF2LDSONnJr0
JA73jQkT0xgd3YSejJql9jlN9i2esPG4odx1/ZyIOuzX3FNliVbvfbjVJspvgx4b942ZHbvGV2g+
H+F2rYCHnrHSKFGPz7WwOcAXw6c1horRlcGo0N5N7grmOWsoZPYk5vPORxcgLjbX/FONx1wUTLEE
xPUQ5zH7PixjOJci5bOMw7+A8kGJe3vgk3sBXPWBbAcfULE7QrMtW9apgdlFzmibyhdUGLlMrTNi
NiEN2de6nlQRUc84FKZZolnTx8x5Gg8FoNbzm9yLBYbeV2G90x8o37xgIcdnNk7zHvbvEfQ1ELbB
AN3ZWOBq9kYYQWin38ipZ8AJ973Ikd+r4CVXb9YwiwUwJx88vGyWiKqVyLhscDlwUo7h8PWdfEF5
PhcFGMs04cUPB65c3hSHwVTUx76i508wZF7axDstbZvkk6eyasA3ot7ec0kkfGGULPpPYmY758xl
vGCTMdNtn1O0/iyiaM16adgs2wpTI/aZZgMuu0Pqell3H5GA1Ntv24euWmKG3fcz6YhTrO5K0J+a
/ycAqxX5YEDi5YCgRBK4QadYgO2puSWWhcNL3JKyygH5XSQrPH1HE2TwD3wlY/laIEKWtNax8NdQ
1dCdt8+vVZB38JIlywcE1fg4eognxKJTw3R2TMPnBJ5ukmSc9xWoRORJw3ShG0Dq0vVVjlMOx5BU
0mcPVjYYYjQpxGeBr/XNWQSFzHzBeaqKwlFcglslEGZ0MWoc/uFfsQbB/WfdhkjrNmUNlUTe9QF6
gJso4f+URHaEzI8nz2bKt7VTYYYoBYXWfGGonY1P6gLZ3Q4Ruzg3Ib5qqrfk/gD/dJQqiVte7qu+
KyCKFf/3WeykLmcyPT59ICjacBmJKIOvlxJ8UZiaPkbD+5J8Kw4SF/HJFcorP0Wm0T/FADViGRJj
q+UF98ZiVFN7hHgfuVXA6cHGDqbsT0piWC2mMoqbA1rvWZNorPLC/PoY9BRNyk5lMu38wbMKY4da
IyMzH2Rc4ynt/69CL+fQUZ+BIVwysR2t3m8WzdeJ58jIl0pLxKjX3Ee/VE0KNED7Ag0qu8KLmpFZ
hPbBD2Re90XxSp7JS2XnK9cno8rg4nAQ3UEd9tfQ9GPFGV3dcPPmD9OKJfvreK4PyI7xaimPiTEC
xRA3xjxzCb7PC1NbgGA2LXoK6mEp+5RbCOmP9WrDRyICMx4JvDAoVKiSswtrTAnQZGdlzbzXtHIP
HBsDyDdIf8VwNN3rAloG6gQ25oFibPhh92cV9jH5i3lxrAL4iV2tuz50rrV5QrJqpi6EedceMVSz
N11bInyHOwSb9TSE6/qhRWdk+/95hvXoeXAnbOhKjm5pU1KIiAkgVBBGkshyRmMDbW5Lf8I0+XVe
x/Z3PUiYqwNXfS4iWGJJJgV/aUVjJ9ytWKLmzUb6N6Mz4642CwcarnB1naBqPPQSO5IIXzWZeIBb
Q4/Mx41wS9uVlsiTnHeLdqlD5dbPB6uS4PQhP7E1LpivmICUFHPJ4//Vzd7IFes6ntmuDZ0Vp7oh
dwJZmbq5huZaIxJQCsMcsmYIf+GzPNPzYjgz6mA0mm4yfoAkHXL1SBhjY6NlRWl7ygkMadsOKrLT
xq3XGnnTRKZBkODV+iT6jk1oWdQondAsBgjxtCJS0BUueeRuBB97zO4CIb0So7zVmwR5A4TJtWcv
G4Z8JEFS4JemjE+lOOn38ERLG1V+Kd3tFj5dIypYDfH/iuKZJ/cjnxBd/9emezztHcsNH2qy6d+0
pXZTiEV8u7AUA7wOQKOofVmZtJ/oUa0eelLCgq+z07fw2klkpyTYogD6J3hoTkhBFzrNlr1312CA
JOEl9zna492r9LGBLkq+gzZilw+9eXgT+H9WLgGxjWeA/ltG2Rujki0ogiteCFfqRAZwpYm/ZNh/
hA7KMxv6NRAwfmysdejbNzAZFRXTFcvsECgyHgWC6YqklJ2pC/NHTdltGoWrVaEIk3AzikpDchoY
QtF5zw/5BwzwQwMOYvBJucmRGNayzl9E1WcENbmUt3d2SFKCLsqfY18s3Qn0qYKN0MYWJfVtcmdK
cXsmxulsMPVomVCIOxk1P3PtOKlOngnsSIxNTH9qGdrlyv20xS3L48nn/iyIsT3oiU+Gmj9x0vLp
rsAzFPHG2hY9MoAd2zNlUtoXO01rx86NCs4vbv52CUC1VQKy1U2QqS/huxxFYHghzGSth+pxQOP+
xiZb266VDxyLQPGEpUwPvjy9st+6I9wr+0Fi5PTNChIL70LuO2Zlx+3ELf9lkgoeNh65t15419CK
5fTwNkRQhuDevIEFApmH8c+Phc/roN18MKdrvSwARMSVn4N9sJGU3bklFGAZSyXYp5zVCjQHutnK
XmsCzBXQJHAcR9zcvuWE9zuALeEKm768ZWZ1eolTJilwSgIjUK2PvADHvd8gXo1jS8zG1gtnLi4U
owP1rCLfLuJg/ATk4x2nHWFZeTDv1K7XhBAhmjyvGTPGmeLhe6LNIjvqETT7owCpPTgoUYaA/nSr
cdb50Fg7zBD7fztJh4gt3AHrAPXgg2tW+V9mgX4F6KdFTvAucPmrlHTQ8o4fSSjxftzJd1gPLQzF
28rNGqQCN1ZqXZP52E2S9Oo49ZeRZ2jL2mcFitsjpswnKiJLzv/nHPOhDj6N3kcWRO7BlNvQBbS8
DdK1ClsLeDa6KrauxUgKTJsaom9TM+Ic4xapGI3vOOAdLZicTPZEPs9BnfeMtZ78ow9Wx0nKvDPr
H2y2c+GhXbjC5i5EtuQUoXD824ZTh/UAirfYAfXAflSDXN1brHM9oDZVGMubFpHGDYqXRgLZZh9s
FkOOJwUs1P2sDTs3agVJ6bom2mT4UpZe8IBq9lDhgIrknziJHK4nE4yzz80oSTpc9BpVgpZyaSzI
mle+WTB+mytU729VN7yqIgJ26pKuPXwVmiajDG+HYAzWn+S15a//uZznN214+aoOA8LUUnAWeURv
jnFzOsSWiw0mEWAOUN5PvWKJ3igG01FWBhDtsfzDekDAgrdqvhVQo3e0GVzNloNYuaye9a3baUi6
m/i2J9kVL1ZlEBsGwD4kTmvDkIm/BBZXSJ5/Krn/ts74oJMM9oNGZ8AFi0CM/Fk41YCe45Mnzu/u
uuCilcjPEe5qmSRBS+CubhQ9PGic87THYt4BA/xKazQp11czfG1BGLCuivxAsuZp/1llVHbz0no2
r2UTcHjJCo5Tup7Ot1TiYqFL7RPLLK15VOMW8giU4UZqb/Oq+kMJFHkvVX4GzMeu+b00z2913QZQ
LxyJBhU3QbrqvGGog6Ui1pym2708YHYfQNKvzKHeup4Ujoji66MtWihZ1ABcs3skKIR6/+5+O7gQ
+dzMLUQ9tvKOBbO/eiGlaIxGg6qUejrx3Q/LofN5bzesLSmU8zP7a+hLql2rHh0g8Dg47WzqfT8u
4TfkHeZIumaeWdUM4dDkxzzE86HDcL4fyJqLHK5YMKRvVVI7xS5tAGClCvdws4CmDAAxNVhlP94f
aTQ/HJxW9edLWjyzQYU01J3AI0KOX9eHwRPYG8DIOw2vJZ4XG4XU1o+/B0tnxIATj7OknkifA+ze
L1scj/mXzF4JzmN92QuSaD9mvKCasHppOa1C18S8iKEyeNcHsaFKA5ypumR7vmoiReL2P9a/2aa1
KxwvZu3SKp871DyYA6Bat/t11NIXbRXrXlSOruikuMaWtDqcMStEAOQp9SDBQmap2/gkTFgZSyun
PeUSAmlnB5cq96twyF4saT5rGRFo68ebHwj6MZD34DrCKPI1Jt0kbuClqAoIzWqf5orRkkX5MHuy
DNg0I2X3YSAToCAqoNdNG2wGGiaT5Eqd4QaHljq0QQygeTNh4zvTroyBTv/YYUDytZ4ZHVCHleFq
ZhgbhluUQmrPV0wwPchkz0jVUCmqoTzvPwrxU6keWsqZUevnyWiia6+17KwbbXcT8Tpacx2cFSYS
onlMJxKucbJc8U2cP8zC5gd1nqQYN22+nZSWruTYjQdHs3z/ehilaDgpvEotZUNZyVt3yW99mgXM
LIsydq/XE3lnJPXFrketarS6bxrqKU0rsE/uFWRNefB008xFfNRbGdOG/ZGp94ULrS3/TKftK4Om
dT1ctvGQvR/z3m5rvShAGiYyvXifS9gdGFkH1rGlVz1NyUhYIgE/vOlWo9V6o+9gn5z5Vz7PnEYC
ANbQBIl+M0ehFrIzhDPhaxtPIjYRt2FNPQjxSL6aDFKwjeTJ3LdXvvd4P54ahRJWdEnmpy0tnbHc
EXyIV1nUcHz2Sj4eB+HNF102Q/mjb4fLI4zVOZVYtPr9QNZcNIERsBZdlWPwLc6Xd/W5mjNQqCm2
6DpgOxRSdiEIEjaXJ0LMANm1jcf/YL1J1KQ3nd4HRkLlKUS4Yh78eVcxJcx37b0GSp/YLjNlailV
uKHSLY+HThL4ysWpCbYQo28I/z9dJgW5Aim30YEiuvdhkHACZndD8560DV4V1YpYoellHiU7FO2J
Q/ijeGwN2N/Tf8AMaq0mbGXzysMFBucwg29+e5pe0mrSx8/LK1VWyH5mWE7RAaH7iHdKnfj0X7fY
Hy5Okhkljex/UomfMPqOEenEjmV6L+RYRdnTB77CWachpjThQsJyk/kG1aSOPpeOFXUoJRRDKGB8
GfScJ5A6xTR6CGXu2GXsQiYTnVtFoxir3Z7L6mI2Qfv9Kc68Q6Xj4sWH+rqLQ1wMgtfz3lo8iy6H
Lql3yYLEIsDy+m8EPPqCbnPMJVNT4Lw0E9yZ8oZGaPjJXZFUCVPLkL0CuU+q1O2Ca9p/+0EYrihP
s9vsDLKK1n5fvgzds7J54alSiYWECqkMTI/sa48WCCZysGzYMzySiyLXlc4F2fOn34sJOFhihPL2
vZ969hGreC/ZYgtCa+3MP/GjPXG2o+TrRopHWZpsmIcMfG5eATAjSxQQuSGOq+6TCrpnbp5WBRdL
C2xu9oAG4s+L2SaS8jYkeTgwlW8UR0n3D9G6FVShA4qA78WfsYkR73H2QL0W6nL1I0SuDwVJoBLM
ultU1k2UAh58jPBmry9HOioOIJUz4vj15jZQApLYB9v+TdlSUH6WSedjZ5/CHOcuOcmpNqG7ZIqA
QIj1kQeaRQDkhFmHWWgjnP6FpmsU7qLGkLcjakFsipJAIpLxZydua+6nXcDiqWcDYT6Fh7jHhjKg
TGfF/LHt16waOfEVFaa4cpy0nRlLj/NftAZZLiJXDPZGXKg82DF//z9Jhp0mOOSIgEug9DiRVI8J
7xDakuF+blXsyLi98RK9w3dLFUqfggmGb33SLBdbbEAc8icJhcb31qRSp2GEFuI+jvfVx6OvWzGq
tBLqQyjr4FDTl+DVooezONIiCln2Ww5ur1jP1B1AjZFwmF1wNu/fv/kUJYFUh3AbdkSOU9C7/B3v
YDg6kHlYLrQz+mjG+S1xYnfjwZ3H8dyZz6vP/JbCFh6UZDssFFUrPmNR12Em6svW2el36irLOa5J
nXIARoIQuEH47W0x8IKNDj80eH9ufkSFdJomMs3QnnyLUUBxZoO9eDWtnjpr2Ngw+ypCy5faaI0A
OJJKbOk6hQihjvlXCaUxXeqtYNsED1Qe9278++Aq02rQ3Hp08pnsD/AB4jPf4dF1/J/aBaBNm2M8
aJgJopT9s6stc5+M/xtdodKAMIDCr9hHQ7/MyzpPydE+l7MdgSGe2sb+LUnMn7YmtgexxINPe3qd
zZBQWRQapFbqCayT3MvIfVZeduQeILqrHQaHnIzOIfi3KwAS2PUdN5pQWdEwTdL6Ipm0cnfURcTc
xImkKN2r+m8G0T/dd5ahKjZ/IgOCFEuuESDlH0ZevtLsWhiUykGW86num7sH4okGmC+47L3A9P7x
3YHoPuesFr4C+yFEWl388hcedEuAoykgRQ8C8qhqhFZWkE7QZaQroGJzXAA1NjMmXPmJqwoO38Q+
8G5gdfSE6L0OVwymCeD7al1YENDmDsLizOeCYnTtQTlr98zsDFdnEoKhugR2aVhxuIx+E5jGT1Kk
G3aJ5Y+zIVAK9RFWYuIUWn29RfZjJaXkVmyJUexol/jUSFS761ONkNa3WglI4a2b+cX2e0xYoZoW
374IVDsFT+J408Zli5jy3zXV9DRy91MbywrUZ2vBvnmeJgtWJmFbBdN6JzC+iAKerLTMllb816k4
qrSakGO3vUMxpVFtdHIaLh/9zhjmUrYPF+iERo3aXfqA27kIt+3PH1jJKNun/wflD7/rRrSAqmmE
ECKnYGjtGvOUkNNaL3MrsO9Ae8X5mXcU57qf+TavfpbaisZkPo1GR7hrWPndTQB4Jn7aW060xUlD
0WrhI8cOL2mRmrz1N32vUqJHEagPHn198Up2jRmw3LbryHWr49ISuzvZndrkcz967DheloE3xFTu
VBOgIdbRbZTPhcdxDKoMhyBdz1GAOSDgM0x7UaEDnpGvoQfXzse/qiXJnNOa/zvKHqRQA0WfgW9Z
FF1gxvQn8ZapUWsGclAlzTOqQoAv/qaKnSxzjRhCjHQjTr1GvmxFeLMg9oHA0+djahrN2RP50oyh
ZS4cAmKwdRp/KKt18u944Iud7+/fzU5ECh+A9QAbdWifH9u94cLh8BGr0GQ9voDzsPdb8+95TOml
2Rx8QKJ2OqD5xu1R/VGePxWnWUR5wSzJeR8i6iaCUxgKjSVdlPsNODA8I0N9GDWGaQjGayoNJjmI
3/ZaVG/jS7Ulh4BB1sU0C9bz0d6a5qdUqgtbeNLycseplMOcMWv788mL77vhBE8s6HCh9cMMfFWW
/jxiOfYQ1g6MQ0e1YlBOMjYqAR02ZyTGN5YusoTjdU3k1GgHn/HSB3iqIImbDhpwEKkh5ajHIN9E
I16Zp/BbwAa0YxtXLpz/qZDSY//7hVR0SJXUK9x8HcVK5AbSkQs+0/PkbUHHC53fiFn2C+xPBGM5
scqSh1Upr6mXbXNtP4gRHU2XPKVr0hWtfcA/rq1Fkw3AAVbVVCjHPq6mXJnTAosyF5iO7SRTTMQ4
dKQ5rWIi6MdJluHCAyc0ddHs9OLUwrIOtC7hoNZSTiU5Scf0bg06M08Ih7Cmh2k/ktzJBrM/j4Ph
q1/dd24EL8IeOmQr60sH3hHlz5L1SXfpCjh9axN2Yz50+U7r54qqHPBVzbtRaSMYyGdtw10SJo2k
ze28EEWkP8c009xlJ6KnLKFuYYsuhWovWy6V3LkLLv275+AixbomEPuP20wfhz5cOi0rhr3QsUcG
Au+FW6FPN5vPC4rp2KeYbxltWoCnt1XLVnLn6Y51gAQdaUZhXAoLevlsDXxckMbPCBuXvkeaoNZW
3l0QOplLQ+LQdnIvrtiXzqV0oBQrmHc7Yn+78QRbtbZyWkrcuoeBlSlKtqS5YsD6hLxCgTD504mC
LrlmBtOvfOxlwgYOcSJOMgpsMlDrqPBz3wY6hVvILiK4vpawY5UmMCD0pXl00yY7Z1gzbSpGb/y0
gN9J2xZq2Bz8VZfFBB6yOMr6u220UCR9dTkNNqg+pCBMj+a2fe6w2jqA04J8YtrYRdVw0UDAd12v
Beqwx281Nr1329cFHBFxuZufTNSL5GjzlSdLEwj2OtekYP9NPbzR0x0aCKLTL/8J9Lce6cxC8SKA
bjfIrER9qlWLiCd764K1Z8NwybdC0T81JmniA5up9fiiY/Jd1ITtb8986BgEIcvyePbp0Zf6jjHt
JDTDSpKYZUDolTmxcJTmlW6950AmjpprvpHpHTryFORqseDqm9wPAsZoxaUY7JjvIP+i52w+Nu4f
vf4ZEp4GjWcG7cGZtngMI+djviqJYujqehSIHkgJY8/7blHT3TN2TN18KR7e/MLxBz6Oet9k96YA
TdPxF5b6V/50txFoWhZ0IZFYwLQ59j/dJd3xEonGUEC4vSVDDZu9xhyM44UAwzUk17MDHIJpHiwB
SOfWNaujOOf3QPONayGpvacN2lSy5WBelhQMAn1iUXDCjNrYxD7Kk6+6RvBwNi2SkTfa2ewmCeOL
QvqS2wmZfUEIBp9kX6qeQ5+TUiyJTyTdH4U7rBNguArhEYWI8nRb96II3TS++otKIQy0g75OJBjB
mb/sPaUdmtCeaeDdSJCgaPShAEHIBgfrReqKX8Ox1/kErkWVUxAOz4VwcHL2L6BnAHBN8SpVoraM
SxdplWlB+5Ig075n5D9CWbOGgo0I4a1O8AK03zaeplkj46DeCuj6p+xIT6bG925J302cGiRy6+s/
kqdIqJhNoNurqo2568jf4eSxEjI5QGN77Y446BwoFpz/du6HvMCExnNXlAbMFpAj7hLGCmoApcwc
rS9MrFarwdX5UCxibeAfMDsVV8fR2ZLbIatGfw3cr5AXqRu7wfes7l88dGUjUSHbpd4xzzbgyuke
0hrhdvw32Ndz4VkvTjE0dI7+09DbWeS0Isn3MBGepU7LMlTOecvrbBfFiCkA3AIckYIcHoIo1obt
xwdOhj5hhjNplkF/pp8QVrzIBshK752xXltPOJCs/VhwBGVMA2j58BKCWxPJ5uMH2FJq5RlrANnz
cjo46sVZti0pY/Ik/fvY847oR22weoI7Q+n0z785jfvgJCz+GF4VSRpnsASZZDuHvbEPrp6Qhw56
hnXwxJv9hby0XREyjO0keF7GovGTSUdGY2iO6aWDFUC8NHV+H+Y49I8EfudnnFz+j/sGqEVpuVL6
JKeFIl/MDBnxjwP9zDk3TDw5zstSXlNt1gbRsRpR7IinYMOD/xmKFEH1kn9+EOE4ZYXoW48BkiBd
Thm1Ktf4+yUBHWaSuJUs1b8h2VAWyird40QoZG5eRfj/AW/x0D5AZbqtoO3u/bP/AYVSfWr2gl+E
rM4O+4MaG21l5SQDYgfNDIPYsHrSj65CptsazfNQNOkrxmS6zQuTFf5JeBt98aiLCeyCG/Jjmtom
9KsFhi5IGSPMGy4oIbR5PE+Sj+TmDAwyZSZ8vb+tjdh49sJKckCsVOXVPAEGRg4EDApie6iJl2Gu
vtaK2f+zPQ0kAVtAhA4L/sN3tjSp+ywi0hcXBpGuWNF6AVU4i+cBZmH4xTtKGTJtPG0Xe7xptmIy
lDHlCbYMthuGlfTu6gqyW14qmqgSracxj89jAPfOH8npsfsElxXgMAiPzctkdqcnDPjuSxVlqhN+
s6pr1tfcvBF5eCsLtJcfXDz42Ny0p0GUr2dekhcFh8nB7Akieo2T+DG58Xg6lIGNAx69YCghH3BU
GFzDrOCqoYi0FmXFOE6ALyEXGBL8maN8+DpNAh/JKS6/QWFW2p0FdT2AqSEhfTKfrhLWm/WSdS1Q
g/gVZxJkgefuyx7XU/1Yf1ZhBVX4MxxRzctVsaCV+oqRtqZRnx/qrIzZoXnsUKAzLUaH+QN1fNNP
CLQYmTPIl2ohPYrxrvaaacMxY1J7WwcQOk0zo0ZaCw/fupzonOa+MfJaUkX05CbmwMM5SSh2KwKh
QO6T+lv5UKEufREf/P3bqnUYPZdMuV816+ENLNpW3rLVO6TUdVhT3Q6NaSR2YFgfkx3eWyKZ9ccs
M0pmUgGHvMix0rVsD+IiJ7BhK3yewdBCNrULPtAsZIxrGTZWMIyzUnCUJCUkCr8mhOYHl8G427Qc
fYYklYwVWAYH2iZU5+zIcLlcNOVPCjtt5ppoZRHC3ccxYIo5wSBXf0LjhEvculS+I7Asn05Ho+rL
j2j9W6XVz2V3pQxom7/rZGfdutl2eVQnrXB5OhI6OjIV5PGvGvww4QvQESCuji7vzuCU6hzmESUj
bka6mNF+cxb84hWGOExfN5APHdtoxvnwYGS6nEnXfRn4ZGzxQsleBRTK12N+kVryon6eQOIT5o14
XVyzTV2b1f9z33/jtV7dpWv5ccOZ49j31vavqle+VQFqFZyC68OTYbudAWetF6iCEUFklHbbq4zs
/KAgFXsTJwJaMVHLt7624VtCv19lo9kgmJrI+27JAB+0zW9Nb17+rLmVRrb2CsTQzAsxV44ooTnm
KkwZZEHUox5BFMPuRjrDzGHQGDsvlYe0Htq1/PxIHEkXyglsh9G87reXDp5a7RqOBqKib7u4Qopk
21gcUjhQTtrcc0FagAsGq7xk3+are9bdJYRpNrhX/xMGPlOAqI97TMWqXhqMK1MF1m4yyfVKsoke
SiKNc0I7HOVVlB0diRv2xJT3mqa8unCcUj1U7xjH0DEcWSX4LjAZHRQb5g+vOzD2idS1ny9X0VPW
QooUU42+cAwJkVX8NNtlHI0CXGw5fr9bn2nmbISfFRqZIkp+KV7izK5lMisGM/NP2G6J9BIEMZL2
KPhstAvFJ/9MNfNfptntnpqm9OtMdh3U9mH2T7RwdbUecd73ZUwm53Jju41rk/ECdsX1I2L62YBt
mB5plrjXKXkoauTPXX4RERvu2qdeBXMG3Hf1SLIFO8jyqcDe5SUj8QD23zD/lCzBCCmOIbeipSSK
V3qCEgMhGx0AFNYPmzlbfzgxHKlNTgqvPbvy9JBkcVvAdY6WTwSMT3iZ6y2uD6R+yCbqmOGyo9Gd
PzJLN3h0Be6qH8fP+BOzpsVjjzrqiSv1LjtEsvBrguj16F9bFS8HTWufDgu92AGUdDH8fw0/Y+5G
fGZbmF5KCE05zEtX80Kknq8sjuT2+8TxDFAv2WUDzRLVojqx3atby/zJDN9ZgN7ppmCnknIZeSLM
cGSBDapEZVvI4oHGzZycgms9vRGdJ5KWqZ5ig5ufPmdU7OJff+1A0S1XtXtPrR8hGpPWDw7Ci/pA
a/KmaGUKg1QvqjJQD188j0TGQoPQ2LBLTVPMK/K8bwnzL4NFYUSwEBH/k/ojpJNfKIasnsO1GXCc
RfW/yHt9pM038g0j55X9AvmEdFXqaMfFaENJvATEp5teqyRKgqsYoGRcf3s03RuT7TVwg/2u9j8A
PnCmsaQ2VvMfqi26k3J4zF+WR5sFp3HXl6L/KUEcI+BqYDJfII91GkF6PVp0oSFnP95wsH434v14
SR8hT+7AJN3SIdzpCABj8bXor6k9iTABKrew6mEnyDI0UxsbhPxei5jot2Qj2WCc3TNlWL5PeYE/
rDF0J2YrdpQYeojwFQt/ADHOAM72xg2k+uiTDWqgBfBk/eAsALvonol9qudy89tDqZUC9xbszuwU
cx+UPb9maXm40yqEDjBsPqjUeun7Zd1eAOdtnkEpw/4V7/RPtJjLwlKlwZAt9hEf4h7SkEpD+ZfV
dNsHe81Ff5XF3i2lk4J/a+x8+1Yd6D+EJ04uAMuOR7H2w1ar+RsYCZ7X4aOtef65Z8pdq2HdWS0n
V1ajH00hIV/ksG1ehVFnVAHi5YZ5dBJaRJhskZbOf+qjtcukEmoTEOUs/pukJYP89Y7vnbS7G1ct
BC9esZUFyN4I/y2lnJX8rZvpe+V2RX/WhFBiCeVL+becqHUoBKh4YJLyURUYFz8UUJyUh6iE/Spx
dGxPHHhK8pCARJdmelatmwCkzS34+qIAZK6+SjEKD+kHwPD2YkBgmaOa3pPrEve/AeBtnDdpxeH0
GIWtL8CTwFfQFU8rLxDK7XLvG9U1fxPCfUQnEsOaySgRKTHwabBzn0rJizg2CNfe4TD2MduYJ264
HX3JG04l3y8qmMpawpuaHsRQGVEEWmi5uE7pUmepbBldBArzMigH3u1++LJk+xKGGw1Ad46Ce9Me
2xDeNrfDxmNXmzWQSSinRbFIa7ne8fLbw7dKxP8R/J/syYHxgFJkyIoAyXDPY6P/pmD3IFLqiZwm
+yVtCG3kXgN8oH3vQSEg3AJIlQU9/YokKdRZfhoZH9bFzTfpTqoiF/7BXy6Vw+Rd/F8TM3opmWkA
N3C8mYBQ5hkFpDj1V4UjtIZ6Nnryjna+hDAyOkoIAKWVsva1vbewjxHI/bBc1p9OsZlya5W44Ucq
4qZCH7/RoS9qILXLWgTdLhRI5Pi+mxKl1Lh7hm+UL8VZ4+2eo392C2Vb2urQnJ404EEkzeX6QDId
xEWO5s37xIRP0DzpRYIU0fdj3UYQ7kWxe/u7Bvp35m8l2RbIXyX159+GJC5WNTNkQMi3ZQDa+gUS
bN63hekzLpahdX//v+XJFI8HU2CjyG+ZUZj6y3qTgK+ulYOr6YEyiBlK9OTJO/H6bXrqDXBfwlW8
5A1eezhip2nqallEhGDV1OARmnDFiBuoYftfIDUebsf4V951QHqW2bc4EdAkV0Aw2mHz0uvy3anV
ZyTq30Zc7bUr599rFxXEhtJYK4WhV6O+FLkwr+ADdqD6x9WnYJMCON6wG318wy+2H7fpa0+kca30
49JudgP46mYXUE13Opr0aamL58A4MSghPAJHFZAvOwqguw7AUg7xy8Ddg7sejuBrI3BDcJScbNXa
JeU0z9bGuv0zN+hlwPy7mnH2nnUk/knrBXEMmrXYs8fd44gNYxncsETHNLOn+xzijOpS/NVIeNbL
wG/bYRwDMBQ9Ifz0CMrTw98cRwJ4UjdKn/F0hRlX8BCFc0lA+sAVWnoTSnIq/FjaLwxP/fJEFV92
rKwbbi4EVsrNQ0QwCZNlMi0XbyW/a7tdOK/SIWgpmSE2BlqkDdcZkC+r1WjvvAFcZJ24rinVibOe
fE/7CTMp50k2vvio91fjGYHmkM+BcZfSt46h0Q6Ysipcl1f1s1fr8FTv3xgf+GFBzk0zrwQoW+c0
4ZkenjflKJAXxndx9KL5aw36GYnJvgcZV0e0jYoclQTcr7x4qkrDCpeMnuTPwaxwjBKTV6lUXuQA
HrrSy9p/vYcmNii18SenZ7duu8o8zXTfU6GaykR1hIZgMEFOO/QV762wz0KHdKh2Cm0ZToLllqOy
4+HQlsi/sEOjd7cYxIvvgkScRMivKk+Q+f5Yi2ZrzZgjVNZTAjctLF8CSVHNGF4MPiRpWtyWcgRl
qP0rb8IG6GWz0h2K7TpHZD6pOcNKLr+6XQuDcxvsm/TGvKVcVeqw24DFnoqd47u/kNErHnezXV/u
3Qzu5ZgWGU7ZtEB0d0eE98o7ECqc3GBTyjKe8DvXXPTqiW2IOLd8xyPxxSiNcC4fRvOH8Q1s1F9L
ReRJZNVp3ySeUKpwDiMTf2omuAn2mMVbVQzzNfQUy39fLU3cZ2H3hDBg/b3kzH/Wwl4MaD6m8/pF
YuMtzOfTpjdQ6aLiDv02wN4xVdqIG1zAg6ZeVfTpZRtC6oHMth+HOtDPyUzRmhfXRYr/CmvvPHhn
xtw6cVpf8W4csYfydVrbN9SKl1jzURqZjlKgqb+lEWNxUshKd3locEWDI0hBhHwcI/nMx3Mz0sln
yM0wLGWubI6kJ5kPJLh6G2G88qB/RuF+mSzeBTs+dBqL3NI2gPyvjT1X3b+fPhfFnOWf46sYos/n
/QFmjd0wjvr5d/22WKn/hdrKM6oE9Ht8CFu/7oMzvhJO+CFDbigc0gqYWaSO1eDZTv2szrf5u2TC
8FVAPm96fFOLyWLsqy+IAengc0RAcAA5d2isWAv0t7jkrVt5S4W8H1QiY+KpL8CknAPHdVAKATTP
2goxYs0y1UPwayAk0rNNZGtrJZ8sX46rWGpjCCo8rHcesWx4B/rz45RA0AbYDUjU3itrpWS1S/PC
YcVDbS7wtSPZhQx/4AG3nCGgJ0Uj6FsKCNlb4f57IIb0szBSTOu91giKSvypVe85KZxE4Pr+CuIN
ZgKvchFkF7lwDoE3hQi1oENqt8YjDNfhzTHfq0Fm0k51L9idQVqpASWpUu+89grPbQV18S5hHeLs
MSVJ48xknqqGpeHm8fIP1paLXpU6Bd2I7Xa47BT7NoKFnBcDSTaV645rS4sUiK7v1pTgfqmyuVoA
ao7HCMfI7SLEyun6QGnWOtgenDepzNCczbqH4O++9HMtR0vW3GaJbs3aQVy2whFijnnc3Y8uzuXg
DX/MhtbT7uov0h/qGB9jIxY8DEQiDlqFGqLxWqOPkPhmL60g5ELgDBADJ0i7JUOhTgpF4mz9vFcE
bjc3SksFWjaiH3SiBH1FNisy+hZMZ7U3W/ioDd9BSKrcaBQL7nPwqnAo6xnrCPG3waoC13C1FGJK
RRIFXEUa2Iu7Q+2yGco078BHKJCFd4OFkgy9l9Uac9p52fnjGuB4o4tjlE7y2vjviQV7fcq1DvDy
s27l78GCaEJO6xk2rJZCd+EfVtuBEF7h7+pYwVWBRy3t28OwxD0QKWRSf+wbI/sCQ0Rj+yUYsrmN
g4ziuoxUr2GeOctkWCx7u/DE46tqGhHs0fTkvPJe9s5d3xp3i6xL2pQ7sM/f6QQqKowR22nUo5tn
g0D0HYHFpdwpiEl3BuVi3Xqal8ZGnYdYLttZWTASvfrLDV8PuL12Z0nYSZtaqQo/UO+3x3yLSzOQ
Gc0FDNmMz1/czUq7NATN5rZnXqBxmKbFA3uvB9YxUsjwdVdSwOBiUqaQ5omlvxa/OBfU6qKrX2MV
ZtRC8zFGNCAqP42rejEQPbtcRR2hj1WhxYhAcLpoN0C+uXqCVku7oWTvy5kgArPqzmypKUeeRfJG
B4U2bd4WJfdfuHbjgr1aK7HBOs1CFAMevzTOKs1YJre+SJ99Bp3f44iBf7bu7xj5Uf9ZVSRI1sRe
GaQxdx1N86u5Fb90zRgjq+4yMMURNY7qN46uUztMwYMCEQIYpHgKydpSHqccuFj4plg5N74ABrPx
BNWcz4HcsNL4Qvzz1kuZI9g8zJ7zDsuqJ12smZyKdtA1WRDP2AJZMC/QoB/cccYgBOiX1AA6FRcY
iCu2nvw+m2Q+9nH+dp1rWwKcLdtv6LlXhSiGvMvLfmr1DzinacevxB4iJqtlIGOP033+LQDvVvPI
mrV/W0NdR+jVd5+GdY6omW5PK4YmcW9CMP5zqvLodmeZiJ9HmfkwaiY/KqnppUBq6Zm7VW148J8P
0OhUDjBMcI4sgwqE5vnTXKyM7wyRYt1FscBlFP5L/pgrWuK9/C2GghIw5R6PphUdSSoYG3b3zJfA
azKeu7A5bVHVyL33iRLgZxWAWkMp090nmHgd8x88RrIJ0TKrE0A1LCOnypV+HMIhAuBAOPUHVHot
JujlqjnvvI4uBkX6jYQ7BNbP+F9fr1DuKo1QZtAonjrpwAwxPs2CsP1EU/UURyVmghJlHnE+Xnz3
agyWWVKHB885Z5mPherJgh3BBlliTdWC/AQGY5e7nlZvfUrz0yDGh2qroK5eqxSVz16wPBHKqY6z
5CTKblN1/46Ioz6cfMzpr5mUafqh33tl7Q3xYIUvSQ7Lqbd8+BeqMRxaMfBcuMETEXvHepQzfI8A
3Of2E+n7C0KZe6nW70zDuPluVKRFzIxTMAr0ZO5Pr1wBx1AmqLTQnwl6bjD3OemAyyUFUx0t3hLx
oFPRVLWcopZW9I1i1ZuFQl1xuATffm6ThoczcoVwtL/dRc3OAaM1lIOi+pzYI89XrKBYNrYzdQ+R
gIvbLL9VR8E78SCzxmB06NaKEVT5Jzkgg0MKSsK3RsR/eDJm2CcHawV26bckLc/eiPA45MVM1ZI6
BpjktRwirTThT4b8GI0tjotHoEZ6WwHvPQyL0Eu1pl2qtiUdv79hWH6IH4BW+6IcNMV2Wipr79Lx
gQali37D7SWtJN36FbmViO+UCNcZXnMgRGKHNCiImmoMOK02y3ga87nxmnLp4KJM28t0yi978FM8
S5MUROkYIknrpWZVNgAGNZrPldqhS65gaM7IXF+4XK/kAFR/Ini2flZiRVI+ISnF9BYKGwFFc02N
ezzkyaA/2prVEc9yLGhu694h6rM/Np4mzPRXh+zCj5qid2QOaF94LVxMSS4mo3IbXduNk8i+Tlqi
oQFuWuvGaktnnV0wdtEXNpeRVMcn5l2C+Tba7hDDEDggIPdviQg1Rh0aPl6mSj/JlL5nwlBReboA
QXgjAv/kK97Bb/pfTb7cJAfaGULMT/h90sGEkAr6RbfnyctYa3Nz4g9Kso6jcDR6PbkELxM7ywl6
7TQTU+hc7UtEyWtcgTTfnjqao87vm6gcUu7MvBk0916ebPv86Wx/4yDs7bWG3FwyGl8Xntrn3Zei
CWsNflX29lLOomG1RmhijCL9w+bgXfgwzmyV6fUhdwhWCZpUnCwnPjqn3KLil/yTjWTd6gSAoxTW
HlOBNdblcP4rud6030kELh5cZ4ch6yZJA0du5HN7JUnN096jOqYLOUPiyv7cOOuaUVuGBDGKx0sF
xCPubAVLA4Aa2rXWjO0VVca5gteJu+UAjRxgKcNAWhsNLyWG5O2W2oBWx3cxk6xXu4yiPRpYVsmT
lMnwc7Z3EqjKSggkOjYRnY1/ux+6iGpsI3mXgzN22bK3z5MQJaoB4xJwooOTf8he7Llv32dDmz1c
yLCzzpl5eeYTDiyxLlSwXh5jPaStaSu5aRPU7hRaFICTh7PNBf5a+Us4QnvBkcbyyj31Fd8uPCeK
xMSpgIin56cDQ5mEHzGAOItmM8mqR9xYn6ESi8ayz2glbwjEDXiRLKrE1xQFrmSu6cmVg9Ug4oOj
F14IjCrSl3Y2dmfJqTcpC7BIjUIM37RDyLL0eoHo9Siug3OVP8sJkET91ziNgpkW06wwGCtcfGPC
BgBdx41QAOVcuiqGG205QKJ2m/PuLS7LGaJATwtjh7dFU1nYIOF9I7QQN/n7uCTatYAcRexHRTQj
FborC3oBv+HOAp3Uf6ghLvBmIbfEG941H4WNby8erTPPPvO2nJNWZdH5Mhi3/gqQ6SheQA6AFEaN
TpS+GVrMEbtYAC1H/y+HtTeSD4omD9KrW10gk4kOx04x6ZzReljTTX03y5sCQCNOZzGsiuVdoIRg
6oUiRoFBIXX4AtvaLpQiuRB3YBfHCHYC5qdY19Xvw5QbrTzvaV49i2tzDteNYVwMQ+h8/2+foSvx
8y9zlAH5K0ymPVFRyX0Be5BnTF7pme3MwGrUTm7YZJ4KLCtZpxn9v728UvDWMYtqAIpS3XZ8lOAq
oIY8XRa3C6TSBzYrlYgU72M1ji0O6KivSVJsRszwK6NfApaNZpfwl4ORgLKZc8faq3Zoe1vi2H2l
/sOIJcxvTcIrPdjeDbenkLRBM+bhGuH67IIJ4frxe1Yoo+RDnOwzI1awMeRNRTBiGvDE0iG8a63p
Im195jUF+vjpd4mgFIOTD6zEDEkoQlVnUpN7noGZJvAP6Nv+B5U1YkrI8ICY3lLBJAGTpg+gTcsC
HLS8bqj22KueksCPTuFqsXCyg6kANWjePAOPSHNY73u5lp21bZAAKq8ejDV1dY1VxDxrxx22lwSt
Snm+0WZmuOLvKkxyu+Oww0YQieJUe2XZm5ZjUjCcREWMrP5SwMiat1A+okNxrCuR2mGH+CTUq6gb
smq/3UW18TDtmDs2c4wFmntSl4UV9MNPc5st/pdg2DYTkjUSQ9CWNIjU53rTLestKzD7xk+hknsP
8o/eAoXLc0aNc6UXyv7as4tL5SUoPlZaQKy+XNVUN+M0S2uFC8+jIWP5CzaXP13tsKw8M3m6SzEu
xB0xIfO7KmxdxW03CHe2dH/8fNjC+XumhCUR4CcUSbptwXv5kHfACS1ElOvUlb4utwsyAJMULgZ3
wL+0v34FizUnCld4Smglv0GZZ0naT9gF8oGUvZ6eHWnIKY6flQoz4/lEkPA2taSDqH/IxEYbt6Op
x1SDPUFmAEYyD6+PNnzdiVzFWlxv6wS3llUayLcK1IKsNsy2t4AItCP5QhcTpzf22CJubdeFjSpB
ubxDziX9rzMioO9ZNsiAhc6R4qjbnj0ueqZeCnf0eOPIjDVMynEFUrQeSaTVPUHqt6A5tuc+thqG
5ycmciEHyxUgwAwdVJEwPklBOMYqBCZfKdoNq6cPFPMcs/3JlAnwQSRg3Rf439tG+csDGl81FRag
hHT+tffKW6PtEe/FQj1rAaxDVDVBH4QnGITxIRGiwq81mPdtPfJf+HQ54crRhUaSyfA1a2K5FqtR
lujj89lF6wvHBcJpZ1dOfB2F+hfUyVG7Aj4G5pvU1G/DxTShIwncXv7rxwbnjaPCM6plqjvQv6d7
SkOTg+sif2krh+NaHuj1TYBf2btbNwCNSpSQlZGbnOYbpv4LV7+Iq6I5eysskIGwBtxL7GS63vlV
B3aJCXjApRaN42bDrYDxkXTWuG2W58RHuewl0rCy46O52aah1rTSDqQKyHiBwBhG86XCl1TsYCB4
QahEGKDsYLWJBM3IKQZQ3EaKe8z9IempQT8AOXD0npRmE+WmduM/N9xYhIpnLwKew+r6tu8LkzJ+
8h8TyJno65ppCHlJolWQGyXzHzQTcTIafmPuGIe87CPDSwN1Y5i/aWc4+kZYVGCWmxsaMQLRZflb
qpNQNTe9VtASUJCz6LQF6xLk5A+wGw1FUSDDUxUEqJH1JT3zfhT2o4474UMHwtQ1fQUoh/F050Hj
XtO7aOPPG3J+S1QWD//SGdK7+aIiAeYsqVX+D6IRkMmYvYxpGkYfbgNUpE0vCCBCpBCupPlTnoT0
NR2cPZM6Ptvn0nJgvR8P9GPD5tvx3gzjiuaeopKc2BohEv+vroDLj9pMiC6KVCrl/mc9069Lgwch
u2CJ+2Kw4wDvi8x/qcHI07puS4hxHnFc3pPCF7hdArLgXVmO3fKbtmrJ0eaCAdAJmChlQSS9c1y9
E/ZtSIlepWRio4H0I/piWtxi/ueGQnpRDjajJSQeVKoeDc+4uyXeuWG9y4GpgQj2OzgohlXYjxdk
5hAlvgoIj8Gu/qA9412QFEAMgdgjM4aiZk3wkFR0kuKgWP8EXoACin6/mkNh7ISrH0QSLKP3ezol
3AJLu+M2xJCjrBB+/ko3Gr7LDesJ+JvzRV76h9eSh0BM3/3lAfAjGRJHUuxOi+m8eTdzpCVDoVld
qJRB0QvRTXuqnfyP5JAz58aboa3v9ViyVgaf47r+YefKLKbbD5+bFjvA23odNDdFcFMhou/Pp1oB
PIr4tz8dcaFDriHB2nCEl+VoOzfXtajd/eD+WMzxYq9XmkhZg7Zo81+yArkgSBkydan7AcOvnOG2
/jhi5wcezyDOfXuYPok6CyslFSW7txh+ray0UxMhsA8DJRlptsq6Y4kI1MVrpeEGRKq1Ry7w7Zn8
FWSxbUUerjnmOoY4gAc6Mac81pKmf5cKx1Y93dvD3QwaI/mj8tPNE5sQpYuhQAEVWIqvz/+stkmS
a4r5PyF8BuufJFZOcz1/Y1Js7EGmFXWY1/8a6fSx131nmS6KA9vFMd3qsGAdj5YX8mV1E3MpxTgV
8+QjwPQ73FTPPsK/gD4OwYpxgfjjXxtrVJSYklkOfZ9j4FSx5q5ZZqbBwLpa5pb0vT2W9ZhFWDEc
fs3ngBCuryeBMwRjWRHjk2Gf7zaipWq+8WA8yQSSBgBB5i98IqQTqokRCUCZvzyAp4jnf6+7wKn7
UDlC/NzhEYxUv6lt+t2CejwKsgdO6OCz+9tM2v4+PtPC0hNS6x+iCHotxoE0qaqum4hpKwFL96KJ
fHmkodyDAxz8Dg/BrqkcBiGiFtrHCT4XqXI22a81owIyWc79jVcqT+yAfbszv03zcqA5j1sDN0B8
nCRmfozTHbkbX9seSGHM33YWZ+N+5Zrr9Gp7mg3RSOO15tq1PV37BpkvT6og2R8TktAdw8oa7XGl
q2xNz4ZdvAabCzBRLfw0DLSszO8c8Uir7a5RLOWJ2nVPbQR27FTPj87LNxFr2a4ju9NYY1fW7AjQ
NoS7f4VklXbD9EFifnH5DT85TlZMy1467COlGT2+nxN2chW8YRn2vesvPga4R3ZB4HoBbvbNWfqk
JSaSk5OfCN4vIJ9mRhIm7DLiv/KpL+TPFaU2br6o8dtRovo0Ctvkj9WO+UYXb879e+I9Jr189py2
lHapfXolhtHo96hya3Zw/arYdfg/4Xr8HXzL0PtBdmmiobq84oh46T62RRZHbiIzuwSFddlkPM+j
/SUH7aKU69aNGC6szI+CQlEM1bs1pGdrNr0wL7A7BPlL7lsr9gDPKhtGY874EyrDk3qHa5CmL2Be
+dqNQ+AwhQBggqqoZ+p1coJrH62YXH5aNRwTNgX5P7mAozc/mqd0JcqmlEZNrrsxSPXkafuDhPSq
r3CTu0RTLbhb9QjbF9F8PtVwkdKQ6q7dbdbvzYiXDL3sBLjeyuW4pIRxlpxuCqV5jCJsn9A2zwWl
1z1jK3lCis/dBGZImckMMNs5P9COXk59EwkJPiIeFWHsJrIRDOljNGhln/xJkzm/KUfXQM6ra3Yx
L5K3K5tWKaEHs06XYSJPTNLbAxmBw7A1CqVlE90RSdkxzT85p7lQu/Qe91otgKQOWpccEVKhCUIJ
A9kUZ57s8uZIvxiWoRh+Fz7GM2oaAGeLLsErYDLv/JMGgyPw//MyWHEeBpNAc0hd0hgwgMFF37HN
bxh7FDcBJtnajFMo8xZ+xoLCn3RVRopStRHzo5wCVQXjUVd4U/Fl7I9pMI28c2xY7Xu3TXOPWD62
1wqfd93oUo8S2FyX8MPmDY3p62yQsRvxQAZVNmcDdnNcn/sikGfJE8xeRtx4yYfoI4rJEzACMipr
X82+BKwmj7vHzeLfVSXX9K4Z6NF9t9f1t9YKVy1d74LGRr3ehLWomm9B3RrSh8Diftl4GIerdAbq
4tzUvMwmRaxjVNsNfC4BT2Mk1O9V6rY9LvfhFzMB4Vga269c4NfjtcChdxzeKWw8fXaUblxZ6PHy
Kea2XXIc8D22SMuOx/iZnhMSQCdwiPbVe8pkoRX2KRGV3/aXXp0tH7GcQSRUfkiuC/JVsAX7AF0B
U3s1r1900ifP+gZsd1oM7bYudeT38N1oM2l1oZ3cIIE35ZyyNKSKXnxZXxqiuBQ7yf1sPOos6Cs/
siX8cBN+ksXjxeIMymAUZbqO8/lyVY5wKjvCcM8xZuSxVeLs5HZP+a7kdDTiEx61RcAgdtHhyaCH
5de+mnIRJN0gluf+txYhf3j7ofPugmq3jEKSYj9PptQg65YUpnMcxiVtFJYlTSdDVOBmguIzTrWE
Tx5H4cqRu+K8nZ98tbo9MLlvSgXKX0jQzsoQJs33IiidhPCg+Q6E7tZ+NfODUmH8ADwyEi6ksLBn
XQdBB1m+mQho4ljHZMmBKhol/1GJmHrtliyUdfhrKCMdBsz5StnmFQ5Hw1xlJAI4DEvbWcsfk1go
ejVAmTcdiVKz9KWM8KKnX7dC5Xu4atWHj52XCSZB/vzhyzte319dDRPmt7rqsJHgwpb0fWf9GuP8
7LSReexBtV44tRTlc9fD9Fx8YzvEE7CFyy/E8ZpUE1ufRVSaWtrOmhqI4X0eRBdYYWyFWL3Ymaw4
cbj4RZrNqZHZN0rEK9fQm3UjWmtYfpOzI4IbJpmP7pACTKp6VTo2eKdXNeM6NXDCLghhbu3EN3c6
2nqQoXhEvFyrAdRYr8ZRvLXxIzkWFq8FAng2AY/JSwAAVO0afMJzNqutiRPaa9BU4pgYwo65GIff
1wJQdFUCwUiFFZgZypU+4KiE+h6pN5tS4lk7UD3hfXQHq80X1pQGFTe5mXFiJDoRnOlAAwtXt/Ug
QNGdQIgNNHCzeb1HgScMuzqdpgdz7mBuEOblIjXTKohsbLrcAQWDWa59cvBLUyFoVFIRPc3s0QyN
9LB/D+mDyW4DbBVUgLW0PmkWlxZuzSKL+nFkcJ4xtZsLxlp3pINIvzKTCrz0DkzGbNQlFRXy3qYy
yUV1vyzO7P0dGAp77t/i+zoPLfPgT/EkFDQDk9j8ydlOtdzzOz3HdKEb3RSmm2huhUmneJc9ipZp
qgt1sIyGnbKYc8tSNJYttQWAkQ5NQP6tu8Dgm5pYkn+SIWy/s09wPaAYMQO9CBJYkgX6/COPoh7m
ybiRWrPq5hVdLPQz57S6g7AytCbbSMiJseq5dM7Y+Z5V5o8vSf4h79FU25zGblomu3UYu1/Xr4pL
mjNuE1M8dYubAksqFBtPHghNrhFdS7Sci2pFbbnEW3WIxG7Ck7pFT/Jho+Ql/9DE0Edx1XUh2sLs
kp+l3kieYzwT3Iv5UBTA72Fy5ejMTQCnxPLuhRld9SssIFKDY2Nsj3lUwBPduXXks9jRPXCrOHri
KSPBzRyef1zF98gIztWurLrypc2YefW9pQpJWvakpDAv2tSKYbFeFeTdRfzpALPEHcyffQgiAu94
uwejS/gd8lEghc6a1XTFg7uY6yB/FzmZisX8JsWhVDqfXKTXhsKfcm3gmdu44lGBeGwQl57E1psv
Vob1N/SFYTvIO+gSFeO9/LQCFIDod5qz8S5UCAjSl+5djKa8qbjZrAWHRVMzRONtQ9cRbs7cZ+GN
clPseFWPHXlpWXqxYpE8jk7eEmp7t7Zi+Ip7rloID+HXL5zTVo5R5ci4vyrGFwk32BbXAz0Zkr3L
3Wzo/8rJ7RLv770MzDYfiFC9qVziZa3UsMWWFq5An3gU6Of+9RuOf2Iw6sqauL3JMsrcXJJ4hTR5
wJJgm7y4qKhh4SiEAtF4dG3Hlr3q0Y1znZw1g4V+h7rTA3eW9lKEedDRELUBnF9JpPO7Ptlo16or
tPEf7/jjOXGEumcbhvT0ineOz0Dih8h+N3ZD2tZkVWbAjNlz2SxAES8iTjM9+/caH7TEZDaTA0K9
DsxLmEEw+sJWa/pExuBNoOqUqHSoUiWFulaL61XcdWkchjb4o1/Ai1PXrgIsDDbuEOs8mEbEIynK
8nBGZ388EV5UtGcXCEuYtig9UGDv37rFGcZ83Cj+Q2HsWrA7vz2VHVkZeAFZMJ6qiZb+f3mcOuCq
5pUsALM+ajiWgPPmlPSKCuQNw6D3HBbEJ54Fiv3tQqhrz48Wg3ajVhl/pcNr1VWn/81rSf/+OXOz
NJiUn2Rx0NPk7WkWnBdxnjjtCoNl8vJCRNk4jdXU1q7A82BdeWgIEyZ7Ez0r/1qlduR+qMie4Mr/
hBNCW0igL4A7klYBG1vAl17wchzBAvn8hBrgtzDIKW+KLQDdOijvuclj9ZKBn2Bbn8yO297djJe2
U5T2qjf3LzLc+V1kGynHOOQGJ9Qyzw3UtGFKgNMEogFzMCwMan2bSTMnES5bhJJz7/aE24xI5twv
egzpbhLZpT8dGaNWqIBpR+/FneKCRqrkPxXKef9TPGmKVFXyfhQ62uoeFlIc0qhQBnJc+prw2o2l
Yt9jya3KZtdduEMckWrvKDCsmX7fiP0f2qKBRb4n6t+dZwI2ExhLP6CFsYW68mEAhYK7/ifXOls1
Bb57C8Hn7/C9gR9kU1S4civEmpii3DGmfxo2cXVw5mM8rXjdG+LYpMSXVZnxNyFgg0G9nRvXygVc
1XEe5FnIgxY2vIA9LmpqgfeDPawhMpnGUeYR2fCy+qEg7zNFnmBAizjRw+1Ocyv7gXVdbb4n0rhL
R1WJgk1fzz3AKz8cM5QikpeHtrcFkE+cfLwfpr1OQwfXhNCXXuqF5Qpj9Zt2AvEo1JQRkOyM9OxZ
8hr6ojI022ch22X6n/QwR25GFp3ce0tTpIwZGojz2OLlYQsYcmAsAxVCuu/4HwvwuQQKsq5TLyYw
IZvN/esp/W5BYWVvkuYSWff+tiX4HI0IRYmNDe+c2Psi3aREaScnnonMg0QUGMbsj9uJLNLaNefe
Aja+BZ2VegNaBDlgkG8BIZgvx/cVsDpoKIHPuT3nLtCkv0MK3R+VMz9fY/NJKTuR/vKChEQM3uyQ
mFHGlD2kBwuREr+sWZzOSOh552NSzKPW//AyoIKTb71mZImv/ZnSqEo3G7bKcqkudAW6D6xIpy3l
oMsWRo0OBA+/Xo0UW83NRnB38dMUqQreMmD9XHi6LbhdLI1KpTmw8tfcEDZFljYwVCf1NBX0NsR/
/n5LnN7nqo9Q1w7AFJsy6wpCm8c04GZgpssmooXrVpyDDrg9blsioqPZG1HHujFZVmHLex08xhfx
TnkcRc6yNEJrplyBUQirzilfaZpQUXjfj64nT4uG++uv0W1KMuKb+c6GNu3VSHnCqzzcnMn7SPzo
8vQNFWuzSVjHQ6Z+vjRUNrDiBju00jXzErmH2QlxsPoGXMeTMrMPl0chw7JRjU+SpyhvDoSIkrvE
e7HTkUolazenbFrb5gawcv2V4LUKG9NQIlE/seoaLJgPiAa5dpSifpaEduKGzGUztd1YNLiORiRQ
LRADoz3j2o87WLSkWAulOhS3KChdSFRdNAmrOrjNIpxjvHI+6oPfmqBE5wp4Yy1XjaVttAwLtuLP
+cHc/B9Kg1qnU+NGRbjShgSL+k6w4UiR8+GTW7puD/WeykI/xFfdQsPvz7zydtNVOIbOb7Tzmd2C
CQcLbANg819HlmpBd4Ivp5FLl/ncLJtxt9tXfOctEpLWYkjy1qf5VLcp1T+ziJYUGFtP/+5iBdAz
S2mAqu81rUYXyKXX1inUhXlocG6lcLLvS12RfACrFEaIQWMzD5KR5nv2re8pvCPh0kSsJMSdkYgh
RFzml1M5cJkGu+EsjsOy+l+cVQ3xaqkg7jcbad/N1LE8U2YDFs6rJ/ey8A6oQAelfnQ9ZIJKjMTT
ZlllQZwPK+pXx2gzzKAQXYLahV1/3dwR/+Qf2bGsiYkx4nYBFpyDlDwkrpi76g+PAWJg8oBhNrQG
mTRBcs5U5TSb8ESzOAY0U9P7YbhzFLF89lNeVdnpE8Qm5lj2Cz46g5XEcbYKpYbZx44RrwkG0wOM
SxRr8J4YOUjGUA8PbhSshVOBIc89nl/o+wIoY5iqGzYoP2W7lCSn+aauPc3c65FUQmQ8Qsk8wr7K
o8NdCYKP+cA3yj5zNV3NXQUoaEFcbZG3KRiXYrYDVPozII8CP5cMyJ6Rl1LAxUCSm5gMkFn8v7RI
py0QS2VVFLNV8y00m3Iv+gScoIen/0y/6G4arOXWVHNa5Ahisq/d23yTjyFyeUH82MmF3KyWzXGN
flOXxU15Py2Z73AfwamfK5yXA4KL+yY9IUV7Hsto4/ndaBMQ6IKKE+9MbqJUEP/lAiacoEetY0+8
QpI/CeEH/yLm23BKLnKz+0of2JzAd4Hd50KhTuYv84Gtax0ayUXePthxp54jA+Y2uaUYdvjwYOeN
AbfufiKIG68fhbi3EtM0rGNKLwQcLXdRRQaOP/BVHgyrxoKhFPiW3rd+BvH86ijNc0eVwkKG9NZF
iZ3S6C6jAGwh70wCVvauHSJuHuI5JBW3EI3iaURuiS6dNAyA25MeOd7EwBPRwnNzZAj14bvMSpwh
RGx8KhsuPFyKqZRUW8V0hxTW384iZaynMDQcvBpHWYvpppnmHTBzczsXUab9I5qCn5CEDN2d1WVn
58XeYvKM3KUnIdGlRsIaYxL+yOxF67s1SnUbnMiychCn7rN2ls65xu/iY9fcK40pOZwu1F4NDoKH
X5mTfcVX7ts8fwWvgVAV2MLD1avXo1kP2OfKbuKe3aNfSnQBIfQoQbdviJbg2oGsNHmGO7TbZwUE
r/a5GRN7sejSNKcXZ+DQVzGiab8GxScUm595kckm1AGY9Soa66gliWjlRoQQhXtKqMYu3HTJl4TK
fsrmTTEwxp3UGYyzCsn7kLISmrRT9TN10LvL6Cnx3Cqo6IT8jviUkpF8fH8eAzSSK1kmRX8si/BC
mOTR9o7I0YximVy2bhJodkEwynta0NfwMjUIXZbHhDZrnYGk/c2n1Zo2nhYNoomUHKi049xorNNf
XVdjF+ZSqluetppV4+8Cg7l1NY8a3okG3Rn8fCyihIM5HaMC+dXqSq4yhvjhWIsVMxwwVEZ0U2vE
lusbbR9XuivUyqY3p5qe5/cS2QluFGQ8mS86vrGjaHyz4k0SxJgHE2kVgfOacXGmSMpbvPdyAVN5
qF+V18fGpdijzbqhpMGJPmSuAtyDUCzD3hcaqbg+OowJBTrmEaOtPkPCVkRJdonfKEYLDJ9fCfH9
6qVOLedZvtsnJ5Tn5Q/pZNyuBA6aX660MBI/Hg6jiBu5zxS1gIN2HmMHDAhc2Qa1Oc6/xm2d3Bvl
WxcYqfNcta0Mg45OqjRlN08uTeVfQ8KsfQ/hRgdLjj4ad1vTti9G1ESkw8zmOzZfwLXtXTivMm0+
rwnGQTuDC18KQhIPqMW/vvip3rcSPm5rS0TZ+Mj+xME4E/k7ZzCYW0YrQqk/g2n5DcC3gWPN1yut
LrcJrBGl1KAMymVMMBoWpPbLjj6hdveAYnVAFVkQKoAxgGJ3Y/Qw4oKqcwlSMo4Cjbuh7H9TUg5j
wNPlCumr34ia9CIAjp9m/CospgSz/BuwqNxooQifZfh2DqihUTFntLnSGXD6fCDGauJwg21o1X4x
bvHTW8W47awDiDFbIVu9WY8yFTcWUqWtlGwaHdrdgnyqfyzuIQqIiDIgJ89K4wQF5YQfbRGxXiWB
W15k4yko9Gjd0ohMqzwfYvupjoQCYefFXzgdLrQI0fdDcL2shIEjxrWiPmrvPwBHCHcreATrJ2au
dm7EJQ9DYU+ROGgOfaYTstcw7BZUG3RK+u2GCc1f9jLOimXwWkCU9RJecJNdKkmo2HYq46RDocSL
tIxERllaIm+c3A2aNe89RePfQ8uLMer7m4qqRTFzDMMemJMLfqzRLYbOTzplvY7X3hfxm0X5RBaa
syiOeb8Iu5pjXPqDCbjeKq4ogk/XCGpKoQlVFBc/Pn9NZE9+InPgQe9zZLdZcX8Z4q630zEdKnuj
7TuvMB8YVi9Dzltj+XDhxXocOsx0vCOhGUjbaiXC9jw89Wy/XS/wIWbGshq+kG5eoZMmQgXwuNH2
QvgAzuNYs1jBC/c8L4JBiei2+vd0lRGmCJSsK/Du75Ytq3Z5ixy5Od2oYdeikZO9BBRpICK2mKlX
71MPPfSjP9RnpFmgw8NI1+kaUoHL5k0XM4gI4PygIcRwjnJu1ofpiAgNIOqS7rSfD+ZkP/nYPUOo
l9yRD4qqXqpxRuQkUMXX9CgMDraWDS8AWPaKimBifhK81A+r9cbIk0JhEQNY5ARj2QNTAKBhH0u6
In+qSxjxemO1SXabyM45wNZVT+NiHMZuBFOKlcspkhmkjwAgbBf24TJ+kFcSR+9gEdLuBkt2jAwD
EO3+dyqPg9iJMSVIH9cKbg83H8t6ZD4R8GInbIye53adVXTVyJ3zCyEc6T0US3267u46l17V1fIK
Tcu7qbjWDLGvov0RzD8i+++QU2giSFZltRiCrrsM+Ibb1nKFSw1FLvu3XPWjz7c17lLGYK2YfLLO
dzHE1g9nS//epurtJ7Bwk2MOVgYisIHWqwa6PCZ7wuSaZQGuEPGNoimld4RVa4rEa8FNUIGTg06P
jf5dW2NPHlYocvI3nY7CQ2A6T3KTLyhvf/wLz1uT1ObTYctQq7/2TLxGWqo2GBs18i1IpqhcMXAG
kYpzzT92kj1jSv33VWleZnsOAg0Pf8X/sXh9RIgx7Rm4xW8PfeY61SYJyVCFYmZx1B8/LrxNcFiE
h2dW4jh+t0P7W5J9ZAVIsbcfMKkIbaw3sIsIh6sh0lciW05WlaxfmtfqWbRUZFlWHkFStKnTfXZL
+iYx0mJi5G2krlvz/YFuIjUn/y5rffUS3lNB2PJcdbUPd+aVr8ydBlnrkd/fxgAcENzEKxangima
7O/3aempnMm/6AHAe1RLZyaNGQseJkUnhf/dqQ9SYOFa0ya2J4CaTE6YwGOBjLgaI9Q5X6+kHsdu
T953InzVMfXjJTbsWhQGnjaF/e5EE+JAlIStwOitj1avX6Ff32YLItHEEsrcov/1WiwdJrg/rCjG
k04tBbJZj4bA+deF3revhLcbU+uzHJXDyx3l/G+NrqJ1rllaVnsNpPme+VOKafyxPgLrValJ0eS+
34Smihgfhyb3z/nqZpCIhSDPQP7Q2GM+wNtbyq1DP4kDjqKseJdUdhlr2yXRigfCCatr2J7Xzp3o
B+wzvxotxjM2mM3qKP9ElA0LdpR9pETyOF6VKDHdP7Cl1YQliHQaqW6eAW5/Af+psE0TsKoHNOSA
UUA5UBaBNwu/VVagTGpK33pRhLIf6Ny/mJzYTddb1TJaBtClh3Wpzolv6VMcMBIA7S1+Wq0QyuLX
eeXtE4LUOhrPVI8eTWgEWagBF70L8G+9e3FJlbB9YVARa+ITpdo3Y10TAvDbNfA2mx9ap6akKBQh
xfgWP1xu7FEXQVdSRwyNYcNU7M3etJx3vnyQAhaQXDPo+b9eVy36Of+BjjFqwLe9OMtTvDZXYT4u
k7uqXt2F8IpvQhQ7T3G0DrxGMhSNz9jCuhp7Wi3+Mee+qWDrRjqhz+eCQP5DNvT8g6ixKK1wkp3R
3rBpWB6LEYbvFF5cWxvXhG8oDLLz6GZAGBANN8rpdGDfNUM4cCgVQ+z6OneR3MLebUKMwygQ6PEK
lBPtPXYO+g4CI/99Vs4EO/5hAV2V6tz0LKtrU3/gaRLWhBDoJDNxjeAAnoRMBmqUfcfEhWXurRFM
V021w5VTT8OmM7YaxcAIs4Myl89ETITKQLgW8CAYQGblqlllA/IAZLoGb5a7NpnhZpUrsBJiYq92
Boy/CuRJOQfwTPwg2tbYeuBVK/21fmr2eiov+U5WUIePfDkIZ3e0YwGPidc995sk3IuqIOhFI3Gl
uPYABjPMWvNEMaRacBlv+2/ODr8bArqPs6jTyD2YFfpUBH7hsf4Q3mpTHV6FdzW7mAP3yBBoZUA/
6tR16Q4TrYRGkPCtE1h3Pu1UEuTCXlJ/7G+HLtfNmC1AvM2DQ2GRLfHZzZNlwvQhkHFp3fOzgzr1
EXKSeqT6L/AJgOQ+ewtSMZk8myNmj+3YKDqv9n9zrAHsIMmtMIvuthkLr5S4dp3cFfYu2QL7EsdT
Xy50WYF84BB5HkWMqmyXeduM8GnWii26ZGNuJpSnA+O+Sng0uYETjOYmQPVQoG+DtX36ecCiBnQw
HfpMEJBJ+XNu1a6fecFQ02gVRussvkuJ99f490ZOPIxgn3j7S6m2Z2w6EeKwGBbWc2cLqQklAGCs
LUDmPrS89oiKHkF30w8h1Iny+PNJPvvtcLUy4EVsLdsiidd5D03Bzcx1SfdCb+5bKWjcKIv3PpR8
E58OCCZyOdy+doIhD3k05jklnceKLwIEaFzQdRWRX7GUQ82sC83X3XDyCxZ9r6OysRbQcGivafEF
Jri+F1oDj5acUC+ASd97yiQUxOrT2S4r/dJS2WM85wnRPwcQYeoeBeo5Apd/A3RckDkuSSK7kdfc
TtpRzvS7NNCWgU0Tm3Npkpo+ggUmzcfucq8dZiY1VnMjH3cs+vFH9zDS0GkvxZpFZC0iKd4xliyy
xxBfkmamrilYcPNGfheJfzKdBOnMvjPzVeFX5TT3sXoApoD6IOnotzc8e5RByKP1BSLSijQCtetz
vfUnPLH0OKnvSu+Ma1jsbBSVWMpTPYO3rKrrTpsm4MsRQg4UIWgzB6ilZ4lQiiFg5unxWi0CV7yb
SKZ5iPJgc+fleyXFkwxcyIN5ZGDqlobVhYj7P6Mjww2VqyNlZIb/sj7U/dPRx6xK6g+FcJnuKs+j
nxTRJhbbciAV7nnlpcokish5q+Xh2AB8Xtm+pEkyJMe3fsa5jvxPaPwwd9psM927uuVl8AhvusLF
qjLnxB4I+vqaP5Yd0851IWVjeegjEFE8jZRAWJvLu4u/db1DKbHMmF3+fxZs7hzz8dptpfNYJe2B
ioqX1S/LO27eNNvfCQLpcqbZx+vaxO8JQJKK/6NaODo40LYVnhPqebE0swI5oGGmTzsek3qZgO34
1JUq0entuR47XiwRRoLNSVZUg/UG6m4keQd1qaevJynplMO3F5mN6G1NinhvWZuglFi8PprFQBLY
Lh9iZUCG+gF5KkFnKavuEa+sLTTfWjIdObyz5Wd+FVFsbDgd//Q8fjF5LauYQ+i2m1rEyOFHstgZ
lRm5Hg4hQaHw4WDK7GCRNN42VOBPUqjC7oQtS4qARd1g8bnn2IrFgqni4bGHGMtRanJbbDByS3sR
Jl3ND1hHkjDzABxZqheF5/fMHwHU/kYLECPAlH55IyE/N+5CsJB9fUsgj0lsCyHjTMOe6v/UmuED
/yJGV7qBg0gU96qanRREyxNnse9gYPSvAK/SBDEqiXGeeHo4uayiPn4jD7MjYdzgTiu/4XavfvlA
wATNGEk3aIjYYWV6QRcKBgOFJe9iwsvd/hEuGBbE387csV6ufV9SiqsD+Cv4Wripw0bpZfNSZRWK
0ZHdmkkGUtlURLcvq/ZHdLmPvUK3dI54EF6lZeH+JcxTD54ZZl5DqOd7/XIksK3mwd0RAbVwE2c8
kiLE7Eh2t5jgUFuGCuDcb13emBHnLC274oaksOlr44deDjG77IbaVjnN79azRG8GnxGZpSjrd+/I
7fxK4zB2pnGyCho2Zn/yfqrHSDbmt5Y7TqwGpM+SSzCSsdt/yhuuMBeRs0FlqinUQ/lZDrPB6uXg
yZXKIoe8u93vNeW4S42HoM+58tVpW2jaZ6stUyl5kVmcCJPB0ixroo5rFpAh6KZMyfxstoPLpoqY
khHEI0IQiqPuhC9pd0+i4Eu2eLdto7YlrJDkAXiLUX527gLWABt9d/mtVmL2UMqPQ9DYfqJoIREm
AlWKGi62Qfuy0VIxKsz/nac39ZN121D7XhjeFqxxTRYmmUfkJgS33S+t7ZJjazmTgdJtwCBVqAbg
wi1OOhXXYRjX/n5Y3xhmrO04rFUMPtDar26HzfAIs+gaLD2qI7gJsqrc2grMVEldn3mvEtgQ/yXd
cbWXVAY7mLAcad7QH1qZlONOdQ8IUtObUfGT7MgI9l2t6cUkGjznM7NGLdKyqFBR3cgfDdB0dY/g
hSnAylrbjVvMAYrySW/VQ0egQl/Hn2Fd6ehcZbGNy3kXpiEsgc2ztLZiI5scw4h6VmffAzbIXBaQ
RNWCEhk7lrVHxZfEnj8HctwGDZZ4sE9wQGvtNVNoqXVDeujHANLR280lFu71T3ua7ajkcBEiHjIN
tCUkOQYui+l2lU2vb4D0TOEQVKD7SFiy9MYjvK+FqPrmMX3zGbzaD0eqRzMgQP0j4IYiZeJu4qmn
pmNVgYCXbjpQorHO9nIHk7T3gh0EpnQK7BOWOmKXU/qVsZkShfbyJa/AWv6MhrRk9BxT2hbwBtsj
gehdraNLi/HpECrPn84agwGVWNxuznZ+eJmdG0aAUhU9swDBhTbQdhSsWPEywnqMXJwH9BLOUSkf
BRubsaN5ibfBUVf9TcdQLjxJWzjhnGb1FM9s09l0sXSQZ2y1o6DpzoWdR/TjYAhGcIWXXqwe2082
g1TFeER3nNpw7yX1hugc8eB0+xKv99LgpQHtX8O6zM+XCYtkCiA6yvg22W/XkKEN9aGPgGN0XUs/
kHxI6SYrb7YLkWPPOWAaJkhe0niZXUQ0dTqnXuhnvAo4bTzLxn94tGPUefED/DwNc+tUcAvckUhY
RTuJJW2iSk2UGERYiCR1mfT3tWwDHuhejABe86QqzkKOs6W3wv4Nd8QS4mqkAZBfswsWYYTm/vyZ
JyKvyGVr3fGh6Zbl9bLg7ga+me2EZeAnND746i5HGBxjdGKpn0JFJZzbNLoHSVI/90F5WE+Pvwi3
xyCrHiV8HLohVo2l9PixFk5y2p9dvRbAg+TJkupHWEfFJwsGAiHGQn/Jgn18ENH0bckMBJNiEVus
wFtWXvvb1jp95gSABns47jH2fYc51n+m8PKu0ECY7In/nCPn+xf67DV5ri+gscDofxXN3eJ98kE7
pD7oceC+35LgLRcAyS1ysQQqb8xAOlXpieB3SUk3517udS/azlXCZwKecrM7Y0QKeFDcw1zg7HMX
Po//r8K2ZpR5jaHtPrFDIO+iotU9M6gOb2pRnDpdb9zwic9iPNxRPu1T1JGY514KURJEJXiwEfMB
WCPwaTpvsvPun3H0dAPe4jdP7ilbFcMJg+q2eaEXJoByqSlywEjL6gTngg+Kc9HRD6AOccUrffYS
jJgYajB8emUCFdWqgeRlBliROW1VwiW3LemLvoYHPvqyLRkrRORkXVmqhxB270iyZ1JVAVMZB2F1
cHrXD6VF8wzUozMGPZkYzNzxJZlHeuiOmDASCQsZHi0mfK76nqSZBZ7I4nJm9KRIwVw6XbLPaFRh
/fxPwSL1kp0cjA7a5MJ37iC059qsrebEUvrXkhoILLqwIp8fa/ynDIOW8Un6tLblaKObbRVvpPGx
GKS12rUuGOcifhKQLk8G5wyzhAfQx6v7FUQibKvqTYraMwmpgdOVZOTjL/e12FbEL01Xwl16v7Hy
txJc83awmqWtwRWv5t2v1mMx4vPLx96ESu5vam6byf9xpkEz587sFPTgWOQx808lmJwa4PZmwtpx
d7DesPYhbkD3KHbGBFo9D/eAx1+rQyV2suYHv4vsdDYlocAyrYsTLGX0EptDTAfXm5pDdZg1mOIZ
BxD7TmwhJXvdVD85c/PgiAYC/oJRE2lq/hPm6dVF0uYwNO7AEN9EA2EzRi0BAO7xmUqi3w8OvuzM
je8I4WCf+oLwpTnR8tPtKvUmK7KAjsjXkvFhqeimfKtD3Cw+ys8/VQ6dvPiaS05ACpS/FoTmfYXH
HKPZECxO0VB7gapQhZC7/M+SSmdzmCv5KL7N0XHZasIO9JNcpysgHU4B+rYKvzXToy2wd5kLt14C
xdpIp9HNomOk432P1OLpOaQdBFExVofTWyWOHSN/WoKvwav+upWT+YpbEsA71fJHzcPrGCcmZaG2
Fk5UYarVUf6ElefvFqlhX3h0Uz1tMyDrDCtvdQ7/UbB5A5UfvzYKkPuCyvUrM2GnYTJaosaU/Txl
x9e8kMmjjSXl+ufTir3yLnVCNRbxwOt6v5NBCQNOK8jYgGTOp45704kjTzK4xUQ6blFGT3bftUT5
P9kWosikV67Kcb0YbxZZpb9TKf0oNbdTdt0VQUn3uPli6ChmdxnUk8Wb6uvPmVwn9b/Xe76Z8xTi
3l8q6gqb5xU20owhfgySLTblxkQ3kbnFpuO+hu1FdnBrfktzazj/+ZqLqQWzg6mKPlLW+emdURo9
HQKkFJFgjF6jliCQsNaS+upksRXy/NJeyE07Szv/OtPpn3Mp7mYyfh22o4In2SX67cIR87WiDVrx
Aoj4phEsPWSsjApWIXMOqmUam5XvtKAzOqkpX61W/dxKP3kB84zMwRZ8r7nrQw03QoIG7cFZ9lCV
e24/ag2hWQLRw3p/0Ea9B4BJM/gCvNC3lDnCGHTXeLxiu1/ptwI1JBRNBLI4MSQgTpTsQ/ztQzpl
bPEWNruIUKhFRkexGzPSOKAZ9YkWflFzRZCs49XsIcSKZ6ipqXXHW8KwrGEV8XTGnLz9Q4rj7wiQ
i/R+DphQkDZEnfMdGqCboUDEhr7VwSBGXypeKh8iNQWyycbd/cN5yMQ3SodKDxFOPeMQ8SavDCjA
Hhph/FX+441adP7RMh8ESI4Wvn/wz/uYda3VrnIEBqKqRpeyr0oddrtbGpMJeHPsayuogPfkcZ4D
RMspIZg1app0sEfhz1rQv9p/bhaYWQ4TuYtlkqt74EXGn2dewRszF5anwPQsxyoIFKKfeIr8XBl8
dhFMigIJBkxua3+fzvCtRJSL+NcgwBogBNaE6dRkn0lNlK2RLMwO764DoUUUCsvQneKbFsFO3OUZ
KM/adS/YKMCo6Jz7KI2NaU9ZBv06fbcLWLq83lVF+eNbsUBejCF1tIVHCeFBjVdvKmT4z4rQ4xrb
Y5xUEayLubjOxBBwFatdQMi4ZMNyjTNf0Latub69/nIXLOQ0dTNc9AH8R1bHuNKHWjzIc3u8ljh7
OSpudK1w5+km/tUTGG3BrQY8MQ474JblaGBmxwi18DlHfwLzVt8xTAwHch6g10ZwxxxwNw9+aGxj
YE7r801okzLK98OuPvgcnH/t7cYnaEHbKF0Sj7V4g2OgtQhQsALJEFiE+YA8fHl6jd5H2YugcyWF
cnQ9yLlPqGafMsdNO8WPedlGy/pR8EngUuJp4jDY7oVq0CezdEv1AaVBlF3g5NFjJeDMty0vWNI8
Rk4lCC0Klp/DcaaWt5WBPm46cawWdo41hRujEOofinV5Xh+A0j4PSfw1dC/poIP1o1b7MYpdGoEN
HUbxpy0Jf1NEGICiu8A8O+1eyLP+8pJGGFhGW/T6OFJ6LyTENPj7HhdiCOI5DwIy3628y/wbhSn8
5Fved7fdGeOfgfZNo+KzI4C4ZC4K/9ZYE5gqi70KGlqVx6QtHhNP0Canob8VFguTYyMeWv6Z8WFS
SftsVeeSoZ0adZsWHnfAy+EEhZzgHn3Lx9HyCFaNg4A+j2Xky+MmILwk6tRifYjNmH5ubBQzGa1t
RVU5o3qQr1CVkG6ZfQv6VjYyxlb3l3/dSh2vg7/3FPG264+Y8fN2XWNPKrOUmPJyTAFtv+9nK5HA
B3Nyw3C4p+rBOYF58h+cK3qkFi+JU0wCaHgHI9C3hw8ZVW2mjSpjp5MSvILP3gk+ckXTXsn5Z32n
fK2fL9KzU6oaz1l0CxSCoFLIgGqABO8hwLah/vf1fwV90Gzy6tciEeI8xZ28zGeKxtOH0UVBYAyO
iJBMgjMdpxaXvpI0ZKMxL7M1OzVvSvu4YhUC6Tw6Uk4CsNuZAzQWFhOs6/Ejcprk9N3CE2PMYkAT
J1zh1OZpceurKguypwL7CriK/f1NHTxKruisR4ya1NjAbw7UN1QGx/HABLTKg6xVW5sH339rPr+t
iKV3R7mhi/4XbiTDMgq1UEJlC1OdOBoc+7JtC1pjTzm4mpazNtzUUYWWqR4sbKwenXFgIGtMldKI
np4TDu7A1pgKU1dTjtb78+kFjyoQrmsn/h3JgLOA9NNOp34Lw4wsQ+gZSFtt+PrfSlutWPbfXAsE
9KLAWNzlerMR/QomjKHL/5x6QG4ZDd+ieTXn+ga1X2dl07B7QzAyeFdHMCl7VuPA1JsDXqNd/yCi
qXxiZ/+b3II2kcXlaUWHbghordH3FTz0gtpKAhEo3GiaEqZpgn7dSNsIUIwV+kIIpYQgpJB9IUS9
7GBJ3q5i0eBRabXonSJVFcvn2PPK5PqavYlbf2c3GjChqAPHIwZCokampxeQxJFqA7Yjtf46VbFr
m4i61692dVnil2VRCcqp0qpVwwLEPYYcX1DKdbTdCVUxfrRD54fZRSKaGdf+4R9EuY8LHnT9N/GW
B/HalkPONRfCXamvOuJoF0AzFthM443D5P4IHgu+Sj1rOGgxzZjtRGZWL9xfFY+1khdtIstyUlcU
G9tf1Kbp9iff5BqajmvrY/HRsBRLHU1/JeMlE0LgKN9z+FBKxDDuTEQwFLMP9Bdyk0/n/YHWTVX2
NpVz4xT+GZxaJ2MhxEq7fvFKmXTl9a39LuSr/0cPaWlK5sSMrl4F5g71U2EOOmTRQoTKA8JqUbbL
1qWeOecgEz/fp4kRroGbnxrhtafk3LCHhFnbdcIAwytGz6uJDsBQrJuoSHwurfUKZBZ+/B0WaklZ
/a6L+pZN5nOKa0UxVAGuo5ApDw5xx97kKD+WBcWnSiILJzCk3BXGwTBkGDbp1BQlCI5eE0Jx/vp7
T+bjyJwJ2F4ANFLHAg0OlUgS2LmwYEiT7Emu4sU8KZjLxkIn1pZ5WaJxSjNTQ7rd83MSReWxhsbM
fM9fmb9Vka2SVouuIgL8aGdW+V5OD1FnjRYrXy/qxldUAO1AFKOu8LtED4qpFQJcoCTMcG49+pLh
RizE3MnSYPg+PFA8ulLuG6uQ0p34oapWv0EmlwvNX1YuSYKdGcqZq4bTFJzaISvl48oSDh2KiE1i
tkep0aPkflP31ben60BCXorcnImZYh/eT1ji9oz3XUkZQyNrJzLSxyqxYUUktcQIhK8jKRKdUiPm
3mhKKa+eztscsCpdUtDCWLBwGFAI/d93ZPqzKUuB2RjoF3icJFKAFanQBQU5yR5BCnN9n4VO5zY2
mRtI50c5iSo7RmGrxBK5Kfk7Ism2yAWU7HqWcsWlzAyn9dtW00DpFyc3XwKQcKM7OwUy48PfaFZv
Xy5lKaaMrtkalSFWRIIZ7b3s98cp1wvmaAqKG+53AF6Xrk8VmqPzzJx5cKt1NeKPW1xW+CS6MYFY
iaeKmR5NepB9+MV3E6wNwCYCg3rjWeREdEyBlbxI9q5sTyyTDc2yh8YC8U6/j2cqNVyKeSVdIeWd
G8/x/tgoFHvAnl0SaTq6h9RR/abyykLa8YjGS6EmsfkvyXCPiCaeQbTD27oLObUWOo1oKk+rpwEK
AlLQZdWwTunvnmY10jQvlHs0LGwBkIGxpVzCVflJTaSF/9Q8V+ogcJXCxQfPVcrJP4NVwsIm4C7Q
P43ca1KMu3/hAMMfB3tyNRJICuewzVMIJLBGmOjvZd8oYBGBJwq/z50gwGBEaNCTH3E/3yyJ/piT
WZzKMepZTq9HkKu3D3T/KIwFXEWWSlNf8+ngeQj69EzzosHFt3gOXYGrZa+sx0srphycbePO1ok1
umbfMZSGUHcfdVfd4C9Fsccery04jphU/l7Vm54nnz8YhgX9nLwMLr622u6v6yKRyJ5FManv5Y+7
YA5ijRK9S4fZ05ikuMgMoX9Xc+WuMsecGJ2CrS1jsG6ciFzUO2+7xMyERenxOGxURmj31vQhp4SA
ki+jIGE2R/Y2WnqBWGiGHBhm04oO/Im9nfGD1rcHCrgc44RZ69ABLjL/mdEiiJ6VsSzouutRF2+R
6vNPIOLEqnVhTtLNxq+50thPQSg2btAp6QasfwiKOCDZ+di5c6B6mK39urs6Y+geR3foIjdqH1CT
YH3jIJYV6p4QTXcAONCzp/aBvfp6PXBBe5ErfLhtAaBC/boQJTclvB3KkJrBpTJzx28c4mm/Niwj
lJev4G9BMZl4fQcom9XIuTIhap6fiyg0pI2gOG/AH4h5Rqu4+0/1kXvjtz8EpPprPwhbaz6AtkN9
H31pkQFjRRrKF9yX8327IpRK6lcHu131iqAm4+paxlVt2p2Lazkx5bqnLrv6wGJ1xIlxCJAfZh8k
EEwv2p54kl/qfEShJuH+2Oz3sBYrZj8YyfL4ExD4+C/qD93jkQv2PIUrranYlPYpFyVnJONaZbzx
tADDiax9R9gqg26TW6DfrgvpX+DRu36iHi7C3L0DSqYD/0H1DoigfbzVdj9SegTr5bGXjpS1EDuB
qZbsJipFm87qowfgJSysQvN00bnkjVvDllVVe6IqCxL9cuaSQ9rKSPrwl7Oa9NK2kJXjl8r4dKCC
BWbpWLzZO3Fw7YrHE45lpKAA94LXsJHMj9GNBXJHXjOB2BYC2tOv2vfHUDngj3Y/meMhk+QxoaJN
654nEAn0bCzQxi9zdgOC2HU0NQvEeahBvKQ5YSJAbSCyQzkcS+HR6NGcHrRlOzZQ2gxYfIeM7vhd
RPMXSc7GeWhB1OmutxaVC2/EcEQM8bCvMrNqNh0+/0Ht6Eg2IYaBvsBj/1wwrHfcRrf7cbcityQ1
4PPn3aigBuy1sC5iuSa/prg8AbggmBd+LcR5ZwTWH2UhDLPTp/1hKbthvoO9mF4J1y3S94zkbIWC
+xWbAET54Lg/iTZKanfly6DSGU8584zAeJTfo+jtoE2gB31G+MgvyUDzNOip3xsnEvuQvRMsO8vy
LQ/CHC0nLMT08DyBHE0+71ssGzKzph5rvMGGg7qwcu+VTqfditgzgqwIBl2/3Z5M3LUu6LrdNEZJ
2kZ6o/5octncrZnadm46JbZzn7HVWY7ieastvT76pZ/Eeq9sllZfvVn8z1dODAef8i5MVAw+ZOx5
T+HeTLEFfAFt3ibI8WLUA1H3/GWgvZkUPyGrWHWzSdip1BIKq9v05vYCMvyRVBZmE8XSegWXUZpw
QslKJhlLcuU5cKsG5VAD75A4KYuWSp79vAXSpgei0xlStR3AG0tF2LSEX8QbFZFXUwS2iMQUnwjU
pDjb/lA265IPHI6sMt/Esqdk6Gq1yvV5Go6X/OdEEPiWNoKYhxHCKm+gHYX8y6R1AOzuJnnBez0t
zxpr5YVTUPEkk09ncY0E/zWzAxQhK4GSpOrvq3y1M1Q03Gp76MA2942LR3vsHoh4BuXqw1x3tEuM
0oMYj+fBZ95Ej+so1eHiVSNYz/NYlq5eyJFDeEeLieXQHHfpyTUgTNAyjiu+tN+OAxFHpelZApLm
bOrelr2HGL5lSddfpsGZ+etED+qw2x6iUqrxPpLfVLE7u1yfXvnQiOtPIugwwRe0tL4GcdsWw0Wp
/QrzZ24cYp2AvGSbc7xuCmwLYlIYx6GMXjgF+hymczJ6NJylWhUzG9+a5mHPrewN7GFdTEiNQOK5
uikuotj0SpoNDAooKB3VHEtg9uiy8f0cFq0QC2XIiwlTvVlyTCIl7yGbjHbuQLiWlnxy8lUBUs/t
RsjqVy4cDHBE+FcCc26CWkjDt1q3U9LbGXqaYyKCWhm+j2HgAkuLMaYEt+/eypmS3kOxrptbkDaU
n1uZhpDASl0o7CupNI3NXG50wux3zdbiLtdYFY0llyhTs3nO4ic5x8/1mVEnitU04IIUdDsmta2W
DQ/+1aDeCMKDqF/Q187ylgCzz/ZIPzvJTTLxMyGjXS4B6woYkHMaKbwZRtkQ0Q2o4/eg+1Fo0d0b
1H2iJpovCkInSMUagecRRfeJWBtq3k4pzrYN4WTh3cCsHruw6YqK8j8qrBuX/qlEKnCEukhvrTqw
Ub+R4d/MaheRN4og8uSHYwzDhPzTVpKIZmlGJkfZN2NXqRQTjgCXZQfwcfGmq2loGohIWsE8zMFt
Eig5SDJqt1L1WuqAM02ZUYbdVKlvZu+n4tRfBs4ymw+cUingB5qXEPlPr+L7U0X/pcs/Jz+DQ4fZ
L9U/qYGKK5XqQERgvEE7yCbse978G4neCHXDHErqfTbmYD5FeAFdZx5rn3BjvJuPCCDjverBLwXv
bduSv9R438plkQqZMhynGzzVwS5qq5uC8efG+2CPf0pA9DY4wQ5vG+DapB4HlMUKAXPLWIm/aO0C
M+YWKLWHMcFhWs3D3drJyJ5tAx1iOsxdub/b4MXTwyuV3YgZqytMjMtEr+MhWpp8PjmBpg4yTE6C
n56d6uHQAhBLA+n6ue2X32FfTLhVEY3Hetx9IVoduAICHv06kB8wjq0BERoonS/idX/Lof4O8DJ/
2fRaAKU8rtjE77wV7JI0d7r6pL5pqipAAzqpeMIcJ+GIjRdCRNtFA2WJ2a/3lUs0Q73RcG4dIoPh
8hRqm85OOlFZ7P951F7MW0z2KW1Eyqr6dbX+6YizZT2U6e3dRcefM2KlcTmYLBKjIvr3whnKhFL9
FWobq49inUpFMiFHiiyj7ruQF+eoO+CqNRqJyJVicSGxOSChDqx03BScaMjF9LNUFq0y6KW2g8rN
nc58RvBqtJl+xzx00rQjBW3K4QgyYOioDM6g1GAa7bwVGwLBlmapJ8EuzZrHYqfSvfy/dXIkPorf
jTEBVu7Ca1NAt7mil7D0HkdnDm7Pjrg5hV7GoPVHCs7gBpxjJmxTl4tHaIN0+6W0SZY2FBJgUiGo
LlDVv2OY3XmbfNgEekqS3SOzHftz60jmR+yIRJt3Smr48jfVu4HkmHt9YyI7LhVBDHEr0AbuKtXJ
ysztm8scPCQp2qUykicEKbR97IbsJjfsIdhKCkmuTc7RgE1bltHGYwhz7Nw1LDAbUMKF4Y5YXCkj
4+1kcRcrboeVgJ/JcWTWB6ueOheb1BxIMs9au3VpUGozJzi76LAd4KxMqQiEW5MWzMrOdAC3v5Xo
mVoL4uGfTdFfAV7MqZY+AwxZSugG55Hr8HQP8R1MQZs9JIFXmCtPjotR9hF7k5iK5xLnZN4Mdpp+
2/92WoK8dswnwirRZ1otUByK4Rv/74QAHvoVX9WfXXzjxR9lsgEjprx5dtlHmhq8jedKeyqzxhZh
Icp/jiLQaoPk1qmuaeMzvVFPNE80Ie8+/dXB7XQk/ECr/hSL1kkYh+QTTPuTDzPQbtU8X4EEp+Rq
pO2CjBBlx76dul/jERAzHVYAlj64eZHSdgqzqElTMhkXCdQddfzhykuBmRbrNsX1bzeSawitEejk
vPQ+TZhBDAppOIjaHw9sRaPo3HPmKJ2KI8XrfYnbWw7/zFTknUfwJbkJ14ZjoEe2oAR7LV0CZ80P
ubjvh88ct/c0ugvR53E5vw68e4XOlw4JKxhcMvAQIgJhHqhM9inUz91lxLD5eRqTagu8eyvag/Jw
rNVbq/q+wsazzvcTzOdWyZpUeS8Q8NQMZONRhl6Bj9KO4+uUEksC6LlQdZQC7y6dC9bFwHvu4L3R
cO1aCEHwUEgPPScLJmn6pq+YoQ6iywe2Yr+if/wZvHTfOdzo5rkICR2elz+pX1XkJln80o/IWIM=
`pragma protect end_protected

// 
