/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
bc4WnAkqx6dlMsl5fn3cAprcqqxHUHgVY/ImIQQum+cRAB7ouhGGGf7iFZf77q22uZ5IUqV83Quw
Hyk2hoLyHV1tsHXgJxRTk+FG0z8kNO9UiseME5aOM/+f1fcoxpdwoF5Nb9O6O9ouJZW/9wU+cOBn
deDxs8Fe2cl/gc7w+7aUoFn4WojygKnIaeby9NCvgShnH90A/5GxWomjUdPAdBRy04fmF471qpG3
rcDSX8G6arFIKQEh5UwVCLxQIuBK6e0cztUh2ocE1tgu0ybaWCTYOjp5wNkYHxW0TxCBiXthO/Y0
21pIqRWTmcspQgDYTjUBBMfo4xnplJBqhrkXZQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="ASJKkguRF7cNZtn0GfYOwaRh6RbIlcvsA1oAuucVfb8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 307280)
`pragma protect data_block
Xy3DKr6jQ6T4G9Vc1bujRtqniuPlr6GpHKueZJ5VKCbUfUEp+gyDprEx2xCJ2KwthNgRxy+62Tje
quj+Hu6xkrUM3z2T5gfrcD+kb11v0J51Xel6CnpwLVAhblGmhWHLkq8gjbSK5B7yiStZ0P4Sfsrx
/bvGqbL7Qw8Lhu0Og+A5opUL9OwnNil9HL2yQpHG5QJonFwztvBQ7m9OTbR8lYHDRt5oCj+nluKg
O0rFt5K0x4chkcrMTMoAtUghfSP1ZLzcBtg9G3UZNKY4O6VSQbvBYGU9w/JmtBfRAOZENi8OL5G0
0ek6fo+OYmNen26V+5vuhJ8tTVdT60WonVU+XsvzamcygAPBJFQbCqdlm3Kf14NSJyyWB6vIFpBZ
nG+2lLm7cUoaACbfXw7LExU1YID0MNNlbtnCoZCtlrP9k5gdWEjvQtegnDe8NdbMHvjoUjGsrEsD
g9AUAtq3Fqlu0bYW117CLbJ0IJ+/3YmjINaiDaskTewqCThtC2fVv2c2S7e9PwHKR4XXtSsYLAD/
FNUXdwL3p6p4Khp53Vb3owqiMiqtI/EV9AruNgE519D5OuEdJh7AH9DIyf5G5oKlzKbv4eg+wspx
Mu0h/J3E3siYiZ3jRB1SCJxabvxVn/Y3qZYk3kYBVpLhnBm13v0MugSNFHPje1yJlPvabbESUYf3
Iox4YJzvV9IO05kD/3XpA9iCTkZcY81oQRqUjjpFYmqMYnPBBv0H2QfKsDotcOm0J4V1/wegbps1
CCPQeJnSQkGJlgl0SjcdmvxPqxyXLEPuGoAuPHzokHWPd0Nm51ZiXV0UHWraZhIlzjc6lsTp08dj
liEn+pmUltUs9yb9mxi8dlhHHpPfY9mqg5859IpFBHwufBB5+BXYQZZzHE3WagwRSDF0vfABBpdn
6OpOTePMYlwdRRjUFw6JAjzBtQIT+ho4mN2zW8ON+jXrmpnDYVMoN8D5NqjXooK9Hnfx1JCVix43
Ej6BuyFVCPtt3Uu3thwxEgjsXEY/WozUo9col4e1z9QXtQi0t0n9pr+dL41hyO52beniZufv/HMX
uEs1uHuSdcso4mOoconkl5aM8QJvO53LzJC8Ulr2dl9SV5ibb+u38REgo2e6RiY/0fKsWMrGaUJE
poQ7s6jWHYJKfeQc7L/aQ74PASObTDoemdaTVYbVgOtQLZQe4zWAV6mvi/YNvSjCxURz3st2xhHN
OKYhAa6bCr2QX2EKr4vy6f90paG7GNPPmJbezoPHDNQoSvL9Rtdcm4wnBXDbT+KKjq7LXtYsqmp3
pMlS7sY2IvnN8KGeycT24Yw6giG76pdZcokmRIDV0dMBQH7Lt83ZEDhz6QPna2Yhqft1kHEZTu6g
ntUTOl+jX9XVtepL1zEUTAc5p1JRd2dmrHlBX0KWIO/ShSJEc7vsza71SsWJKo8e2NuUPZ7zgYZs
Vi+N7NMjyPoapbsgnlNTkbdXU8SsDtryiZaZLL3wJCtvqFENIlsAuQAelCxxZYJ0m6wOzV9SHhf2
egn0GY7mh9xKXnNtDx3/zHuZiLtRYVuIt2OAjDwm6lpw6E+hqJaFDqwJSZ3Dhng3qdQ2OXfXCkQW
gOW31rEWWyV0giLYOvR/NJSyi5l+KXQe/NvlmeBaTY9AEA2dsOHa6aMHCzb4DsMwFbZgEZnS+PKQ
33z2TBRLzCSNLDFtA0ZhRPOIasl00ARImNIvtKLtmebxJCb9or+CwoM2qLJW3XvI7YtMSBLig0vp
vK2cIR2DjBsqSyaiLD1Pry2vZkjc7EHeCC1o12oLTJJ6LU3Cw9QZaMkUidnRM6qDsKkDC1Mr6GdW
JKbmN4HlETXUG8U+LX3Pb5zL4XnXqVyS/YnPSAkHdwQQltGJ2HxXl+gvAqj5XxNrnbJOcnLnR3Gn
WvPnZMMuiIW7SFY1TfnS4k806L7SHIgPuV0RKeVjkMuDt5fFFksG2DGb3FSQqgeUE6ny6xDFEXme
EwQASWRTiMcqcNSFDl34CN7M0MeuvLpsep57oAdBq3NswniN4cbDGawiENLQ7DKwvaRT+SwU+/b8
99TPDSfrJTSWllM7nhronhQ/NbxnN2LVzmb8J5q1SH14a/GnwBEx0nu3P7Jqaf6u+4klTgmqTsHC
Lx8tpM4riBJzXj5pZg2HEscHOnxLx15f6uC7fbqdWbujTVrBJV7sTRVTGGFsuOYC4/dz3M2mHQeM
ciONhNINsq+gpKAvvzSem+PhFmM5vxlnINYGGtoYxH3XkbYLyTrcapP5Dc2NLmT5byKx3fSerj+E
6KjVxSpgpe49y4b2hizx+3DX44wmxA9vVW7spBpAxiLn60Cuc6/Lzl6JG5gZoeULTpmOXQQPLMCk
iyjKSxGea64n8TFidgw1AzItI3aFguF5qbNr95dfQtbMVO7HnYSNQ/r9kpqN1d2k6ajmRR/ExNAL
CWpUnk9LBw+9QTNk/HwWkZANp56oOQMbcE7ZQ+yqSei3NkWTpgYYfr4bBkwA7LSyzI8zTRPtMZTg
eUR4lYJRgV6WagFND3nE+nPHP415+jU6mBlFo8oDhs0nKUN+d0mOlaV/irMQmBgQNeA+Iv/Vp5M/
734p+Jg+GcZBD2RGrcfW8GCI9dWX1X4sHGW04aRlKUu/wRDZpj72p8fonKPzn5WKTSIVpe3T2PWO
tDh2Hr+y1ZI/bgJinm/noVZf8kt6ErABK0KUE9cocCxoOjCVei2n3yqgDPMZl+TB8IH4/ljxObLz
ZgxehDjMoi4apg5/fGXo5/PYBDtrUMRotS+H6sLNZYIGOXjY2NveR3YMnixe8jsZaohPNddlXesS
E1d/UQ3zAzuopbXDDQakZzPACDfYaa3wG+5Tv3Fb0M/cBQQw4JzVVBANc9m7pFljK9OiWOi0rLPm
XXGtI3GHcsmu0dvBm8JbVluryDdiG5YsJyCkdFB9hla+bl3l9JWVGulqUcfSy3mv6I5yNVQQtx9e
YHj+zw2lgPBZbxe8Z9RR7sQ9fCiXwMCdUSVAnMm8SMRizhI5MOn28uQF1U742ARxMLEVZbNtxPv3
aH0jRKvdgivFvGYJhWdSJ9VWI8fjJLJbaUiiIQ6yTPX9/O/Trop5WdmyErkR0hazo1STrLgJGRwq
6ZXs7n6xtb+qxAPUWpA9dFU4ERn5dG+JEk2GbWPCTXntd4A0uAz4HIECwWUXplnQdJZWYZOw0lm/
E6agfhmBV2hP+Xzxq+TVg00PDk2fI1tMJaB9JrXKuQaXeSS/4WvCL6Gw/fMZn4txF+9tdC4TL+/v
3wPS+12NMu5B2W7PKlb2Z5gpF19/TIoXW8paFey7+eqYCIQcj533agRIz2cNNJux7Ebh8DODJacv
SO2LgFhb5tA5tdplpW56tfdETpec1n/lkuB1ZHjrIko/0w2ysy2Qi3GXisuJ3cAISjhvedpVxlvH
sN658ov8I6/vxZWEhLV4dwmBHb+nUS5BM5zvyhZoXRINwU9QplTs5S+uT2QaI83yvjIYPxZHySBj
9Aox+Q0ZQ9Zrd/dEivM9oIc8Am0m3PrVrvgTduK8QoKK+ro9Cc3xLy/lTy/ucH5bgb/weXnIpvXZ
/AwrsAzwe4ziuuViSip7MK2P0knyo2FemPBm5o/W+Qmu2WLM6eQHosjUd/RwIYOQkN2KJf8eqdaK
Yt3nxUYYBqvtZ1er9TJeHXiHqZxpfVTcQRwL6zXFfQsDSGnqTNlSIfAArii0YXlWOpTTstjy3iSu
z75oJvGISbEEXR3fj/KphOeactQD6VwwMn3Ip8oLqZjX1j/K4vz70+SCdoBaCSyDKkdVcu0MhkcR
+0wRqrOmGmteTsMbsTLZHzUeAf1BP6wwiOXS1htPVj7yu8kSDByAkYbPF8wvsVg1U1yl2lA8UQk8
CZCucz3AZ5i/yToYxQ6qQ+YEfeTZE5CQhtBW6ziGi9EnTfpNVPrPrA+zsaPKWq8mS6zsFo/wIjWK
DmLfGuSSfSFaLCUibHO0IFpowhoogJv5O3PDKZgAckSIXpzoMYnaP0q9YLqjr/3+rebl3mW8j590
Ry4SUz7Cd52hCSXPL6LmbBbtsI9m841DD/xqb2nojw5vhFTYe+TtbbJVHL/p/brTySuf232wcuss
RUwW/GMkf0mPk/lilUvq4ujp/LNVoB476vzh/RiUXUxLGUXm6jbt4FQkBhVjjhvSAJ2Y6Bn7PiH5
LUJClpL8bFCfJ7/iP2hGbPVBbgSs6EPW84iOw1HOfgFpvDHnARsV2mKnjrJkBpdrDNua9PkH0qQ1
ef782J6liFnYVMFyspvHradv+gyRjRXOLf5F14H9lM6rkkdQ+EmlnPnmdAwhEu/Vqx4CUD+yfGQG
C+6sXPoexUOaX2NxplnWhAZnU/rBfTL2gEKZjAZzb7wwAl8iA5IP9az18Tf+vqDjWmsjk4aYniDw
A5u5YPMSXNrUB1BcfsYXmjzh1U/VLrTBSOSEmYLpbnEFCvOwKDDwb+qB9MqwtVKb138T2xDhROE9
FktUsBT9D7CnOnm/ENQZyeG9jNmqrq0Cp3OydHL6NGeo9M9v42YkJfWORkbqEm36WFXH/8dIRcmG
bDXkO3m+e6K9MriP+C4gPPZ8JSKXjbMpUoIx6Np/7dYvKJ9fTOBKXBQIHczi2wTX2hwvfxCIiF4O
k/5AKTC1bmibypNFEF0hOLSqEnl+1UdcFbkfniCwOyr5LYJgjdBBj5KUGWorCBBLM8qIibsPB6Rc
caNvR8qHkWeyBXdJNIgOLIAYc9E8logznLLDn/gHDRl19g3ZsodJRvF87ZGSEhZjKWeZMTI38T6i
835lgWNfizEG6zlpNBcpcAeVJbSUFc72p9Jr7wGAJrx+dpA1NMg0ocNf9yuIwl+spRpg1oXegJ2Q
LVHrWq+M6IGgMSJ0YHSho648SKkgHi+QwPGMFTHENfp/UYfrMZcJhCJC5XDm6nke5gt0PuhH3oNH
L77cWdVhY7YM5lWgyd5UiGTovraj6s7l7XzSvusyT7a/iGGv5FZyF8JMgArOUE3JH7pz1hep0rJE
sDRkaY4RlDRcU+1Qe1uYg8HAtaTyhuTw7pbWv79BRMusfedKGB4t2q+2VYeNsmp2xFZKJzv5DHQd
cadZc+eAQpQ50K6D+NXwYl8fA+S2Vqa6x28XSkzWAW/kKBzXSkqezAau/0PX5e1s3HnsB+lyM7Zp
EH6ck5W6DlgPkY7wuJNzxVqOB/gHsmqmNBUV4X2ECXWayfuCppyXF62+teey9xWeaMlkOFhzdJ4H
Ijbm5hu6zr0DDh1OJWbS8K0wgwP2006sbLw7I7DPyv/K6lZ7lEwTDvl7YE1ASUHs7WlqfYSs3exB
cMm3M+0VcLNDDFNsVRjR7NnnfIP4uzOmA6/LkGHshhXby/fMtfGlos8PIjBH/wv3gbslJVQoXSMd
jOhxGEKG3KZyeCoZvrkski45VjRz19pIbEILPtN5X7MMl0Hsy09GtxshmO3sV5OWAQ9gF+emGnl8
2HEDUti5fvREgl3OL9CMgg4qQcqYJl6nmi1BYzKc8hD+xHiBt2sUGLUMIpXyO+gc/4SG3e3UsNpe
1yGtMRduptw8rnprzypBpmluugRE/SdW6Bgyk5Ko75HBxn6FDarMJLfNj0bjJI5R52cMRVMFxzBA
Jl/uaxAe+DCUw+UzYoirJ+Zyh0QTaUzuFx1eNQmZiw3DacYRIzkOcljAVXNdR9cbzJdYpo5ZJOBq
1a07/LohWYHBzilbI6hRTB5farb+giIkLK0WwP8I6ISGSLkYug+EmK7kBmFQDl/oYVqmxV4shVo6
Mx5IUNBmth87TZg+4W+cZ3H2+ktB65/QE8tn8h5uS89VhgJnYrnfjsqxoDlTykhB5VOuxkzpGKip
tbSUZsxiI18jql1OU6E9cGBM/wafrLr4RhtqmZe8enPqt91yXnuTIejGdYr7r4zuaqpa774kEptV
QQ6QNo3xhhzItNbe5LUiwOL+1r0ytbShcxO7RbGf3MQHD719azngpg21LYezxdsjy8Hzgr2Cmj2p
8O2PIDCfAOWchu+LTppc+GzBRRZb6+o0GLla0lZnl5xmaUBx/WzI8Mfe57sf0mFrUVHxu08C87uJ
uAlgUVtaoA7nBbbx2E0qQJZeu1qh0dh9SRfZsqRzkaihcpgDY4NDJUz7G1tPwmG5GQMQLFbMSt5n
8DMs9HaDnF/hk3LMr0+fK1m30BWhU71QpA1Ju8lm8nklyPd8iuBdMcpbH9xstMB1gOoiGKOIGEBs
3KZaNaZh95vtsO1s0/N1Kip9jYTc8Bgo0XDKLyOM5YiSAzBv8U+Sa2vxeHrE86H5C3sIUbdN52Eu
WMDpWm6QI8IKwjY28l+GOf9KpakR9z641caKSDmq77hAbFDoJPD02oHt4siRNnrIx0z/xO+/9ujI
rBy3XRliPe2fMvZbDqMT+iAX4BA+05/pPapaj9lbS4u87XoWERjIhIUX77qH45KJ6JZVrv/GhkNU
RALIyPTHVo7dH4ISRkaDOKX6AdrS/4bi0IWFTzZKZDoEYmZobJ0D2inoh7TSWiBTvplD7guiWYK0
cxP59KCtaRlQpHnRe1+I08hKjWRO1Wa24iZJEDGHjDqTYnpVOkJ5A8YOvAyuxRLtzRmAbXaejaBH
Bs8fDhYMExEDG+xWuC56B7PR024uYQFxFOCyrdV5PLUZBPzsU16q3ApcTz3M6yRUUL0AfHBrglYP
hOePdgNYcDVapVltjFn8xwRqV4KGRdSyNtGdIgUnwy2AdYlNNGKb8ww+COD0za9UhOvn+ogRSvaA
mCNno69RPWLcG1S/kJTyBBXA9S+Xp+MQUrAgsRnyJOQSqtvnMCr3AFw+jQIFLwmh6lespsRgv6u7
06XQXH7r1LBgFK9QAhAZWGh1fqYx/mqkio/kqTpEfh/Zz80L/Ry2mavhv5AcE5qkTlpSqIT/M12f
iXKLCel9uzZBv9+fya2e6O02Mbo1qAqWoawh4quJ7UeYoQyzy2pLSG0ldDsfCSJxGWFx1UIWIULN
mAPmsGyyHDm1RMvSdaqdk+2DqA68whCBTQ6l+ucq0Q+Mp0TvbyoHUMWn4uDDS4/xwsTMJ2D1iVqX
x585Di8LBZNv1uRsiqaJtGzvMVGSwjuIUIJYTgM498JOcs/A2HyC/RAL0y1CpIXrVxBoGUe8/AVP
3/szz7+suD1bjE4yXJ8aZyyGLbTdROQmOAf73UC7Yg1/6bdApFzK2eY4+wcPC99O2q0SUCDN3WNc
ZYqxlT/+eDcf3SVHpq3YYHjoPdRMzRSuTZ+5aTcPlSMfxKuP6bdNsKWODI5ulEcwCjmrLH/YuLyE
mwujmwp1t+9Dt5Szj6sJQWXwHsPpF/a26mPJ1MfCtzfS3Nf+m7WhIu+4G4hubvdguwnJKdwtvVqO
ulWgqIkdd5miv0HT86HiT0CGIvwT1+jMRKWoHOnYXycv7m5Yl7oR1I0BPYbGgPviOrdI+QH5k32N
D23ZKWbC89mUNG2A9M2/4chI+BQT5vHRp/zTjdosysihCPfmb1WkVboc9BfQ4OlwQJP3jvW0+XpQ
X9I5rX/RXas7eq44dRBz1M1vVzACGzs91Sl2DxGuUG2A2N+/PQbsVIhXb/ib8eZ89OJsONH3yUUr
Mc/y88gB/883DhGNd6zSvU2lK6h9/ph0Uaa/7UqfXTVkduz2CphMIT449eJ6g3KHGMltUQpYDD7p
J2U6Hlp4DvbHczJGlrc6+/nDZkUQr0Jwr0UDaC2OSWJLVPaDxTj7L1prq8NcGB4m6bYDZZ+BZd8G
KK3I2mt7yjbRCTuwAdxlLsoEEqPiDL+md/aaAvr34PFHCOxvo/1nWcBi9lAQ2KHUHrfHS1D2lUK8
5lkiX6XHOtBY+YJxhHdKzO3pa6Fep2VIfJRCE+8eUU8lbmFNnh6/jDdQCGQhX8RaVuPRcNISDi0q
lQTzDiwujMS/MXkveNSOsbRPpybzctAaaXPJQvEErLzWivQA7+OJuupccFbESgVk1RJAr5Lp65UW
/78NggA58PXDzeigXzGq6y7FHtvzKM4U6WwQPLY/QSeqlvndu/AXQn/Lf9XtUHxOwvpvpidRGLQ2
HmdSlGNTEtWOMdPcpp7h+D2JO3pS0FXzeTXm07Iji1bv+/MpZ8Hb66G7za3LoGmcrHucFBE0aLJx
WothznJB97NWB6BHn0MiJ4igZIOnUr4E16Mli52hfGd0fzJOq2C/2bbyMU11qFXTVskvLjyhUXXT
nvmr58HXYZ95MIzDbCY6hYuy8s/EPpL8IzMUMXyPA5i5dhUUz0R3apYRlk4RFGeojXTdA7i+yS2j
iqS88Zu8XshKJjWQ+GMTKTDHR6JLzLRt0G9zunSZRhjVj0QuA8HVn/HDK8C2lujXr9qVUmWl4Flc
HXxp2W5LMViB/R0wdvcMt6I3Z4VVPfTfoX1QmE60lkzcbAHv87DhEq3eDVMqrsiYmJjKqsdH0Fty
mLTHeMnKf/Wj52ZtRtWOeu24GwPpMbhq8p1eVU6OLtjFQEXA7oEs+nj1j8sllz/ewym1wqz+k7D/
cDQN/zHRuUaL0HN1au2ziUd6PJkDmGcxDtm8c+qZUkmWXb7oXaxu5Yt7dttZdqZgovfi/eVuUg0y
Dh4H+XvxElGP6iztj5or9nz+OigNXa9BgLEiPFa7RTRloxeQ1jopUNfa/4f1evwP8h2XUn1rGYiZ
68+jDf1LdZq2aPgenaDTqHWaIu/hHYoGKuQRuL/KreXnR0TwR/f5t+ZfheYBGEiYrIb0zna7D5MK
MznDLhgfp8Ttm4ksgoklDRaeoasoOE/FOCrMeLnkATlzpPCCNEmnWpiAGCtB79Cy1hhC3ZYvFf9U
yTz/jrUqRNzAgzMom7TB4RQoMVvz3JFUKENc4RbRdVsaFB44IrcTQSYG7DB+xALVJhdkPFDXssty
fWlCpk5gVXzUKm3x3W+qaQyuFuadN3QtCe8NdxI8J+9PbBC1Sh/kYF33MbEGb6zdTdIOHah6xoPn
f1n6bPq6vElrP4aq5SSd7G+e/I5l8s+Yisz1zj1AYUNRmcmvzzZjn6gqLHKyM1544PWPyrEtdsb0
JZB5DNLRyyrsXgcmb+omxVWwVAO/jlJNgQOixB2QOQi3ww7YK4kinM+SPshOBsv1TcfdBAwQPu49
+9pwtIJHlCnC68REa7vQKOOMXUtwS0zUuSYMh8vZhWowpezzPq8T1X9o5BOCqdyDJmhLlT4t1KET
RRxbNrtA/9zOJ05Enm2Xd/DPfFHMGHSxKV60PZghqlgD784H/SAFWskT479vTl3MDR13D+lB7MPp
qyob+Pjf/manfx6Y7pBFvGgDBplEPc94N7mPpHVP0ymU4DFqwvAtBI3Xafh5hhu3CQKRCsMBOHGX
OCDSOSOL/ImBTtwdqFCs5HYeCojvHRcRuExwTbS7OTzZY9+b2EKJaykOiEaqdvcoZpbsq/qjp+ab
lZkPp3Aq4rTJ/Nq3JoyIPrN0d5MPJSDdk2d/7dFFFHAoTIU/qVdffEOKS3VjHdIxFatoivg6oGmf
KE/VTg9J0XjFA9RhB27vYAbnahKOIM5F8t1Qv3nJHJ1Pm0psInsEMac1cqKdL/+57YLxwUx7uSTd
IF5Ggj7TUZgLGg/0nWMmqqQtw66k0rWD0BPCrDsFvD5AfwXOdpuRK+StcpfXL8Ywzt6von/BKJzm
4y6gDCnJfEHcg6uIP2J0PZr8JRVaBGXT7JUcorFCLT+U7Ub6D/4Oo7KoYJOgaBJqNwNFgjUweYAA
81CLNW6qsnpGf+6ZOqkv94z7snK6T5XDLZLW0wUJ10+ersaW/43pxYkaN4tM7AoPQX9sriyDV1Eh
pIiAeH25qN70LztcWlMf6dYohC6C0AAMwo7jpJyOU7wXqoVTN7ToOU0/xdBQVAD4479r21IeQ8rF
jYWLHgqEe2eLVPCB4D5zffU7f2LxhC/6lyixhiKNMlzCE8g14BwZMhkbL90G9V7kr6o6h1sU7EJp
J5cEy+6lgWgjOJXNbC2ROy67J0hoEKdRUcjM3m2oifQ6fN3Lqr46Z4J9bAN+kXibEcXjjYWTJd6j
6YCLq9r27kJxV0Ocq0yhl3gQnUj+1KgWDAQR4M140rwh8sZOoLZuvTWmw4ymWJ7Bj5DHKAjgBxgW
P+z9vIZO4ZKzWpC8WH0UxU7POVrC9Ulk/eJwzLOxbzRnuFEo8h6tgTCqKnx3EOubS2Ak3YgTAdNj
jgazkTcLG6Uv2OxaesvEA5zEHiXdMuatM+j+dFIX+pt0NTEyfgCSXiO3oBPpSxpeS46e2umr3aMl
nYx6Rj1mOZSvbIy+Qs+eNywZTzowaiIrIyIXISLVuAJgl8NyJIuvmZE464f1ngOhAl/4CTQm8//y
jnUZnHp6M0BDTT+8f2XKiXWG+s89HwUXsH12UsE85zRcq93RZnMWAqHwfBx4WOe8cM+JNVqyEm6c
1XNWRNqPLVQklkNY+9LOmdkcSpFWume4NVxsK/2SC4uWtB8qZRzmm2jVHxvdvBvUX2fS3zfGPF1o
1xbe0XCsiBXegMn92GQXFgCnEhfgsM8RkX9rBWhU1Lz0sk2v29vYz52bCPEX+/tlNC7NhNCl4Tvj
DdyNkwUVt0sSJDXcSmTnuJoDDcfyd9AkqZlI3NauPrbbMOvXOZJnWlkUceeujHLKq7ECjFZwNhSR
EVuRJtcEopYeSMSJwmGyO4icHzNvM8I/NwsnM8nSksLOqWwhkRJICZsw/On22YSXwlB4W2+1ZQHZ
jCmPilvVaATIr/ciCYw+csvz8RdwDRn956pk8b5zSP9ksFwTQReRF/8/zpxSoAsMaU8qtpRxvsYZ
9rfVrKktNF6vtrColr6qokNQn5EBEWhbcYByS1C0MWcgftvlh8SvfiC8BtQPdqIi6vk9JXHFB/PL
G+HVTqneP4MJ80DVFSWRcfLIQ9HdNcCq/NodeLhqh4vGpJnshU1IZsXq7mamn+wba1cAwKxY0Upw
iaXYsLjcRIfnWSjWxbfoNzm5zatdkQLL/WAQSauSDM+w7pM5eGD2uAD+TXZAlz4C05GLGj0sRcJj
c3tmlW5njJ3rPWiXQr48HLFbOm1XL2BCOilEoJBAHPw6wCqpi00VIPunfnYMP94S6M7CCES4O4LI
yn2yj9cGOpLPIEU9tC7rxUaMGL9EezBI8rsiVWIhjOstqqWx8TbXRE1KUbMWD3GD41DQvDwYSvxm
mTMZWfW1Y6sz8iUcgiSmd3tjMF9qKDP5Dq5CcbZ+lQwFIqo5fTrSkMHWP/RKfPUVjkR5VuZXl2WK
NY/Vdz3UWX8Yj7EJJCZZLNeQ2+nvYKcvRn3U9bhudUO+7AWKP+F7XB1NXOREFAHHJkLSpxVrBniZ
2Tu3uGn1TBXMavuZSwMUQU/MLXj/EASQ/WlfOgkElUj94G3+OXe/nVWKruW6w1YT9Zj3OBtz4Y8/
5k6ENgZrG1UeaxMuqs4MVY2ChxF+kprWUnbCXlUjcs1ivWRNe9dqpaGooorvATdune17wpjNLGZL
/BiAmerM1W1N3RXYDnz75q9AIoXbc9ZEtJYkew7x/Sd1Fp8tssM+zy2qQdCOI6qsrbUhAwaIiuC1
vbRgB/8+erCZbHRsmRpPIufrE+fUJitBJGxQ/svZpg5QQrBbdwD008FqdjUW/iVtooRKCY5mWTNp
SKHer9UGLs8x8fmqdKlGmp90DZFcIuTstcOpwg4GLg3/OwljRL7KlC9MCViFxpcIckv2O/lk89dv
dJlf7XCdXCuaHb1dpBUFuGxxU48xdMFUPTUSSJOP82w5g1GeifdPynwsvWCAp6mZemKJhKAEjkZl
lz4VRIKHePKQ2IMWQiDTE/l2lPANbH8imYuP3JIQAfPhQ43Y91L6hXhjUkcAMp5sakeRpXLgI/Z2
NmM49NRBV4NdbmuzPEpKf7sI8eWXI5f5m7xwRM286ORzz1uTcTZDKD15WruCUTKPdhnrbEMNkDRx
jpncCzsb6kc1BzSF+9dFoiq82PgpnmGw+dyENANNSsiTKu4w/1pNd77Do6Dw20BAauVaHlTUqVPr
jgzsHTeaAQ8rgbZiUSdetqbYuriVD3coA0oYFrsBit9RvYKMy9sv7Vm5I05B6i6odqe98TtxqKiI
eJ1Kq+wyiDCp9/DaN6odSKtefzQpm91tK2TSZ8QkiGDchusPYd288BLCr9PRcVhElcQe5abtzbL+
E0iLz1yQfZMfIZxudWfVsNnYle/axdgbl7UxfMX7goaxowXaX8NHhT/OpegExiJvK4e1oAHh3OhW
yNT6/V2GgOFZPhWUr3q5/vGvDUh7c6Rex2nAP1NqgC7LtSYwvuKDAzWWl5aQjXMp96Ts3l4kdvbI
lsgzPPRz3sV+rIxzan2r4yZAg8X3QSs/NjSFkPp7bQVlOBowILVDsD2qb0wlc310ogcFR/XW7su4
vuokX52QFTfLMzTNcALlDTKVoN7Qa27Knp8/fwykipJeaPbK90wK03ga4aLRLxP2qvFJp88IoS50
+y/RljE3dj2Pn3uNS2951C5AkJfwYKnWxXhhY92k/dC8iCDwY/XwYtp39Itgf1Nlb7hcsk03a8qW
S5s4JiO2fedv74NeC6yg9BhEfL89/XTzbLmsMeSdROySJGmscRskxv+ymzPMFTnFaeZueiJ7BXId
H8JIeVoLBaq7a62TLOeyUJGWnU2ox7AgdeeWGWjg2i3UVR2fh7Wfpjbi1xbRE2QPqICdljxDCGPO
4+J5gDjDNvBxBaeh5NDz8c3o3s5x77s7NL12+Hm8Hf6yXqDFA37GnXLVvod7EJSzwXaYBI+VpJcK
ZjHP5Igy4AJoLQUF5lhjS4erbkIORmMX0q3+BlE+jyDk8+3Yj5iAJP+iS5m8lzPxeY3Ry8osxLx2
YPtQx1wPAIrqJFKuTuGsu2na0YqhITVjqS0w2KSlT7WLxAUZ4cJUAtJ3GlLUwNqF3iRrARtMxAPl
iZZ2gUxxaTBs16ya4Q1WxL9uBMCYu9OwA+2QksXeJ9DWwYWQ+I49dnn2baw402WdpyEGedyyzloF
+b4zhSAr4RZdI/YxGLQ5NsdZqkZRzRLbtMJJAg6ny+fNH8vgUMmWnVzSdsUt8Jtohpyv3LQfFu8s
buJaiaPT2xK2eT6f17J1ZkfzmcouBS4zKVJ79Pg/9i2cUKm5bTwuD9Vo7M7u7SyNj/Q/0Dg6D3CS
UshYyCTUuEqCfbZ1Q7+829/cvG46X1EdZXbaQ7+TUD9WbwPCVXT+QNm2vQOM4jz+OHLNDK2q2Usj
hahLC7O4cA7xdG5PB839yvWBK9XM2hpGSWyDMpJ9eAaFSZhbggXvINpWz3EAzWIeZhME9wxHUnqu
/M+lz6Tb6h49IX2vAMmyFRdYdo/qVS9C3VcdMtjX3UHXJzFiWFjxtShfXqRLObFvWHP8asi1q13g
ZLGwNthH+eC4hSYNQ8FDHmbjjHejkWTwkg1PToi32j46uRTRdWhjonYnk/6dgi3JtLYIxA2iS0CB
vEgmOtyjycfypTUTD4nlMoC40ZUhCvqXJxA8IJ0Vrrwd3m6uro9FTREfO2M9hJcwTyo/Co5G356V
OoJv3lDdpeCnRs+4HuJBi4pJtz2q+v8Lh7C/94/aFg6psi6WMtaTT+IGcL1CL601ya+DtYb6OSla
Yg60rnKF1yZkpX66o/4pHGAfCgp40p1yfG63IWEG/wIKZQCuELa1lAQXMY8iGhUUPHejkWwRyzfp
5UdzuMa8JKjzmrvPzchVxG9wIBOENQzQpluNzhnyisJiLb5h4fglVlAFVSkvnHZRal0JlXFEpjfT
lLRYecsvQxqUUy9q4hWi0oTgXMeRwmRUjRqJuB9c/m3JeCPRhTjQkZwuZpL9TgChI1CfeWZDB6ua
7eyHfAuHPg+XzyfxwpxIR5Yx8so1f/N+9KtN9tYNjchGdwtwUlLb1qAmUzFQjAYccHqH0AU5NjE+
GWIcNDnrxhHQHyCih7iPIS0jZQyCJFSg5QhFXS4PdHYX2xmHj1V1drbf8Awj6EFdBC/PJwY/bIpf
ACt2lU744dTfPGX8zy7cCfhreaOoUsflRhO07Vdi69LzwVb3J25FigRocsNo4oQcdVydnSQpEiZU
RF8s9OXgiAX13esxbST2LZE/oEvn4LgRQ6c92Nx5tYQo7YYdL6wrm+UgX4dWQVUFgnIaXyG/Q+xZ
jmXTopBYEq+GVe1sVdye08FDncTRGudjoWJb/NTo/TxWys3oraBZJNPE8uaFHbJCWlmp1SdWM8wi
UK4JygPK+HPQi2XZTyS2Y3FImlX4l0LkCWmH0H5yboW7L15FnSaBjGnEngec1qlThkDjQGKT+DF3
LVbR4lMZq2kyTHa8cMbzkGWTeq1NM4yTgRaKv2uePQtgAwo/2U916fzZRauNT4x526RYQgVEKeJR
Jo6nOl8fX1yNbEFZblE4kk9C9m2lRUGxtVBiYdorP49HKyYUwQKzSjeMkbkTayKTw7xFFAt/sk8C
2zkLrLdtnnT3K+30t35aPjFfTacfKrwTRRMA7hvTrm2b1KxmIMzQBDCkoCbNeTlpETvlcUVNk3iM
kg8yYwf/uxuky9QrgBEHclNSnNsGi2kt5j/+4kGAY/JAR4n7lFcTqOkGLKSZSjbLXNy7cRqDOvv7
NCNQsq1/MUD0bTsbV1d4MlHj++aW9rm7NgJlSZXXuqrwL4o1gPgmDb4py0PtozxkJZd21IizeRY2
tJKcQEl8LREYyBvSre9lTQBcLYK+cgQqfVPFNVQ6HkWF0QbooJ2C88bSpYrwMloS62WlfetZxOX6
pY31d8h9ekKdfhpr/S1Yg1MDtwLknROBB1EZkDKNygm3GmaRkvHzfu0iRRxxlNSa/uzdkvw8/RWa
1ZhsRN0Cmzqd/92kkcHtJB+JVdoQ+hhr0KaAGZ9QLQA8kCNIxJ/7xeIRFiwDuuITmXJicUe9hulM
0wx8a8NOcSfIlePOfLblIwgqE2u+VNUTBO1SZNgZ7UODHGUUEmP3+dGln7OncI0dzajiesN82UDq
Gm06OAW++AXQ/eiC5zXAK48AT9U+AY81T253OAzVbMSCv4rF1YQXtwMK2Ghaz+CUlnJM39HNdtpe
cxJ+aamqpUmvsq7OhNOM+wGAXRTwA23N7jqIi8vRRZAkQbhWbwMryqOPAk1JcunIteRalQ6hPT4E
skhoiS9yCknRQVGO2+QStOfKQBdnvkk7BjdO6SO4othSepC15PDODrg8RrLt41yw1Ii2zpidTiuV
BWY9OgMx5GVq/dcwHgoJLIxPZEEzUt9KF9pfIdafqEJcPJmssWUuUV8OL/t5fwhv2pCQJJojV7Nn
igph8Raf8iXUor5RJ8UwcRZZr9/Yvd5j+xBCB5wx9Rze0N0dBpTX4fjdEd8ma7aR0SgKJBpfAcKC
dAgp7ljtyq2NXo7qxqdHKS/lsmDw/x/KNgyCTe6a/UZ2VyAJzWg8ig9Z6i/lZ5dyWMFrPYiMuRJZ
S9Kc5HFhbBLSDPtfaE2sL3mdiAK82akMRokF3fKOS+0tvWqiIpaKn1gtV+Mi+MkQoanop7iFzqYZ
HU6WJicubgD54JRgBD2EOjOLDjFkXMFU6DV0H1NyqmgxzsoyT3CLd9IIUXnyRE96FHW8GG0ITYiW
71UPd2ZqSVG7dkjafAgTVzSyS4VlroLsuKkOFLogG6pHMdzVWecmGthOvx72HIW1vqzs4APT+TkA
JF0mk0ssPcBNkIV0IcMVHDhN5wbs339V2ptlALGfI/dvd+xubOSfpRDIidCnzQXbJs08DWoE+qTM
Yd7B2af4+EX4S8Fn+IKer2RdVTv6vRFstc0BQasuk4Y3n49w1YAFBcVvEi56rstkxCOG3ZGOawl2
8DDpYdwaKn0O4G/FmkiA7S5uF/NTQieGhSFsrb6iqv8yZ3WDN9j7ITFgSP5tF6Y94LGB1yvqgA0w
beBCY1bjiAX8hltZRLW/cFQFCcLWK3FzBhOQZQv5JXC48o/yiBTv31ASXVv9mDMPWnIR8u0acVKD
pT6LwoJTbzEHi0Q8HUY+ub98IpUJuAEDvRY/jtuKmdquYG3qUTpyqfcglwf5PxitOLdLXD8PF1Mj
0LmzVxOnJdsQO56XElzCF1YqEr/oqbKD2/EK0oFlrrKlcY60GQghHwgnZUx1fDMuuhAR7zopt9jk
2cBoRvRBPyAGAJdpDwbRmQ0hgicZVs+yEbev/Crtn/+ucHIxknHh7qXNA1OI4mw/WCRhrAVZutaT
JCStB3yoL5AztAvhWDPj9m9AgxhRWPUsJt1T8wl5XnAzAfwkIMOfM+Aayetgh92QlRJlQ6ymtnLG
9sPbzx/dtwYH/JZXcpcc7iE6T1qQBqaUoLhsLjy0kNwEDSgg72QxbR9cIppA07CvAAMCqQ4hnfNd
akzyntHhhf0bgYAkfXI8aKGE8DWw3UU5ozmJokK62e2mmM3DdZBwGNicn2UYc3cX/hsm3zLIliY3
kkDcosJSgDyOHcTZoDhAZ4HZRAdeeNQhFMFZHpsio/fVgBy209i9giRpKjlX88Fhf/m9Sep90fHw
KqU3nC/+Cwv0THhNmrS5lVuJwK7EmEcvJ2zoQ6fkyqzzkblCYU5BB1Y1Iu3APWacO0bMiiM+j+Hk
ILdDVyg/yRotgtubYS0gVEtlMbaTvmhZIIj/hQs2y6oK3/cVvSXpoaXuoPfFY7fRORCfq8zwNnH0
v7Fa0rGFOcoYZFbMrjTjtQULcPCkwAETwWsCO6kHHJHu6ok3CsLAIzKa3R0ZYFurok8RxY/bk4bR
O14RfsYkUUEP2aRvXzYoa4lSNxH4ZWO3G1yBITh0QT4NOby2+WgMbERydqS22GFkaWh/qai90z6t
cMisGfTK5/8OAPOXpuedFI/KL2MveGu1PbWwQhCV4GUHMxInvEDkqt4tGUq7Lzqd2EmHDj6AAqky
E0O5hU1BN4oJOaDYoO+ddWAO5HcqcvtFAaEDsZRXH/3j4RH5zr+mQpdcJnhvAj0D5PQTynapcfCq
WZcnORSYOVbNVcGpObhxXw7zcXg0ZHjS1SXGODtlDNd3QcfqzYN1urpMJvmRRspf8VbfE50ighDk
59uJZSg8YroRmU6uYrNPjD+muu2Kg3oz2JUY5cZ4VEQNRNJCiE4UTknbqFwRH0FUExLTv3PhCEPK
Du6XYhM51nPIaY48MLRLiIynx9DatUWZaR8fAgR41R3iwThB2Cq+AjR2zGpaCZHdcDJNHLWrIYZ1
TC2dd3lwv9rt4OA4xGvBCKcQU7juH1NUvg8YNZwtmsVKQIlftlGYC0Lu27wKSjjaMTQdvc46qc2X
r8K66n+22zm2Yrmllr6ymWcNqCfT6/4lKaZre9sqVqQ3uuW009fkKJDuLFEKQf52jaRR3g3NWaoK
vklTz7VaVWtl1yO+Fl+WYRNMK0pywAuSYGq+lTmienWoKqUFBRB1qXvsgVWjy5BaW3B0mbSyphqX
nNsb7q7/E41PW2gZe6WUlmFvVuERVCkqgzGP93icT901tP9c3C84WA1GbE0ex+Qu4kIusrdCsA4R
sW2c+r5qJe+iwLJyV9/OIXPQq3cEn6hUhK+fBQwNCcXF78nXZ+YKFjdnAWeRd84GbwfDQy1K63cf
0wycwbhVPlFt2lVu8JlalHwLMIupHVyZv0ESEREtaoDDEaqRH8aq2I2WW94QMNpqWnznmiOt1GyX
FGRyQwb5848DTd9TZKJs7lsS3K83vV28Nu4ySBjfDz5J6JnwaQ1p/uZg1uHHJo7em5kKe3uvVi0j
iDQv86xmvLubkXhluclNnkleLLQ9+ZcMVO11Kj2nDVAiSp2LOxJC9bFH5tS0labA0pUMdjzaRhWx
WfODyMWV5bvFVnaHvNQj59+7fPzz96kQ1zsV08hLLy1x9XSrmlHZDBhmhBMdMjpQDTwsZ7iJ6PVf
+5V98feuxrtOT9y2x3Ub9Hmjn/W9DDtzxCgXIYP/EkD5sI6kE3qu4/077Hz+lVZCuEdD7djfgyy1
TRcKpOjXcz/jiSnQubaOm/0c30YC8kV1YNXdot2tvxQKER+TTLe1WhGA4pxifWOtZvx9FezNZOxk
lNqmh1PVDWpUorM1p9eVog8ZIpS6E5xNPvImwkzZw3S4gfigSIcmOlQlnrXgiaJthD4HEEp/aAt0
HeX0qGGVFih9mRknKhHAc/SOE53YBBgWW0wPF8y0H5PyZN+hZI7np/4o9579PzngjhPUci677Qlf
044d5avLX6XRW+2kxstCP8zCd+S15BXNKQOaRDFyb/WTvrcq+NzFwjmiAjJl1DRtbRRWkSxCLQ+M
fa3oayJvaOACftnPAll41eiLpdUr/UpMdQK8CD7dz1HgBS8MJxkpXA44yLeDgaMMW5t3h1kiqrYN
Lz8dHN2tLI8I9xWQiHw90I1Ak57DDF6Ua1vok+6VKH+VA1MbjQZwy0ALXN8ggbbPzrEvyzdVhKs+
NT5j0E95c8wAt17hAfiS7/ztnHV7I9IbdKcGCNlhUWqyOMR741tlx9+uGzs8dNUje0gm6SaitqZh
fmRg8xLlP5MdcbfYjZFqOvatN7jTuEWM1e9QLRiM29WwaDC/25ByspcyxTEWfiu43i6QcXgTPhJC
uFxFDQ94JbGf0g1RH8sQv+5xkhkrwxOHDM6D/YEIU/wRqCHssa8g+slKfYOExb4EFQ2ufwT4sQEg
tYXjVhyB2Wj300dvbDZVRFTlCYV+RXzpV9qbfqasRWaEke1oa0mFFgc6axLGgKcgOLfviqlQX2TA
rDlRHT5U/FssnMOgdy4JPUV/UIcSkVTGyvTkX6YWWfl54FTTdxm1yJezFGCQBTMrGuHjt9nucn0t
xqTaPJUBZmbD9nI2cJ0vldOoIVOO5tY4i0SMCjiOPrWf0AZhJUf3uSe9N3IziyI1WYMs+EuNIziW
wwlS9G6KOOKacrI+BxY/CRxPMN8odPdbtJWwwHQz++Qfg9ariwdql/jB7N3zZsD8WDVwhL+UgKd0
eqE30sNIQWPDdCSsx0OVQGCT2b4nhU85uUcXDMjxBXubLo8VLQy1+HuY0PO3hUVk3Q0iSSYw5IWO
Mmjp8qhxlJW3eZKtmeQADPLWpVNeSM/nOh/R91WgtoOBTAz5NKfi5bTqLxntxIEAEWMidvv6PMuR
WaREjaVzONuCwQWtjin2HzL/xrmfi7QkTmE+l2hbqQcOQcQtpRMRr9HNBoUZsZg1A1klCsaOvzMS
Lm8jyQbtRgEUGrl0bu4KcW6If2CV4F5T20mVoqME4/qzxII0/v9h3FxDfHlHzy/WJHg2v44XWmqC
qKvz4d9BZ5o+U7llqr0ZisdbTY/dhsaNoF6SevAkS/P3EXzUW+vyRvzWylqHbb+sRpQEJUOj0BN8
oaMVIdlLc5qsgrBplInEp4bynrtwuISteafaRMm+/4xdXlE1qRGjIaIXjKihHKq6BYZGfBYzFCdu
gNX6ksSx/GoNa6YDTuJ1HXbaZjd6g2u5/seDngICMw8WPpuM8fE0metnq7z8W5nypRhN0+XDzXqu
T9f6AljHcvk3muSkd9xhXhaNtgz49rMI6srEs4NLb8Vos8Xsa+kZ87RhHkXX4klOZsN5TSv1g6dY
rXGsjSuwM5dOTA1x5Ti4W8TfHWbSUMAJN9jXfny4d/YfhLWx2/SAKnJCyejhcThflnsktNAsemCx
gPbiw8yyAKBNQV1x/ztUZVBqn9Y1/6jbgKa91DTM16a5mP+gVoCxcieyYN0Pn3zu7RAkgGDW07gD
tcC3t7Y3yhDRY68bkWKX0i2wwft+jmdqRtDC+BDDLU5R+PqhNmfgnZfDN3fQs1Znsj0R3b7DKFY6
Memef5X13WMmQH7XXmpm14wYvqWZk1vY9/EzF9RHDDt2pnxYjGbuoLn0fjehBprI2/VOPC8Yh2rk
RnI1DMOw4k9F2aIpmdQqGTmVecGl6rcK4INKahBbCQnezQvWPC+JW8c0MTXEqX4M76MeScGieVIb
d3JAy61yErVtDVroztDZTHCuD2hhNGRxdrav+nGPzmaBCW/kEi2KIAfScit+eiO4mRuiMQ5eDV4x
FkTmwI4jEceYqWfoMzPeqldkLsAHT/mDYp5Q1+nf7hzEPJGBE0UmtHGxB1Sg+x+MEQlkb5b7Y7FA
v1Q8O+zq2usyp+F+mbvmySfchSxyZFeQCJSDElLA13VNcj7x2kcZT9cxLH1HxPtp1xYtj+tGN8gI
IRp9ftVfQ3hJ6TRCOGGxxvMKChtbVX3QK27/tkyGslE6d0tJIPPOiSUkEnnUMFN201QUpTyhO1Wb
tiQW6jBVJLOZvrnpUTpOQ1tzvysvIGQzeRuYtWSRTkC67s8cS19ZYmodcctDbmnhiiN+QFUGlrrV
Q5atxvkVtrIVv5gfcgwAMyJC9TnD+wgfk5FnqM0QJbqmRQpmJfCPNKc9pMRAvyL8/rcx1ci1BmDz
2Dj1SYdFBzQ2NgRt2y/up66rkaedMaJ4yFTs476AJgcFKPL+LoT0B1ntJHLmwmv8FuFt8wDYgWYe
7cRRjMC7Ta7TUQiyHy5hPVIfIWaQAZTCZooj3rodc3pxa00qehlWuFTMLxsiLmc9Fbe+J/ERDK75
5rcOs9dBWLwoQrX/QmJWLD3/MwkZJGkPKZetUV+m5s9TpqRN7eF+BCnLIBuKtT9Gv70v14nxmYLm
C1SgLmMOGFiw+iXOPdwPcGaJ5KKtF/uHcpV+1L0Qnw6tOKd6UhiPWAwo4MJXaPU/VECNIsVKbc5+
bhs1U/+nf8Zgy8dxPT7Jes4QOeFRVYWWWgSAntPtPaPZMDfRttWqcrQXjMLr0gI257iyojWY0NpA
rO75Jmx+JmszUADSTcS1uwCdhc7NDGrv4UdFp9zDpsywwhdXrGBQqEYJLpSS2COqkolELHShTiY+
FtnDnuAvS+GLh2Eyoerot3E+3J67OgD+eVd2eLlMraIHaoh2+bsR7S98YqNpxmQYyqH1B4BYAJGQ
pV10rfzKS6awPTRc1ShcRdmOvPJj9r3fv0PQk2/DSihkmQHReOZGn6DlTJl8VzI1n7DAEsUnlgEy
C5CC4i0S+HGLzLJU0g1BiwVqnnzctw4G+8ZXpVJ01EPdJwcha1jTxlFBAQ1EbCZSloKzl3E/kmEf
oQuJcFxuymBdZgpjjhq3vI6gU/LIHjsDFLoZgT4uzY5Qx4b7W0Yf0g8gf82/2nbQMdl65J93zUOf
u+ZuBgZQJgq6PfjozUhgqJ6jvh0yXRLqsjEUQnGuSSEEdbNCBAjnDJ0sdLLw/y5zVGxfIuxV6wiI
myuK4JmCJcotRoOi9AVPmTHXlBz/sdSvq69p2ZJstoB/8loJcK21ot/6EGvZqWH/BplqSoPJHtq+
EOykMZwSBUyEh5PE/FU61Sr30aXMs72BzfczvVNS3zU3gJYgs1MLl+ofCIfYOIqffdFgNQYwPKOM
TU/iIwJautdVEkJAKt8tNGdoj6Uifw6KDc1Vx4/8lI4vfHdNskKWs+UEbbTJimNcjQ4I9aL3kYA7
oWSg7ZCc7+AeNmoqtsgos3jL0QhbuvXFqdjbi2EeR3P9tBq75ydlIc1uLPfAq9xmotQ1ei/M89IK
ufgcaObIgLvZuaARhnMKAE/WPZYZUv5HrT3+HfepDcdPLKpm150IHnecR4+zF6bOEBl7sx4DgP7/
8Ttn74wNQ8TFxslT8B7ZFQMQy0HhShAwUZgOTfXaUiwAftw3XQ+eGOFNDdnh7nnmPDkaFQ4XaElA
KZmo0KgnYQSxfnedMjEWNWIfyTSHLbiI8tkLkOk9jmcK5G5dKiautndGO9Vvz5xrVZGboTTniz37
v0hcTX3ixLRRy7iZ+AkXGcFGlhBHIhUkRqRukI8KhJ59KWLPPZI2C7QvzocCbUhg8YI+V13Qae4D
Ser9D52ljiEtvwGH1DXILBYihHAZv4HRHixKpVuozAUeZLcxkkcRKc9mU8jk6lk8+zz1iy70dR58
OARnuOfm59YLsniNlaZ5cPGcl/1J/qa3TFEHYF2KsO934Hsc6Nca6KPh0VImaniZNM6pKxDBXZLP
PE40jgVn6EPJJDyd2ftl1SazAI3LI5+PcXkz0nfjdn9Ob04HENZL39Nxh2tb1x1o9EgTEItr2oin
PXlxS3YchtlBcCRE5oVEbiovkxLuGhTR+WbwljGWbUEvx4li09YMCti7RbOnlU1Tjn0uY+Oxbn0q
E5GkgyiPezJcrR5B9Xm86MnaZHnx9WoPcWOSI23s0IxoDU+XogayQlCPBF+LgdHAx3y+gF4PT1L8
7p9Yuir+OCqKGoOPlX5O6/QZ160557zNBA9dFFdJT5UHgZsPz1z40GH630emXr57V1h+wor9srEO
+zmHBA66jGtrONoXCbDxP80Pw+Hz7w4dhn/3IWeRWmx5JSDfCfDx5y3YZ+n9xBJF+vpRmZX6p67R
VYoCK5ugTWCwGI7e6wCudyjhvr6ZO7DOnxPWfKuB92uQT2Nq/j2ZXIP1XqSwKyIk1v419xrJHYbK
Ka9TAsB6GKXscIlDq9+zd4jmChJXW1X4SJ4n7THbx3dqe+gvHmYXLhpmXtsgt8g0r9ldaxuaaEyP
FVZw/zjWqqhyQK51Z8aTy1N8UbE9NHtowiv+t3vZLh40PJ4HWNY1U57T2MgJ1vHA3sZEhwwJ1txV
ZD5ZNFlCuqzp6ifSR+zRml5S45b6M0OCNXWOFmxlJlmGNn27uW89RMth0UZ3/B8aN19CbXMIgV5z
Hq1eX9zHWVt27bt8QTT0+nhWceTWnK36u1hacopROlPUXi8+C2rgdfukysiZa1DZeFIsvVBDz6xd
ysXJm8TdTMxnDl1LuYKmlrsc8MZo3e8k+XwMvsE2wfAj+rLLvEBvySvWh0/DSnjoNUoUAZIkmgKj
wRr7DHfwb+BXF8Vk1A7roXbDVLvAWg6Uc1NO46cfdbhyF22id2/VgrL3AadEd9nvKSAC2q2vc2R3
g6XLvwhqM7IQSYs/aHx998/uLZkcjFcFD1kz9eEab9f+H1UmcDJgvBOJcZfcW13mm4ZpNCorCyho
kyVHUI4K9YuTolt0OFWPvNrsrlzI/jeXFYSiKPVgPu5wqvMUTsIJdhq4FAeKQxfebj+nQE9/d2iF
R8SzrkSgR5jlajWSecMV5S+DcOMpUJPzhGCSulTnEOk1Ox925SYi5wj5u2WMxegKxa0SjtIAky8j
eqFif2uvcwkBAkFdwdHOaW6mYOGhzClS6fVOFH8HBgC0osnlGcS4DdTWaRMoQJJiiA7blZ93/+Bc
fMHnY/UD2Qznegbn/UlJ7regBvKq9sV0zXA773dBze/uvO8htk3VwXQ42fRSMk8r4+MuBQg2/kSG
rNUgUkuHG0le1VzJRffsAo4fVdRPfsaABj5qyZBxkcQloU8sNJ/xuvFwZcfZZ7USr35kpSgPb6ka
5c2157N+wJralPGa4slbRLJJvvKALoWatg0XpfOANs3jYc35AW5SvbnQ3MTY6tE9glrZnGOsDtL6
TwiO6+Zm9jlmX4axy6U/1VBN2g2pjzJJWc8Vb2OCYdlr/Gbc/fGMVMvM+14+WvkCKh3Su5M0nNh3
wnq39HAtvBLqqaWAeLkNyhFsrRehamkDTiAqnPhFon3cFgtNNXHIducGkd9NWAVpzcBV6NMVIeQd
qZNp4wVB7FGu7buS5ctY+yx0gDEU7itB+9TWgQKG28wb9bNuaNrZXRa8mc3gfmAk7Z7BzJ2H4uA0
mG0hj700lZGw4cQmHeA7BjhVVlwtYOpVdxavHeh9CeqHyM/tY/iiJmzXAmUCs/M1/DC1cd4iVOg+
EHdt647uToCES/Tw+js8jks9jBarKn56PbqwanqIkreFj1pykiWQDL6dfSLwUQla+huXresmOGdj
okyLTbZV3tK6a8c/D0xF3FXW1w4IPuadHcuWDnciXSn41g84lrnSwNJNosRHujYSnP0fYDO8El8i
7EPgCeuso1fBPZp1cis/+g0pLVS3bUSNNcy9GTlJtM9bvhbSdn4b1JG+3e6tN0LGHGOEN8AOTONy
dEiYy8QV0/wfMAQypqN97GQewM4KVQj3+TLAJHvCOIM/hOYbkwOCLYkmaUtAXYOefzbhAvRdUH3A
DZHPZskyxQhc4IQrVR533LIzRx2eEctpo5d5/oii6uL0Y6BF+cIKf22+S1eFsEWGTN8KLeC1k7gD
vJvqakciG9xP0Huu5o+Yjidx7YAUyBFnraBXVbApQV6GLTvbdQvdykDV99bYkIMTMbz3Ke8JCm7m
14o5n8knNAgJXSTwm+lVyOumAicO8SbRsB9lQpavDAGaThv5gC3L6ezKT6zc80DrchgL4NPCIC+h
gK3fNuk7t+SBsA6VDcbUR4PsMdl/n/xC6KQewcvLVoqk/vadqhfh8E99x14BX7k/8PZdCPoIO/En
N0yDJXtILpcCs4azbdE6/DVeS63O7KbCib6rmivSjyG7b9N1XnWXHgMNu9sooeSSrpHFLaYlQvV/
tr0REsy7OI755eUNDyaoC2JtoecboVTsyT8JAa4OnmPNn8XUgAgltiJSQwKYGlNjfdX+17Cir+jm
YezwtzBtiKlzb/ONdCUTSWO7yoouodtbxXZpimL96gylEJzcOJwru+jqjr+Gp+Xc4r7VK5d5tObP
IzTlLo9mdcf3lYkxGEgRA293t/Ct7q5kberQo3ofkej8L2cxMv91oKgki+YjS/314gQumlGg1160
+ER3vfKVPqcjj9rGQk6IJeDrrA2Cwd9B0lvdOhIwD7T2iTsrHgiLws1AGzdnOGznJgTAsxYiItlM
9LuZfgUzup639l1WvStVFU2Azg6lQZl4Ehh/Hg0zLcOXSh25KZ/Z8L9V6EBNh36oh+S0HiWlekmX
tajIUWp5QTVAYod3bmsU07FGU8/OyOkIDPWixC8iH0FI+RxAaEcbn8dXwpLW1F2MyG8+xwzO/7LJ
oBQ8ZSpjb9wfT1Bpoq8GBNeKRO7wQq72+mZYmJeO5bcOMSCIAg6+9rjB/3PiaUmtw/Czd+3Uxqj+
1ldtDjuBEuhWLgOlCRZ9cH+ufRFmO3qHvJyV6HDNSEB6odyyn84501zqKFzXR8Z6tAe8pCF17d3A
xVnzrK9/OCE84RoWuHiFBHKrZo7uoRHKbFVtPYqqdTGQBVN/boP2YqblIuI10NyTf63EWMgvMVzy
SRfJrr2qOgM/hi1JTOrhPMaQREBkdvG1HgzfqrjV8LkdpbxKE+U0asj3aj+GeoTtb9YDks0kOmVl
1V9UfPD/iLs2ZxoBdmvYmjphxeh7rvv/1Jw89aMSEdHLue4evfrml61m5u8ptSrehTJcCWP49DOI
VgYuj9KyGNBu1Jqn5R4fm1IfN3RMcw1ZuULdqzOMCKtkNEwkpVq7choSWl3oj10B01xfwEQMIsnp
Qv7oKmcjkTCb/F3rP+PwnD8e0VIwrmuYa96j0awpukd86+vPfvIlF1axj8VlB96Wyt88EJm1gWqx
49pveUuEG5vylZIwUjZcxYWs7XKqlCBrGpx5MMrtzaLLmN2vzS7h9qFUPP5dBtawpGPlx0JhRm8H
aJFEU3rlQYRA06JdobuCnMsJZWJ2T1pD+rf0lhuJEhZLZLCfa1Kk4aWbjn4oet0YcMAsgwRTgcB/
xPRfCzjqIxVHBY8k93XkI91DdUAwHVFbw/UY5Y8qI8c8Tsb8WhFyKDOSXBWC7+JCuAfUByMBxIU7
4s4Y1074wH5RqDKcoCFjiXsnt5uRGDpGITS/jJQUBRPmewV7uDAMxyHlJDfok5ZmCKlWZ4i9hl18
envCt2JV8WBr1p3Gg6VSE1aFuSTrgwMIxgiSlsiKczd543rx31UkJQfHhcy1xxysw12jHzMEvjuC
/SgygEMEZwJrgeiapVtDc7m2R9xPgKK3Fs1GtbpixpMdvGfa+u5EvTnfr3igZzxpDnkPJgQxW35X
8B95YzUb5o3bFis0kyVjuCO0uj/hen6i/1/KmHbYqBuqeDx2uHtJVodxQzqXZHK8PChlYaXhJXyy
74u+dyfwaW29kviTENHdxk4WQbh3SFUEMeRCrk1r+hxoLa1OJWm8MpQHY+AGETM4sizQN27T2MYI
LVPEbF0+Io4ZqdRUykPE/HQbMIBL6oJ6jUg9yr4gKzeU4lsLXMCOqjhsmHp6Zjq0HuPXtwPXVj6a
h6ID2qkb5v0U2CLOx1aZV+LtcwqnpixKeSvvw9wyl0iv68/XBZPkN5GWyLWdb7Va3IFstsScV8SI
4E6DiQnPAEI0cxybFCUtdQYUijmxuX90GHjIOdYJyxdSa+RQT4F5NZmDGrzQTmdXjj2lMDvszVq5
3FPQe/z9tJekN8CeXJ2qUxxw4zlBxa7YGbtNU+F6PTqGnNuYeUdXqHY/wJ3JbwKe3Im0V4HYIA7c
/uxbhEF+4DXnG9RMtWjGiWqqdy6VlIzQcFAsbI8Dm3ip5/kiylc/VqyH7Rve99JW1w/UmGK7W/rA
DoveH2hSVLjjxR0pD+ZJdUtDzg75WSjemhmVwJQqdHPrrYoqsu9jATa1UaOqYrxEKBv+j2lGNiEq
wrVsdxnkWeWdjj+LGRbAfZzXLRwJYeMntHzixYctIrCRgpLtCb4BaYeZ/vki6Y5bztxVG22v/J9u
RAfzJ2gYiLJujUG3fR4hyMhL3e0HPXswTZRMCD84QumvBUyOVOtWkPCJhnhzdnNtBT9iC6wEK10J
a6a7Cpf0jD/thR4AzMAdMQ+nwmHs4zS8VcD+X3nCLh4DBH7cTpzqaZivoZkbaY8JlqfenNuU5iTZ
prvvBh68evVyMDYXWdTwC1V6oPZ7veZ+deFF68Exf50/fn1Mlh4v5uGXsWmIJjSIGjax0VXLflYf
WlbB/15ohtfUU2xaq4Z410bVyOuX/IuF7EAO94ZW6+I0BiDq3yOT73Aa7z/An/e7LOqlHeVPXvnT
l2QNLcDWDWsqvAzp321/04gv0CYtAZoNVJUlqbXAb7HA9qW3wpw6Gx6wlkeiDgqXdqtKzxkSAiyT
PQyjlK0kSO/RcMbbeuqLSmf8jyR7TC+BYKOskmWU4Ce5o2dnlHFGPp8ycl2I8LyykAN/R9pQc4/4
ZeHIX8FhD47tGXVXidD9HEufSODVjGEAgHfuAfTgdjKiqvChrB8Z+tSyHOWlN2o+8riXJlGzSaU6
p4Lt80dtz02+Ce+L3qOspWjQDgQ7VSFY2qD8Pusg49gdkaEH2cxcd0bQNSrvQJMAYd+MikaZoUu6
FXJRtWR4vRuFrzQKwatj33ZbYw/XMhMAnb1p+I3b1hCZVSsbp6N4v008TleNiX7rok7NSlmFvyfQ
nal5BFuAkkLu2lNQTWX92+jqUZ45k1by15rHSF4+OhZfgYJ6T54tjCHg8bcJMtvvI7bqT/Gz+TG6
rV9s0GoEWkHSfzPBEjhYd4FZQPECkfG6UJ5g69Z7Ge7q9/hP7Ad4S/oyb2hkvl4Z/6VWppqoafgN
+zDgxIIMLJ+uZlcclZ/goiHKHJbjJIh0JGIs9oRqKz9Q2npnTS4l1fBkYL2XM3+ClSj3x3ffRLCu
aHDfODHjvIaAG1tx8xY/ntG+Dhk/utJtGIof4o7AoVa6PITJS05EitkejJXa3fYAimaKVfs5MbBz
t8GhLVxN/1dGXlK6wDpA5EtQr0JyzHsuZa4Zezv/8EVxqublkMLIxbKzPxS/2KXTR3uBjHPRrBHB
1F7HNVicLZx61adXSJj6ScqGao/GrJ5VY0F1PfRCOqflvsnWfzXak4Wd4btDgLMXenztp75tZMp2
6xqk08smxwsaSZULMy2dtFbvutiTydUh+dUZ8kM8x8yjatnzFtWXJIgSGYbucrBtZiDK5SUFA+RJ
G+X0+g88r6xTna7WRN4mKg3e2AK+t4WkHmRerLZPBV1zg6oyx4076WOBusI4MJR+YgPrrnhlCK1Q
cli3OwA3m+q5eWjP+DFGLYKrXOk+Y3dGfGZ+a9cj30W1Sv5gwLW5tq+7iI3ktbMzRYn/5WXFHqCQ
84m/pGJZFiBllcGz8pG8FWglEhW66nNcT8B6pGrFpscuLwGxkbIqRUUDvdK76uxoJYXuiKiQwF5V
A9nCMAnTpiSipeCheRI/Tb8RPxANHUR8HG2C9xl6+J76OdjtvaP/n0DNo2KH6APXX/g9fMF5n7SI
v8pLz3ov8NOGrDcCUu5ojSa6hGB2qOJ96xJDc2nM7wrU1nBjQpNVI3ekMER81nXcXGIdovh0/MP0
Ae0ZNGdqbDVon2FLqcOKgLtkLTO0DUWnmFNp2BX9T+I8P5mmiCgYjvZbzKHU74OM7K5xdQK4iREV
pltYMghCDchP8+pcnKv0CQMw0fxx7Ql0R0ouvY92vVQDsBQqOFGSkxDmrBuMUPI1BMdwlCXQDjMo
PxJyCsPnkcfxLPZWSto3pN/e/8yvaEz4Kk7iq9vWM2lwYXLdRa06j7AmqmM63f10n0BtjOuj0cHs
rX+XhhP9R6Fcd6YHrFPlZ1z7rKkMPb6I5CP56ItWRuvo56xzceB5m6lorSK9TensVSix1y0WjmDr
DXaPxkWvIOLim2nBiSuGquH9W4XdZ4jaObDA/+eRsDKG8L9L01aMPF1oSNTEfoiyYvVspttwdfEN
RSqnkTjy1ozKGWbyloFbJY54t6+xtQNgn/4jzl0O3iFI2NQp2vwNH0hIPWsruVoIoWQEtKzqZ6O8
3fMgtCi/ccWb6xpMiyz3JRK6jrOEUcLegel3ine9WCRcP1CJobMRr+fZwE1eILuYmYbNAHJa7Pjt
SbGE3b1mccKqxgdvrlv+DTK2/Zns0UM2tIcJJ2I6AAd52L3Dul89RvNCxvm5SOii/2jNONBqXSgy
nlFT2ZfVztZdltJZ8DMkmS5byyA+sfB1eaCNM3uiltcaxXQOrGCjyMVhX1suivP2NqT5LF2APK+/
PKNoxOuVsebgPX0UHwQmbyHho4f0oV0kHdDRbuWqHr5Hgfxz2IdsDbx36kbQgQz7w4v4uF1sNYWL
Z6HtAU2tLfn8+D5Qst91AAuw+TOKrbB8Wy+FV26PgatYGaNah2iuLhzDe1BDROhbm8R23vbi0Wvr
6vnDU3hn61bGgaNLGV9T0MThu9r8FExUuPcP6KsNkH5/jkxhaH3uiw45rmf5LCWYGCZ2JazkwSzX
nmh6obEl1efABfQbFF3wDgTwnUXo0LymqtJCX4/g3ZCyuBBO0/CgZ9xJioeELUE2Khr53HZPCsXZ
fGrDv93u2JxOsrzOWc23NXSeO7nw876ZGwy8rtAekH2/aHg/Po+7ysmq2mMdfBqsAKz+tnEmSS/7
HTYuH59a/+mM3DIRnotPnZJaKr1JTEeNsLwpWACS4WUUY+PcRNQIsHNXqKdopKeN9rjyxE9Ds2io
fYvCdaGEHEfP1VzYmkWpvuCJC9EIfE0UNfp3+Xm1OrN/0hdk3SNmsRRpT/WZKE4q78GgWKa6mvTR
kZOYiuScfV6p8zWfqn6tHCUEaih0cmgcsyW1V9g/lMUQynqpJal1fCEW4dDx1EAHI+byeIZ40ZpC
d6ewSTQ/z7QvQC2vYAFPZ9zy3wW1KPDXf0Pxd7y+cdKSJmLMEwtIfv1T3tHUHJYeirmkIBdOJWqY
+V0Ei0DOaED1f/NW5e4yZx5bD+01eF6cFlkiXYo0DHwaqLdWBYhfAFtwPngAZLAGhKz8bV41bNj3
oJRiW0UHN3mtoxURXT4KSQDIITIjxoLhFi6z+SFVrJkvbeqlVFSbx3rlrTnpoN3wj+o0dVHKtWpg
mayyh6P4MUO60s6T75bdHE5T/xrOzN/Y9ZOAhvibTgiDw1sz5Z1hBIfx0DY5DXiSxM3sYsMor8fy
vegdy5uUzLf3EnU4PkyjFrH5v3QngPZqapDEvgED3u8CyUJhDwXAkSsvAhAIEJc/CpEePJpvLOWo
AqtqG4mkbQtTB455H8ByXIBFWPBQhrAO5naMkzbDDLAKgcswjSVyYEQKTRULTR+xSRtIp2+BFsw0
8+uVMWyYlzVkkCIFrypG05C3al10vjN1RPbD8j8Lb9dJWasoEHBtxES2nisoY8OsqIkPWzFxTDy2
GMe9rmsRop7ExKPzWzOFdgtQKdANnZqf1msrbqId6SjrY8LYeOzEzVLWSTsAu1nsutg4k6YicURW
0bTBa31ve+c4hzu5pAUzQgdIQ/GkUfhstflNQlPFac9xHuiKWTC4X6oysgw9edfGafMzOVRi9Vz/
VnSFGZzPagiXx6N5xqxfqbTm3MIFTfHbNDfeX1voMBk00MbJOTcDAlW1aCKVeIN3g9uYiq+PwQFf
OYD8iIgieRrxM9Bbyzxc5NBDZaX63cnWAaZn4uH+/fF0y9X7n67SBwUQJApiu3+2YqiYxiBEKLup
Y1H4P6ASbAaAXZ90G4vlk+N6aOHQUH1397+DkaTcUv0wHGTulH+2aHR24F0fZ9LlKDLAqH4WZDdf
t1hT2vfSi1nICndhHmDeiU9WqW2Rhnc0kvRKP9PbtvgWAPjCtvf+UrU3IzI7PCQ9qdZq6EOLkXQp
ovMwdnIMxSPowjJSg+0hTi9EXlwR8BzOuXdwuGKg+gnhoRBezQM3lDCAyu7Z7Fa9GxTi7v+3Geyl
9SbES/i982cb+ulU8xGaZlsjjJ56dmMLB6VNMUeF4YbgM5do4+sqJrJ+8Z/L4y1aDNVADdYJb/c5
rdEk/fl6JHi3bLLVbODv8WL2wJBlYQGbj51R7RDf4KR/TW0H0ohQ6PBPtOV7P+D2c0HMD3pTVhZ9
GnItoIDAGgzSR/k/wIrGzNmWHNN1D09MlTwcOZWR9iNuOLeh4sNEjNUWYc79vedGF1kbkoWe6I6U
VFionIZMhUCXYuHslF00j3//AVaF4hMK4p9ziw0bwdcaLIraIvrOQ6skKJRvxip5R//b9r4wrpZG
hb4hwPiKSWRlLdYU1ZgLT4Ohlsy6KbBaems3Q01Gz2Y+jddu752QexZ8kMhKs0RB6kkE+IH8SM9D
XPNLtzRWtwbCpLznBlk9rRvaRkg8hiZS4RdpRHMc9hMGMor++K8MIo/lYLV2mTX8zSkpT2yqnGae
cyn5w+xUMo0Nb1OjAHniVW5op0CxYD2CEcwfeJ6N8nVukaBa/VHsvNTmsmXWO4Nsd5wrQFfZuQfA
/KSNWojPPTBd7JpqSNIRN3bqgVq5PHwLDZLwV9v3cf9NVEaaJfzB21vZnp0b6SZL7LWc5flJWZGi
wMqUtplye8Y0TClvYVkILuihIu9lNXVoRV7t+UhjdV9FH3M2bgt2/DS7uw6lJww2skuleUMbWAJL
9dMukqCIcfTbNASuLDbmS64+6gd9VjMWXEq9x940gk/9DfpziUMSC4TiJzwTXvFCdTiNC60a/yiq
kY0D/L4cXHetPJxxlunYUXd36ryt9MJWW26JCiDPcNh+t2xkPWtDn69mFTaL6w1bT0qHVaUYXoBI
a+42ImT7fvAScdMswzcJSvsN8/7al8A0UVKf6YlMxDp4lVodXWOe0ysCNfb0eWM/B7fcQjcmFiA1
eIpM6iLVfNhEExRfKCg5yi2/UrzEtSV+BilcABg/OxecHJ2XKF3NOHuNBlbjyBpBv8ZQXvdftLE3
YPTdPL0H2VphL/YLjD3lmUmnXSbJ96ZbycWPo8qyErhhGWFY10TwYHNEoyyj55p2Gibd7h9CIhca
nOTlbty6GLQUEqQccJcZ24kyP3zczHZwQXz84r47mwqSLAXymZDa8LYnAD+dy1DweJel5zn+icBT
jffyf5vTgl3QQf4Lw/sZ4zJQT7waZJnl4dgxDaFfTMPMawgkItjWAPD47RKkcbGs7PrZkeNym9uK
Umh/Ps5zpYHfOHtm+Dcluc68QWZyMmslBsgKV4p6Eoc8i+QoKRNXBVB1lIOcsDJ6onw9dXjCAd95
WfxFOSfK4ELB7i4YV89czDpMpcmmKiHefuwdrAZnpdHIKReL5PCdE3RUBYj+XOshNyGix3fA262j
92YBb7cwNjtlFbBt9M/LSvaYYjA2100Vfxm1KzZHyxwcdGAFZ83fqg8cy48Tfqnouk5ykSPutIGp
XV8i/B6iPntYXlvhcjbzRWVqdzRlOdvysMzkFLawWUsncRCNiFizTSmIb5DOVUhlcBU8hnDJW7f0
frjiAYKAZWBJ7tgM1iI3PW2tHaontrBmf8G2anePNzrXQAuYGkVE1gZLQOxpKc1SQZJz3cYSa1VX
yZZV3N8SpMerugm3j+1ZFAKEQuk82hij3bm6aE9Y9mk05C8f5z1ZVcIiJD4IQ14Cb69fH4coKk2a
6F+wWzi8lyJ9Jn7lcVONiNMvGuK/mPng7HFhSPOG9AlKfjT74p+/O8Nv5xOxN6fAsgtSkueqoMiH
KbFdt99c/f7wfvuL6/Kuci0aI/5qlNUqH0LUqqtTrpTDNt1SV0BCZxs5lpuuebZC3OjHWNu7b7mj
M0SrS5lZBIdmuyzC9xVUtAvsiKNc3Vh5VFGh+QlQ0RZV8qqOuLykAmhYfmFWKEASfzA2VGURVQNy
andryxaV26dSGcxK3ZOgRWCZ5/D5Wm8TIIudk2y1rXKXCwDQbB2upeu9+KObvWK/mb5Qr9+zAMFX
S++y7/qJoa8X6C5Ob0tMPcLz9+oAR8tnExVI0g1FxRKC00j6pi4N2RjlH2uuw31ZreiFMWv3PfAi
lwhqaxtkiYgYpyHYf0Pz8f01/2c80e8lsXX4f911mG/3eup+KyMVslx7TUnmg2UJH8aTyB0KVmL5
486xFZP+9cZVTcGd670GJ5oICLK4BRiZ4/9E9S1olStQolO/StOZevB/KqAYjW40m7JNBKSmJxlY
JDWIhfV6H0Jvh+dSMrl/+H7h2MDR/dMSnNhHCdnEkCLHyWCuu4dvTidJIU/EEOSWU2mzZlRgTi1E
yovFS0nCJvd1hUK0KVZ0S+aNrM31efmHbXGVIxhkt1r1VME+vUrMqpvFZWemU3dywwVTIwceLyWU
atLJi2BqfOOnRSFIJ1hcUDKSa9yD2kLdhQ+9P3LAm67kN2FjvDsIFU3KbuxzleQOd+1VS0A9+Elr
FOfnSxhSOi00mIGPOEjx/eMZtfOcNmLm0sFfYTJDFcrHziDuojaiNAD83HoAqDklEDT9rCqsTgxV
JITJnKec/Mywd+hCN1Dmy+1dOe/F5Roz12HqtSK8LJmOrqwkp5G65sOTQM1tzp63/O389/Pg0JU+
agid+Zppl8UsU/SPCZ8yEE5CfMUjdH9CzIK9KnIy6kCz52KVHcZof937tu2DLtcq/N8SaDOVnVHj
j7TRPLPZNJW053dW9EjQsIGoW0vo6GKu7zaN7qBsDmYFYIkWa0jORm93IFriqgu7HJYNuf6RttuL
0E/PI8tIYxoncRalYBwo4cONMgLU64lyCQck7XsMqg5nny0aJoV/fiyFTqat2DM6dXUUUvRfl33I
6YmKdAeRtrUo1bFo4zDFRhGEeV5E8WQJmoMvCRIpnYFP6qBgtD2rYQO2jBWJ2rdrLn8NKePIy5EI
3kmgameZiW+8CiSsRbxMouGSjjvyZVq+08OPRG6QIdCgdG4/h+PFF3tFDZdKqx8KKVROlaEjXEvF
wFBOAlldmrsOde9j3ORP5FgVyUN1veAX+ic9BrkuM6EIqDBhDqEXSJRTxMLsIt5gMsuegxxC9Ed+
o6LeCJuwmDUEAON5BUDDziEkLcPSWHhuqn17AneyF+0hkOF/PBscXwJbxYJSFvV6VfOGs9aMb2iR
pjq8iPY/y6tljgA/CdWCoP0gxQyFkz8YeLIQfFEbVBoOfJf7AFNJmlJsWqySAcVTErEbDBrga4k5
DOl1V9eLoxvMdjRM7SQWZ0001pOuDZXf+ubwXp9TTilB9OcWtXnzcAFSlxRTrjLHmwHgyW+Q3xHt
S0IvJ/vzQWDFtWe83CJDjGf6muvEUGLQ53+DY/15EFyab/sixUbz6Iitcm+/O76ExvTEjmisbtqr
XTinrcDVzY2kPgmYufQ2JA9cvGkM6lHVOkXyMcLnPkXPUKaY5bW2AZqCbWtP0F9TBeyoW36EWibv
Obbnljr4dX8ZPOFQrgmnIKq8TCpjSCzToLK5F22pcxnzTt8TBoF3YTbsoR/OWYo3WJhvjTU0wos1
kK+sGj3ITLA9lhlGfyFF4WYg2v2qRtjYtI6DRgLEY85eRFk9hM2doAeqhfcWaqRk05eW8nLoqwgA
6TuJvNE3EGHvjgZYCKymOBwFtDp0tf+SKq7xk5SzvrL6L0qT4eiMxCKZKcXJrnl79ezwmIcoEejb
YFW42Ts7OnhWs7U9mEwzWgL4sZI4pmA6IWK7xl5oh7Rwz9i+F6F2IBZ02mqRRaD/yQ2ZdXc6cIBM
RTQgZOo+qR5rErK5PKH73Njq9n41cZmBnzwezFLZQq0YPpE0gWuCqxEeZQw9Q9LgwP/1RpD/Kot8
stjDpC9j6dYeGvixYtzCwMvilfCGT4aoTurPOtSeP9DYUA4VWJTQuUIIfMxOox3WiE6HmmbiK/U8
TkNDOZTov0mZyBksku2dA7BOFcXHHxRBjzbb15VKAFDrW/j5Lr0y0xNduLexre1pZtjQS4ppWj6k
dGiAkYbheNEvgJD4FYMfT78jNEq6iX66lGvOHjcwGCr/LMEYdirPKPKNDp7gKACUAbF6NkQ9ipZI
tIU3zbsCsipN+nbsauB4v0/faw0Nng1EI6OlDjhN/UglJ4heT4o5bUX2RjhGL1C4Gs1V55H8Lcrl
l+N0W7VN6Pe0sNmAOjVMSQLVgyC13WCTVwDJP4m4ZgfErnJKD+2LUmsfgPmEmDRV1wQaAulwunOm
8xlAO0dSDwFVdidTLWnW8CN2zWpJtgG/o0RNFYyL/rgfWx2vjpHEQg3SSgdC+foVbE41Pm9Jmlyj
mGjdUK7pjBD/DL089H9qVxAO0KoY7Vntpi/xdbOFs5lXi3XNos6ZNuwvEZWGnh6sWmRc4bjedu6Z
VseDowjYX/OZ9BgdIggQfLeyrBng5gfCiioiAakDhF2HpfbCKKfID0G7R0dnU24OaruU26UKEIoL
jGLAXpL/fvVBXUxesyTJ0ummGKAIfqRNFIsusmOHynpiIBLKYE6RI7XLD7KCusfEjAn5J8GzSo+B
O4Ex5tcH9csiXO8DvsBO9p6zgszhjLHKiyq/XOhBiRb/lEPelQylbLlxP9eBl6vO9cF0xdYMEqjZ
mdwwlIYGTZgzbI6wMBnt8K6ACtpUH1/ImbbzsUcVJsUYb2NJ+bnQjVR8PXHap1y6/GvZ4EKiFmLS
a4Z4rS5h3t6YX5ryEhKYqLfg/sM9yl6pQvlUef/4UAn+glGiNyNKH7dHLAzZKW02QwaR9aA1RFsq
VHV4bKimHHP2fbrgTYfhDoRKkKK1a1VO1j7GCdj+C4iY2db5Aa2Vckw7TWGDB2x1ojoETESKkxlh
n5q8FGw6OOE5dRzCTqfwBPo75HFQNKavQqMct6m8OlYpVOm8zxufdycm0Qur2Jhvcrn+RouIBR6B
QBIzbxb8jTCJYIqtucZadHb92+ZvxA5hTgddBJ1vQUnKxc77V1C1m+5HxbIYhhIhiODMomMgJZLG
/eyg3InKtug257xK6m270xjYfdZrEsH6gDR7J/52wzkPqrQm5WvqwD/2JszjomBcpHmfp6kFUN3t
4OHMh7Tq90C8Az+Xmd7adg+ExZ5uOOz1hrjC4tvwJHHK4G8YALhyAvt/sa5RD/+TKpTXvtooEEIN
MU7CzoCh2nmZ8R3oRl5Ip4rig6tXTppbRj2M/H2kwOnrpaFr50QBp719rGq2wB0HOVvHsPXZHLtE
s41dIw3JWi+x07CZSACtVXt6Uu1m+d80aH2s8Rf6SyrJeZwierUjI2m1HXn+/aqFCXXgH0OUhAoK
yqRmPWkf7K8rM0H4086u6R7ucp71EWobjymexIOBAeUCU3Zm4eav1uojyvOVz5FziwhEdwzlq9PV
4kBK4hw7tpEiY8dgK3KTddhwXU7tBNMk+XhnfBydjGte3nDU0cuyIWGrdSwc8VoZ3wcR1EaY5hwE
XjroffLiCCr4VB8BenAS+dy0C/3psn0qVn9rmpmNoAmwzF13rB2DeKwD5CdNjM/Pni83cCo/LlFb
6dqLNlTbBMGkAtm3OW/uSjuFPBMuhPEFnXUaCfT7HPqoBNRspBZ6m4YN81xtYAvh1SWTYw7IxjpP
xELYvn91qpMSueVgCx5BoP4K9REXSUKL8yNXMGkvZlbzQtiiBbFyKLIksGsqT4N0MHXmxyADugDO
cVIZQ3PLrc+mjm4gBX7rBJpX9r7Xk9CDtsNLLJEDv/9QocT+Bqg41x+LNeEIRtyX0q3aAib7rFvH
VVAI4SBhF91xe55dYX3AhWvTwcpO6PkJBwjAZ9oGvJpn/n6rzUgwgNsFNZsDgIBsSngDk+K1gV2T
HQnJkdVkPMcsXo+S432yl1IKDqrKQuU73AEryit20MJ3EWlKa9rbrus8JJU7euM/HQCKPkAlbH8Q
QJV5hlHuX09CrvlXqP5cWvKVan5WLHtKoyB1iJnk4he1MztJ98IBziV9RgnGVF2L//swDj5QdqXL
kwZoyKFsGDsXKTNfO0ubyiPZ3D0d1N9aqDxDVfOickvoGT+J+bs6Ggo3zXuveJok57htWuCbxXBH
kas1kuIC0bN+RMO0NVPsoSaEcBRHSUvbfNcpbrvwukbAhdhFSxu2i3Mw4dbShlcDs6f9OKHIlKU0
bUHkTBNb/IeG1SpDjlESRAQhXB/DaSlabhnqXmCVPti8mKpKuN95xxVY5x67IjeJCx5RGmqSkEzD
3cct715ugiQbXpgSNNrn5PBOfZasj0QqHnkb+rx+JYYoUwSURdjq6f0wPesAPXpmkB5InJwzyymV
74/ir+wagXor+6wW38AyzP0Zn4OI3QA0hhtik7i00ap8qPL4QMcF5DGbbkhW01DGROWb+9wKfGcA
uY/6L9yzYoZ62Dyx0H8KZesJJNbhZCJWG3NqNHS3GxOHs8FM/9UWLWLih/CV+imDpCudjmpxdxra
rQcq1xaKCsRcK0vfEee5ASpV7v2mm9RnHPHn0XH+Lu1eZC+2ikUzGGR68mBbzeZRR9bkDY1j3dHH
nYo8bB5bQaMjA20uzKu+g2hOqwCXAqhoCVK687KCZwnPtnu5opn4Xqz/wt7gmglhBlJcDVzqOgZR
K/eYTckngA8Gq76Lc+nCfS5TzGi+wSONVdseDmAyjs0gU1yAMvifJ/Yc3oERCZX+jzVew+kEVQ49
gydQR9DsttUTNCOooCEZ46oSSckZrZlAGF8nz22jxHuHmh77sAPoFHRkYV90bf0ufBGmIf3L5isk
CfPu/RSF/1xmlCjkKO1dN0Vaxu6l46p3U2C7OkkQI0NATTaxAcFMXPqt1L0D4KLnQQKNkwR3faRf
euZp8t4OfJtq8WzUMTx0zFzmhm1Aiu52piKT+tJUpaKyZGa2HS/BLpVd2IiccVM+JRJw7fpMW8tp
EuxvitZ9hXr6trjLyuVi8FLkLhl0y3KqxdNevY3FJPqRTcpqFW6cD1rzOFL/3Te4DvJhfKPsFpAC
hMT/77bf7nKwnZywz3hD15Ill4gXDb2tOZ/u71WrWhSRxWY8KkwUZIrsfB2Y68F9hj0/4lYPH6fN
5UYYtfeyCrWamAvCl9WGMRr3rAdjMfo2QLs44HPHmWvGjRfkO1CaCkVPr7WcT+z4KZGsJtjJZnSy
B9/BaUnOuOHdUCtScKMhpdXh0Un6r3nzblzj1KTFz2uZOg2/H3uiTug2x9f3iLbcV88o+h8FMYEv
MR+asyeCr4cQ2KCAFQWs/R4BdeZ5W5lTkFu4RK8eo7tGJ07gD4VdWHnbRJ6glsiPZD9RGMvmXc3U
3+bzrLZYfUD6ouPsZMrSJjc230GzJw9kKtWqhzfvwXJ1aF3mcAwwZ/b3x7xanbBJE/3o3dJxk9Rq
+G/V2glXfqT7FzBS0Ytqr9luxt58seTjUAuHpnsnGDy8ZnXznqSyCVFzz5vW7nccDlGAk/qpR8vF
pduEp9txGzVj5Kyhm1EcTjPQ6UZe2n71DWsFrxPEtH4sCpPCIFDxCDPOQ6vR8v18i/7xIVs48nxk
801WD9RRBxYsnwdIee+hQp+5McFdb7xzi08z9/JlOpt2ImoY+Cmd7XodXAmtA/spgm1ssVK465QB
P9y6GtfWYFJbFl2qefVpz/TN6ujj28rus420jLmLHCq+4wkcBdapBqPwRM3lpvVrciPVQxZOv3p9
AcCH+pTlqg7GFFWbjp+rx1X27I9K99qkqxh3HL4fSttuxHy5vYdz/YhKmsoZcXDsTL2XlZc2Z06F
AFg27Uts4c4B2E0JysdoQPf5/sddYsOn69Y8llEhUNw71oXLN4s6TyHygqwVHIcvOR3semZZ7G1M
oUDUWcKgvsRxp+78Rb/yCyg20n645eb6ThBfTPyUB9MyR+hl/6HmOdgl5pPfVqPShwAS0kaWTcNL
P3Vxb3t+C8TQVDdH9SvMB8TpgXykCD4qkDUZJR/KaWEGugVOJPgkKrZSbfK/FLs2tJ7wiW3Ny3AR
yLW3WJ/tC+s7JeWgVBLZfmXDbHixKuHwkkTYy2Wg+7ySHS9RRH6FI6jwdaEMRCDiZuQ8CRjcqxeF
+KWBxLIgpPVuaV16LrQhN9kUdnllbC3jL3OM7BzfK5J9SzE9ReILgfduJHvePOqilwUDY/zn4csG
/S1eg4fvoCo6ENyei16sg4FFhtMmlWXmXwBdIL9ZLa83IRJghI9565F8j11yyjdelCApTxqUlO0a
CzJULna/ZEq9ubo+J6bJJgW4cs/XnsU1xcf25H2p8rotKTRHKEXxZFBDY4KwKbZBkIlH9Bblbhiv
RcPVRWWmGY3zGmGv9AkB/OQAsVUMAiCvhKhOSTg+7ixA7/LENXNaS96sO3QBnwQNPU/tG12Lq5Ku
mXJ6nypF5t72ga3MFyoJJVmh18ZfQJp/J1fDw8tmFScxoNdxD4UzO765qZaJalk8794ZuFluXdyw
HhYnq+YQVEJctmv486AtnP4nFulfea7VtijBRmtBPWlB6YFEwgcJhjcBUcMwBbK1lqw9zPY0BYO3
ueQkWxg+/ZbAmYvV3ju5byvAUx2nXqv3ubcJ8kYVQh2gvyv5+OQXSLaUhFHb2H08BRQVmdP9B8if
/NakEPnfcp5N07coa/hPaV0+ZS8tZedh/JfzQoLDC2Msrl7RbtGQ1zCkJRmu423eWrrhgNf8xK3t
P5nBrfDeKvX9gICZpxfndhQrYqFqx5oiv6hj//BM65kPlQ/9gFbHVAmJzwocC/YpfWoBj0sVHruG
0937MUEEcs3eZ6Aie+4qN3DunIc2RFrwmE04Jx4YCbvPhACqhKcuXbboqiRQfdqK9KE95NF5VaFI
pHLpSNcnhb6UcCYabaJv/VTmsnM9wMJJK7NvLGM0ASYU0wfWHopVDtqIJMDv14NKg/O789bzkIED
br/KwARLGUTfOXgNKzUBOA8roNsKDDvfJERRDLwy62AbHNh+6U2jtptbWEn9fy4ZNhRm8xYpGN6T
91Yj1YU+NFxq1tEyRQru4ZFS2ki8y1uXCKlAZevXHFCukZ/LwYbC8o7VSf0gIJtkFM8z1Appc4ZF
XsimFWmZf4gdovxC1jVtsn2yu115HuDA4sYEpft1dBLdSGmaviN75cQRYouMfDRMRT/H/TY2k8vM
HFQQduaZyCRlQXT3Qr388AJqI5mcpAHck1MPviv3wOdkETJij2sR7OuamCP309sPk50sfHCWu3TI
toQTbyKSeII5KuWPHslpALS3ofNYFwYFMcJ8uekqwvnO7y0fbTMJTf20Yip33jbsCcBe4I+OGts9
vVlSe28cryqEZDcUuKJOeWmSdTbRZwgktUdOwf+BBNgQozPLdi+yASR+Tna5cFfvi9XEks/MuOG4
WD1vIM6498de1Y21rjRLXlThRjVHEwEpMYoKqG0J/rKtgiEd11a9FUoN22C0hFX3w7ZVfVarzUDc
yS0cJ4RFLqb6LT62TACiNlVrP1BTOwMW6uNjr5BfB7VuO/3mBSAK4bqdZkhwEELmdjva1EcA3PFu
XU3NE1arSC5hxM8pJswmWiYGieFgMNGl4QOwes33pw+VzbfWsFpP0BSOQHeCNV3pQwbm3G84e8tw
l3z49hecNrQl1OFHTG5R+zpx+3vv9+f2Ebw2sra8q34l+TPEtFEuesiEZP7yrg+UycPnZCMmpriN
LWR5caqR/4J8W9E4NOKn4lcwdQByIGW8mwrhgFcolaXmNu9N/E3prS/XhdwKMb/H97JRGubP/1uJ
+iNGo+qSAJnKvmyuPQTbLgP3NcU8ditpo9sJGzafx7r5YpqFrcp36DA8jz6ytw5ARFo6vcz0ijiB
j5trhZSJv3OX6KeTrNWuUz6vcYHL+rzkC0B5/u5Q3Cf4LYco0S2L6vm6dsHIolO+zs2Lcl8kYT5O
H2wNUbAj2M2d80KrLMr3IGoZlLweY4LengPkH1G8reNxWGghw+g5aNdjttBT4fGt8/+b2BvZmTs8
JVBtRyY6nTf0agPCZ2GbOnqCTIFfLQUg9NMw9pq0lnQGWQCL2TrvLuW+yyHvWTPkMpVKnSDpG2uV
tX+xVic/CLpY7fW7Ndp3crRBlWyBNzJakVU99wwFWrkC5ht6YnONP2dC7wawWxMcEq2F3u4gVmKz
fE2Kt4eIvdxbVuZR+gEAitJwBcNnMqURuK/cxoDS561H+yeCFS36y5F0ezbx9pATP+9BL8/twOUu
99QjuIDZbuLDqFkLA5NuBZxEXkmFiM8wKGyU8hHNfv1UhAl/6i5f0GPXzjOYbQWRu4BjQZOiglwQ
TTCmyVKwVCq8usRWWOV7Q6v00W8b2dStJNVVdf4l6Tk5kOuVvAPM4tPZbXaqEvkqU3VyqoWaHxUv
6iRKvCIK3iqutWNNm0NhZBJIMhyxsrjCioYpcuUQNSE+suWE0vF+b0tIJfA4PlaRdp8bJGGIqUnc
WJBR0E1KPxljhGBX9nISotJFl7Lf+fPMnwKS6G8wsFvdZqFC/nJW8nNetLYObk581gkJG2zNt9Za
OnLr/2HVcFFzKd3CBEAb/QSaZu1owS45PoPDtADxXjCc2oEG0LqST7uvsu+qJxo9bhZTyY9Qy3lw
hopTX6k5DZi0r4AJzWRbOvJegCce0KuMpmg4lrgHUfjCyoP3AfhYfd4FoR92fOs9uIeWgdWzAtug
NMvjHrjkaNi7caGFuo64oOLo99eHDAvmrVVuTiwWM+dztM5rWwY2EqAaZiqCs3g5ElyOmpa/lldt
dYBN1dUfE2A3CBJY9zDzfgO/ok1NlAVRbTXj+EHAcx74A8BEi7s73IvMFXB6HzfnO1OAW1CUdlKv
abozX63nS8qaYounB5P7fzYS/PTLnsy0ySwlG7Uk7MDyOBbJXYpnnkyWDXL0gfPS+OJw128BLv0P
6XbCCnXiTJrtQYmAiHX55xOR7icMA+SA2ZAnS6UEOq1qmLLd3CwtDr/mpyPCOxl7MzR59eOla6hL
X6stxwLwKIieghM/vOJlZD69V7bRTuDB/Hc9ppcwuZghtztx1JAG+NG84LEHxNnBWcx0G3YCLv8c
CPHi3WWRlly+TKqdeNdLLmG1A0zniDkCyX1KHl1llm9fg8u6EBWNjGItYxAEHS+4NiAXemQFH5NN
sr/gxKWiRhRBUK6LCbROu8kiariUj/WDNxaN/BZsOqE0SpNj+SWMD2i6EDbqpijwCieshXfacX8X
kWRSxV2tXfVoKAL+pz4bMYQTRD0X+OPTXhqxKydBzrV6BVthO865LsSlTlfdsIPlWZh/E+nQQpwe
0wJT9o11yHbzkcN8zHnDNMHL6a4zRniiKX46ks4rTTMrtWw00YIfNfG/O55vEymVGAOeESjGksIq
ZIt8eLavl+i1T5XZPLqYgIE+LSmK9CBluDBAPvXpYSbfb9iiOWrG4nmL91ux1GV+uPCb8jWSch/k
J74mZkILJXVg9Qk16kZf0tOfYH83oDHrZ41cKyXYGOTD6miBMMOqszMJIquf5/bgb/D94vDzyk28
UY0Bz190nS5C4WxdcyHV/+tI2I/G6J5HXOwCP/m/xIVsnrIn51d6rEJIngjRZV0mBQpHVSTnQzy0
BkgoR5DLg+2KMS3fg889TC7Np5wbScbdQvZbi/e9sZThaj7zPDf0ZLetnYFvyqd3MRRbdsoZ28cp
XL0VLN8ljHEtyC6qM7Ddb6F3+ibsU/bbkzNdY8WiDFQ7lkyjZg2lTq0645eagcKwSDfjap9X9rdq
ZRA4rjroFdCwoCkjgD42WSnjQKS4Q99OwkxF2sBm9hGeRcnMxK1UeoOXkTkdoB6Zw0xSY4f3tvfO
WWXagie9jV1LDTKrEnwKEtAfMWBYFdTSj5ia0Cf1XVyZHGuuEsPdNOjY4phjHYBNv1PM5q0TOlol
q34b4bxIYgGqUktGmYckBBywPZIkqsChIOnKNoxMDsz+qWUrOI9Fyu65tsLnVRJjX7Hb6tO97w4Y
i9cVBQRtZvNbGZ/WMvVdsOmScdg36+Qb82d3UXRCxm5nDS729bTO3nf3EFP0nodsdCXMB0CtnfcN
9ujtCNVmAY3LdvXVbvj+qnICztTt1J0BeDC4SFtfzSY0hUwAwJ1DoaOyUSSZIvSINArvVKL+e/yP
3OD90BIfs38amZjbdwHvPVRPg1bPv5CYgxa7e0Qq4y1dPhmHQOiyNIexIntMDbS+ElYqn6fObdcd
7xnXgIW3uoU9HSoRL6mYtGLY801lzWicgaSOz6LZRtiOWtfpU23l1gCWBo5Oc7sctTdzLBftc1Go
7TMgweGMuXPLu7m+KVPGcYZx2mpElxVvnqN/Va8X4ehhmDRbG0jvrYeQ29SvWP2jn/itQw/CwMZV
p+96cN+WmHgEHvjI7Oz61IKdpSsGuF2DbqmFMGLSxYs6rjcwU0+F28VdqZRWfp9+fqL8jaWl4xeF
+7fhBbuAwvqeZIP88/qv8TjtEqSgQTVvhiKrdxREndhca4L/VV2OFWLWkShQHUQQjIt9GmRxNf29
s9R269U5jsjCNq1avncG6Koj31PjRfUWDSoE51pHLlOS63Iqn3bVTjUgSPAcg8HyvPM4Kwo6uj2X
pzRRheMPM+6/dPPr5D0VBJsVMDVYEysXEDicHDeqi9zSEYgVyd2AiRo/gG+IWY5ddVkhcfexwkdU
+KwRSCQv97NtEG8JVRKbZVcnAFJp9HxHlIqChNyjFXzzP5xdV2TdjLhUTZiUfqyBhlP18qQKcoeI
KOkNKV2whsT/W3eqed7NP4Fn0GKNriYYZd0TvzqaappuP7pOO+WXlUtEjCLf3q68ZfjSafGRtZxJ
P9qwJqm5peSbAeEf33h0aHvWGb3FS5n7kKd2GBuS5Rzx87owmOY6D9/5d96ORdM+qq1EiNZsslMA
xW/GvvdO4tpTXtc74lWC1ox0NO4fgWENvlmXbyeSygNqrgm6EQZq9zr34p7bmsBUxElZatpehkAo
8tlix2D/H2AQ9SxxMEyA3OBNdJLns7GESwQ0qaHADWuuKajQYyI+5GVQ4ll5pz6x55uy6ZsWW0lt
Lvr5p60/eIlMagw3p/b2ke/xGmZ0r5DZabDASG8OMu4bzJohpihkT9mnUQpNJo949e+DoEiMXWK8
+qQQzgI5RrSWisuSbrHO3HXTs0e+XlE/LF0OfA1AByv1IXcY+vpXZIwc5b1026msimsigK0m8pQH
NTmYl5cVs1jcemfFIPDagTaxd8e7VGbXpFqp+xVv7DZ5YVR9tyk6nxaGcYjOePnI9trcwO4Qte13
v7ChZsd5jlHvURQi6Aspl+KXZTSC9XSHTy25SngZp4W72eK2yZqqHpU/O/oAymXBXtVDfg3muFno
G9WZxmQsP2fe0Mi2luZsxh55HHFawGhbRxlZcY6Aa/xsu92K1shRmnPT3IGT0SJk5c33CSQPkq++
l7MN/72xeHwSEm7j7IDJMGsHrPcLwECMljwv3F8itWwh+1fpXzKZl0TJQjznnUiGUt/XQWoCUkjf
n/eM/ifDEKZtdHjaQwOM4/pR6aLXdfwezHMp4E2dGxMQQZAY9SHtPtehKoIXkCg/P/6PTjWqtIB3
4VAv7GvFQbxFo7NRlijEA2LRnIRVIOSVSInOw0nnODQGZDWWnZmzUN1zcc1AQ/q2MzDdLjqGwlEQ
DvKErp3KRkCI8SsdNIwVme0HX4LLMvkxn+9kNFQHSJHNYJlx3pjEgtWfZiFEB5mdPRuql3RVlDZ/
JqKIfkgjih/wjneG9c+nu401OtPc6GXWLXV/JENsMW8zTU/PtkqMiBpiMxNKB/KM2neG1x/iCLFI
VEsNQ3GntenNPiSH6KCVXIIdBfDwmwes7mvNNH0+nP2/GmZ5XZQKulHLUUFtIbAiKNbG8cM0zYCH
IcssZgWHVgNxSfRgZRV6n8Fauv9hmA06+33P1pJYRyqbhhjDVGifVaLk6809Mi0T09Og/bB+FqkV
eCtZOe0dUgL2kpU3Cs7OBV0OOSqLcmN8S61KzWorceT3wPRkkUW4nHAlzT4N+ZnLOG+Favtfae7S
3OWy3mvje+ffwxDxeyQUGIWJwu6OtH8ve4U76vg41w4wS3+/bra2CZjZ3JVAln3Vp8tbYeH3M6MC
fW8lxQBdewiPQP1dxYDHQuhsq1IcxhLPySiN4xOpFKhw2FiAfWCM82LL4LT7DIt8bNGtgcWQ4KTr
10zjrdD/tkYGgI20R0C+dXJiQmI7MQ7zaTv1VCYPL8XM73S6U1SblF2knnAltn1lWeiusRMgHoDF
EiCbl+r7TKEihvF6Ep8/AFnk7pL6wtIq+c3ma4TexIUsr20hM4gNsfWimTI9hqKXg6yexNH2VgAH
UB/Qac1bhd1vMkLJGnvkTajkbBIC03PFu5ELfmbbIHzAWXTQZnw/iW961nSQ9oTCSb0Jq31NyHEp
Bwme3eGIknDZ0SwKYL4OtlOJAbZ5V5rO2FQFVEloUUKVky/xGuOG9K9yMDLbdvP3VoAFsW7QOiIG
B4qAK4KjrJVklbWtyugm5hvsgySYPXyU8iv7215AyQ5EUx2dgVWFGQ9zU1jX/6qgtgbb4yz201HL
Ro5Z3CEina/q2+Ojb43Jz0n5nioaz1ppg5QTak0oSXO0bDcdjJm3HHfg324JS0DfNCpR+vL57sN6
ABEaZxmL/SyIKFsf/Yb3Uu6SN339IjcFSD3bo00b74SpXoxWhnq9aNsJOo1HkIjEkoQHu4D5fP3w
5ItuvNECJ9v7TCIonZ8hVpWz39Wqz2br4sF4OLqYtWYW/ulF6aKB7PzZ/hzmYdfACgVT6l/UtCwL
5xH+LggBWV1FBURd65Okol8mf60vhuI7Qh57W/byEClcoBf0yFm8FOFEBWxvOD7CcZP0waALynpC
69midY/HiFk/gJcnjZj4vP9mu2PHKlShbk/b+e5Kwfw5k2mYZzAsFveZZ2jz3EXw7yWjGgYprdD1
PabrPj09KeMYPw+gn6hAgdpf0/hpbQlX8XbXz1vvXNxTxOmtvqcdDi1FKgdQ1a+xk23Hu4mhgoCS
nYO0L7jg8EqEVtxVaffE5xwIpT/nUKpzUY+0yfauDbEI6HsiJ+dBgoPEpzya9S3aHWXNS/PlAZE2
BAI1TW0Bm31D68knG/Z6d4M8r2AU13AowSZaZzfBpxWyoRzio/UTIq7NUyjV9CSZ+fPrIPR3NWSv
RvL9CEGBnhSKTZFlw6+qnpnF67sinzXuaPbWuPm2SbuzrDgkKejhOFjEq4f3AAxPCvllznpiflc8
t3A2tDA+yXXQmkQIlhOs6xUlhxIbLJy7b+Jgy5J99GJS/Ph98pk4RdvwFR3bgLauajzj6yn2iP62
aldDW+8QjyqoCejosnWKoUOFvRq0fxDU/JgC+kQU4fv078QJ8156xZX3VAc/lDDAqEwJ2kQEkvl/
MQRKC9002VVUNEnhjoBBAWDHKbaBXjxHfBJI9vewElfO3SbW7r2Luzv1Qxxh4lqf1gGRKWp59R7H
YC7/K5wCQObnmssQ4xiazfOu7wJp6+wgNq16i11DbWoYy1hJrKRoibci4fBUg4RlujSnECaXlj0X
xlbflFxXt0Unno+J84RZHaxRHlhU3X+12O4PHUhQjS5PWhQKqD6jXjs7Xov3mF4Un5WftyKYBvfW
aGYg0zuUCTPyJQAuV9AXrelczT0sq+yVgzjYRGvvHpMz/gJVF8FUdIK3AksZC7I8farTi6NhTQiD
JwrKneJuUR+/ManAzT+IHUeDmBLNfRhprlY7FUeFO/B2ltuqFbmxEyWx9TkEq02JVB/RMrr5zisw
TeDtCmvNrVv3+4y+g9JZ3AUP8BuJvScyK0MN9tHfPO29Yoc+Nt+oOllDp4GvooGor7clsLE4F9IU
k64h1W+dxiukBKgVm38Zntg4BgPOEte7QsjA5+ky4NMLy9Pfm9zJaHwI4SYpjNILwjPMrd9wrKDF
lmBYzbXh0Vc0G/tDah7X9r/9UKMSSKPfNGv5cA0BFrqco5GFas0IMsGYhn10fHKCeL1Gqa5ICULF
nvVOJzEVjRFmHSRI1A4zqYd5hK26PksYyIUKAVh/hHlhM7ftloj186bRmRABMTsqLEf/TS7C8HjI
zregChFwHDNgP/AGnQkLC/4Zhze7U8Pyxx6oA9h0NvIIEKUdqSN9CfVt45Lp8pr+6d4UveE/0RgG
itvBA1M35yA0/Irlm2YiPDbdGiUhskUAACaJMTy4O6O35xxheMzFnePa+sMY64G7Oc7ig1BkrigQ
bQGjdmztnXUtTmrmgfdgqRLdXrT7HIIjYa/Hx/6FvlfBo74NfKU0NeZt6+aBt4DHjRsWx+hVrj3Q
gXv6ZTBuNJcVd7omvtHYT+XrYti8dkd5Hq3FXNpVnj9ZwwTPJ5egRP1Ddj43x4yPPWULRn8HpEY8
fapIrWVrZF8YBP40nMnWgVFW4bxeDxSRLRXzUbX+NAg6IbeTZc6yGV0RY5YNlKT1ZSDTZytDCUgS
rPMcxn0hVRupuUPOp/Ur3pIjTJDamKsTPC6qePr+lSvh/NLKLlZE7+/xt1nJCKJKO0wlTxAq5cRC
5Z+8jBy6XtnBWE2mTB2IjrQ5lGrU4T+VsP2GdSO6Ei9JAx19GJVL+97S7JwLhEU15iUiclHwHv9S
ZqZw1MZKoJ5UHJ1IhKPL69ChWNApik8t+5Wy/LcNeGWTvQj7TXq2h8guosQ7M0c7NuDnyDWzu/2e
Z/XE6d8SR8Z1CZBKGD7MgiwqGVyQz91qfpWLE3kZVZbrUdy+F4nIJLacux12DlOS9NjIFI0tKcpi
r1qkZWVWtU8aVRjj2y3DyAkaEL09BEn8vpdnqUKAQZbJJklUuZLg+yCg5Pl/iZqnFxLw91nLuRc/
5LZy8RJBBUcAqO2UI7ETFoug5OhlbNBf5Z7ZpQpuV14ryPOhsrsd62mERCZaYm6h7YZeBrBbc8Zi
lcUf76KFUJuDoWHpfP8lj5QYK9Xln6UHywhjQFxKRdZQNvUD4jeZmgBrQ4cruEIYpQh8TbSnsZYr
qUHj//oEczfZdsW/lcTeGy/B72gY2HNQZP2uzM93hiwRPS5LAtuGachZ4c6sBXu7eibtsJbCq3qU
3Z/Ny2zPukbuvePDWQRopYJAltaa2vZrAqthaC3YTcJA5eV8UAzHtCjcvNjh0yHIecMqyPqqUULb
M4ZDZN/7EKuYVOQoxxeAuoTnaaUddUO/US5OBzsV3xymtiFuz+wJmDmag9fOsD0Vx+T5U8ztUG9j
soYRRcV6Q6MCu23laam0bETvorQATk9YSNQn0s2TCQ0ybLx3iz6RaR9Cr1pLsV0kGW1PrSDHFCxX
aXPbx7wvmhb92KV5J6mdoS8ZfJ9gkh5zvk1IRQR4OZbVIhk6yOsjsYRjFosuWB2GMgGTr0pNsxg0
5AQnvOJKUOUHu/OOkEJeDVjjLpFd0Do1Qm1IfWICkyATWCOacVWn3yEiMPm4/TH5gFUoUloOhU/x
QfBf7S5J5lMKDCJBe/4vgh0urmnNZnA4/sfI9Nm1qcRCCg11/eKFUhVNpY8l3BdALYoupmLKBi0V
0MX7F3poAmvW0qSidoIiHv+lxuN1Tg8WofhzzjLBRWqMhkIwZP0FntkzIfRxGTWcbL1CCCspxEMB
JPl9CF1SKGwQZmgGr6EgHPVWWLSHWlYwb5c9k/vvWCg2AKwl+ndGNhrcg6CNuJUZquLEL5rE9wts
X3GO+wh/BZDOoIn13ZE8F2+9vOTzz2oKfDNkvn8VoSB6N4C0GqRKVmG67QmEBV0HLATvCEhia/gR
N3A9FmxY3CKy23cxrgF9WTywGlTbsBvOevTejimJrw7zLdwRTcKCGnszaxrrljJQF/LdOtiYW6AK
yuNlgRTuxHCj/uy79qzDnFJtdvHFmW4v4KuJXnfXPAuFLkuUn54yJeSeSgkcP7johuuo17xoCjfO
0ZWLqh2o9KvAqrpI/SRNiWxjtT1TLzxu4jntgeTt8H4hCKayAhlMGrfZLgIgtHkUmNZywrKRfRQj
+6iQdlx2h6S0Ti65HhPIaHlX9k5EYyTQwpJpfWoZlRA0plN8/FhUGc/PDSIvheqppESnn/o3YefB
P4O+DEwI1r4Hf0XxroGMhlHPuBdMpyeMp6wGLHR+PMUWNMNN3zsxQ+CNOsxhvq1EuwTJtKb0T+9I
NWU1j/kRLaQBDmdX7RAPjIXd1qx5Qf9qgqhLJPeTK9JtKxpxDWsTXAzTYr6eWRMUFV1sIxS8IMKf
c71YeRKuaowEfkwD3+QTXjp16FhE0fDW8tn+rD4JWXvGg5kD46MPNvOcDwfTFvmX5yc1+cnc8Rpb
XQnYud4WV4P4ik0INoU0IRd80zMto//Dnm7k9tGZJn8huCKL1t8Fqm4G5k4O7TIVk62EX85fAgoE
zvVTg9Mg2K9TczdI9jXMX6wmA9r5wXDV1eqV8ZU71sbWL6vivQFbVr4sv+EiVXHtIc1Buy4KWjrV
MkIGrjKeQ1dNIWpiFI9BF1g9Jl/uNsWQZZABWRe09a7oKxTpz4gOy6MRgXeNi8NgWIzTYKpyEm3b
eC88sMD7AfsihovCnPDI24MI9izIkXkQggDk46xeVrYFOheheVRkGO+eblc76lxUoLNZT4LFmmKq
MAuOS2H5LgeMtpVxyM8RhrvNvnrLt/JIkcHpT+4mbMCgIuRFeTZVOslzWTp8zh17OGeLiUyKGEc9
CARj9lsYLa6tW4CGxoENy7r3C23OWGUyKfOGd527ILUiJYJUHbHHfSCwH6y2jd2wFN7rh1RaITtI
vRTFG+IAT/Bu16Jg93nYa7c+mDWmzydrPI3nVnBwrPSpZF1x+vzKU0mEuFc+b6GNC9CfnpEgTnZW
cELTRxLiz7y3eHhQFrusJxFsQPChKyYk9aO0UZWr3haCzxPDR8tQyAeY9jqb6WWaU/jkPDuqrAwA
4qxOu2c1+tK5IaIAzTTdblCePGrjQkmeWyF3zeMrIFSeqALRAoTt1P152Xxp2guudaxz9ut0RVbt
YKQbCsuiBzz7xaj8h7Wke6Qo6/kyzJ6wjXewVqzghGlvMsj9nAfL8FxsmT1Wo94wJlENYmNN2Izr
+qVtLmWfcApZhd4IZBN8Gdt1EYp5Bh8eC552g4aw0kEV2cvqtPXAyrih0OqHpRAyEP0ScqSKWPAW
loswsjygj3X9p5KxYP3hsUQ426SZBnrCErIwJlMRfO04We8YG/UsLswtivDhPFUshqQfI39Q8Fxc
x80dL3DwJLhNrxv3yfqM2nrJVwU5SmA8afOnGT/qGgYPgf3o87x5kOFszqcwMLB/zJCHA/6InkLp
TiN8o2IdNZ/QKDuwAX/Ix2ngHycfn5i6MiTdHWPv8WgKZLB2rCDHuPpyt36oA0hTRyGh1KZVyBSx
bve0f6DvaDRFWPysqItfHGc99zLMcNJDbOzmICHFqIQ97TBWMl1YRUG30rwcUrrN/+I1ai9N1rYB
iGIbGn27LNcT9q9ZuFnoDfkq+hjuOq+gMnrtcUxlS83LS/rNMGFCGW6y6UQF/eCDAgyrRI1JUyXG
D+Z9wZvz6jxIe3Lxv54/jwX5gAp0+ap6E2fAMPW3T9SgPdAmb8oz+Ft/0n7t/ywIoZS5I4wneMY+
kFGdzbiBkLpJQemH4F6gyfqbyFuou44d3VzWl6ub1cHz7BLCzYG2cP4hdsjViJNasqZU8p+sKp/8
1rAoqhaoS9uDGZTRtUETY4Rqmbfp9qd7f2Swfd8zd6PSGh7NjOqMPiYKjRKkMvfMyV4l1H9M7ncA
M444oaK3O+LvUmHAZUn825TTn4T1Y27QBm1IZofhwyimG1olbybF+UuahkoEPj7IUdUltYIqi4L6
f+164d6zImKAGMV9Om9mrmQELKsepLzFGTnxzcdxs7dy2u5q63PvOtcM7MsoB4jHvie/34O3k5FS
7tqF1ENxQo8imekFNfxMK885+Nh/1iGP/nomIS0mgZEAgervBPSYPDoxOBrWHzDqAcdCeyo7WFi7
go8vpMJs+JpYKn14ypevsAqO00TPX0WOXvNObDQN0p6Hty0EJLbDIxwtlhJLbsp9gZ5shibLQu/M
stbSmOrvYNPuph5kmr+l9sDdGuzAjNXHVfyiUWev62cA50xi02Kmkr0aek6eXhSbhWH6WUo4w5AB
fkWmaEduLVo9avU4A7MCjufRQOp2pBAfOmqtVzkHG5orhB1QubjnqUMFJNF+ujit5zzJVxgjC4F6
LDNkRD3TREkq9BI6QlL0sXBLJ9Pe9DzSbO0AEKEt9J7j9tSJMhvVXjsAAWApX7/Paq2WzdXo7+b/
kwAFb324V4WvaL/jIwhe4r+AGI0CBNKXQGEZdUxzaCEUfLFdEgt+IudAeOfgNv2KRl0ZGjb1zj10
KVeaIOfD+eMc1iCJA4hbeDa8YFOBusSdqrLS+Fdis0GSp8kwXpcIBgi9XcMPunW58M8sOXEVobn5
LpdEtOMI4nf9bJb0Gau4xIXr+vi4mlYFRcH40PwuAQYIdYH7HG+TqJCtcdSyecVI5QCHxdGBXZft
+lEFdZ6vVziBBTgbxIm8ao2okQsHl4NRCavjUu1T7rBmFl4L3+2zQYE0SaZ7Qn/qbaSVutcqn0v1
+Mw4gF1Owc3C+LSY7LLYp2hUY2PrL2A8lk9Y974mV3TcCrpUzXm8xULnBOllVajSZGghbOv5sQ9e
3d5Zn4SyoujgEQKjyaALpnhl0Y4ITHcqvu51PnZfZ+iLgBwsjeiPACpW51l92ZINSTalnZsVpLq8
8pNtqeUarXBoRUxzPLL6STihceIX+gqlvOQIz9mi28r4mrhdmU045MX8g4+VKfjTfheiy6W2UMw7
bKA96hEcARiS44fq1jCMgqHBAo3yW/xNilU9R3CODAvUGW+iSC5w2q2K8m0MfgQKX3HTiSo+57Ac
CKCtDrfiMbAt4YwyIUwPlwwP2Yd/LNkt7Fr/l9lpp9UF7AEZjCWPUXNqfj2bd4t7a83JcSAEXAXR
BAGb+/yjrCNOH2kEXilYTo3ahq3EJAjgCP+IFdRNfuDjfS+9e6gaIJkg+KfzloQZTqHakgu1ULp2
H2/DNaniBN8uCM/a1KVzSYRlVFui2NnMrS2VAftViqkmK/e9w1IA3QcCeM/WlRwtXBzLxFfgxmmQ
lBpRtkIsovPz+pO0arjRUa4Wy5WBdPwYcOzIFcCcj8uIYBYWZePGQ5RH2kNVgF6+2DMcZKOzgepr
/hpUzqPdGOtK5rrZnSQCKhdBqSy9Nt6h6FWQgy6NqbUHeBTr2mJB8qLo19S5xFiW6bB+CsESI8Sw
u3EF3bQdrsTgJNqGtCS+Rlop4RL+6EBCdnvtbFlLFLJh5U+xQt2oWkG6ahRjgbeiyO3G1zi6Ot6q
oBYXcMerJ2YXuKMQRdlsIYkHvqX0ZYUiHPEnEw8ZJ4AK4p2EQB+Kl3GzIhM+/Trl1yYiScI/Z030
K64u8ViQeayfbLX8+WS3nppmJs/Q3Mw1hg97ynlc3cb8qq6OQEcztAv8MneAjQ3zaUNIm6DzymT+
0HMQSjFnmoeFXOLP0Im5/C3YPNET6TNtiZCgOOPmw3Qf6npDdM7Vx50XebHAoIfs/4NlqD5mzlJy
q+itbm97P12cRino6l8F8TJw6DI/zjxogfEs/qtElUznJ2R2V4jxYE3I24dhoBQbYgjRL0098+bU
p0tEpsSKWh9cIg1d3kvEs06L01EPZeEwYta696uZZWTMWtWvDHJynXO+cd9QzIyHU773R+6aiYBB
+2wHOUySVoBjt6c4oh+/7h/BlJG3xonBsGDGZZdFmKpR6FdENGWEUcixVPVsuqiNUOvJiODOVaJx
B2GUtgvK89eRnTOOf69Ex/iIBAwkB6vqie/FstuQWLKrgDOJ91e+NnSCgz66GOQXDzB117UB7O/I
I+8H0fyGCDgV3Nky/NGiehvSQPI3VM/C0963vekmikkFjsc0YUP0QDSdEgOyo4LtaKiGLjjPXJVE
UXXEodc/yRrrWcJ5CiOPZqDNFhjAro3wWNQlL63TcDSFhS1T9b4Zg8Gsuxh2o5wZg8ILvF/MkSgD
9ePslnZPT8g8LATC1l7OOZxP56DapHyv502IqFewsSp6w7KWaAdQBaFKO0aT0Rqqgt6TXCUaGZuQ
sfWfzzkB2Ks5Yoh72JkkL2q02LKsNk4VVJ64SZkq9UryGq8PjSdiMI2+kZ1zBApDCWMRIIeP8Hdf
OQ9NSoi5GlVY4tHPGPxVwOm4/ykcs0qcnhN1BRerHYYYmKXQSHjHKqZxtfL/NSaDgU0yh3zoBa3y
omVQutzX+GLlD83DX55RdBO8obznxdI+afAOz2yzkz0g80ayZUanFdzEWpyKB2+LN0j44AdpPUxJ
2zieB+Pra+lWim8yA4bPg/5TMLwD+Db2vn0Vmqgj1bgE6/q0LwVw8m6gM8pUez0mBRUSfQTfWApN
xFKAVGnMa5vH/0eEcmQYLzhGi8audeizYvHdKBJ0UbVnxtJlanTE5q9HFpsFvTpvtY3mIRLzf/ND
esV6XO2wrXZ1PWEa4JIY1y84BI/OPnQPQMR9Y3FBTnaEDKJx2eL324FLkgDfKrYR84315J7WjLny
/AU1l1YtX3HVpqgP0Gf3BkW0MAqZABmzpbUtJOOE4NdGXpmrB6r1hdraLLvfU5KhGQnd7ja4iqdn
xNNzlzSHjMi5sgiq0hftSIMh2Mu+xUQDrb0eu1w1VLG27CPygRC+fTkNlRbSVK6iKC8tCDmwLQ6T
YV6zsiFiRmzZxvuhhYFm3u54DlCw4MFLjpalDEU9h/cRGwZY7Wnrd2K3BvxpXNdE4bJMPvnUDqBX
xqxfmHQu4KT23vGASrFBliW+TR+JQX46OHkkz2O8yAATHac2YNw3Io3lZaUZdxFwDiDVtOjUdNlz
hx4yI85X2GFPGzQMd0DQwWObHGg8RsZ3mdDTQEGa75psrjux74xFr7KnfRZ65BfdrlvNnEvRA2n2
WpjMDW7GjkUMYLsARsV+rsJyXEifyk3CO7BFNPd3wLm416JBDn+18EfMdrwIVV8qk674+4Qgx+aF
M+XeIRQEi03DFhJU5ILBaW1QLwnAXA3tdAdFWq0N6NSFASw9lDHE+FsF/A9FzQXeexKEy/wgCXEj
UmtjmzYCX6VaKZLgO+rBe9MlIfUvAZ/IxfQtIJ17LP1cexooeRkbY+fhrRIDPj9es+Li6s9DIZdj
Yp58DE7iNxbFcSNMIE7nfMbHxWhwuSOxNns3kMs8dTi/SsFHuhAVkqHZNZpz6ngRLllgNV8l1pvo
KzijKe451mJTSfsH7xAJJOXpVCRAlaGOzEhFET1+7y6Vp8X0ISTsElcdFzpWTRIV4dMqg6w9wMTg
TLTfpKUchCAvzTYzqU6OJSnmVjWLeWZ8yU9ncO647Z8DROwyitzMQ16QL3n+bTMHR/3G05HajU54
vpn1PQq/sPGDMuIpP6WkLkgfIAKeSXkZjYjp4ee+KmoxKYXZiguUeNW7ggn4GEHXymPDIwwrxKph
O7Yzahn66a+dNwpzwsVVU2M1NYdNYSISweU0eQd/JYg4PWtd7/DNmaHSdGhIDGrVTpc/Apblm5Xp
YXmSMeSMDhFo3eAtvoyNfzcGHlhGIu+Bsei48cKTrJ7fgEQsOEo7ga6fn0PLNmpkfBTfus2847GK
+j+sMTdXYPtgpPxTyWzp7VFEIDTrdzcQRVdjtUEfercjpZpOYMloZ7Is6EKWpVGLDtVV9m/Z1Rwn
qJlENSEMo0cX7jzoVvGpqkqT1qKHMSHdrgYTQjr2w7s5BBH7hrBg4f7ADBqJP2XTaAWK8bfoEBto
sS0t5ltX5JV5pn8d1OBGy4ecNrYFdTb1K8IKaiA/76i7EgSZUt3N+1vXixtcReV7Wv4LOlTug9P4
ZkyzC3uNJoTymbr1T3zXi+a+MMvxc2ZicQSR6QnM0/h0TZp5w8hTuHG8gf5horSPOWyTqH4nVZ+A
nOk3XJnMr3WHfqI8t5ODncs8gUqevMvTCHgPMS7AVc+HzfeSGzKboWP7UBsBdSb0547q7d+7aYQa
I41/EwvgKzqjU1G6TKJVlr85lMC+3T+lIy4MRxz8WYCTEaO9+D6m0ahrTxtpTTN1EHPobbTaBY1G
gXdywdZB8ie6UoG9iDVmLZBAzTyJxN+HUSm/0sLYMM5bvtPBGdtH+wr85i/cz2BLVFAik6SnFlGI
fI1qzXrOCP9DE9TSLqCjOJeC/MTU6EXnk0Xy+A0QlYYKH6ZithTHTAKVn3uJX1gcXrmuklAUD27S
8vk/PnUneWy0TfatklI0tTV86qbkRG2BMjB+TFSklTJPezXA/AfCGaUQlOY2ofFMNriGGbCmyV+7
uobqz9IeCASss92OvuTB5sSNUjvTth2GTdKDI25BxDwIVncjuELg1T8S397/wGgTWqAKts3/JMRf
xyEBCs3mKtCvkQr0b5+DcgsIM6A2OFSXMfl5GU4ePDzZr4+ytfzjk5/EkPACy4fQMjpDyWdQ07BH
7beU7UKlESQLEwLc/aQAeo+FpqpFwwsomBgx5qBWaeeyGE/c2OB/sZYK1CcnnoykupQl3d9CZAnU
IIhD2eyns7aphlAbG23dvA/KmHfQ/LEy0uOEb4QC5WvfUgbL6V0z2KXEu1Zl22TJBh6BsGfH2/Ck
nJSRBiYsnn4hXwGBV2KvgkvEL6m0Pp4NZ76Inc9pKKqSstJFJNFqTarB9rtiZS0fgGeGDuvZlYxv
wfn31Sdj2q2+bUCIx8jdWPnVEhUVD3Cd398hf4Gn0IPHUgK0Ztpy1nPs4sAh6BLgfYi4ctMcgL6s
c56uTGOghhhsza9LcqM7qaJjYfHDDTv//cFIjAvM4jclGi1rpxJp5jpspLmAubUZzKlVCsSLcSUB
ceaqJ6OrwYmBGyCUMUMKYQm0zAHUbVmws44gu/LY8lv2BmEjllWWyDK9k+FS0xJHjRcoFBZXPyOh
drT5k8X0mmwhkqxP143FjWDmzCZHKgm50eGNYm5EPJmDoFMr1dbUFSsI6jwiJqy2jn2f4ITN6tYx
XBy3ffD83cOVNgq6vIrmtQWEluGjWBHXcXa0Vef/bx1gQ9aiRezY0a02WJb8lTGbuDyZdAWUDoNR
LpiFkAOGhHVwRpPktxS8vlIOecyF2TKDvW6gfxPL7qAbwM89KZSqYpL14dlrP/rh4s8Kpq2/r2pp
giN4Cxnboz8z3ZfGQxUF3zdbL0nyrggZIq93S92jo6ynUEkEHbAPLcMoibHqmY+6h/Hne4/TWv5X
gC4cJvTuvH/k8s6bFQs4dnv4xppQhFcEg3jUn7cUbtyXoIA+eacYT3p5/U+vkFKbio3XdE1rXJf0
HOenRTmBQk6V+H3yV4U5G8HIJ8fUyuqDkeFWnl+Hfi0iSrUMmbCX+VANWu1gjpamKZFWqNjVvjxF
0sNytDgHR+M7PbToInGwuXBM99AET4WKhmQfNrpjtwewJOm5jIb9DuX5n0C5eul89+tYp5M3ticZ
0nqx6uE1UgCe5Macpb2P4A8Dm/VQcJp9ihC9DOpqO8IT9ZLxVFaFyFRgk146VjQr6k8gA7q0fyh9
fOxt9AElu9Co8W0Qrdpavi+yrFwRJbn+HUOGY6cUMtIzBm71bKcefmMPh+SY1EBMJamiByEGaZe3
onXgw48rB2EUfX3rGX/bac5B+0EI7lip+BnGHSFF2yRp0QFwTOpM59qW68xM2LhnzzPG/2MOhnP8
sYAG6wz6A5SykEPinOaOjh9U3fEeqd65zK6Eh0rSUorwSNxk0ZFlgfF63li9/V5aRHrr/srq1cdE
8XUDb2Qpre+AkIEJuK7vca4AZOFz4lHglZb7wu6l1PT34WuM4esIBnBl7kE1el6dHGYTyI4Vuea0
i52CH4lFiKzLrf/5p956NrbnJSbP5BTkoCJN37bg0EwQsiR1oEE+jDunx2ck/3HuiIlnRkJF+YAs
su8UxJbYE5boE7LwNX9Lb0L1i4i3uEVe3KzeOaO1jkEsbOs8B1YWt7aFSKaxoJGn+dktLdG5hu+f
oWB/93SU0eUhxTtkFcYYa54MsawXazyrJOpT7WouvLzEyfFkHnkishaqQiRgMduy9sHVk7n2oSh+
yis20XrZU1z6Z8jYmwRRCyIZoA6Y0ShviTfiA8Xb3knmjU/qy18WIsHg3Iz8En3TNnOH8Ook+vBy
u2+gy7v2+txGpDKDnUPAc1dxF5RVusg8ouCaetr99lu8SIozYgS2pw0X0nCwl2/LS0AH2aLYl1wK
BrycUMFuqevyzjzfi8wZQk2KcBP59n/lkUoipd7yx5pF4RfuS+ptk+OJSjRBwCBXR3cd9jpHGFZ7
RGoQGxqy+3SwElzsu5Q6QocyFE798Pd/uxQmQvpAq9Esp5ccJC5oUbFzFnx2YTSuM67jsnyBi3rJ
gES9TO0FinPpa4vmfZmkCYBVJSxKTsnqmUIr/aZ50vG7KukkUQ/YU8Wrnz2gD/xVvLNBxUCS/a7V
DWjmaAqrKWGaYGRbhP0HKNFSFGono+hErV8b36pQNflsfy3cgTLx6DdS6e4lU4j+Rllhh3R9+2wz
bLSTGig6dgrN4I74MyQUrl1rH8S90MQTD7OTzO1hyeVjfqcYnjMPKDPhNg6g7VRCYukITk7yP4Tq
p5RoSCHkoJ5XurygkQVXN2KWcmjbNra4fV8b8kr8Uwc7Aa382HxQ1/dvWeuqj5pUCitTwwqwiETP
6cCfHeQDmrvFvwYw1P4WaGRv9gw24Oe9G3mKrVTDAQRIxEm2xhOHfDcpkAYOcvUCueLo04+XeeY0
9Jynjqh2ioE+dT3ITjULofcQ+UvvNX9J5x4ADXbopzbX96V+hqhCIKxMCq0JTSpdGpproK//oWUe
lDK5xdDa142fXRnvBDLkkGVsdzs4EsJqxQocPXj1e1mmnfVyuBPXh3Mp63Pq1UrA8m9eiHSOCv0W
wDK4csni8GstRDMdv3Or+qgTXJiKKqEWpcbeH8TizA48CkCcF6ad/7vr/CrCt/TnT9ns1sZ8DoS+
PQT+noMpOxdTlDqqt2OLwmMVZdmVVnnc22j7v0uRLPoX2Ob4TovggLxaDQ2wc435Ej0tqFOrcJ44
qsu2gsgdvByLvuyGbONJDdFe60BvO7vSDQy61CmKWXSUCaGxsFS0T914Rq8NTwZK2nGAdNXzgi37
ZSMg71qxLUNsDVggcXtmvAQlpEM7PL+J9K6ZKxPEaf6DHDQV8jcscrdXvce1BKwpKOe2gmDNer+6
rI44QIjfSS3sCNYReqpYR+WIh5KFTAtz6QgXX2toZf00t0W/eqWleWJOGl1XYVHmjE5DBKvl3UHL
cwCgpklNJUf8mV5hsWv7U194H7jLp1ZteLFY/Lggusf91b34VxShhJ86thYhh5+VDD/C5Cm27mb7
UTXjb4C7+8Y/5HTKlktRLquFZugBqXHaJaDICzKX5s4412oVR1QsaYvTyDL7hAYDSoawuMEVW/1b
ourgVZufuWi1W8qAsFRGjfX1zf8cAbhpOFTiZVKXMN1R4eWhk75F4MedZkDiHBaBKMq+fccaE4H6
5Y0l/t2369zjZBPFTPVxRNmMbW5WJcOFB6liOVatnjqFVSzwtNueXbgub9rV4HpXCzFmgAaMyY3x
F4Znw8EEfqbxQxQGrz0+X4IHNkp7fmHhFV8tyMuSS+VYTV9NHlcTN7YYvEYO6rD5J9R7Papj+/Tg
B5OHHS6dbcL1FbOpWUwP7vhi2VXsrr+StGmD7oIRoSVCDnQ+f1sQw+n3NuYXWML9NqtmIrYJMyUr
wHDIrpsO+GS6eFYewpAsozuC05wbO5vk1AAs0Pr4mGn4UAC6oBPHRm22HxX8u1rYUYM7Nn/TfJRf
IBrISVSYOSoIS+4q4NiTBQerjDtW+oP9JPK96e0ta7WJgVv+e2ixryc5q3W/jmxKS10hbd6wZd4m
htgGMbN4l3tkyhozMgssXm3YC7M9CN1wv4OtRJMqy0fNg3h4pF2fahQlpjwMBufR96GGw2d+LBJM
tbzufIPjWwb+/CaQkhMTCOx/Csa8hFwB90wNKHkh6bcK991wmpkdklTvu5FbKAYbdcQqaTQPzPcT
5GexfPXljvHfnutTfhs8UIC8iDcqiKqA0MdYhWrpJnh241BTnq4EhaNkg2mDdoIyAyMiVLvyI/0k
KVM8lrk7wCDVZFN57gDhS2txk41InzEswth4oaY/9ec658BpQp8Zzm4fr0M/MrFQUraMA34nTkFT
lp4Rv6n1LdP7PdQlSNrP2wnpzAU4ipMDc1TzuIk2yVN4cB1O6lZSzPNO1edf6ILjDru/Morytn20
g2HlJLdebX2zilWp0591ZCFelxjBtYALkGMrPkgHrSQA2Kk/XfQ15J8hD+0dP8q4lwdfglBGsQ8C
WaTmlV92MHTV74lqMgH7Ry3DmzOZvB2VSzbB5tZuLdjO+wLdWR3eZtT1oDvGxn+sf5sYdlDD0j0L
KKg4GdLQmxLYi8rtndcZRofvtq1z2x5OzbtA4E6oi3C4HnW+jMpvY/cCBiZ8Un1PSB5DJOs/gJ9S
Bilk45vhcpDqVqxj2V5xEUN4CTDGSj66pNY/GPw0PGPCl0U7FQHhu+lb15jHP4Ny0PegJ2cNVhJr
55ZM2QwcEjiRE8IezQBq5cYfMMjdA37BcCkIJMUOrgg+JLTg+WIjmkNJQQYIvoJNH3NK+Zi4Sb7e
3AwUXTjA5dc6GxwvN5Tmu7OHTl6QRUxNNYonbpb33G+pominfSCVi+zyQjhPqmdC6VGcYHg1pNpl
RvwJe35tZgB9YOrn8T60v6uWaPLYGz+M5xRaxIIGjnPmIXy6pV4dsHdtSk+Be5SfkHPCCDrZZspV
qChjwLeELjY1+Lcf0ufF6bIH0j17EOqYdiV1KpyIv3bJV0EHTC8l7kgake9DR+2+5JZ23+Vdkh8B
edslFs/5Ld5IvWq1OMcpHiw717mmcQJ4FNPRc6JxArsygGY0lBGbPLHagfqXs1gM/8wcYdJuKG7i
vko2+FUra6I0WaMgQUckPErkI2jUrlQgylbjrcgD/imXLJ4FN/Y1o1XjhzRlehMwtFHWrKQLKRBk
KihckpEev1QZ/d9UwVpEm0zX36Mq7bQ5KWuE6UnwNkD1gNFHtsynxNd5Gjy1NWfCgXa6d1CzKycC
ZIyo5l1Alir8xhp7oHn+HIMX9RrceDamd/fWTB0i9ahBuzDaruW86ioIk+f/o8SjqXiUIwOyz8gK
ij0NQLq277hNXhjVdJDoNoy9Lsgw/BfX9iLYb3shtVj6msNNL+OoGhJhNS2HTdSLX2YUjYijIUzb
KAKPIEuT0f5vmfucYQe6WsvfyVgngYtqJNiKAYzS5t3pCduMsy+gnFBRCjqdmiS+gOhRWHwIs78u
Hj5LbNw4STHNb00P3+h2pfH67c5gRqmXMye1yWdJqMQQFwqaiin5tYH3h/zVnqIFoFHAA76oUbJ/
jj3LZm8A7iz7C6lqZ1xYc1UqgdrJh2FzqB27YTicKZwkM/DjsX4DBNX4no8RGEfFMGMd+gvRXUL8
afH84q829F5WeZmOCKZzvG1FZYAsk8Be6rxksPqAfTnR45D804RrbRKxDGmrFfOHNZXpXrtOKIJ9
HOwj2xH7vYJ9Cfyn+ss5l8FcXtSUSOAG1aq1cP0OIUYjAzeOc7zlPVVJF3EiQlZDOyKWp7SqOicR
HdI+eZpompu1w5LXtau49hX5SVbkOSF0DfS/5U4cZNE2maDnJs1jyk19vRR0nimhJarBayoGRJ3w
vPhsz1VF8p6eeh8xNBNEy3pyYHBGK0SPcsJOmAvB/PUCZD7dKyU0eL045qZ5P3XIsOhRGgF36Jb2
SDHOzf7J1V3u16xqv1g8LjQCMgGukosL+9BHfdcPSj0pFtwO+bM9pkre2vH2zavaoNYupGdEPkre
U3MT4zYyz6Y4wGkXDUG2+y7Jz+20PeYvRBRMYkmLhYZCvwY+nXJRPdQWl0W8px741SaSQqEr72Fi
I7OaRBIIz4zW0a9ULkAaRRgauvti3Zs1/Tj5raZGA2jZN+yvd1Qs8CeJBmbXPN9wK4WJvg5coZV3
ml5PgaGqYTMsZLJEOVrSqCgq6VuOdmM7LKKAXn+mDTPQ4ntXV1uhCmgq7Pl4cCLkx+EaXPTeIBlo
HrRHEhIxcu5iPcFBnGP/+k5Ln6+XcL4kg1UXWeKrrZvrpvU77e+U9uiuEtpMdgwEDGIBv9BgA1Bt
0tftaYbMi9nwke/d60hsmwgKGgEXO65g7huVN/VXrbrOXZJWtgqFL1z34y54q0VORQFJ2A1a3yBR
mZTC/rkCqt//Z0iPH3ih01K2ag3s5tUdF2dqUeME69TgN99AFfuEYYpySJ+nn2OuPaTC6BtoSqXw
7MNBHx4zPfRtXYVRCWlbjmqVlbXAS/+WHUxbZuKReUhkfYC3J6oYmdP0vOBGR6fVNjE9AKA4QykL
lGyhlyO0cXANh5fGEk0IjpmFGMf48I6cFPjGixyhr8lLuDZfxcEYCzMHqN+vmcCGYIjj/EfZuh+L
FEqN4ylKHZ2E3s9lCVVS0lMLYLOBaI0Pg9OLrzOneYyB9CQCRazEaqNdIfecAU7fiEJWAzT2eu1o
6OPz9Lm2Se8/LTHwpgGOBDab724kiIk0HSx9GAMCNE7gLj5Kl1XCujBxi54fHtQZNkGDS05K6bjG
nw0mojcCA3RNmjE6uCgz8J0LThV8Ynx8YH44mt5sV0kpsOHhbbGJjJ7cyFm7bws0doXPin33cvrd
DP6pVgtgGDh0uN1yCxXixcIRqbCg3WLCHsuwK+hcO/p+BnofSdMhwmEK4kxkGgqC38BLRqZybQcK
AmKS1uPZ1M+NC0CLOFoK8JrrqcRqhuoDZHe/N/4Dqk7x0m6Mkm4+iyn2oOJoDv2U6Mfmo7F0DVPr
HzEvHH4ys+CJBxj1nQorYy6VsJ/8ErzmZIFJ7bAiaso5Vq1p4Ojf4rDYq8LKwzsApR00L3ChRKc8
cul3wl/+qk+73Ik0KZC4POMpn38z98pGo21LPi97vdqFRRfbRrF3zAB/pbGUOA285DFOYxyhFeus
2CzJzaLE6J8U0gWeNgw1+ASkoP7lnk+jbY0IhsywTLsNUmaE+FxP0+LSYQu21RADwDXVtPndjWk3
gTZxPX7N+WvKFzg91PNTwWIEApQtZDZk/m+I1pOQmO/E7PwCJoCVdCmyVVonh1MAxviuQkPzhkjN
ia2KXfMT54J8axJUFM6OSbXwJFmdZXtvNeIcfWo/jLJdqw8rU/WiWSmjHoClptNG5lv/ukNGxeTI
RxOF8UfFRQR0uFZ/C0x/zE70urrjG/8GEKDlr5PcRVyp0Xn7QnsRtyyyBI70TsritZYN+x7gIhCs
QFFnapODBeTlbqV8GtHAUq02EIuPfM3VvudLlIFKo/8H1HMwXkzu+/DJfdNjLx9oOFC2tU5Eh4cC
8Q1267n0G+lFGcyhQjrhrMo6GIxQJ5So/dNzPf1otKYp0P+btZXABHws14JSIx4q5gG1bWYgbi/L
DZl4w6eoA9+du1CqZNVE4hlepAQYZ9Bg0zGnpsiPuMfyThGZ1UbHopsk8vFq3447uhHBF+Q8quzI
otldnqABmCY0Os4Bsgi3UMulI45cfA40+KcwGtU0lHxx5QXQ4Rm88TPU9ah7IrsVdJRq24Qm+Wet
37eD8DubXqhyURYop4PZuFhWUoGPkrJi6uKkyVIPNFAuzGJ1sFoV1sNR1SVG/GVsnUztTvrnFfnA
lvSBWHeZxNhflRE8fFVIMuR1dkBd6rPWmfR7alJxjkzWO1lluJkxihmoH1q5/y3DYhNDEwoC0eRo
pe9YkgdBQ7YmIX6pNeoNSrymDC6pL6wCbNmM7G39oVGRPQFrV88mrEeQOk3moGZ8Q2chp0w1Hk7B
e1dxaqIsjOlULJmYqFI64FbpcmQyQhZp93mDE4IIgmWm9MSgGKcEvVTGiDLSxmzLwTRwy3rLAoxI
N/4aL8BGWZRS3Y3OmPq5z8f/adcmQP1CJQr6isJhE+oTBShgKWhnuJkbPELMl9iB1hzcR1qhKUQz
2HF+sbWXKlrpsqxzWIvsV8mrGz86GkHBUAjz+3FfY66991GUU9cyujQgU2U0/v8ODoEmrok+ldAS
mPue6agw8im1P37bD8HCk6KIDonUDfDPYlhQwOrCfLCNAt65dbZV1WDq0PImDgwBKwYRmjUnJVpG
dklKralZgFCur6GNgokzu6f28clnsIxtQtlC0dIOvT61fZ0ehrfYL40Ui82zWtGo3Y0IsTvjt745
85mzgyI1p5adyvyDmqvLcjtghvsSWL80CPVKuRL8VlVTMomdnrv6F8hvSDIGH0ayXyND+DrZrVYc
O3FXzQSYIzsPlEtQ29zMMmUdPuFhaVGRTeYsxcDwssBVC5G4jOVdNsJeqNe7JK5mAyivt0Lsze0U
codv5imlanpAs+M5JWv0SwvFaUZKunWC29Ej9Rn0QiTi1OKww9Vz1IWBMZnREisdLOvRnmBQhpO6
2EWKadjwegUCrrVJqWakgMiMPu094iZp04m0jMifj7wOQOLsm4cJLq6fK9ss6P7y0SNUqVSDE45P
vsOtxZMcUYHygrKKdHRNlQ13p5ua7L1Q/xF0a3YXAvrNALcRQgWdhtaDhehh0GaNIrjMMdG06cw5
e3nOTtW4FiiJgwCP0fNMOZpVlmdyoZyKgFs5L3HcxwNoeD54AT6nm6wIT4Q2OvbCiVxnGOr8FYZ7
qSaZ7fX9h9KYe+4HQd5n+X+rAkMVqfJxqLk6YjowQiieGSydkDrkHBBLkd+Zrf6lCd5sZV//V45M
DxIFSC/uppwV3sn+mRSjwTk0dmhc19tzVaA7gdZdi5odqZHcqhl3LrR4OYakBhCRrYNG29KkBvRF
t0z69U0H6u2NhIOnQGA4S8zbJ3V1DKOSUOfsFYZFUgdLBCDtaYMl0PxweBpz1fvkzLuipRzOcV1Y
KdY4tFMVxJ3IOFINmqOjssMcsqqja4+DJNqfQNrMLHK+sSOsit4cLgxzB8W3AeN8Xl8KzcBfj123
PPxdm/OCKP62Dzzto66talGiC2kVzbkx0qyIsM/bDkpPrIDWmjjB9Nn5m79O/0Ha7iz+u9Bj33Xs
NnHZZY3OpUb7EJPURXODBiGqa9rXUb8742mNqhh/BxeQvK43P5V4W9DCGJaOqKLC5eAMlqgkP+h/
wfuX/hmLoJ9tsXrUXxVthQ+oSPlroyV3HhNWr+ZYfVJv7dC3SkR8GIIvyiryjycmM2i9nCh4zo29
UiS9CNxqkFg5wRuW7GXsgTckL1xSt11H5ZDCGa3JgpYJ8Bn6o7OpjnZMtB6BHBzpx6YKVs90TpA5
bZgkzMHUvKRKcpBhy1IZb84NYQWh9IlCT1Lbutwvlyr3cVlM3Ncx4wxYd1qfQjair5x08nB1dJu5
P6+Yk5zh5F2HvHtNcuLhmirabfoV9l+bmhwA5zJ53uXlPsaR2TcxZ/hdsc9q5NkqlNnmwQVgW0AM
3xHrY9tPcZaowMMWIR8xEua63CFjQQbac0zy7wvcfHyX1diJl1B7gxCeMV+MAMp7QHNAa4ro41EO
Q2IiFEscNo4cW0X5fw3Y9ZJgZ6rBQMaFZ+TZnm6A5MGwCuYIibu+JfeojgwL2ux9MAQTygHqNdXb
SVlY7m13ogwFmyuOyqeoOV2GLHNd894H7Zvs8k6eOrHrkwvyrZyWan2QNeJc6qC3bh2Yl/geH7Qk
NZWgCngE/lSrV7FzkHHvVEYbgAk/K7LByySnRS/uLk2GTgkYx0zJbzSx5f23Au9gNgZlAvmlZ79A
u0hwJ2c07UXxtEq26FSfHXic0gjNsENexWTSjrGVMDdM1+RlQwvV8QnYROr+aTmXYbEZDii6Yx4p
0rDZoQljQFNWhv0W+ilk29COob8NAJOql7Y1P2NLhveMEBjn4wqFpELObO6IB1x0F33hxKuiOb1M
GSr6KIB92OwvHZuj2g/Rs4nPFDuFqF5Y58qaJK8DA3VboK02JT0/RNnlisDTSSRbpfYhBnY49k9V
GrIqBfwUGRL2a7pMsSJSf7daf703X8K47x81TOdBQ/nctDs370BEJi4TdW3rQcRSiBp3/SE8a12G
oY4DQbiT+MxrgzbWqlqxTOkeVDREVEpDS9/LMMjBoBfPmBDRIbKpKzeceDsjiPtVwVy0RT7OGaWp
qEBlYvOh4i+NNIHWx+9q6jThMmRGuFYJDkfISq8QiSdHwcpLS3XJ6uIid2OaC1magm1zUBj03LRx
iD36FH8tckn7wtLRpvotlutzlLN6zzeARPXdCLojb/5jyUgj+M5xbue4oLY2xj3uV3Zmrcv5/K1k
5v6seDxahXgx4VfIdKxOuxC4dNYhMlO9WUSQ0hUQC8anjIsyXUugZxc3XmDJU9Wc893Fui1gaqf5
3gPawWYhVi0oc3R2xoRgTEQ2rnVG66/8bSKrGv3JE4qKNW2dkSPZmoTidxSDOzAKdxhuOyGBC6QX
+QDetUm8OAR9BO7YPeGBqUFidDrkGri86q2pjoQNxRNxLtehMuaByIGiSbZK6iYmm4+gdmFQjzbI
YwEEAgjW9LQKcZvv2XbSWvCKOXNAfo5ymCN1c3/Om1Cjmu/keeNQmfW6NsubyXqLefXi7/nwjOZp
1dAXcgG7Bk986k2DmKXp609wraxbHuW8RhmJ7vmGb0kirUHKb2WQJIZPzK2JUsBxAZyTFHAty360
u+T8DgqQ4JYwKyh1vFc6kl97R7nR2z1Ao6yHxGRpB7nz0aOFJE3CVZ7Kq5t7bm6HCcwNzTxu7Qg5
tGJYky6Pg4Cz8qOMRXkHkTtsC+c90jRLjTdFXhOSS6QthTvlqFzeZhrAJ2cKFzlOJwO/hRRoDkuD
0ffiZjgc6gaAbgB6MzS+xS6Vb5rGlyXbIzZdtz7rTn7YfENBjd3ruk3Hz9DwROPfLKPLHlqwEX/k
ZeYpYxXJ6WiM/yFp/t3LQJcAQ8ywjFy00LmS8AJv0ShOwd5LyTCb+lIQqrj+CZPvpvCBnt4DBwQg
FEMduJEr317+PvGvj/att+bfPRbS7pZT2dmF2lcw4Np5KZR4AIzkbqbHWDHIMYooXNM4adUTlAvH
ch3FiCt0UJjPK2+XhpolA1nOi+q1yBX7rIYV4DhuD8v9jRmbzIjMMO4yUqeqIDTSVP2FJMRl2dW2
LSpXnksCT09DJvb5MMG/jgaXyVQeMyTEbzXOjZnwlT6e7h8IUtGfy03LXM3Fkuf2kAG7QijdlYSK
L9moEVMz9we/34KLKW8kfzNjSBglvItJipWvp4+2TcKMxCac8iSJCXxD07997zkhwG88UbfZ6ebO
cKpQmwwXzqTdS1/FRIyECJk94tf0NIW0e2SjzyHXw7lZ7dP6gq+Cpp8ed56r5SJV3MIGaNSoo4HX
88H94TGtFLy0Gca/VJyblE4TL1YOgKAUYpctGZU0C64tUwsNhTl0/SkrPR5QgJzQ8WP+PkOYYbRJ
7dMDTvBXCGoh9LAHqCTtOH9gHopkmhsGTY1dqdCaAOT/pkABGmzbBk8wZZ+avBfJ0oB3AVpXCQbM
guTaUea1Z5ywDqFOFp3yX1nMf4UkFdQW2DNZLEiQVD7sIrlk/ouSDwaDJzftLl4rED2yxF4cqeoY
YxhbQLKvAXQ53PWZhyOtW+LgJ1dc0Mo2tZUHrW4kZLvfEkFpg7S8nFwXYIGgYP2GtQ3uQRvAKBle
+A53cfUDZaBXOiUPmiUm94i0Ir8bnaA3pw/E/kVeME67ncxWR7QinhdEOli1VDBwrug5G2QDRnvj
Tkp7BjmJ4vLQECNT+4MmsqWIZss1SUt1KQ5AuGZsNAIvvPVAoYUnJdlKtiGVJ310g1soKHXXiznS
jKvQ16B9BwBUQ4PkQG9dNQkmEGQiw/AnfP5Pw6bcpPkymuLjDlywyECKFZMkbySseLNTDRHP54lk
CYTtDpSRJhENGDi2XLuIdWzkGRlz0qVe9F/v7J3uXPXYa4ZdmToQZJHZEz1THKLICPE8AINYq+5p
4eCgjXUB6hxbgsrB19cj1fbRVme/W4agsV3h2q47urR/+yxZAwmqOuh980o4QDffbwChU4XfhJzq
hXCtMWXkajKWMrZSQlykgULG/D6DGxnGyKRzml+zHNfrGY+YBf9ZWltPW1XsYd6MUhEtTfMZnRWx
y4aJ93JEDnm/STEszwAUHNmccekpml4KagUKpyIo7KpfS0okq4Pg2wcbO7sz5WHTgxY7dW6GNHpD
l0nbKVYH96RZ3tG6DPRD5NRbA5WM1IFNong9DOniwpMNDrZ50p6cZyn3Y04jWnVgo3itrmWs3Yf7
1bFPi9UPObDHTgw3EpoNVdMY2gjCInGyCZwPMM4HlcFzdgaWc5wVhGnDCT6eA2zkIVsyh4WfGdU/
jc6kmJnG839xBwUDest8/akRuuZ9yKPzMzrXNaei+I9YJTD+HwRwpjRFhAqZc7NEhW+/sfFaEviP
Cp641mqez4DwRGGOQbgFLFZ7yerD2pE8dHufAJ1GS8iqTH3+dNluCzw+QBd2wFNf8m5YaT9Xdnbg
b5ylF0k2RSBX16qE3gj+7TfwkZVJPXdQt1ZWVD3qVX0uQofEwR0hcu8rhwEbjn5Y2+1VJBRjzTtY
slufMpjRkGjyECrWII7NVrpbp1u0vwlp8UErQPAX8mNehKJ+mm/mxgg+vLCKJSCKQF9eYoyeBaOU
BKOGB7QqRbz6rGblYc+0qjf4NqGKCfFi0py43J8H2+Ncmeicot9YilH5HScPX8lh86vCXME62WiF
7tByiaOmOn5SlgN2yh2Svpnjyzk/37NVs0xhPWOhhRuQTWHtt27maWce9hOz7y3jKOEmElBuloqJ
1tNFn2+0RuF83h7ptLl24Gawk0OPDxvqlCNg20DpNeuoyPAEFcaUJVFLmecYFSmLLJvz0yxU4W6f
TzsvIabqO7cR6DFKP19+g/18x0jHQi+hPMtWD7Hh0K3D9hu4Oe8WXe/AR+cXgiXIXSYQVkZxzkv+
Itu70a1l8AyrdWx26LplJBzc2gkh4M7rq2dbhLbeopbtZ/rMBWRpFneasL0zhyOEMdH+DO6y7xWP
CJM8SRNuhwQcDCuKJWRdA8twOJJEZeaxZUx/g3ocn/bUergSvtRAg2yyi2I+ciRDHAgFwJZu3cVa
RC5eecaSlUvK6uoG7GDlzgjG1oHQCno3EsyxCPFo0+Ku8+ad0GB35EQnxMihpjNwaOiuciXbUt9m
CY/ZIp/qykoL6ZlZIq7Bqb8shkZF5XbFxA+L3nGphThQb8A42hTB8WjUgImZ5n5JrKQsMR9s/y1P
1UARcIDXjv6sNp24hNygo95BQ0c05eQwAk38fIwfhHEx9l6KXzE2H4gJV2W307qRSUavdThhNPKA
JwCRZgEtA/uburrcD3rw8PwTqKSTzuetR2HPjSP9PmMa5dlEUylBf5D8JzFePgkg8seWPByLxW2z
2L0B7C9nNF4frpdjaeg4B4UxXVGLewEg9uTHUFoY4+a0hDnVV/TsKMiFBPZySM50Awnl2QGgEjU3
cizY3o3a/5kji7k80ILf2Bf06aoOUZELX7cxUGfnvN9yEYktRzVcOhRl0aGfk7UmRkDH0G4wJiMx
hux24deXOF1d+dTGP+cJ+TAKNRl5DfT5ROHmRTaA7pSeoPFGXsLo0hrqO9xJFtKeOmsIcCFR+jPx
AZX5dOn1e/w3/TicYhuqRMukdHKqJLCwvM/xwXQLaAHe/wNnJaGCzfqNoxF+VLBHouRjwo/2R2LP
IOS6IVvM03z8vE4TmnLTeiQFeIQ5lgc3lFXEMKi31+v7tQTSQdj5CWmYhZj8PHax7j4Ulgh7V59q
nHxlINBSOmDIwuRC6VPiNQEUMFdHHck8kodHAqg+wgLebH/kYcaKWcjOwm7qj9E8n8hx2PEaVzx/
6rk2Kfx9aQzRtPD0BG+C5tjUglGft8R0nBR4GUhK6UXqy0sOz3Oqqt+IU+IecnvxYz0Za9COlZie
z5drArsmCp+p1+AVWTy8/m6FPeqhS1rtYN9N7Kq0uyyA/ulfyyOOrwoYxGxVaChh0ui+VXaX1zIn
+yWlKm5QxFb2cowrmYmzO1+6U8I/pAoy4h0PpIUEBvGizXlvw2Xsg2GaiLVZrKX1V0pK3JHPF8jK
zpvSBzXxCqPCn84uHWRQLDlTAUk64hXMqv9qBogQGCd8pSkOjMMM7U32xvPoLHbXRckGa780i6GT
1n/4Lrah5S/Ha00AlNXBjBxY8DmdIJ54tf7DIg2FO3MZcRaTQFKln10NidrjdN1+ogQu0iUKeLi6
uwDEQv0UeQPyBKEQPv1Ej00ewMAEsCLvZ9k9crOJ97zhf2kB+adpRpT0yhU2sJ3ASUPUxBdYqok6
sBl3QUxJx4e5+n+8bjn2jheabK8ot8DRg5d/jr7Yn+r+Ls0cY8GvUkglwDkRqmY2wpr810Be43EO
dvzPWWndDKxklBnziDRnC3RkZjjqAdq/4JN9FY9F82s64fkOxbfIMREp82YS4RX3pihtmUvb+9lx
wCWRfuQrIiugp6zfctBzzr0KF+Lf1Ct7dGa4kmy7/pgHxFn3IW0NXPdQ5s0BK+ESjPso/kfEqRHU
zBW+rDD6n5vP+djHsnJFbo/yr/X9J6SlI2URVZL4SUvMvdnPWn/77F2+bnpclSMqCYV2GniuPe9Q
WhLhsfdQvoa5smensIUnANOWx6jjkurkTV18jlN2KmMgzt2HSImDOgERVlFZm6TLcKsgVlu/Bv8p
K9pZwX+Wjd6jvW4JzySl8xAVgHBvDNqZfZD/JRTHM/9yShyzWeIzr3RusNJfm/grXIBZkFUBQ+Zc
gVbS3m7fViaORRpsljT4eiRMQ/NRiJx0pD+9FHTd43UlBFGvbDKLv1RYeM7rbpNKzsoLvWKmO5v7
M2Bx7nycg6DwcXvNWR4beaV9IOiajw6z3J+zgJadWDjeqQCCWJxCxp9b5tuWStXF5Gt/JJc+I99o
dPheRES95leeB0gXN21wPUyzHv58i0gKGVk0S6f9FOC2qme2kMsQcFjoxQjeEfALpz/EYz1gudkc
eFPtI91Go9Xo7K33/gS2wAjFbWC/69/PcnER9rAUE432LZFzmxCrzUKBrur4x2JnD9En3IZR5Y8u
QhVJnyjWjpwR+/TN6HwIKJuuPHLwwzMIV75ziDvLiqzdUXzCx03BnH9UKuWLd9Mu76jWtUsFNFVu
HKsJozPRJykpJwd9YcL5fbEfwO3q+e2eF1R0tbnluINtOU8W085vaHcwy2LxRDl4B06qrSaH8bzr
OoeuuYYhjilu5skOBwxxtGMI2nmM6l+CWQmmdOga4HK4xlTt8kUCRzjhb7kJEITceC/pgO4xBio1
yXPzvsOyBLQy1I9Eg4o0j+iTXTzMPRTVX/8EBNICYhhcn/3Boy2b3IZ2SVzZmQ/0+0hrV9r07rAB
8yHNkVWiPtqgI6IFwmqJvCY1WgKbxAXeSSrRaFCeBihQePvbyIuMOFHG9mj7XIpklUo1Brn0Ei6j
W3yYw/EJF5Z8x/TiwdmteLxMrRadf4JF6ApwipSgV81WDlyrFKsV5um54bxMmDgdcxCP48889pei
Rpd1Wqt0YED2X1pX3qG4mQJ/9fNzKqtVF/jXFZymwS030s9FGFQ8Co+6Bur5VK1aSZISgHbMkpd/
EgciG26rvlg8hMWJLQFXSFu8Z3rI8iwKYhZTRuIVK50uJHenruHiB0Q0FRYa4Dh2YqI3nbmF3d+v
xfPDVYclRSRwUA8slvythZJoV0Mo3A6AclRFMGAEF1HH0XC0RC+bw8tiavlqZgVjOsa5QkN7sC+U
AF6uVoq+TGv0xEmPgDerNAezkWDumOMljdSjDigjqmtHaM/3bUjn790LNFGn5eIgX8Qz5c8sUIFM
j0AeB0XPeNcn8z078KJ3L8a3HACPzHZAj1YfDJ3ShZOt/8ztZDlhJ9wb59wwgdsGPeqlUxg8oWZO
AiGnckY61zphbpqmm+d49CQQY4XGuC8wVTn5t0dilzVLVKe41L3lGbG1YdRdlZBbsAD0d8tQxujR
Db36xOZcBwZwl/k87jiRiCrkHfTlj0Icip4lht/EAWGylgpYD6Y9jhVsFpsC+ce6r4stqy/H2/bM
kJQ9gneAisDCYwKNxcYzSiMNH2I8fMi14W5NPnwMSYz/YncihVrVe7UHUE4gMXwjor/yUUxPsugw
3cAXzMbHMRYVT3VcZK4/zLHsTQwpOLZhz98su1NKKBPpoaxImzwQ01EM9hVkFpX/OdUxRHaru4vj
H+GXEmfUtYUqONRQ1ZweLK6YFkdXJfqZd2w+BHqa4WFy/lLmfEbkop5qNKHT/HkpVAp5gMjzZmDL
mAotjsh5GuqknxTRd5L5FZ6V91DUF/+TKeNJgOV/fGAhcD+UnlJr7hW/oKq5J/QZLoMLeeTNb8Ny
9BkrXbbFyle42EPL1NaQJGhfuFC7kPM9rOQ3qQYeGszx5TqkqUMH9X/4G6Nv0D5F8+YPQquE9lBG
C37XLi1KJpJmj0iCaeTbrVhq47MsHlIOpUnrnErlp6O7SnFHD0wwTgro5U1cpOXIdZ2HWkmzi6pw
C6KvESiNmOofkaXd1DerN8jiSODjhpQxSsCycvj8/kG0a4aYaH2Nhc+Eg+Z4oRrVgE5eWNwaHWNf
CJ60b6g2toB4fGxA2sBG9caETPPtks8w293UtOZqYpoO0IyO02SfjIPCZpmxK7Pjrw3DnGoX23q3
bSGGa/F/qR3w6LV0tcL2XJj5Rs/jX6hNUikKTUJtT8ZX9JAb7LGYE5ocBwSEBhMH3kS2R46Ec+Iz
oJeUeftGIJPMKIzzFGQdol52IvEYIgY/cuLNFsJNx8XERHBCpWPRxy4RLDj8zMuIxDoaGw4hA3Xr
BhDAQJ09KpJlT3swXZ8Mk63S2uvuBwT1+pj4VvjpUH8ERE6hmsLYD0J4yFzuiIQ1/o+ByUN+Mwwo
H1ZE2K+ho78iGuAkw05KfcVFbOVe4o55U7TOqHrTrnGJyAYRIxb7nfN0BzHCf6cFxXL8ccXFbQZ4
4BXeZf62I08RTxosWCM/JAVH1V2DN/di8advvJtXUkPUQ9evCTBe+EtbL7xSqTqxrWnHgR0dHYjP
pJ1sYGQF5ge4K4VS6dtOBVZba1qfrELkglRiBjAFrWm2PpgAI2FMaYEhxJJWmpKedAoEPCb1pguO
mk6NUMTtWvbgQs/ACONb1WW6DQsokVxAftXGpxH+T4JhNrairXoogQ+UHw8Wriv0cZ3RuFen7RBG
KbN66qAlmFQ47U7lNRlnPEG/RYW89rkVW/QRJBriuSczGkBeuEjStquCIkSoz1NzBVARQ9vF2jAU
4N6mtuw3W3AENheHwR2VfbaMtKtBnMHrGv3NtLTjNLpHm2iwYRdJJ3fanwLGsa9xzpevJs3m19/q
HDrJNedn2uRqCbAqEyG69RnCxXE86K7zI+gUeTtytRTGHMGOOGGp8Bhb85P90ztA6DikBs0ix/ML
dHu+IKkITa82uGUraIc/L47E1aNbgvsGi3UeDjFZlL3jZ/GnnGDyD3V4mwBzk+UOHKJfWxH6emZc
63CooV0bY/WVKGoUe0p5No/wrK874bf8EMjC7ij1dUw/izgyDkyDCsvVPQuzxKYoSPwgl3DAHMpb
tLQaNOAloYhuBLTRielZs6XOwgp66OQEP3PTXLuhSw6mqMXUyfAaLjgokhOZaiQI4ri+9JnMtG4E
bvp3GL5afapK1GyhEPwVPXssgEQ0hQTcCDYehSg/3stcwm0wbSSAvZLaRke9MYOvfEzGGeD+QlDG
ck2WJREf18CNfQR38rFTm1DQ3l3S9dT7fPI/ElR90dsaciJr8b5sBoILLM1FFaDUFSRgQZvjokTJ
1HfCnUsECBx3R6TtTVXUzqp+ksblbmcWSgLSJf4xailjg/6HXAE/q7YpHuN2H/aCslAGqwLynS5z
BhOPPrmujMQpbWqZfMHIYW34sfbtp9w1/VRxJdztt+a1pAhHtesT3hohm551K3bisWF/KQ9XduwT
oNbYFkTuJmn56UoL/2CG7WMerwpCz/9Cu3gEjKHxJspDF2I6bSP2nN5CyLsERoZ1u6oq5sj/6EyT
RlVTHQ1Q4WwlSecijYvk0La0fmYaxA4oqiZXX0cFzT5uZhb84AUfj+B1JYPqxcYsaxxziCmra9NI
GCGZUyyN1Lye/C3JGFfmW/Qzdi3wyMaij+oG/adnE98JNS9VST6ys66LcZvgOTY6rBUBvCgWQIbj
fdrRdg/peVOKZuhY5VB9FvoGYpSOiCJbcpv1UtFF0V5iJIq6uohjl2210Yc5HLVJaR1IrO3PS/fZ
hv/iqwEf4gDhZAFDn1qpwKdfznfAV9HzSwyK6z6fuK3qXTXSrPWq5w9Ut9uSmSllte3aQz3p9awf
vZn6xCEMxo/X6mdhzYDA6Nc58jyAe4t65tS5n9UPaO6YOytEnU9s3UAgrtjliQbENenjV+QBbttG
vSSGkrUwqvbaANjGInp4KtBO1gOlV3sIxMUjX9xuESP8nOnUJjrg7h44Qkiodn22OgCul2brMHdm
EtJnM9wBwPjKkCUDzOhAHrORN4dFTQNcsPEKcKNfifZPPoq0kL5e1j4nYORaWbT8QY0cPwm+i6iU
VrngL13c9rQLehuHowqOFNuTmh3C2Zo1NTMov7uj3d82AH9gVqXH1OAsioBA1Fl+3j6AgYR3r+Uh
Xdl094kpszcXqbDrstL6LAlrlb45KTYSDRjQBAiBBgXmV99b2MlKsu0irajCjKhb/F0svkKKsHmS
GHqUipK1mUxsK057RWtgodHWDwv6BBhs5XtLu5bdBX77q6xq+P/LuByvSoSPo2g24W5rMMcBDLgR
5uW7SQ/m2R1gpMcvhVQCRkyRIyLhHmV2Zypt5fs58WSsxV9/slxW9pCa7YWzbZGP18xQEEOoib7/
bYEjyk6T3i2aYnsZxSSHW+4M3QbLX7FFi2TIMDpf2jAxV/ffZsC+wOtwxE7Gn7FHNScnnhCQIxcx
DAiTTaR8Zewm1AjT4sEv+OLHW4egD7sFybUOcIIShjiiTRhPHgF3NZ3TGZUs9aR12B4vkxh+D9wF
jAAExMFMv3H/N5dU4jyvMChZO0YvdH4wFwelA9YOsNPAWjkso1GFPu1U5sErAr4PzGLQH+nIsQQm
MoOFf2ViXaVzcVnncpoBqjf0kOqZG1ZoijARIFjUc0ZSBn1iowU3RPN+n3hDVYWOKr54CAJYRiKx
ojrM1MJ2WkswPA1q9dmc60uFDjTbkprUbukfUoEmHQy7XLCrvtBowLWi82kG4JeWyL1tz5HGRc2A
N7JIhlYqx5mm7EEu6OvyuaLCZM697rdpiICI3di3a1SZV2q9qCYzfAojcRiZRaZICzGTHzaRAHRp
zKuvM6X8K58XhsrNbDU/TU5s8KZKeMAaHADx37isLtwxxCmgiVfI1CipSvrL3d/fU2kVdkrL1+eR
EQPmO4YpKcjYgSRxqAElmajNyZZbp+Z5H0aQTzYL2NB7YeuguInMxNaJYJFwO1/fV7RK/lkY4DUM
nJU1aAXa1X/xkQPOrkaypmFS1qFBf3hbngIsE8OGNgB130nAYESvf80WDkGhi87COzICmR2NnQQH
yO12xIjutjKJjmupmoPxip5jgMjD8qBQ0OOvj60hSHwxNe9LVLE8itQ+v+r7NMa3Yn7INkssQq4R
Q777rC7qXu1nKhvOEYXtu4Dcesl+hu8/HLePAQleMWA+LvkgtUzPNhhpuZ/l+YRGko7XV2Vd0eyN
oOLfHQ2gBiMb8grOw34kIOkyMhgLng8QD3A5+/ANcWw1MHI0djMOb12xPv5jWq6tXQnNCVhYwEp3
y5NHmB5F9c/ypOvN1AfWuscfoWrZYcxYftx0vQPKaHeY2ujDPruku9LBWWBAOp3q5br6wPlMBOTy
eA4v/wJO3WSIeU5BaU0IKcv5b1a9wfgGKxXBvGJf5ftUZfo6O2JqTKBHaCwFkBLB6tDBilUgjMWr
Uz5k3aUa4Hz89RfoHIwJMEeBonik2EMp79yD6bGL9a1SOOaVGuhBDiHu+2qsPoZPE/TFrvZr5cmx
miufnyJW40K7nGMlOYGSP0rWmbOKaZgDXlsi4UjogNOX7Aibnimk4bS3vBSsLUopEHRgwrANhjrP
B4nZrs2WNejpG01SkAFIYYf59rzwUY2i5qSScdZDUmh5kBk2IZ5dbADQnSWetovGrmnDaDpD1QRp
y9uMMOAcHJu4wcnlhPxzbk4t6d/Zio2kTZmEqF4gcNRyT/FXwdxwskfItjezY/FpR4hqYcg/BAfa
6/6UdcjhobcEM13YB2+XLgq6R0LyN2T4Ks+MwvFgoo70qKrdJNoWGFZq2JhTR/+1v8q5Sutl6jAn
+3BWZLKDCbS8M4PDf2fAQUJkFsn7VBbczmN9bAbwY/evkR39E4w1ePAUkUeV7qPU9ShUEX3FzKjb
xyX0BjDbZjcXmewFFs29WJvJBvkpdcfLf/rqLXOK0bDaYMa6t0HjfR4llr+/m36iAjg1dToagGnK
0iC6E8pjUMgQ7Z8zChFuk7z7gy7wq5Rgr815mqqNa8b/8Ga1NRoRm1S4X44Yspgke9luh8eAP7Zl
Inxb0dvD+5PTsUpPgccbNmUrZnivxd0YJ6hu6awlXueWj/YkhsWgplfr2KFXZ/xTXmAHSQQ1SsYW
EUXpjxXVMp4MpM8yLTQ9GpVQCaRMugppSvhjABS7WFH8PnWNsELXJRXivRdxgxvQMPxyofPW1md9
A5Hb/wH3tlVz/tmR6aZIZVKLPdGMFNZ+d771rr2PBSxy1bq8IDLOdjVzN6CfTtdZ1IYCDrTi+4Hf
uEg+uNEgzgxjfjM559gEuoJLsTm5FTAx9FcuvzncuvoSfpSIMS946h3PyOEJfymBbx8KmbvCwJbT
1+682ikbQ+WPS4hvScm+u3cjf9jSG88Oj6qAtb4T3UbuLR/UduRLUR6ntTFv0oUBTvnFQYYIB9om
E8m3SmjjWto5RiiihIxFFOfp7YTL/vMH0rKoo2anb7qDgZkNVi9Q2EQ3c1jcylSCnKezJS7ae4bM
0qExv2CTdhSUMAw8b1bN5bhU7ne0oOLLmXWHQoq5OGhRcKobBcqP1L7Lb3byt1LK5vKURH4QwBMa
LKdDR/p30CWaqNI1rdOxQA20nBAITYHSx1S1kVRUIh6CCUmkl6r8YQKkPPArvMdh5qFMGvOBu6X1
QMQBNMYIhdr0099PhgusXyKYPo7SCEQHRoM5lD71oM6RH3yk5GShjfbNhOSbej87DfkDO/U6ggYy
MgfwN1ZzN0+aOarQsWw2BQpicKa9PijL0UqdTQKAIV+0How6BM/b3nArtbWcNlmEM4XZKDThblgR
Q2t0bk9zKsSXK40/kBescK9Hy1iVDy8Q6Qw46iz4CnM/maJgSKIKCYc43PBgGkq/xEzV0LoBcYiR
XqtoregAzyAmerYs6hUCxborUJcjSr6j7B+CDlhRIc73yWKGfGyzNnWmGaQLbTSsvwliQXZjszYV
Gwp7psPIahKGOiDSR1HoRfBv7pqzU/rJMj/lTugH61sN9uZCvEqV3dyZJ7U85JuayCg2LmL41wDR
Jhy8AYlDKMQ2Dq7b3ZLaGKux0T1lQUGL13feoBfS4xQlOKkD3plgG/a1gn3EEgmR2tenqHxrzq3Q
Iywve+03JITbgBOuuoXs5vjol7dzx1p9PGUgtb1jMdEPiI/44//gkdk7CvTA3nrv7k0KtVEk/4p9
V7Blt8Pl2wlGJxWHUltpG0TZmTNs5a15/DzvkFVExJoW5OI4SY0aY1RTYJGtN6BPpbRLmLgd0CBP
rP60IL+NvuTCGdosJ9WPnL615v+jWtLTABQW++vOWHxfiKSnK5LZ5idi6VvQFsPlyjKS97dB3Hi2
obfniafMrwDPz0yDLW+fwOm+Ac+wKNh4taL5G+2c9oF2d7JvtpYt8YZs241fBsvz3mPvPcIBDTia
vOTQ4O56HrjxqGAgePPKsMzOBBEyfSdE1xC0/nlZ3dFnRlmifNXEKwL/FaxS/Hl7aPe5y2knEPF6
iaYRuTl9u7lcafHRuQyTeYQRxuD7Ik3YDashvI3MUvmz/RhLbxloBWpT6wAKVN7XSBNhqpEJuatO
1JLsNLtm2+hFFuA4c1D7ju75ZCYQW0UQopg9Nxr1v+bOXoSyI9PRR6BS1Wr/gnfwrDhTdsKBsBi0
RLb+kie2EpzEIgr4o2xlsSXheF8cLhCHRZFbo6A0py1nAMj7L4wPSsY+1iMZ6RDUFfk6/+97RnLE
RaJAAdcGF8B0TeyeWJkAv/alZE5w3jPqWuQWnS83yNPqGZOI9vX1myXnkUYbzQhJdB1Y8PDNZ5kg
+qxIsGSl/ptPtnxTvUMGHqo1MY49tqIaZcokkXtJ4jy3HKZyjb9vr+K6ks2SCNjKB0nSz9KWm8ZF
GK4CfjqbPFF4YlP0XDUl3mqMV5UDMIKTMcgWftGr4G0OB5WAJdN+74ktOPwH9SJfqNQzshq2OBh7
Bs3KjqdWrbWKGS7q46uRY8PuLUR4uEZNVnRp02N1KhqWA8jkVpmMlBrOhA+T+jtR/CerrhPPGI+y
qrEzqclIe2Js/pMebUPj7mfRr607+vKcDhZj700XQK55xJK4XYbXgFOFho/Uw5mKlc/zE3ONDwHJ
NBGh5SF0T1viMIPSiWh2CPMEvlEGgpb/lWmjf8m50SQhul9tws/nNOyA5gB0JsBKF+jNG2E+pb/d
Csm3g6PlzCYYx/uGpgt3RfObHygO5XYtiEcrGlTHyzUx1UUcY6gHZyXdbKWCW+e/kB2e2bJTdiez
C/pCdDZ/7fqN4+EG2sQBROYNhnlAxob4Vm+VWAFXDesoHdfwUGpsKVSFWLgyGJqqDstPsbgp+YKm
RrVfdDQWWFA4F0RnOKqvpfMJxWJMgtOZQ1WWa4GxWMv6ot0FVLy6b1l93+t02W576l7tp1nx77AD
P+DYJeGbxp2VFnBcWRHSAd2QJCM0PUFx+Y9veL2TmIQckOH1id4V7R14Dx+/HGd5ZKzhJJywbGUb
BjYl77rfo6AlqorNnergVwdXjlgpBXbNORb8oCNwvrsbbYv6YIkkiJgpuX3TIbdCHwYs6Uhjuy+F
xj6icHgVqFUZyZovbXgPeypxGoE4keqqKo8EWM1XmO1RLCp/F5YgE+xdBZ6PorvW2+IyC3E7bXyr
vLdl94zPwOG7jSDkKjVFGG52jWkdMhNfFzcCchsTzDtoWs/EqZECN1Axm0Yoh1H+KtPdwBhG+ztq
reixR9rsBp9QvGYcjFBlilrgRZRczNWVuzDrBTQRF3gFT697ac0FbM2rfOVOTGy9YWBQm8rPV0SJ
jrbG4HkIfiG+AW+PdfQdsXyG+Jhx4KDjyFv3mfo6F5uVEgwajuFPIxVS8J3HL91cEFgwIpMDyANm
HWpbjn5LaE084hK8cq0c6B5CJ6tKyNRuDrQtanZTys33tB1LjQdkp6vwWNYm7E2pUtW4Yxs2X1nu
FgIi6h6pS9ne7T0V8ft11lsuQ+WCIyROWFjKRP9eE1E5Ych85VtHCWsY5f4cLg6pq+eyVAjfTAf1
MkxP4EYsTqjoBYZyXD8yN6zN5DKXChB/xDFd7fWhbPb4sb439ZvPOoTJnqdjt0RYoIyRQ80gLgrI
72ykMSWl9vRNd1KRh8B+cwpznl937dmBKlCIKTozctnPlA4LVRw5AzmkTtjU22K8YgAtg4A+B5nZ
BKqR287ctrIFOA9Yz9hBxKb2V87TaabTZq13IS5+pEdcUHCcNP9rBPG3EOJNq8YJ7WK0cp6kalvb
BXP96lsbl/R6IawRjMe37wrwKAAxt9GoQSam5+za8o6pKimSrZbOrIyf+OGfGKIM4Vi8uuRCkduj
2MzUhhlJNli/DNAwvte4AJay9I+xJVEdkcWVnRc3oqqagJGBAw9YoMRPVEpZIRb2kMI4zcqX4ctM
mil79qcB2PqUyrzktF0LubZNej42OBq2y7ywLhHsQumdjvsvuLlYI4dGBk3A10toUItUxKdlr+y5
O6ScRuIzVofChMkObgpZa6K9vtvt6y6SNNdWeKU97G8CUpF0uey0yF+fsuFBAgwoO2CwfT9MiHlo
rFpE9L3Y9jIsFkR6KcYhaTGnVzjcD8a6i/G5NIWWPh8ti9Td/QGKM+aPU+H6c4uwxLsxAZqindsm
zpXHnV/xEHen8OW96bcDIlD6dgqkNOFB95IkSBvBT+pqklKb5gXYw/ujGhCENgG1NCuYZPe1V36l
Hhn5JG4gltRREDrjUic5vnZy4xRCqVqAhB/Dtnixrq9G+kIlViTVIhLHHVuaNR9boBEeb+63aS9U
+RFi5JXTgSxk5cGStWo791FRQ7t9ite0ntxUsFhlX4syFAAsOKHP2rICNZjGY4S9AlELGSk/R89Y
3N9EgYONwy5XqOR6udylyatak0670x8o0lrOQbxZ+h2VO+w64ZYF8DvUTYFuNGLG84zGI9bG4mea
/CFEyh9YbDR1ludfrMDscl7T+yG/ih8vnwj/PWhpE9gcPkKqrraVJublT4nazXmP37XBBidw7Baz
kao1PjZhlmUQgnhrTUoedfeu4q2Z3Wf8IFTZkiaSxHN4sPNkf8r9MFnbb7lIHlGlvB4KJazr9fSx
RawwPB0R3uRRw1qp2DWFvD+8nzBbNNhbO9D5RWvrH3fP7OZTFO1VCe2DZePRyw5jAtwnx6VeWZXW
NH7qIGMDmCSa5QSbQU/V2/N+S4M8FvwRPhbqP1eUPHCZjG1Wd0ej2+IphKixpiSxmR1qqUn6Z2c2
JxwkPslgopT9ysdsGdRNRHX0WBAJAdBtGj2vtdqLmE/00PplUXt04sT9C3dFqxXXSg6q0o+CyFE0
I557LKe9WdH62LlFziyVSxcDA3QvtI6Ik72OV8aRgSnPbIucuqC0Ibwbms74ZhwjsFaTBlaDk7SJ
bpgWQljqrTLhHf5NVuhG2p9O2ZbPJhGobLAgJDbjROU8SnMz9g2ANbsTSjmwTpD1upAeupORdnnf
fFy7C75IQFq1VZfApwsNuK1SK7S8JZ0t7W15Jghz9J3Yn0hRSMZgSJMnoEqcwPtmpuKFz04m5DGR
83PK2CCBX0cXdsedGV4h2C+UMiLB4L8IHG9Bs6VJZMgGv7Tr4mI5oSUGT6IcqlCy27XKBLjx3HXJ
7/BOWBZMVWdNx9OzN6PuYd7SStvz7RM4nCG9HtvyjBNqQDLt6DPBRtJ+vq54++amCK89jWzXOnxM
7ncq3rVOVwNW1hTp31yskcjTeNS2h743Awwzfu+qqmvIoqaAaoPS+JQhZLp+Kk10fltSHr4xyTdm
uL8gMUpKlvC5UtiwlO1DkqhjnF3uI9OwYmTKPdHa44awxd1l/QHk02xaorJWrKsWqzMaJcghWzXx
46DtSPHdvghXY+cDSFZSMnDfSltP+crJ5QH/VYKs0fKNHdRANwYtabyZTWVfZzITTU7nIj0fFLl8
E0K6E9wWgWe/C7+sLIm+Ac5JMzSacbfaPOpiA4ZWvLrI/Ahl8tL5kUh7V7WFWxBh8qHMTvo+ygZf
gp4IESEejAv1uFXTXWLs3Ro8QrkShW+eTY96Tuuqz50ok9Y31N7MIkz6YBHZ5bht5widWLb6ZHdK
ZX2tVCe+Q3lmZW6j4F55v1zv/iGq+AMUAQT8WNR1qfmztj7ZXMUUGvIZ99VPX/5KlXauoby/siMZ
SaRWmRWK6rOFjWUX85BGeR7ooz8hGtC+zJLilzKib3TDLTFcpk6B1mDMYp2M7dTh7zUNj+z3Tr9d
LhnFxM0jUrTmMpKsMH+zxQQweRGFM9IgqXJCcipogA8WcdLUEuxTvqriFS1Pe2AyGbgsrJOCWTd3
PuyFR+BfXxoGQL7u0ODOjRhH+8KOdZHg7dCOU3uHXtao2L4b/9HwF7vqS0o226TYyih1efgrfXjo
Lz63r1fcnuqguFtOH8qCkq9jfiGjBRsMrn5wAqHPeMcpdYVuQ4p38ArWTNCqhrRhBnHt4znRJGBk
W7SyWQnP/b8d8Y4k3cB86BHyyli+dCuobqEgBxbyIqypMdlX3y+360O5cH/8UHksPFsiZ7dMMo4L
fJpUbsaPr5dV9ah5xdBhwlG+uACwWpwLpfTgcKod+X328p/wFagPcwst7eGLixPi2LMcWuXgqq4Q
hKeO4jTK219ck0XCnPoQZW6cuq/aY75LPZzyUmGxfuKOz70fVNgfrybqSu1IS6WMxjsbYw/FSsO0
zyALAtX4V/gqqjT30TNPIx+LWGmDJHvkE/imUfAkO8xIDwZYf65iDY4WeFbz5tBu7feT5iYCjC03
hodRVT0isU9oFTufWROpgZID7wZ+tWnGVtcpOZljhzWdgo/TpNbH2tQiVNw2AkjxxQh1ibMiWGOz
0P3iqBBOLvRxeK26p105g4OZ3AjyvX6YySoA1hscNIH+VbinZw6mKAe7Y2L6OTJdE+IcfXtAmnMv
2Ze4AU6Pal6iw5xgpjZoYyzVwS+nfxN9a/T3zby955lu1aCOKU61eQXjm1oWUkg7hKbWgvNnmV8e
9nQ7X5zDFhFrL6Ghx6+AlwPrwZjdKXRAHLMwsqTEYQtPHQMDfZMxcFBAnQ9PYYUW3onB0nSqrhGk
tZwd04TSi6mjTDOg7s5jrPv1KXzBjjxpXVJYUDW5czOCIAcfz3A4Pa0knTY8qkireWn8/vPUiEw/
GPlkjrBqHvo/nrLUPh5H05+AsXF9d7QdEJl4OrFUIZHZdVEyZ93T1jY+BNTs1Lmm2WtQTFoYEey9
i07eW8t6nWDqrvviC1149qBaeYAZ+Ff5Rt7NX0zILf5NdxntgnkKP7EyPW5BZpLw+0daL7qnc1Fm
Az31f7zyFkpKbb7SrGgAjV6qJqDfYRoqfT4yXBZ7K1GgmyHpfJMWGcr1gEI4dewWyZhIhxR5n2Rl
UUdXQozKPoSPVTK3s/PGiAFtHC0/t4+1VPj6sA/xPR/OQndtU7gWyGDRq22yHoufHwJWzVWFhLe/
MEFx6n0vImOaSMP8BcIeJfUjEOyzYRHMT4hGryBMCZywaHvpwf7C5jit0HmOsCibel67dLn+eeDR
BI6PirK85Z9zizcbgTcDM6tdYMzIR0d/Fw2ejm4KfrWhFj9+sUORoJZDa9xaEN/8UPQONpXhvZO6
PpKrE9QdvIiPDwylC16HPZTl9SfV0JJk6cKiH9iiZTY+7WVzGX/kYz7Md3fKh2ZnGkqvqoTdd6PQ
9EtDWH1Ma0HgQTIKFVjWBxS7q7X+gtaRhuh461IHGcLzU7B0X+MtesvTEoR/XIrc9eX6CksEA35/
beK4dTT9c0MgFTcV63Rn0CgaqQKrkJjLldPMn613WLr22siAgohF6ObZ4oJ68Qn7ggfm+9Xo6Xf2
U0PDpsPnlILcfhpJN0T1nBEqVUAYxomDDzNi6yGLxhgvs1v2cvzBzfYAP5Aqsq9svW/Xq9y/PCSh
udkK4al9aIxx9TnMQWA9iZuA9tmtaD/QGaRnf77mwmazDNzVDo1XgxY8uIAwJHQ0zouzcixyMD7h
oduBiRh5TifogExneO1h0COKYQ7cMMWDE/h8OGwdfGX2BmbWxFj6bX3eSTZouSQDZkCYNV3MXeLM
F0OuMRQhz7UQz+aNhhf+6csUOp99qG65pgM+7sUUKPctlfYtrYfdNeyY/z015lHEJOHA/PMSPmag
TqTmI7bvbuWfY6ggnvd4YQZjdTBAthcrfmMB6eRA9+APHQhsESmZ6K6PkSSmDCDuAoInhMNfpD7M
fEwoQGYct9c1r+TMVH4SSl76TVgwguA+F19be7ur/sk2r2uCtT5we4LkF5MV2UP1MDZqFrHm3cZV
NjAxL6pMM8SSAoerbO6w+yg9/vY8pEceLGt0JoEixbotslYelH8RaDH5n77O9QTVxxlcLBmqB9J2
7eoxA5fuZ8bRyluJP5HRrdszsl2VCC1zBAn5pfiNX/CqDmFH8BjYf/zWorP+W895jkWH8qLSQuDf
2YCRod1FJ091f/JdMhNmcOLF5PrAhoMLidmi7GP+vF0pQFMEhj0kEZCmv/DIvQjXiHAzBsTYJMj3
C62IMZZft7XqqYrODKQ63oN9IIf2gnCIaDLwNBhr1olGRAu85hPLCcei8mx15Bcssfq9U6p+WAo1
Gu9HGy65nT5dHZ6NFMfTo6mXvOxP6uameNabjuf0fYi/8Y8pIYtCko0UkQQsMnGzNBy5cs+WABjm
PYInx7Un1h+nSZSATBwUeiXpZIkEQ2N61DPaUXop+0R3REmoMcyGpWO5Fg/o/CMJLmJBXlyfshm9
89gKm9sJ1xDxaChEan1hsTNpjdxSRPADNFXu0E4KNkOk8fZhcoT2mnv1k0HgQBChv8/DcAaCpT5W
RMfIFKt6TMNqWcEj9icTOnBTlE15JchR5E3aT8JZvuEWuA47X1+eTPXfapA8ZEFAQcklqsCMuS7n
tdEl9az63ImlvXsokMycF8IJ1qfRgVrmYiTZyNJm5yT2Tshn3db8gTbcEQhUUpxr7djnjsDYKqx0
3bhO34/ugLtUTx9ng7aAqAseO5U9Q59ZpA5kRUVhf4D1z6J6SoNEzztR172wTgSLntfcgfEvd4NV
gnFhlaWPU6yrZh9G1LK50V1hraHt9/vvq5UZPhVwzksQAs0hXvW5yzZ/Xt2HI9OJfcSxqbgUkkcZ
iZwlxqTLANXVn/yWN4FGut9z8yximaYGndiGrdHssr0E8ufTueUxh5FXLQ033kxEgr/xQ6dTkgpZ
AZjX0kByPZHsdgQeSuLBF+ZdWGdunouWKYBBRVnFMk3M+znaogLSkaImEc3Ub1DwybwEhsYsMwtR
1LZavhkDK4PDQoikMPi5e/aE42RdWshwTDAugAJ+M31gS9IIdMy6wLruN/oKHscmPRP55DpJW6LZ
+cmXod0GL52FY0K2azBkrzD9ii7SXshj6gzv7IMvAFx//SYLukWWTxYtzUNti+SwJluoVVUy8TYL
fxRj8Bzs9APsXPRKadEpJFHJ3qzUamkzbfxF8+xX1WGw9VHYxPaWNC6wF+Gvv1g1YTDz8qnBKdTD
TxcjR3W5QJc4BLKGxXr4rMO1uGD2ozVlJWRdk8VTEcuWHyCqd9N+hf09Sh6QpHoyAZ1NlBtEosJl
n2Y0iPYGIXOz/v6vGtDNSItiAnPza6nG3eAgx+i5HLXHefkO1AXjpK6HAvvaYaDcN3ODzbsPJw3M
lpoqyAnPICRELO7EoKr7EA0EJKwNtwrmz21fCNnMA8l2ylEVwkTN0g0w76IBrJT4doLWnS0UHgZ1
hxFg/LiO77pmzzOi1R27jD6BTxDUR9eDUeHXXBEe2udLgpIaLwj5V4/KW8q73p5DuHzja9pv30D1
Ou49stGvWUFHcBYLMFbjVe5Fe0VLGhXqpAtehjfVs8/375n8TI9lIN/xa+CMznpFnW71a6S7OzEK
DiW8bOPSaekucKvgEZqaBcByxy3fS4rFKiF48hvE4gX4ep/jnm3iE16J+o2U2oaVYAkmeV/dIw21
6fKeBIuuOrTDbBJ1whxEVnESkyg4ISVHPvWH0qOMXUPyThrVXdOy3W6Z7VnwF+Jj5IBHLqW1CPbY
/d/p5RysdazAHfycBeXNucOw/aWFqIAiWCiMokGmxX/FO8/RdjW32OAphJtntcLxbvVGwdG2W51l
SvdC+yXWHQtaMtCqQKCI5sc9x52y6PHb7osVLosboNyBX+xuMDsTZm78LOl/4I5UrZFghBm+tqrG
tEzSriOndhOspwZ7WwAwqLfrfYYh9ycXGIq7ENq5TpOWI+chU/KCOoVpPTuccdez4lu9xCRPyFbq
I2Ajn6o8/7gMgZ/HpYv0kDoCZZiMPS5ITlhyHpMFbwvrWYzR6fHljpPrE55beZV5h1sC0XhA1ykB
L9h1e0qmlQ2OzMQGsOT5X3XYn65rfX85iG0NyUNQ0wNDslPHbAVt2C/KovINgKEK5366gASBXCOn
3DqwujCFmTFuE1d6bX25+lic5pm9/IVYNw3Ne9BxQm/Oa3OvtjJrGpV8fOpfNQSLC+zJCQ+udrgK
AkFbEgiDIbgMm3hFabb8H8oGFgpObG1yJ5NSr2tWbDb1B41ogvKJpwg9Mhdv5KoQbFJMKOymPIPl
VQyOLqeaUr38yZNBv64Llv6gx91y4S5XjrcXg09acVG/CH/M61qBiocKSRS465aNFIbeglgz9eXk
tEUj8jISEvWEIshTYecdUaaDHOAEDVdW04ucEZHZSHBWfwmQKFnYodSZICo7CRHiZeQjMdgNRMiz
r4lupJSqF2ppS05gRyvhrvrLuQ1ayJ7zNu5J5L5enualz4pGSNc+D4OblWIcbIFxN1Whd2VwNV48
gRVbaqU5FcVqYmNVzF5qAP3Hy85IEYaIjWzgXCsyBmHq4EkH/OTnMaUhBjeiEK/Dt4W0hDIt+L7b
wjZc62tz9eS+p2RrhVpaXv/oeqsGZJm/KpxZSntMhUp3UmYuzw7FNZ8lIGgAKOq+zLK9sIm29JbF
fzot8DCqfjQ2dhsHCrxIK0uy2qFIc7jaAs51n/TUmssD8u9ZoG9Na71ONJpgr3vVSynlJ2mfp9oS
FuGhJVl0B9cHwgOWFOjfzK2DaYfFhalqIa6EQs9zQb+O8ir0oLLJFBiXjNOv7xq9+3G0SaFCQULR
D0Kb0V1tABBqD3FmfntBt+q30hLp6gj9WyIEjnUv5DLkycc42nmkQNTd26sB+5Arv2z70GI8k5ts
I+SstiwZ3wpFW8wjRwDFchzd9yA6lyhflt0SCGePvt8BYH9X+KrxAMxA/QkNEl5Qnj5x3cw4Tuxg
5bM78uwBXOoVf/mQtvHmBUXYmY6o2/fL+UFvq1iuK/2sa1CyHZBcdr1pj/4AymariLlQTeYtoolc
Qs5bg8NdSNuZlG/CSQzf/Lq1IO9ORYHtIvze3tMpQPXUDEwp0J2qeRDEWYw9fZ/RWBDM6Hf/0NW9
GMsCj1OR9j88kCj3H9svzfLmv9ZQKFLZ+YFHGykKufRtOg13c55kFcmYX5eTJ1Vbas1WmtYyE49S
BJq+0KMNRjdtvqk/BSkWE8pdPGDAzNtZojz+E019RErazacydCRRr5LB7MqnAs9ss92GXp/tXRYf
Dg1jxxxVwLTR9k3/lnjI8UGJosuOoW31BH8yDFXZW6jLifGDgH0ZevcqZOIACAwypyEyKATbUtNg
ROyotWaVALMsP2gb0mnoEZ3ipH2qs48MXRQ0geFEwFFUXG7AbOGxYmFxXCPzIOblB8xXR4AC/xFJ
f9R9ZF5PEAMT1cxYyZ/UJR85WhXEbkvyo2FKD6b4chvnEPUiInNx/S7+/YHnzsznmsbuolQ7U6z5
eQUpt2NZ5eiPDQtjFFKdOBuddHeV2En4dl8t9AyqleTeKQVVs+/7zrvHESCAjCEM2ZEoHAgcIRdA
3rqr0PrGkw9mUX/xhrg44M6/ghD4BuDwFvdOYBlrf57LdocspdBtgcrIdxivv2rrwxJpRDY5ulg+
Kj5GtgJWfrOgQu4pwbXYLdy7z3oYXSb6s0ejZg/KDczcLe/O/iXrqxdfkKjx86n6jRQgrKj3Lnxk
cmuW0+oIk6Ags2T/XwLVECZUTpzd6RxBhlJTtxGyZmxywxw+sW3UFG6WpUDHn7rRtd76jkQsXTpp
bN0wlvqzdzrWBJrdbGg9eVL8qgDG+4KjRVr2vc43iE1JrnSlG93Os/XnmDNz2Q+oTzG12jwYtIC/
/wqfbRNHtTco61ivvrUrV2I2OhB62m9ptfWRIMVVvlmnNdKExw/ihZGtugUSclSk1L8NJ3iNlYbU
QaLUwNyizskREIuD83E0oTXntlsLl3erAO00/cvF4Sc83iwGmAC343kK566aj1/Ylgu3s1pU2aC9
ihlimxd1eJ6xpRxc+HBQF2+o+Gh3STI+yChwxaAJ4UBkffg07sr77Od64f/ODsHQ7eMFg5r9vk0y
ou2wt24NmCAnx/3lMHU6XX0eKyjuVYUYYGP+MNnX7j8t+P/OYaX9i3vlD3zLkHuPjbEQe94eEEn+
AbJTnH3twG6p843Sp2C44Fhm65EwmqD3uBG6CJ3BJY054+vtQEHoewkuC3E/VjzmO1zBBzpgOsXH
wjfuHleB8bh7hvXGkUmoPJCl5FAUa9G9WoBf/gmfX3R4004aw8Dax62L05wBiv9eX6zdTbPgmlos
CRK15wUutHRKEInmC9CwZYYrFF2TSmggX8x/D/fa+c4GzjjZCF+8G4UisWDTYoWe0RMoD8dgYLTM
kCGsq9L1T3c61AmAdoxH5bPZLKElPP8lyBNDDkS+VqKRCZbFvNpaQHFPsIl/33x2RDF0DOA6y/PA
PeosG1Da1C6QWaERiHIXf8SL0Tbbfutk1qZqvHYFdjbAb3OjoV6mRUva3OEPypGRd9m8oW7uNSlV
/+wCauekOF143HszH5W/hgxxSb3RUnQMmgS0Vml+ZTZYFaVaMijqLJwgV7AuFB5J43MF1+bUSTIO
mnOVuF9UHwgOCzd7eWadcEhDOUtA2Yl/atMUDUlpOOeXgrYgS9Lo9PQMCxk+ON45FBT2Sy7vBt8O
KDi9akUpTETU9+QvCKqimYCUJEbICA9FGzwGR65m+J+NssQwoMa+JcAM2Dnh3bQT3KhBLtJZk0kg
AepscBbTiVi6LlAVJoqNt32BdMZbU8nItCvIShDbkOhfvVHmnkocAtUliGllCQfftb8PhjQXgEPF
AhHPgFuAVGwSy//ciwZSyqZqOje0WCrWKkGHSaaUaxnGRhLRGwQh1GCZtT9wqFOAIxveQ2gjdFDW
RTcY8dTjOd3qWtgZIkv5nZlGF+WjVSXdJ3ZvPCiun2OyMMkTrsbWvTX5PeLTBBhUQSUMaxjvAGxt
xnqdDf2tVUsrBVtsj2H4F7Dr/Fe/fNKC4jXhzv8T0S7m4SiDctpsIznUaeANjhf0mH9okyQyljdL
tCFDjirdjpCO2M0py7hnHNmiimW4KCLfzJ4RZ2b+HH3sPG2F/7+j+xvHmXEWpqrrzQ3MlvCam+IW
fKO55HLJCNN0zNY7kAXZ7rMM3CBxcHee2X6UDgTYLVDhDRMQz5Br6NBU1hUFp4vPpDNoEzWMrOdB
1AJcVxoP6ZqZTk5+TPX2TtsOo2HejT7D5y/6p9W1s1x9Ae40n9kMaZx2yLfQk74uCBInJ+r0MO5M
If2ypxKxdinJTZLhC7YRcKX5kIsg008PFKfsg8yvp0R2X1AKG4qyQtSQK46AvgJDeEhBB2cElm0Z
bPB562bMmmjE0kYlgz7zsoQFFDqHAVvlxLjNyYNg2Zbamz9TiK6qSvAcPD6A3ddoz3coCbC5Th1v
Uyp2KqwGAOlRTgvOR+mfYTV8mHxYwonxPtCuyAYXnS+PCSMl3oqV9Ulic2T1QnikctjjTlPvU7SE
P52T4x+2D+WKcrJo5jKyK7T7I92Ui5LPyYd3ge9MFSG+vE0/QjsXZ5PbfU9ZywfbYtteHfHi6PDf
b/rvt92BC+fJqRZMCE/qlriK1bePdj0mP/t6Mw00sBt2BlsPdOr2HYcZrdvPZT467NWhmTWybxe/
oaSbPjoUXf5Nkl0PDqT/XTQiQKO6POaKDOkBB2kYpX5eXpjA5vVROSW+qZPGJEi2qH9aV5gfMYyC
kgawWGkMyhUR8YUUmPXuADlYfH8eSNvAdeCFP5f9QqVr/V9GGx5y/IwA/YIQoA4ilqpQUpoyLlrm
EVmJsyT4xXx7zMmUv/g3iTPj73VwMog7c/BcOaBS8C9Gg8dhkbW6yMIg8/K3dDgboWWnN9eya2Eq
aikctZDMzKDKsYNCt5ksPw6IL/dOeKmWLLYAUlckhsnIsytA8WOFslNNZIuffxQu6ejgxTL8l741
v+Jfp5bTDnIVnB98o4GDuB7kvSZDEzbIp9BwsTZnuD04+DjiQr0pXnvD3unxxsPWfAQna7H7go1v
xkVSW6nq53jSccAM2kmBRnL5VNkmhUGoklEx0mBHJjB4fPBUK7SjepFf5KISHgfRoq0sy2v9Cyt2
0iVz6FYFhG3XRrjkHD/xDYLCv8QBcrJlzNxtirQiLcJFnyZYCroI214Y23XJ4U5iabyzOj8KJiZM
eNrrgl3vbOiSvgIcegwsDv9WjupNGDhtdCO5QERFjDQSqRNVEF8Un96DENpYe2oATqPygsQZVQtz
wQfNCY5zDjdlx6xLk92KTKlWL0zyofFNFpskKZ3j462wNIgM9/lZEIO1szQS3U0UcjfxHLprmaan
AMa3ANQJcAOynAT2nF74WC2ky1n96Io8OYOrrsrNcjjb+ujYRLAhrdlh5rIuR00Vv4oLOkN7uo0z
+jvxm8iM5wngv1Uqu8qLvqAtoT7fldO0eUvqVL6IsvToewSAA2+3lPmoR8uVhRip+DkFWMy6Dyaw
L6gB6gZfmhMICDlYii6BZ3olZB0LFaDrxFf9iPPO8DgbQpqILUEk/+1EiYk7OsIgQqN6hdBxV6mg
GYf68K86C+TaZ9OgWWjOnKcd5B+xIh0uhRQviP3ZXb+kbA/0smv01qr1sKMiKqPUD9np1h2f0tdv
SDMvwfzIvu1cxF1yE6dGs7wSQPrVpB7xHzmIbug7zqiDTYGSj+KwBBxYWy2rubbriQ3lh7NLsJQr
TOoilFjplKZ6TVvtCxQas4vArsd3/7RPC95FvKR9B7Z4CsIdFpiWoB0LcVVw0Iv3wy3HPukNl14D
dy82Ih2E5w7DkPAvl1BFGp9pspUCvYaMZzrOhNTezyU3PcnjfxUTs4ZlTNDzO5O40nziWt3BT4PH
gRTFTfMYd/ucNPK7v5nRT3nFzAPQa1Bswq3ulOwiCRHdKZyZjuiYUImWV4N8J1W1yEhXUlG7do4r
MalJ6+SlUG8nMuhVSWGmUtbJUCvNfPJekCw8BbP1H9wnJ+re6UR7rs7tCyXcirZdaDs9NMjIEMbw
8ShZ4EJ5DEZ6SiZK8Sx1kMYYxMKTNhSCSzehzoA2EuWC9rdvTZJV98yXomVRy7zg4BZlaRyaoAuw
A6H8VzFHycNIPQ3lwdu6oTNoeZOY/cefzb0u4gxfSL1YGwFKdtcgGeM/Jk1VTkuewC3VEJIfOdIQ
rTIjrFjVXfhbj+NwzhDggYkRLmN+u5+yjyP8DR1JhiV93M5QIOZHI8jThFraLG60bDb16SIjdbW4
ZpVAxDsD4IJUjSXJU5Ml2Xh1vjCSETU3jYFRmN/4LDiWt5b+cW/iFfjid4Z+tBaiQZgndJxoTdMC
3qsfJQLTxr7oi4jc7p0+u/PofPTCcYwixG5jigF5MUqWzTEl52C6bEv21jIzbk66BPj7oUiAhAOq
iO2VxF46+Z09tEec0thezmVpw9J/HtLbryngAzxN7dXRSpGKRAOYd3WGaLVH0ijir176j0q+1hb1
BdevH6bafk13Wm8f/EJnLsrI+dc058CkgzlBr9VdVLwGwELGNotcM9heoYtv2ooHHXCLFM9C7a1J
SufPIAQadYLLMNVmK+tY2v9wnVvyKXfqspVdrhXoXi819X6ANi7bAsvQwOyjuDWUva2qsEasgrJM
y0K5BeyQXVD8w2Ekh5rFkTICrYHVZ4HIHHDW3H8SXC+o6XNZrIkdAFTJv+ihFEV/jxhA0MrRhzgb
tRP0P2WX+PHSINzrcTsptx6/0svpjsJKjhshkCZ2kGW9D9JbW2D2Bwd7uoB+1dQfDMLUqIWWL/Fu
De7mIsgrHrjlArTeYcqq5EnG/ZzxggLUOEnTk1HWK8R6ZSmUbU9uj/17i/XcpPmcEmgMRtQIX9m3
OpuQXEOvNccKCbGILoVsxGEshbn7QsRBpHnJ6tIE2p7B+w7IxzeQPmcv66qpel39pyeL1FaXukwL
FdNVosS3ZPDtmpuMeMApgF7WoJzlFCB2rPV2yJwDf4tP/BnGF/vCzDenWimLNawDw8M9H9r3535z
IEeQ0ukaaORDJB7MZfVCpiVxT8KjvhVKsrBCBLVx/TtI9Bk8hZNekCpMJzin70ERpNkrwRpJh6hC
9YefWRMCWiT3H5ZDeV1SoV8p6p4NTieY8v7NMkSLom7DMMDTXthVNwZlyj1iwNy0k/0RkEZpCAYg
7nySHHBaVoFaIn1nh+R/eHdv73kgOn6dUuqT4S5w43FMCZqauZLUAAyj2XxFaSZNmFkUHk9hJ/2E
Q+AwRMqkAgOfmLTShQO3Ex4ojDAMCNGf3fGrQunVL7h4JA9cj7PU61Bqa/oiJ8t0bk3J0JrJWRzt
YY/mYGk+sWImIe6umNBxuw8EsJeE1mvALitia1XyFKpjJoL5bJgdrTswZ2wPqeRVM1GXnJ+dGqtM
9XGqrn9BXgNNLK9qCRR7M4s15Q0JjTfiO2yX9io9eT065qvbnO5E7nEIuRfUzDMo4wBMM5q8HcUM
Yqb9kBX4HMvEiakE+pmIbBbLFnSaivw5nrrZTvX3NI9XdFt2uwhMaq+opH5+aBD81MkWFh2YcusD
4KwgsE6gf51ReYv+eurSFFA+229hniZBQJb4car1lD9xuJkdSKjOeOiYyHIeSMqRJNapM5sGlJ0M
cyzY6GguSdDBydRQVV3UPme0ENRuy0iZl83Wa97rKWSAitabiqTcbdtYw/AqPeKTK6E3gU8QOIT+
OYJxx4w2vRQEal8Fb0GZSumvX2lcRT9/ASGEXAdIDe7vf27it1OfOslx8P1kbghBujlPiMb45/zN
iaNkn8Ltjplhg+braaez3EpEALkmmTK0IzQ/K36w1UHebLftHH47Qbnl8DrzN7y7xF6Yxa6FvwVK
0urRSAsciDFPwosWAINwAwdQ7Ea1H7UGyDlGOI2r5fWK7F/62oBjk2kqMKBdmZ9p/CYJPNdouEB9
KTVtSr23n0I1y9tqa5dKXBjp20Nq5J9IfRREf0J885EoAZG3X8NtoNwKN8/SD+MqW8aMx7xBtQxO
8YzbcPMKIQDmUS7oxjw36lwwePJJ51hcUDTmAkca6dGXMKUDs2UqUXWoUrcYHSvxrwVLGd0Y7qo0
bX2x5w5SZBo/zp+CEu6hck6DJerSGM1gtXlYVyNv/AmOyqvNJ0jJn1W4biFxlztpAShAzHjUJNRa
QmlvZfoXg8EKPYvQcWLNMxXFsUgGPKl4hkobHh0dOyeaWbjN7wCGjWXRXoRDIxrWALlAypuCTOyA
BsR2mLRE1fULHgqWzBA/ixCC2sYG75stc7NcVGIMR2TekZ5f6Px1DoMePMleVw7xLXhxifTDCHj4
cCR+IRymHov2BPhz7GP1Jh/wVOWyB9rC7+5KKPXg7h6PFPfpp8m4teKwcj25a46byiFopJpUH/bT
2HwkDDL2WEA2klzQbNOD0p5Vj8YsScLGLz0rwZhhl4/qUwA1SO8XZjZ2MBlyEoa/x6utiZWCPmSz
+ExnlU2edSJugxvJ4Sb81hTCfJWbAvnVWL9nGmKvllBjXhjdpLcaekPjjG7rx6vp/dj9NYnM07eA
C/E0uuH26GUOcaSLRfHla5HdzmNrkeCY1sv+pgJSnJyAIRwQTCJNyzvrzyT3H2zC6+CO9rL8UcHU
MLBSFWdBc9pdT5pg2tQMZAKfA4f9Rd+kiVWhHdkoXFSNvC8qADCokODLlkOHBLEubH4vbhGEz4tR
CItExf5KcqBMLzY3ubWYdTq8iLPnhU5rji1IEhACUd2sXt43h3CwUgoS+g96krYNQ0NFFLSDfr+s
w5t59cHwDzF9BVcQUDaQ069GH8wmA2CChwr3F9H022jMHCQDbemx7j3OfndZxgwMq770L7GIWEQV
6TTjXZsqHT0f3PVlMJo8LVdfX4fqclQJPan5q4Rd0ncFzupxegVlY7+ZLK7YFPbn4T4pFmrq0Mie
oyxX8GOHgahH43DZ7RhwEmHWrNfUboDURoTA52PD7xk8h60B70GpB6MgwIn67L9Gqbuc9JoaRcEN
jQlE7SxLbZmUHlIpU9HOMKVLdYGBtURxS6NeakSs4+2DsAMJZkRgyuDCFGZTA5jwHegTKeNZqNJZ
FoUMSzYuenlQW7EAJ1PbqNq1CRQ/JPFlgt49aBnnSjpw+GCQFyTyeBlGuUvEti13CwMbjmX5iUnS
Opmm0lAHtr0XNQiJB34XhLc36X9Y8Fct9lSiC2Qr86yWvtRCKavuY/TwO993O04S2v3eQQOA2qiv
QJI8t83q4rprrNMezAE9cpLuz67NiK+lgT6sChL/kyTztFKGyUA6Ih9WwG9n7dpfIJfx2OMm16qJ
ZlqrCkWhn60saqiz0M7yCC1LYip9f2qAyLJaqSDekq3cjXtpeNTP6QYRiN5A2BWW0CpuG2gkXAJe
k/gnwnQjjOws3Kdmh2S98gzpg+fp8vFlZTASlyGDA5BOB15KDvZuLgtuN+nMAa7RHTzP7Zj5oKAJ
T95ylMqszyqb8HM5ji7ycvy7x8Cs28f3qTg0k2BhtabFDlm46B5yJe+kBAeEvCWU2iberGqXFfZJ
I56h/okaxRZGVrrPJzNr4nM5hFjdXrJvBQEI0iMVwraSDqFnuF1kmRM/pnXcNwAZEf7+glQyzH6j
BzC+QcrKPaPpubPRL0RtrLs/k00rIaBPnumWWMBUL21m5lSjkDknIUGxuD2wc6O2hcMdf9DBcPGT
1P+k2Aw53J14szF6+PSYil1ZDoLdMRwqZNEQj0xebuV3cSz2eMF41RP/uaQedzsQys7/l4wftoLA
EHBKHsCiNRHS89a6jJMr2hh0FPhQp35rDF2J6Tn+gCCw5Infksy07tx4B9LbG1SfUYRuqbVqktP2
Q8squUeU0gyXxARD8+1WLTCHaVbOFz+Nr9/SMPEOHA2FSrkc5gD9BRLT8mOC+39bTx4T13MhL48w
1HTvDmPPrFa3dVCc6kCLnJ2U9yslCuK0RxWP2/W5M2bJUykwojTJyjLgk1JsX61bUeAu61oAUdZa
d2ueS96sDYtH6rDIHzMHCPW4E71u2v5NUPZFwFnd/MFbjNr6095weHkaaRDkVHRM925ZpAd27mOc
iW9+tKHyYiyD5KpWK854d4sNHkiHfaVrYNgn4b2aSDNNXP22R2IQ4K7rlos6eW+gREDJ3ACA+rYZ
jg9lm/Fw/GV9RWVIDG2lnxBEGTAAs9hk8400hnJoRtU7WjKm94rfb47sIeGEYU85tUaxapK40nbh
JyJJ8CpfUztbJ2c0wi9n+JwL0x/kwbqZy1XW8C5UyTBFyfD2xx85PwxJaWdjPj3tMIWAD9XNeRWY
KKFR66BsfbFO0i/OhUEvA4pPjK+8c5/BC/ibUFDfQii33jUPVCfaVMlCbTY1P5wPmsfNNYLsek4L
IODcCCTcNSbUbXA07GyTNLWQMB8Jns6+jaiFdDmrEo1Z673xEE0mBkZBPcJhQ/xF7+32OhyOOp4b
525dLm+SQVso0dAQDgltyth6ZHs/lxu9WZzpDFQPxIJkGyhMxJUPybgz4sF/2zVAWp8Q+A5g9BIV
NdY3WV6M0vl8rOHL+DjWHdvpo20vChUjgXujdWtcYo+Z1sJnEWK2b4gu19f0R1xVyBQk0YBGAHVy
U1FAzEBIDy5Nbi7LXQt99HGE4PWCiZPbFIsHv9+SqtKsoCWAvnlSEHifX6930UEMXRG2hiXZnBZP
VP1qDJdSAFpWXEMoh+DdKCRKHqM+3VXUkkCZsQPsRX64RfeCjyq4ANuaVCsuBHD2KUmfF+GGsE7y
dn53IwkQ2fxvrfAlVj5FaqvZdeCwgQB27w8Ub6lh3LND8lZmQaoD5gSCcCqeEIFnTh47rvR/qNqK
WOs9GiaBhoZnDbN9qHgkEqFKQFsntEd7iqBOdhNwHOAKNoup4oxzgrjBNoVN6ve+Sw6F7RV5M+5J
qOt+Yej4IIzhk990x/uMeCqsQHAZWfHeWVZtfweVvAfn2Iz59Pg/5WnuuwI5C1GGhbtB1xDQh8LT
zPEOkgSSnutHzFL/XUNQaRyuSpkeo8OuDvjRWyWGgSjo/TfecxxCISSaazaDCiyVKSlwY9PKyhUP
KPTZq/VQnpqV7cGBu/o1JkQxqPNd+R82X1vurSBvMb4Xpz/LLFmKdko9JHWPvlcbFVPq1SU+e0vG
vsNn9vT+abQgcmHXI4TNANLs2+0AAvz4VLifP7LrvCvRhF4PO1wmdPS80JMD4VDFCBXHrn86KI4M
WZ6h4BFFXo2LEon5794R9kAkPTq4DqxMZeCZXI2byVKNbQt0cGuNH8j0fbcZR7UnKRlJ0p2wkka+
wpyS9snQ8j7T/F9D3ZsCnBi6snG5EEM2c1Wz+1EolIkziaJ59j8Szj/mV+Zb2frHMvZGDen4bncY
fwH7PhPzNkKJQ2X3cSrwIdInKWKnF7kGMtgX6q1eM6QH5t/9R8VQn0yoyxpYZfbqvn9EvvwFlZcf
CB5HryRysovK/QkL7+b9Cpnc8ZQ9t0ed1pdk0EwDbegb3kKEv2ZbHANwScTHP0GIC5o5E5cV5zaQ
EK/w/BUpUmd0wDSiPB/IYGCbHcACupgmdaLheVlsiX5LZxldRxuaCRFYOPtrptyS2zsKA54qkLJC
xz4PWqX/vcIjUxniUoX0PGBKk88lOoMkSrRbYGblXjxzRn/FqmhIO60eE6TpmmJqQBsp7WcRLt2f
kRmThGeiodtlbW75SyYnI+4jQWTaOWLwlC7pS1NRqf0Q11UVmzknNJfo/Sk6KsV2ByHuEr0w43Yk
dCMpIUxPAeygoJxPF8ZrV60eEA+f2ePgpjyY3PI2FK53B/1TsQVBo0eeoXBTS5NmPIhi4eoMB9u5
50jS38bXtU/NWzo4MMenVe+7JUzbmyPBRrn7YcOtOa87mmhUGXaWu/rj8VQGVzJZhBr9KFZwpxFL
q42yZ+5aIVjJ2OuwgFl4tjGgHcOdnZRW7XWeIlUPYmjSwcuc++ombDA+FygNbJWJxuvZHH8dAaZC
srGgUf/U/vvPliyKGXvww9Qrv1Dn6jgOeh4//1N3gR1kNWAtjhdFP4dynqtvRHrnCIqfppPqX8Jz
CrifkADhvv2hz3m0VbQLm4UkHTcXuKwnhFcrYgNOTC5/3Xkw8HNWYE2ic+yLAfFZQzIODJioLUwU
4u3dJZWXijGVw3ovrzeBttL3O5V61ga7jGqNI4916aGU0Zoyp641Mxmuvo0MiVeh5L8yEZPkqc6S
L4qGBnHOSnmsIQvK4cvLGxvFIxhLI5SnIqVNyvsKSc6ZqQWHJyyXErJpKswDpe4Mbd6LUkWZn0K9
jfbzFFpAx5FWXd9nQWUnEVPX1qSF7TAigrMyZrWQep5SjRx1YnLBpoqMK+Fcppqd3QMvWXBD6T+U
tEDPkCdUas78NLDBEAbOyiNktYpUCYty23WFOy4Ge+RYssZRYIFER6JmwBR629O0OrByhlCwedbM
TCPHrw4tQSt+sr2kQhGybLB01b2+9+pBIb/GGbmxVHEeem2Wmp6z2O03ubk1OTiI61vJ8R2XtWEN
Zf4Ii7w62qFfbK+DQrfjJjfgz9qPpQ2LmnaxAf8JNKA7JxBmJO2/wDq6wC+rDN29DQ5Hd2Fx7N6P
E32NAR3zSAG1vcA4kGeMEpnGxI6hAPH5qokp+yADV2EY3A5HQN36dVQBpW+wSSDofNMUvtKxc67L
RPZBuyMqEN6buViZ/TeJjUukHr5VCsSX7kXr8GiWrnSYREKAW/Xje57qnuzZeWO04fRhIuqvpRtl
LrhPVKCWC8+UahWDcySue2NLdgDIE3jT8cNo7/sRi5B2zrAp5EbCVW1GEucZL+4L+Gz2WonS3B6C
Wc/Bd6PL+wYOy7jBiNA+TUOUmf6LPsG7h+gvhe/JJFst+RPfZspfp3+LWAgB7m7xrQy2eW9X+Ze1
Q0nZwLj/eXN34hVpEQNzNgK0fOkPz5Waiey5FwjIRJwk9di4gfejbaIRjyNRMFObp2gvCNV7cjeA
xYyR4EnOxT5zJQQma7tur+iYnw6AsPg+i7tH0zM798CIWwD7VLkFVF+vb1/8U39V5hkxncds9clJ
RZ0ZRSMm8xceofzpOXwtMeWMFmhN8D3BaGjQz30l9SfsCqNJGxD9ksTiv2M8s3PsqQFKo4BfW9mW
p186jvfxbtiNgEtMsXUE10D+dLi86dct3UgUoTmD+GCoK28DNe0Fxg0ZnEeb4sJOQO2QnLYeuxhY
BLD0zes4XDZ28ZlyJqCH4UenmxdVJGusst0SCCaekE6zb6EDkEGN+jAi/NUdWTx9i8hx4fOgHWJ6
Y1SL8QAFg0rDxS5bicyjZ/zf/FdHjVY8VLfsqnAjxO28x6nhlkY6P3tNHqLXdvJuku4ucXJHuznV
gC2KZD/Z8mvDPUFKtPwru3iUG0A3RlXk34lH2PNQ3V7YwyUqJ1sLg7CkBszobGs6r0EsjBMzfuSn
bufzxTaXhmLTmAyiO3k16rU/LDSs1kPYv7RtE1PVU1JQBPgzDmS4Gp1OhuSYYGaWQTWQUvo6rxLe
4zDY5rOk4D1CHcHfpwSIvB/1j0CYp4QhT4ujSCt13wN5fe6P6OeIJwbO5opbUDnIVv3etjEGeSY1
xQ0ZqCCGNMhD8K5sZbMzzW9MimtUPzSEcLZsWN7jUpSLSa83jIrHc/zlNP8WpKL75ncnXJidyWd1
rnb50BfqOVP4yGwpmOj4PWTRMSv/Puz6z0s7FOJS0kUDHA3ttcgMB51Bt3qjx0rqNDz2qQx7PoSq
ZfIsGqGuga0QtkvIWnCX6xVxaWatAT+fPpb6lJxN+0QeDz27kGAJxm+esSbCHAts3wJWV5VHwe8T
k8KIL4QaBkxp82B24FzvIgDuuunuk+SqtORF267KfnsS7ES/zY+MFI74qu2NlzXpOxzAPb8+bSMz
Tn/C/9wIKRlwxFVaN4T2KzntxR1KlQT8UhPCgokQSZxLXtn9GdF+d5uWz0PGL1mBRUq7Q6w2u1AQ
Fm3L7hFXFW+oNh5iZdUueuws/hfg+vLQZ2zYjN11kwMYe0zQ7mkBcu4BgV+Mrh578eFZD6KTBjrK
mTBnG4MfouHRMrrJBmnNc6KbO69WvLq/x8J/opLuO2yUFzCfLh99eJ/UuQ3X9M9PyZCQW7CLctzy
E1M17UjphiM8JnkiSOTO5j7UXpQFswDtIg7XMmn8fdlQutZPyCXYVETuvm/JZzBhji5zFgT22Vg/
1NFiyWwKd7pJrEf1kpdahSXAZcXkINR52Bgqbdiv4HVGkRhc9+hAMCNbpPjjaZEAzAI2sOlIA1io
5DGrdXcUQpR/BvYu7iCaaZJqHbATUWg0wkMJPwkvRYMBEqWB3boHdmf6bx6/Seb7iNZbETlwCkdm
3CZnGj8/GPJxQb0R7WpsPeFOOchGhpY/sz+9RF4tMAnnlGJJQN4xezIUMBLMBzG8ygemdU1w1ypR
AUKoQtdRcmMXGvjAQgeivSE0sYir29TxL/nprI477bt+Wha+aTUrckAmX0vL8iE9YlIsEb988iJP
Roz4VZWLGR2AsThxziwv/209LPHu9LA8CiWhaKuwUM3LJLzMOTRho71o3cJPzJF+KPHdWtqkhR56
ky2rx2v6XH2XGUZRyb3wp0iDY/pUEC93uVdpskEMJKhdrJenmu+7C/+qKIC4CHfUyZxVT/+dYM1A
n6jeYWccv31H6gP83BZuqcVZoslDRExkYoqYnVP6TD6FZqIZVOtNJMw0d56CFriwYioSrP1uwJxF
pQEojrubtKZhiItBVfR7v6NB0Ywz86UirIgABR7NuAuMD9kliqilGaQjZJoawFkcTS2d7OsvsNrA
YrxBF3A+Zd646ZXl2xLuC/56ENUPrOB8s3HfSP08mMgcZgzU8Y9Ji1sChmLgtS3uDO0b7eQWypQZ
SD3ap96GRuyhI46p8c99vi8JTFotpqjc/tcpspVPnGqNeFt5xS5WpXnuRT5hP5inHXwsxtCDLpuL
bBwNMHBCxcTTlGumLfMrlOZA7rl3Qyg24b0s5JZ/IYGuDlBRmzrvi0OFLvAPTv9WO2sXE/UySPMP
o/Muf5mXA76EJ42ZFYgJRAyH8ylVsQus3htQRxYdEY1fqScm87Ayf50pKf1aWwIsvHSh9UzkAgyJ
H2rW93EeFYgIb4Cf9PmvkALF3xaEpncBPi1TtgDJem0QDndpP2PiRhUGvvSkyr6K4DMdd7zxiZ/K
qNXO648opXMnvOPm3huzhkBco+Pzxi93zsXHzRVE1xPzaa/N4eWmp6sB6ziOw+r1yuJZSMEAVmlq
4AEnfXfK+Gb2zggFCE3fjW6VWMaVcy8NSQo2zZ8YwcCgLrBLpFr+oOA3P9oyKKaCt6w8gDttaTcJ
TQDUncbUtc1Q/wV6nfSn4DuR0/2C7dIcOTtf4+d5fWC8p293M3KvxGwAvVM4fjApdGCThr+vwYHb
rS/ZYdPkbNqn4+mk1F1lTINZr2VrP2VxA+Zto2WvOhOQzeqt962o5GBvfa7B7asYPoZZN2mqUePy
OSpMK80GOs9kWLC7PYRuWR4KSNtuB8D9GALNBuOVtC8c+IBXdSrlraYYfFilI7gA2kRmkOaodxl8
M7tUvnAjaFMAnkzEltvFRLbFxfAPWOenSIqjYKOd3D9RO+IXrqEaw0gsfEa9FCcFM8Nb51q7RYjW
BmQ2HdLpCk/l393TcwHii4XjqFvItkqf+0GwETrAo7CITuG6YRin1L/0dn/WgnYIBiS49XUmKOqs
aK/SjY8v1De8hAx+tWX0DwUDLRXPNhair40Q9Hex4XQLmZT5/BGQUGX4OAwEkGZV1KUXUAVIdqDm
WIlg3YJXDbkK3ZVXCRqy4BVcTiBn5+9H0k2wUAwJmPPh+xvAmKzH9pwgrYpoerQ8bYsXkV5TP3fd
7YEMXHn3hnH3PVyp88Y+cbpJIZNNPWHFI1ubhY4EkAmRioFtXpqbXj58nmKTl3p/UdVbyhY4foh6
Q1s9or+EqHLXkWR+TCmcjv3qQT5jHJEez3C++c27Y/f1hSdxGmJEwIb7jUTE/zOqdpz/SvFU1bhI
yh6ouKZ8Q2Go+QNot3cORsItiZXwjNlZmCo7Ii3pNg75YIB8PALopLLbSztaWGYgAzoMAxINMJUs
pCSct2lb3hVpVX1XxOEEGegHGKEPeHTyqn/BfD4aoLruFt13dxhwjLn169WVp86l+D+voQSltMpF
KJHXwBye/+ti7JyoRl98Px7u9b5SkfllwnLgJF7A1J/F7YchG/j0MGAhr8OxVek9nEe1eOPEC9WJ
4jnmlMWtVmlY9QQuRA8Zs8dMfYp/2vPMR7+BPj1YSFt7AtSgiYSjaCflI9+3w2wPl2waC+30ydYC
+uvlVaAs4BtCLmdI61nbTgdWRLsCAuGeaBZdtJNs3dn1wsNFD9efRvK05DWI0UVoo+Reive9ZFha
qvdLaqInLRKdfU+isopSVnCxB9x/JLxQQm7g1lc1TgLQM2xpROPFywogFYbRj1DTojCNQ3EgMuM6
8agrio5FkBbpj1plYvgJd/pPTIjVT36nhwHN94U1rLo4RqqsgIW5HIlo2agEUUXQujlTF8QCCROB
eTtW2KvClz4Ts+XZn2itHDW0SBbwUWUDlmpBxjWGhskW8vX2FlyIHeFgnucADL4gNuQ3QtTg0YBq
KZvGky0v2VNzYGclE8R2opia04COCmZFQP0P6wRfbjj+5XM4KM6/zo5B/EuJAsmbup3/FUSjFZJU
WCSpPLTdDiQ9rwCMI7YYEyVAu0zEF3CF3+a/liH1NPMZJwaDAsEJoBFcXg51q5bfKsV7FEyD0a0s
r27XvEi1bPHYPtl+dyNVvXefuIV/qhsznaexYGtuXsSUHWgI5d85hvEsKNfI6B6Ny8sAn037CfNI
6M/gwpeQ0W78BbazHzxA0oBNT7C9nxUvb3Jl2i2MzcKc+WCozpeK9t096LGNNJ/aj5qnzzay5Org
nRktpzLYbvl2j0DFRi68xNeqcfw2VCMkWRcymcKGUr88eWU4ssZzItMrCRse0ZazpqREa9BUZAgr
+BlQoMu4R3s9OrKoZF/1d+O7Ud/uUfCbKtQER0UdYwVlO71bH6h5DKatmIRmrqZ6Pw9gaPli1t/8
xyeTHQFOcqxhwuuQxPNhiiSbK4sKic6EcdllJ4SKr1f8DbT3ZUQiHqHS/SfsKxWuGH8qDo20QGAf
bY4Zj87upX6BnIzJgtTSwuIwW2xU6ddreGq0E/b7Zu0Xz4ITiQTjoShufv/gPcryKsLUcqp2MhPV
O8avAmp/ypsWgBQbXy4UcVZJkXCs8iWyvji5UGBETPes314g7h81TK7WW/+9UK/wVwGt5xo92E3p
MbmJ13LDby1IGBp+52CCUWFVeoqdvhYJ5CwUvdTXdDT34p88MGeniIMZl1wwuZti+VnERmxl5g6B
S3KtPsPJHJubT2OEmOw28Bwwe5jAy/bZ417xeovXi0P0FR/Hbz01R7d8O4LRkvwnuf1BuncvvtxZ
KbfML5V6DVDhlUJycoH8rCJEkW7TGUAqoERnqdzV9Np7VeWpvlihij5nDsEnJAeZ3HfqRoIP9dxJ
eofC9n74S5J6zYMqTRS8iqyC6xfWTnsxMcoHIHEwAYxEhufWGvnQRMBtBof7Zib/ZZGAy2tdd7uI
vqfIIVd/crzta/7N+XCS2X7EJdWdq65vtd0jn54bzSYD3eNYrkBS0azMlUCsi1zWcQuKpTLDTADd
pBFy5ZjnY5LoKyqZ3rxZUoS9DPl9dihG+B2VJ3BAjgLNOpnW/Zmvo9Eye4L28NtJJ78qe+1rUaA1
e1o87z1KATTyrid23JvvpfRdBi2LmPgsVRvFih6L8726dexF8vtxJAmPWHXuCuamsqdb8aHkOTFK
D18pSd/Ntim9k3bgk5J7vubQWqOu8VN0QVro+CmkA8dAwPJ25RvQReCHfZAqYjiTHj/uwVM6WXKP
F2Q5Lcze1z8o1Kav7LlkkNrlVtcf+SR1zqj4nU+SPmD+G7DyXT4UQjzBqV62MyrOBO7hS7C/p3oc
ozbQfUNdVhQpUriRnpF8/GdCMQ8WgHuzWbBVrMzTay7lz60FHw8uHQ1zDPTA61ongutDW/3PZ1/b
urs/X8SUnlrO8tMNkW8fxRz/uVpBd+7OwrL4TzeVgmSBVqLrOqsvp6/dyf0cOsp0wRHhJ4BziHdn
yS0O1CdbOWqWJsRu2ulFirZNuftBZATxuGmlAbqzsVXA3pXGYuGid/ttCjXALe9FFefLDUrGoCN1
7JWqqTRMXV9ega5YGsfbOe67LE4fF8xu+AZuUsCxyz2d9FHS8JJR4kqt0KyUg2TUPBhShtRfb3YE
OE0MsBBr/5Nq6TtvfAZNiKusauZHWMBPxCLalNJ3lnUMvxuvSKCZY2+GowqjBmN3PZN22U4T8ZuQ
ITZcR1bi4ru+juROejJXvpfWMBqUnOsKtSIRHq3JkrcJmw3VXS0urYLeE79Cqw+MJOfR8emhM9ee
7mgzdubnJrPTlLCVBbhGRgm5UL85ZbfBkcwGEhUb3VVOW7F5a/fbbxvCILo8N246HsFA6uQP/Dz1
+b3OI0ZvKHdX0BMXiSv3a5cqU1fsFSNtEDbmy56IJEb0K1RlEfL6PJZ7K34zC95Chnybm5YqnBFX
kJrCDx/5LCYA5LBJtruDgZF+bYaaMmk9x9WQid6QuQ5U4Ykepd50pPob67U8KOMbiYnRJF2/i1Ra
82wIM/mobQSCzGrVVb1K+urNA+GIhF4yop4hxHgRoxNaid5+hzIbCj/GoNGJPF46922LpWbgA/J7
5NMybyZOQxWy007psvKmuNzo1FG9bFVag6DRx25ZaCs2hN2aHfDkkq03/3pY0rOIdgASd3QChOQw
YMsxRtxywxUFHMZgnZa4wFp51GV70NwGrexxGdetdttLmo6W87Wc5FRT0CrutP4MekiUG+90SCzK
9FCNY9M+Sgy1u+0JGSi1It/tXYWUUBscOJhZv7MRjlFbvzQktLcrOJP5KaFMyStWGYJdbz9PHDPW
YbiF3iOnSQnXUqT9Nd00K0ERDpbvOF5Kmb2HHZ7n3c2RVvwImIyUeXfelVpPqDvG+9FVZeyNCcrt
nLznEDgLpnrx9Rg0lcsP817QDR+qBEzyPxvq4/nYJiAhics65j++14MyySIJg1I5vomo2wELpCsy
UO3WlQXl9n7nv6At9h/WyHHpbJDDFSNntNZL7viwVm2OkpxDgsDw/vO51PCvYG/Km00CnFOZaT0S
tIsomgDSGVt8egnL2ybhQAAdpaNOoJwXXU5vagr1xL6iCAbd5r/TNVhVHl0mbQmgRBBuPtsPimGe
uFPv9FtrhWs9jjx8vXLkTHArtkhhaTUivx8B21ISS9WPhPBsQ306+gp0ckNiilM+B1pGch7d2Ju0
8hjG7ZaoiAZIr0K8M/yJZ363vPSFsBp3ONhMO0Lbj/0iBJCwxheEssAsVNOJEn7S+icBWIUeenSQ
crphaU46HWd/YYUvodjgNcu737broG2xKg81Qy89io//U28FLlCAE6F+zIK0TXhl4+ZFQp74l2sX
bKsRjrj4daSeM5KUbUESIexJFSJWgQ5ZRk2ZddXJMf8LQd4YQZJ161kcbMwUuC61N6Qyh/0R5QA2
inWmSXdr9O3cQfWWaMat8D8LfavAibHM23vCeO3EMmmitZbowJxlmdHe7I9ZI/jXJTjwGCtuY424
LW6bkoN1Tiwj957QH04vakUB9Ej7pyT5TPJAyx/C/vNcQV7v5b8mZzN63LAWLU86+huknlGHhi0J
JlMj/h2ADssOpapR8lSgQLzxvVVhhH1DJfkba9epmT1Gtt3TMviJNtTnga+ofrRnAZCerbcbOe15
F+oj9pakMpdY8yuB371XsRNrgqJlt6DJHO0/RmRi18nYJvpbFieCkwU6flTcR3if67GlJAPGrIUs
g8VPYlAMP/WEcFY7ys5th/tY8utaS2o+3z4hCEJYLJEkBqplASSj7Kypi2s6/i24U+qqmFbR3Do5
gTzb3QZT4PqeLvnISZQjWdOVDcUhebtwLUOR/7pbvkCrEAKKnybW6peT/mzrxYlEUYWZC9pPgNbn
2WjssJa5iBEKjFEsvl/xHn+GdZgN+08e8Y78WcdmHCkYTO/0xbqZuWJFRdTK9IHLDsjrPyzuqNgz
b5xerB5qLKkSJTY+Up9HzLN5pCGr5EVcy/dLd8V0OV0BqU+fgZWgfwhuHN5LjQaNFdciFnqbvfN6
owu8clN79oWaUf2rl8p+WT2oMJysc2MmeE1BY+vCATnuR31L711hbqJbrCmmrPB5o2EjEpVuBnDt
xpkaXDRl6DKgSeZXHeJot3AznnDmyrvpuICfG5F/icIRbV0Z9EPZ92t83L0uqVKvFZDw6mbKioHE
jiHifobNWquQFSR6OYdcWTQEnpSlCvF/QziofnzAu56pkh+kQSUXIYF1rSl8Nyq50ZVQBKPxD6gc
USlKlgK1mUdS9MNNHDZfm6a7mXj8nx78M88qLZGmk/7iHmJwHUMg9KyLNYUiVby8hQXDmsdU+sS/
0Xog/4SwmNQTAu6fZ6la9UYeG55DKf+Z1vVEdzvTrEMuPKzLRkMlDAM/w5r1dEoamJaE9jVIrzu7
AGObqEPh9ArEuljzazyPf9kEzw68W9ESwLVUpM7TyI5ho1gU0bfnRiJ1L11/6Qw52vOf9l7C800l
IGOw4xsBTCUpKo8dqu+2dJ9PTu4x9XA+nQ79erGCaFBybFJ8uGRO+pXWP2Q17bJq4SYl8w4W/7R2
izFsugJrJRlI14SNv1UB8jBNy6nXzdO4nnN8o1LGvYSsy/s5s/cShXIMtayT48orlGqkPmFI1T6z
Eo0C0CpfjlvzBNpCJtcPvgzwEBBzH0Q0520C9dOBDmGNjzbE74qFoJ2e8j95oWIW4kmE/ABze3EN
Io68UqzQWevXMTWEtEXA0xYDjuHBRM/sWeSK6KJU/7ZNVyDg+PnnoGtLo0l40MEvAs1r7aqM72Fs
qhVkc1iRy6YNdB2hSpwTncd3PDmRAbJfBx4RDLyfydQb9mfdJ4rHe/12HR+D9qqS0xXZUWmimtCR
ZP1Z8QAA4kagrLaKcjUBehGo5RtkSbQ/97KBT/zRzdQnSLxS99Moh/SIsYKa0vrTu1HGXbHC1kqQ
dPixoP1d39aUpoPYYnLsa1rPognRy2yyskoZIZxKMDs+F9sxazXW6YsPOSQi8QObENiaUtbtzqFz
/s1tEJW1q/1vwOq3VkQV9nQzU9auQN8t7LZlctjLE77s3iI33A2ZdOATe/ydONQGqb0fDP//liHR
WQzBui/fqJ4vz2J+CuXrRHh6GThBA/BTe6MrkOV81BqRYghbpantiCg+JbzkK23CDq2l595lts5x
mLDF1Iody2+Z0+PRsUfIS5DfvV4Su8titun5daRzVWs2Y4kfoIBZ5gY59aYtaSs9zLB9vm8ANd9q
W4euOd4+VgZfV/EL/P+X+5ZbBcDlPplo3SriNlv5KNx4KgwhShr8hgW5wJ0DcHZQ+xsOjuc1y1H2
EY5gH9+K2hlxPYOCBsj+sQXn0JmfaL9BhwzRnKq9JS0Ekx3NMLnsmKAbcAOSoN+6RUjAjRVj7Uzi
zsN0/j5dg+x6TygL8o7q0pmfRFPWU2tj+QBPD++sIPOeKcZwpudF73LgnqccOnKsM3Q+hLb/blLX
/m8keUwk/UPB+fNsjEdGX77RJ4BuyVV4yCGUZR3Y95Qwvl/eYb6we7MQWWPkhILt/sJOp3l8e/zE
IqOS9z5ThakE9dxcDh8mayNaICNq1xF+VQ35rtxrjzmQDSMSzarMBnGh7M7pET4SBCAZ7l6dIfyJ
BFZXIzyGDsIZ0pBAGJfLsQV5LYWBJ8xmIFKeAoOyM5QRKZYtAwnorCoaT0QCZ5+XdDp325spM5oE
pD+ixy9B1r9jpWMLiOL79Uv5Igv7KXBRWqy3a+65azb6CZsj2cMlv/sFECf9QNAxF6+zJdXSm697
T8TSjECUL0gtlUnXmpxmcFGCllWrx9v72n+3FZD7OhwokrhycsFLawbVuZOJNe4gbc7xo2acYW0Z
H/nJTwkQbC2g+bfFZkA6qbLjugWV4F+3w4PU6el5hMo8TTUAKCoMxlgrYf+cf1tE9/siYoKXd1dZ
HsKkrpN3zFHK5AAIPXXXPb1gUPout5cL1xlWQjSjjMLm9V66ob6cWjPrpygX51u/Qws4QVNGn1Pl
zxAIWPlmGLLVPp1kW9XUFCvZL6lBPA19PtHwqRBw+FKZ0wbATj19D2Gzk8Eeg4dBEP16RbkYvUQe
LYR+5gw4RxprCd32nWkHt7azmGesBUhkZVOYI759vsXqwUCFW7jqB0xtPZQgC6KYAr4vUv/ZFZ9K
4k4hJ3DClDg+e6QzT0klSZ/sRX+MOrXfe5BGPMeIveGpCP1sLRPZA4DQwGWyANlGudwwqt5ECYSy
Heg9AkKeGc6qL1w6G/2CbPZqutEHfOBCFAb0DZttsrWPGSddHYfBlowPTXmWdKBfpZgHhjjJgH/k
bucL4lxxv+QQVew7U2JPz2fGkIgzd9/Jh5IOeKAfkXGc8VImFYR/hswHyHQkIdeUrxb7OHQmJ2As
pCSKGBHPiZLBbB7EbvY2AAXr3qNymUGPtylrzt7+OcVsAeGv4S11vjRuCQe4GBN/BpBzvcdogHY2
o2fF7p4SYGQp0VoTb+I721MnGzJXcN0K1MeEP1lLFxyL8CdtqnnGJb/F3paO2sDVEK5SXDLtIkaE
kLpDFJZzD3Y8fDr7tb9hnxAcc0IP8U+D+r6wVGpDtSj4xUbr1eH9LZFmSNxnDPZHMKTnbHhch71T
wumLxpV0mKwv1vyzT2pHpeIqkaWOf658EvMSsq9d8dz6FEqkb3Exi3r9gSTLl4CKVJe2Sdll9Rr6
sNK7QctUAcbDikvOYBdY60MmYemucWNQ0LumpCOL5nP6uUZak2jvsRUYn93jXNTa1wHvOvB3Y7p0
WHMu67jnwzpudDznwxg7aXUo41ZBa+fjV63yECryQi9qwfgQ0ZDYCTE3Tmrb+JbK9i5eOb7Zn3ao
jMxVS4m9fe7Lm4+Ih/j0UfitYxN3pHR2m2vhxKZAHTQXe6SvNpzokG1RBiZ8cGKEj7e2vZfO4AnF
uJ4UKQIga4o5yLUnGRyHh3Uyc8Vm7EWpyViIeV4p6Cc18kwpPnohbrBaK6WupW06N9ymna5elvr0
lAhFETJ/Y9eXGD3ND07YckUJzF626sOM0mjpyRK+1PSyFeOMj6E3+P4FJT9vBV85L18W+vgGJnA6
1/p2QLbxV+SsLpvUY/NQCxwd2ec4qYIplVeiNGZHNBAa1zbse7hTAvCvf0/GLyzdj+UYpIpUD/BP
+aNJSAI4XPwiGYVHcqSGDpuUn6xL+DsbsluO5IeEupIg+e6YVelxcIlQdT0PGUwXWW/GEsypp3VI
RhXjYM4CQxCXgZT4Xxm/r0ZU/qpCjLkOlzzwgHEeTKXI+MkuM9fW3gGC857rX7mpwapPs3tJ6BNo
vZZ4qOF/vwP5uoiNkdlilN0ldwUlkvC5hYOlknv3Cu3g4mTvFd6dmVMSO8dJsgPZq8aomL8ds6an
2f1VLc2hejCk+tyaKD5Tc7WqK2I2fI9u2+tYl/OG9RjLb7j4wQhGH1aj8dJWsNCeEpwIvTldH/yY
wkTEsLC5DZPw5Wn8DmBDxsf70gv4BXSekxPoGp+tHaa2BPg0cqFMHKP48XKnWnQT5QhnUrYYF+P7
rIzRTLs7GhvWA7CWGBcVstA2IEXOVRy1bMKitTU7fPbCDicEM1mSy0nunk+oRT0qY76qtyUO1KDr
YR/CDvNvnphDJakvq0Fr4n3WPnt+PK9TLrMHnUCe0pq7WjWMc4RTSm2uMVdHAVJOx8l4+ULf7IiN
r8p/B1WPPijTIrfi4Hm7GT+EQzmI1thn5FDM+sKG+TXZXoA5FSFbq3RPPBTfFwxmwx2Pv6+HVLIA
nVzsRi3GvNdey+5lOcKJtuwAhuLvWaNBK0VLC4q77KSYU/7BHNyjikIKRCcCFt86mYvkQxygJH+d
VJwWLUZQBYGCZ7NJjDiROpOtbma4Ccz/Pbl5cvwQFrzrrD0TDqDYfxT4lBS9PXrNS7nDei4GEWv+
FzNHAE2ZZ8JM4i4VRdSQMK2Alj7+IQ1l2/j6Fu2z75K8CdN6e2UM9Ir7TpSETh4Qv6bU1gzkseWN
nmKtsJUmCPRl6UQak4iLbXLmJ5lTVoahvCK3yBPh40ACyCvkVVhfI3DF4PDgGCKZZ+boqJhW2Zbt
4r8pVeFMRsEuidc8nJ6VGnyFNxZe82hfyCzs3gSwXUlAVrDZIxAR7EElsP9zEZmN6FL7yLF/8BRn
DNyqQxC48xcDurkONNfWoCLKdc9XkXtH3g+QkhmIzRa6FZUadY2gZc8xIlPIhzR+cOH+eMPRH25b
1VSr2icCoRHSzRGzSFxNkyHekuFNPg6QrCJtTfWXuaOcKTgNb3k/yc640PwdWigQ2IVNVkgV5UMP
X6lgRkJ0VFd0+5A/xPuHu57TrxreiZxL/t8zk7Dma0KMqpHGgHjI31Dzf/PTunoYP46FAT4pbwry
dMGmAnrXw2iNL0qttNg61F3ca55n+sbKrY3NTBNA/1kOjcB5WHW07mDzdNauX5kdaUbSKng5jRIb
n9j34i9d0inMlgf/+FHxRu5gcUThvsNRFd/5PshtYd+1k1TBm738fJ2PgiUjcD0qObE6hnStCozR
Cxuth6+CayEvL/mV2OcO039bVXn1ZMN6zjEffE7VQz9FdOFD11gt/cycmBSqhIsS+d7+G2TtgXNO
cIUAREV0uPyUDVHdoDiufdZYC4j/xLrNpWmCYJx6z1KcaS3IxWegPqxl5ydvgOnEPfUIo8BNpzRw
Tsgt5MppZr3AxBkae8NQJo4YvrA+4vZoggKnbNBSHcIUbmr4AJLaBwLLJdQGNgL39+N2g5UE0zNr
W0xWgy+rIXqUsUquEoMB3pP5RsaTIPGtCagxrC7yfJituPZyNaJ4hpenoTHKv9n9vFjd1QW+yGU1
DG+aacqHqN/gVkxvWfwURQJwJ30jGH7PB6xe4zIWHa50mvihEwMbbb17LWnKUfloLJq5Qza4Nmas
wEtn9C8pA64F4JzUyh53AvyNOb8HsLI57DYhqB8cCVSwSbaB+7Oex1xqTdRX/59erdkMoIJy9fN6
0Qq78FnEEqSbY1wDMzFxyVjcUvbvxEZIymQI5lagISkPgkuwxS6AO6gNpcmlLPix1Yz1ipBS9asp
fswXcDuwKvQnZKbUpsuJ2AFf1H/qmKPCVil1sOW/VwSWRNxiQcE6+IAsPuU8muG76Yuav+huhFhH
Od0xPdjxr5/AltTvXBp+xXXmQPnj0Fz22WkzHz07PWLfVG4gA/7jBYxCWL9ZpsWmFPt1mVBy8poL
Vrpdwh4WlNlkJ9yQbYCQUl9c5bwLRg6F2tElb2FalGaJsCnJPBvt2l1bft7a2G4LyJQ8i3oTo9Jb
E8UczPAZmwi5VMM97ML9PqQmtxzJw5Nyo/rAlqn4aV1HVMRDwpXX27t+L/+QmwJ0QT6kfApfiHNe
1m7RAz8pnOM9Qx5AXZLdTlOuSeufqvszEUaDK4fStPeS2F5xeBv4uB7X0vzJeelalmzuSRulNp4M
pVdsesW1tVXkvDJSu0DN0n2L8takGM/OyQzfJKCQb6BpfdyDTNNwO23QIgqJb6G/vUC7/DJ6zU0+
BE8BKIeeu2BFQeq5XozvJETJO9qlsv3j7ouqVtwwEVREVB/YQwP6OKRAHtHt/1WoVSYFulEmNHBK
o2s5mesF6P1HlyctFQSkROSDGhkokaUzuHfeoWCd3LTC3mkcngySRtB1cvrt4/W1AVO7m3I8E8fM
J9anxhVaCxJdPfxvsZFD+OTkuy204Ml7aV7ETXYSZEanLVddUtHY795YDiTIomtpH4PrYoi1l3Oa
3Rf5MSleNbD4Y2KcBXvbT1KVWqYkix6lc1yBusoMP6xmAY4YKH9Y4dqZBOT50Bo0FWmFINZcx3li
86thCZ4E8nK5hLqjes181tke9EyCnROwTma0VS/pdnb13BAuuppdGj9Su8lqHVSjIuKHhEF5Kk1M
uyWPNd4cKN/CtXJ8lDOTjahs5whwKQesBYMbsugOpQMcGapWFXll/qkHsvkwoouLytIKxPIMBdYV
ki+Mg4Wtjf5+CErijy8lZwrcOoJbe94XLSLnIo5jvQ5sOPvNA0lM8ourd5KCGONfUdKCqPyD4WmW
8niWCjuLEM6oqyNl2yoKv7sVgF2Seek8k84ir7DSOtOH8Cg8N7K6oxRB65hed7GewJA259KtyVhz
EM0FVjZhRX/OIXQItYUzBHSPniaOjQvk6y34sAWD5TlpfUam9DoouqxSlFknpgwCmUDpuF27MrNm
T+ArqUqEiklqA++TL0l6sgO3j+YnH/5bGuuDnKjfiFY95OLiYcWS9p1qt1vJ4/Dy+6Uy+Vr5a4Hj
a1Zf3e1v4hIKta6z//XAvyKucdqNxVNqrJq0ms/MXk7d5wzN5lY4NBj7jIIMSK9Detvso4+RTyOX
KlKpzXnYjPTRyd4XZuX0Q2vf2tJoHYwZF2dL1gIeLoWPVFyMEO3axrSUZZ8cH8BsHJFBubfMPnsR
xTyLSmgrBfGkD9L7CkWQqJYmYl0kaW0bYtXtTtWyHHvJIyeFdhXyg/a2ZOH4s/mFEXuSsXXKN0N0
ekwshvdNfx2/Owd4FLXvrbwXmMnLQKCeAgRhvaAFl1B5VluIzyyQc6MyDDNzUrYXvKiMdh6S7Hj0
xfv6nkforhDXjMXuHRdTBGAbitguS84RQErXKxI7PvyN+4epfyZvokG5qLj8j/G9jYPYrE+ok8tr
c9lbfulQdU0qUgEUlS4GcPKV6lHWmbVR9u1ykgFRwDzTLk7jW08+vP15EyD42rkg6XO8F6JHQ91u
udSLYm+TCzD+3CNJRCm5c7a+vzDm9nGeDYKuBl6IuFCzsb0pbz14/Gt4zKAU+ltwCN7l+NKDXZvu
gVV/LpbxfIhElAq5yr+NRMBX7xH9IvF0NhpGyb9fcrnJ9diwlsxP2+Yp6CBgkVakzlTN9yHqcxN2
z8PaBZUiLgz1PiyD0GXDPNLtdX6xneACd2/uOB056nI9SWynDHrcjHIEQwZgvt3yewqD4jew6Y69
LpMIlybLrkDPyO+zF4m4nCNvwiI8K3p77byKzFJ3NoYTrb5BSA61DZnMVoiWXGRuhLBMemWLaY6S
g4CaB5dizVIw7CzHc7P+jFnFKaDQ3nKDY86JPpCNlEADQMo9C7j/kgo6gpt2SyXIECzgeaEbfFKu
9WwK9vOAV1E3pAUYyEXHoW1/NE+ELPgslZpo58QynsTjQn0H/Gpqor3xF/miuXkYajPCxq1lFbRJ
/k7yREb5luer1juxVS4o1YfxnYrr/qDYlPxUoRVaYJidDksJOAOTDfGTsFgW/mLclFukjRq/AjmN
O/Z7jpU8XQp27lw0uMUrRYTSjY6XbZD1XsrnUGwq6lJn1jndB2q6i1YdR6ss4nr0mRm49jwAYeJz
ZFWYGV0XFEo/B+6WvzixxTeh9i0mCbAstF1f6soju4S25D+Fj8JU2gJroCQEsGx5f7hN2r+WJp18
4rwmujid3P0ULj9bdEvwx5ukljNXP9b0n+kC+XIQV605tQ3z6+E+6J7qcZhCeLmayx5vqWt+QlOn
FUrONVQ8VUTUhuJownkeU5L4R1HGAGLNB9OY/nrw7jm/b9TADHaI07roGTGgI4KzjIeTojnCeBk5
605T7oCDXTn+U9laIjFlu8Neoom+dIy04gvr/r6vgJ4hVw+Z6I+1bT8OYpqhD4KGAIyceqdUjJ8w
mKLlesBhjlGpv2hsDJDgOyb9jjxf3n/Euzd3ptn27mL6KRLx5t3EInlUw1JndWhruDkMBSRq8ea7
4fGQMCNA21Vw+/20MwnF2v/CwbcBPhTJo2aXdUnsyFqcRskVPyVxCaP6wAdens2yBcmexT8J9tfF
gdNOJHy5fL5HIl+9ToVruj+rZUSf/Ns4PZ2ps14eHuKDBdLsRgLaeA+hYVyE0LI5J4uFjJRz52CG
oDD3sruV/bdYpvCPGwTNnEntcJ0FDnYy/o6+ylZB787s/lgCPdn8zQvb6OwFCV9gJJ84S7VgGGV9
Vo9Pvr1qtazB6F5BgXcaYVK36+UFwayZB8poKdfanTdRzjQv5UuBjpzkrGkFM4iQj9XfFQ/B8ECz
k7JdWnNaHDBS9yBa4ucVPcv7kPrM9pDUIaYdhX0v1ZaLJvYu/Ip3t7XoIMLSbs6eI1mzvwXpVjS5
q3kLMezKIxqKYpAUj98oy4Bha/3jpSlBsrC7JW98wtBw3eS5PsNVCb0GQKu4MwBA/Bqs2t/1cYca
FX+aqt9/++xoOeWbTXiU0dcP6YZvomJCG8gAWng9nLUOFKgYxtZGpRS+QDRp0ZF2Xs5V8kTUuK6P
SW2q7oVC5UCITMr9rxJ3pk0f6nOFu4fVEEBQklflXKwVw3E6NacfiQhBfUatgsJl3v0pPv9keczz
5rKT5hvfp5mghF5ahwdJGzWZIrQ689dKIHKgGdjyl/nEbDWZGaf3M/6gj9bfR4+AxL9HXuhABGrd
oL210BHN9BJMSyy7lPf+8HCMVE8q0/O2DoLFACLy2YyNLX4etgXwVasyHKfeQxyTfhwlnjKdsrGO
Gx4//olXhbL2teyr1QClc9uXwwaaDXCDwTXtRMccP0MTFUtV+6eyez6uxfgtIR+rZbyO/MrekBhN
QEy0gmaDUY7+wgZSWYnETxtd7eknvXtOsK/C4U9aL0xR4eEJbNr6TzPCPTJTAX3ds7qGXkMwtgv3
ukeQkMP1eKApwf3e5qJML2DkR7FJLgYH4UkORbpaaDANHFddmKgmbR0Kw1cbREMdvRHBh6AARcm9
fdZikEoC6FvMEN1Bnuzm8DMGQRrybLvfbChx5I4TGUilVOIlhcy78Qr0YIHNnYkZHF4vJrdBtWxq
5JStXvNpQiKTMusvR2S3zDiZsab8/emRY5BEWozibIRMkgzwOMcHRFfIFQdDl2H0TIXGQGy0IbEg
RHgG+nHudHBGZm9tUtOzO1gLf1GWha1x8xosuAOkGv9fr7hbjnMBwyt+Hjs8Xj4EISncCOVIbjxN
rv2jT1Q3ubYbKs9T3IOAwPbJWANh+0uka0m52MAyHj7Gk3Yatf3WB/hwFHhpd0VvjgsG6vhpuGO9
PwCLyLv+PGwZPrh3HJKTfN5LqikC3Er2D83++r/yYDFl28b2xRQinHKuJ5SLsFGkXW8nGMtngkNB
rV1LdyRdPXB4oCWcMnRVy5hofSasobC458kRGFUxkYj6gXq+N3G72DuEHkR+FH55FuztTNmjG2Z+
yb7OGl6DNXZkGd4MisVWV2eS0x7GW5PvhfXFGWtzFIr2yMw+HiYCA9JQyLnafW7/OSmaS47pjjIv
W1G4MrRejFpS9OAR764oOKkVtzOwnV+/DG9FCB8hjFXx76V5UsxZy7ourE6isUuyUUbEo1z5ytd2
VOyJ6syZxCFSqeO6YRQvFZP8KkR62tSBAxPfe0vj54atFGnSaiSlIbFcL+d0thci6Rbx2iEpn5qu
Sd6eqyDQHl0WfZi1mXjLGrouu3lRxsBK3lBP/L65CGgJ42GWZoYoHsiD0TN7fR89AqPYmvP6tRyN
IGBLrjSH3+EjXuSGudzZnlZKzgGraP/jWSLn7dy1q9nR5Y7vccEKlFMSG4cRCJzINGV/HF7Di66I
6tVv6/GE/HRRl0JoV/wSUWxtxusc/PlC/u7I/KSWJLYP//FmJu8A8T7RC6nBeRWVWQZIhkNaCUod
iU7oDiE4i3VAJst05B/wr3XFV5zkM72T13HXW44LBhdgojUr0TVLUpNPmDfbRl9r+Weqfj6Zy6AL
/+MFvTkDMi+LcjW0TpOj7SipcXCTmWDiVQHxllQFZh5yWdfn7RFhFZEvat7yOOG6vWbuiJmCcxpA
ny4znTx6yjXInYEWyJgu7NE9ezL/zz/mxMxbbHlLImYj9XjY2hrCZkTCFaE6BMaM+UWeuiREgL12
gCv92SyN+Mrg4g9nR/pOkieB26R9SfChUa37gj86b7qTK53ySiX5jT5XabZ22dRQ1rKtqrVF/Q+6
ozBcV9O9T+u+q8mHWTBYHjdg0vXmF8ewNyordBu9l51efNz2EBUwCdE2kBZ4+ExTNwDDLuKUeExW
4SfxQ/4VBg7qov058DfFg+ioVJ6alZRdYBft1fv/+nQ8HoYoJVjqUZ/pzIkeV3lFzYow3ylfEX3y
ZpRyC8X0L/R9q0COAmvUA2HxMXvBODHE+BbcZ9Aby1GPw6stDm3eszu+2ZH9RLGfhEmSRCAsTGhn
UsvDlSTmaTinSbBQ6xSeI1wOCihQ27ZhewcEb1J6laX5SVGsg6qCyGD0EAfUtIRmxGdFN6Ya16VW
RJyZCcBDvMZmoKqG9k4qWFVPANDE+1gophUYQ5Xnikn/+JapMiB42JZzMTsvn8BCawDyjEAJJQN/
krhgftvXl/mw1KRsJ75CiPNdKW50oGrbMnelOhYOnrNAD9JS9GQURH7Y6ZmMMBliSeOssMASTZqy
yMfRLR0Kve7wjWAcNsG38nsDFyuzvZNLoEkmEnd0zVYpq6Shq93gqSNFB8/g/lq5jfbMU8/CFq10
cj8USx3J2mTy9WwFNHKEimjE/BKrLB7ukCCrsvG84OO9vRyqHb/ki8UCvX5boBEBfbPSFcXc+knX
1mWzLIlERpQwOjBu4ob2YBRk9wcyvPuRMR0Z5Jpuo4f5bM65YHp87R8As17GGvfvYTFizDuBqu5f
6ma4yRy0gjBPRDBgQqRoqqNbtq0p0XAUvcl+TOhe9J/ZlPCK4aX9zHW/tuNz1lThadEVm8JchPav
/vudkq5vPSmnWErIMtLwRYxQ1Zqvb//yjfD61w0SI3+2yTLgQwl42bgRj1pLfYJxHLCXfdxlXlRx
Kq/S/q58ScoWBLIxKREIkZJGFD664AUQ32VUurGeixGN3PMyrlpm++qNc/ybtuDPiUlj4yzDp0Uv
oW45AGbhHyDL9RgC3Ysxnm1ATNr56Je5xEJsI46c9qSHFr3qbR2Ufqr7KqNkua3OVvhOssAsxAS7
PvMI1PvUles45m5K39eTo7FF1kEVKlDbmgrh5uWrxFB+/TFwEpcD6lFUDfSgegzTioXobDvLUMYy
aQ7US5H95kM7DFhe3PmMFJ03VOtktjEYhNNnOcD9lEC+Yu71Q5IZNIp1tqjie7SemlnPBeU14vc/
HXV2HQoIFG+EXZBIO8duYrLZDjp0f5RmB+KcJvfA1T+MNpDknNa0WN11BKJeNgaSJcTH7L/SO+Q4
xMfnbUPfaYJ7UlEvrkCrhkKxwhIHB3J24BQeSUuqO47/luSWZZtEeb8UwknMn5gQKfnCQvpl2cGM
1SfvvrXm5DfFGOFmsat+2OGdDqSP9EIXq2ddCH66uZk5QMSzWJ9/TmkL1WfGqyQyRXDsUHI7PwQ7
hUxmLmhhkjXiSSFpR5gWwR0s2p3dxMnu4/vwL2PBdzlptSqPHCNgQZ9KBl1b/azFGESslqauDvX2
oCoKLE55DmEedNqRCEnBxRYvJO4AjtRS9Xqdu9r62iF2DwLdPlG4Jgo7gzngyCtULosOkoQzZSrV
PRpW+w6LiSmtIBZQX8Z14btObVj58MqgZOlaQpV6Q64N2oLZ5x0gRBvrhQbVLHycZc2o/lwN6C05
VzKRIoJq35h/1X3t5wFFaXXATJy/d1lHwlLMKwmOr+t1fss1dZuq/FsYLAo72h0JR/zukBqIoF4p
avWfX/uTWZBVeweoy9+hbl98DvdlsnvY+jSN9vl48GBugTwKA9iaBBgB0ovRQxZnxpLgEADVl7qv
WWaLZMaqTf7CXLLNnL9CPKM3Ihb93ZxVojHRHHweLrea2RdGI1MXWx25vxPh4itAks2yJR5sGnSM
lxMpCQKAT5INDfqfSVRVGfLhBC0Li/ujy8sY+3r+Z5LJG05BpnuVA6IX4KU2NH0MWJ7OF3hKTxHQ
ZuhB5o9fSirU4fgNswCqsTM4bY+WrdjaHabkGR72n5b4WUkDR15pNfAHVY+b35NTnFoCuJ9D1B1y
KzLlJHvsohDUIcYtDSjHi9l5J5tfloVNtaKxsvFU7+ZPVVDKTTb2pu4eV//lfSCHXOB9mF/nWmCz
BAwS0E1/S2KsJD6rJ5dO0hplQs+eR9sRanmTid2wd38ymr3/wEJaI+xp8kiVdrowMGXcnuvJzSUz
ETWbDBK09j6MPShgJUALv3nvif9fGM1Jao/XgIG6Tk7QqkgDR3qUdOLxfSxY2wmzrlFAg5dYVuy8
TLBPx943eNV4S354p4cYhcsd0s7zt2wxeccrLfYQz87Di3YxQCCiNriJHMbC+BZSwljtWqrfU+h2
xCeT8Xr/Oat4JAc0DqC5MN+kDFStMH39jNQEC0WbjE9p/yI3p9xPqZP45P87YErSU+a9GBRDieRu
Z3TlykZ39X2ZCJlYsrgbu+FS7F0NHkjNUZ9eVC51Tj7EmfAu6g94lQp+QWS9KJxUaunOdBybXFDA
jTHmVIVRs0LpZGzf4BWx00ahsMQwi99FnvEo5Sav8A9CfAx3VQ2/5IQcYT5V0n/FQFuEDKQEZ484
JMMYtjApgcb0JpzYSng3f0le27SGJgbdWRi7SyFrNm+PzC0byC9d/ZGCDDFUf5PCv258QmhEWjWO
TljVDpvnA6JUWmIdRgLRGvwszrMSVhRc5xpBikC4r7DouDkB1Y0oAwmuYqYeojDt6xmHqcovICVs
cb2S0G05BohynbJFg+uCBKMJfSxAeJMMq7Jdhmy7X7BEBYx0m6ULrhjmeH6OwAV2edIDB9HBSO4z
qAEChQHyaOBfL1yjKqcLSqcgVQC6y5c5noYqKPntRgcgkBVO9t0OYyuWh2jwtQMiuyT0Om0mrFIk
IAi+iWPWa3winOqmWKcN0/9fUn8N8LR2OM7qqPMEIjvmOK0s1Ywi9fNT/9XSOY8m2YthJePHJpof
z/9V3Yn80NLXKSQfaGr87BQPMpzW2TGTm+R4Fcmbr3kOZJJiE55s0bJsBJBk1JtnEF8uB3rIjmzC
vyTqXE3TrLZBhanPHr683JnV2cHLwr//Zsu0Z2I+VQ7E5Dshp92AIT3lVNY6XHRX+7TAZFzGoMOy
vLx1hWDKETWLPIPoTa4y86v9T0vSVhwqW8+c5/cAqy7QQYS6fVbP8B2ILoYz45joIdrUGZvRDIO7
9kuzK6Oqb1eN9j9SX17I/sRvW0uEdQqBG+u1fAu+xg/2tqjGqqR1IGkBlDlAhE1h9lmc5j2Nx2zg
tYYHvfCj3z7H5NFhnXlZfO7RV2RwvQ/dDvfMuv9O1lpJgeFHHzhnMzGNwJQXFoyENZvCCpSN9X4y
WJeyaDKQLB6JQG6/tcnS4fC9K4pZvxdfos1nVBoTogpJrypiveN4YY0lGfdo96bl/B8TaFs77RpC
mZfPLhcJ6n2FGeZYajEWI6WzPHgoeCRe4WWHtqf7/GHmRA/PUf/HvCM8BgTuMnLQ/w3u/V1DlyCF
7Prlal92Eyb0P7pRzQbvV+XaGgtfOkVmUGBGuNYEnVbL9X35GIFCrmZYA5OyekOvzlvMUuZkuFaL
S7H/A31aHsg2R/q0Bru+N3iCY3OfKDT2Fb3AOU7cQ2qUomGbwPVTzRM06ZCe6BW0YR/n9Tw75E9E
GdDFBBbBhu81xdJ7S9xIPK6YMuSdyh5UiGYDHNMUSr5ktrZzzM+JCSFfQXevEsw1W+GRdmQVGcD4
ef/iyBhIYptkJhgYBKVM5iXrhNlZlD++4n1KW7DW+c8cSx3E2abSP09cUuGo05znqgFY1zqV/Zum
l12bE/HEGZDceRARgWk681BAC+AVxhx1iiuvtlnNzB/C40DR9l0YQmvGjIZIQuA47t6HqQ7C1vKi
DW4zKVUtHSb11y/MC6SfvteTRxPVFE/b5mHj1ZaOkN4YzrFYayj+ZgWnOuT6qJ7FpUhY1B13cl7n
PxKK8GrwzUdbvMrEmIV7mZhmnUhY2GmNlEpRA5KkrYrPs8sLGvzBrtptlr8KRsK3Yu4H0RIQJUvO
aADGfxQIys5L/ZEu7/Vz+oK/84xpQn1N+tWovu+OgzwmAtwx2INo86SFmKBmzxyqGafWyW8G6T4Q
Jyqn1osdQH9628/XTGUBUKPEf8KA245wA2Gg21Al1sjcw9eK5Ln9uZQhJoZSh/KdSXU8Bgebw9OY
GSMDyebc24Z6knZOpe35oGr+H7p/AwEvAtBgkAbWy2NY5jW3wP0/n/y5hzRb/3V9E6BO/dELUdnE
qjET7rgX4iua+Z54Rg6M3hXiaeupcBmyAvtgh/nTC9ROX2Ia2A46b2Rh1Oi38V2C+wB6Drdh8r5M
7IeVbnBXUcbH4T5Vc05mhlPmw59Lhr2waYs6JeTd3/UkGfwEQg1UYHo94oE5E9ohtvuOMdlNDIAw
XmviX9nOXwU8/bCdOp4+QphN1vWGgjIl5F8NnMtbZnEeoWyMUIhxcn56Tr4Z724YkWBDstlD5NzT
9MHrDyfhkd5f/1PU7/sX4Xlq3sh8Mp9AYIPM6Mr5/Ca8H2feTr1dQu8g/Otj8zXUWM44D5oX6/LV
NYXadULGuvHhrqLsowPwRM3dUChic2ui4q2f4qBSQHDEGdIUYOB7MXvN9s+DkUPJ8nYKTyE+UAAp
xsIKc3kORVsZrie5GlhVt5ifOMM/Q3j3UUEg3CpDqoymhyepRnsCNGCsEtrzTCEBGvNTw8VMcqxH
kKbTKICmptdrc2jjmX2wr2spk0QmmlE7ASy+Q1weC84FHBicITrLY9GeDofmWkIb116Cke4w657M
14wAvcTTtK/0Uf+a3R0ZJ3/wTy/3MBiTQXb2MU9PABruqMh4fb1DruvpfrM4LYXNb1u2lFJSiCgx
DXcvb5UlMb/V9zVFqDah5SkGtQPD+0BFK7QbClqCt0K1wHBGFfWwa3xr0Ib99CorOjIwuwo0HLgb
t7gZ/dT7vaI6xuhgZ1VS1IpQXmMJws+GZPSk4TLras9HfS8kFJNEJeBQI4Lv339txxGKfpbxhcCt
ozokd26zCv6PoigMngsh0pf8iKOHob6FaIAmhIgO1PVl+puiT/wGak6DmSeoBrZnZZNh9GgBISKc
wWBC1RrKC+LnQVuXZmMmVZqCyWN2x1JnOQtxKlbzoGDNZVSblEncz5xqTxATBgbVveU/XwwrgB/t
604/32tNTC5C+7er8B9iIf7mUNNck8Yd1RJR/KIBrTYg5UvUq6OoqgnGiPzIUypzHLQfJeoa6/eQ
gtpVUX5ucCLj4qaEOohMNrjHoITuD/fgDfblfuQmA5C64z6X0RoeqH4UWmLVL/qfSJ8z/3Yzm1QS
UsyCShAbSjvgENEEip00/Q0LsHKSHKj4dOYiBkXF0xH6LZ1ndfe8KtBbf2LptexiXAaDSfw+Hsq4
xHoMvIgQfkzEGaOCzBqCDmFr3+pdCQkbk4EOmKVKsGa/QY9SyPWmwzeW9vcpnWs5XsJIIQVA9BPo
yrBOKpVrNkwB1Wb4LdXfAvQ7Ma+zk1dOLmJkm7K7E1J2JLXyUxnaG7v1SF3pfeWm1dmjBOYr0typ
w358TuVzHNME+YWcU+o4Yl7nW3F7TPYEYjOI0I9QxPHTJHC7NEMcAKFlbPfFmQnttmAbtUBe0JDQ
H+F9IIPf26p9qNrLA61/bbR1qAim0NGc4SvtIWOOSPu4LwnqTYEi6EQ/hje7nOnMGh/faWIPwKLE
EbdA+hlcHhDTyNzjlv+Wj7tuDLSPialur6t/Mx4OaTeXXLZFMGivEO23S3dl99M75+kK301uqXGq
9r+Tw9BJ32lyZs8q0EdNzou8ThKYKQ4Yv6u/1LalMPHAVmw3rD3L8y42Ox7yQKr5NrbFWXvgquGj
nxxivwOyJ2q8fdCo/gmA0OTvjG5N/5M0CR6/hPIMp2I0aRw0Su38WdBO3uQHuUxsMsyogcvuvuO/
v3aOvT271+62uQjzSTtfkljGRTExnr4eE3NsSCoVfBisNYiL2Ll3R7YaMJa03pdWLtUlChGJnU9G
ajyiJAuA4r8/iK8XN02ykkI0z0FvXmObGUuyCTeFo4nbLkD3GwCfKqOKyj4sicKO2sBKKscBvhJq
uKmti2xEZwF/vwGYq9wPiWWmz+1nF6sElbAj8YI4LE7TySj1A/WFPy3x5RntExh4IBSS417m1Z3D
cmI6Xvk1+hhGnEMvLXVnx3CI21HIgCGxAK6Ypug4p+xiqP7Wk+rFSDAXNFyEnqR5Z1KJFziOz0Rs
C0PlZ+hyx93ojhR65YZiPf78VrHKyGnZ7y8rdQg4rgyOw1RMA9xpk2/pOE9/Tr5g1WS3JaNvkTXv
7Vybj/SjVZhJULl+RqCaxAnbiANDfeEjeaW4KeAz2Sadj/8H+FjoArwUesnOCEz2GpaHIANVwYMP
0St0HO3AvsrCSpCzK6KiwPCftZfDbze7auRsP4Ka/IERNgF2QtJf7FmGpCw9ZXvow9FOurdA2gv5
Ky+4fcFbHnfBNsGwlQ5qfzBl6S3mm3Zosivf6zjMOkqymUMKhGcr0Qq2jx2TpBJ00htsGbAt6imo
sNOo7GRRapOT+hCi7s9VW1ZUhPCLTJFjhz0wojW8++WERqyziC2k50DC5tpKWZRWpyi8zC/QxpTz
PulsisJdkh11ksOSbyqhuk3Z7WomL3BFOIeIfYTYBxeqvJJfUyew5wBiHRq7Rp6Hw4Qy5wbvES2A
v1ILM4S/eBopaQxePbqqkPdyHQF5JHs77myKvi1r0dz/1JTN9Wnivhf6U0dYiqdKoqAposPhIHiu
uQ5vORVKpGg9g4hnaLzXzkWEwgoiCLrdHwG8qyz7L1DRRFSa2nWGdW7OY3/f1bA1eq/Y5n2nYu4T
xQsumGBpffP/YGpyoyKyWZYbCgjS3q+9i1YN4itfctOlGQivVqIsQmUGho8jQYD1wKEsF3nuQlj3
AqnBa17jpczVGZ5VVyyWsYrjlw5YjJTMeqBbtst1fFRReIJuCjbLTpOBu5TH0A18MeV21wuXoWgP
KLSUNqmQYm3m6XCfNgar+J9zm/Yf5te42aIrfoZsPAbD6Oz3dIfSZCSpIXPHebm6WXJaMal6vptq
O1iL0CrGaNDM9Y3u2CyV+vHcTZmVIkUtlz+bBTRt89096mDbsBx5NkS7RX6/cN0espGFaB0ml0Nt
JftuGvMMiW1leB3MC157TwhkZPMgAuv2mB0NeHDcEHq/rMOqahsHAIK9m6pSCEOH0W2ZSJOUHTOM
B8iNaBWGGwl6ZieE9ov6SNhDZd7JEwr7ZV6bvCsqybvLodcHkIunnsM9UtA1KOsB2rUd4lQ7+3Sx
ctAKAMkZue6qKwHZwNo8rsSx/E5mHKMvXL0Ge/DttyzyGpMjeHJnf14Ag0WhF5ckznZQookXV1LE
qYYGU6w19WPBmmq0Fw1WQZeof3gp5ifem153zV/oQajNvdhgo8QzBIq3adHverAJM++LayS+8eH7
19lbzej/yiHt8Bsp1Ji8tKBbgR36zg02pWC3CIDeaoJMCI2v49qH/SdjdtYR6d4Bjj2JVdVHaNLl
gyTKpsCginnTHSZA0luOA4WmpbruL1BMT0eMPtvjUavUSaD6LdkcC4eTOCynoyG3eVvVnrqBcBsF
25RMv8PA/l0RrXA5Unc3IZC+nLFOxKjvkN7aDxGXw16OybyBSCpWayT/Dh1RvDb6v01nhm1KP1mE
X5rslRqKmXJmaOVQZXeg6l+nIE1zuNtSkeAsvcmPvLh41f2W8qPwDa8e6glcfcR4bTawfR/kUwsO
U9iN94t0m0FU6k+uUEVczNknulhkqtlKHS2tcGtoCgcdiscuborkdAUnnMcRJJh1p+IBe3hqDT/L
LzzwtefUdgSNThoQesnwJ/AC84ZMzg2XJv1wQvG6Z8wyqWd1/Fi8DgkjLthqeifkmuviBD60JVRn
JG1rbDmjx2IFbPzhYjIINxzi603oawXadfkiDgDOft1oV+jPMeX84NY24aV8pywUgWyE6e/1cvyC
VekoSYNYtwGCyAB0iO2H+l5ITRrkqNP98d6c4+dxsBmGAT6WcKnPJGw1dPTX0mpEVWNcRi/ZPpQW
TnMIG2Jz441AKH8RlNQNQB+MNuhydzz00xKnvT3g+YhPHjTeQE5RM0iYuMIU+PTp/kMBDVrG9kBu
21PkttlXCGljsx9tfPC9K0x0ksL3bPZC25qm53GSDjYCxiH5AbvRGbqQrbB9yaoRwKMVdge74BLM
0KHrSTyoMX7fK90fgqQCmK7UkAOiWpFbuEfIoK6bXijvUfUlBOYAZgT3gfPnNtLIHh+w55myzchX
AOqut9KR6rUwEjOH6zj0mxwUWI7vFWKgQwETcGl6MdhYznt6LIwK58MRF9BzhRHGxigHaw/vnKFQ
wM2/dYW3ici9Lkz7SHtaD4F3PAUWBUXJ47nBlmtnrdu28kDu74eBY+JjoWRpqbT3h/J13FV57nZ8
dnM11Hg9Elvc8Dbk+VzPuGNL4ZVpT+XqRed0wloR1XDm+qVDoEPfRsUU4Vp6fGWaHq1Vm0kcRuOH
M3lAjoE8RJULKpmtUVZzysxOJmZf7lc/YhfKx3bUxA1mfAlE9tPznNsueCW8xy2qyHgok3OyqPg0
fYk/NoleHRdj9GHWe2ry+mRtqpr8HdTRkdTrittuHP0L+rcOALY+Wj4/D5m0Fa/wBAwX5cuRQm+h
72DnezNgGWO234b3duWwyxzEJGSDwiT4X7dWqG6uxn6/FK6kBQConOpaLXlpptUxrHQiUuRaFuSb
DMD845/roRlfV8rz1DtpZ6yUreO/qOAHxeN+bCm2iTJojAjIw1Oe5cZ9hXMVKI5+CUS9B3EkoWL0
psH1HNdJaIvGqZCbbKZO9tJEI/ZAK/odKtl7ntfhwiwae2jYJ1a5i8r5HjM0du10V4m88r/9AmlQ
QPRbcrSYoYsWfFxSJxwKeXJHf+eAdvdD4Iuo+c2iGN3vEIVZzc5/eZgtLSd+MIVGw/6F3Pu5e6y6
5OkiA0XHzBG3vmZcwPY3YxZpOEC66aqEMmcGPablknvJnpQEQ3scbAPmHjyEolo+8QsOm6VRjip/
tl2tHkGDGlUdW/lII3XlsHSTEXQ2NkdxROCsxxuTyYQqJf/AKaRQjb0ySDctT5Jz5mgutG9JRC4n
AqqSwNX52+46JBTWPJpcwwzdyOBt+1A6i4kJHRQ54ySkGLM2xAJUhJuyTZidBOQZyPYc4afIq+aQ
mvVr81BgPnvykqHQ0RNSinC7dV2IG8t6L4YkBc5KKqsIjDvDSZVugcRzm9lI3Nbus5FduI7CZs1+
cUJKH84NIi+NrgljA2x23yqZBhLZBn4f6GBASTNGNZUOCAba8oCCpHs4ztCXfZ6Vlswo+lLGaF59
Fdr4OrW4upLoTH1SJZzKhdHIug1QjlpsScC4MMZzrNC8FWKfeDGNKWNSVguc4ycvLnweJx57eFeD
XlwdEyMvSvz1dgko3xuRmOj7pU4eJ3nMI5nOritanWkmO8mLZpH4iEBQKwUqTg45NmCL+SBsPtd8
L76C+G98ojSJ924ImVNjXoD5FywR6WYdKll5Bs/UOXFD9RE5U7BVPNiq6qrgAlzMjApy9Yon1yho
PwAPAke9+2orp3vff3wzMSQTQRCjPgATSUlrVHCiCKkYCOvO4B5jM1WTFlWsfXZJP0kK1iBoghsw
O1iBTNMvsCpYl4YP88snckLrwf7vbbd16aTb9M1vfuVnom054QF9gev7ZfntHeapgD5IbJnmcf7U
WkjDDC4zqyPyHNI64CPEtsTTmTOfH9TTr8K3/4LVQvHDwXlJux/MmOK0lhCDjUm+D85a+d9rH189
Z0Vhr0qsvjbeH6YgLhlga8Xppj3e0GwoVSme2eIV1/9aAMr+mOdWDdOQ1AKWWQwTtqwJOfDO9exz
WpwnubzZax0mPZ/H+ZO29ujETnYVk/tIE6hdA2xRAmqjffL9kjOj26Y0nmg5jD5DCXXWY3mnoO4m
NK9N1VVDZqsBkAPBSJwx4P9F1FfU+6dRAmPvXirbHvvJMMsNHPylzO6lZw9he6VUhRVoXV3h4c4E
wdJLqsVoIux4DdpeNtu7iex9RrExKt4HQanRYrM/MPn0gtVxtP/3LFnoFiSJspdvsL2LiLtIT4TO
wSLiL8UVnkY9HGrNZoqDrXltLzu+1QBgGPfsZbMHrTKk7xCn1Db/a8BNXwaPuoXNfUqdzcPj83oX
MhwvkdYNnWQwWE+lWDNNNuwN5Px5oo2XC19rScSKe5/XT+Jc+ijggOtbeFBo99ztmnGLghgqy5M4
1XNeBOr2XV30lgz2+v81KcJNupSGQq9Z2rXBbDx6VGKPoMLWmcrtv+gts/5+8SeOfrDQtgNO+x9+
s7lS3hm55igQi73asqN0GGLufqhuG5CftQ2oBHN3FmWQzO9rC9swa8v+NE/lq7vys1o5Xpjiqrgq
ReBnGy2WqmXnb68zjxQJHdpdiY32U4XmdRorlEABrLmqvW4muShtwdXq5ZDSFKh6MO84+H69rHSn
AYgW/2vdjnhYsg1g/+xBTXLmL6gc7pkOHU+9+93K3z4O+90ghza4BC7AlVONxN46nYG42CGU6ElA
MaeVLf0PB8udh4kOHKzQdIX7TvOxpDVXozwXQWVmUt7B/5efHWyveWOy7P3sojhd11NTpSJcVAy0
+N/FwRDQslW7F9bD+o6C6oa8chuUbZfssxD9B9KjOTrZBt5Wn2ImD6EJjr19Q9U0evAcZ+mFUe2T
XHWzkliGItBiuXVLjoQszJBHuLrxzia0RcMcGIfLk3QXItszfzzWJ1htBajdLaBqbRsWzrCE9kzs
Y7x9YAASub3jU+kpJpyf3Y2zB5z50XD643cCKBxd5KS/89jsWa7rODwwYTI+Kv9ltu6qxsbNojMM
HEojdmvKD5kpvYIAcNO9oqHn38QUb4g6WOyka3nIvM3hzjEVX2DEso5O/RvWyMb2JVHEoLG8N5Ei
LiwAMmvzOwO7i9WrNYwp4eyjxqdKwVWBZV1GwuohycR8r6ATSVXGTwSAygtpYFyI+kbe5/ppyzeo
KsojjkQoO7rSyVMGIaX0hAHeO6bk5u/Ga2X/+dVxTYTQowguU/5Ji5TgUQu7yYgoxtMhkqzT+BIc
Rea5s6MM0Zx6KMlZNe94L8dZDeTbS2HpSVhi+I7imIaQkD2vbhm3PfsxYN2PZenu9hH54gnyp6fh
TlFVAwAZO2T5pyAPnpLLa6pJbz8JlQQmL7WaWQNvub7drQxC1DoUKoIg0P9NOZ9b5MmTmfuy0A/X
BogQD9KNzYjFERaxXOLUiCoU2OGr5i4Ti7KVCfAhzop8sLhW1Bkvs2JV0NTXE1NkPgFb9G5shmL9
HG3TgZHDoRKJGcqZqSZSMUzvJMg+/jfRZxLG8UQhlSsoY2eEOB5bpJe2B5ZNX6E9ZqvH/Zo7NhEP
de4/ugncORxr9rEkUxCP2Yn3WBFRwGpz6JFRUOzPF5m4TyKd4ybg13us9ycaCw4J34nC6atFUN5N
zPzXUYa5K4SB7d6UzK1qCLg7ZwQKFKgsExC8fub+VTy8nxcvvmR2o/OSh+JvMDZtrT0mbV62ivZu
hsRQ/+HWkPUPeWAMJZxfKVFfUcBgKUiyCffYwBcDMqhBSa1BpLgXY1GBHVBN+OV3PjlVSnlQKzzf
IcQ6Y8J1tVpbRiv/5+cg/kzEkYmRyh0hHl/LWfCIUYdkR5bONP7TMuPf9nUHMqqPkUB6xTjXy2fi
CY4FTAdDR2Hmww9ITr6/WcvzUtzihozEGEiaisuejpIqBv3LkNY4bm2s3GgWzl7dnKezLP5qY+ax
wao+OR1aBpzMM2qpWXTE6maXLniXhi/dAGl6xSEegQ1+/9eHS8p8q4Wuk9F1QXRQr+61kAG01MPq
gNRWTYwi3S+KzOgQKlTIJu5uvFS/pZD+O/9chpgGD1gt2OF+jGauqKNADtQa3b4Fp5W67fUHF0dg
JnfLXSI0/4QQjmNQ5npBXNBx1YnmEXi3igByWn9G6MiiQ3blF99z0dS/KKssr2CT2+M0K2aMj2TL
ipImQv1wcgqP5UDufTacuZEvaDVtIAZjWyViWQ16cqnyM8WC5/aaDAt7Tku3sjPWxHAnjKq0C/UK
CHaiRvRQdBZt/chD912Ve6FcakX6hwV1nIxce3WU3Tq0A8buUVliu1nJNzEBAaDNCtRfHlk3CsfX
cf+F0OVWcL2KY3Jnqt+hl8X9Jbm6ltImMtgpFlCP1+9s0QaCrnfTviwreV+J+DSdFOrHntC/XQIB
uwpMEcQCg5ZxdewwfUbM1PGsUwF1OO2uiVhOa3k9N8G1yKhfOGGm/nmDlyGNnb3SfuVKqh+gEZhn
jBNmT3AX2zY/9Vi6xpD13GxHSbt/1XIjGT+ywC2CpprEsh4uiWRi/a26hOuPdPvUVhIwA8Q3RhRb
e39ZqQpdNT3EFvEhA+9QVd252SQgXXd9xjM32aqQSQBwT9Cm+S3qXC/mwQ7FapocV7tpDf07NRZG
olN+RMzaQFhH9jxF54zz+o8+f/wBMNzSfYvHnRmO2MAt4AgoLmjPhDEdgcEU6ck7EDMSCN2ujF/G
uNpCfXyHq8WDRd1aWyC7w7AxWixrhXF+I7vqA4JMQKk8DYOxewhXsN6DGswWozGnQE1LYuJ04+2Q
SPGFFF/ekpeMQrCR142hKiISZxo2PhWQcsT7Q7Gko5RfIdprFKWOUvEoKiuWifNlDVe5fZ8fdK/B
B/by2oaFO9wBx9tYn2RhubaS1Sb0CL4+RcsDO8Xsidr/PxrMaGBXPS8m3KBGU6rhdVztbDxcnTEV
frWvS4Vz38mb8HEOl90VUxHHVIAVrqNjE3QIesf9KM5RMjMy7Fh6vWrZoLKfFVPMrjmPmx9w7Ky+
Zb3ta3GH2aYqLBxPPnrzn2sXYE6yJHXwrW9jXi1toZbDWoWFsSj/0l8fSdRrv68jkD/mtL6fHyMi
IVJ6nEBujowFvHztOZhbonpAqt0NcL+mOBPfx9PcFuTdWkXaHAe9T6W7K03cKsX3a5fcLaXMZfXB
9Yrjf/U4I5jbIz5oB8oSkN+iagTEWYRDsJVg6RihMQfwTANsrHYVNUf/JaTTpdAdev5Ggk28KW3J
92CETqLazUlffD/HOF1kL2BXl1C/b3O0F+zM9Yy6wyOXhUsFvJSyUBcxQpzxgOKnGVrvquaY30X+
XKlRKiFniDkIp1VYXHam8u/qOoBTmP07yRjqJVBZOKb9a15/Y9SodHpaNjac1oi5eWbFRex+FK2L
l6nmudsqZwmQ8FALWLAAX35vDi7gJoz3wx0C5xyaTdEyfu6l2eKEzIrWPZgMHLeemtdQM7FXzYlb
mVpn/blhiavURkLNZVHKvJ0YvLQg8T2X3MRbJF/RSEeZJ6Y+bz6YOIkNp9DpGNoesD1fYIh0lR6h
5E9gF27k8swmxlGwBrHFFwst5qLZqbHdXP+WEHRqTRWq93t5McLTmDfm6FfKCsIpO3qIul4qlI6v
LKJRLFagqIL0xlU9cFCQfmpTLiiAJGcGXh4+GUPqLvUHf1A75YgrdIz8G9/awQhh1W/7YOHWyE9t
S347RoXB0oX9mt5tK87fC9IBfIziLeiiY/c1Th+4Yo8DayXm6/bvKo8xhTAMo/b2YQzlfaoIhqDo
q26zJWwL9nBiDOogkvA5SNFQrjqtY7t8To9D5N2FQXughDhv0bORwEEkFXlb4esNsdxpoYOZgUQU
LCDRaeJeBcLr3Qcu/8NV+iBt9/fxus1B4qk3HPp8x1UH+lrcum+AZrZuaS5/UftAVWjoTr8gRdoq
tDCrC88VaDCtK2ssQ8zO+2CCrUt++ZbKqkb3uyxchMHVRKjlo0ZlGlF4yGvUGr6yPHImVBEk+/jy
bgRgzUvDPzBdQnTmPc/K7sCq4mmO9YF/QNMcsOjLUqZEM33z5EilukHTH6zcT3ly3zxcJNJf6A4i
QCu5J+mrrY2jNkOwSrMCcHQrXOZV7kYcEnMXrSSsJFKdM3eEw2N9nkiJOSQyKjjnYGhkIurPQV9Y
3RfFE5Rb2aUi4VzijfDkCU6UX1JKb7+gDUTies2/bA2fU+f8UQjTi+XkmlBA7ofeekp7eCsjUmKs
mKwZtA4T5QTFjVOh+ixzOwPo8SseCr8HK6UtFxrq1JAeGRzS0/WZAZ2z8p8RPLurQntfE8XjO9Qk
PsjnNlMtzcj803j1rN5eKRW5AXAzlGcwVs5qhpI2wG19IBXdwOa555jJ9zZuhSzST2kVVj09ODr1
R1KJumcglKZIKy7mzPWYjBS5SgLh5yLYwbDM+vaRbnxDHzmoa9/aTxR9/SqRpmhZeqWSO1qN3wqo
Is++Uq97II7wKkGDg6NodDXEuTOAapdLFF4voj1ND+XVzqUYR5eCXpcsyJYWmi3ETtgEMi/j1nPx
AyzkVTbopoBmQVFQNIt7wfDiP//M0yNkJTvWoDpuNzJnDWMqQAWVt4Y+6IF4H1jgrp099cgk7Hw5
xZ54Af1TOPuCtAiTlq25Pz+Kj1pGjvhfdm6+SOnCRkWcvdh5cPb8P+xGPJHA9RmS7fsPs1g7ZwW3
T6LEfvUQSmwWzIaq1Ei7MGNGAbu0IWbiSI60gi3u5GqINfKcjqmvXlaT6M0FfqmMIGNH3EMbvBBq
Mbyosihx7WZ6djiSKCHVcO7XS62u5/23lxvVDZkCqlPhx51Z0qu/odTWnZW80ttGABULDyTRB5OW
4ZjmRYM1qwgQAdu12+uCwChrnuxREkzWDx2FQFF1MIrfapCq7L83gPm7AZ9pHqQ5zkzjcHPiJu6d
Kz4bNwgk0CdNzMsTdjDWpNUbgpuAnDxYIiFWQBA4TScVkseZrNbZUOc0FE/RoPkLELF3levsrtjy
xjLxVi+f1w45rA+dnvuLRxPG4iTOPAQvIujhBX4vnzleLRhSY4DQZbQbgDrRGRumw1nA+1uek6xo
DnXRQLrXrxJGsrLx+AU+sVs0bok4+vQNeWfWbXzwIwoC6IYD0DNl9eymuIYtEVZDFKOf1dRTwCEv
mGbAc8iiA0YBlbUrXKEGO49c6luwYPV6HDosEm27p7Vq+IQDJhcuj73PvbwyuokIdsqx3idpH0ut
UeN1Nmc8qLIBEPvd4HbpX6zkIrmU9RfC93Dxw/73sb5J9zBpsZ+ILSeUDcD56EGSA2rYoiJSHlty
673MsvQmSF0M2rYRkvRA6ll3nlVN91pYdrwLLN2uo566KH/VKZXSJFXBqiUAaDhdOOk4/kBR7KD2
MvdUlef6a5IsWM0pfcP9js0VUhRrRe//xoubB+hIwn1mK3+P4CHul0a/OUJF4ZX6D6qxznkUOpmU
yBwFiM5cUcKgPFHrXWHhgmVe0bRMDUxdoiFDzI2rO9JaO29WnY1lRwn074EIE8HlrPyC8FtB5jYW
ILOsisQV7RvDO89Q5QU4qGmfLAUWuS+gmT47PUgmdaM7pUqaZsMsXk1f7r9UElMFeRnSXfg1NkET
nF54a1rOp/RpQc1Ok7HBpvzYULZ/JF/oBfIb5zG3jq07QHco+9eTMG+Z2z+Y/pVys+zTm8uJ1V5K
jA7TuXjK4z6a447NVnwwWdUuj0wf2Piu/SDzf3XLH8fQcEn/brl9w+t7Uug10W11KpeRNyShLALt
1pBWCrWRuxQUCObu9QKNOU2nl2dT4b9sIPMsT03dc29VeTKe+O8Fh76zp1QQN96rZfzqhddMxSSQ
wh3ZMsgaNMMVC3ZXyO+w4oR8hFUEruUqfJLoAD4a8zYoFTgrTR6EGnC3UAhZS/F8KqWl3A5r0mho
FtryCDrrlQqeoi3JuAOc3aJ3jlWWa+l+4mHeweFcXJBv2FiCl0GuIAPtuBTo4go6hiV7R7i3EVr7
gzwKc6mMqcWcxSjVj6cFG4C6Yg8OtnIi/SZihyGkCqeHk1HsRwQzMUlcTAzNd1U0F6ZIlaDUFbqV
UTz9ujiQuUfGqORqxJ710BfWSjuAoOOucF0HE6VVkV0oXemkziDbPhlGcV876GonwtJy/QlzI+CI
eSHJ18Mu0IlyvKIz2L1/ujjCQ2UmDzjpJW0OWqy1GQnDc+bYBRfX3fWOEIAp3afFFaFWj18OF/Bz
pZK88m/xfpMKyL4cnh4puWiGP9iqqDMbWjzR4c0ZnOZ/A90aQzsplHIR0IN2tv54mfJClwDaXu0M
zNhCR4wH7j+SvEf6QXEV8fywAXwfA4uVKVR5ZtmSzmw+22Ayw4DY+aEaI+igQxPtV/XwtJ2rsj2L
AzX+dVMfDW5v1sUKifZwGmKUIRPaGzoLWWZyOiE+12fy5rtv2M+4/KaNWgsWBhM3UUn9xwRnH88B
8lWcjpc1d9DPv+PGzfWlZhT6xEVHl1mXHBb9rDBCLS2SpH5FU64lnyYRcovx19k3jtneYbAVyky4
CFVvDnq10OmQNU6hk+uPwAM45eOr9FY1J7puXN59zKd6UYGABl5Lhs2m82K60VuTKpY8xwU8xFPS
nXzGXhyc4O4VaZzsqabwHU+6yB91iFli0KlOjyzCoDxu3xs7dyPl5v8P90A+e6Z8BG0cIoPxiFvN
EY2gyItiNaEFkXAK7v7gpuoq0yFA3BJzqPKX0knZnRzhh00QB58FB4BKmnkuf4GiHVOL0m8sjfCm
YitMwPowaRvYxfQbhqxaXStv1ROzriBvT01G2jQkORirIbKH/sN/E+4hAsjKpGPnq8eIwxnms0AB
wUflKDAESWh4D/gMs0RSZn50T1+SW8+s+h/uNF6Nm8PUcelJQ3yzGDRGvuZlRsvOHRfpEastD3Li
F0u+/MQo7rNhW/90LFgFVy7OwL0XJmuFce/ncg0kOFbZTikrlI0YSd00h7v62WS2+ITC3zgslNoU
Gc8YrAMLoBcPnaOnQ/s6UiJ9AyLnmNZoOarptgWutUgxORXy7fuC9MwGahmBOG8vYvRoze8FHvLu
O4zbOSlJLmqgKfFK6lu8daNAriJShUBFptc9GWAZFXU1L/i8UsFhhiu9haR7nS5BYwTb3O1jQ7lL
HYrRPF6wnVDBnsKfBcG1+xNiXIWtt11ft1DYqsBGtLIPzmE3BDrVnmdKkKQfI3UEyYF6NB0gLLV/
RB1oCRo2fYXZr1F8MtSu66V7yV7weWX1rRlPJWkQ5DzseuJo/tQXFDFXX0BZ0Z+NxaM/4Xecmn8T
U5CXRu8zAzJwVqPcHoCvDdwrhYfObnpWYSu6GUwz15HOJsViXHq6YKSMse5m0DZbtNA4eAnruAYP
BbqgYMttrE4HoljbbHga4UZL27jugsO0Nl2JcASgXURaKIm47izvH8/Ds9r+4YZnMtzf5IqE0MbK
kp8WlqbLhKzqLdUDcdEZpXwM7e0DK0A4Pp0Ia3Hgbe1JQ3MxYS4WZIeXIPoSWicqDmdqN+mhrd8v
rNDUEU3gFUrCUKTyeafj/9V+6wh/kQKc/qgTm+EBiArKVRPgY0sgyD5U6TLHRJ7AYS+BhKwkopwq
JIvp/cob/oEJs2IknWKlpBYkrtIQxhfWQ4U3rLdxrmD93D3nhbPIq6d7i1kUC34nx/DAxW9zS35q
YCT4oa1a1xAQc2MO1YDcYr/pN/ZO5KpmqrDOTcoVwDwU/S6hAKqwc05GRd9KG7Yj4XcT7fG1frwe
XCx456jutZvcaDfYttm3rTyqKYzvL+TRqCML2XKaf2BgxPM7Y+R1ddiO9HJzKk4yqvl6bMsugDp6
zPxO5gCMzNM2uR8nwHhnsNd5oiIBkxTQHjrQvNUyNGAuchpm3Eic1wXoV4hjvORb3nv3XqNgEX9t
w10qKC570gAWrXBjBiPobHwiswYl7ajBHB9f2PiKLpoP/KdPV8/oKOfPxcLUeJU6utJErhCTVKUj
v1xc1y5VAHJ3hqe8CUv3EtcIFfD21Yu+YX1DCHm2z5lwPgJDTxcFeNHUP6e6wJoATIxPPIome3Qe
lr5wVF88CisKwBRLZLqvjucM+63tRRxm+t9iEm30GsRBvt/xBarDqzkU/9fsTPsakjkOiIHUUmLd
uMi2lWOpqcdcslMbNe4NJekprNdWvfrMnZAAy9CYE3GLBci7cqiC2vwqlWU7gjty/TYDI6eTJ0UM
Wmd1a6t2TCiRxT7d43l5d7JxViMFH98jTtXxB+lc8AFkMdzKdWv1HwxK5/OQLjI0ejhAMl+7F0GB
sxBSPpCIzdtb4gCWcIupyTkre4cxYLjvanLJyxkqFg0OZwahIdDXw5a/xxmkNQXbq5k3lwqoxyy4
RXIYpfqUDE1s4yTYZ/BvgdYjr+b4Y2WD9JiQ9YzT6+gZz3tWzm3J5Lrep5BRR2SzR9azzb7+Hk3e
Zr6HQMImH3zq8Fw7JXf9+JmgOTWVO5tQ7cII2mGsTCqN39ttLxeN/fsv+CEtl8MiyyJOtBtUGSkr
YpMJnvsKma0GHmiRuruU9H+w6Hg87IBrIfHCMPPe/X5sLwIno1v++KoiM0ZlvtRJJHRrVSOpgGmp
BFN0c2k8k2lRhZirBy68BzkRCEkOuAm3GYV8Q2Rm64RqLar5iDIL0JysDjAILRyO22d2GfuhWEMo
4bJDzXL0eDT2W5Cwh9VhtR1dy26qTsk768ZJo2sLsEJbp5wQ9hewn4oy9QX2vn0b3+g/0NqbXgZz
au+EFoG3RBNnr71AiUt16QZdK1f9+itjuRmikvc/LplIqJIVi+geTOf5uIoS09IntLE2kErC2F3i
k6+0KgrVAomSwsV21sABX3nRm1AVzh7s5fOmUymvRWaXdBwajiYjqGCobYofF6g6boapn4wg7PTq
TNPF/wXCj1hD04NsIJ4KlqNJRJI7S+k8l7tUytcHzLtq2qN9WuAtp+6vyiGjpm+Y6XNFZf1xk2Vp
gHLYoaVgSFQqSf6Qy/kHNDOkfXFWWgnnkr2gAgnXzwqiMWd2Nm5I/MrItt/oagjnd2Dzp1WKOzbY
qJ6pvbXY7v6G3RdT/L4HB5cmDQtR9C0FkPBE44t13QcYZNA6eL763E93Or1ZMYA1TNBeX8vWsm+r
gytx9x1eNA5hnBFZEGIXC2lGoaGNiXe0o15uZOK9xvocw2d6u9gm/KzzGby7O2c+BTJnXHpiIAul
BZD8wP/fIrNXemFmBmy4hYvhaju3qlcpHCkrMlAFVTeV+vg1CaRRVKH8gYvTgLayG7NaExvS7SMb
011BZQU+ImEmjuPHQS4Xmpm07mXxbb9gZGLwCD38inXxSZWKJtdOQsbwVlsg+N0fvqNHNtPhGvtD
k9Nn5nB+gCNEXvh1Fq1b0RuGdU3QxezDJHj+b2cUlqMJvyDDZ2BW3BGkA+CTjmDVi55cHD/ynnDe
nfBCrWmrsmBqdPMnJne7aECTOsSo72VjzDhyXcgDjkQe+rOZbxB32ucLCOyyukMPMMxiIxkxc3yE
aXexrcPEWcQyrWYB8K1oN7wTE5CEVsYmCj8F2oFPeMoosIv+TMuFcr0SwWMAR7sb1WnwCB181XLA
c7c63gkE/TdpPrBqjdDi6u0qyzLZ7NJRSHK1hXRhEdszduEd80O1mDHmxk4V8Gb94sV+L0WTFNDT
hYNEJRGeqHetNpe8NOewnQjj+0h8xn/g26NYSUew8hwyalM40r2T8/5On9jWTF4+evh8QIqTfVck
VUzaC9tPgH7RmkKw4WNC41ynKl7TXTCubWvCJ2dgB28UDmtWbdu1wCEfIczhFaA/qgK7R5LGYVcf
y/MU+e2FXNosgFj80bjwA/XkCWw5BLHENH1cYfcY1uDI2WdEZL41qbZq12X5uDQ6zEPOqjcAYi1l
/HKCdf5WAcJF8XmUJgWYRzveVKl6NE0SM/suExv5B0aNTzfpJ7ur0my+HJ7RPQsEiWE7uVivzZuj
jpkRchK58JiPC4DskagK4vBK5xkibdPWsdxA5+wZqY8ZuMegSXQUeL11Fhz0WFbg+BrvK/5IL04+
hpywuBjHcmUPD4JCzoWaITD5T2KYu8l4bgTibUpr6OSL09b61eoi9lOYh2JBsJJPUy7Fla/IU014
6Z0dRThYAATu9Hn1e0LNdMVqHVSbiQVp8SVDSGgxgLH55cvqlgb5umCNhdZt7H53BbY/+KMVNPTh
6hMWG8L+FrZzFKwSDZEJoMHIz+tMJJXz20XH+JINw4LYdbr5km8TnwYGPuBiNNRxVZCcRnihW2sZ
9NwMwI7k2VO7Kfj4rY2aO1qQRCipK6PLkzyAwesCh2BcPlCjoK+V0G1hBUdO8HSrgstNrF7xyiIT
40CJJQewZJnHZKSWAAk265M+S2Jn8NiGzrCmTvdzq1Fl3h169ih1y9uqKCc2Wck+f6fu6KPmoHZY
dpFvnntnQi7XToK6CaADI2chfoPv5GDbtwpN6VixuiWMa9YFJTMXheRorRRH/6EEc1CO05iMEz1j
kfIkfecb8ncNbIMzDNaIZqERfYQHI2jIXKUygPYby/2XeijInqF2ZTKefM02dcNsezGSgzGz30I1
DKYEUMNa4XrRTDuIgG6yOt6BWCLJwxDXDdAiuYc1GnaeyVfiKsxJYie5RAb2s+NkGi/WRFcUgKhU
ArUim4sCNvmKGbLq/YpDTF3FDEtxiKUjcLUOYN3Mcs4EIGfbDSwOlAhbTgewbF3z/NiO5tclhhU/
ahGvUObzXaR0WZaLgv8rYxFngq9+QYk/tSKQ0UFuBTbBbDPBasC1tBjhJtxIW4bMiLYp0z8K9Yr3
qAJNF6k9ZT6chHtagGEWgcUTqCEjUbCyg52j7MLuVm5PoyAnwiYHddPjFFF9WN/8N0tfN0TBF47n
hBLH4pEJ4ZikevUUqM2DOf0gW1JIbC/T3EWUa2PikryF+Bdwptr/VFIBFC2IoS5Imk68mXx7DgCk
wkmpA7QH12R59CNiYFwdW6qXssFkFoGhxI7qTNtJhgdxPQLkTwPtac7wsUCmTz2Rvu0TESr+Ll3H
FEcrCmgfuC9lNU05+8EssZ0hNeOHoVCy9lFIN1QWhzDOM/kAfaZzLNmu7GOJ53I6aDnC2ZLAHtvo
VHehx1FklQQRz9d0Ip1uU4cAUhdb+uARRrluXDuhNCkR8mcc+gSnVaHHcweilu8oKzV9y71ofcjV
2TvqROTEXkkRmbAuvnKdLSg8UpkgradsljjLeJf8Ju3qChDSR22jv5/R2rX5iwP3xCG6Kj9qEhXW
6viJ69R6fAsNlidLlMvNbwf+bBbfihSC8Jx67TfNiv1Gm/bdqN3U/mBWQrlClkIlemlDY3uKAsWc
St6aFjntD4mo0zIWwhLaJv/JgMF1A8YxSd9RM2b70+ITm/lJYAg3LQjY6Y4nKd5iL28p+acbA826
bmUklPTriQ37jKdQ9PQY9tv5Q7+XAaWSgzRL6CUGTLCSiL5gw89ZD6qXFAxT5EBQZ4DdmOwHJ1jV
88e0L4E8CgMqlchB2dCGa3nCuITe6W8yBjyYrK0aB0KfNXSA8YuU58Wcvayh13vH9bbkJjCgpL60
dzOwBo1Sf+FVn0gE6fGGYJULu2xfopYsdbVozc+X3PRWdtl51MueYbNgpD/SiclN+MdBsAbLYtaI
onYEj0yNJTL+lZ0J+QUtmbgFmHCSldtyKhEGM6ZIVaf5K85yRGAyBrlrnXlmzKq0PA1EgA49au/T
SnvdhA9jAdjTCPwZM3d5SrA8qLhu2fH9EBPl5UXyjCQSZhIMcoJDo5p0ArVlP5+IY227hLv6Zm+7
HhrT8PRia1pukBSWqOBRDnFSCOXcpZLytK87FAht6IyS/DnV6itT3m23QeXeX/QOjX9eUH4xAmmT
qJdsyJooK5dQovt0W8rI3nvkemTAM/AhrzbULayOaAC0zSdHTrx5QwzGEh2TAV2BXOWEapCSg6l+
GJvb5aZq+3O+X7+vQS8xPdyxwcB8QRfBA4U0K5DVtHL7Uh8KEP8QbyeabG3uVwmWynoS6d640Eg6
s3LuR8hmhzBZG5qqWpLGW7kTJrj0h5ni8WXwDyQGKf39iP89Pcu+2LyAE+H5F63K8oZfwUvwNN0z
sHwcv/kFxH5Zhv+UbEEjysYJ3nQBoNcEvpfmadhqLGFYWlz5ridQxjerCYsP6ja4wKdYMycnoqHn
gCUa9/KHDlWt6HWX2+Bc+JZ7nsiRlUdJpQ6ZNejROATgR3UUlM+1s8odIkoovZfGczZ9dsL6P357
NvS4AS1DK/j1+51nVfYDudv+cR0njUPX3HHr3gh7surfYkj7/wBZclD3nEwp9+UUI48fEDm/1FK2
XG9HEbhyWR2PUlPuzrnb2KMOcHIozpQtBH0MjtuII3VocC8rrhE/8M0ordEaOERzoMLUMpUOZWJJ
GNsAWRCcluIK2DKZ5+ihCYrG4RZF8pbCh31XHG3bjjKkQM1RPZjZuZ7N2Gg1La7P77wbLyK2PL+3
xA7S8FOoWR4hWkwN1Iu+IDApayabealRX39oJao8jjGrwxF7F3SkuiAKLQnXE+eODuuWmI3nUupq
r9GpV+b4KhR+xggyl9MnonvERc3GllI8SDkQqaeIjDFP2WshCHggkS3VPaJY2AmfoSBOvgA7Sx7j
4I2QKaBejP+jR2ONwUSpkxeJTqIyCKy8mwRAGrQtGkHVlnxuPuqSUJu68/W75wihThqZtNVwl731
KcKx++wiSB193OeXPfXji5tSnVDMTLkVnsh95qcghVrmgB4/Z/sW1WLfL+xx7M0rkFgH4x9vqEN+
K+ldtlcuiIgVDRfzdkn5BzGZ1J2TS4gvnaij+ALAm8UO1+IMHsDL+b5oYPCbd8n0HRb7tdorCqRf
OddEpojNAlLk1fpjQWHWkYP+E/aZo2IcIM8ductKZFHfHL/GrGD5pPN3ixv3hfa3UY37YjpIvNvR
x/k8vzkCP1UqhS6VGB/5SfdJl7XckCxsUzzco3ThyNtqeQ/qArILlOzJRGlSFhRLSYK+Fb4WVGaD
UWP/OeMLiJu1/ArpUhCQoqY+Zgq8onxkHpHzbzbVx+ChFHaIVgbALfiRZG3F0O0zATvWfkQ7Bhee
/WULyAteuGlN1E35jSt50pVQ7fDmAxtuPvCxKzhrIyP8axPwSiEMaV9uG6Nr1JNVVzhYyK6S1Ed0
KGlY6dRfXgxwCoeAIZbr2hmr3MvxI/s/93yGK5LXT2sgpEb4Y4dnb3OVUnJ+V8HVaG1+Sib0CjPS
3bJKhcam1w8UqUaQgDNW0276P1LlhzYxfzBGx1v9qBh4WUOPgXwf4ruyMZ5kz986uhVM99lKNOYH
R1JRGr2B3IOCF/ThmnxNuH1MVQDaeSABssoWgYKKtIX5XCOTvOV2Mg0W2lpU0+xrCj8UDQmvjehJ
m9ihiqh6oKmwQ3kr1uefUX6IW5vj2z/2RDNnj1RVKchY85M9St21UvwCYGlkv/5biqgMoWh68msg
waNLWSVjubs+F3Q0ZZ5UYvD2oyDR5hGoHWwcB5OWZsnJfWuyrkWcUJ7K2MRLVPpJw4NbCjHhcpLc
dgg2mO0mZdY00AQgfmXxOUnxOfXgRKQQuzrRzowu7OmNMmvYNPhTtABofij9PEm4rbq2KXxtMrzK
SMEeutvEf41ZV+4NHJG1i4Nvd+Kz+WoRt0hLJPnMcK0BX/D9OSi44sZTb1nhV2wsKcuS/eDNiUtG
cgLqd6dZFvtWcJFJcELvhXK/Iq+MLnc7+M84iSArtzbtjLwlaCrLbrOe5dTVfgWADHJOsZumR7kZ
k4jLT7qTCHZqEYT2+qmBW8VEZLjamC29n9MegeQcBLKK+ZSE/IP9iE4caWzDYMlxy9q4VlnjiXSP
V55kF3JgBOx+fyVSqqVu4Fk4dpk8pAN1WgkBhLL3/j3cAIm1/W4o0usF9Fizzm4QVOKhGmx4TKe3
ukacn7vI0yujDNS6J7d+pPtibHK8X0Mu6eGhITNWziE/unl32f8OGz6ij1ulVCjNHHlnE0OzFl9K
ONFIk+Rp/geagQE9Nk5wfSR/ay5R4TA+zxT/QJUQdYMOcm2Xsc2UnnFHS4mNv0+KWghraW7KfA78
pwK01dJLCJqaznqR8DHhhkvvy/ukqi/7in8bIwULuhkjKPBWqmt48MqlHMt0KDAAq82r7SeigRrl
KCV45YggPH2/uH5MU5ak65JtwmemLKP4SGq4BjozeFrQCZDKEn5uq5Clx660AuOfctuwNxYl2wFq
xGZLET/9GZdgiSU+SYms2yUI3uv5d/Yp7YFymPUpDGbNPziE65JJPXg/J+aPSUwXAmakGBrs7/CP
ertrBjMH1yPWfMyOAuE0EXvrxLWjXYh/dtA91lt9tgfJgpz8KhNKtx+XMMUowqua48zmBunz2XQK
8DPpntd1Bvfd9qrKd2CQdC9/Q25n7VMX+/f5hZsQLjs74c3IsGVixTsLwfIrLPqCBxTwbpJK2ALz
G2269RM98MYxYEWn78ujbv3lzWyj7CB7MeBamJJOP/9AFFuMJkEDsEMeFqCGgybz2f/DugozWhNy
BlzS7983kmQkk4cxvIx8VYP02vZJDY4m5QtDQDXZRmwTUJPiznIXiCB81zClLJSTAKGo4MHUncdE
pVBnWgnwM5bWo9f3pWq0MYL7bcAUggxaTHu6pDHOstm6bHj3GVY39CJdfA+3019CcoggbkmvTVpb
5ziWkJi5aHHcvV8RGofQ0sMa3L4tgvNXRH+BaGeNwRMstPQaDoedsSpjnrGj+IbjKOGvFgR6gCcA
ne4tYGMFINJXcPPfSZ/crs1q6TO/VO75li97IIdTZoCup7ZnuDm/NyrBDRkMbmqD6fBaGqP6tKVG
BS7Vk3TIThg5Na2sUyLbME7vZOo36KTO56QUYAVXk3DwlkrS2+rK02HVy6LwpiBc3kVIQd9yNBjY
26WrBnCKAoxlHBi4I135PJe889w/SkRyl3kqMHjpYA0cKoYPjOoE+uydKlVh3WogEa77UJh83TvK
6U8+qfxcFykC2LgYO3FtF8cdWac4zojOi4RE7NxaJ3Vjlaunye5EbX9NYcAvUzYxK9o4SXNLhxad
v7tbW0FWiYtZinfhd1M+sPwBZtQVMaJH8A77TEGM2I/HghEt9BqK0YqJFJRaKi6ouBVVSPqHTWf/
oVkrh6W5CuRU8lcP7s1SFrYSd2gH20EQtjNnTuVs2EwczYqLI4x8u1Fd+29UrhrLBLxOOp5u3bbB
dCNCV8UrDL3igW5gVy33HV4zZzB5ntZjzwlQhDKa0qFSO2O4xIS8+h/lhgdhRrPBPr+Nk2uoLas+
1+W4sRPAx0L4LCOkAG9z0exZ4slUOf+yt7IhT/Qw7wIgLBNkncI/1zlVBtzgSGtDq0aG7hMGNaFd
OEdrmtLNPewQx9U3GAyCzxPZk0VLntCOdf8DgjddTLCxq5LG2bYPcgg7NFBuP0EObFuoUw4GhtOW
QxoWybieQbRpL1A1goMQolA3lervyJwuqUG8Etbu7aGFXkmY8gY6n5xvQDIMc3aRaTd+1MDqVSz5
USeV/P5YJXbkYGtfJPpw5rfAflehSg3X7Ore3xyxpCsYFQ8COOkn39LvuOXxSDJAQxJH4NuN9RaE
cr8ONdrtRDB57Ot5zp33BV4vC45Tz/1pspq/F+sgxz0nt2nyAYMer0ibOqkbS/0d0vSmjtsB/Kcq
+Tp9b6BPjWH0MJH6LvHUcLi4rkt5aZLjWsNH32KY4ZPhDt4hfeskxgGmahl0gsI8WcKFBtas5xz7
FKXpxQG5pfHDYFzq6bV16a+eLthVsa40BDETrDnYQ1uSREEViZLtWNy1zLoVPreAcdGqQISfaO6z
vpVk3iY0JLhfuY9DUOkgbDwe+abYW9+7qspWmJdEn8TH9lv0EQui+zmTaEF88t9YTlIdiMYk+WML
iEc1Pcfu7GgIUgJOzCIa19HSROGFCp1REmWt0ibAXVuuA4ZC4K8jFlV85QAsZcH2CTgK5mYvWWPF
aDdJ5f1eY/uQJosSZUTP/LWQIV60Zj1VjMAHK0V8K2mERZVKketxUr9+I7yaZ5OWa6UivAfZFe/w
Zxu6WVTnXBKsC6Q0guUuNMVZFe+1l+XYKldwO2yHn4PMjXhn0NBa2CdIabm5OjRMNy+WsFIGzACt
HFsPcwnykARGWSa/aaAk1K0Vwy5voojUHzhyUhfTeleWZ4JcNd8+bCKWiDLaVgukZ0ks9Y7e3D0x
CYSUVHyS9DRJEJtzzu9mN1U56xZFLGMpgTJhmpYrT6V+/aQIkVOkZKd7Ah/4v+2LSqc6gQ44NLdU
VoHlDBZnCcW/LvSvN+mNTOe+uvaEX5nyvRIdo2eai9BpT41RGrbiH8HLGji3a4QDe67fieFgqSFl
0ohneF5dopIJ7q7XZ2wzDZ3Rmc9yba8L6OZni1FjMj0nTvn0QaVINKJXXP1QQaeCd9HhFhbEanwa
IHGXsqSV6plBg54ImIsOXqKFGGgoh/yza0DXUBX1vZntRmEaI9yIaRNp9QunzdRaN3RtnQYr9mZI
OOuiiiXBXukqfq+TihHhMLv9A5fo50VdVIP4hjDrRcnYphSBUpOVPl4TOce0vKuVBdLJVvRfC5Bz
PV1DDO/5iBVd+N3CQJFPp+4fkDrwx/Cq+vX3dNAVYO3AojU/KupNTNnup2ewdU2XG5/ojbvNJfnF
6LL1P8qFVnklEXIWeDDLJfVkZXhsAmgcQXDVEIZrb3QncOoivCXnDt5Zk0uCqmjui84dD3UjODRm
/P2lzf+iFVtp1IOeM+gkheIVAiFIUTFWg2mxBioS9jc20072xINGy/7BLel6ygZXl4xmRdNSNmEl
K/nX3AiNgIp0pxlGNQnD7Q6UOQPZdgGcMhxQW/IM/2KC5KDs7MNy6RDfBGEJPzTZJrAfvxXEjQ3n
M83dnhCqjwiD+xpYawtTqxKUoXJxXtaaMfFrbh59knyQQ14BFD9rZHXo353Pz7/jKN3mygYy+Qzh
GVnU5cB+9LqcdeJplP1EWc18Winf8MQZrgpW/Acm+t0gD03wMXUnU19Ftv3ShuRSKhY4BcK6vh5g
sDOPyRJdJd6QgyA0Oq29mYtUJS1ekMfFMZaLSi8KdbZDFMQQOBuzhI+RQl3CzhL7lBvaymJQASt1
CVfYPm2Hugu9uDaqE1j//IbrSqjP9LAODvceil3dpgdFVrc+2c5Xv79JAlqZ0AHB2BFeW7LC1HBi
LVyZdnLCP7Ady/0+k59qcYMvMUzdZv/Kg8lE3VP6ixLenqjs3xWOv/HqNB+l+7cKVHf42MyfTZiP
ztmYTeMEsEQsSa73YD8i+e21XFyXcuRDXIy/JIUQ8c+EzYjJC1f/jGyvG1eOplz42E2/d9R8EBpc
43Y4bQDNiXrOWtiX6HgME5faHd7Yi2iuNjYIKw4lJ3Vfh0IK1rAfVNz/mKEd74o5LrvwFJSBbj3g
Vme0Df4/mBGcWdyqCij7v9V7u0Kt0Ro38GIIwQ9HVuA8CPeyBIL9qg3I/cGky0dowXmWWePUmr8R
gnLh6lwIFDhh/pLQc5rVHUAv8pTP/LAsmbU9Rks6+VXd38+dkJBNLe2emjIhDs1n8GjdugnXWdCB
aq4V/KCUdLJUSKivK0PMC0O6XX9Ki1oAIVY6MWLlLI5dJK+g71S1AvH93Njun8LxlP5wc5ADIwtn
6vkPvdTGaw5inEXn1jOr0GcXmx8RYFAjCTT4f+0e7VHhyLEoF2FebDKSL0b+bsYeHldcoBoV8sl9
ZLfD3xazj/jumWdZcdyZ+SzKVTvhgFxd88ZkgC/hbcI3OYeZsfVD+cqkj9qgDRnGPWu3d4u7gfDR
/Ql+EMCINi5LeJDBRke1lJPfophF0k01nkFAk1RBQ2L3Bw2Bb+XWT7bZ4dgxDnnlzxfq4ZzDnI+i
QXpDx3XWOq6K5c2uVU7RGUBDIbuwUGJoR74eIxEjJ9C7QcYdosWg7hXBCnBypECrJpHZtDqOrbaz
Hb5AUwngqVPIBgcQLEUQ0kjgQy53NE8f7kbR2BSor5c3shphGjmA/W+omq5vzwvSQeAe6hKcMcaF
1XGcGidXwpLk4AwXJ06tFBQNcBa0RRl3bnizv2neoI8VifjgHslXjLvNAnT4lyVH+tlyZ2VEbVlm
m7ZeS2JBkHH2svSs37mKGG9F/nVrJUNEKemP97QnWvbBehN1pwffzzU8rnjE0eGKnTTddBN5Fa+6
j4tuZTUv+NCaCgSaCawtb0nE12co9CfC1c5dtpZt9CWN04xNyWYf9xVeqYm7uTQntVKttCvqop27
cq5eqsq0p33IuA4oeDQuFjZtzFBdz+sdZ7FCR5Ut78TTQYbaBCZsN70V6RQkcRB5d25DUNBgV3fe
XCJikZX3QmBSep96lwpEF7N/QU8gBsyOQzVhAvOnyUvjtst09wFfUTh7o40ctkJRhsFnWNX2i03D
q6pjCGQglr3DZ2MJbGFIvPAk+fcIIwCaPPs4lLe1wpXtlGI4ztWEi6cI/NEys2KcqqlrR+f6iLOl
pYVH6fulPlkz1Ddt1IL2aLMskjaibAKXbcay7mAZpRFMfRbFoJ/3zVW3vr2sMkelIajdq/jTAkfA
L2PA9dlmGHJHGxV84xuVaNxNH9oBvzoMP7Nxo4b6KdT+3YF97Kien62CQqbOPmMpTNqt+FIkgH+X
JxS/D6N29vUp/j7c6ZSr56S5/WJcR2E8Bb7vK5DYwDJH9uBgL2FIYLmg4DzQ639+AWKEbKeYKKdx
qZJK9/g5Ssng6KFMdccRA1ARU90Db1vtX83XH23ipZeX88ANbWnmT76cxmuek8MxzI77cTv1MI1e
oie1y0Fpa2egc6B68ln7msHPjMjFlZadOcLmBVh3J8mMUslIwhFivfTjBXEDSp3WYsSgYj6ye91/
ghKyt1BlsWJj0e2W2pt+wC1m9q61C3PoPtMoz41xPibc3SOuwTJpUzv94SQyXL6ydkzhTvCkS1Zo
97gJlY3ouye0AixhZA9JZtJCSdA6OM4NYUS/qRdq6xy3skP5+c1tSpasRhqJNdvRn+SOQ5zd03aZ
s5bwffYZMfJ5qcfWrCta4/U8q+l9QzuDFItluCfOBTFtqVxDQOapPXCh4AQfztr0sT7Nw4qp/pD7
hGl3LXylcsG38WpdL9u85ef6D2Eqi4azaZqQRzYnbBq0hXMKaRZFWLPn9WhYVcxYDXIPunihc0zV
Pr7azb7ClG1amKx38CQKV3s23lcfglnl2TE5t+fBVdLSpS3wNzysMYBbNXKD6AZxXXHWYqy+Vtrw
YbmY012r5J4QmMIUZgMZJs3g64+16OtfWwuKkV45wK5UfjaoEfdUHfq61fThdMreWy3ApwsJ2LE/
M9bjyeJMLTW65risluGs6YA06WmVxRLeA2WHuX7Na+FFxQDYK/6Vagr8cHwyMKnGkgWSd5pubcx4
g86VgRUvFk+j2MLuXa3y0/dREMUWyrDY27LLO9x8/FKAJoHmggCmZMr8XWK0XMnTgTsQs/oKzTva
L1AzqnaBi5u/Wm40RUNheynxFXzyq99AcJvC58tMO4DGSNCeJM2ACWaMAEJclzktJXdLcqe4VZdS
gm1Gr9V+nL9cFdnoZDsujSO0Fbx1niXrifreTB1mSWEo0VES4xxdirXlz7lDe7oHZwsqzF7Wl9mJ
qC/dXOe4IBXXw8lIO5r1FEOwxK1539b4GqyzqE7W2PevjW7C1Jm34Toq8pGhYqIoR8T+JbSOcBEP
8MZjwtSlG5gcX5BAx/DsR+Nk9dDhuXgZ8IhZHCsQVIssIQlnMvAPh9dNeRi8RHpwC8Hv3K8h7Ipa
csGNk1NGBxntqPycVpneeJne5xDW6HV2SWTgypPjcbT+l7zLdYXLQeCH/c2zMNM4IZzp8qxsWx/g
r74Rjm1TVZOro7J05zJ5/IGqg7Gpa9I8O9+eTKWY0EN6bBZakEfPGhy/85iaNZaA/aqsJ/E5h84j
IzZTs9LUE0zgeA8CEooKPSfYQLAQ6KJpsqz5nWJCHoYd86wXJdhdogGBYyVyltMBxMNkElR+P0k2
oM2inFnkX66SF5DXDTlKkMOK1X3+jR27Qo9LcHw5ZV3WzB+xyfayLOpZP4YzgaJa65JyIyDmLRmV
Db448rTFpCTS8YFlRw2lZuNKCAXnPfRJ3TKtQFrIeisf1FVenptjfeWRSQ4e+5zdAnkmQSReHdMx
fYf6It5bhdsHx9JveHsUxnmJNIrpzNmo3StJFe+7geijLVFKQj8ldOvdeVFAAJWKVdm8TkccYD+p
6YrDJqqVLLvTv/bDhUQJTjKiUIfW8onaTe5DxaMFq9MTZpdIEq7FP3uxJUyZwKIFv0bQY/UScLLt
gfxP0co5yx/t7YY9VpzwbcDNQPoABXErrmTsywK8p27YT67nJM1ueBzt74RkHd1OGarQqIF6PpLZ
ObAtugqRyu6IOoVr/hd0dwmVSaFdpHn7G7119jGxg2wHjDWgcP9UlXj3djULFLN7ZXIdLdR9H/7y
NbrDAhBLTnnRQUjNXnbRHAlwZ2zPx77l4SJNrUn9UFxx3ssQyfT+ufT8B6ha7JSBERIMgcsXHcBv
YucTf6h9HAetWZ3MdFwV/0Elet3nMwRtyoCwbUwbWpFo7/VzmL18+PeLxkh/8hRmvTxI4WtVDmzO
7yYPamaLcVtMvxSTUh+ywWpmbJGL8EiOmsAtJlDr0HK2XJAg7usCv6F8ZVJxtFN6xEFA2U9soCW7
Wb2vy5qxg72wVfUFEZSxRpe/C9DbgAmklI0AMu0i4VyTAIbGnReuDQU0FrZGkhBT2p+Fd40sxFEm
EhBLXKyE2bRMWZihIsZ7y+EI2ipGGRkPVkMFmF+KIY3k+xbwcbdEzTnE6hB3G7BoG16tCQnkWI/d
btZjpL+vsWdwNMcMqBAXjoa3W+aVgAZCHrrjcXUfcuy6WGwnHrOWHBmRn3ytG/5rAwzGjZDUAsSJ
roVzTVMH+vh8LIgxYwIOdEw5mYnj+DolYlefdK4G0mtCzpMtAg+wu+i16fEDN+DBvQQHBb9gS2SP
+wr3GKSuSVP+s4DYjGYD5MMnwxOsMAZkNhTspwDdVFeuwvq3bU+rABc9HWCNplnHSNTUDjd0yxVZ
MAdVQw+NhgJnlvwAU7xZsFOnrkIc9K/bLila8ekRtryXSTRgxWV8qqEPQDefU1Dcdd5cw5cZlIBx
5+hTLOcpideVxxTRiPMbQehHrjvCyOWPGupPvK+lBHsbAG8GjBpXV2rNEf/YD2iVLgBF53oT7kDv
iO1x6b5W/3u6aq1Wpvxluw1FIFKkA/ueaC3UbeRpH+TZ4QnRabVNMYxcXDVLDwEMMzsYOTaXo1yb
U8ESrC1aWVtoRzSl3vf8zdoyWeG8fY5h5v/e/hIIhl1ZqbCp/c9tb7QcSamtpdhnstqM9hdAd6/A
l6cke8Okx1/uEMCbawYl1Yvh1vZBfjyP9hWnrnPZyb4RZx1OlHt5+ZESK6iT3SFqSrQ5DfXNRHa+
YnwVYbQBbf4U/reRk0JEL/r/gzX2oy8D7NHqXdqPv5u0K4iEh1EMxD9g5wA+v3B2fbUbqo8aBEu5
GcaEYJLIyoKx5wJVo834vrhLHWiX0WWs92bq8Z3oXddNo4dl3DADFg779S8RU6iz1pI/nDZRLwX6
kvF/C+luMd6oTDyo8FEYfBsYmtLYbtyU80/B3ydyjrIT5gB49eTROWioCSvV9LHtH8VgpiZJU7h0
E6IQ02hWHVJNcoBoua7Cj2jNF2b0aTrUyI+kOWBtFMVTzp7DAHhp0wPnbRxAHkaDL/CKj8CL53lR
sN0+ei6VLVQhyjnoHd+6q9d7XWAGdJJfnG0b76TsLtPTJGCZZ9uN4QDJaeRFbDJKKewBUhOphTqv
qAZTa/VFpSRO3uV6W/Y0ziyC2/0i586SgHRoP+5b2wbOlwqsh6wVjH0o//bSxadenT9+W/3Dygeq
3lT0nbOnzyO0yZL/bmgOtxn+owNzZgZycQ+gJo4anet2gWT0V83hInhDBHKjU1D5t5VL7lo7dCN/
9d3rQ95B9eEdI1PoCOFRhEtFtcddISdAaQ1UM0QSvlko3xYW7nwU4t5xfEYpd7ZVcLHCKOrpqdiW
eoRmrmyxKYztTPqp6cLqvDRGLWfnSlKbW2rutIMd+D4MkFPhnfN5doEwV0kjvd+7NkANt4incKAR
A+l4Nfxd9FVKNECW/yWulRa3sWv1MDxpJK0b1ikh1DmfOwzMULK331bHAY2x379vPnqE0Tz9nHvx
vrJWnnIdwAy3CnteVp09AJ25tZOCWOmM0s69dUMz0lHd3A/zGK6exbJVV5+koPmDH8KYQYtGqRnP
cJxySY4jcdHh0hWRx+sTQMUtGJ0LXLKDPVOZRgbQcbSJGK0UnP0wcR1z7155aupReQAnCBh9oKwD
Dt7UBmNEk8xcTglOc/3WKtFMTxKVcjfR9UeiFNh0RTpZoJp3QcDAbCrJ8tgtkLbowrrPiPjDoiWE
aX2BqLXY+IphSQsI2/6mHap+I1f8+FKZxGJ1VDPPvE/ytyqjuvHA4zVaf8hAylfLY34pn/hxJED+
134V9tuXXfdwymkus4qM0+0x8alZGPgJp4iX1IE8Mgdf8IhmZSUznbI4Tv7tnbM3AnWaUSA0CO28
7gFWJ8Tl4c+C2JeVNk77XOylZsv6mymHSPcMkRwqW8yoC7TPc9TvNT/K++ez4Z+n2CTIOUHnCf2K
Cr+Vg1EdGi0iMvDHkqON5NqxOE6PqhF7BmzIijqZfyMWAZxZzM8+vOSpHKEzrFbOkpYH3bca+zpw
S8ZWSUEzbS/yllHhe9RTSPXfBiKPcGN35BhXfUc4joz9Qh+aJs3a8vOzkEQtQXDEyH+zVeSyjrsN
UpToZswR725KEemHMmUXY9irn80E8aa6WAWxSx6Ww0tuzT1jTBszODENFmblR5r7Wal271N6CLjG
mN4NV0XetxidDsF9ajs0TgO8Oby37sdBYT8gdk4XYCnPg79v2lJZ9y1WKvfXglcBTi+eByfH2m9u
jkplu3rtFT8uEU/tlZdvDt9+ui4qM1SKdGnJCT3MfB4rVO/g+CYlaihd56DOjvPky3CW7gAMY35s
VwZWpUtpaumUBIUz7wr6IJpQ//phAmclXBAcPDwCowWS7REoBBUJ5Ch2gvqF9uwUIFBhZDNNNCrE
LwZQwpUT3Z3/ZlMxFC5n+PwpUw2u5Ebqx5W/0pVOIjikfJi4pqIYGYJkLzfIDo4NKS2LShqjq/w3
t+rre1Svkm2reo+LiUlOl12KU/eUl72//HCCfUC44nzPY6EnIXL0OXSBkuE9oCOygVZl9XBmMY2b
v8aMiedfJ9EQT7laIyc9gyoAAF1aNEvWkNktlzWxKdL7sSRSPZvqPyAt1mU3HHVhtwkS4K5x7+Op
9DmVeHYLcdc1Qr7IYYidUQGgtFQ0S776+K3fZ3RquBDCm8gwUPHEXQcc7OoWJ63R0aV+8W2IBnsw
Fz72QqCyeywFqgjXJAffF6LxWmrcu6buX9UYf2tEg3LUM02IR2kKzkiocpptfEtbOFYkCEsIaJR2
cW8WBNmM7m+fDwSO77C+1syDvK8l+6qYhZe+RSe2IoY3DfYQkzBsH7a/BDMHLymbBxZKuJ8STCT4
uUSMVDvZHHWPDWwxslPVnC76ovtn9OejouMyRvbTFCEWGxzT8gilCpCKmgsEDkdjG7EuHOlH1ZYA
Wu3/rcgGaTcjeWZ8jbEBGc6XHQ1NS+slohao/npDzYosEmqEoSLfGJ7Z+F6u0nH8lR0au2qN+1hK
8nt/0zsnq0RcGTIuukz0u+x1+HQsGbXWBW73UVP1EoKrE4R5VyjTi8vb5z7ER5sivkE+YCLSwL+9
GBsMrWyEbiW+mKEa/n+TJBDatBsWWdYc9x1BXxU6Qgkr6IbhjZ3vMNu1kUqcqt8+9K3rb5PNZ9pt
To/7w0JTQ85481HPbpdyKzhGliiyimYrrCjWOw1RbdrFXLVL3eK3C6kVaDRks1C6QORNf5V4Yla5
wFQ/StYSnJB9r5xIK42ZejPS5RhHhUhtyCBEH2W86lHLQqvc07lDY5VNu5rFrtx2RycDHKXaX27F
CZlC7xJxhRmYlHzIORPiUHrVvP/pkMhEbmH8+XplbnN5a9khuP6qjkzAtbKYMxiaGHYuNYp8Tw4Q
biZMqGi8b1BJTHUHtADo/m3s/whim5/UG2l7sm0uF1sL6hE+fBle8FmWEDwgfIF0si2/QP1j7D2D
P1lmCgC7QBmHF+WnQZKhy9J1iDUHHzuVvEbOch4lsrVkUUE0Q+wWuPiG0xcuILvMZnMZzGjzODFb
DprwbWDUcSOxhvIMJjl79KlRWmo/0/XOwk/m4RIW/m4T6yFR4/DAbJGzjmkGghFHjBUg/WbUanoU
bpGPPCRNivkiGDbR4EJ1FETwiYUALnpDF2NWd5PzaVNB4wVZOfsn8YRWcLO4sne8uyfDjKLYcef0
7wm2SNKnT7F5eclXWyhmGMAMz7V25jNgXwjX+B/aS5/AGz30iAm+xWOEvXw+ihou2/B8mh/3iCUP
XybLaQGTr9m3D7mR19VijIIy5VY2WtK12lvN2RBsh5o8+H+EjlG+X3971i0/pEaFtOEx5x3w6MZO
/3BLwgKnROHHrlcKUDx5+yDZO88jGQXg5lRBNm41bZNAmuRYxgEqS6m0SrVE9oc7GuUfn4p5OqWD
lMs8hk+7QfmRyHd5QBCjRL4hQCQdtB9e6kVvHQbC5pAYGoC/GxI04czRBfzlngEUIkREtM4AhFYb
32nv2sSTdNNpW1zmbl7gkLLJpeP2xLkGu73nwpfbzPtRvmbv8d4yXQqlG8mUGGGq71KChTNRS6zF
dV7lSZg7DtnrFjWQX51Co42hh0iQLnbSDkvzv4JAljuRbuIeL6XJ5EDuZ7BXrOfiNmCuv/srKLZy
1ZHawcIno6CE4H9vcT4iNHSNBXXYsnCtizhiLWE6UQzoVdJYH3yv3w/QBxW4a878l49nAqTPetbI
YetVDebO1aOXFAu133PrMf9OrfcgcEz6HD3Lmub88zxab0VIGpC373knhaI1lpeFL6pSD2m1iHI+
j58bp5JbL+0eLE19K9OI3fPHaE2+ov8WOuDnmSxi62TqrIVnpx3I/WDofFTZiGa3LZvWkm6OJer8
A2IBQZZll+j/XS81N7T4XuAw553JKKk+Wu0ctXUj/woWzzT35g6HJEZ9ThdX/ujccnEBPWCy9oZ9
Fs5iUaLtJ9zZ/V8dI82OpQpTsMVRu++zN7hWbOwQ9V4SKL5VCb1cwdkaN35TV4LppDImBZMgDVbe
bg9Dd2CIdDi+MUPuAeYkJ1FDMO2csR6yOYvaH0+KbRnJEpNq7oEfRTiimM0usBsXUJ+Zz3mUGWPq
BJ8rLnqw5Ca5erqedKefxoksHKBFGgKJJVcdinrtC0V35AayPTHfQJxrULLSNYY/QxIVQ8uVeM/x
3eEGRWxjz+DB6eWtfHlgEipFU1eEiw9rmSSEAe2yjyMwdt27bXbpNiHN8zWBZ06fMQGzMjwsOVvZ
E+XEuEs38FUSJkZZhKvWySbPkb8cjYzRH5ic+1UEdc1x2o7DtxSRlKt7ThZf9XkJgK9gBfh9/ldI
/Hh0Q22jIg3wFPIEW1tXQJaLSGfnfAvzkZfclZE5RxAVyNMLJvmonHAcqE63HpbEXHzd2MdYHSer
w2+/e0oqX6+tcqJ0UKy8G3Fe7BnUwPV+3SLJbTnDu4C+/D9bPolXJ5rxfgce7be9xru0Z4/pQhBF
5L49Neme3Q8cHF3JAGqJYQ6zwrwbcVOdSV860Jk8B4VmqNPp5CG9AnfsMZTrvDcl+DtoqwLlIWpH
XmM0Kg+a+YE4N/k0rtbWHQ8cfoqUr4Chw0hCa6Oc10pcQXkroidkKrPHPQtqtVbevIYCUmw3QMUV
ZkKWWg9CARpu5MqT5/pq8vWzFzNWuaBgj2SaNZFOuyywB8D2bVi6W5w4NEn1VVkSbhWzDX6Tdrgv
H/wNE3MfqrDeFA7jCdBU3Xr4/JRL/evOKotBj0XNeLr3DDkn/05I5Eg3PFL44GxfCmRKG16N+1dG
wyfR4oFs+X6ItDzUjvUAZpTj23qnLYAv6Qb0vHm+fBsYp6G77mqR6oQ3YYGWBSTuTBsjDSFzpvOF
y5Fv0yThU4MPmuabYR3LjUFPHXH4Hdyoz27s/K/q4uoOFlX2vcxuCOdY2QK8JWNF015094z1zvXe
GFAgQKG8xDBWZa43UsvqCaBc6Sacu0M9VfEfrS2zs6cu1FXyTBrvV45NA0elQLnsbwdhnzjSzNvl
r4tBp5pLCOozyOZvq8vi+Uio62zL90dlX1BXQMQpr4G3RZKAOAFq9uQ17j9eDTSJGyC7CO9fiJmW
qizydOlNV/yF5L8tertf+zAkpPIA41PccD5U3yfaLvtbyoaBFfYx/KwhmWZfUc2HGRt146BqqtmX
Yib2A+9Nf+tKjBotoZsjA8DPZaOZ9Ncoxch2f5xj5hZ//pbhwQNyiHlaH0I8jUeAazOdn1GWn/9s
Lwo765wWmWs6oL1S17DCid94GDBffxiW+SxmktT6e2g+3Oj7ALHZY2ishQyi5AJWQ+RZq3coi0cj
NkwRwc9WDd5Ni7nEAwk03wGHT9WYVg2tpPCOFU5TOyAL294W59PxbU0dezP6d40uqmd+xka/ptSc
Fblzmow3uOuvHR8aBpQI8ZmAlAsIF8QdEPXMgjeBLPV+HNd6+6HDVeFH8HJQ4YD9SHm1i7N7FjHR
xHQDDz/JmesULCGwh4aWVQO8tFCjJLuNBz72B+N/NbiyiEFYSZ8ntaWpQKBRxYBB7wgFoowMFqdH
eRhzeZYmyMDl5BApvb8MiJeZfWIovQn0YA+P8fkos4vJpUjxnSQ/FPBDIFckm/oB11n2pAtT+N0f
HPgLOaCtIerm5rBoNhFUQV3N3f3MaVWOpQuY2z7qMsAi3ZKiku7DFGSnO8p0MupBOdRadXOepaKM
YEb9IrLlgTditmOWUqvGn0GUZzkibX3PjZ4sjZmbTm7kK/YJy3p9nAqPyZamkz8k8W1oE4npcPW4
J7v8Zw/7rJInJWOp69d8KHIvZ8WlU22GLN4fG1Udni8LcSGOTEO4nyvj6F+Rq9WuvyUIf3qCzwxs
dPl2SdkkiS42T9hjKeDTa4o9sl/6EN0bj8OUz2K2qRmH3RIEBi+5ko0DnNqWgz01MEdF/jU8O+XY
PgNz20WhDR5+cXKl7rGiFL+ZkcQ76L7cj86kiFaAOq2Jd/x+gdPJl1Kp0h6O2AchRtloUrtnMAKb
5YxPal6ZOnse+/6FNKmt2zdv3QFcJh/NjEu7xIjQ7+YnvKVlkrYqyWz8OvGt4ZLcnPMv5WJS5G9I
nCMCUHDJxZ8Po06nen/+xIZTKYhTcj2CTh5SQOqznWVF5bL0HuKFXQSciSLMPqUjyQMW2kt2HAI1
xWc4Ol9rC8AjG2/DWKXbiCThoBUkQkuik6QxnPJ2svx/59sU5+rf5Dc/8QLwO3XON0PR/LIpb4I4
vddTdUEioIF5d20YQyStant+ydqXWcmcYTZSZczmlHifMjn9mCceerPNIJ5bjO0P9e64Ov3X3R77
DnwIaq8XIaqN/CVjFxLBWAW5pzCD8pcVJzWSYbregumrmyJOENXdDfOZE/x4lQg6rgO7k6hxEQsY
GMUNAonFDfffwS6V9p0cuMUCMOsILy3GacvlaLM2JuXRtVtWioDV9fkGZUdADgYaYNAC1xR2aDIt
96h/WY713ad4FyVBRCGjK8TBsr9EHXdBIcDYcR/1a19MfZdVrAr/RQMO1TkxxWSHCp4xArVY89gi
MsCbE5s6CVO9RXenuP/8KR6rIUpwQlyn1SLp1ximF4pRFwGDuWv57JbfJnRMk8knDzjefvXa2y9a
+b5AdJmPhSbaODrXGdtfkHEWyWbhPGiMq6V9quSwZ/7pMmDp4jfjw/YKd9OVnKOlSgEUKwB7Axcp
mTjgbw9D8w0Ep0l8jDaUh1UxkFfy581FM9JS9zWPLzuTuHAA23r3wtC8XMAW1aD/Y+h7iDZoehyT
+T5fJVbuJnuV5sQK+GDQmU94KXUJPxGq9gDDz/qXqrrbD/m+B5oMal4CHs2MNfVyHx2hJIipP2lC
frbckagcv/+Qzatg0cvOQx8DeuI/+OBq/hsHp1Q0LbmuRO2uaFPnBXfDv9e73R77i/wfhifz2QK0
BrPqoy5QP/jILlAS+BsWrBa8qa4pFUFWbUUhXzhMcbtrGBsmYIlQGbp6YFL1QCAYk2vibFzneA9Q
b4ebv6G/sAw59wv553WzXZOp60UtafldSsnSzc5G28lFIGeKLsJ4IkLDvf8jH6DJ2WveRvcSuVST
NNRYeGxSwekoXvj//zPLcybLb1C3+WbDBrqYZaUbO6JEvizWTBDbZVSc5QnOjw6nx5exe5p9K0+v
qUDZjqYA2FD5Yabg9A7p1kRLqKi8F96FL7p0uE9e2xuzfl4aFaUTlIl8jh4CPrwLVovnVm2q07Yt
o2k64RS7OPDCf7kdBLnyi0it0/Vo4pKMDM6SrFt4WRupenogoz7kpSxlBbZiIOJPpJNRNaPET8fo
vOv6UBf3k13MxHZk+QHwxqoT9dRLKUwL8BUB7WS2FnIy/6F+zrKpgZBVR41tNZFjafTAGxHEyT/5
d8tuTJU/Axx1nLIPXyk9vEn8ZEA6qdJ5fvQUSdOP+OKX76XL4PcgbmfLFEZaWR7HRIFiVEdFGrw7
intYo9Jf9hD/X89DmTg64YIwuWpRskLmzRjcYhkm3jAVtOU0s+1kSqhUa8YuyzmvDty4mun7a3zv
mHURnuRlnxQTHCf7/HwIBhXc70v00xMynp00oHGbtKqFNiJhlOwCsjFLUg144yAGw68mS/tOf0pm
muAn+hNeFihQhh3nA35Z+V3wRXtLjwD7vwMg8JPl09SknXhQDzcjNWcYnXGaAcjJP9VbZKPFAsyT
ue6L8t2y9IEZvzAVHqxA2fz1fGA5HRWidAKEKszL9hFdcKDkFlAu/ARElCJSYhY3M/tGCV630Aa9
IyMQKYdmW48DZq3Uy+yuJ8k0fbnyvZ/BmHAm5wkk2/N6qwMahuwnzQxfMnTiifLIhHbBjRnpgTCL
TRjSYEXyfCuPtN9G3c3kq+aUssJia8GOO4cNJBG2M74/EsWuW9LWaFUpn2KDC1Jjotu2xOT5WNhd
yMgdB8gLQIjxMsD8JxGDN5Z6M538DLo3NFwrl55B6YARPBBz8qH8oKy07+e36VdUkqwYlQduv+Eb
f4rl/8cA8YAvwWqo0dTYRKbCAJC6+I4F3381Ym2wEBFjvnNWuQ0cU9gSqNt/n5wYZH8ZMIPZoPyC
U0RyBBBwrUTWa/+OsQPNrlkkPy8Dk48a0zVJghQ0tW72Gl0SVaVQtBM3SFT+LZhN8w2bSLMJsQG/
UUPEpTYfSOJsZrDAfVXhFIu6LEokMui0SmO6K2FdtLtTbOkbF2YBp4v1XpwrC661rfVZ2zT68EWT
yXdkABF9kP8CpbQpT6+docz0KAVER2MR1kZGuwfFfPwg9jRpB+VB9Q2wocvAlG1TD5+uZ2YPSbt3
wsD3DPxHj0GquPeObB/OoH2OcUVUskWcNegB04tefnlCXCCO5+cuVkgn4EMJRoA4iokhKs26zTSB
wV8bM/Qn/P1nQJqpA6oTzyKoIhxCbT3amwJIiwu7zsaUXNyQU/E1ijY+2bLWNPMDx+VND7oAU0u2
ZKCnNu+jpu4GqrZst1Y2mmOxt4sZRxz/xNkKFQr0VTtSNvb/2lxau5AoM4Zb6+FtrzoTkRg/6QAJ
C1WAjlSl1pi0BI1KE5g/7GqCGTNNcD8jK+KV7K4oTJpOv871+xyrhJQue9ImqA/etIua2WI66a/q
0A+VkSyQRONPcEDQdMkXWG58AwbtwfzjSlh08LaY7/oIev7nh7pCeEwdK0UpjZ2c9XElLS4JHp4U
xBa8oyvL0Gz/iZ0zQqnwIiQ6JlZ8tc8qJY8NnlrjNlwLQjXLBOddcKIJ7scJEYTSd3BMNKrRhwhn
hsYRMnsuo+ikPBLNASz+DeuIZMDDul3ljwk5UG/mO9sOt77MrbT9dUVLz/sAJ2B6Ojt2ZrGZw2e5
AI8o0g3fuMsTy5esaeRMh25/7etJkM35d/lAnLvEmCrzWdAMzNGvrFQO9Bm0sVbcuWULHIlWQS6U
zrtmDyvTP+PEKMorCT+vpzvLINk00YkJdG37GWC2l5HiQsOIjih1nE2e3/ExFfnP+t1LkkVidtM5
rlvhkeKznSnGr/LwJJsS+fJ34//+EtsrU0/OBWT1kBZZ4h2q6o5RAOTXlX2SkzaLaQcuC/AqjDk3
0kSwBFfWtqoYwbLDe5u3sVbZbIiDQ2TJ9YcsVvsDoYEjX3ERV9Dqs+qhk8nx1SckvtFXxdd9L9Tq
f719btopBFqS1eZMPJkA+bfVhtcbDiyfwDjeXv91SWsGOJ61m9arVJo62Y/6Al4kvz+kOE3NwQLd
QKgXQn33/EdLK8QqPg/HATNOFZKBXNofkagkS2HWi7K0pa8x5u+I4LmtmxuBMG3GJY9E8S97RPWZ
3EMQFUyED3jiCUsYNo2M4o0fvkFjEZe0hcIuVP04NDZZYE065JcTM+U6+RaQ9ZmPQVeOrGutJepm
nZHlktrMmJTtmf+yF+yhfJREWyihKeaLgbnUe/qgU0P+ZLGTF4hVmml3IeeQrcQKvR3Z+HdNEe8E
k5p8zxXsEY4u0fS8ihqV2D0cZw1q7ZUlCeFMFpAIiot7y5be1KpBepQ2YWJkOIZi8nuIDbUVr5zv
93huiRVUiFnFqpUY+YfKtMoo1WNnrZlGQRVwkHIPWpAn/JEhbafnqYzDK2GYJCS1RrUXeDOnWtQu
f7OEMFnv+gVTzzgNv79vHME8Sn+duNvanboaMlO1QeOS4MvjwC9OFggaN3kkQebMP/bBz34zMzRq
6QWNA4FlvynuZcdYd/f5BUSTUIu/i5SgsDq0+djCk/OSVoR+AE3ZOC81B7J+sjwpMJcd8+HPCdN8
9lURqWI5K7abgFbYzzEaqz6aRJ/FL9nhjPixrT3XQwu1tt8rk417Gij1D48pXrOupdReEXhnSYpS
WmCGmKsopag8/EKH+4g0fPu9N7yOQlANMU3ATuMUtbLMOYpFypwuEZWm81hZfw81SDfpGG9L6yT7
UXG13vDtmVIu9VRCjDshd5CnS4iEOazJp4RUq2OrC2DEyX60/PpIsqRB/RkPRqC+Ttvi4LIv9Z1P
+0Z6Sm8/go+rE27RQcn4Cifbf98bAZ2avVwMiCwvrXo5k0uwonxU8A63CxsAcLgZbS0dslvcPJa5
IyURN0Hju6yoDTauSORr3YQJok58yX0fdhqn9gnzolLwR+c2CZQ90xoLawpAc6vnuZZESGin+bij
HYYsgfc++3STEbSvfMyYT23voICNM0/PaelklfOVaWxw6gF5C+M5X31Lnukd9sMWkhl1hUwmf+L0
4IDKjMjkVzXcFuesBf+xJfyYOw2vzJXiGDi4oQL9k1HiLJJ2CzlBmSauJFT/2E7ixL0eNwcgDknY
rHM3SlI3t//B742SldjGQjFgvH4PtpoyeiZ0thged20gLwymVGRlZXv0crefOmYvv95VQrRbSfTA
seOkreH5HYnE1WqfIbnSZJrWkVu6JJXay4y97oYt/5eRUSM1vYNarCF/sc0S/yUzzREtjCO9SKWV
Jwth5Kkm5np+Pi06F4o1vPlxMHLg7lNw/zMUMtt509oH1w64TYt0tDW1dI7oyvUPdtGmJIrwIRy9
eZIGswUZMC+BoINlGDUGLx0PidZ2G35PURQYfX8t55gZAUBUs/n+aEZwR49oP3bwTlhahmZmbP0A
WxDaSDuWJgzpo2lRPa55GrfaI3z5UwnNis5V4vNylKncZCyHo5HfqYaKT3Y367TJ/gW11AnA/2ag
EnHCgBSFxtCY8utfcplmFg6RthgqDmOYhSXHDLdY/qoUNfZi65RlaKc4crGZVC9vd016yIkkDYeZ
BhrlLjyMRF1ef1K/1lq7lqKdmf+NVF1nOHlqbKV/ZrCfiffJQdg/KZO9IlJcPY7PvcLUa3+whysB
zY3mUmKIrUGVxNL1KmlCbfwuUw1NROBvJQsHxPwoQusXCoqzzMvw+WLioyEpxolPy8G4n5Fo+s61
vhTcwr9wFnRhOQ8RiBx5GqBVDWeIWquP8V0KFaAhGloILUNNSM8Z/iJfFWJ0EQdaW/BLEc3u8ccd
6WXtD6kzpYV/qc6DLT5oUgzocjUTwP0EODw9l1yvc9mZ7TXIZevaKDh9du/JcnKKvVS3l/sM1J2B
/4Q3Ikj1dq8E/xYBDOD5bJA35BTiAecGT1jGdpJDlUlo9T6+jFHhAnIFIEi/LbT+KocgzE0pLbXa
iaHUq5TvGueSi1EddH8776RPB4Wtw1j8xyUsmZ2gK4kXmy+7hDnvyqd/JFzaWIqD7AfPdaooEmb1
dnWwWcfrkuhXh66WzDN4TVo2BTBxLy/gODAX0GaAjUw7SrxbHliwvkc/NNDoYaOOs6coYiPmSzWe
fBZE3RYNFDA3tSp74mbG5zSqnDP5uvtpoPKhAIGPfyVV15aYW6vGXaJ45fsqfQhlZEikfzpQ4VbP
T7+NPOVwo8BbhbJSvanF404CdYvCTazIXNqswWmHPTNkMqHljipNjn2iYHc05M+FU0H4dMxUoszZ
TJ4jVau+oQejRS14jGgl9Pt67B3kIUyQ1Jc62BX0IdVDkcHHSTvyjXb6LbvzEKoplbycspiWVAFi
jVh8BnOCYsW9nAZfk5TdeocnXRtNNho/HDcaKpg0OGn04r+qVZ7qv/hgIsciurCtV6T5niAUBUFj
cKNpcw5XxogE6IgdnP8BEvRxRwTqg8arPnttDJXWOLUZzh1X73aHmFvdwqrAEvUJyMsGDe1lox5B
DqcJ0QZ+sTmvot8SQzALu54PyUDiNcdxE9gAsJuB6B5t2vYiZSgsw75eQis74u4unOx6IEFBkABh
OJg/NGxjCHMsxrTvUKHuGCMp+aQgf20A8FWJD2mNB8oPXLyF0i/M6MlLdZcnmMbWlP6Px0QMxAdb
rilXqYQmGYhpoP8LEPYc4F8WuCnqf8dkqS2bTtIF0vBU7rBfZfuCSjc8UX1WNuUNZqYbcAH2KC4/
1fReprQTV4GPCPaNQYRu5zTsGFNDj8U3R/ivDgBeSc5MXeSohz7nQF1XFKT7yDxL0DYQzrzvjMtv
zeV/4awdwIS7cDSfIypa61rDQdypR3QZv9/xItHPWe3VMVeP0sMyBer/W3FvHjbbV4XdQnP5vcEa
3Y/QjLaShY7CTUtG76Dcsu68hfm0jdm5we+AFG4b7++w2+I3rTyD6/gge/jGkmQH9rzWSxCH8u5i
GC3oEgk5ZhX2NrA/FqpJ86oltmPzbQsI0h907Y6/7vWWyqbD6wVXBx5gacewIHcxP0wqXzBxRTiE
H92kxug4T1fGtx62HwoQ4DVbU0FkKSV0hxC8L/DX2+jQzYuN2zj5gsslnCaWFCCg9uBaJtbNQFAS
6DXB8+Jro25fcYr1a5zT6XtqZunT5IeZy7RJqLtOLAVqFEyOA9fMi2ff5cOMOkP296NrpiuktOD/
M4bS+t41IkxFywBHP4ImlIspJV78Rh/2GTVkNxwTcov+jMDJq6wZzwG9bZqitoctMtg+G00YYsz8
HQVe0VFnwJxCj5Q9CUSZLAzdLkGxJvgiJ/MuMsFA08Bk2LSJ0L3qn1M30IAAAgBkOwGz2sYA08LA
/A74HV0VTdNDPonXG6tyiRaLEWXyObBWBRr6iuYAp4MFA6lAQuSZ9HnqX7KnKL6tnAH0RBWQeeo5
pu7W2TsA6hHEOFA3UDdH3TXSehoD3y84NsgD8j3zOn4oW8Uic+C6NtJa8NFPX9hhs5ihaDoI0o8B
8QPPVKfo6eIl0l/Ma6C2Us9YZdOVbg/nE4sWDn+ZIcK5pzcExvGIh+tsZEptnvReoGMFaF5EcFRE
ACMfYbOsi2RYxSZYGlgeh5hHisf/DfNiSCJaPPbfQcQXow6CWi5Rqlt/hQCaMWIXm/OjlQJLkRVh
kzdOfj4UIrD9U1PQX8IwbM8Tnz/URwXWashD/qjxdhdIIF3qj57n+82Fjz6rsH0ctSvHUY+ri0S8
zV3rKoJgT2tWnkvuJXRLZRoI/1LUXK0T1HC6ZMSviafiVNfYBi1eA5B6D1UH3XsNZqavxSJuaRQs
yMr6BwQbiiJuQzt5Cpylyt25t3QW36OCdiFxT4WepZRabdDz2WOB88pzOFZ0Syqfwd2cNOb96QZq
47jnVep3LSs1c/sEkd8HDgxY3cxGwQB774no65vTbthqRScs8YYIWjnF/vTLH1izVzBbl9F0gRsW
iXqsQ2E+87cALflIKpdAVA6WUc29LWhzii17dRfPAj1F+ni8Kz1qVWp93K7T5YxSoixr+xMtSnvN
M3gYBjhbPBugvyGCJi/5tHo/Ko6qGvX3wbRwzEG+TV6S5SsrXyFwB7f5ZokvhGkYKgERbd53fkwz
A70VT3997LSv9gRSwEUORubuPfp5cpyEaEVx3LhkLT02obyZn5yicecwRpj3DKGaKGvMuaB+oiEP
p3Ncr9qA/zBdgAC5D6l949+EEEF3F8sWNZyYnKF/LRrsLV7J8ZU9vUG03va9qK4dQWs6lzo6Iw3h
Urt9kFiMEVWwtBmi4U7/nwyzwjT7aNfdGieXnc4vjEK//B7RzwDXdIIiO9JhFuILMje8zm4msdPx
zMeSem9EoMwxa6bgVeQzuQV3ThjVLL9uwYI6yCR3xovUErtcPT3ZsqE8VbwF02vOKeXU0u14x480
AU+B0xne1sLgw4dcia+RACRHatPdwGcKo4lXHVF0nygjcQMBZrjMC4xE0jSbhHSISxqTp4MU7W2n
bZCF/ZyVbSQjQRLMMwuPBs/SA9uUEErs6tLr3wProd+xwE+Q4tWuzvgP34fLg0NYPu63GUVYTfRy
09UclvLJ+EEokWmZE3sJLdpYFRSPeWdVznZkFM+a5ATkQTg3ZzW0NvYsk2A5u4ArH1e1kR3W1Zyz
1oeYDcdxhl3ceEyLHiw2aMARtm/gp0myhuKMKqso0Ia3/Gqc0i1rVJzayFWgq+G4ABb+F+99SiN6
AoZK90djwGrR4scIpF27/oImz8B9jlR/h31xBVzm0wIlyLP9V+jqXqKPFE3zqOFfYSULSIQ7CGWX
Hg7IttuZqUhCGZnzXCUgPAcd4zjnoJVd4tcdaPW9wsZz0pUnCooudwR8b1JB3/wFaRQxjVarCk/H
A6GoFwwZGY4EA9KbpoN3/DHDwvfyWKL+4e9tQpyjoXDGuYcYEZEw9aShrbiXSoyUf4IRI2pQuIMb
kkop1v4FDsKFXuKR9uJ0VZNnZ3ZMI2677Ox7LIzlZG/GLX/A1DQ8ppqAZiKwYOnqwfDvZB3/J/tL
FVyZHSDqBSnrULmcNncSVbx6q6N4U613MlnsHXP7Mi/TRJSlVWUad91vkcwyt1RaSIrCJQX/+zG3
wHnGhAu63zhXOEq5eWdlNSatVy9li8C5v970qO17OvDUVwQpd9qOfdu8jtKRarilHDVFfqsShvGs
ddz6avMKqVKgfsZeEs04AOfnImWQXkueg9zrFXLMJH9/UnKN9V1PjPwrgA/b95CD++jSrmvsGXjI
eR9uG8rOPllSN06wi/IXzwThTKsmjoZf5OdznE9/bcPzdnJROwy/iymfFWmlLOzp20damUIhCep+
NB/r/2JY+xj5qeEcyDJg0V8vwgm6BpaYG1S7fsVRyMU4+h9ALHD7jYs3R0NejVjiF7IHiHlzIDTB
Ywy93zTNVm4c52zDyaqqG5b9rpziuPr3nfnCIP0qUytoa6ATFT+L1SEoliXPFbHVYk1EYC0LHcfG
xk6I5pMlnxyyIZbL2L7kgmuUbmGa8jG+g7OCB4aOkc3MEviUh4kiXnePVU29l4SzfQY8PwsZu0t6
1QlI8U7vFFGLy7SkfC74b6CR9Tqko1bzFtZPvXXM3yHQzdMSlvXNNapTW+5vYJW6E00CA/kqdhaL
/uBAWcsgAXzDZVC6JcWM5qs8QxrENbM6TcLS2SdtYBAK7RhZ+NxlKVBaljPFeuTe/wUpsTnpOVWX
AITvq9TVfJi9Po6BPwbLf7XbleaHpf5pcJsBvA6OkV6qNZJvMWOY87GRmUcPxufADbd5bCu8Zrpt
AX+pDxoJ+rpbYpJtceCh28jHcBO3IauSmV8yeN4dqYhr7zWpkaSGef9/7gr7h0V3lo4E7NWqICaF
uNIDE3rnoZo4OhiBCc0eO/W5oFLz7LgFHRZWaJRuChVNqGAfzR/KOxiqlR/dPSu6R93MhJoyD/Xn
/7/1JhZIL3fsv8bcRj9rnNUb8b1NomONEqHb7IDyy5zlwyJBv+p2sL8Uaa+f757mLbPyPjESNucj
rB6gOi8wit5OXUuJgos16f7v6mKT71Al6NXFJo6SmE/okKfZ+3yIsAbktgWKj81OCZ0PunVJ7j2C
dq+emVua3eCfwUS4X6fdrTqyizqvS+QjwOFlTHzylXjunPn+V3uAS1eUmlUoaY8//2WpG5xYT3sg
aLyUlN0jYQZVmQeFEvA1IbjgUc2nXpD8dP4mkYbERRijtclBAWtXjQNFsPv2HAPeoyVuJfuJVdVm
Y98VvApERnQeJnsjjZ0f9cpTmft87mirsGN/1+kyNQAhqgJQdIyrz/Wy735cATDW5Pf7k1yfbZN3
TiL2Rj1D/UNvSNp5toPeW+cBi8pU8xeVjeQF9BUoqhUpBb8Y5L7/DqDvcllFRyiO/cc2iJjXulI7
l7FyoFnY1sm8MZVwJGno0tgog1OmdL8V4s2aj0EF+CXpPGhReUTfZQwx2jXGXSZfRjyPhrin2AwV
dq5Tv/1iu3yYVNN5dVXmniFLSvCPbwQT5fpo3i2LaNeo/IfopO0oJPwTgCJjZs732fGAmQ5R+htg
iR89GFU3lRrv/hLWFHSzhdfund5iZgwx2D7kqN6lhtsVMFO4a5TnTfXq7wXygYbRvr8qT+qZ6CZo
+HuO2pqSGXtuVHOTP+FPwWgZdOe1Vh6vo+qZHppMyAwgD9I6ZOnaENVcwIY+vE/zcr64Y66NL9X7
Co2R5X9x2pLNk/EqzI9m7wAXFd0jMyItKewP07swEQ9TZ2XEJl5jrxxQ/d4eoEbvIW2CTSyvq/qV
pE1JCpGvbSQjQTL/bjRIWVB/F/udmYVyKaG5AaCp+BkJXplnEtGUVXI1wT8ITS0G5PLs28dyL4kT
iXmtBgZnkqXHd6mpVB/BtzxgacT1EcRHKLomPs04zTuEezBZbf/IHx9bm4zoHCsxeSpsHhvBl7iP
ffiWhCutU2KLLrPHceYZnuEDcivoRWd9fd+83uq78hB4QI27qY0WeCWoEGMPpQPQnpxl3eH/EzJT
9LPdBIWxQ3uVIHxompjeTyySoqeka4jPgStHzqZVrEXy19ORQgqKbijKA/Yw4NMsK75Kr7sX8TpC
c3d9ccRdGYUc0omIExxp9aKH1NIIb8fYsvdJBAPxK5o0mYeZLXTQpu9/2AOWUjaARzX/1CIfs6lu
OJYASvb9onri/AKqeyTW+hWxo710fiqKB+crD87ePKEQUkkUSPEwM01It0mApx4n/qlY+ir9TLJa
OD3J1ehgObe4sra0FBFOOQ9VK7xAa2s1tFz2g5XExDAu+Bo2Znxb+/tfYq0d27HjPSDRCNAOUSEb
QTcs3aDnX04i5lVsBnNKUU/uIj0WCO7Aq6KJ+xPHMz+5yQo12/xaDU+OLCm/H/eCStu+mAWuqk6S
9Eo0rr8PBWVGaOEMgTnjza/47KHcPEcxuIpklLqpJRyiivcbXXz8T7jwsm8IDskjX5yV9Kj5D6Vw
2CsFVBQ5YT2n0IPxnDEnJ7BwSapE2jGhH7t7AIwRtDs2E9pvjBDyLn1eScVEoBIKJ1aLPd4TUDz1
0yV95ZmqBmrt82R39lP/Jh6wEIgYGz6OFuQyyi/ksDuXokR/s04usEMIhTQS2/EgDWY7U5hVOJgs
Lw69GObem0Vc88Ht7Xc3HEZovPWg0GF8cuZOMw4XJN046pB1DEs+xJBme+JQDP9o2s5WIrgXGbyN
heRlP9MCtQkibRzgWUMt4CRUCSVnnMfOEFD99vg7eveNXwUhVOp25oeLOXjsWuvyMkqBuZ1iXGn0
xWw5xzfkSIpOxDDtk79Q+zMUVAOpTFYq72yECDrNGdQD+YyINSNk9JEbPkK25cILajfYd4LkjPof
4+PFthXPz7ncZ0N+hw++JicV+OOMuO84Gzwdam+Dq5YnPAesnUSu9jDHLfV3aNzVlIcQkefpO/OR
Oa+98+xygHjU/D+DvVXkGO7IchZRmt19Bd8OfxpbHD2UTIC8oKwXouW+MoO9vKnLfpEqUnyIuILF
v/WQDMBFXgUrQMqV6fY2zuUuHrfbYpHuDcit6DQ2NVNXro5tXISQuY7E5eECXB0jJnzaaK0cK+F5
JY4EsgUSjIpAIzjIj40RJfEaYryS9OoCgNYz1Ssz4+lOt2NU3on/HMK3uyyFe/OdzEZd6WC9zjcm
SyyMjTahQSOAERqJmFyrc+bXvdP/yP0CEVq7xGF5vTSR6G8cKvjPzi5FCiXBmSxGalJxCNrOuSk7
RpPAOVxiwDE9PDYyb5v+svYmRiOzxHDtO917GT+VsTVxA0o0f9e8PoimMgoLXd4Z2Q1w8yEQfVva
zBpJiApCGu1a3jo8rPbndCCtQdwmkiDNxkDzo4kLduymQHPJlJvuk58VeHrSsoQOkVP5gyCUZ77K
ZI/v3LPO+09wIUiJ2/oiCduQs9sl+m1iF88nbegW0Ly8dMT8LfJJHVbUt+Vj99QmY8Ygmtnhyl/K
kjzKWtZg5mzhebXN+Ywi9ykpyfzRlTg159uyp4iOmQfWhvFNF10dX6eJCZ+m/zaQdQum2urMldod
N3AGUYKk5mvzyDfBbGFd6NnlE+MtIXwJsuk6U72HHdTFZ+r1MaDHWXn4tfuFX8yst606EUprWz+x
aWGh8FkdYLvQz07DgbCg1HxIvRlgJt7W2LT3OYJqZDKO+RDd9LMTXiYxreSmFWe8z+IYfBwwnyKU
5uEMXyxZtqXer/bX4BUGPMEibnyi29Ow4upqQZttch2UZN8Zsr69ZI1ySxg+Ek9DLUHXOm8Hwp5F
PFoRuln9KBTbWYfrGsRkakpwcAGaLmMM7VMpBI7zToyF2LRiDOS5nQPfQjem49z7EX5tXasX7lcH
/I+t9PvHDS5OwFMpLGeiqlmfDGhnjkgD2KeJTUtOCWwwvLPIexSFIWM5mwOIaeDVY9HMMC8FSud+
himQ7XjzuvX+tdkY1YeWp/HyYM7/Tdqb4IYiS/Sg5lPy72Ax0qyXCgAbR7E0rW9cJVLnftEu4icp
Ux4xOj6dC44MbecwkQpU+8+i/mDuMVD9CEPGCwq4YsHNKvzYBZnG7gty7xsMvLfS7bLsaV+fSKU8
Ty9cLCB683yaHTBSgq5kfmwEYWhy/TyPsW/Bx3HJcaorJfC8sLzMsU8Lysp7N9iayUBJHUzjYH3R
hWqgvpib3J8vGShcAFzlMfARTvbGQfSnvGmDv5t/1I1+O7twmdmH9ie9WsOzsTRQ7lhbT9F3OjMZ
rxqjBfiDS4pkK5D17SQa2le/mzdCFGhV5wUFVCu4mE8z9pJlEJ1R5Yp8dEW0V3AmvJjHx4+gcHa8
mT8/9PzUrcORNQlQPObVtMEhTD3JhWgOH8DYuONGkhNqeH0Figi2uGTJtxKbU6vpf0hwNoSHlEj5
GIdznthmz3t1k1Y41v9Az02t/gd85Ksk0i6vqC4Obn+5sPfndCIMSxPjx5raPqQqwPMKfjnzP09Y
fiDc+Zp+tZqUgu8OTxYz01Vzju1bETvhzOmqcQoAtx6HQTYo0i3lhusitwgYZlTxHrSSrVuRFINt
pT1QNfQUWEt3lVLAE+hvN8lH20LyXGlbcsTnIgMhPabvae250SsmZ8qocjApCax5ScyAYWDltgRT
WsWBMLvo4+swEyhKlnVqOSdJ3RqkzaKkTynGJgzm/YyHteoviBlgga7St6/bGzpfX0J051HmRHW1
rF45gej4yDaY+3HUZnD3lQJZ24DwArSeDRhMdsPZf2NanajcqMctBrZslwHskDuXP+Qj3oM6NgnE
3lFFtHgLvj6ApAb9GjxsDe/D75sr71R5Yqob/cpxE+CvvBp7aiSafR+gsB3BwMGJQ1MhAsH9meep
EAnhhteq/E5NhJifZo3JN3bBor2OB964QIGjRHLtSdj1AS1JY+fMgukz1TAF1Jd5cc1AJIG7zHE8
AM/hDRIU2eyIl0LZLZ3N/TlkLOYSy9FUwENaTYamPy0qvkQ32vtWMjiEhZp0ctZzwBlng5V/LzaS
G5RTIzSOnSReuMp7EMbokIVf7gOhJOJbC5bXRZbBMEOdeh34n2Gh6bLtk89anZx/PxUvNkKhz7xy
ie+XD/a9QLefw0+VOvOIMN+ne/3JkSGLVye77z2pG3w5+/LMAPdz4VJd2vPQ2kA9zW6eQsZuTXmh
lGaavp7O+6rcsDxBs3tQPRowEr9EF7hugqOMOxXQ59edzjsoIYM41xk2htyEiIix5a1K1T52D87v
qnlEXz/w05roDhhhDJOYheL3qNi6UzXmIEzuAb3mjWz0PCYU7smTZluWTr6aEslHm5yogK+ZdZNL
niYKS3VSeyhKdLNPdGAClOxjQGjQ7qmtO4H7aWzZ+60kcGAVN+NlzFArnfvyF7/LvOHDCNFS1SGa
i13EthnOUhvWuiCXpKyc7V2rp2Yb1m5XM1l3DSeqhM+Z25LMBpRPnudYrkn3ja0sIrqHFS2PXQer
owTyO9HXQzSKBJ8756wh6qxA6hDC8M1Pzvt+L3OG5DfpwlUSGm1Ats4I7zwjTBbX0V2KqSFGxPDE
YgSAXQpegEjAeKwTpP2PlT8bQpqozjCNlfGYqROwZ5UBD5u78Q+VTGt7z9x7QueFA+G6zEubNz2M
S9NQoYJlqx7uOIQ6cgzuPf1by8lKSJtTfLpIk7bP3MjQj+TuEhNicR6RZE6oZGr+Wvtd7TKD0soF
Mqqz4lcA4W9rBLTmgY0EQO4+ctds2BnFpimYA08FaMAz/vAZ+WtjQG56ShWmEK+zjFYP+zJfE7Vd
T5K/KOnyaL4xCXzGzE+qwrraJWfC6715oWm6HdffxbTgEWM+wiFXeMmNvSmgaYned8g9jOBgTG67
Y5RrDNY37ctePyzmhg8QrKyDKCwynJThFl4zom4oGhnvl8G2+kNSYgL7CFSeQ/gi31BRlb1+WMSC
Yn2NHCHA1v+XF6dsvsecGlrJedSYT56IxVDMMkS++ei4mkp3V3k4mJgH+TXd2HpTv4SWaaxETjkX
+uP00I3A6U4wp9UnXAWBvXG8EXSjIskMWCwh+YZFa3ZvjEhPMEyhF5f/YqaEdImYP2/vZ7OmmUKP
ieXhUb4aLxOtYGxt2bwCydf0NU2ZRpmwwFSBdYsNZ8L0IAlaCINQNqbWQVJvuck7mXJLk4P94EvI
nAjdDtAn6sVHRF5LYxmfH0/ONmzxQUMRxcMLFNmPmnq72g4HAPIEbisW2cgBvwPOSNzUWCm6CaVG
9ezNVOb5cNQgjygQipIbBfTE7ipeiAVHUY+e0c0kpkarfqTpb3xjOJGfn357qsTS81wITD7ymf42
Mn0QQqZwlAUs7fT6WdP+TQkGU0X3qQFj5r7LMVPRkT1jwYlCSFtPxA5Vc+1odpop2F+lFzQr6PvZ
ythuG93lVqJAmchGP6t9XjVA9h9dMxASrftdKHsd2OF9W3UUZcvYKC9N+YKmgLs4viczkk6k3BBv
04zbqfcPhf+UXIIP0deB9Prqyc3ehfkElOH1gIKXPVPzUn0aFkeB8ESSV6+MVw+6K6kQ0hBEhQUx
AJLSa6N3MketT9EhhJzVbLigZ5bQEuOV1uYCTTbW+4AsC8q1VDeCfVEu1z6f/0KuBDBbyzGO/ich
6jOP8SdiaudKL11QxIw3tlKCb4MJlfagNDkoFU+Izn88LVel+hiqyMF+UGkFNEjcIqD+4mQi7Zbh
X4pMpF3r5lwh+F/P8kUU26hvgeyxClJrOaSs8s1QwQxTBwDvKOSi7LoVbK5dzxQzG/YpVdUd9bYD
eUualoBXEsaXvncZnLYo0Qei7Kl89EMU/UUfUdDsClGA7cAS9sfk9g44knI1M+dsKxpf+rhTl3hG
jPeDrb3S5zm3TPIVny0ATMuuhfHgvLm4MsF7rTMq+yjQOzrzkF6olwIWWN9FNYgozV7oFMrizByL
lsaDyLC7YmBGZUS7kp3M5DGHMD6/lqv4MnPY+WR9IpIrGbNeU8vRKxgR2dXD6UqmvkSkJTWUBeb6
x/PKFYuS077jUEUsca4N0nYxoit7zZr/4YDJ0RctHFyKmaV/gY5KyPNEgO8gsUOnxT8lLLy/fq/h
mcwlp5l/Na3t8xK1drSuacqWBVnHb4X07tt6tzKhdj8AcMpY/uwrfSPd4UlTqM37FGTAVDfD+nCd
PBDnybsuozqsCdeSzJCPI+zVGVysZziwYVQ5G9hS0/doyNyc5eMViVZT1p1E5ehNFAlkz3A3V2o5
II2Ingw/Cuuqs7MVX2gJzIXN15pvn42cHjSqdzjJSVytoIjyj0tVDSkoFnauQD+72LQQoZ+aaId7
qgE1QCUGnGOp5gy3KE46swuPArX7CLSvfRWfc59A+m5RmpNeJaxz1cpmHVFvcJyQ5Sv6tP206xVY
vQrntnuDdYD40Cuwqf0R+cOsOW4tLe3HMBDBigHjYbP8i0r+HULfb4FDaNDs2QavFZetEVbaKkEJ
9mHFKybXL+hzot0VseaK3HZJxptSKkFDxNcdP2ZME4wxZAm2GfdMaN6tZ+G3POzwT5x2ylQqwFTo
vDIUWmpS8vkbpWygyx9NGcMzaYGj+wOevxb8uuZlLrDjz2DoRUYj+78OZ6/qTJBo1uQI6CiChWRA
k+9lWpAEH0Gpy5No7pafvIu4taBQA5XTTc2smcOGS4HS7a0zTW8WSh19X/JrvceyvAAma8drPOM3
eU+ML6jVYY3Lgb+Iv/uJCVc9nlRJHgA4eI1D/My4HF8WaUpD5NsivUEb9nQYwqxaEcL6sLrPkNRS
ok6D7UliaKUU/cmGLPgWVxZlhMOVHbjRf+ZH22WTek784dtTsU1mVl5130MXFrDHjPCNJiZRYRb3
sP3pTPJGuVxFk8GPfuI+CO3WLhpJUj7b1+3b4FlmIustrUYxHtH5sWVVr7IugS3/LxYynNVCsSiZ
Xc8NEC4Su679qLFzfmKgrFpcb0ufkKqITWhh/8eE2HmQuPj2CUfAMgW0L5CL+KyZDPOAJ6UrJOEF
g52TBMMbbLqX5VNc58OqrG+Bt8yaCKx5kgVNSeSCxcYTx8ZGYVfzIRtQphSHGWHmkfdjBOfxq8pZ
w64tfGya/Lnmm0u39SeVUYo8qqO4j5wLgT3ljRdqkhJZOwvMaAJ4i2/5duHj9O4VSZRcrnQ113Sb
5QGEHLnD7R8TwnZmeNKwyiKfMatXr30oKqqq+Ke05lFc2YRmlD60nGvASX+s/3TVuvsKDFgUjhD6
Ez1s9Q8HkAcdLaDg1NXV8UibftNMj7tYAHgHQ3aZ4swO8Gf998Yeyv+e0zJDCBvHC4t67bpOJwN1
GyZWWiwa4xMSifJrvySApbSiickYZk+ZjjRsiHST5xB1sVr6dRHaMLACMvQE+/PNoRNbWy17IZK5
7/jvdyDgXxN45CSNvjJcug3/wmduQ/nH09P5sAZOqjoEwcHulCZFG/PJo4gHwvQuV75FU0KjWrNA
hLvH9Rh+ILGAnZ4wDw1JDf/rMHKBHNg584LyhPRl58Lr8AlSHq6Lk99cmMxDsDwvrlZAqqLeNNZr
Quz9/GbF9Zu0Wuq4/Atr4IKFxfB/iw/l5o+GeJsGWzs8f3xcMGCv7nP7UaaTKbu6NjVwe0WRoiXR
CjAiswYZxeJ43XdycvygLTHhwThmB4zu+Nw6RRYPj3Zxy5NYZLJ7Dxzcly834p2k2L4TQY9oJKKW
0Q5RZu559dQIZYsAlnsqQjTpkhxNBpE33nvXpxdDbwqXmtdZ0c8UagllASUKww1aPWbSuhuTZyYE
mS+cYZjTMaiMqPljW1u9llg0cbFMkms2SHQnX4ZJMhQhjX7W3lfhNEHQG4+1LPEaO2rTsRACVIhR
59lEgqGr1KWyJy7nqFU6jfxtBtnzfJvuLceWckWx00SO79bR/KcZ51pY8uwsXKPbvwhiWUbNNImr
Lj3Oa6S4Zp5M1p5EPTy6sVTWINA2V3HtzMRntGWSBuz2+uDTq4+i0CloQyQpVROu6a9ysUesGlnN
7Fcr8uzE+XCCCfWELqR4pxpK2tk7sreu+WfY3OwpIip5btN4KRUJ5kZp/KK30vz1xjUgc3Wu10nv
te1S1cvThKo5ysHxffA5o62zf10sCoUE6TfxwPzSwLTMvfhhv3tbsrXPK0yJn09SrbWNlEbQ8/kW
EASnNC2gg8ZYz44Vk9lbTdqyPF5ra/8cXs1y7fZA6nBxMNzqLuHs47qd/8OSffAxedJh/242zdzN
yhDbZjoXAEyzYleynYKVKM+MREAt17s3PqgmKfgnjSxhFFGrgEs4U9IX54xDjSpOKgy9goWcxCa5
f8Lki4oToJ4CvHgTnhf6u0/j6WHY3Yc7l/I9fQ6LRm6Y3G16DaDXToqv0lioPVotOi2BfzyCwjOa
7lOKdnrisBW02Eql9tb63e6xUuzhS7TD2G5aiQkQMOdc6JRlvilZhMhuJG4c6UuI6lsbhh4Pl90x
maJqTnD+OHPeJuuXRHhrAo9RSEO3+NhpOoye3xPi1WFLhqsPbhOHcLu6G0cby1ZDlbT7XcJVyD6N
rwGoi2SOCjpvHCd8uW1Rip27FaNgAChBG8XiM6D5LvSDHYU2eCMGIcwfncUkUByDBqtzCdXDPRG9
lmz9kfK+dmDM4grLS14R+F8ZwzHpnOlvTpL7mr1uo0nWJ7g0szjuOLprk5gHN496eSx9+pFmGUSL
2cDWMBRVb2SK9K5aq7mTAujQ//lsEVKM6A6guQ2YH0Qz8jQgOOD0UbG6yTZ8vXab6RHSr/IbSzT4
f2ownsOYa2GLUK+197ENFYlfDr8Ghz+NWPI8YLvukX9H18HMEHJ8ju0/RHvYDFbTr2sbZyhZ8Wfi
FRBM5iY/efIB11KI5MkZg1Uql9XN1n6Tf7dIPRouD2TC5tO6cfVk0IAaKIIOureXQN5Moqi0A87q
M/jOEV0bp7oIWWWl+yweFQIwFKmFiiaow+UVI7U29K6SjvzlcUmiEraADV7WjmAMRbgM6MFyMg/t
CQtmS32ZPZvy3FVJpK95fd9s5Yowd9/ufKYouMUNy3ufAY8NznXSEqGgmxFjV2KZOyknXt4XpBll
IjHL+pExb8aWzsFH9C5H89wBZyiJAhnxnVKcVNzIci6ZJdEYBTKLb+ztzLQZ/FgKLwho3IGxb/cU
QaX3pg6DZMc7vuE/Eb/q2Ab9neEGfAT4IWx0Zzr3EPKE+OaQTDXcbixHKKmQAlWoZOo+SyWMTwSj
2SXVfRLrJDO25BDi+ZJGaFFEFuNNi9qPTERAdtVVLrCUm1XD07eDdF+l9SHJU9k/Y1c4tjBaBwaK
ncpb1Ea5lAjal7lfeWuK9eFsMd3LPwD0GDWZ+0pumzTwpmQMPnIbpOHsq2MEUf5ZYm6/1ZAQTLVn
cb2ZqgiVM3Vsk1bOCjANKmK481tkkqiajhniBX7JmaxOGcAaXEMCa2VuwlzNwOYay1OAtIr8W1A+
9FFmZzC7izA6vEaAcuNp+hBrbeV0d/jsecND5JZntZCrimtviiqxfSgWm2jPSUlmopdlZzCgJLgz
cxD5FKeQitN3IeVb8amWfQyq9BXz7/Z5QMWcqD+PAPbrjomgKsbDmHhEZ7UN5yMuYs3rAQM1TgNL
pxr0E7rVFhsht2hQlmAKuHomvcRKtMKnVtj709m5cVRd3jTRxGS5ck4C7k3brEFQMCqWxP1ArtaQ
VHOUu6O8l4Jhyl5mER+ThgbwexM+Ag92cHH1e+EY/7KTBXyJ3GU3DR1sXbFf94WCkiwlbc3lyI3L
GPQB8HPthLGCJx9yUNXKvAZJUXCV+xr2hlP6Yh1JkEpaHI9BQp2QNx+6ElpNsEfttSLu1enFYpo5
ZbEG6SHSv1mTt+XC2ZxoNFMR+lhSlY4qZkBabIb7BVl9dNb9NcdvBIdqLkuPCAMSzU3XqC8yFtzU
fPq3k+Ms0nVxE8ZA84iFSXF7cP+IHiU2UUmHE9SAhR+McREXL5t01k8TEWsCCYVSwjmDU/F7QQ+/
Q3WJ6yIuMPFwXjK7MulAL4D46vPbXSvJsP7CSOvmhtqhz7OHBA6Ac0kpeWM+VvBH0c9h+LRnxp3t
LwK1xP1lq9fb3a7cnIiPwN3M9u9zci1e89UAmQpR9Ze/lI8H/gilc03ko3o7riMhNw0/EobHp6UY
Tzwjp1r56EnSR1RfQQ1F2lFf+tTFKJ/nH8WABUch0NXD6iB2R2suaRM0q495ZxLI3EWDZq7pn4kf
/xdlhGIW28qs/AfkoCgBQAUUZgO0aOkXKBfZjzyAL+dbqM5r3S43GC/Zab/ybx8ckqbcE/6//hbx
iguzsHTah3TLOkm246TD8MT4yGccIZdIkx2g7JDgDh1bHn06xB1jmgokLkHXCAmwidA1zZcBFiYp
rS1GCoXHv7ouNDIZukVNUeTph9gJLoyRVTiofG2t7ZTfPAnJOrgygovsoOc3nZNzo5DFgqFXXgcC
SsAytPSs4vRK9+jvUif4Luhm/0Ou04PO6BNQSn4yvNmQcI1uCYz1h8EiI77saBqM0VeInFXeUPUZ
O1ZP/7ykRPfVPK0UR1SQv4uNB5SSYqemJGQjOG0JszzG/W/XtO9lHWBVCaSb5rIR67V0LfUa17ZE
WE1HM/NZd8l5XhMPua15QYJE3EBtRbgMPsn2MZJ1XVHzvA8WI3VaeJkaDLOvmS+JVuDmhCErx8vH
sqxhRo8cpkTJZ4IO/CMznTbP0FAVjFacxB2QRBdulxTwOSKIuBtaHUV43PxtcPOfP0LSU7GOzgdU
KeB/JdBkA7eRUCIkpUL5asxWEarIl4hDEdjFuTlOhnhT7lUgGRalxXrjmjIqWhcEAio5Srdspb/Z
iuSICFxRmaByg87phBlJhu4niu79jL38Gf3dOxVPIPk45uUlaSLEAqtJlNs6Z+v1KlHJIRvH70iY
6Ul73Jm8XAImOy0EjQPtZ3xPejZ2N79Pj83IKvH/28vGKY8h5XGyEM8qDw3F3AeytnJy63+0dhAx
SRPIzk4L9u/lMWrEDPZSJU63rmNWiVnr4qfEXIUw/9GfJgd2w46hTxUCNX5Lh22TxJg4vEwWO3HJ
10tIGEkvDHDaSdKK9uBAhbEwyDbpVpYxmpOkJo0Se4kpkeiot4hUAdPMuvEksH14b8oBksBXX+CI
ZV9/896av6+Q6FpkOilAhNpqi1E2nRRh4YUsv/UO79LGG5mVEH202JEnUt8mNtcqwbe7SGyLPDEQ
VDHv3fXCCdL7u/Rm+eQC/vA2Pxt4JMRzPaiXN9s4UhO6y2NRgd/idvYgUDDpsq8cNnC6X9FuvkkN
MSwV+XR3Kf72iPZ/bKvpxJsW4ksnSN7IFlRB8z6ed6d74jqqZXpiyUs+Dma9+sYzQ/xDgZnKFsqG
EE+jpCGLWLruAeeLJdHuPnGdA26Zal9xNqs4RwJFfuVUjZk6UJkDfTcrEA36100b4I5t8ruTm9eb
+JPnJKXxVxnsmjvyrVK5zur+tPIqw6JS5h7lfeJrhbdkl0H9ZhG3v3elAN2TeaVKZwMcw6XwaCNX
5Rjb0ACujb9Y056MFtCOsKZL6xUmGs4KqfEbitczCn9+7W5PfMKavfkPPOLCoK7so2M3eIK33nLG
GeeT1CVuBNEXF+OrXSF8217Jf4sdLFUNEGC2zNRuSksF7oughZ2wRKYW2CFm6mQFOJYApddLm7pT
RBEYj94LGvoWj5VUGUTTKvPeCqKK/QwrKf9YH6RugFPpUdAaU4W0e+m/jum2qCYBVD4RIZ49a8Ky
4zb2/SVOGixX6LVFmRw8t2NXThUNxpv7u7V+/ZYp6fjDEIwi7T8oPxpkM5b0koOLVpTFLtN7KyOH
JNL/80/KB8YLUe5eyWR/egsPis3GQOHufdI00tafrsdXxLvf3pgGZi9cYcAMeiqFvU2nK7PPyh7u
tQ8IgBjXaIg5eaP4ryuRcx5IOz8lPPEMfXRl4GW7WrtY5fqR+Au5CEpsDKdunQr7Ob7ineX8k8rk
IZhSiJjnJr9jFm4JbUq6V5I4AVx/IY2GJJt6YlWRX2ej4WzrEFqF+DUEsZAhiorgrdU51tDAeOLO
ACtOhnjI6ITJgwL5s9XBkROzAY6VG85nyaodGsCPfebDCnL43k3UJO3679Fsmsl/fDQTdDTuC4Tf
DugImspCg4ghCorZGP5rDnXmW5G5HmAbljd78cjBFD0OvnJAXq2gj4FO7NfVuJRpMEz1Jepy05hY
NjLFcohkVPtOt4E4hmg/O5L0Uu8sor4cAcp5bLs5uYBAIGp7jKAFFzWe7Qs1HiU4jd97l5X3Ov7k
35Ljawg442eOq368WCQgZuyo0GaA+41QXgQCPEqsqZVgoz/jh+jcAcv96UFs15ajGtdav4Audlk8
FmK/ZR+Fi7KlMJFOUacmhXP30sEoHfEgxn652FVGc1/PIfkFuIMju8pZdsuNgYR8QzIekZl5b5c0
uKvq5K7fcj8HLLozaO8vYoo9Mzk9onnPKasllqBPrzjA79Dizbj6drEDWC/3bh2Zai8HVTRaxZnq
h+ofQ/lvFctKl7kWpZyFY2TsxdUj7IIHpYILd6qc4HWuCQT0sqiz4wQPSrpV06m8Aq2wc8LGMggc
gk4ozmSFqbb3dS1ZSxTX76D0IImWV0ICU2thrNPkigJQAbU9aYjrtCGTbTMnvPw/WdOqWTG0ekfS
Ri+ZsGE8wfsXdFdSVRwNvetuJaboZfQj7FWxH8pTvQ+/rH6nm9p7/VrKtXBEm8AJVkYevvZYtzCg
+w1oSA/Q7w+8FTt3/JhqQT8/IKMHGTv1BtX9ff1qHuZOG0VyOW8G3tP8UPkWoLHOGBxOklLjE3m4
zKfPl2AANdj9K7aUs2Dpl90tq47l8Gqj9nclTitFqnWYCUmwatoULAieQyhh7y0vaD/OuHqiAjI9
1gkH1khdA1HUU7OFmde1cTBPrHFdVnDW18NXq5sOqciNluSf+zTF5aaejWfslKKAWV6zXtwopK+q
TIClpAY/ke5AJGqaBoIzgCknINoA7eld7z7nPpbtVL8kwoMpZtPX8W/DV85FHLbQBBkZxosrsBPl
Aehtx+UQaeH5dUnXH0R8jDr5i6Nl+JvTHcBOE47NLNM3ZqIdHOeRWvhAnYzes+KUijEtK0Wswovi
KQt9ilNOyl2lPaQEIOMZ8I05EZ8vuUKUVpQqAqvhqvGJyxKR+wtd9tYM24txkFrNF0ggd46F7whw
jFLcpRvTP7ztjaunWTtS+Ud3Aob7zGu1Y0Xo8ud64cdmSiySJCDmgwpahkTSTIiXjwHDWcE6d8BS
MyuqrxNFDurqJFUEZlKE6kxk9JCrJzKrW6w7Dfy8GhInBQRXL8kLs7OtcQsB+lZ6TBGZBIyQG0EA
v+97qQvIU78Takkr44FQ287hg6bw3l7zk7+xWn4krLLJ8wXWAz4/OPyjXUX3EN6TSOabuiqxZ3HM
64l8RivuyYtuO7dKdF6Nqk2NcsOm4P4PjdXEPvqfVP2oC/LEBbRgqNkKaL+QlMlg5aw8zstnHvHH
H0nBhJfWIZLda2HSP+vJNI1rbuRzFYOhllyjcCSXoj1XfjkVK651wwFq3Ao162RyNPQQXz+/BASU
h3rmedrRLOGVkPmi5AvbadQibUJgZPTmh6PiN6zgAM+NkdEW0Wox3zpUQgjlCC8JudxjyfJM47BB
LrXCIA/7VyaGRI6yER+X2znDzWm/Rn/E9hKB8Gza4oIXYl4Ji5Tu4rAOiFiq7pYWTXkmxG9jiGm1
3me2Iyuj42OHwdtMb6OBFNWEjehLROk7RmzBVKY9G91lTYX7vzIuaW0fcQXSakWzK5eFRSvAYnx2
e1XJvyEgw5nSRiisC+mTqBKGZg9kMK+CXmDM5+lCNn25Wo/NC2LHS5hI1Q609k7g3Sd8RtKFu51b
Bl+1FrxHBmZbUL21OKqJDk11czvLCSGMfAsTTaOMN2NmM5CfCqGvm8BFo+DQEY0aHfZNk8EtKgXf
uo9RhyrUbE0WAyLQpwLWyHWGcVbYdAZn6Zd77jraw4P/f/k6lkwYJu7JRimadX8Y74axnCxAlldj
8kmGygUjFtW8HMLD6Ix7GtTsKMMmgFkFU2alB8ldmZ8mebwUkfFkRBIWkiem/94jY1Ge0mUZAqPr
tWan6QD6xzMiBtYD8tc97ZGeRH10huMUaW1puXJxtwg3eO4SqQ/Bxw04CsmYVlifSiMUa25wO0KH
4Mx+B/7U2LeIDE7ac7RE9jEi847a4zjk2Pos2mvK7HwryHX0H7i02CLBSe5Mj1KJEQiF2hSGKnSC
CoaTDbouXBvUQUgLKV+4Kp0QcQBekpqs3pS+aYD4d+ezYpf35LOlQ3VwqTG8Saz64AYfsFN9rosd
15bMCXsmEbVuCVZip98WpfXrXzenzW2BDafbvpRnb8P3k5Sw86EG0PMM+RoPnUYcChhC6WSnRfRR
/ABtxjwBgLvTRxsvoi+d5ppQzXKHqCF8Y42LGAIk637mSyOl8Myw/k+kksvnYLHbl0ICkRszsHHB
fbf/FQWi9E+pQkjy6H9RNW2g9uoZI3j/N5qE+BkdL8GFr4K06G7MFxWtHqnotc4IpiUBT3iimPoJ
OCMEJHKfFeTtQ49rJzPevDbOE5+vwVJVXsGMbPpcnktRC972ZVeV3NJxgA2G8pRdfFqm9eqmIqsR
v8C9IpulIvbUWgVmwsViQ7EQ9pIyW0puyFZ8Of7TRqNbE+exofmo4rnHjBZXqBCF4Dd7xeuxYnXI
UVJafO2+Lav7TF+NyyrXmDE/rBmqi1ex2t6AzJfd0lMpa5HYOjVoykZUvASldyGxDyKfh5LaUb6M
we4/xGD8Q9IpKsCxeYt7KaWlA1ljLGPPYuRe1WnzjgBZg4LMqDYbBU+3bvGpYso2TRKkdIU692IG
6gMLh6l0GLsKxYyc8HAXKMFV4ZzB/6/cxwZqOM5n4IVicJrFXvcWXZ5qs9KOo1uVToUJOZcL7RG7
Dt3WfAwhodsGUelGR2zqXJxb/vamlNNAjCgoUAVgsLbuvgi+keWSaqyZhL5aB+o+2yamC0snL6pw
FIkmb6Uaj8217c2VvTw1yj5uzgb//eubUuKyjaLRT4+GYv88MeUn3wUxQ6gdFzrOP3bCXN9kFtlg
ceWIkVmynzk8Cw2ZUkJt2ypGDQwlsCeyK2aQF5Y61z+C5d/P1seD7L98Hx77yp3VhnxpkfO7WRVv
vowN3dVh2CtuSrNjHmDSdGUgBDJs8piUCCZSZrKeP5dzPOQZG+AxkevcPxnbK3lKYquxTEPFtRNe
pQuaAdPQa/oxZCP3v62Ng72wm3/T++nzSfLQOtBYCN2VR0GRbYMtJ2Dyqw0+8ebi4ILyPiplENku
WnJaBq5QnU+RRaPmjO8EOLRvEr9z+9U8oljV6bgAMANZMi1/aprLWwVLXV3GUCbUDd+DT+2NSi+a
NNZLBtvo6AK+DsPo4hyDQjiLpyH10qkuiHaovsuH/efgeNNXqCPgJfPkeDl/BJa60roP9yPHwAZl
XXOd8RRh1BoKtfv4C4lzMwj4ADKUJX5ch2jY5AU8H0zY+i0ZJhqQbt1hn2/mJemmP4QL+nKrGd7H
Jsa5g5R+9TpwJbNju+Aym7y6zgXntyBukoOdLOjKBWO8lF0nHPKrJ5piyQ5GGmfnVR67Aaud1TyO
LnSfr7UwLQHyJ6KxqCSxjn/Aq4OP2YaYiESRIRsy0QRaSmfI3hAAmJB8w4LTJgHaRrhDE5dLKxKz
BPI+Yy9cd5Cj/FqsvGC2/qBI+9044t06E0Xhhc/MiJqr/Rm/c7IPE0XnqBgHdGz5ZOH0Jwab437I
WMFIogO4kRaLZx8hfYdXY6k4a/n9/dRZvBZtyl2T5LD9BPvC92WJyM8loTlT4tEwWCvXbCv4xv4+
bKBTw9DM/xTwa6J3qr+X5WSxow7tSbjzmzQOxQiWWi/Rze9Xb3ZXUR3KRMpBMiIkUnn0NQ1JlTgw
/9ftWGm5bXJapO53UnDHQN3Q2JolMWjdB0PIi+q9zbt0xWea0LTAkYW62hppASHl9mrsxgk0oHQ3
trxhAF6peye1IDosf/Rw3V+HEaMqNxn9iHhx2nae80CxVqI97hzaTe4Mqswc+6QoDT8fVDQJvogF
yfa29ly1M2AWH7taHuw9FN37IexHwvd0wUnTk2kPKcfCe5f3xoV8k4OxVo/MsFq6DYKOH60pTvVt
kM3R9zbzd/J9uFbB5R2KOkmAJgqvP2XAZG05F0mgezlZFC4/V8qwn70YMjtobQXuC44SGpnC3yzX
kuR6SJC+MppRlci1lrUUFPcu3Cpu39OblvO0zCUOZNY/d7DGuUH8AxdXze7YPYGnBJJWxNvPUA1l
Id+yTqzxC73yz1swY2/p8byToL8uCSWUdBmbwQKOotpyZPBBhRGZfiKO2ZrcLN/J4JsM0+LYeDPh
9ZGFNb3+pnYvy9WwC8vPFq03HWMDAu9AveZnAP15hqtdTrmRo/ZehtAYxUjX1512DSGaxEaPkwID
LzR0Y8q1QFGXgyPl4YaXcY3quaZWWYp+xe1IZSsrDITlLnNi0s62CTxcV1vVlYVZJxj8/nDSsVJA
q8w5pH8GfHrS0z2sspAR8rOem3d5W/AjqvVbCwKcz0w465lqZpV1r+Niid3weAbRDr7BLBTjIOoi
mqMdZLJ+1CVWPw0eucmm0NO6GryFjwxf+u31BFAZV4EezQbTjwVq4/4WExfZpcZEi67Xp+hEQgP0
UEzl+Jh3fwXKNXEye4zW5qnApIwTwN6kO/YY7LQ1b8V8j/WfZaaPU6+VHRkm7P5/feeJByzKPboi
hS1Gvla6kqIiSripxaQ3IWxBZQM2LymVd2C1hYgIdPKhCqIlSQ9kiJX3/5K8VgSk30nR8QDDRhYJ
hizfpijdCUNjNHFWCu/Q90e0gSZWb6e1xiX6mjOnUPVYk6+/XyEwsJd9j/0feYePvxwa+1t40uU9
+DnJAs3ofPum/9ICNZOSA4XKbiASdjSEAYWzNFqgaPPOUhRDJ/r7J0B0g+2OGkYLTNCvIPjVldVe
ZZq9PZis/cxXtyQwGRBmx+d2klGuhXFBtZxwldWDIWtn+3VBZMmsRaWZ+3p+miqQtW1gtMMaLQbU
ULUipNw2CzeFnd5Jq4z+9Edp5miyrLL8HmCGJdUX4rRGlhggl68AXH1CdF/VUOc6UwY0RGn3aoU/
KLhxywPQuYNlGOeYVf5u+rJMvlMWd6alAv5mX41sCv6Yw5yzmLWgskX8k3Ek/YzX3bLGT7Kfnn1I
ZbD9tHu/iZM1QNxqC+46tnAovA6Sm4Q7P9qNTyjl1yxgQc85aDxZ9OBiWA+qdI4hKMngRPIXgNLf
pN0KDl/ZM3yYUjtok8rsUmkypwK0Ppym4emLz5LSYl95IIGZaD1IUTbH7mC6izYVki8anJueAODb
awkHlTlpzTXnKScwVsVIYhHwq9L7ktqM0jWsEdeMEVjPHcCvt7ZPZGFRV1QcXylSgkee1VxeuV40
bjeWiKRutuowI/MZRRJi1n0qJ3pvUUchP5o6eiRwoyUf7nygRjwb6SvnhvNxG5mHrfHA9NJued3n
vCWZ8fNReZIVjUi5muIGag8V4TU0FKEK/Nt8y8PvvvydXVz1Fj3d9dM0VKHVYI4lzH/YgDv3Dguv
jw5o+SQ5nYcHJ7FwA7EJArxkxKD1mjL+ThhAEZLTMKgGyCQ/DgarBr3hDLNc32U1zAqt1RfAToGU
dLWvi+eN1Zf87dnpckF0xKAKslaF9bbFuVYneCMhfdd0b9OZCeO2oViecEDJLCz1enIxa9pzyguW
3h2nGvrGSBI9Kwu/iqPDyR0OyZyagSThfu79clvs6wmwLDqYTjcitf9fnT0Q7iN2/Goa3oAExXfa
b4jTMbo/4RXMVN9nrvLUYHJgLo/NaawWXlxJ7/SUhq4shi/RnorTuqsi4Doastmo83KXIsx9XERK
zNU+z32kr8MEZ0eEDv1u4Og3HovCh6Zw9rnoFZ1d0gb0DV5Qtt/qknjN8Pm3BstUCpmzEJaMl8JF
XwFzjNkhRu7yuvKIBqAd3lb4Q3FP6osmJokKDGlTi6qsxxZgdZQqcmPfdwf7UCiLlqQug6PEKaGV
tc/j1bNhPN4LrmxO/E6SEmYrzOEw/pzIyD5XSfdN4BOmdIn9SCDsATzAPytnye0GR5Rjnm3VvKwa
FuXgSfM8qJSYKT9TsllcYiI83Jch9TkDMO7xLpHlIO8E7ic9P2bUCs3rEoscUvtNV/WR18O5ipF3
dOWn0HZIuZbdMS8kfZP/lLb3eXgalt3uiZFVEVJAiHXKrZO4As5UFPhWWqq6vn9Tby5W+oRZPztw
HvdwHu8Ogqh6fBpW9QF5CIfxnSsbKmCt0rrmusr+AGjknFv+whNG7pOoyq3OJRfc5iva8zNs2bid
yKauytgKGXUZHRFIdWMsJ6KKmt6rSnMKfucKP/OuH4IhVznGW1xTta4ODOtqQY4ijmLkxMS1tc9q
oBQfFbW6YqcytEe92TzbMKYFwRvFprnaXSdkIEhE5J8cjpzAGUXKsa22pz6NUqmZHDL4uRxf8zvn
G6e2I9N8O3mnr2ycWcR2+2QdSCoGAYrEwnn1wJkFgWyAGbSlBc9qb4lxvO4GnyHPz9p0lxRahl+v
i21bMW5ORf8bbMUtteTRrnJ0mkU0WDskhrKPfKEh4Yo4EC3VDZMrqt/9RvHzzb+UoAnNuc3L9sgr
OUVbxgp0aNNRLLE3UiKXk9JNnH1rVWzMCInE0npQh0UiXvqCvXLsDhAxFcSZcwx308dC8WpjH5Td
cMwHK/VNWKWrnE7AHdh95uudsMYdwcc1KxuUyyGDpHAjfDxy937VPS+Iz7eVwVHePxgWp2aXS+iI
Aw8RO5aphOMqrfDEYlbXygJqstSC77qa2YbKE9Q0H65OMq1V8XaIdznsEOJBhjkAhJERasEZBPpV
JL7KezG9EPW7rdwzIJQz3UnOQErCU6qpXAYkf/1Vp070NMyRDFMuMDVySZ+nvTmMkj+KsYLhREYL
Bxb8cCyYEVL4ficIVpfvhUQJ/3eoTlulq+tkTwaPvGHtADqI1StwemtjeRflq5rE2N8ftXloaK4r
P76lyFxCHcX6U5YLpmfnCX+ImfNvl1j+3ugg3Nw7KX1trwmITfVxyw47mepialLWvq2YNVK2s3x+
2QqiMeYx3HicqSXYk2+OFUnHl0wy63ANbiixU/HM+ACLAfDvw8qfT/qdWyKFHm1HqganBxl80n1m
n/Py9gZwU873jEcjR9mUV5nUcvMF2Dpin6JwD458eo4S0IGDCNEY1DM7N4TmcIz9yReO2/ECoCcw
/7wVKEF66in8wdYysaVxQFfhsSqexLb8JIN3+m7Jz+g1k37+TXehqCefETV7FHiiYGhUh8agzTM9
aZK0Da9UVvD7/4uEueYp1p2cy3/HhmnSXUhPrK5MJrI050FNecinlC8WkSPR84o2/jvD3FUYI/OK
UV222LRox3PG1lfmc1eQgezO1Z0Kz8KlKTnD3oJqrCs73r109vpl334nCpfflqebsYa1Ymetssft
63dMlXc6R6wZJYIxQhZQxGwLi7LrhuCYdnH+240efUIASj3URcSMnZGl4HeOx6XWyqebhuzInQuu
kzODIREhv8Bu4ZS37RK2O9l3a/FXRPtZFFjmKo2B8yrbLNAv/f8pt7pVi4dGqZJSm0pEB7DWqYN1
+jYfQtpLT2IsxWDrCiw99Mah+F6imtwy3MsD4DPtZhoa8RYOJ/KeSUnJSy923xdXd/xkro1DaIaS
KAefBXQwhaTLNc+gFsxyVpWpp4hZIhjMKbeiIlvA0wlUvlIOwXfGeoZeIBFi24GHi3BKiPFWw7ar
iHtEAvS2+X2M8x4MsXmCGxk3vGriHLTBOU2f+x+3iuLIQOL2n7gtzrkoveY2HUeBRmnQEM77Zv/v
0rzt9Kaa6Sc7zg6c4YFRj5n317BCdv7VMZlnndgRDYuSyH9O/LEsM0ykd9w5mWVmd4ki7E2WgP69
BgW4ILdOShrHlQuI4RSPZYYsPPUdrN0CL4jbvWwjkhhkvw/WAWbyZIvU1fc05f362u7aU0bXMw/q
WothM/ntnar+BAflc16K6SO1nqJJizVPDe+rB5FPYcESm9DhZjs0w+UT50Q2uzMMLay33Y+8vsky
udvSd7xxaQF5jM0sFedE6g7Vt8JWbFwCZLosqTvd6gJ8QNe4HqtLlPuO3lMM4t66N7pm4IuyfXlh
4eJ4/n3coh89g+7jnGcWJY2rPLnikmzpyjjo91cmUFn3DNkV1vQgtofX57VZHwh612YSMCRUQJDy
J4bTtyUi06xnsdmSGaf/mdPmvIKOSUXhi0e7cerVigtAAPsdV3rNXzp3AFHCz2W2mhJ3XUSHnj3S
cdonuebwBhmJc3XY+Jjjs489n9gNuuADdbuievwkASl/lSH5P2zHJ2/hg4Spb3FB1+F5cwsmZkdv
lqopRokTRuu7ZwB3AV0s1/+44pqzBCrmjJe/x797c/0A2LqPHnoST8R9ZgRsZqY3/eYcDQ3jIDpb
2e4CAF/I2c2Kr2zUltY+1r1I2RjBAwJBlAB/13PmzTynYc0DsjhXng45zRUNcGwINpvs17bF8Gwe
jKmtNuP8aQTZpp/R4zfDRSXYmxKNEtjQxN5qHnGyFgAavdtsOEJ6hHh8SyYcXmJ4km2Zl9Q+7ZDt
580P0A5wAE4odBM5bk9Y2nzexnxI4j9oJFYdyMhcciD+o9mOhlW9bqYZdaE+ivnVu2ESm0Xr07iA
teKJ96+pOQKiQXr3OU5UFJqO8FOQ5kc7nM8rxrfu0XxtgyQVUKsn4KDprSoF+TeUh18KPpHd3j9Q
4e9UU3DiciRD7VK2bYprp43nqmUvho+Oe80TrtQjOt6esoVbwyNaGnvCeX/A1DE0/56J3p9XmV0d
H9C8eTjnQcyQAJOj/h+/nC588J/rXmvRWyvArJDrdczHS+O8MQKd2qqiD7VbYLjMOKWhMOeRZVoq
gtw+R5s/iqdHEJ2Laa2Xvc4fnao0q8HeHxvZ6Kh8WAqjxwU4IKOWU41USNktj3DuEuz2ovgopKg7
1YgT0rQycUfQTmik3NP+66821HmbRnA7UwD2IReAGK2Nx+zexFpKAaFdYLm0/f+skq0c30M6evLl
X+CVky8JL7nhEDfGQurBEKWb7ap3NzQzQfEW66mnhb8aM0Fyd2LQ96a0MYjZxUFmczPZCE3Q/uOe
ocBqVBtpEF6dEqIU7J1M9dXBjuDK71SyuuvO5CPi0R+6Tc2gwWmzXxSgKKOQtwDk9sAc5hOetDBj
MAgE26B6BoX/LbmKc2Kg+7XrXzpj2iRwx5t5t0WLTwzZ/YUZuXUvYCwJDydVA+n4oEwnV+ksahx8
NWBmW8keqkYuqyeagBD0TyyYiK/jlVa0da2AO4rdUd9gjhs6hH4Rlvb+CxiA6QjCwJ8wboOxv4vC
jxPvcgIJY77FhHrf743d9zYYzM5pQh9yLUHWd8zJWmwT3aMSwFqP1LtfPLUBEnN4UcgmX21gxPna
hGmb9a780y2XAMJhwNt2dF2LwJPmwhHblSXJAG9kzsB8Gbru5bj2MtP+Eh/V9Aktu4svYe+2CSCK
B090/f/Qhd+GCTQcVxS2q/BD5EZaITDkzr9zshIe0Uc7DgOA52gAD2rKzngFdO5XeIJMrLQvzg5f
7fZMlPuG0AOOAbo2T2RkhMmv3BXL40T/t0SwfbDsgI73/bzXmK2n8RLkT56qEDJH/veNhy0W/+UC
ky9rGn1l7ge8usHJWz3j5erhbpJiNsNzJ6e2P7OfbXaET/48tnHUGYEItorWKPsJXROfAtgUG49a
ziwfq9iESugtGJTpxJ0+LJl3R8q2p9WtFViczTyMqOQwz3qSCdQTiJaOa0vTilGYOmYuYXHtb+Gr
nt5ChNojsHpSHmm/fhCCKokTAuQNBLuZzDZP/61/fVPLlfK1UINgpescrEzX5asig3/Dh8uSSJnh
/s51zyR6MZ8qBVQ6Fq2fmsqa+OCQ+K6+ntpgOGzKY2U9F9hBIc42j8lkBHzztLJpKKwXLKy0fqy4
w0m5oZlF4WQH5w4+2xkQIWXgisjVox1M/93D/o635uCQfehHxsNcjUK1xYVBmowjxOtU7jWx7Hrs
TfvyFPNdMzTeQm+SAY8ZmL2OBFvoqTtsKJ402UFtND/Jnka8qaZln/Os55S6kTF/43eDZ7Opr3s8
1vmDl2P6APSuGTZgCn3Fn82Jc7+qciTkLaxdLY9GigTOPVi/s8nOvARun3nDjPXnjCksV4nHWvyE
iXZwd+xLXUsLm/KCgpFFmp6BOfL5dnp4jPi2tREVeDuT7Nn4uBBSfalxp/eNbjnmT8mVfSHQqEsM
ksOLKnRp1RDlqpiREmFHtWxSYaN5qYMJF1OeIbIcPo8eGeTuS4KLtR9YqE+EXwA6Hgoot6JtJ9Wu
6aCX9MBrlWDzC/Dza0+zqod1OKpEtqqsO3ED+ZsY9fd9PKfoJ4/1kBOfGCATw2bZp1itbh54oByd
pzGUfCcedffQnEvqktR+ygT946TX/op2qPNo5iXkZT0v+bYLSUWpVploccKm6vFacNi9GjxbN/+a
IFmv7uFD6IzV0YZNJgHkKF35HdTownNJAOOX1ums+ISKYBqWwNcSmWZg482H4vSmKi/J4wR2ERHb
70hggXr8/5y8/Msz9BHRJV+4IZD+eOHZCockjWcm/9FC3KNuzMoJTIzfcH/1oP9yX91beoBpS2E7
l0Bgc2snQnXBjtoCTDrvZRZCyQldAosq5DaVq8HGJ2dOCY1cart5ds8fNJHrZHm8Xtk53flGQTj/
PTw750/aKAD8lZdRBXcXk2oxAMt6ty1ZIAwtibGqm8nBEF8DuxFM+/SVvImLEdNf7zl7/w+2JDfy
8tZqMo2+DRc5oVReK19q2q1zRvUJT3HmCxJa1BbAvIgbqorRGil0UXUW+Q+Htgk4i3WEsV1mi7rW
5VNv2JsyTySfU9gBjGeobPLs+S1u20HKkrlIXaR22WEsJmVGplHMpr9BDMp8++Oadt+bW9uCz9m6
RugUKbJ9U4DdEAv0Ee5X1fiWJhc/PDZQRZ7vZ6k1+yfZM6DxevE6w86CDllnJRVHQxqYnAfWS+6F
ugTB7pfq5S0j93bFVQxfUGvypOw2gjVNQ9YC5ryeMDXbTsTXeXbadHMWEKvc5HvfmaJAQtJIhe7j
KKlGdgVZGh/uSqqZO+lqzURSyGrFxeHUcD8sqfXLZIK/UkRjjGLxoU0JOQc45JtMoAowJCJSqade
GPfBsKP4LsS/io/ajGMgYqBzfu/qenxJD+DxpRbn6n5ZlSNsugCG/y8jzRLzo/kJZ1QYLTfuzeBH
F2eGYaWCnfsm+SbWDT2UIw/tVB9Z1Aq7/02MaQM+uYJwE1APKSBn7ZY7Nf/L/iuPgikUQjnN3GbM
AZzOvEl0HqD84PFLTIWhXv/3P9+Bw6nYCA/Orhocg2/zsvyuZOQ4h1lNMw3mX8O0FOunC3wpKV3Z
cWHl5ajhSTEEmUEBG5dI1eh2WRLwDepnIeTdS4yOfGx9l3xXU5rUU9we1GXhENJuvCKDgdBUYzfb
xTDkcNwWhKJ3hG5uryjbFb/reaoWWufUynyw7IOWR0k5wlDMgHgQrbLrTeXTycqIwoUW66QYG8KH
LjbQqrB4YFVk8e3MVZgU73zqhAzjNn1mAFjIl5n+K/vWXEUcGv2JnrhdrKoIg/oIpg1tOCq+A76p
suE765Th1yC49lQ2IIJvlKFtXCScYODx/th9TjXlUNikpKxift++aBHIhCLErn0QFVl9G55cdA9/
rMhpePGD5g6/aipycaeYevncUOgXeqFV+HjqB52BCtqk3AyBqbszpzHGoJ6lKk44w0/EZ9Zj00yN
fxtyKQ+RnO0baaB6w/exkYYEjScjpVv+NYVlVCpZzi+pWEML/U+HxjYZuXCfphTVIkuNUzFZ0rJ0
piuBFBNgc2M0zosqHgABfMk7JDiZMiZv046q3EH0yhAEqUg1S86gX95RK71JQsnTMj8nzotB0mlC
B/JOQBG/STzdWMpJGMeIgqRXdbQ4yw7eGg+hRlN8BMoATi0FzAAQ9J/tmzF53KA7r1AWQF5TGzMc
BGwQoNBmKDV8WFDSSjq8gZPWM+y+SXyJB3tRbqKgSInlTxazgBszVoLPyP+dhxSW15TT2ann+qo6
G+kufnmd2cwcBg/Au8L02yd1xEDu0qRTMVWy2pfpqHOzlIh6ieHC7gPU0HnWQJdxTUgup2cDUm2F
URlQrtTfjtdetpnsEOawzNpxtSJE31i0JIoKs0RVRRGQiczdbqfGq5FIvSWzZAli0WtgeUzRl6cY
4uEaKo2tTJhQUQG85NpmNRP4nXxBUlyxonAqg4pYWo9EzJzYQ3kvp101mO8a1Ff1gLTPh3p6Jk//
fiFqzLtoo03LqMDKbki2tpXb99aXFnUOuRRBEJix9H/ommYqqC08eK93W8xSs1FtifFVq/0afjcO
YXQtJnfr8HyB+FRI9xvM48vrXoicpzBvsD87lG+9BHJrekIaVRMFW5ggdxhLPeNDO+LsIQUI5aXh
xbNNAewSQVzsUWzkvALfk3F4TXia33VtXqJiPZ5lf/yipz9TFgOmyVDZBVelEE+xb4BU84RcRlO9
4tcxcc1qqG6xOcB2XSuKxXl7FTwGV62fkLvt3i5zkZze45Psh3A8pnlNqzsTfDs5zsfibVAuSLF7
Wj625N0sKyz5Gdqu9NZPErwda7DJfsPBjCCwJFvyawZHdMV5WSvUdDXor2jhaAk3jcV5yPhNyBLO
rryeErtpcFqhM8g/QHuOvM9B2gmplMk/AiSlsOBWs9pvVVsA149pvFa3d9fyTtcJI3YZyUkmfiFh
gVyLIapwTfSA0uSygAfUw58mwEmEIKlAonmaM6ZtlFsvfAND1oTR9XByqPy9oSYIeVNefUGA+4uy
oq8DAgqO4rnyvcLEvZTEPuVOCxo5MtPQmW/cGNxbB/4forLhQN8vexVUV8wdzg6/y6YdE3pG97Z0
dI/tyC4fAPEBKfxxd0tXrlripciy0HGJk/j7bpYQ0/8SQQ7FPiJea5+v8QHZaS5COAnWzFSiZkbf
wnIoLEM8a9PipC3fQW7nGM2Q0ISqhyOry4GjI8qVNj9QFFGllwsWfui/PsgXWiyHLNJvvyTvQAX4
AKfl7z+E9KESZpJ/Un705ZGNQde7xN/ncTE4sYFs6DnPfFOxdqNjpPt982LISxEDMn6ecBsg1Od6
7Hw14wsgBj2/TJuPO0qWaQehQlSIuUznNVaTX4LYgr/d75S4wlH11B7X+KyN3YMDSqIuvmq/zoMh
DZaO41YeZFXgPDVMyLPH647iG4n9EPVCSTIu7B4rOFAD0BK5Ho8OjxYPTJHtsx1sGybObq2yJORG
32QtEyHX2MUyM6WRRBhUon92+6cNts9jPuxaONRoDTDbo3na/NXyVv40Gw9KxlcTs3WoJifl/TkR
XKLldj/zZrECWi4c/TzN1b+cZbYpwK0dg2PZn5e1/s8uT5bXefC9NhldIDfKT/F+FHqiIxPCS9Oi
/venqTwXSxzqzHq6TmaiLXj1xIPz8m/oy2l5gmNsc+Wp2zq/s2oKCjekgzmSBIQtWAEvdOxQCtlF
7FvPWjzsiPuRbb0w1gtdM/Q3c2wMjDBbpK/eSy+yrIzU5U4jrtKr8ul2Tu6y6+28ZfPSEZOZFmDD
ccVfa0Fhss8bYKALbLQ1noyy+aoUd+uWf8ueTMzsCwaJnYDreQAzI4sJJJuffuUKP0/mbvP+Vq/O
IdWI8QHKwElcpgRnw9OrWYJ4Wuy/VIjyoY/FJ4aqhW7t3A4ByNJ1d85skfQ+Vz6p1ZfFkyj+0ctt
o/QiBK1dC92y1Ot6BvlZpLtc90K/EBMADA3VyHEREhyQ4iY+CWfhX1UstbXWyYR3gG9qBXF2NtBf
8pj/RjQu3ZVVG9Vg2iATf0/V1GbEMMWGtUowWupSDd+73BSBAK/2GmDap1Om4b9vh+b/470/FQXz
wM8++GRELb4ktOlqSxaCl99Ms5wkGvO1hTeMyhGTv3tb1Ba14TMj+6zYn1dsMgpO2oj8tNxjdaSU
smuhxMK7uvcJHc+2v3xa3KiBY2evrJiPuGYH9uo6ZyZypfcnsbKZslDXmpF2uFkKEZ9hwL7vfbHR
De3x6T1ec0yqpSriQ2GVgR+dqE9DMem2XciUy+XoV59C1MXPTyubxD+WE5E/qXSEE5/JpaMBhwrc
6ctRY3fa/QyOWjjSKXkOmkGVgOf9P6GIbD0RYSbNr4Quo05eS3Gyu8jibAFila4JkqOFcYs2B+fs
oOVAVy2KusU9D9F+x6qutwOSPZ7EV1wbYN1AEECrCHATrrFODdU9sKq6XmJbTf/b49WrZL7ne8l7
x55dE56h1uhlqgYkNxGNdime/EgR3ZL1HmCr5BXbUcqEVQX7eBgNCWxGk0/AopGJaush56oQa8ET
Fj3Y1DcUxlvDXngS4lhO37XsgTOvXDS1CH+rRLq7MdNmbdUxb/pcgWBLrdcy5/hniDyhX2dkrEFu
/iKRTp7VsSk7bi5Kbp6U7l1LbIU5TWctGtwtBssK4wRHhc01CkQ4jcauKbX3P4OyfDnw/4rRcgFc
a9Lqsnd2rhn+fTip9j3NzMzqOeQy+5aRfaaWjioWnkEPxpo3mXJ+zsGHGukSHAygLWzj9HNqqh+q
HnqCDgRToFKCYM+qBcHJ9YjfbmdLnYjhDHgsNCQ7NF5L+W3ccbtogIJSnP2gj4dNx5oQ3avB/aWk
hhjcfbgUKwQS0pQL/g5lgFFHWCPcGIvhsvZbLoqv14sScL7UVmVj2BFoSwadEASYYo6q1TnH0q94
bn9PmCHA375SFHoh4FrJdB9Ki4K7Lc/oNeoUNj25l8FkEwKy1hrEmmNkcj7tLO7BjWfVPYTYXT0V
p3z8bQjkZtI682/FYOj2IRzQflaOs1/GbzZEyd4yxI5eemySaHAbjuDHEK2NH3iDbpS6ALQwJAvq
kDgmRlkFeUhwv9eZVOmY+pbmiVWY/jipLA7Yov0VovM2miYNUj8Ahhuqm4j4Pa05hAqnJD6jG3Pz
VSYXhLRk43NEj6Czwm4T6v+EV/JeXUiFw+vw9G+fuqhDEx90J35DLSiaRHxaEXIypNvn8RHQfjbX
yyp/MWR1QdQRiyYhCREGAAL1oIu2mAYlKMDuue/9s135ejbyMZPFjSX/ReFUdaiqBgzllkSYSWRF
R4+GB9kMV/4AEwRIpq9hAp40qM0BwBTpbmB4B4HtzfQY9bUb90Rqdon0r7jlDQg27yEHcgM6Iece
6UY11BXIFwE7NsmRs7k9AuEsmnDJ9JNGqib6ctzdFbs3T/7kW+9dWhqsX1qNzuVaIpiI9wIR2sFS
sbIbEC3DmvSfp8pC4cUNSxs2+xOfYOpJOvbJuhsWj8orB6ei0CFXF4V8zcYKKUNdlR8Sqk7zbTFB
hA1Fv1N3UZZfcTRC7b1oj/8VSPQRP4H9fbLxE/31N9PLrn2Vj1e2NqVcQ4gklgTtkiSuC+4c1l2G
XNmfR97Bt1nA2fb03lkcbR/P703Z6BTjxGcCXIlQeoE0KCzMe5g/fW9LTWjLZ41qFy3PyEdX4yhM
95ClmdX/jP4snQb5bNVmTEJjFdXDtR3zZHJ3kRQUG3yTvirPE8UnCSxTmYNKQNlVxF57faxuoNU6
evYLzzA2YquUVwKEe2uAy9prFSqbtth4O7qeMbIC3hYcE2gfz18dEucVl3OT99loGYFM0A42KXM9
tx5RfI/dE3WnWhvWgRIuMi7tV22FZTimJpUXv7zGsXR8b1eAgbu3azhM5vUPICkhGUMLyH77NfR9
tDK3bHbXhjKjtGGAFTrN35ZuuXGXFbnN8ToIWCXzJa4ywncK2EAuwGQ0cQ91CXVPOs2MkWoljN/C
A+PzN20LAsSQl9T5KtVVK5My5C74btrwDCbW96vO9YUGUnRdT8VGlibWHQaIF7fQTn+lNzEYdPZq
l/mhgGANR9bt8AQlYXqXoRiDDh+yrwnb3/JE1Mrh45P2ONv3EGCaDqUHvmS68VT40ffYzVtVkWGR
sVDfLTjZgU443J+YAG1sfylljclUgNeDd6EbCrDoJ7c/Q793xxxEWvt5K3Aq6S0PQkHeBgXQLQbu
7ep3V8CVXiGXa0wuchS50AtnZNNyVFAjxstpy84zhFraVcKighAyVr5xi5nMRmWGmFX0SRuS1BjT
B1mk3PjEgyojTwst1M7KFUJoDDqznRb0C+VRskqVDQ4INjXReAImxDYSmeogVBmiu2sFnDtLPDgo
2QhLR1dF6ytl2yiy/F74HdTrhum584IZcX0S9fGY9pC0WLdW/pvxTXaqWRQE5v8B3sBT/eX+2swy
IjbsqEDqN0ZwGCycW1qD76rlfA2jXyau63/7FoaUnq2uXNBMrmF2V6yAOBYrRCEeu1Bt7631o/qp
cLOcykwv0p+H+AgRHaL3O+YpgEg7TeJkWF4ZSOW5R0hCQFcVj4MdYsy+kwhbE9MyVyRXEglxFcgD
NZty7UY2q88g7HCsm7IDQ2wI1nieVmEuHI3FVcdLmpqejPLshFyABZpu3Eokdck/XtjB8OIgBEh0
sqq5eAh6Qg0JIGiCleRyOhDIFKcqa9w19U+EkzBik1tm3Pcws0VF2t7obMgga+m1+rhn6A1eyzZ7
5ciIF+OSEdmAFdhqKQkvRaBg/2EHUjVSLAPwwqCwBdoWvn0mL1E0lUyMQvhmT5kwlOb+LGKsZqMf
q4KJSEEjzsrpj1S6MNFxcrc7dfVmfRQo/+HRueDddkqYdEX7EPq8WCrHyxJAYuLTOGaSYLgL3tzy
Mwi9EX8wQk9phP+puD6EPETgF4HrPEQqPsZ0Y/eL36VyepVXizElc3Depc4IA5vKt4yPkqH/Tv94
+JN4lzqTGjLsKxuZi9lhiLmJuxrjzlfaAO5rH/QMfe5m5gxG5beQ8K+30t5YoNHKIALW/DU9gpe0
wdcMc5UJf9z3paMhzduAg0dDDCROraBaQODllbHMvPWh+Aq4q6kQrgpe7+InS866w3FwRznWmign
xzuqqwiHiiSXDUYzK1ULnWLvgt/NivF0srszsYv7eWdVXxTdLEugyQ+6QGUlNRPQkp1EqA7u8Xpx
Av1TVZqSQsC6r2SAd0A0seZX0JCoeWswCC60wdf/NKz08VW6qn9UreX38XR2K6t8zzQYALp97t36
MbmrR2NLp87OvOXF8TVJQUohQjwzQPWkrbH/O5/Qf4tri3uVO4RYp0QN1y28sfCL9MyuBpbsnvG6
VBplXVBDW0AifejWCYau2Nznre3sfy4WyHfb8TgKcFEIEmxT5EiJjK44nkeUkhMmseuoGbv0oytE
+LNhEdtTvLbEYn1A9Yfknl7IOddi0Hj9kej+/dc+WYiK0MGr7Zem2uCIgeH4UQ8nTPtJRbpVNWFy
ZxwH8TKJXLpG2FfYgStWzW5GL9m8Uyt1ziSgJVIv+4krZ7g6rEfWIDoksi9BTarsg4ZCWC8+wwsY
LJsPtJ2NreRn8Abtg11cgEk8DOhPpBUbvWDH3FH2a5o8fIr/umB1PcIsX9CN3DqyAmkxGmwvYLEd
k/9F1Op/kAy5badIVTuUdSQiE6gSUm/HqvN6Qenjo2hpU0xXmv0nFpof5iOKwWzLLXKjCiYMNXVR
Sb2bsn3XgWtS3jpCwCejrGY+KReDUPI/L7adlKkPJfDRI/tam452AersVUMpW1aj7HdlNI0DOihd
k+SFK58GTiIDBOP1HNs4WlIZLGgOj65h1JkgIm6vUvqJHdwwov9+omXJKt5NNtYhzdeM6e5U3Ntp
LBn6hFjzjXrAlFCM+WS/LQWXOD5WsO1mokxnM/Tiz69zvMR08tNcl1uSQnFvBPWmhUqNAk51UQ2w
GhlHP83kLwRzZiW9P/Q3FZln+JaYnjT8WF+dl1X4UhaOMcpxKjNzaXAxggIYGDVD//JvtmiPzsn3
5qNl0rpI1y8r5I2HvI3vNJKLKBYEboZb7R54PS9QBozw13A+ceELNKrpyKv3tPjx3W5HaeqvCFfx
Y0eVk4PciigRim9SnKOcCwcBjtOBPsKnNqW+9RQ5YEpG+mcDoVieadIYXiNeoc4yJZ/VljwdV1JJ
v3l3E7F8Wtn1DJu9phonSBA3Lc3PYK8t9XanYAshlPPbcfMyzWCfGEecJxI9q4tlNq27hQEEKID+
f8escDHHTf6qbc3DhnfXCCLt4BkbVMMfW6xCRey4yuvg1zOgS9g78Isq1PMpsll9KVsxP16d8fel
SOTx1AwNDk/iOSdM41rm/zX6kYaQSPWRJ9L4AGWavvCu0mvMhzc+h1AsvnqRIn7tNiEZJiEMzVvY
Y6MKUmOwKp1XctcPjRptrzW8dY7v9iw0o9oYk5UIOpemsPn3i7VT97q1X0NyY5+Vr1GkqeFP4Ok/
BJSktqnCx+BO2GtRGo0ToBFoXdGP4Rz5KjRVozoqQ2T18hQJ6OPz22k+t2mWCzziJnucHLsjKJFG
3oj2YbiUHHkxx3TLy+ooIBGP5p1pDcD3cXxnBPTPoclPkoeFFc8oLxTwoJYcKcz3Rz4TkdwywIT6
Y8J8fLYGJauwFlIgO74zBlE7zqlPGhdA4NQJP8TjsJsVSLSo2vfQVVE3Q60VUkXETWTY4YMLOLXn
KS4EYiieF7CDWB3ND7lcg3/9xw0udITUTsqcIlvunox+dVrS62C19xEwlFgDj2f+d57GB8GzJ09z
XMXiigD9v6q740l7b+I91WBNdbhc5vPOKZWRcd07v7Or3qnJ7pJoyMTFgf6p0yYhMn5wdxpFd497
G9+SvT8nckFvWwOplmWG9XQnTCGlR8HGsMAg+N7TxQJDtoL0U2erOMCgQTOgnTZ8IUsxRZL6ssaV
f2ljdIrqkP0uHQqKin0M2odGzZiZKtfYnoohpno4qgZp3qypZezllGf04ODZOhWG0G5dv592zaAB
+hUFUvD8am3R6raOYCNNBw0P1Z3poNy5HzgTAnGismbJ9vvV4LPOfYVu4SK7R0KPuXB1ISSZM48b
tDSTy9veznxqjSFITw/vS4Qsx01I2tZCxK81PD5NAYHQFkylQRhsrNtmC5jx48Zjt99bDK9GuMRh
EZUNJfi07CZLkiy8mePgAIsJZucFqDGT+dSi0vYPleZ++B/PIXbGQ6ByrVzM9t6mlavCn5XjYBjw
qleeo7ePryyrEVO+P1TBWTK9w+FxUpedbi9zFtxCHN7jiu5RIaO53m/FFyL/HqAcVHMIRfLrVaog
1LYsMGeNHRAV3OlYQZ/agNZ7xvEJrcRq3rHKhxHKWWj0l8Idp9t788eDX2twue2fFgTjZ1ApdCSJ
NQp4Ft8z9V7WS+tMp/Yz4db/W0j4rzx6uxrJpnIVpis2PUqUKrxppl11M/nXlglQFAJQip9gQSD/
BERGusUYO+hsAQZFpaD9F+iXUCcGK2zHXwp3p8JnrM9NXUwtEKWUCANEWQuYyFdIj1ENhjaMuPoK
WrE7EIhhuS/WW+VjSJJeWjwnl4Es7Tx24A1VrtpAEKTLbcvqZipc6wrLM2XWM1/dDu2JFn41EGoU
ft1GXRycBPHD7L2d3ba1KX/X4YctQQSn+/srQWpwjpUdfjSulGrYPgojNUWJjgvxphKidDWS+d5y
cnW8hutwjhJNkvU7VlQl6v5RShTnix7aMPLw3vFRtsvMeAkJKjU8oeA/M3ltYf0wNSPkjeIDHAkJ
CRjvoIDjgobHLnIqvd20PxXWNo5stwXvfNh4FoyF/OroHcGf/f+ulnobTl7amtTUyp5KvTzW8m7O
VxOhOQi7zshbobMLA5ldbWoJhkSWArp67ul5hcejR8Y71YUslposrQtRHote+c6AV6HhS73NreeX
6Yca6mpO1b4rIdcl8V4pkDOnwMy++X7C9HL5eNsDzq9DZ8yxcTXSxBw0MF1LIaUBgJZ+lZCsbL6T
jXmrYt1CGeXQ1dXlVwAiHFIlEwCndJIU1L0D8kjwV1n8DYP5aI4J/TVcIzxZNNlvso/ksj7wdPSA
DrzTB7nNo1oNLy/8oQPToxfhn1sBnI25+qwLAMp6D/yN6OdX+5SrS7Mx8FaPjfYpviecWylFQOUd
ackLQn+Y947G8E9GQFLBfnP4hZL2zZlnjdX9Aku6nsSzMZezmL7INeg4oI3Zr79ntTDftw12c6sx
y8CHjZKMVnS6FQbH8R8LBYd0itUCJAc8GMk2w6AIZcmsYxllUVt1YWGQ7xd83lYVR3wHHmKYyvVo
vFIzzrC9cIvxPCB7uVr/g5kX9IPmp+C3hdAtzXNveymwNroxoy2IMZq6l+nRXZOhkHvwm+oDuj0/
jHYpyngGiDMxibmM5HCHyq0feNPsKQyruDPiovBjZ/QWq+z5rioSJReIYGYjkq44X1pHIuVQqANQ
+HIQFgJFwnPvmIJA3Y8HewAsPPq4jsTKK+J2Q3PhCLmWwbDPWKouNblFcsucGHWC3+sOSWUj3CeV
Xde+PDc1iM1xGDDDv3VHRyk/6hZj1h3M6+EU9lhLCJtfMk2sCQtubDi4/COjKbjGlHiFXr0BgDBl
9NBPppZdIlhyOvcvJbBSLulyHxZgUTsEX7tCZfL7LXOslVH1taHTcYc9R7h9ilIE7le1MuLrgBZ2
kqKZsfYeQvCHcoraT3qZXyH4+0uRdkK76wGDJ4yrS5dsobVHqN34Vj9FjDitEdp+kpSEpYHfrYgh
H8phvRUpLqCDsQ/yIXK+pNQiW10RvaKGtsOwgKOrdWiCMwvQIQbHYCHs9pjeFsfheabH/DXTZ0d1
HhNREmbEAinLx4DlAG6m8XEWOPy7xD7+/dh18lCDnnFKNKBqcIdN/rEGGW15Q87XixcbLqOvBYKk
DxLaCK317ngB5Fnyqbc8BcQqD/DH5CN1ZipgivAC3SU+CJT9Y4ODeFnLdmYQc0GqwNQKt76ITSJh
IuhK/2Jbot1AoXv/O4y3ErALBkSEtnsXijUsGJBuZBs8UMyPWs7uRg/rL/UuhpQGDjQlAlGHnH59
c58Aa0GK0bPCAeOGc9I5Q/4EI9eGKNTcaodT8gBP3fottBsyzp24S/6qPrrR6MGZCqvsJB/nfFIM
qHFmA2Dbtg3z7cIwR1e7HOH3O83pXwctYUTLESwZJFfsTdheepQ1ABYrnEJjSdeYUf627SkstJeC
ktOcLznPfVWQFdt1FcTHmQkfCH1hRxJC7/0gtp/w10D6//vzo9F2tgTzCNurNoqBr6yNRWJdeeiO
a+7FAyU7ZrKJUqsDJlMAaV/WhZE5FC5wYu/s2qwFImwQwi+VqG+UiafgUS3fhQ2mmsP+f9m+JK/1
OyXCbc/MVpumpS0fi5KfTxNq3FFV2lSf+cPFJRDprV9oYhtQSkKfENhu2hS92yC7DGg9n0EVtCAI
ANxla7x/rShnX/CYYsd+drZMzxoVFvS7aP1ba4pbQUeuVsi9geikgn+Z/ffUk/Ed5+TO+aWU22wg
AZfw2C5iO/wcntnkdPr8WEtDZLSNsEW5+vsNEi60QwLbttbCSXE8M7vWEg88HVw7QrUT7TNs7uru
UFZh/ZXLHP0HYCbFwh4dHin3eKyHTobACDDCbaRTh3EAM1rlPf59ZxiJy+Gscu49M4/CM+uJ/lXp
FFTC1gxm1RxX6OSaBBkJ9bmsvJxYjlK4I1w3ytOdjzlPJXf6vMAMi9Maz+nNagWOW6RNBUHM9moI
U7fZtG1KhvnHV1Zdj6rN1gQmFCe4WRGXK7GeFAIsbIdJB/3tHYaqUnqfFqtbTPdR0U6K96KvlD0/
gCa35rBSC+GWuIStHRcvv8upJJBzw01x2CHgUA7cJ37CYtD//nN83Yva56MLSbZ3YDvrWAW06Mfx
UDkoMJNp/2QcqukD+z8KEchYC0mS+iwY6jzHU4aBMs+SJSVf+YuttONuQXPKCNxM6e9kLrnD0uqO
MUk3qmzwsZCUjrIfeYUn28ed2daTQ20N3Zg6MH9qPM4sh7Vl05BlNk1cNRMLXT2LQeaNy58AHXpg
s+ogAswGbyrcwk9UIdk30recmlCRWX/iFOaWMkWm/Nj7zObYBzwlzvG6EwDL9vBAjwstTdgP8BFI
bKNjBpx46dhCSKKiDyXabUTsAuZXlN3m924CuMi1ILuoJ2UxUu9sJFieCD3qQDyPwk+KlpwFNk6P
Un67LMlvDQ7fhJOdo/snEpeYqQLsK6dfu4GFvNs4DBwq9/DgvDKHLa6iKoLWcVsipCLD+vBCfeTC
8lEfMIf1BK6rcCG8lR3+s1NP7EXtBritrJympCUDNKGxsgiLYVLcT/9HR3pYRmqti1HoUtAAAzyD
suhhzI5uS3rLPJV/1RnVFXgrvMB4xo29bGKnavJO7ftOLGGKefteEmPJ+mnd7ePTC/jdH+rjdPnk
Wt6uTfbqAaWstvw7NalenmrM7jkoIpzTaMzMF3P1n9wjrYeSCxJFm0ydoqtGCZqZ+qCoj/myq/G2
67WnptI1O2CMX7r0k7k61xEOWZ7yD34gzagl5jQfa52I2T0usfh1C1HSdZWKQU+lM7S2r2GoIdTM
ReFYYLkKGWjykVrY8pbYblpGt3sfiJyOcG2CX0GKeUNWX00YOWT4kv1YQvUP5G8nTPIs41VXnsyf
M0qqQAJQWvH8sGCGrQjxS1qAaOrlOhBktU9BEK4OSGs38NNJfmDrzbo/e0lrAsoPvzME7WCDqSaZ
J6a27y8k++e96oY875S0jWM+45Ci7FdBdpKHpeEj9KZ0jExuOEget/kTz1+lbcjoXNIh5gxXP6Dv
ZxcnyA6NTC/ExgZ8wsDu3I2+cuPae14NSt6h9cGLoju0iJUjaPsi3E8OdfHXK5mywJmIyfuGZa6z
2lkJHZOufZNs77hcZvXvYwQuzFcYvTJBAsUQ/f9Y8mpmwfmeaY2V0X3Cb1ZivdwEWWTrQWHu09Nf
VaFVR1jui+Rk2Tykd4KKcDTHaQSWxlO7iMZAnc0KXRdUiD7RG2Z6NW8RYx0bSP3ffj/HsAE4AjLK
QH5sfafEs588cvUXS25N6wE8Wcjgof4BpqtIFibADbBag3zcSC5HDrEZdaVy1vOrr1ZH61LrcnYC
iuWbqoNpxrFVeAtIhwMHLvjdmJLNMwyvkSeX2IVc5Rq0znpNuBRSz1N5Ejw9kA5irKGrQvWOVMgu
ohWtSqURsqruJRQ7CTHCQjDaPPctYBC5yaF94KDUKMjQU69VEZPgtotgjhem+i7l6Qo24eA78xae
Id2J/GQqbe+BRvYUlhbZR3MVtNSerV+5Ct5UiGmaj7ATMnmhiPzxgi8kWUBpUugLi/PxZFnTI5Dy
dTiWlASvOfziwRerNbd3wwviSEx8DGQqvby8SrciHM1fT791qzhLG0V8rwu+0L8KlVMnd132jX95
Hb7C/c2cSBFu5rTUDPATEKEWCjCRFbkkqM/P0q+4zm3uxqXzuQY5SYL2aUp8gSakrPkVQnlD6zRJ
Wfj0/ikClqzS0biu0UOVwyyN48uLKlA4rk7IIt9ADzZErItxW3GsLyFaAKSEk1MQbLjrHRl6FA+H
ur1GRmIfeHr29OOdd6+Zp/NrDRQSTiY9eCRzkBb8w4+bRTOgfk2C8Uu/WpM5luNF0775/uozfZk1
/JH5Qt6UtpxEogCqpZCv1gel+NxpOqgH46SLRjk96wAQMhd/6ok8jSP+7i3IO6ArNMCwyk5vYlDc
6OXGKK7kI5YBQmXPgY5yGdWRSI1yYjtNd2i+ixW3iMOMFIDQlla6MINUayQW81gPS7ikBlpbMERw
Fzq7X1DDyR8Lee2fX7ROhRQv2Q2iW6Xd8QzkSfbzsDtHs0S/rFnNLF8CJNTxxyVwBCxZ+QIQx/4G
6EY1MrMeOqUpVAw1aFPhNB6i7op3tbgIbSzRan9nbskl3HhGLZICpKaqt5bMpEzlMa97v3Yxdl8D
hjKIogzjKpVaWzChHHjm7iEH6I5e+0+JQ7WyhW7WOh286SViM36gQLpostQxGC665osLsZjJb9rH
uo88ytvMOegTsd2jNPUfCyMrtSBc76n4epFsdG3TD/Hq2HJyUunoP+EHnp67b7yXLL0ubP4Rbw+1
gIkSLqnEd3osEKDwzrxr4qccFDBxx8AikLuRx3IbR/6jbTC4pRYB0dL+9K5z3n5IbdTaVSQV/EdY
juRdeY7yy1qzUhGLDqt2t9KG+/CsBep8mk1Au1A3ry7L5UkSW+AVK2JhIbA0KTEgKbT27HIwP8Ca
irZcTCbyVbooGTLALLqH50YXQtpiv2TUstj4V0tj+JUWBEETRYNSRsBalZiTYZYcws7RDUSctPJY
eT+i5iw2ZFjr5lHQLH+glNz/behZIsimLSG9fVYuirxeepLdCpV6C3M2Ttq3Esn94k7aiABjQVbj
j9LEFWqvis95yhMYgeUqN3BamTdMD9wcZp6pXIZAbEZekW7B0mz5CxhBqvWZ7n7FamjpZ/j4z1T4
5my2B1p88NduTdsGjFdOrqtjE5pTKU9pUNCEExTSMoDyLMpcpt6JKoG0vdl2/xs9Hx19DCVfLWsw
evmVS2gMa1+Su+qSnVcN4Fbi2Ll0nbe+51bwmOjRiNEBRhy3hzVuso3Xx932sEuodHwjaQYhpy2x
/mlZ0eQP17ZblaktSaFxO39OdkdCMpmAhERsc2JNVLAxCPt700yducVYELO1IIE5wbvyiXGwRXFK
eRxbSsndKbIK3iXv8PL8bXVFg1xhjYaVnS3ba00JIPr1pnx9eAwzJ0hHzJKOb2caDFamgJjuo/Kz
/7y/I7OyE+i8EJHCeQPHb5dlUaGVfASgFzzIDbJ9xS/Xu89Q2y+NX47Be6HgsQvCAdK9CbECrpTW
rtfmTTwp8wIZYnkw+nXYJGxmpMAURqLx12mEetVUYQeZFCZ9CJRytqGTgnQ3PmvZ+GPjz+lQ3k04
cb6jcsv40ANdukB/kDtb5ljloKhBwd5XyBeYn6mD04ZEhjnNVo4ClAaWlEsjspnIE9KCP/1/pRgS
7Ve8Ggap7KRnUOrHP6uND03+ATVDYgH2qg42KcoM2zaZ3LuMO+XPzJFoa7blijQ4R9+kdmDr/pQv
SOGf+na4cQs+B6iPOaqa4xGE514BCZ9/N1SD0yAE6SZm5nghbNAZ90zxxAlsoUf5s6XSSs2NNGme
sYeSZOAZub3YAGxk//rz70uomQ6P2VX9sU7dHV3lCjWvWrVbsiE/cl4/Ee5EoGQv+p36qKiUYdsa
w6eYcBcNmr5T9bBTN2mGMHOaAjvXOh1X89jaEYKz/3056TYnv/O9sGYd+vejkOpbRUlDYNEBWquT
1dHCJYtHNJFfzwtWz7P/uZUYZ2iHDnrApG0hQIIk3XZNfEclvJuFmES5zB4DjkSSRFJvBUlKFe+I
GYgonsGpfMBGBi3abNmNFmE3W49dLUMYFJcPruBRTrxH5HfQ6um+0IDxPEMad5XE7otxaSoaehHN
NWlPR9Sw8433cE414FAa4kvtKmtH6A+PBWnALvadvM7zV6NlkcICQqAqa5f434MNl8s5BqVQWwVY
J2lodQa9C1e1pSMrHszW+ZpftuFt+40NmkM6JmJ1Slp/BLKzHlnFqbQx5ulgKtmv08NTRdD2oW+7
VXknBL4f2VKpb3y8hGBL9VaT4Menzi/yZTrQN44DSkvgrmviVLST21oOz+dHtGedjCjqDee7DWQC
axIHblHKZwHTJsavjQMkm6I7nqNfbUJ7Y7BeQS+Y0lWlNcl14HjVCJkXGqnHLe28/7N2RMyKTsjo
GEvmG1W4SYzt/kEaDuahG5ykajen47jBCOJQPLKBbAY+WH87QVsd6jcT03Tb19LGTEEv7Rewr2N9
dXxvW6sczAtBHgLbgdVZw02OCN2crgBx++sVb/PLLw/ljzALzfPMmR/YsYWncvos3KSoEhtwDk9t
5fxX/cTkNq/yYjvf6WrmNryyTWaD33MlLTMAE8czBv4gMWlR2aLgzsDHi9Tc8NGXJKaxXlWhd1bx
Sv4uct79wKJNWXUavDhh5ocaUAfxBwGSiTdtx8r6OSQWJY+Ae+1cYqFZktH2POoPNSQs+AFbFjXz
nmPbrOZNnZDdbrDk6vQjlIgOOJ5lE37muk0BPEDsIpn7TfMThK2WfvDCTb8hKpK2ad6s/nZ/c2eX
VjEAI8XlBPyLe+l/z73gEOgvsJpxGeK1w8Ga+n8+CHJzy/8Mefjj1LXiYPb/NNVmh1D+LLkahJid
fFEdrv0lfNFfO96MHa7nWyGIIiSdHoK/Qkv4hhBDrrQSnwDJWtFHg4DMSo1QXngZrcC+M/Tu/nlo
bSzYeqSpK+JpiMVAWZCvnd8Hqi++o4Vyb2y5TOvoyzbmk84IB3YodRc8mZkn+BLsnFU7WbLW8OEo
096QUUg8KF9Ut56ATWglj51zatcn5ux7C+2zx4oJ3G6gt/Wg9gl9+tp7R9ev2sUu72U/ehta17+9
VJnKBLH9KeZ+N9B5nC3AECti3VcLASrIZR6fVDQuGVKGUqk2IyjCeSIQ+wL8pytw38D9DAbU+4i1
E+2DaRCOfxxLVcRTYYnjO6iL4pZbaB+fN9wJmxbMPUYuayp27RkGQbhNUNZGiicLt08zHQX1W0+E
aWpDQCoPB1OSnLeSTEmHgawoTankiy19R5mw8UTaJDCtzcq3+8GVxS07Neagq3lyMCpWsq3VUa+5
pTEzebCSllcpXv/2n2aODGt751O3G0RrF8kY4PhRZAY2fw2Bcz7zCncGv2yJw5iIrAEfCh3YyEwt
e/UH/NxZcU3FqpU5v55crida/hm8zk+BD8uPdjS5xBSRiygxkWH6K+D/3ZkBhy2SGU8g+qoShYzz
+4hA7MHoJCLWXuuyIG3nOsCuYBrjvOFTIXwRT+5o/wRcp22p1HO8SnLnUoFQpZQhn0x9wRym+a3J
vftA55FuT5EY+egEOha/JhOqZvBpVrYkPHqiQ5QyNRdTQxX4MW6LHYAGbuE18pLllI7Kfa1BL8Q1
BT+fb0V1SAmE8eLMV/1Chx97L5k/sxJN4aVBSQ2RNv4CgRL+U6rC/qT7FPiWc7updqDQ1OSyzxsM
lHwM9BqoxTtFXyOz+KuxDYoTz/oWIVtWOsUSHx/QekODZIcT81wIiv4ObYdJVDNRRFjqaT0vZ21O
FyC4z2Unt1Bl7tUDDbIgF5PNwMKlnOTEYerJrqdi+efWxzKJ69ex5v5Xnl6wPlNFGWNH6psc/Kbb
6U010BSpZrHL4ExYYbYDXOOTt3QLSbBnrW5LNJXDJi8KW9nQU28srYSOaxfC8Yf6zbzfQNtNjeNP
WG3P1nT03Tj7wHUnrFHNnHijnQntylu9NQZTDkZ2pbLpHIw3IamEkAUSO6/C/JVT3qlmN2uZinDP
HesL3MmwDXHQG65h6sfAt70a6EMMlMFjzki/+QRVWN2khfgLzyzWzTyl0uWLYjvtkCq2aCrCoDsM
nabT5RL15+apgZNGUINV8+RqxyU5r5q2iXPCdiOgdmzK3oBLcZ/IEG8kDDkNH5N/M6AbwJyMXvaa
psQUjrMoXPOu14/9saZ7StU5UOvG8h7OVqVibtGbnQa/U3OOE1NO++ZxaGEsNgdLWu062M2579B8
TenIolaT/ikbalPp+S0ftoiJlqRsRrKaK2D1sLAqjnJB/vowdO7LqeanTb9Pw11N4OfLNR3sNcC1
gA+BMNVaDwb68LbIdNaPSkB/TeaZyKrXRt0b/iUa63Sfu0/lPBvICqQlCdIL65h3vdEBO1mnzi6Y
s3mHer2N4Rm3UOVb9MM/AiD9b6T/fRH2Kf/gtZo9BTp+4wDmA+G0SJMxLlWVumEnD749vqyilvWF
26qzQ53ZzihxpxU9LbT2y9Zdl7YnGx7SH1n509COZMwOwd7j4hRnN2qFa2E1zDBUJIdWEThQhM/s
DvTvu/xf97ONOWFfQ6Wnb1MZhqDku2jIzr6Ur7d1snm2gww+XXDY7kd64X1mrUEpLnTI72rnG2xA
bGRtj1t5BQJYw1iNHmw5QXRLlYiKIQd7NjQ5jV6KtZJMHewIPNK0mTV6tyHh7riswBt2OejPJhK9
C60tryIRgGb22koKsBpK6s94cNmbrc/ysP/HS0X0f9asFjJY2DS0xjGzfzsSL3JkR+F0CnQZt1RU
Be8sa3fr4FrCXBkTXdz+e0LV4FbxQmbDpyr34H7mdPSNo2lwfgSUJiSOgiRcbV+YtWOn++XhyL8A
b/eur4PduANHEZaoIhQqkBSgnr1KB7lLdeDrvBLeJVCPSNW32JMycvr3x+sq8SXwc8xxSn7iMo8I
GIuqz5foRpApwoS3CTQSoHJQtlsl1nZubWRw0YLwHPgPb7isV1595I/W05OVKeUuAYTQI3O9bK6j
YrrWdjtYoxb0L4cyn0gNxjI8dV8+xyUlUSCG4NAh3LKlj6vZdZQEqURK8DttMvrXVgos/ijv+BJD
dj5EH6EPacX1u4A3C7g7Af0taTJklfv3eYbPMPolkVXPlTLmsvNXtqGlu79hCtpJoK7KEYFMxdx/
SKe2XhRLam13fsZvsYOf/LvMdHoSapvY5nxlLwXmwxnc4pUhND0d1m2aNXw1Ks/NO0DqScZtAjaE
bZzhCkWbClYz4mJx9NzfZDFRd8ifb+5EV+r3n4mq7wsYlxG7U+nWkX4gzN13nCJqpZf/2vx/xe47
7dsuhpNcFk1LqUO//nazTWeDy95lgmrVUIrob7d3Rg/i2MYegb/rfhHV0IWHLYu32VfVT12zjFqp
7mpnn3HopdxmB/YMoNJSVUXFHVyYpRIMMm2UDVq4ImcnhtbUjhEABUszztFAfqZrp/4zqtIGqgvK
8zmeyG7KVwuTkR8GcAffXvFSd82QzbaPynIoO7IVMb4PwcAtZzsmIN0t8Jf+gPIKtH5+QRtZpnNm
2ISxc7yXtHdc/C+Ujfn0ut3qxaHnoi787q1TGjtveJ7jWGH7V5b4+ZXKY72D6vOP5oJufCLUSWvE
Wrm2uscPYn5ou0/kBq0wQ9oMQJ9BuEdb3nt8oEle01zq9e9EG4/SIaL4O9M99PQrnXwJiTTUNQ32
6iah7BzY8jTb1XBU8ThDU0SYE0Uyz8xnuROcEovhFW8zHfatHeNBoVtn7CwwT3FT5INi1DIqGLPL
EAfEKz9zbTYdHaIizQPD1GZf68wWRdh1C8pMTPn/dHi9fQEeq/012rQV1ndbMGNPDRTjE4y8JFZ/
3Eay3YyDfOYrlazNI7QELCJDnnCPtHAGvDH2+TOMv64GjJ/cZPizTUwqzqd+DXZoXUOh1fczrs1X
xa6SNR6YTh8OuCYtJ9KlLg6qzH8y0g6hfKwpXw65MtdFQ8VmaSNvfJ1csl4qopXhqf7wn1HQ2Teo
W8gAOxnIfb3l3KRLzHx/Z9DbDZXyiGV2ecV5LO4oZkd/olU46GgiFf8fMIrOPjWvR9fesXCL/m6n
6g8FB/NICI31As8pX2lRpI6GUNEc+P5y/gpwQyH7V2QyAA07EJjs/ddPm6SbBIAOmLyKhspKKgiH
d6k671q4bzFFWUrn6k5CSb6+ytgyDbYHlrkN6rI6GLZaVH5zMjk6GcBKw7jrbN6yQPJ1XXQPh3Sm
A9xP6YwqD9oeLbmtHWqjmAm32a7fINiUgZ2TAg4t6A5E+/X1sGBBPRZnAgqnfEJbOH0YQp5dq1GH
mc37aJiq/015rLmRZBTA7soDdFxAUuq98dsa+n60wr6mdwq1ahZGAJ53A58irow7gX2ozDrw2N+S
eFPMP7bWiWEiXA8AA+9s0CRG5C1EEJTvTxihFMNhBm7HB3pYmU3mXCs5+58aOXkS2VhDQH16xckj
o7jFGAr9nAhsYfM6k4MKnhw9ldtVsIPCxI13AfWtWtS0dD60PiFYeGc51wcB7HJLgWsu/6xTVMzL
ux77KxbR78kW8tk2G6Mt+IyeVDs1AI5Gah8ZDOFs3AUWQX05hISH/TEK1Q1LKlvpBPVsHMdkBw7Y
sMwwffr2tsPAxxmUUkUwR6qmKX9DL11AcXWn3zgs074YEYf3EeJfqbMEhWStXdkmyrmzliHSg2A4
8wi1s0RVgh6M6OVm4Rr3/sAMrcDl5e6vrrk4Q9H6wVFgJFEII3Sdf9xeMZYqUhv1dYIc1z6Dgged
t2Khw2bovHL9Q4BYBiEGTPS9+eujJPiCp8RLN3tUPucGVerclJQwG56bA75VP60ivZ7J8CvaPOdm
zgixxoFfcGyjIteMsWmiBVwOzNQ58WTsjXv5n8Ghzm3pNWs3489I9B7hbQ7P+4QLdYX/tqM7/BoY
G4oaCDqiUPTtUSB0ZENuOFM1U/8gfx48K7Fd8sMWYGap5h7EGSVCm3+6cVjQRJPp1FVcabsTjGPY
ErSBPeZ/JuFJIUHt2xLwhn8j3ZApFSVIE4hY5UU2iYfRqsKYq/s8Iqbh1juD6xzJrazQrZsTHfAK
p1NsDRCed89JkDnIOGAQcjJPqnHi+Z1nBzu7tvlrxpGoG0K/GL8zpUDhcfeqTYM6nKjTDWb8Eufs
qiBIjiXEdohs4diiInPIyr/071oQRYtqEU1EwEaGeg3qENlfuoAvRkzRq/PerlgrKVxWQHhPXTTT
OaX6cOKZHxKirR8SXHZKlz/6QCXasim9I6dSOVY+PUoGTcha2zYp9Mtgr0E0XVV4fYnHydpODJOp
cdWB2Ksa6SmKXIOQAdJSD3NeMg1ZtV2z2PxY6wl/BwQEdR0q8XVOTtTnSp0o78+lQ2bGTsbfvBqn
sE370FzBd5FBV+Rxx+djuzwuQ8FKCmHoqJhWgr/qvSvC8vBYJ2IhoLSKwFnuFCd+ci12iEKzh9/E
YcWErELw6sOGAGDPEbRoCmF0VVPRMch2WnH6IpqHSSXdaDX6uCshyhDin8RSPp9F+s0jhwTKRpFs
xzv/883hnoSUKf0008XRNex25+GyBOaYDtaJVL1uwY1B6KBD6VvTh0IzyaggwmlXX1Sh2sRkgysb
PDt0X51H4IAcGupUanIWL78PYDSKi1MswaGswU2f/XNC+7FlcL9VjiHIWIMdmSKcD5yUEAktTNwT
X8QpVgLiIpYbwmSQPsgTmGkvges0Z9B6w4EnyiRa4VuY9TVNumVB/mAP0+euWCR91uMCZNpnJ2Sr
0fFVSk/mSQZcYjavVLsbYZFXFY6zoOrI8XAPnXuF5GH6Q7dOq7uDVAIR+cknYD//xIM7AvgpF0L5
Zd8O1CJP+0COmdxoLjpg8laXNy1rQj3Q0+KbeDoATCZvmIAQRu1+xDR4WV/QtZg0XyS3ZWdAFw+Q
v525fKqiZtNYuztqVbP5EdpnfVs2GkQ24atM0ZrkEyxsDPRm5djhUxKoTFfsrx+y4lGQzpb9NQCx
XfUxsaQa4xkbMo4DxeNdwvBWa0hH3kDlWNS1Akme2SoWfXBiDeb13TLeMrPcNgbjHFm4zo5omCm/
Uikj42iZa+G7pKNOZNbB37e9IC/3iruPxHYqA0IoIEdmyFL2OXHNDiXW09/Xmkfd1TAkqsj9ihE0
ODX34c4Eam8IBgqaG4k4/70BDstYLQdb9P5Zl6cp7pYVp5G9S9evln8H3MB7vt+ge7qrDlO0BC0+
SJ+TOuDEBerKaoQFe9QRxMVXqzDGFfR1PnV+aUJVpsYm+8CAzOMP+uTLoFuZNBjYGYD3w3iaRO1Q
rEYtC5HK9LipkfSwGjKFT8zlHHsLjHPWxbaxav+8Wq7l9RTsGT1JOWfbBNsAlrRSSGOg+oEKFOlR
zVwitB4jfNr9pBHhrKp9bZ3zAh4/cd/Cd6lAhwZxF6gqvHmd+7duLohVdOGk/u/auR+7FGo3/QaB
NSblb/UwstocWz6fmjWjeMRN+poNh8so987eKhh+aUCYC61/FiVePkdCUhxolIrsgTJ5LUTt+omz
D+D/u6BqKVNW7K1V+yOoLibl3weoczAe3X3HT4ZmF320YMpQmCDDSaxWlhywb+O+I6XHxXcuDLZk
jJwOfvc48IaqKWWNliDNaQV84rPQm6n8VKGJC57nOduD53aSBCe41oTtGjneLVmuHLJfysJyqd42
wJkrso0aMidoKzi6GGb7T0/cpo+iKW1nwT4tCpVBdhXoaCYmBa7q/8cgPrgDki9YpSWx/s7sqLBp
5b+IkOOWyDGKnGf7ma8D+lQtxRMB8cGC7OZtnUZt4uhTiF+A9W1taa0+Vxdcqdd8KXOOg/e2n8IU
Lea4KyslqMZEDTsgrRoLdV6WYys0M3oE+8SQfCZVHzN1uj+mxs2wGbKTduIQFvhdu084/I3oKLcg
cnk4Aq+9NXQnLexIB3iWOJb305dAeXFmJOVkysxyNLi8K1fr/0gtCZeGlF3Lxor5ZT+Z2R9o/QK8
pB7Q+g6X3ArbPiCf+UpwdDaCz866p1m3pCpzmDv3cFMUbgFQ1W8vreauM2mtCLegweCBY3xfp98Z
FkLcLsnpZGx7QV8qdFxJ1qtca7ubaDRq7M0g74aKlDbc8idaMo46EARbqxmzXrEwwtJpR1rDgF3Y
SRLF6V9T8gveWI9w4OQnqMlUXN5NB6CidrU4HmNtSY21hnZkD7KyQ0qPnxpZ0AoSa4tBsr7i/ukl
4b8LTT6hnR/zZsomcT8KmgS+OKfywlJ5YWJDsPzdmN5kcOfRu+jiSV8rOgF94Tu5FKth5U2jAvib
b/6/cPEDIUZ/SqvpDfeVWFcf+3u8smCILMTsCCv+MNBRmPjmMswD1151L+Iizoj1jSTnvTbwjMTX
uZKCd0YAyHp+rGIqpzfYAS2D74ze+nqa0xHKwrPEb+cAM8Rf5kM7RFgTGRylFaR9+U4SPVSeNTDM
Ulr5pOai1xJ3SB++enmZ2KRQhO2RjBINrHL5Ujj/5P+KRV0SPm3ySaLn8XD95dyr1b3KAcuLXyB7
+WYayN/Iax5HqPWT3+f36+tEJ7iqg5awcdEVWgAhl5nedbj6qnJX6nFrtKNjkpzcD5F8PVzh50DO
EgqdpxDYRfynXAJ/zTc//N+bsUI3Po41Ymdh/zgLRsQHvpKbtkkjoICWIH2bK9zq55YB2z2TA+S5
4jx67U0NmIJh9kaK1iEgQOXqlfwkgIfTPnQwiRm05+68+o0AB2EcKIZfgznQj9Ou97svZdMR8qgO
BJIjqtPmAaIGwL/tawpWPCTDUp7uNpLoAl9WcPOpveinnUHmzk0l10/EkRcyqnowbDRgsW7H1m9u
jdiMvI9nB/rZCsItzUTeLhGlhZ7GF9O8Rx0tuLRcMqJK2ZO1xgP41coozDVeqxP6A40vjkAxYB/V
Zj6vQxeSKBP08p8vphJzAzUYeoehDkiYTzaGDh4/mXVlpKLK4y8J1wDlhjHxsMBLDC3N66vrW0Bx
XuUWhdQDMpXlNaUXTdg8xLLeid1scr0QIGTsQo3w7wXaWtuAo9JK5KD8PkkGuP3WyV0m3ZPSwoYN
JjuG7Z7TPpV+EIfQBhrNGuDeAs5ewBLICXK0mPvfA+flTlWijMFPk6wfAsNumXg75YOj40H2fmup
Ud5b45nYRfl+rNW7dFHPH21J2TJ4cNvX6Gzh6gBljl9Xzl1/zkA5iC4bvm0baFnRaLduDp1nhAqt
DZvgUYuYt5/JQwkPH6IaIxIk4CPX/Bk9/PJ0aHvn8pejhaW+b+jjgWhS+fOVurzNzoUytNysbOYP
2Cky9tu9NyROR1XMyvVP73c7VMO/3UJ6AbYzknQB1wUK+KEi2DnRI2CQDnm9FJsiwCV4kuOBrqJu
HhyLoWHb2dZ7Uzaq7UkKGMnoBpICp8M7F76Z4Aekk1sKMp+tYVh0O0rb5OR3olwR5vz/M9KD96gy
zoChOpCIX3W/ilgusPPQhBVYAHebtGj55Yl38kJySl7GzDuf6oWs6kkB8ML20BbsTGtcgP3+uylT
8F4KewfDe2nWHPJIJxAJnK5nxjTludQTn6KudJPq5eGA+npyreKAz4Xw0WmIusXtVhW3ocF2tgB+
Omd4KyTeIR6uTG0TKz5D3sRbKKD0Gu8PYR2zUul786as9v+9qFPzdoC4sPG/lpOmTz9FI0SBgPcX
ioTwwAGiluyxeR0ucKPxEqlB2F89n4GRD7i37JcR2hSynyT2D+NYk2elXlrS+hGuPYX7hNpjQzrK
IPYmhnlq9Vk4xtwTKMjibzIfJTR00OmUqzgeMQhneLxAru+pbpRmXbl3QxEQioFbcsii1APOW/MW
sileqfCUWo6L/t2/mDcZOmW1MiPe/XohtqDRWC+Wug3C71ELX1QadGEzdCCW0G+nQVh2GwT0dqkY
TwVkb2pThYzz7O28Q7kmHXHTI1KYA8LdIEnhOSE0C/GjHANJJ/MnnPpkw5c3hYV3KIY4C38UExrD
Hsyw+5B8fiNfqv935rHBhF4jha2UaTBuQmJnh+b50rZe3kpZ3FXh7Ao79IIZD24+94zcmM7UW/xE
R2rba94ZIp+YW0HKukUu/BFqOAuX/VsASW34hmlaTs4PbG6xaQxgBxVXIdyJanGUPFq9YzabcZ5z
rpAnie3rkAS2SsexBJILMWfXiKOcJ7xUHBPtWYGpQCcgDM8E2ic4g0Wu3+gKY58TGGexNn8BkkbB
T3tlEGQI9v9Rl4JI5xsIi4OPezw+T9lVwQb7ZeqYv2gLaRMj9I/7uRKuDtJ4IReYL2VSCaNwWis3
RKbrSwHgopqWwKBBquZQSoWnxxAxfUqwNSn5JKeD4GVav2Ypqs1B9cXDIl19O8pYjwUQ9jgGQLFG
82RDO3lic3gIDvm3I0GV37+DFv8+zxFPgo63HtwlsliA3rUg3TyEPNTNbhFGusHr3IOOyUSIusGd
WIDAntCgc4/mjb9tOQfgke+CxpBLKVLIHhCy/miQhVsGFrteMTDJONKfbBpMMnGcx/Dt41NA/t7n
1KK9jm2IISzEZ8KlbDtyvWBNcSYqTrTgUeYBYpFt0UUGm0g7IjhX/kpLJRMdFUwlaDa6C7KyHszi
BV4NL3Fka7D+kuSVJj98jY0YZsuLCP5EjFlp9Nhdm1rrRyFBrHurGzPEuM7PIYDrRsUziWs8g5Q5
bnJby6eHOA7nfFOjx4r+LSvRcBNLUtipnc968KVeU/YF7Xg29JZC8h6+WvK+9FlkIWSi8gos/h8k
b8o1RENZHQceENFjFzUJoqt7FxYCT+wrAUkFFnsMZI/1HGIT1cSRNtsXtZ8PhIkXwisgQe0hnlLl
65htwGBcZc8SZPUvIxFWGJL1Y13k62Ws4v5bslSHY5mwvOUoi/k/EPIouxIVExJ4X2Z610WG8eO+
CPXPQU4Ef2rbECc5zkL6g+Qm3A61rsz0Z3IaCpiCRaPg9MbZP8rbSvxj3nYofhFnrp58D6+RgaQR
ddI5pGIwp1yMuCn7XGHCdITQSEZbhRh6UP7kUj5NwuEpuED3SKVzK13X4y/qpl2fbowDxxjXul1O
DI4B0zZ9McPGkZ87sWN4+hCLMJLf0iAwOzak8ItSwG4SAwfoRs8huhcwvxbJlA4602uy7BuML8iw
7kOfyPzezVDtXbXNHt9FlAdZBgyct6O8KGJO2hyBa7WuP5UWi4LHWADoPVEx6lfPB+hq/rFG/z+C
XKwGRGG8a+pQlR0J6f58UJV1U8W3xBB5ynYEv5Cc2aZ9WxIj4c/iTLb0LsERrY8/BLJ5b7QMN0YW
WL5B6tznhxzBil04DVE31OEZ3IIzE+UVbSxkMRLm0nTv7vFzOr0ljJq4Cp0VCt+qJV7emu9/2hZC
QHGf7p+wPyw4Dv5E/RhNXwUG3QWhJRrB+ZbVQTcHjUn0rCtd17Kfay4OJmKrz7acEOGaFIrlSwrr
N0U3rZjmeCMnNP628vquVLFOC8e1YO6aUIuZVYx5gtmxmLx23hA2HhxYH6QfORzGubtoAij2VzuO
w8FPVIJ4QXrCXfukUJtAgq0+FyAv4BDYmbeen+XER1qCOm2usoFNy6FJS2s/PLH3ZpuOD+/9aFwU
OCBRpbfx9qaCDckMgeUXRdr5aQijAMQ1GYVBgp3QMx532dTPWYKMFWrySxxleA1ASYSvm4ua/jdI
+EvBAa60nxeSFKjjjyVmUlbd0ud58AFsN+FvtsCdWFaY78Ok/Mr7ihErosBZI0eL/98NG2FKT4PJ
u5UZ56ZoPYQLIx6XhZR7b2VNdXTe/0tj3eKIwimVTf4nA6pA6EdT9/hl3LTyqm1uYlnp+pL03Sxh
u9FnQLPpMEx+I5ZzqKaRHWONsm+zXESD/DtxdTbRa2QlJpOr2e7kSl0/Ezl1vq7gI9an/8o7+G/S
MRSZvHbk4+vyFubP0i5s5wXClycm+DLMoICGtwlUmwX8f4TyPVKxXhX6Vjaal2BaqN7jipqh3tYu
TQFfFdzeu0QqHmmia6WCTQRsu5Fm3/Oew9JKJcQZBnuauBLnOqMz304v15x2SuifmX7E/2OWJuz4
vVmntT9E0hnPtsYRfG889kHsA3+TkppMS/Ov82MvzWqY3CNsizLboqYTXYArvKT1bt9KevEdhrDp
uaVDEdxWTMLTpsppDi1IiWa/auLzJb2wH/WxTMxMtW4kxXtDx5sefPIMjL76AUztPKf7bu+vrtx9
pyq+xvW/2mxiLRcq8mvX9+AYQlJbWGBGvOCyj2j4Jfez3m20auE95Bhs3swepgaIIES4kMf4meiC
ax4PeFRyjr62df9sGjXYH86IviHJCGk9qBNZ3sMiWDrId35z34+HMmxfpiGT/AeebPrybWLU8fbk
sLRvL8lp2RjyYoRtgKTm4lxVphgNoDQMPtFMZgIV5Y0iqu1mIiOiuIB02pY4mJPINfwfT0ALVdM7
u0KCxO9M1vBt6I6od5N8GolCFKkCqF5s87jA8TltxdAX56amPzRGysVpZe7T8ewukWbcDKCCNLRo
NEMSB5btupnJymLQYoRC1vgVd8jKwvjxzddcGXKnNDDM1apH16qP9uKKzl6L2O/KrYjBPKLLkaqf
v2n7csybLq+2onboK4xBQcYrwSPpGrzLBqmwZbNrRDX5V9VGnxm+55kzWQ0w57uorlrYdXaDA05r
GBdxEodCiuJFhvzDY/kFDH3jysjwPSTa6E5MyEZ6QvpLU2VNtQMuYlJ+Dnva/l0iaeAh+2sOD+jz
yy1I+U0F9KA/aB0RHxTaiqwufYINgY0RU9fAuPIhEHdKCQeUHGmBYQy7v10Y5dzWP5vr7onRBv9O
jPpCa3qJnh017UWEDnhup9h5rqrHp+m+0oTPfKTPHETBiqqLkImUs39hYXgCb+GEMJlGhBMiSnlL
Y/hs+KTpGftlYUnh0oXw6u+4MPawauRJJaniLEcxujHtMsPZ7dNsV3YbC+64Bj+1PSsUEqlGIBHp
J+ZW8HjOuMA2ULTsC4o3oO4R8wHN6SYouj6m7pzHVbST4ZHgYa0GndAiG84xbe90IBJDe8DVnh1I
Jg8Bs4VH2vfcWk0zI5s7ykhAT9s/Ib//DJoqoXqdYhf4IEfyAzBuCmw2OXrIXL9no0HhQ6kLqXZG
Ooo2AmW9SvFQ3lNv0ypUozLO2sAQ/3zkXwHnKMNzZ1fxiICAW1HE3p5YXZZAoD4OK2BSlAKHHyps
3kPblPBM5DaUUAEArZUkZSdiuJ46dxs4MvWBjp7K1MqGRte/vnafmz/QPMb9+3i23X6qMCUdOGac
E2ZmeAqZkA+qDS1VW/+82C5c/YuZmEvFSTLRG0KD9AgVzXSst9oaJKf57aub+vpSAKkCOsysxPf7
7rBH/NX2jwzLH7BNPch/akg3u3OvGjarMI6+6oP4jWtUW0uvW2AoyDDbbEtqBtvLI0WeasgHVXtm
mWRiCemiUAQ7z8036pjFym+f6kx+za5wdnI7b8FlBWHiTcqypFCxRwIuGdcxL+13Hw9fgXzXvvlN
IldX/hDsr0POO14lcvXDcR9lqtG1cHRUteTZ843cQcENW0TlWyifIjBdgSGej75P3xOdGtTkFqsc
tU4L9WyUvlrkNMyQVLQcSYgElXTbYEJCbjR6TOmvDwh+SHoSY38YbpDLz4NAsZlu9/5PGLTktByk
bU0u2t+nI1QCHFGFD4KrDf/t/WfWmSORAzOG5qLXLyYUCbHsFwA3MZKteDxtMdI2uZCv2p331tuR
oYwCkImS8uq0elUJOlOmZ/jTMl6KPI/u+9Zt1Se+X8b8SXlI27UIbmCUkayuIn7J4oby/438RgZq
Bq8KtGjsi6uIm+55bvde22r2mBUlG9TNPMWzHGMUg7bIhh7hEVmAPfWxdomuLdu2vu25vR3WLpxj
gkQrjyEd4Wd5/7ldAa8sn0WdLS67wJ2jFe06BN5P8VlPgDhgpwU+AIjRbrDGBet04P2D4SZMyt1m
yRlNWINQm97QuoWNUgGEPDUKpRaW1s1gHZRAeSKDiddQ5EBwOrwZMt6t7dNzHHlxmUb/YQZPDEBP
oaiHhd2K5nJZIXRLAjC9fvU+n013q9I8Ih43hSbl8eudOT77gNUwARMuzsdWXIYmSiD3g/WYYIzH
9tFCZItVcfHWeXrMMKJdBrKtpihZN5zVF2VvqYECslDReqLNzNKrj708w+/PHevHxCbEYsoufNAJ
Ygz7VLozndNsWQfMjZY4o+CsuW9AG7khMTk5C66WvDcLocNapcHQFEzmEAIxt+pkglQtbLFxrgtb
t6f8TaoTbKm8h6Fr+NC1T70Y8JpeZwPULjbj+WEcd5ALtTNRcPSEDQq8YXQwHBo2+jmGZxMPbl/r
30NLcCkGsm4522NZQOrvmSmBXE3KJiDklZ7SC4MgalNJ/twbSh0cvWYSl9joBSMObATNaYlrMZjf
xWL4DRgTFMFbWC1qzJo9vyiantpMXHecovwHcMJo4/dvl324vJ6FzuiTHZ/vv6mGSUqOka1QcdP8
hr1xZNFLG9udeO91TI2OO3Db+vPFf3uSdjpi/BXt3LBfAmC5WXpy8gDSOpiyIC10hrYK4GaIiHL5
TJos24MarYGc3YeqefB5kOFlUKjRgKqfIjWFx2C06cIsfzu9DYXxzdKXyIHdN2f5ChDsuw+lrZ6E
oiJzuYMhsKjYtNjxCHioE7IH973F29sDE1OIH2fgaqVKzy5cgTRhSfA/aZPWis1WGO+o5LS4bt60
jjj4Xc4qAEd9LalCmIItiM1Kd5Y/v4uki/Ckms68G+YzRJAyT3eOelGSvG5kR9hUz2MYr3ElG4AK
nHUivusVlZwVMKhRRQVjJBKuJZtS+0fiSoo0mvoWytHtr+LVwilOFwoqh8eX8JCrNyl0ZNVGKIH2
Q4cR9eHDyk9Sg6BttW/VMgt+6mmQzefx/1NEsb0h3ricvaVEfncHf5cVF+C2TnE1xwyWqh5T01fN
uOrc+mZjBfMqxlLUanA73zJrldX3tjsIKndEBT/altTMaBiHdhA3xwOXClgL+nfBKD9xhi135WC/
Lqk1pWfwUttZ7zmiBpiA4zsNx6jFg0QxAby45FiCGQHz4P4fWR25BePOEjrnvtuMVMbgqdYbQEiR
Wl9Ih3hQ14pzhM95yzsxaAx2+xcOlqDS23hDBDQX+jvJIsHqHOXCzscXNNN9Ij8R6Y0NxelJsq13
IERFUajYlV3HWeooK0S88tVZr4kZJXDDJ2CJ2aXbXoKt5iuz4pgkr+w2jv63mxvVQQ6VdmyLui+G
Em1tGqvOVCoIJwRnHYUnqjdAY7hArDM9CDy78F0JY64w1T1VKYQst0fYjR24TZ3VDm4CE1Dg8XEW
h4p8AGYq6LVoFyMdmzdMa6T0xQj5DV2a+jfZ42UnrbV/F/R2CX7QiIj9hymoV9XcnbTH5flObOeZ
FrmNUe2jmY33qGzO9lcjtyjP4I9Kyb4U6kTjFbB27HPDqNLwB3YM3cjOy9BLjO5tmnLnTvluszus
QkWpedTG/ffURI4/pKt89hCu+V7wRskJ0Aw9sLQyWMANg/2DM6KuBeqIcoT7WR9ocTS0F0XsRVJR
CwxcYqeCdNQxD4UUxmuxYT7T5cwAvyFocfKIAMWe+aPoSluH3i8P83CholtMkG2trjmk+YglN5uc
nGTdVT664Hw6w015x5xT1dsfBhSIR8xQT5ImGdH5IDQrETcOnzlPorBQSEViPbxunEOj612LCTQc
hptx0Ud9LLTsqzU7dyIy4f4QrkvlDU8kBfbdN66pbphPk/T8Jn7ZvVdH5lwWUnZpkdMw2qc8+7T3
HfmwzYOEELgqzLWicZ0Z0g4yf7Jbik1fUCgoyPYEvfGOgnHNBWL9QJoOaXC+hiee6KYC7lTFqa2I
18D9mz+5poxlRZflZLU+zZ/k9RvGsrbOl22d0CqpWvknpdboi/KVqCaUaJgKhFMcVthepcexXsY0
1+FqrXzBo3MBzzS/pLYzpnq0JfO1PLbZHrTr12N1Enk9CqsZV2Lbhw0bO4V3PzM0yprWy6kDAR8v
mQKllTckGqH850jp16k1/vAam74UUNNU0Q6Zj+J9+D+vUYLh0eJLrog3hXuEwRTywUq2R4hd+XDn
rdpxwkcgmo1T9Ni3MBrX/ZbfnuQxUHZQYuitGqjovFp5mVkXXve9b/5Q4KmhVJpxj13RfO1kOiee
jm11TfnPLTMBX60mmfWasJ5hpi4jZODQW31MnkQ4MTCPYBG5os4q5VWR4hCjeeSOyJClxhXaA6kK
YrYxBwsUkjMmRJ2vRgWFVf6F4Ux6J/3r9BE5yp5w+sOLhUDPXgOyZumK22mo5Vv3daSMzHehi0kj
dIW93MCF1YFk0yMkgmOrLFieXCtmIr1sOKUujgrvZoMOHPBTjfDo7W9W8tZq3Ori67sSj7OjPBrL
EqdSBhdiWz4Ef6YT1NH72PdMSx9f/q9Vtm/v1I+H9i6zL6OwMQ+PP4s6rGSL7hEgpZEU/tTN32D9
33NxnQ5ZIW7S1dDS2/quCs5arUn32jaP9cjIIEVFzNSB1BmwriNjuLph8k0skgcOMFT5HgbPPS7v
GfbwgYgIrWJCUOljxFCs10LfmxSfeptPBtHOUx0SacaX6DuMZeB0lguLFA4QxlPHOnspyrYZFSDy
7GvcRsgx6BIFmrJAg9qYj+xH7rmIp3eHKIJUdVT+mEi4JyTm2bwpl7sTD4VWMXEDhy1kNF5Il2xe
SRAVBtcEoBQWT2Oqw86eHOzziim/Y6i6sosMEPsPvfWAf1U7zWK7+8Kc+s2e8ijnPWprA+qJQu+f
8Grzk1pZ+ZcJGtQ5xXZyt8CtaIQsVBTU3ymxeyYk87V3eYx/YpRUi5SEFPR2WvEgweI4oVJCea/b
ESZ5Gj9HgCka+oeoLNWYyojx3QEXdGM9xD8o7tUCRfjRDhIpUWuFUb/TQ+0zeL3MXFEf93BGLhsM
duMdu8kx9VwyFaCUtCFclJl3b4Ky9/L+0H05dTsl2ifxRraJGwPz36Luj5K8ykNq/KKn7MHNteCj
/sQJJVPfr4E/B7xxzvX9xKgg+mxPnVcKDgk0qzr2bd6YK+2NnA2ylfRIaj8JHiwoQFzYu3cvBqks
6e1kZJdQd3YY4x0V4zneIg/z02MtrX1ugLWqsVbnBPIkQvyRy+i+osngSJtbTIiMSXprdJoGDY+a
/LZW+0GXcd2q3b8pLg2VG2IJuuIpgXRjDVDBQJo6sZCVmXLOV+enyeTs6CgRtR14UMSQh5Ig0v7z
cCziazGad/2XTjprrOhkJ8Upx/A8kgirnujMOmwExomh/oNL7I2Q9gUOW7UzsYF2pSw2gEQIc186
J7/Lv03SOzVJd2v0hHCdy4A8PlIjzBhDoYsjfVNfQBOeLNoma3cCk66d8GHWZQta8vOXGv2y5z4N
UeWGV4Ej4od8/Gv4q94f0d3y+H0tnqa9/G0DtnDzadgAhlUXdfQdpGYzqlZzj0XSpa83+BmWi3cs
GRwFK97CYggCv36BLBRIillvEiD40r9CO8eJwd0qoSs+MHS+Nm3oTm8C0zwJHFk7CR/YKWwFLVEk
N+ewnmPs1N8/BnY/JLphYXnkLZCdEj/fI26mNvai0N1uEsj2CWBl6AHDtpkC8qvhSsjv1jG6IX21
gXXgfjGrv1b+9mr4RJxVx0LzNDrOEeK0tUccRh/a4kVHZpRDnyOQoln8J7xETneZWzvjAtkyNQV1
A45Zbowf8wJGi6CfFwswVON6XkaDDS0ZJaLryr2lu5aONBG5/RsbscVLrOgYDB4/pJnCsSH+5PZA
qdct/ya9f/kK9VlWtvS+FnvbkAZrHAG9A0dXx3ssWLVcT76rPcUJlz8JFWYZm9vqLWHbU+ezH5jx
Xq7eRcPe8gpdu1qoF4JsFIgczGoQpmZaDO5n4wt4p4aWOHF8cGOGtfrLKFdrC1HisyWxK0uBga4c
8ZmuDFXZQiTUQMJMNSAIaoyd6aY1bQ/6OMF3pwfNJgKUPP8GcJvtVGw4iQ4DHK1B2K1TOg87Ogma
Z5/L9qXt/4QwbuuIoXl0Rc8Z70wprriltcRuho3s/UevYUV5BnrWRbw6OePChMG8skYKw5BSGcrA
hBG4u33in0b/ZxRk7GjHWhGxoL8QBUIODLVtoQsSTnPb6CF05dLn/ivBlpWjX0UdR6gs09k1VPP+
uN7szre68FfUHE+4VHjoXWje/sHq0cDkcH8B3m09IhYzEE+8YZOyPFbS/2qSGgQClxkap/9MRddw
btOSJk66lLRvhinYMPYetdcLRLD5so4CKhe2pWVUz8PAOqa1F1mu+5rLlKtLnexDxgZ8uQ9zQX+2
iGZ+pw8ptJ+7ozJ0eEoIHzDiRtBBRBPFhRYIRwpdNel6am7ZHaGFVRo9f7Zhez1K3LcULoOQkAQr
wCm+fgsk0H3YG54JQg1Cpyc4yr6dRw5YO2jAZBVaJ2QeBrM2zjfxn3C+M1QwBW/qN+CUkPmB2P8D
7zSZc0Y/ZsN73I3gzk9s5MQpw1kIO2WASuYwfWDh3AqKJwUJulCRgD6GUeI1wXnu5ifNkE+WN/Kf
8eaK/172P/X+jTrdg2d3wnBx22hFFaINCKdAPwy86qHe+zevCTtienSUTy80qXHNbghBtqdoNpfR
m8TRV9XXI2+VuyGYN4GGmY5BWHp+QP8SDmOEJ0UZIhMQP5W4XhkWepL3NDB93ANarXkVYtQXoLqL
CwZmY2JyRh8uWAKLBK7MfWIEc7yGms6KUYCRQAdrt1RqHZg4VtAQIePEXljlK+4pwm+ZN5e03X+p
1XmD0GHMmyxNcUPpE7iz6ZPDxV5cBk6bgJgUBer8JurG8OgS8qcmW+91O9Uy1bhl90u7Dw+unNLN
k6xih8foQFgI286ccPVQeM9QoTxRxVDBb8WIH3qWROLV0EZdrfgUGOkZGUl6dGsu9SP611rxGfXE
p5WxNdJDbg/mxAAGNcAnQQDAsf2GfguwTLQytlwcByWrXxCwHMvaKZilI/iM2KdMlO5MyezJ5UU6
Wpp7D7abYpn5WSmeu7Gyr6OpQm3soN/bRzhoCsKpIum5xqbQhE5ehWs3aHwYptZEFElk4QMIgsCK
yu9Zn6JA62WwlmzSq0KCtgcR1Op9m53uPcTpcZK3gHMMI4p9pg9G1NQdM19GqPKctDgmj6RYpiRk
2F6MLkitE9/SmUGFoG5eQNceNOgd01C9pbBMsGOydDXlyZHwSmNCO4yQfkg0D92236u0oMVQqiTO
PyOUOzmGd43WSD+EKOxMJnQd0CFtUBuGcpanf9o5o2hLRL53fjG+viSRtvFzB0qTLK7EPmydN/OR
AJkdWdZe0W3BHCPA0inj7mHDGQ8ZBrRGju2eISSRa3xZt4Y1TLdkBv2W8xsG63oULSUs99yThsg8
kbMb4fMPFqGqENV26KEtpTLEy1E4Tr7vFYsOI3l/wV4prunI7Jx6QTW4GZKYLEHaJg3MoaAyrGc8
GaYCskkp2LZgY2oXljU3z+kXLgDAslOTtZB16yomzQawlHQeG2/LJjf4kW24M6Wo8pwGHp3HCxr6
mWApzzGxNugukg6dpRXfwKAqp3FkBpRU3WQvCNnxizMgMNrRXIZikTc3Hgkimxx4b51WVYGFhGD1
xgBuNMuAKBnFiQSRpniA2xSx1zXXlDyguJlTYAENO3D1G8PJJidpnIqmJdNpzoBFR2o0MCqGweYa
kcNsKcnDzA6TwMmElEclKWkUsRjCrB7nZUcwOUm0zx9XZCXr8ftJfFwLcZ7aCxatE3ovkVVarsnQ
02aUzqQkjRwQpjsA9xR4ntCklA4feQBJHwWETxg1ZcqN+2l80U8gEAUuitMlLDh40g46DDQNpwHA
1stLHYwdNVUqjXvZEbeYtam2VZtIb/yUB0CarKLSuZirfq8zcF5fowY6w09tlpziNo4hIu6DNeWO
EcGhgk52ggABhvwRun6X8V3fOxO6xesFnGa+DKOFWvCSZMAZcqJXRa3uPfyLjYmTQqryobDT7wR6
JiB2+IhfC4t6wZ9ZTpVgSSwOTAz+k0Zw3nlSRNAJt3Tv56uyroa2MpaBwRehbkmcVs9nMWMKrk78
u8AWu1syNtnTeD79qHJFCLSHdS+ro2abYeDbItC4cVvaBu2zgRhClH306OHv4gA9GcW3y/BhlJE+
E14/NF1qVlAUMXMJi2aBUpA8FX5bL6PXK/YhP9wSzRhwqH7vQVObx5mi5D7Nd611/Dmt75Dl6I/n
BnzFbNryXcII+eF31MvYkaWTnnS+olaEjw4VGmGCeV6R/48eFmQyVilbKzZxlHGqtrDuvl0UmxfG
hRpunTFPRRmQ6rr8435kcyraG7JBRG6QY4AZ2H+ejL2odEJTCzMlz6tKjxTYl0JRlKtdXKkeUCOc
f/+7D7BnanuNuUmiDxM3Y7C9V/7JLFxaKwvLAQaA6AtijhIVHxIxYCxkp1hALgUgod7Cfxm/YG6K
/XrlxGuMRexF//+SMO1Ohr+JHMiMookQ6zv0msIvtg47Ez/2xGes6lmheXt+sotF2GbvO53trfki
P+6llh+oZFef3/IDetYJ66RmYurlR+oRas+6Ir+yFxjkSMBm4vTTlyhu158e5DxCFa7vuWehh4Ou
Tm8rLWgAlCMm+mSI2Kin0m8fblSR0mcO5aPyjVCZhDqKGFeftEx7G0lAsb9Nywc9E5xxPb5OVT+B
j1asCvMMpRvwNLvVZBE8iPKrbxRatRX0lqgiol3pd1h5LV8aItmhB6JLDrqmXY/VjShypUIht3Ho
M3bJ6SAzKriMLsitHnuldYo+nB48+FMujf0A2prad3GMhV3g/wFL6cNjmRbCDGYCkg9pFORbO+n/
CRUshjsyPwOoTHJv/+a5tEpr1lBoTzAIi9LhGlfUEoz3jIbfO/Qz8cTPEEbnOCPCoocArdpisk0V
5DkSUHtcgUoCgxjelkFRUXJVWmaI83EDGqNPxu50DuyR+TudDn8PmMhzuAgBYab1wItyxYHrdPfl
get+6uZl8fg40w5MmcB9IYIprJ3VpsZZKXlNV1LmH0uH4ecoAIfpvrqqxkTgzUFfbQlXWJfrY/eF
fSxe72PRBjea4icIl+o3cVx3SaWS/F/Nc0Ycnv3N9MJPT6NmQEp2DgQLuDmKPYb0YED1DqqOcHVj
+vFs1UGVmq4qZerLIFFqnYWKdAactTfjI7/9MiZibVU6bVtOTMLdcoWWTp0UWXmIzaCj563xRHkw
9sDqFW/BG9gV/bR863iMCv9ZMWlXOVKRmfqQgvqUiui80PL15e48Ybo3YSxjUvqOILYFOir62pKF
E7VY5ZERKIit3zHauisArLJtIeQY8oUF1RpyQZzULPamkF0cRWmw8D/Bqdffig+ALCRLUXlECc4x
TNLfyZXkoFjIH1boprV24EuiVSNLoTwPFFkqZh8o42dWZOnUiKqpMtoA90bqKnoFRyD2z0mhj3xj
afVOJK7jHTLFSEkz8B3oc3DlpiGRVdUmYckVL+il9Ng+udjafkcAXnJRv8WoY9YcM+x7ICks6bBh
QHZxkpb4o61GW2foujyZQguREUbBg9Qxb2CQ20xJjBA7jWmeEot9fOqnyWBxXdk4e2Zfev+a9j5i
Z+EGqxM29TyMPrTGIAKCfQW2yoZOdQOMKSRax2+UssZMJixlQnoB5YrvED/WnUnsIA93Ad6pfmbh
yJdSAJvtDHNRjhVsvMOvjTa/APF5UwPiZ5aiwvqxVJwYmLs7OkBZeH5VDvhvA8TnazEI4BNFwa+p
3oK/X6uw6mBTXr9mDxoERh9LS6YvAaoHvnSy1nyru+vUb6TTf2374VmFDlbA81TgFTq3Pjh/MkE1
QGp7ISxSlwcpoyxsP99HAv006zrAvtjKlPHGsO1Y7ZzLBaYPpwXcacd5ZYCpTyCLIzett3S0mJE3
AS1GWG8g9zYuhGqn+8dgW4slN1tekmEqoFbo+tXy5XxNgSuxVrKUu6uSGAVzwHGN/DZ3m/zVEtkI
dj8JDpQ+WBYHDPjv4hzGqbyRxOV9kcABTuy0kgXxzHNjKuluun+2PxQWMwY2xGiRqwMKdOwapGKJ
39UaM4hPHEJErFxv0Ev5Sxf2nI7KVPYlUeQlM6QbEecljNpdtPAWteA+ck2oB4zYDvBJ2I8eOt+k
hxBrzysf63I6pTBky/xrrgA2+LqlwgWkvtd8l+VYPSXytuk2cd/5Fdz+3gauzkvsUKE719nr0o+7
4CfdpDzZaVoTt427AALfahwup5qGRRuXtadhtXcCvRv1UbdNPOk0sB3QZRxaPwP41PNgw/xqQtFA
B73QCXWnL2JcV4nSGesh+SicM+EbXcOmvFDVIRV0nHn5gJlPHVc5v3a6mQ8NarArIJpQgL6XZy1z
+ADhGjePTT44KnBXmpkqgfoNq/hCWsfBKkvq9TrbVUB7rroe78Bluk/rmIjUYiMJeQ+8fKy1Rr5D
QRDvzdTpBsr63gSb8eSsAWODKIWdI9T3fWHYp4lzeoJNnBezavNBFfZg3w+ibZZ7p3hclPkbJlZd
8k/vANNEFW2gx1yCSmexUgAnwQhVs/q9VHJGIWLplVx5RBS/A9zxSTdYTEb7DFIIJhhClirGXAKA
uTddmgCKa894OrEJ8KqpPW2Mos0PpPXma7a/qQ2BPzjBGcmMx0WH1pWPmxbaYkfghCINCN8rZFWF
5YvkuTXc2Nvg5zL68NYUreD28u88ezLUhsJDQqkxjYjwbR5RIezoK11HYncR+SJC8dgzL8hcukP0
1C1q1xOTA40g08Sm1MqNpgQnIqJDfekMhxoLgnefhw4fHUnxMLXyR306eiJRTBkm2mxa/FJNM7Qc
rXqQHVfeNwdWfl0o47hR07TmfuQMp8b6OgMqmte/GJG3/NcplOU8/j6oW9mXC32py4i4GF3d5JOB
eBwVtf+GUBKjv+MPeClJtmxoA2g8It4rWqm88Y87S/L2Q+TScewWYvs9ug9LoW8HbQcPfEPwdFrM
cTwX8YMyJHYTq5Mi9JbSYFHZjguX52QA046bnV6mtSMJs5Su77+BQbZGOvvY28WS9hSiO3iaSQvm
hwRt8WNOdX20WTrpT1e+PBnj6rMFMTfn6LeCAfK6+N50H1tE1NH0HXl7S53H+2/sZUo/9gJNEKWj
HYcVoxXGFfg824NVmOldPGJv/tmxE/gHy/c5Ua1IiZfXEXJ7fC7EnMmvpqbBVlGIPC/jBBCQiZBW
6ODTQKxMpHxt0qQ1W2c2eFapAFwMxfQVEGZ+qfezEbnXz/QwgD/Nq+6VtjayDVwuZLrwRXRutZ9L
wCptmwJ1Ns2pJK622h1n0OpkUi9U1fk9bpUFi1ELSGWgBLK75MGYOaBEckpMMdL64Av/Nb0k0MfA
oNiurm9VZeFQONtQFJwB8iZhx/FJbPpdlYX7+7PY3jWD79+vXvUgt7aFthhMvoxc8iYlicqibX5r
aWj9oGYGdCjrPTzqCzOYTXMT4Z0aexNpcLjuTsz5lrZEUVs4LzucCQX1Fw62rJEezXzhBa9jYskv
OeKe8Y14V+a/8uTq1X810mVPF+WaNpiePhnRMl39e0mwLDsXZSFTpI/msx7XVTd/aGxhpM+VV9yi
KybtEzbl40Sx8vS0oJkxo1OOYNqgmR4OGOz4Z+UiQjksYkp0MosEjiKRFk3DWXtBHLS1S/Dt+gee
x/b860mvnfXB0Xua8+O7DumBoOUDvqkwWg71wu35KQv53nv3WTCVy8HpyKskYmSAbxlTYuAKrBDo
EuKVi2rD1EnpPmNuR9ViG9O8Fg3uyK5Pn5QqTGRSAjCPVyiCdNNspoJIqjm88PhwJKZn5Ijo84aE
dwBXJULKFXRhL9eJFo2XXt/EbkB07+iosM9+m2QLa21bpM43sj6K1HACVgZQLlSn2LV6GYLrmh1M
95ZDfXgt365iyN4wo5a7DP5FOhbSXWTXD+ku8JhKcyCS57hrYQgikxA8WtgJQzMSVXK5E2KQcrxy
F7xrgB+f2OQx6sPtYPejQeYk/2xXoB5WiWyOpdepDb0RQ4OYRhwNRF+3uOPTCFZIMx4rtfRYKKf/
pCh5YmDWe9I4gwsoWh07RL8rbDrMRAq9MjB8S6jOFAVTbIzwy0chYINCZQLnXFZeuEZIK6yfQs4M
pQXtRtJH7EkSHyPp08n8xyRm/U9qvLNd8mIxl0XNwlvHLOOydd3prHdOJ2tfPuJM+ErFuat9DD+J
4gp2FaKaIty+5ZqeoN10OciqsEzth+k7OSBEqN+V9qwf8UhkN42A/U6KDmnvJnUe90Fu0+eFf5jS
qUPWNDp2ZGeDSSGOi3iq4KM2wRMFcM9mwc/aH+ehMYFUTgzq5GnaNGrCueHFwA9taVUtib6pzNSw
GUu7czAi6N7OMs8osX7HyCacSdzuT8Yz763bkfvQMvBr7wzHg5iE7fFenmn1VcVoizLl7vy/D6WP
jKNgrK3+rzt3E70jXYY0h6i3eu+BU0FC1QcPDHAETkGE41FvYjC47KNlAZnQJlhDLvB4L8jeIM2J
bQjD3rW/2foA2k1zlf8I4STlBgblzU6DGHeQc8+4Yjm+knKdbd9Ee9g9BUjW/J2m+Ie1cFJt06aI
aK9DWp9WEMrU/BiQ4OPwsXLMSU0wx00beS/m4NNeFfFfAQF8EDoadX8IyT348Tyl0TziVvu36Te/
O34V41p7Ypep4WVsKsXWk+cbSD60aYUo+TfvqD/RMyuCIvbMtzPWEC2y3IdiUZHFLCFnVPxqp7v+
dBwz9dnVUStAxNMfjWRbZpSRNUionTLv/0TyjMPT1waB9A+/nVAXynCi2SJ6MvnOQvMJBYRUHJRx
AOsdcmwqmUyNK00UkerTKtZglL1uJfvZ9UVbfyMNVyUHFRxWSkUrh9CaFprT5cWR1X9m/UJR4Yqw
jhWaSFsDMYhSqlgEeMyXWy/1UhKMggyct2ncHNmhj6airoy6sA6CtTYcM0WcunTlU3ayHcRQ5vHm
PoBSY4iZM+9073deSR3tB7f1o3hChmZR9XVhs2pP4P1QlHTQTXOLOqz00mWQX2I0Qb51z5d3aWwC
PdoUiLKOGTz9FEeY2Nic/I6N1/klWjK0kfH/6fJ4+Gpi+2o1d4eZAh6z4vuHEBC/mW+HMn+w3uC6
F7ps2rxDGZCNH0ykgbGKsVNMj/iWDQRkJVhWmdL8lyafQzfQ+ed7EtAAjlfIt0rHIVG4WN/gw32u
n5kRfVZcW0Jog3ehnRMKdoTTX5pwnCdrlIQ2bcdr3wHzsJ1q9KWw973sZ+93gn4g1BUxNOORSTKO
42EU/6cGGJ769rO+O2he46yOvlaSOT0fNVdX0EADbS5huJczZYDRF5AXGjOJgAknWItgQvkGE7Bt
GXd0F6wdJn3JiYa4uEmPfa/F4Q6MZWmSsFmhd50zVQ7ZPOk5jLlG0CsvuDozQ4IrCaCX5R1NNK2x
If3xK9itbZmR0vfXPuzCq/ja/FDo+3d2YisQ9knkiK8hLwfpGxGExY7W9aFUvQW5NurndQyvNev6
w02RcEAygWbZq4So4R9291O2aY6fnkDZjeSbGvNuqNSw8Js0wDnzy6rfcaIgMLAa74AN1Ugqw8vS
+becEAYS7b5G8q0pn3dbR7PWxbexH7Uqt4A+8V7aYyW36mF0oaMIDVPqj5ElXyM50u6t/kyjj68S
mj9ZWQmIMCTv9GYlv9w/lK0vf0+2zJ9oAVDUqTGqPtLQFJxE5zZ//hKocKh3KDRf8Mtv4yLJQ095
k99FCh0BwFz3/P8TShT1G+G0G7seIwQjHBPM9hRnEnS76//sEQO+qdvE9SyYugssuCA/aqRuj4Oj
DrHRNbmuq7KEZ8lUsm6qG5Jlw8zOwoWNYCGaCEe0DXe9Ibylz2UOp/Gpx/P81n5OlBgMVyE19oha
4aj+KOtua+tgqSeMIJaznMZb+Mk+Ru/yt3IxrjdmNT58seXQulbPEj0VD1gX9er+xomJnB3IlVex
6Q2jF7H9DtwiEJR87n8E7zzblhU/O6xoOjn6x57WBojD00bV6nLVxYjzAExxEu0CfhDZ3F+aYXBL
udxl2lvBzXyAznHMQPEa64gSGfShxqXdn2MzjUM3YNo8R5xcHwAdcaXBHH5XMZNPUHn/qF5HN3gh
081C2NXZm1bT8BLIj4hK9rhMqPaurpLrAakSWPx8FKr1bvcrZR7q0sRBmo/gPzQCB72iQdZqlQ2k
aykhAduZxLyCHuMLy7LeqsZkzhFV0QCEAvfHeN6pK1cGge+hRBbei6KgYT7lYmdTVMr4vlpFF86M
s2AbZUecRFzUILkNCN1/Y+PWnmHyhLuHQyjKThwI0bq46hhhrYcW2l8J02HhSzKkf7ct/z40I0Ex
lhf3xc9VAXp3jd+nkL2y1EpjDopNEakU7f2krF4Dhv952TQaDJe9iscaBBM+fjooH+St3RhzdE3N
8WHgvZbrkOf6KQoWFKz9PivXsVndrEuizY6vYxtZ+40lxbu3WAyJ3aXagd/xqiiGQ49Ak1Up/snq
9/EIOjCDkus3Es8Mk3V0MTjM1r474xxf/VHvQ+e9ItkEr8uGBE4WEIFi+xbq8KFkqhVWCgOuh9Uy
vC4TZNynIaipJnHGz1FJkhnrCS/NAKlRIAIuodB7ffu+LNqnizZECkq0Qvv+nQyUSGQICfEborEm
ADbsX3EPk5Q68C4tnM3Ktcmi62CMXGGZ4xo9Rj7VRSC1wz/XYJ3urPzSne940WWdFO0a/zUmtkdA
VZQkT0kOhoyQ5YJdcXff3f7FyV0LG3EW6UpLTPD5Ozly51Alx3fPyvSbCEhCOz3UO0wGr0mJNZhL
TIsItzffvFQN2LO1DyE2mIRLvy85tGB6kEdrM/03F51nxxDf8SsSX6POYEqdPnuCxzFqVaL9+w6T
IUKLALneTpz7Fuv6TW2GeV1B2jZDeruPWhzqQGdxZ/E23oskJJoFjqgTycJOpumyKFeKSfHGhZTE
/DkeZn4bc7tEcuduuLjuWnnqjGUqDacRKeIy57j48NSgPQg1fUvJ2wkeEW/+iEgCpmTfFKQzcX4h
Fad+9+CkWjgcgGj7U4qk6r1fP1vZelhi9goDTf8pfZOeBOfSJWQXkEJ+NCot8WqH6dSsuHySzSD5
0UGgedPO2vqpn7392l1IZMT30dllsMkVXN6B6vL5nymMQdp8suUWHOqpjKr0XYnu146hwI02pFKl
iNM+VeohW2xc/rPgiQcdPB98Eu2bwSkFo0K2dnVndyrMV6vXz26muH2Xlc8pImV+PL/yYhPE/uq9
r/ZLpEp0+vws+FUXkqySeSzXMK03sfdW03T8SH3V0elaQmPMrB24nC5DNqix/Z0kYtTjuSVEj4PP
TewDOvIgzXcDyof0gwxF92bthPQwOLiQROfDQ5WEWrKoNBnYteiARAq2WcBRDRGD0aVDh280bSzf
I3R4JjM5FxdH1/97evgbhrgmB11ZWfKQ3fiagO1cdHuMWVPSzkt4hTe3WkqBTv5Ea2e/zn99e/7t
WoaJV9Fflc1n5JE1Efb4nJMGBymfI3KyeowUhfgpFC4L2gGoP0sY2UF/kkXG6ESWmnOD7NnoL6DU
59V9OryaVVCA5Txd1jj2evN15L39d+DzrAXgmBl2Ss5STOXqYRh7gTLFKUI3HF+KSHHuceqSg+Nm
TlKTmz1L4d0riFZrel8FE5K1zBBX/epOpPS4MZZcPANYRxEY8KgSuayQsOwFPBlFfQeTDKt8jpqf
Mu7RZk0GPYruo1FVch0LQk1E08gd88SvcCpifWAly089D5q724KVdIxHIqoGhsJYHvDbuejsrprq
Ath5XjvFTg74QzRE7lOULt0X2GyPzqars2jJGMbsVg3eAtvoXVjZrSHniz1HKzykdVMz5KkOIxRm
z6jngKOWvf2aE4TsF7Y5JVu2WSM/h1fWPm0UoYtR/68WkzSaxhWMaKfCdx0UmTwYGA4N8FPzpuPc
j5jS+jWyMYB/edBU/V2JzTcNX3xFvDLq6J1FCw6V9kLppORl10auX1xEsdgSbY9UTYa88p8mb2zK
jBQL9THMiuK3nVOJ5k0Lg9hlyqR5Lc+cNsgEleONJLFLxEUp7NYoSdwMQBXOByo+4J6JQOPWtSq2
1ElS76fILbNBZhpcC1sDjomldMeDyScP97DIB46K700lRe7O/Z3hlRsGmXd3nbOgbbGaJTiz9ZQb
8YeC3TwWMceEJr10a3NbuG0IDr4P8ayzVMvr6spzl7UybsUU2kFBqqGOU55Y9kGpxI6gB6KNazC/
JaUmMJNI2hDTbyyAlxf0lSSi2KQjg24rvVVnihdq6A4Vkpb7kl9hGvTkoOIvi0pHO0fgxjL3bCHa
0U3s/hPag8RBFrwtEboSON7VvFOROfLof40w4dwgDK842QSUfFZeuMnED6AlZBxBAwiUsWb0Z4ot
tLG2pQqr7GAekzwYKbSa5s/iyXVXNz+NF92JTQuxyIEf5fnX3wSXiPGhpn/L0WBT9mB6NUtbr0uU
QufoLyT4vxsXqvfdtwxzj4iokZVcikMkSREMfarrbLod35MIKhur/2skiPLFVub1oYEGnYLHVxTj
e6jMmXNC5FhIgJVXTkSJb60cBGAaKSsuN/xy583swL/A1s+oP+yvxWCE6IJ+Dds5TqAZ1yGr+DmP
cdsfPhpyfsIs87rKu6ofCQgN0OtjJsLizBzcPrOZOnmgXnKHVLQ6y2NG+UptkHlDQ0wgtyOT9bQ5
xDTXEgYo30RkpfzY2e+VrlFh4XfEnmmLGLDWrpVmq9Z/N+5GYnPndjc6WSmXMFqBP7j72uojJEw9
Z3u1FNlaxem3k1Hc1n+YxeHAKqXCndVBEUFRRgFjd/rK06aoLCSfGyDJhRB/yE42DcVCQLKWoxhZ
Wpw/+di96YW2zTeZBcuGdtwJoC05PVzZJMjs4Vy8YsLm5OK3LOUj40teKqG6/oBO9/rY3ApmDB9L
SQ0pCw4VvqzgrYK4QaLnWVpCeQehd2i1LQaJL09dVTcl94I6S0iA5ue9kekiFIcD3QEWQvUbvZ1U
L0qhMxlHzKoTpx4cQNdrFWU1I5saDUbsa93Jt4zgd9IkPPjgy9CcCM58g1E4AO+n4cO2bZ8qFGwD
gmAKRZyRJEPUryibqtTfmBQvtwnbCNYym/8GUX1ytiy3o8e52sMAxtp0GipbuV6++N2XB/nfjRDY
d5qihM+NBKamQZDZ2zJ3ve4hP6O+1zvzgLl1ZbHS2W87cJX8z8yDf2EK10QK8h0ftgnSgXxKN0rQ
Tw4jWMxkTJFEUXvqDRsyriAw2f2KM4Dr5lXWvoSwJtpeC+tILjlSO47BedwA7PQcdrh42ztecGcE
B1BcBKlWkb3mrjkC84Iti102HCofuwfu6qyPZRFC8p8rqpLqAnJK5YNRU46YBLi5nDn4bqcNPNNA
NkSDHEdcYIsPNOUPAawsUfXR3CYCzPRWtw8Z54Jl2ACJLmhO4SQrimf76Tl1MGd+JoajlOUnGFIW
qZvEuPvw1R8XCUkv9xT9u7qz4H5O+nM5JTgq0ZSuOB4whzQz3pXamlWb/7Y//oX/IDsahk5cdw/Y
DaDyZBNsYBeQ2mB+0gU0WBHzxqkAczFjsptCMnCGl+agJdgnVLUlQE9yb98z82R13aMJylTHjpOK
69pAGYaFQvN4GB+BvjWvqebnEtyARZ/UORJb/q/Yrs3dlV0RpyaWsFySr4NzBYYzDYAWL09BV21n
SDgTtZJNoY8/RTDesz5yrUw+gG15WE0UdIwhh7LIyzGXLZlKxVeQJ0K3/WcaR1Gt59TgHUHEg9dX
6UN9TtcJ6kbDLGyV/7NjwPW/lRT4LQp/NrDlgYMe6cUvpr2D35fkTyxI2YBDgkdVpsCkXLtH7KzM
0v/7HNeZbNA60hsJOamI2mtdar+lMaVUM+XatJkKSA0Xb4KZTWLZHYXWXSOtVRgOjoaWNi0iUOw/
TtqNc1Va22cbQs4+1qTCHuWtf67PWra9UHWy32F1yA+1ER4TwFXFCdrjPpYR2IAMn3UQ6Bjl5aP9
cKvx2T4+UqsQAKdofXQHy3HaUTF6D7WLc3lY7bgdkrj39vY+Ptg0Homt8r24RX0qh3rKBDEZoDV1
ZFqN4LUQTzxXKJ0KYpRS7eHEZ+ikOflk1RFZrnDB3uyHVgL9CLy9b4FNyi/funVweEEZd0Kp4vIr
dR/VANQPGTmRWs8IVifB76DALUI4pD49uj7UbQZkp2lUBfRa1SqTk2dxnCel391CFVHEXMzTF5Ky
HR7G1mu85td0kS1TLchmoM2eBUNcsEa3dRx84kux7/AiknUB47cR+cpOSrU5+293ED4DYXXnYp69
Gk3S+DgAJ1cX2EWKQhIUxM0yKX2fK3TcqHDSSzhk2bNznskZmUVmUK9sew5rDF/siO5MZc0TKnWQ
sp1c5T2Uy8mE3/XFHmrDmfOC8R5OJyPxSa06nBp1XzdgBPlxOcPdqvNR3+CAFrTT9Vy+XUSEu6fs
hWpRyV+53zzA+xVPAz+rqN4skCcL5p7yt+jlpqiY/iVwKBfH7unBvyLqb0UTNMcW6EDtZe9ICJ0K
UoFxE97pzs3sflF37QfzlE/dt372TcS5EGF9dkTpOkTwAJpyGho/e+UB/13Nf5bmuw9Mn+1+o8wT
DA6o36vXA6emcyI/nB2VDMztbaYhC3mGalrWzcuUOz468+VEl02nzY5Ru7jEMh5glVyYFC0n63MY
1P/he6Z+npKO+4VjNYLq1bLV72R/QuKSO99Fe7ZGEIiiuTmYPoCs1mkn+h0Zekmtvua7EiZ0NRdg
ndbtOL94/gV0hE8mzGuYVMBsl6QBxxu1344auFF9+u/Xf5D0jDzcnvMGjjUnileh8FG31thz2igB
Ydf7YR8qLP1WIjz01KGi/oejc8aDILLytfEKZEzgzcgxx/+p3lYLnO38ZgzkK8IdrOmwntVKCRyu
glrzCBe8fESOLXXAKz3i6ZUDNW9yJx3c4f4U//i/f29MyqZbxGBlnz8e2Ly8gNwiFk9/FYgF6y8L
cTyPTT8oe2d3yVrb+tYF/F2HKO1gvGIDa3kiGKrAqsSsIBrsLGom8ko4ifMS+2TurZ+YgHFqRKLM
LtZIzyOW0MJcMA+itLl8aryXbYCpDhCFD6ydjYWrcyPKta+o3ggtiQeKvp5ltisb/TDR8jZ01mhL
0+Ssp/sx3AfJo0n8BbJt84xnhytsLi08HOWxFr70Vpm9nDCtY+h69o7wP2C0KOF0w4QlGBLr5LKR
9dt+7ptLkNfmRo8YdikB0NxQWq2QwMXKcJ5pJpnRBxQ2gSC4QLE4IFc1mitsTphvWmMScL9nmVv7
NF7MospBPfScM0ElxoV0L8mVsXwumGtnj4McOEzZdOx00P5UEaAe13/THxUZh6yL0JCqHv7+XfsW
zwX2rE2tDlpSImM95YcrtHhhkqsHGX3X09bXRijpzvWVHnkOXNlRF4OfHWPT2iZ4+i36wpNRCrQL
L6yFdMBHn7QPi6bTIbvj/9HhyKf/ZfoVumYJMQFSromtV0Jk4fMfBUZTBxUx5aeyUIb4DhBhyBIW
fnXIgNWzM0qfJ7cU/xQpcW2rFZ/eeuusoAnD8ht2LcepqEC901/U/2MkrZ6UzxR4N+obxmcw39PS
Z8cOfNvUR6KDWOjdLRHsqWzh41e0LHFos8zVduzYUoc0lCj7k34LqS1jc7hg80//wL6ytd/pegTC
/qz4e51E+FR7X06llWuR4jwNAA/zJFMdTrlXsvVNjQaUz0JBGup4G9ZLaio/Z0STMh7QuvWsEcXU
T3oZk3MFT46qhwUHJ1XxoUGzjT9ifzMupkvO20k+DBCqyDMJ8OyzHLAn6e7hzJ99vMUoqf765Gsz
sEIfSM/B6cG2C06Nrs5LXChHJrzIyu1uCIjuJ8HmIQK4GuWJLQ754DFI13Ys5u1nnFIICe2JxIRH
ZGTlkfFHl9ogYPWPossebZFSEh+uyGNimW/3r29eIS4Ft/ka3hyGCznRaoiXtyxxk1I4xIYcxMay
62yg8B+ZImdQV0JOJ7AZFDoZb8/LISrx7Ag0z3ZlQVy6VQx7aVcnl1BvGsY387hhE4Sd5TiMj3ag
/wj+71mCSrylY5ur+Syor84ZQUMzpIkYp4oq1pWRvhh0GeHrInS9fmabMUC/xJu60HQ4XN6iHDLv
VLMkFiHdH675+jtUtac7dY7RG+a0hxnTZ/mYJ+nDB/5dJtEFQsOJJKKy2+X4FT5PBufMvuP76XR6
PdvSqmrm9gcZIfb1mL0QnNpJ0p5QcnodG9shv/sWydRKkMn3kI1H/IMBaVNDNF89o/CSMlVJSS4D
v3Vh67WTnWvw8iwHG2pmRWWkOQMRQ/S0p16oba0MyOPnesguZVKbYUy6s3NiH8TD3iM2QVjqdMCZ
6mDFFJsahivc/n5F32N9fDiTUw85DXKLcy/A5q/p6aWcT2joqiKy5mGifuLPLvGamuDpvTdPBhm2
QvpF8qGVWedJyFVprlSlGUXyshXuEGDb2daPMjG85rwhY4ZA/Zhjw2DeBFCd7QdOXdTXmAupumHq
AdzpoCBVMIp5HlJPWbtV148y8NTk1RBPrCjkZSPS8T1prIj5v7pUhbb7cY3d9NYFCjaG1hoEaYl5
/Y8BFJJalc2J95IuoImxLmAGIVg0QbamVJh9jEfTD5G5IjsJo67uLyXGlv5OH68osy5F1l12xl/f
/E7QtsajS9FUuJoGhujOITxXnTpIfeJs5CSklGR427oLwBai4rU1tWNn91FZf59EHfjRxpABISfJ
/YvPeAXpQ/gkxwl+HpJz1AMO1VCSlKJd7E0OhckCBG+TyXlP4pLjfb4jBQJCeS6Rksk5WqJAyMxz
ErgaKE6xNCBzqZV6skHetGOB0f7ApTHJeng95pl4gKgoG24zAzMQr3VANVIAEM6rCFrz45of6e5e
JZKqCAbihepgrrUU+2+G+pf7H6NfcRm+fB/aWJnqyzR2WNBSgcSpTQ8red/9qbzlAtKqa/pJRske
xyY2ZSOz29ZRHPqOSTgnZ23WCe4uvWcWo55oRAJTp+nphvIL74a05ZoDHEiBw10ML/lBDT44hXtJ
E1yOGswL9ztvHztficxtVergdz4WGmu+a9EmKyFZh1NoKz0FmyhB6EDqjoGGNPMFy6NFKFrPTRnp
XivCBMH7B7z0jcm2ulIdmtR7pF3KxJCCJDnijlu9tMNvbyaQOutJi1bFGvP/VET26w9aGV603w7X
19QxWMJQZJMLGPIcTtsniZ1JsqikIAbgMa65KqDFsg375N87tD8Jxpdq60ZDDxYXpStz+VN0iV42
gofPjqttLK9rdFaneCSvLOTQwigzCnqy6X/Vi7iOMx4O4JINMHmpCOgu0yDyYtSckA3bDmMCOAFo
ikYhAiB7YFC94vJyeL7Oyqva0VzFqbzHSGW+tmaVr6IYOsY12yOqTF59jmvsBUmKnkYYoZMxEbKo
pWzu8Qx7+AApr8l3tY0sScNHNL3Mgcv/Z5YN2wF2JgfiTGb9dv9W+jv1onkJhYCu47+sFlykVnMU
rDCSnFZycF3ZTTARFZ7AMdm8MCWPv92EzxzrsQ1oKYGHlLDktcSggrzbsv4rgo1llbuxt5/AuunW
L/9YvbWeubiu6Ve/ZNPt72gqu2EmjR6MgVbPf5X8huCDRSJ9Lupl9vqbpLe+0+QdYT+BqVZ9Fdcr
1I8nLTazNvsnjTrYhMNQTi2Zdg+W32d3xUo+GloLOjN/nZxS02LDu53MzcYKS/WQA2wwi8kpRL76
zJMGfA2uokJ/QzwNwcGA1yDJxxQW6zmOpnz9pn4EFPTUOS9SfL6Pf8f5JMgS0h49TJgk6gOq1Q95
SNpbg0POjEO/4qaaJHT4ylWKfwSeqhnkdrgTnnPYZSdYzI5ThxUpAdHfHO6wbDMw97Zrr87eF2xa
yOFV6UZmjCX286kzv33CDnUO4V/E/VxEZcQPOp9xv+r9O/cy70Q46fnV+PsYE/azoIJ2k4sfhQJL
WCV1Ymq+QGeDfz1JhvXimZQ4e2wFwWXhSZ47b0V7l6BMpTk7ve5e41A8SPBJdAC3EbPKz8FuJG8D
hbJM7scp4JjqqDQXkB+dluKwqSlCYU90jROdPhqRwX4rRHXVRQBTl7WhDAih0MjEDGE6A8Bm8UZ5
vBrTT2KgWF7e7MdiRxP3a4mzyiv0MH8zvShx0tnC1vJDm4bnFYN5UGB21tUIYxUz/T1t+Tj5G3yy
Xd/JOdxon+0dm/vPgmeJkEJD1INS6EgCeqt5dQDEME+gkRCjYh/LNsnEedOE/Z8R1eqFqcMFIF1w
Pgwyzfgd1hqp4rh066y8yRv8Wx7hpnr7NKmzfNEJhAUKVylhyNzm85zsLomxIbJ70WsvUOnOwbKa
gqYpL8dGI6sI5XQ74Mmyc3iP0lQz+hZ5rJfR547vTIr3Sf51DrfIm0vxRGGDvfctBTI4kAavj61p
oG6l9Isrb39RMh9P2eClLLXSK1eWESkXbw3bGaw57sy9Oa4Xd/7uGIJlmTc8KQXBaQBYmeXXGE32
q8whwUa8ey5SmYvsjzB/RsFpkxPSuJvG/lGAuknxE9XujrveJXw6bmeo0ozhomfw35+BS9at/Y4s
b0fXt39w4U3t1nkFUNe0PoHgYVTYrbZDs/e6CW6VZYMDDSpREPU1m92OsO4VouBHjiCAGFcio5ta
fnAn0U7/+n/lVt9CXpw7gvEHVuNwC7mll2NleKDdmG5C21FzVmwbpPZmsIhXxFljHZXRm7GE00Zj
UfhNP7b9Z14JvvhVzzrMz3+rjm1VueNqIDXqJGH9YUPMA5VBZi0WBeOdXzA1vn1hY83fXWv016lX
irl4euuwuGz3fXxbNmYsFdok3LX30DnWWXHWboSzJKU/93wBkz9w/tnKWczs67IzbwUlRPsAGPJr
z10o6Qrvr17dmoYqKEXTNw7nGHvFuHxFSYWe10zylb1nFqwbZm+mkyvH8xHtjlgTEUeBJL8LJXY9
PuK4+5G5LV806IkwjL7n+BAR50rYqw0Ku6i47a48sVzXLXkLrdEUBPhuGByPwxv0b9quTEALBLSV
Rtwn/nF+Ir37/DmmWzDqgFDYCYyAGFzczEsG7gaISamjd4wwJ7bkE4waLL/f+FnykbBlIQF6c3Ug
I8k7a6sIL/2l+9s46hw/FSaVb57XHWL/2hVr73Ve6h6kfPin/zM4JvwuQsqma40C4FzTRWsvE7G8
6mBsFYDINOXCO/3Tl1UCrLNGVwXlF1xJXPj4vYqOd/EGPDjRtDh/xIuB7xqVLSeiTJkcBB0bQjnq
NYwovVrQPEc68nsvMgzWEL9b7uV8LFJgFg3x6xsbSD7hjrROtOXp7XGYOTFBJkXNNuyzo+bEPJj6
mMGScnGtoRDvw8t53REH8VZMsjl5j6EkRGe7nA6G0Ranqu0Zpw5n7nuLrFbHVXewXy4KX5Zpi1gK
7qwbL/QuYxtag9leopBhthDGjEwdf+Dg9t4t6zyvulRsGxZmW64Z5bEaQFiOnLi15lq2QYmOkzgU
oUDwCWZm4BWC3Bqt50cG8WzcA+VHtVpPCgvlxA1q3/OLPy/MFRBThuYj53gnSdhJHAE/HzQInv7C
1U6M+E9EF6u3ly0k6yCVXpTIDYeML6FMkdh6zbelkTd+P7h5Ab/o5RkG0icfjuLcfUTEIvtxXyr3
l1rf6f0Fgtk0VNNlO+wVS3XsnevKy5cnPOQjdFP13fr5C2lJL0MdirCDSwbP1dSVZh7cNWUbrk/n
L6FmFyZaIDPpCJzkiNVcE/6UHEcJ8Xu8QJxb3WywQ0g336OXRTQNj5Jl8VtyWcCWiIco5D3ha0bk
6Q4k/dIptOat6k+aznj4CNGDfGz4+1VcRkP5sv2EUC3xob08/5E8JieZ5Xtf5WeYtPf/kyVuESsQ
pY3FHveN/dQKXtaOkVtr/nmUF/hyzm+mKwgerS9wnKvGH+9kdWO6ROn0QatAIrFS0s+7Adkl4aDa
fQ7Nf9XhtgnqINbjQzy/REOoXfO3r4Z1IlSq8N0v32PKh8cyPwK3PhjO5z5YYlM/o6ym0GNxQNOR
lVh/HVDiiLJauYhczRMvmjf9vx0NRErkiFonHjnE5rRAR9hoMYNN6LEdAQNBb9E365xBxXlyLE1Z
Ct4K9s3q/vQ0nIxSwUMIXjiX73HFyLar3SomQnCoscbjgpefwPAQG8QWVr2lWam+LzkTpKfNOBoj
2iOPJSvXTV3Uqq3cdfm7twnqvQnCtwdXmPkRU/NHQnxG1l4oCiiSwJwIgqkAWLVNCKVP/gr7UtQh
l2GpQvoiLePJGRwjvWbn1tHnO6o8QdOWcRVaqNzhQmhZF7ot4vBXA14W9o4g5SGpQ5fHzCQC4WWV
DuUb2umXTYzVI/2QfjGRkkYE6Jc3f4FawzJ/uBw7dbUn+e/ZI0yc/d0ClhAweBev0EBqlIyZuKXw
ArZiPoZjmrOLbern6uXMCNOWBFKldoV6HHn0g1tYm8OSgePJLoRkgezEfdjgae8/ZpHRzgrSUHxD
csxEYjLDU3RqSXUGxigdbt2/WKpqNdDozAtYy3b9ILS7yLxyMO4IPEB9UpBq4dErVYZ1lev1WWf4
Vb5oBBvx74bX/t6+3IWrqtcgbGXzP3Cr0ikkCD8Kc652B2QX4Lr0kDXVCt0bqWC/i3jrXIir5oFk
0wVwtAr1DpwXUsMG1JRBkNSGEusxehgPJH5jBHQHSG2rAnMZk68AXQnS2auydrmjkEN+5U2xuLIf
rNnFDnPO10PSHdHZWgGNAv99UJSa94DIkdSSRZHwpFhj5rW97AWIXoYVjXdAslbHT49HOVbbgF9j
N0tD+elCnqxiHOhmQ4XlMYUnLsoA5chGOeufMp4+V4jsXBM3YuJGrKIfWTKjzC4voYs6qqwvVcGl
IWQqiQTuF1KZky+YSXBW9OYYpQlGL5vCmsg3Mij0+RyYcy2WkXWIj6H+9p/L381fzC6XvKSeeXaA
f2fjSmK61V6862FNovxUkO7UFr0hrAglWVFbDW28YnZg3Yfne3M8bsEhsWzgikjB4So6hs9dXdbs
t0/djb70oKFnVuFLcDB8Rs2wHHmnbkhNA+XB/w5ss24RYoIDJc+Sl555j0qYXb1ASCkixlART8UK
eiWga6NLM58Y/9oTJSPqx+XiTeY8c3qPXWdK7yuqXqGCgsTkQ9YIrFipkDpKmtlBy9xWhyzbCuLX
M3Em/DdhZaFbBmbDx+ZP/XtUpBPB2Pn6sOwZGMjWzY9MrD25Z6X3xhkt12Ekh7NyArvCZlR72P3F
tRVLA+wTiRKpLdGCcwYtx00iphTch3D+TvSLSI7CIFOv7ONdcvYRQEA0aqRLKo9ekFywPz0oTa2L
SfgguwC4EDQEWV0LeAAD8MqzsGUORX4ExuNOlZWhEtWNMGN2dVHO9ICYOAklaEnZWjJu2tujmtBB
3ieHufGaHXSXmFDz5ZREPotRsTnby7DJkJKkggpdN6WOG2YMaOb5TrT5HjKkiCiH125RMF+Jxgyw
n5Tmij23mPQO8VPjPQHCycDSUfBhSncpSIRzNNVj4qphrS0M4J6JUwMs6iDX/b4EZPy3dYKFsnoJ
7AxjEuJPuCPZAJja69vNCgsKgFOb6/52amlRJcBZrxXsbBgXmsmSZDwts9OXUiuWqMrLQaNjtwth
9OjpBrOvCE3lfqKgcKa+dlT1RNrusLVLMmFHcUmYU6F0LMa/MytZbUz9cutjkZoABqEoubOS5frW
J8fc4i8HHpTz3LlTUSpjfvnpoe235qJromfiexPEHY5T8bNzIz0wCnTIQKO98xojWhzZXfzLoBwB
UrGU4HTJPjeTzheCBhLpBGXFLJ7NkTgxOCDDPisEvmJARwTEWrgY2L+eA0eUMK9LajSC8NzaT95k
rWcxoJvmPEx/c3DpQCr1yKw6V5TwBRF6SErpP73YTSyw04KlipAddvVOcoVuPeNwvrpcVhJxjqIH
zeu8tNyPKJ5gz8+X5qTBitefGk4TZYS9OJesW5xB9+uPGJ6+MJNCaYXtW2QMg+k7jhymgF5m7eTB
2PxUhZX/iisiSJ2nnat9SSn1O2KltZHg/5ZrVv/At2HCHvXMGUu1mYtbBWUYqS45krI30/e50oxr
nm+6J21Z02gR3Pnsp8DZmu2PlUuTlsyr0GnZQoyh9MjEzS5+Aq/XNM0de38xS+ZyERkzpxcsaGtU
CfVutXLmD+ljUu9b3sjepIjPieRLQ3tOumW3UkdzihrucmNdK5niPRnQbQM95M2Nm9IV0kd8KBkt
bN4JSpq7ZbbtlLjC92V7FooJtCEgs4QPgt7cky5rSl+kyhyjEJ4CeNHaWq/ZCsGKV0H6Z4APS2a5
868+4rfZrTip8StOeVNCilnXMEeO7oe2HERxxF2u0sFw6R358c4IvMyQJCk8aOtoW2Im5EVEi2Un
GHhDkrzxgPTt2ZDJ9K3uq1X0YAV9eoouzTIqPtHRulDZWtk8REZN6Mf5spkTuu68OQKVj54aFJFb
MTsZ0SKu1ySC+At0v8DBLJK/+MFygFiq2YSZMrUE/WgZ1whQ8IQtTuMm22dKsa2O3Zygnmp67K3r
KMKkPQLa1jittjVgqKn9hiBGPBsvRO4egSKGf7Lzax/OShnn/CAKPqWLljXuSve3UPSaYmp2FQwe
0XKqkeWnp2ZdbQaV4tqBEcPPA3CfgpXhXru417d4NBz4WjPIwtGHjF85ijRB9MZNoDTmEJW7GIeV
EFEjoyfSgwnFkZeWTaA3vbhDW001BlgwOXI6ck0pJfGsOvZRSab7PXk6BNX7TKqpFu8LuqHHWXuO
XjeKYkZHNIvvjsqBagCQYath5DC+UdelovXRFsxC4G2jZFNpcZyd7adD7V1p8B1gLw+RX7Qqxes8
j1r23pKTTNZCNAxt4KSzoHz0awGFmIRAUxb9jL3Bz/ZZtZh9pxd0ukcBYlCtZlpo3bCiqZGO0w4w
0eSF+uX/4Vkw8CE8PN3T/jvB7DmWfjBjC+2J3Vn6+RRUG/H+5tJf7jJL3F014/vRX9gI3xlUHb5P
ywRvO3wQu1C1eW8iJVAqcrC9CKmrBxYlpW5ulJzW7QMckWZGcDLwVmHVJkoZsWe1hlBIuhhez7Kq
/5z4wiwxmyJV3CTRACHRhh1PWZGq1SwCc9PxUrBWdrJxldV3YtRNbO+SX0jH4IaLenoQuh6Ca8Z0
wz2gtUtM2ib32WqyWR0b/pM1omOgGvj/i7uByus5XpTrPdEKH6yw0WOWwrG5/8RLx2+EObEMkdZ3
nxAQp4CbChyahavdpIPAa7ZSKjESfHKIFHfiINj90PKmgANibVPmcp0JJpJyWa/qIjALPPBl/BeW
Iz6OBMiWuTWDq7E+97ypfIam4/1JCJ+D0MNQ0ILr9VED4FfU2t0vhoa1MkcNGsNmoLtXAdlQ1Zpm
JULas3cWAfqymXkdRN6UEiFV9aDkj7iiFfJ9KezGniJIzYCra/eR/MkyH7p9kzj5bESBOREa0QbN
Oz3iAJWNa3szIF/POxiTJ7qhhm4olviXPrZ6HiyA58yrkwM+KoCXifdSpfhXd0c3m7QD+QA8GBL1
ixkLtmE37NXUCUgVMUNs1ppzZmb22EV17kbSPepBelWO59ryyeZNTMSe1qU8x3JBaVrL5TUMcot9
wiOuz2etFUoJCqQl9RvsIgWk+cwtjKGk7ivCLwzMt6CU383Ufw3uP85pDO5jtraj6Y667e4SitLa
CbZDMonN9yYJsyOMINUoK4PUbzndt+ZuTbvmip2/rxzsMMB5j/7eFO5eKhaPFTkdsPs2vvtNzDQE
rsOfqOi6mufDQxIQoTb6a+vcK14FSrerd2tN/r3sMs7dlbowM6Xgu/IcL9om7RW7uzGdLYsoKPyI
/9FqP9N5rYS+hSzRwW0qjnouP+c0r2D+MRsMhFsQ+NqcTh9tC63zacgNgvp2kMbHfSaYdYBoI5id
4lagBIdy7WkUODLu8CzOna7SM95G+LxynGgTUH095h7zjgnpYWImhxJAQK77L9RjCvBPZnlXHOQU
Pj5s9yMxWKNHF3LZX/LCMOMXxPR8uazOxUpUErW/YIULkYQkqwNqHE64gOy6k4UAFWdwwh/Vg9Cc
U/OqL0TESNoh9ZQUmV/pzW8cmMS0G2oNwD1+WOvVcqt9I+P172SAKeexFr7BXAGd76Xbzq1A03Xf
6AiSXQChhhPN+K04Menlt1zFetUThjwwCUOvKeQSONg3c9kQtk4ilOn+r35meQ/njHw4E4yQAOxz
fCXvcunm7OTj8oHE1kijcxH+N3CihmMIRdfuzQv/IIxt6QqtHCYszXo03Z5u3gdm6yhILCZJ6prE
hqSaAkYH1xfepuTnvQgmE0k7ZmhRB4g5CZ3QjApAt95KOqarP8bnXT2Z8KmDel/RRVpIgGsHcpR8
jlmztkVoW8GUTWMjtGw/nCrZ/gifem+Gqe5X+r3NREJXX+OVHBmiACfRpz5qzgwYXeRhEuSDbg0+
0OxhChj01gognk4lWn7P+VMWQ1B4EBuF6amOSExUQxTcIdFjG+mLB9nVtPaLEz4qLuMV8vDYps1T
pIVZ1pcWVkKbhGT/a6/J0XzLJ4DaKws/yxz60bsLk2myjpuuhUB5XK2pm1yl5z8gUjFJqBa3C/0D
HrI5e+Wr59p5dAUd7Geksy70Cq0jP53kt0lNrNcodS7Mg6lVdSdK0b4iCwtJKF5FTVMMJONoJEt5
39i9+MrvzaTIS2tqei1E4XuC42MYI3yXGEx5hTGCkpjnWRd4vRgViogOHMEymzcs6gg+b8FJUzGY
w2tBNRhPB8j6g0d6TAe2m/jbQRIwX2/n1aiTs1Pj4tuJV8UNwAqniYJmCy8FG0Jff52At61bFPPi
yUgaiuhd9m3iPV85V2+UsdXY1QQWg6cF4eBvSFUb+QV/zrO12ZrK4iQcSxopPlskyH+yZpAZ/E3w
sL3yoG1b3r7tsTpylOY9uyQwt3nDyh0Mihp1vhQFdMcfPoYC6SCaEkl9LB0EF31kzlOBc2c5nspl
YqX/U58WgG3Fe/2B15IcGAOJDBm5WyoTdlaMjpnzNiZ9XLTvfgK2bsSS6A4BUSfyh/qQvydg32HO
fHmzRxdwIkMC3XKoNE0IJO9iJxeRdr6z//f7bE4hLvj7SOKBER/S7Ey6wtrxV6OjRJPbckapupoY
0EYLqgERT6X9ZaOzPO8R2FcqMtnfcd6yKgohS2xvbk51y4vS5Y2KjGKsmMCeuTmQiroVo9q4aHp7
OE/vDEqM0OsZV5sMEEKkftvk+EyQ3L8mTV7i+UBMldcddp9kJeFp0jL8RRHWVaWLahGppQNW8wbI
ba5HZddaR0C8OxgDJTwM+nyCHVd9iA1EkDMe5gW05+LAwhX04GO81IPqvUssiXYVlSGUFJzwEj6E
AvBflxyMxtVoi7F7cAfY8Xg11cleTSBPlsHvYie3YjSdFykDh8NjHrRbVLzx8SVYUPo98nGv4G0w
g84DV23VY2ZhyvJYHkDFQYhsjWS5uY9W0t1/bdzVeCdj1MKc6tx8tZTBdVPq50jmph1s+4vP3Ftv
pO8jprCkFNW2Thp8jDLOkwKnNR1NhkWvDfsYhKkdkmH0ja+5A0hA/Mu6RJGhGyQ7DKc9rbzBIoIw
7ROLZ4K/ULF4A8X8VaAv4cCaDCooaW0vtb4BiqUL6hMBWqdAhXeT6+c5eED7h5K5wvRcA3gp9mDa
vLcLXQatoPOd/um9nW1YNEbW/2aXOxZJ7az6f3/P4Z4Bos/ktUScQSwf96JpA9x2ZgT89vfdFAas
F8qYcHpPu4TeZykKA7QPdKilYUPiiDVEVPW+s7tkQM0zKZHXtfrQua8la/69at/aVHdRi+eXCodO
4ZTSIKiiF/2Kfh1LG3by3pBzfgiBeKCIm2IS1+C+bGBzoPaZjvfegJcF6Sgq0aPVenr6JtPdkAnE
2NcLmINiZoe3rAAIpwgNDmDqakfDk47XQ/EAxXDmCnWUB3CgdgKd7coD4pWlOcyqhNmUC9ixYr+c
kifcFz8G9qKMxdQP3eoHXvlZAo0kz9pIrqxDD2EGf/dC08qY8ktH3eeSbC6MT1H5i2daJwf8T6UB
HpiD/cxEoxedW5iuEFyEEAkGz8g3VvcnAThu7h+Yb6Lq8PchGwn5lX94qf9sHibDYnK1/hV2toT+
6LvZ/H5Xbn34P+VmW2KHF1vgOMss7FZTaG6Q9b3HTagppU3NrsKPzq7QVzR4IPiHi0JxKGZa3AWF
hy1vmp1DfcUM6jk4hJmWhc6dzbbNR8Hsj/orFu2HkseU8MaPxh8ow5+dsJJl69HArs6ftp1UqCUR
1meM88Y1y8dj6hF58gcqZaIOyYTF+MFUNR4mYz44AwZRR+t4gGXRvF9gchAlPzhSrAwUKfTAjObd
v0NB9SKwo+jQfj5Y/EodcjkWhoGiuTXNkLsdKUl9NUGYb4+VYen6w3SH8QNmccOyB6jyMNWrjlyp
tXMQABVO4WgniKBUr8CPc3U6ck1OUSrZwXiOiWZlaPNR853iNixqktJy2tgEaLQWU+vT0ZwrtH2P
nxU+E6VYWMnKmvtMZul3LzoCHv1PnHplD1FOt/jhxa2b2l35HskmDVewE1bm5V2ZcRYQWpUDJuuO
/f5cWvjKeNqbRLl7xkzYZCgo6+GheLScvbzp5YFDb9ILi6mkq+0qAQ/cogGw7D75M23tb8Oeqqi/
BD/XJY0jT6wOOS41XXk0tzb3pI4JuKvnJpyo1STfmyAOZ4Drr4dG8C6dwmW0G0ldc3BYcvhK6gim
ZVyikfho2LdHxCqy1mzBx622bFAA21bLLirOwSGXW2FcfVY/XGmEcwuK6Bpk6To5G9WXs3I2IHUR
Wo7E8uZW+xsGGk7eFQPu/Bzy73knOm3IMGUeUPTRTZglNfHfO8AAswbJDwRNcO2FUUOb0njg2Kz6
UHjt02ICxmHVQt9mHgvjXRfUm1ybuAtNZslaTw6LVy2Ayd0QCeOmn3v2Y/yd90Xq6Ifv7qq7Ea6L
CnrIR2YCsDCvkOGRN+SMbX6up/d38memjaJay2uTojavHY/9XbWQeP/Il7pJX3nnViBavkm9A3/d
4VQAvJgaFQ86YNlRyCYgC1o0ASlmf8LlPAgpVCKOAYv/aU9q5uuiclPRZOfabe3lScOPWiwQyYli
BnhncUH8IaKisqNvMi9bxlfjLJN4FuFftJ4eDVuzSFePYf5p8Rfv8CtNyOMdFQzmWZlBXZlyCX4d
aQEKDpTEOcG911h2orPvrftrv3V4oFtUSaLyxWIJ242GS1dH4NbnCRgoE7gqbSNgN1p7wQ06efA5
CyeE/siIByxyxV7hEYrXi08M4VwmPgq3XJ0HfUkdf6A5OA583/cqhhJZo5px59ruGY/hfybHlCNr
Bz5Y+PkGn3w8o+5rb6xnN3lg4w7lGWfnbFD5xdUp8dPT+/ZCxnDdrCFXsr1pxVIB6mUWaVG/43Dk
vGDGJe2odDhij7dOS1CFtXlS/8kVkbEKLVCRcYqYTanq1X/45udWRBsp4gIbOEFdORpJX81mQgXm
jrbtIdIWHW2ynO6SMpOiWJ3TM30sfHGBsQWnfxxcbDcayjJAPhK98ne0yA8+AyjKi5yocGaO43z/
dJfGqYPv5pDvaJR6ExiyoRbJztBDmFYI7FN3N1EXYI5y2CHD4FbYQHi3LbazKsTADVmicRSt0SQi
Etg9cZ/MtAg2f9tHmD5MrIKC1KE4cClfKHCIvGHtkSc4XOgJEOYDxdB+jKUvgcx0AmGJxlcMkmHa
/DTNeUnJW+fsNKqDOIHxdljFbWtH+J70TEbP5ORdol5S1cVbdOBLh6cSRXYsNGWrm2OR0yfXhe8w
rcV7Qf3qvG8OCY6IrBQNlW+Zq0+KSURFIjTH17q+T4P+K0H6OT9j6ttqFpd2yoQYiv3hkgs8N6Nv
WMa2ymwR6evULU8cDxfpTPUQjHcigFGR8sON8qKRxAZ4Y9s8Dib72ZM6UHcqZ2M6IYxHjbP+19AQ
xVSpu8Go7/2CQa8W3j9Jp9viOcRj0Nzn6c9koFrpqBLJHOFZMoVPtrQjHBOzTiDK5gwpxNZVE0Y2
DssiiFQzj7C+bbdA9whieDXqNAff4HKUn1Ma90SWZfwoQV38zWk1gBndMsRNpS0AElAafuAdZmPe
EFfm0GT9UKWncww/VwdT4yihIUNTElPIBEV9TCR4cBmHFrAvR1ysHkJ/sD8xGtUaUoOenorfqBzX
efxKSmDMD8v94nEpzJEv/sifyg7Hgzao5Sb7f7+BolMmmAOMk4oSv3NArkC4hOqC5AWDVIJXTotb
W8CdGVMgi77B6Er/m6yeiHotzHuKFhc/LCgZH46i9CoIyd1bS+Mtz+xaq5RFdWAnPs+puaE64coF
gIZ40xGTFFydagdnTbmWC3Vo8jjWJKphrqyRScAoViLoAOSXcrxyaq7O3tL/9E4Iv0czZJC/wzFP
NiRRb/TWQ/N+Q8UJ2z5X4xIOC/9oMYSacfFpmL1VFX70FIc1kznqCbIGnQxC9cwm3rHuKWTBJBac
QUAYPv1rFhNcnPYWsJsho2a2JjUdm15U9Cj/pFLG+hIVSViT+FcrVlWX9Ue1h/0fbcNSB3H6vITU
ch8jFYixYZLaqPDSmMH+9Uy9dcnlLe51i6bX/4UfzCvaPwOedgsFuNc52x5Xk4WmXZIXmclyNfCt
9BzBSt5DiiZIlQscwekwtvScDd4CbLiuQDdrnGM45bgs9UGgjfET3vCTMoSLt9KTgYEkX6A9GbfB
SSQTnJpF32F4QebrS1Eho4THfPownvqoQT7pboFzzfIOGpOf33M+ZwMDTEgKJZwcuNOsPSSxxAS/
Cu+wLCmgsCINaOEamdiBIp5aeixiUmHCcw2zyziM0+hmZLdjHp7vJR1V8nub+6syr9EMMTuTGGmy
W3QBlbpDlbheiYvnnD0vqtCjsCuJ1AxtGmnWWCP4v9ON6kKbEuCCc6zfgV9kYLRqIHVzrvLgC6gn
t8TlAAQWqtdWRUe1SwxihP4PZjTuLDX3teSi5YXRa3qSB+2w7gFai2crWQx1xDeib70VoNBHllox
zPuPFgURcfSi1SMy5cUQ59SkEJ+0Z+9JcEXKnZZO6G8DQeRmH2O/jdE9Y+Xodw86u/vEg8xPKQfo
bg40ajWiP5Gg7PLsQ2ys9/2IeIlLhSxNfGO9jhg4Hnw/TLyeZ91Ancq6+E+BuGLqZ+StVTSh2+R4
zWcI0bgxfraltS3/WLrGl+b4EEsb5Oh8lZf1lRYHBAj6r6KT9TflrRPAUsKxLw1rZGto5r4n+l9I
7hFohDrU7oJFqkxdhUIDpoP5fdd/l8ZG4I94kqEvwI2pPDoOcKJxBJK0InD22V41/97Xq39SjuiH
Rx3c/g4McUKoco4IxvvdSJcuHOI6f3BpckGmxrmJlu8dsP0UTYZTHK+huaXLhVTursI2Ga1n6lg+
XT7hSv3aUITpXv8rEx2IC7fRdu5eGhOWPuANQXngY+ujwjiGWOoU8KPmjpzyeNsCV9X1L4ks2Mi3
k5eEKdMGOQHWiHX1IhOyRmnIZESAi5+dxAbJHAVOnigjCl2RA9uPNTrjYZTCwfZ4VnWfSHOzsXR9
ddILJ4AXCaggWi28LhK48BT7zegjefapmFIy+0ner5hK/7cyWSJXMN1OI5O22OjFEEQ6RUBidR8C
H8HttMTVQdHbJDoOB+macaWFjHnFwwRwYpQYboEtTosJEUQo3E/9EhqH+E/btcLtE7dW4JFllhqW
RU734zVtgFzNYBsMCOwStXfCJI4Y98noqaesOvQKrOXL0NNZdp0ayut+EF3uHCqFNEpk8iWPRmQ3
WJKSWYQFsciJP32hhl5CvwkEQZ8nr20K7C2A/1ZftSIdBbRgY6C2K+fgeXeGVm1x24+feTthJfzx
Ik8A9axbpS8T4vOeu3nkRdjKqjPSuP4YUEoA3Hgh6vcv5pMyeLIcwngueewHcDbi2Js29+KoeIMm
u76XOKqjOQVxEDIhEfiNyxNL/E7Zwe6Qjr5LkNwPxaYSVxVTvt15f6wgnLDiB/C4+5Zsa3L23vaS
nLg1lXNhyI3oyVP8KWGQqShWuj2cYlXUPc9S7Zk5BSQ3jKtT4OXqid/0svitR3uCYZXOuQM4FAwm
y5BCTK1slpY+4CBype1AbLBGDr3gNaoCbZLqvn9XWo87dB+Ef9A2YggI56vNo1pinaZRXGlmLEaG
ROyjOrWWRXeZ9QR+1hQmrQa+Uq1SdKkXZ7ql48hgf40iBqFraf+Qk2zAIUB5pdmosFpXHm7u1O3A
t2K44+r1ggk7w0Tb18f7Aa0SdnL3w7QGZ+XcETLI/C9UJaumjNMNdkA3Mp85HZy5IPlLoJxQRuaS
vipHT7YR2UfuHoTvVFqHrUpG8ltnLm1iJz1fj18OOAqq7L+k0xXeOBPB3qI42HaDAcCmwhrhgFrd
rMw3PyWHKpoqdltAUjEhvTYVFXzn69ttAjlnAPtdfoLv5bH1tmx/c2t4eMbUH+G8gXjQZIJdgFQZ
0cYPTLx/QGRkUD5NTEW2NPT4IIeyzDjUAUEWLL1lRC+incrqN0x4B4PTM+dxo7MimqTsMC8LrXlN
rWUm+orwvYk1rWRSJt2+tQjlB6oVrFxQa+5TWI2xyud/BrrOZctl8TBP5r538fVzmxiGA1V/B3Rn
N6eoFB2vc/KRKpEhuLOq8y0E4/OqvQtIEQO0bWqHRkDj4Zz2MaX1OdrjDfaugtAuHFN1Y6nzLc0J
2piK9JstycNTso9xAKn2a1EbAjjgxrbHPNXvbbSLsDRt+eqxseIpaZ7VbvKWA8bhmlQ4PO7mfiBp
ErhZqEK0xFodkBi2P8Zu/oTVoHeKZfPOnWXRxaL9re4EXUxYj1PK765ghzdGLtwBtbF20K8wICCt
HfamFQRqF7QDFpd4ewbt6ec8NqYD1zflDoGWUJvVkLb/D353G4ttKjuzl0lGYpzN7cGDYPj4pgpo
8Zn/lcbnxk9xM3cl5Vqv+K5bNBq1dPuoRnkG8mDSdCrRhXYBC2aZG6K4G4J/50punZpA55M/HZLF
Kul8DGo0oWDrPd7aosSRyavQsZI/lQTwGG5zPGnCst90oJljYwMh4M0ltYVnyuzNZyYGhLgEovGT
JtySwbw6WVydIaMoZgXXpS+W0e/CyjyNyuwy5nB3zBVL5WzkZOFB3FFKPsyxPfT/OzZbimYN18NZ
YsKhSRpPnCPk07jqVj3HlKMPBNsPRbtqZ39IRUEhqbQU5+muwGfQm+Vqa9zlLj5eO8EzIJdmlR0R
I0geh26X3pJSQsOt4zp7u3LgHvp/XNJS8LGDIByXGvzZ/IsTsxj8ETuoXTW/8Xts2MKSEwdGKPz6
ILEb66t6Q/C0NZeQp2QkA1Z2/p4TmL/bRGaI6vkfXiIKiUEu0Ulhr+ZesNj/+6cdrvE8EfSVs1AA
pPStFdYlqdNIwhzA2oKVz8bxWq+w/Grstk0o2Ku8nAz6zRpqKIKumo7yH/pqfMORueG5VXr5cfzn
c9N1zpPMMh8qDbHMMDFs3T/FSNNcu8onm7QJL3Ul61ZV7i2QE6cmS8XOdAMvg1Sef42PGC9/VnVV
4xrfPRRH43Ix49+PstA77Pz9AXL3mpSOp9qogjVC/AWaJqehZ3ID7K7RgcFQcLqWYhLiV5SdJvAv
vAMzLfG79vpkGhz/6Ds9m03CtjIsiP2UmONW1FlaOgZsqpXz8DqOov1At7V4m4cMs0qmsWr/9gL8
M4OqZmNXB+Du/8YYFoeriMTfUop4TiT5Ris7j/3huQYa+6vInFwm2+X11s9uMdFNjCre/xCHSg1W
Db1loQUo8Bhel+SJKYGUIgyffajlUEZFoZY700qqXTybxQ8I5giSJ3LOlu+VteDUMMWnerOoQuo5
KNAj4mZ1yap8kIdvTuJH2zC9h0gzyYcTx4F/d1AXz2/jv1KB8ZFmreN3256voJwRp6fcjFD8qFbh
LZKYivUU50PLI6lUFTHRgKlAPfNWM9yus6Bgsjen88zCgz+Y11J8J9Ywn7+WMaGn9shkg2Tu1LlB
Djz/mnYXxkM2lHJY4KgHlvi59AnB04++ImtPszkGfzTXDNZFlUVEfEyFnRzMbULf2+AQBvkAQ1VA
V9c/11Kzf/ATt/gRoX6dV5CQrcU69G+ScW0H1RKtiGP2oKicaXcdMA35I5acv2RbzU6mqoTwRdTX
m41Z/ny59ECw1QZNkPyozCCc36aZtcbqYuOawBioiSuOK0QPqn6Ow9JczNNaVGTiilbQ2t7/qbR5
0y1d9tnd58FTrExTy7eRBnGnk6jlATY97KGfSN9zQyb6X9/knHal49AT/D5w6eZpceFA7aEmebgA
obs3QkddV8xin3cgYsX0aI0yKriTXzwYGtY+QlSWIEMYBxfpNsT+joDsKdyaqkC0vE4WD4wpPhBW
Y79OqYDPtcxA5NKDEm/vZpxU8/NcWi6DzHCzpHr74H1aC70HGvt7Br/SLFJR9ek6fCvcNuhH2ioy
X6Co5lv7666YT9aBwUrZWJ0bIWlUkF5WAVdGsrj+0GNm9uWgobxjyaIdOjsSF3Os4yazSLjYRx5l
7mdHodDL34NzKvUtHawl+Oq9wVM/zmmtcmCpUE5zndclAjwd1kemludZ/IQZQ6CClYE2Bx6VEsZs
bPINMOIUouYv/jgwWEuzj6Eqi+XbSIz+o8UpSSv7Gvs5BKkntUFCexFOsEeVH166FLJRcfmPMdX2
hXjI4H7FHwoM5tO4lmvZRUm9wz16Qgd1sRlpmsHqGp6PXZA4R7mK8g5V8nSUo4+XBZ+zIap7NJGO
bzYeyJ8SI7KFWTNJFYJAlc+OZiUP4ePD1DpnvuKYv2kAqcEoIELoHFjEnCYgIJGWAzHHYIDAa5qr
ksauLqMSaEjXLzv1Ng5Sq4BxJiEdPe0+gsEvVwPf+PxJJ2TTb2NTIOjM/aj3y7pPOugP0E3VbLVT
CmJrRi6izTvZLIhCJdkFIZn+D8OzK8WELfD4E0o3NAaHuFHIGTTIrSbi5WQInL8ff6Sie7/UnmMH
uDH2lK44X5c9exnKtkza1KOeYxdAG4QKntmE7U8q9MtNSDhSltsToF4mb+LB51SyLAl0CmORvvxG
lVlSKhMLi9R8F7w/kSpsub5JYlafNyeQjGYLbUsQtzOpJc4R6w1TyKOPo3PujmMIH+XDvdSKX28Q
2Ybtp2wmiQvmVlPCxjaUNdi/crqBLoyjeumOegJDeCJR/qEWZVh7aUbUKhq17ZsxEia3y4f6cT/o
HWOivR3ECrvGqihGHbbQ37xqcfIyjZjLaVT7Xib7Q2yYusmXgNGPiuJxdMnleKacKVjdUQBDoxcA
XuEJrC8T4rzlkU3KN+TKsDvmfk6z2bW/r2Ti8EwLw0pRWpaCWMYwbNfLF2V/pSh7A0nZx2+K0vYk
swZTQnaEtokemWIUpiRLuhELe0CZDo8/X24dbFcbrfW5VIlYEBbJBZeI3an7DrSkcTAbe0W9SEl+
c0IyeDG4KVvZ6SW9B4OGQJLWl1d6DzDt5PokuKPuGuPL+npHWOw0P/TWec5ZTbsAKXiqYFkGKvCe
ZQer9N9aiBfraKNAuIqrRe3SrYyC8QxPb/78uV7Ibb4G1FasQLlvOBk3RWJqia2jpWsO8cq9f8SI
0t3Cil8o/X5w1J8E9kLyPD088y8npV4jqKIMxf45oVpy7DG/9GnCmAaemcLvGRPmCa11Tjr3v0Hw
QwITiloQLEy7sqYInuBkvzFDjx03fk5RUp4lbK/pXzfEXsyHiJxBZu7eYdtUeX18dF9eR5jhruM9
qJEak1Swh3hC1R4iIixA5aVt8rK4fAEO56M5D9BD5ObpSX5A9UXOPjDTp6W0ZaF1EhTADm1dYVzO
/Q58kmk1N3lEyyOw3pYkaSR3usRGveIFyufXsTACSYLA0yOLwfSCjiK+iUxbrBnONKqQRt9JsKc2
wKI+gPi1hpTqKvih8UZuWKF3pV6KLtUUE/O08XgUiGpFCNp9S+Sih9qHUk+YYeDkpYDknzAHAG3X
zjA7dOOhPL9OvoeDh2dyDjUMCuOLb1/3zQvUfl8mqx0PTmrPGGUCZ4+BbpMudWjdYhm+HDNlTWFm
oDIwqm6v0JJ/W9T3cBWOyRWrmxDHd8toTujhmpWmshseyeXYUVIY2p9xA/RajDGR5Z7r0qlrPQDS
oAgWBUp8NH/I12Ou76mPA9UZ7SI84ttI9xDjwL9JeE0qTnKH6K6ODpz7EjXEz223AmIhyJUW9qQS
PRMPuHRxDi2fS+UNLkxYmr12ubLQ+N4vppWi6NSNuTtSE+iJLKa/6hdNZ9qm75XK1cZfj6S9L+sU
6TqQcwWFAIcQkzpR7ZZNlIAA3Oi2OXGxM/wlINrv62J1VMkVbygrxjVviHRjriZuM5B4AuesyUn9
aQaR6+U8bAzsucqttJLWSMHB/ldKqwMaRBE1uxnVGWFe189NDYjDfmIews3+tsHfZi/ciPJ79j3X
kO7HLvzUeg84L13L31mWwIYJsRKDXHDGSjGj9YiRBmQNS8grZBScyZ0QV43ahPW+nZfNJgFeKVRI
nFBM/JmFa0YaigeKJVP5Tv39fKCCB6pWAgwTxQRHUBYmaWnq9/eViak4oh4lkFGE2rQv+ryJPxRd
pKaFq3WLc/CUZU1RuQCZNJ8UHDRaNJG97G3/faW6ZqPgd7A/SbP3YIivvKDBx2YDgdyt7lV1TKNs
BiMQ6z2Lq54h5mHFpuySzK3IPT7MAWMknhtXWWZsksXgbKUOtsWEFyTnJzHRdQ1eBGudw8YflqrA
flY28aZKpeMVIfYrrZ0KuXaI5iCXFCRlZxHdrFYVkf6q00i3/CNKYZDjLgnLYxhF3VJTwI+tiGXl
09t/9iH2/hqo3m9hqdSxMEIIEvMCMFu05pH0oK7YNcdiaLJc71QmgSDZHVjjCbTj9gxPKI4e27cC
t6cKJFJMcHX2jO/n5/rrk0KxUj9icj1mTNbundfN7FJYQS9nAIlC702EbYwONHe24rfjhi1yi2Zb
nemAvfPnmQ5+Ng3Xo5/4RX0A8p12tE6tbkZpFGZQ9W2ik1f3NwBeco9w6pj9VHstsj0yv4zCoJAQ
hegZB+h1AY+PxuteD7sMckWfcSiMxbmQAUeAyd1q6NUX3PJOUMGEKnsF0GMgbsUwneIOHty46t9W
E7YkKCJ1K4tJ5g5V67EzUGuRBBd8Mf9v1PUP/OAdnR6waT83/g6sn5HpcsGWGRZpQBwCRiran/y4
LQYynFn1/m0ylxIgDm7ZLlBPg4zG2HKxe7vRMPybguIggG9FXJqAVD/954ZZTaTlGf0PWmRELAeY
qX2k8KlypcDEaArhStPDiM25fVevG46CGEDtAc3rxmjZr4KNBMtQfp5ZeCZ1x1H3RUjpdPxAQS96
YcHSlHb/FWgoIC5g0DQb4dmG+0sRmJFZUvUU0JNPU9KahjL+GXK3DLsa0qyG2pRlduL8C63aG5eB
5UZWaWoJwOgW+I5jb0k0kUt/u35Rpbd+glmEoYZ7R0b5dhsFDfv4b0kwe3PX6A7Wp90HujpUpNlh
UuqMGitWZujrYbRWXCRr/wlmonbHwRUSZd//VpFHRZ6aEcV2YDZD1K5C10zHrDgxsoYkn5EOYiTQ
J0ylcpjIa+Vr5cnqSx3Vilv67cx6VnbnX+Ps8RjkCKBxfHEdj9k4QBWZ/OU1X9n9ZSw/LbGqCb56
Vb9tYSs3kXQ+E0F2BYQWJL5Rx7w6lLNvSLyabhjHG463wEVmQ05Dgn72q2duq1BUmnCMIeNq3r8l
9QNUsE31XIKQ9KlLHn6anXhK21QOY/OHtYzBd5+0gY00sIUCFEkipHgZuXuzqUOImCp1FzJL7k8e
HE2RRPhVjTFRX49pguneOxDlB0qFFY+t9XLUwRJzqN+3xmeHNSPgV0pPRXRlbu/yPyRsfisbx6E7
cfka/ealwBKFdlzYGJG1M+hq2H0Xolp18XumAXQMcI2h7Z1lvC2sb4KkjLVSnNAgJakvM4x4AsMb
QgTiRP7QJaISeH/js1p2OpA25QReR5OZnl2Y0aqPleq9hxmAx1qDAVJ6rq2SQ2/lMDcm7dSHD+ZQ
Dy2E4aTPVKqz1qYI2Pp88hEkonGz+s+trNRhfY0k2hrfmqYXFTEYb7rJGylzFYRcGs3+mTSFjHof
XI+iNcm7pCLZmNOqmUnEKW9zZp2EQ0zumQaZ/+rNg1Qvk9xGa+hxJJhiV41Tx+8JN/3/yV6C9TMS
/BjtdFiLkrlQadwv+uNp8Wj6sTJn8RV4/jWJ8jzLA1e/rGesAQO7YKeBDmszDmNmW+7Ppy9O5rbI
91tKfOSvmMFHk2UA4TAUs2tcTuxx0tz26YXJVGFORN6sbEL+sdM8klNN1/Ylur+hhJ52RG85uVHg
IG8z3SunBQE8BXklZzdn8igIPQMClCDTzC4FzcaZv5RFzS6+zqVVC3gS5paWlsAD5jlxSUFxqoe7
DE1lYTl45EaItSSg3YToZwSZEB/psPa5oH1jx553egoIFkiERdZbJkqkoPUjxwnVvWuocZ/jVyZn
vJ3fA+qM7yQXbPnwoNNoTLzJ+c3xvdchC4mEe+wDfdYPsE5FPn4+blEt9LSm1x0KIlG88sfsuKgK
lPU5qmSu7HwzONDNA7NfCyLUBl7lnESmMlfxWzI9EeD+cyt8ILUZA5SS3wsa5c000bs6763yGz22
BRGqE/eRcDFS/8JnI+KuK6mjN94v9+hxmhYDbrBdGFd3AluyE8neZpuvyGnlYI8pSKJFhMu0QOEu
hdCLYqjYp4AxDqo/f23q0l5ItL465wk88woklRIWHE7P4Li9HdJKS2mMO1gfqZKYzLEIjgRELhX5
pqz/5oKJk7SpYGNum109VSMg3EIO9aJQ0nCDtNbGOrba/1yqFCqVlZXbFl3qhP8dfs1oqCpiAf3F
tn3lI3budS4e2WiDE6LxX2NDUwpWSMDVY1NQtaidKVE0t1EerqMS1EJ4RjOmsOPMmjecRVXgCGqE
5ayMlA2ddJafXEOfWqGiyBFPJbAOv4YR09+fMWmytAmamLEBQ7/L+38kJUadBpHoPTXRyuTLVWfg
KhrIjb6hH8clWWBxQ87ah/rgCEu3sBVemweHkF0DfXkIyRT9k+thqrA0SzQAMv0/WFGB+ven2YJT
JFAs7nQuQFYwaVMGsOe8o3HSZnAxNI5820+3TpoQ9SOzrhDYYfSb7gwVGB87C1mL5zqMqjAxob27
vOKd7Ln+bCVhvVmB+eIqLdAU6f6nelq6ZN5PKwiI3wtMTW92kxJo3+Uv2X+uzoCYrqfQebs11iCX
ApVkQ2FgZ+ivYLw/BLeoPqp8L5/M1vhE9CEB45TIsTuNvjBOC/yBM9xNUQRZz+bulRfvSdaf/PXy
wZHZSeC+nq2izMgniw5Ej+d/pJW/4MmNnmjP2dl6/SGt6UwvAr0t+MU94liZ31QnaHPbfgaC66cN
pIcspgishNxneXTEByoUxWU/M0nK3I5YCgy5mitgs2a/R4bM/XH019WYSm2xIv2eyoNVVqYtK9R/
xnGMxkqtE5eGkZS1LJg18ub9wf/1jqP/as46oIgZQlp5ey1Xb+ZbxM/coo6ci9L6wh59zyH9HWG8
2doJ3aRsidRoH2wLzqbo0KytVT0f/BtPiU3qI1W+WFamDqm0lvcTakpoz/WMzrB8OZU5JNbtZp2/
36JduBcbtcWHFyd/s9PNDufEL/RAhOA8FCJA/lpC2FQT95LW1UuEF+a+GFbKZuyPIrrnLIbo2r7r
4vL7fV7kYSgdusBeLzxtroiOyoZ82B3COX9VQGfPrVQtYrin7Qka1rVMgmAHhqQonCB4Zhp0ogpi
D2OetdsYIraum29gaGzptZaRsJeMSS/L1QsAbuzBVGFA8oxlFSvQIqBtvrBeH6CL8HAzVnf8dbMu
maNursuQCgXsWXOo6JM+mOciEwVut/nAWuDee7VkFdkOW2Va1NVi6lRF43KzWDIzkWwnIdSLoaW+
U/1im0UaiIukiOleELT/PJbVWcup1RNFOxFSRgteNMlkkbm2Q0JlK+Xo8dFJglvJWsYtVTXi0m66
UoUvO+U1Mor7JkET1i9SxOVRCe4p9gskXRJiHvBodjrkV/F3OpwXLP0Fo6WfZnoDIm2xQzeMzr54
XpabQkcbTllcsWTNGykkbgTEd5zzE212ynX7Z5oKKpv39aMhdoCy0sTXJ3s/kZk3RaE26RRlMpy/
mATWU8VsHrDOfffzvfk9gzDtsS47dJaZYiG63G6ENAfWIK2MmUCGjhrX3Ou52bQDWZ6bTALEmzdI
Ka8QjABWWhFrKjQJnMWtKpKBi8k1Aj/w8/GonwX93l3PTWv8DkeCTQ5e9vFd6DkpYV3m+Y16aBca
ADKsdiVZDTPRuOtWEmMp5gaindSC/0zBBxm/3was1lD7BZUlsOe7NEyosmarIVSixcsbfmAli8wa
8zC5PbTpJYe9QtkZlea31XM0GgbN3CnaaGATbQ2lK+EkK8Hj3o0Qy+hAE665DaKhmaFWRQ1vmBsB
FdQG1Ov4b4E0TMgHoT2tRTwC/PQ4OTCqWNpnFl2ycPiPfqxJ/z62O61dKKrXy3tHeSr7pPfq6Tb4
OASsqH1E6GIlZK3SCAomGXJmluRDmJ/tRUb7IYoQsK9rLah5ATfUoVAlGERzSQ1LLygjUQILcbF0
qKwFQnFTCFpEHL6ZAoS05x0NsqDs8nU5KLZrvsHyUkNuf9BrlEcbd9Xyrb+wePMyLPi1VOyfFRFj
swQsPmo1816NrdM6nAHSXo6hXdCGj/bX3K/LFga3TbafMuJCxSnIyMtuS9rz1T47izhFLdW/6V0o
1wxaYUEvO6BRHhTHWn0ac2c79Aek3vU0sYzh0hvoYoMJTsHhP6YkCvY/aj7hz3OV0qIZVMExWvtk
xnxx+UC0cMzT1wSYmRXUDKWnU2AgmB5iIFZXyENttBUV7szd7FqKAYYoQ9R/b0r0pmpYh93OrZwb
YfKA7IMp+9089tYtb58OssaESDUIRvPejZcavA1HC1+HPgd5aasPYLpBDcguN6EnhXpo7Y7ZTUcD
iN6UJXcoxl3qNm6rjYDPmBq/PRdM/YQt0kkIjWzfdZMluEw3dl4F/snPmMsiY/Vju36h9LXL/9pk
nzsMI1ldXJCsTnGWzswdLA6/rKuG49SDKH8yXmJA9l1+Y3Jlie5V7LVLzhvAOTgTDtFl1N8TTLMN
6dJwPd6XyvDMvQyS+O+7btqG6fP9aQni8kzUULGsvphEvIFN34lRha2+7tmU/Rw0A9gYH/55KFXu
CeFwmJeZVa9OyUDRSpWCyolE+C0FmEM1FvE38kL6e933XCKgQ6+XfWFvOC8pkifmoqJ1jCRDtdZG
rX8u5tc57eo8C8FHEoHLWoUUr6omJv26sQ/veIi6Gl16Y6CdQwjQ0PiKQZ2Kfkdc3TSZ2umImcGt
njbhO/3X+LG+8pm7sh52ia/BiTr3ZGUxmbAQqh3YLHNi+oK8Ne2T7DdDf08XmJb20BNk4Mz5K0os
mKjFL9d964LHRgOGAu7jx/XIESDCZ+FBXSKBjLO3uRT7XTPdC3jcwvL7BmqeuVkJ+cyAiloGSlEL
56THkJS7PijJJUfD7b9uRag3DLRZjZikSQ3KDaDM08ZUxpUqQebPjsniwq6PpFjTM/nIT6aeBhtu
JbtHeQ/dhwk1yHKLsRhIOETS6wWVmzbEy2GpraxrSmhZ6R6pnBV4wucXkGlvW5OO6tp5Rbk1I0By
LOgoTtPqulCZWUj1I2xF1je5CMFMMvt8fWiinTm9UTu9DLEFu7Jy26zy99EIiKfPIXgOuC8TkdEG
U9L9jQ5lY6bp4FUzyFyCLu/ZwoYpaFcHteuWbHzTpinc+oF5yHQ/BhBbR26Ls/Ug3XMaPSAE29zt
rEeOZwhyDSlU/D0g+lAjApW5Wjg4DFrJDGTjyuS4Y1nMUvhwAT30J4qMqHDXLjfhSqtH4pDuGl2C
NclHyqym44hvTlFFsczaXWz5sz46n72ui3vqd/Au6Y/kB5XkUgGGTvgMKQduxJPS9pwWqpoGaESA
Ic0N26xX2QxZLdlE/pLrL9ZPFWfDltnaeq/Is7OyMYOBbGmCEEsCN+C42v84CbOFvNMJr9GDN582
pIquvQrlgSeB9Pk+MMwTii+/KMJv/N7pSYkAbRT6AJji50axXU41RWrS4rPuJllyYzxM9VxrLh/0
Al73dW3qn/cIJnfHkAxoh3+XV65jxLN0RKz8rICFuYYj8GlVnxGIv/5v/mrc7luU1dIgF84Sz24E
jOZjiZF4tfQb8uyoDgkQsxXxLPU/MAtcL7t6P6OE1c1orYEeoDtM/QBl9dutkxQNNeAHOKDgtN55
0hLghMVrlPWX1JcmexjUWABIyN4QC/NT210UPv5n1y/hcxZhG4lgbXLRAnktQqMNSELwbc9UlKlF
FLX1dx2HO4BCHMgKfz3g4EeQ0BcC3/WThiD6Ur7j57RLfS1OK9UYPE4uRowgo5Viq/tqZq5EeGuf
7mKq0n029NUDwqR0bC0GEa8qM6eN8MEYPeH9wrAKLH5f6ZncWgYukDHYy1v5hY4CYkEBCaEZuy1S
YZEounbyUeSHiWZjxceSZQHCqFJpUYdsZ15iXMd76jtb+mmQ3mwSZYFTUCa3RjOvCV8SOkFu2+Zg
bS1wi3cZXxNBT3S53bUJ0qXw9ATzYgiAM6e+Zi51R6U0lv7NuxfS0b6CLbE28oYPj87uwml2snfA
EaFqOeFzrFLleOuIYCQDA4CjVPr9VqGWPVErsJwplO8LZgvfGV9gZZ5LQAXlIgEk42YcVztNpq9n
1iO1pbwgygHqKYDg//X8GDpVkuT3WM2/Lm2oR3nqC7EKS8iwHttSyqTRKhhzAx8NBnF7P31GZ9sL
zYPsV63HX1MlCUc66IwbqsjT93YdZ/icskcBk1WEmEMv67qHecV2EALauwcdgDBtzXQWJaD19TpU
0Em0vhH9y5DNQ/0y8X9tKm/npONiIvE1uTZyylWhwQU1Fe6rCJvrvC/GwO55fMX2WWWuB8GcPLlD
bEcpqbXW0Rnyp5v2s7RgOGIxOK2wwi7yLK5f5VUSVs7PaGioW3ulUD1qYbY2LIJ4XdEK5mzL128g
3uwwuXVz2WiNjMEQsqO+I0dDmhZ5O4DNKeYN9CorVDqDCY1nY80/nGSSLx8iuFjfiBSPA9b68fWe
X/mbXbHm+zYpbRUg2Sqs627ubKAqAXzXuxQuAeX2MEVsTTBW4NDWt43uVM/sAOPpb3FEfy+Zb4pA
bTS5UBkIKr9knhHFzvT1MhexhMawKqD7D2liHLFGd5oUrVfhegjRbF1JLXmwIxJ0/biDa2EihE1Z
0JfR4o9yVvsZQPYBNG0a+zXDM/iZLtDZBkwbb29FXYUIVnI1Ytcmzta+S3YmbaZiSO+rjPTa7mLe
SSiianlTDBtDiyI0LkLoXwO0SkSOnUK/G0hjr/+IdybFeKs0lHvn9h+AtZtcQ8T4yUgMK0Rr8uBA
2w/TusTBD1BDzA/8bJzHig+EwhS+YMOiEI6GomMrLD03NxRS8hGI+SkZS5woKyYy7eEGKjteOz7i
z7MdbE56sAnUI44y6EBCipIn43RmbQuz/Xn8sNG4ZgSukJU3Dmuzgazwrud30Z9KHSCIHNjyvJiO
EGvMuqu/WBH2eDyXxFZrDsGTlI3osTYDUZSNU2bnJ3XT8MNpbfYAJkCx9/cY/5ybHa4sjCvGqISQ
WHOuFCHvhet0wCXwfA1k44laidDdYePW7oEc021WPjkCfwOgzwb30AeNW9Hqgby/RHLGR3tYGft4
3nc4bp2AI8i/ifJgsY/hZGqRi4mqTkyZtp2FNpKjbethR9AqL0imPbJrO1CJYZB+c1YMg1+3tAfH
O6tiHL+CmcJryRdths0aY+7u0Bem4W4xDM5a0wjWCqQNfsff2iKJrpissA+mUMffQlAzW12qG+ci
6fPhcbs0E/oIlIR1X/C8Dlh925IfNkaHM9lhxRj0UibY7o5zDZyz789NbV8upOzg9fZNaLHtKvuu
5anfzxB+o/tQVRZUnfr+vV8B0UFKhOqV445Vq+DNz+bP9h9YslC3/hUO0f/pcmVCrjZ4K4yjykc2
VruY/NJ2Hm4ymln6PRyDZM8aH3gPod2qYSbG5ayVctPhVbCv8NSBGUH+6HbLApy0lGJ45FZ2poSh
ODMNRW9wGTxA3ViCD39urXFIy/9liLSSutodFxC+LuXW77nnMLXePFT4p3A6TOwFpttm0UEIW9VG
nxhvvFyZr4gLWSZMWUO9AK6dMJ4XFv7SFc0gyQQrkMSy2vwaHHW/tndJ22jXAxCCFzG+lcAetpn0
Gs7FeTlnqA1psS10VUJkDaKcX+L5mTzOX+mp5w0qwH5Phpt0+gxFsmIPCWoAbtaDufPGaQLA7L8e
JCQpT+o1xjMInfuCXnovhmT6FDlAqs4WMvkzQ3XTyvdMmSXVs+3iL8RcDNzHlTSpUFNCSJoeSoXS
gBPQay2os6zopKiwWuW99YB88JSUAoQmuaBit6v3O6DbATw+62ucY3VfoW4Rmkl1fUgzK30eNmHa
nQjTyGxylr1U1GNr4NU+RzsUHqGOpaEqerfz4g+OwRMFU8luLBWnpVFJ97XrJgYFP1UnMg6QwLRm
avdLViwnN0DRZLz7UDE2OsArLHp4TqSrNTONWjK+dCDB0UrswlGHX25ZjEc4hRrqkv0iUh87SFVE
K0YaxsqkAEDI56qOn97o86sT1IaZOwUc9hZyA1gG+N/Y/KNEM25Ii6pFrmIfhToPqd9vfVFN5OEJ
p9NJYgE09rCuDmVIiHqLVGOvFYUMDWwf/l32S4sDVuiduqJkZjmB1dtzZ+cCfcyuFkIhQWtuRKeP
PXJs9lUwaQSXpEiwGO2qV/Tnf+r7wht+OWqoOFQ+tA6a03mAABapoxvvAEz8aZk7xhzwLULajoCo
0LvMdF2+9c2vi+LrZPTR1fLMVJTnFJ9c7t/i2Ohq9Ua20pdaI65NAPTvkD6u56JvbLoZdxiYczdZ
ReHtblQfvwzfeLT/l+oFPLWELQvJbEYAQ9wnGd+/gOyVINBwcIG76ZKqZ5sft/3SUcaUbn8HYC6O
ygRPajVrDM0DaBXWEyw2DT/v6nC4aBirfwCtRq2LnICHpRiqmP0bCwnE+kc6mW05AU/a8EpAebsJ
0qPjvEpWf+qqZ4Wbx6eTZyRfJ1hKTZCcljt4uVElhrBq1PyF/n6KAb0DzqNpxh46giamG2roYuCT
FcfTWcvyKmaK0ZEEVJp487+TdE5KTOgPmxthRtQJKEfh6ZvtRUkNQvuFjKBQvPe3BqXKgOigbFfd
dgLfTGNqx4qvmhLef4r3dMaE+4Ra0MPIlQ6mkvOK5TCsUzBN/8i8wQQw2t5rEUbSgFfXORMU1iVw
Hen8DgxG6V42wqdNLGNFreQqM1PqyHI+FAyshQ0Bshh5ymeTWybEB1ek23Hr8krtx9J9MPE31MUy
e6nL9CaH+0UkCwi5EL/r2OjrQyGWHHS+c8DD5EObYnkn0xJuekDlhV4ViDULgcwr542x6pJEQaPE
g3AnrqqindQ8d/BQDeH3e5V8CbKgUwLl2A8uVubev7kcrbuIbeZn2UC2GPWxPgolYH+60ejnbjbS
JJs1oMjoGgez8elsbjjwKY0YW+GCmKNPc4m0nDtUx7BrhX+iXf1bzlK+JHkBYGqc3e+b9EMpn0LD
e4EC/bgPb1yJu+BDXTPXhHapodmBG0repmgm1cKFcrpod5jvNctbOV0X0c6YKJp/H/EVrn/jhu3L
24wjGOTbsupsdxlzPVoSB+kfFThMRWzvZWxkeXLuFInrSCpKssSx+gXA22d9Y/khMqk2oa1jLmkR
yDkk2XbDy/pbLUhAMQP4ugPqqj0UBYu2s9Xi7tqDLQ87nYvX7ekLM2ZVEbim8gDlyun6jzEmb2qv
Y39xsW3KQpp2TUutzVwNvBawwAjKL4mTrpvm1gF8I36IZj6lj355MxSd3WQ2AIHS4g83GPJzSRCi
LSoXmVddMcJphztcnjV0TqMZ/kPxnO5oQ8Guy9t9Dgpbb1nBG6LZ7j37EBWqzXo4sGIju8muBU99
0Q4zgk4/toqdnH6vNQPe2WHmMv6aJLhOPbLYV/zkk+NYbREHD8DEU0bu7SUD2vbmoenM1r1YPyJC
tfhljMLc13rO9k+49lz/Qj2GtyXC9AVFbznHhY3ZISwb/AEqj+VH9PfV4a1527HC05w/SclkOOjQ
uq4sWsNrxbqXzqoL3rXTed+bT1JMMiICe24kD8QqPjdoSYe/6w9SuvxwxE/2GHTLpefYu/o8e+yk
HCTE/O9vj1ZZcaDQM7Zn6QYSYRFpDLO5PM8KT+9q8gjfy6MoeTHcRuXoyfzOFhiVjsxoGXVEHPa5
52qmNBo6Aqmdg/DO78U8iKZqN+WNL+shZkis6JNXXcHMDs2w5PB4xukxzQtMhFRd/T0egcwwIdTI
jQe6fU/c1ks0ELbQZlJxmd19VxrWbDN7U4zIcMuDA1VHk2sx6PJ4u/ZyxOFcpeyPUIb7mZupo47s
QPnR3mYPc68rDHCvkXP0s3Wuydi3mSNx1kqyGCKxfsY9NY+GLwRZfUtoYKecnYxC+lF7EYWD4JMR
iFPWgby0SGpaAr1unt58IMMz9ew8y9xIyjHbfgS/H7oArDDHC6yO/Wzk4AmZvUfFrcbPsGib7aI8
a1ONrG8KJRBgPV5iCsZcwV3EclXeXDn3HgJtAnbna6vuW0/B+IobypUNx7W+9yifAeTXX4xFMPoT
guSQzkiwQ6N2m8uO5esQ2bgYNO/cLq8JMwqe7ep7tXyzH9gcI3oMTAQ+lD9ptjZjxritJ0LvuqQK
Eiy8itHZ/WxUFJbLz1YBeGFTT/IO6KDc3coo//k+FZZy5pI2uSLO5c0vZ//n5GQYDl9r8fTi8bhX
xgXM0xlhR6z6eBqLaT7VHI0FcW4ukrOUlJzrx8pvz7o10gqV56mXUsCEde4YrU5zpM4S20hcsPVG
k+WGmi+cjEhb1aJ2EQH1wSZ3oKZSWdQfn+t1dx1En/+tm8aycgx6d8dlfHcZzxFp7MTx4xpav9wz
73WRMe+txow8HkE2V3ANLko0QFMNQY7UEwSdkGrawRIPorHCEZHkrEX4P/xpVfaWXjPhrapAJUFE
+ZvvKpOl5V5McM4eg7+5gXEJBcX3x5506hW1M/0WGGYG500yCoHD5YaNfK7tbLE+rMbI0vHAA3nt
PZi9PzmEEWYQSqTTvuvg/f7kLh+igKHgqMM7/nDVBOnXjhFA+r2vJCug5cugFIkNIeLTrPZXVZlS
QUJtfph2kKX2VjP033CgUFPb8QsA3Tfs3GtDIaReahq3qBJzzk2ur20KAiz4IiA+7oPaxOta/44Z
gh6mBJsJGLKj0E2q+Nx7NwvT+7GBlim4u5ogg+67FlXW8dQfx06vbgXpjI9mtN0yGB0XJXPzSioG
YDVCoB4AuS94bG/606MtLFpHe4RXNY6aG6j8GuN4xAL3Lm+eRUM/bujnokUd6R0xxl7OSAv3rPHa
CNYmG6ZA+rIT/BdbDlGppm1yREyuY8bE8aKGvh2Mg/ub1AQxdnEYZ/DkoWtF9Cp+AJi4Ucot7DOf
ud8Y+aR4jFUwpfkLLcBRAYwBgOzX+0rTLvid2mM+xJZIj29oUXXzDfwe7B7HSHvQoNyPWVDEur8V
ddekJSKeZVPT3ZVyuZo8Abot6L/BRi3vvuG5luI05w3dJsu8Yeay6OLDjcXVsEJYsIJg6RSCR2vy
ZyJ7AVP2Xu/FpdLCIJsmEXAvvqlu+AwP6NekUj+oZdCWEJbd3ntcQfpo6vmEwDd5RmdhkqFQYyqX
ZyZLReciDWZ0KYSchXwJCC8VPkRwwToQMmeDW6qDLS0k90Q+4wwMm0pgRii51SnMQtCI5bUG/hVi
ZOjkiZjr7uPCbDnv9d9gGkRynz55ScwmR+EueZEmefzfFbX+Ku+PqBXap8Bdvp66oi7MzgtKI0SB
rIeSaOygNFDMTT49XuSw/+qEhDbDTk6DTEYZ5GC4bWmc+NITR4GFakqdn62V4SgDUMPehXDU+i9o
54O77VkDtn2ex8NyGjeMlhLSddE8heneGmycmoU/QM86g2kX8ao7NsmMIVUgAxvojCVP+YT7c2Rq
GeXsoVX7K1NiJbpCmgcRdCwTL/uxRC8bjZpuPz1geOsCQI1OGp1JfBE4FoOCdEDASut8CVXFQzMc
sQGcb9eFluNtoB/+kAeXy79wYOtaBW+Dt73scqeC2szaTVhSISoqa1Jdjz4EDGecL8h8IU4q8c+o
47IQnaE+4coeMKRL2V1AdzjarZWvV7hP8aZQKz41jwxehHG5U13Sa3QJmnw/VTR2fQLuDF3uOdlz
sPYaa93DAJWZBUdJoptMeduvF+7ZJMFEZHOwJbkTEfi0Tot+QQaKbxbpPsFw+vfwwrJ/0yjRrqJI
LadfYUHcUN0eP2ZOjkqb0kXCRUaVrlDfoHg/p2tVuapvhvoP60hDgAk/Ca3AzawLL6RwBZPFynNr
8w0+lpMLL/dWcS1fkCCfGTdw3NgjfKA5eS7BXen5WZRQB3mUyNZhBYCrcOns8UkYLHWvz3ZAd+dK
nZz3AhqQU6u8Dd9be5XxhFLo12Y+7lcePdEMa7OCL99DVR9CGtFSfO0Kukod/1ly7zp1lmTHfrSS
Upk/hfbuyFWmC6Fg4Og/ZeXql5iprrk/yLl93QAbX0ENe+4Mlkixc33nyweT7Q0YbdeU0fcvIsCG
9E0MHCGFDFl559/cDQhKhv6rn9b2w4rBimVJpyYYSIGGgJCrcMfwkwnTvfV4RnwoXZodmwc82Y9e
Aux8N6s1Cp4UsGyk4OseACML9Dwqjge/ujpsNmO+QAMisr7MGEhCiVP2TBW9zDjglC/9lCujUXdW
SJ32r6avHu7f5uMNMqfK339kTvE7TD9LLNthICpEpnFGeQNB7gRTJSmB4e/goqZ+5c9YDY3i+o/W
BTABCEAZe2UeI9JUwbYp7OxQNo3wm4ZAhviKuV/68nOMStkpgaDbhy5AHD4JtI/BuJyJJoz8iObH
YI2n0KSsMiQyR5RPjG0F7RHfLOZKTR30gXCcpzrIy+8AYCgJtYy/6GXVf+fvaW9X2W1LRGdIJKmU
tTuK8+nKK1kkOpGTSVnLC1qb3qvoLcu3mguTkzKCMn/tbZnxqrSajdSBZ3aLzMqfmo34jNQ3KBt2
K9EC4LhflrBcz6HcIVc99ttljAJKpaJQ6iSW2rDFDns2Vf5qwrid4JHVXtI3t0WY988vWdy5uZpx
flCIGeQPZd+NOcsAmL6SnzSd/2fRNuyFF8j2VimylYHsUJbjpGIyamaz7uu8HD8V5mAf7hDUgGkc
EcUISWThiGn9/gmM9ThMY883+62/ScPlQw6sSgSzC0opRq2yVE3cP+5dyY2PVg8kxUO3QYO52E+l
kbaRAXndwFIbH2/1Y7kScrp7oXicWkdwu01UgvQ011F2/mOEfTRu2i4n4XRawLya7dCumz9ftk6p
f02l2kgU8mUix5mM3cQ89OQcvvRiLx6hGc63+weufjg955cP0+R7NpLfsj9VHuRUj/2q7aU/zumK
n4gfQk5zLrrpaO6mJ92LJSSc8Euhkf9PzMtq36uGbGNEQyzJDbZjkbA3jFLciAah1j2tu1lOZ3vP
/AdzktkRVSV+9FbjNmHw0WfTUfoslil+3FodGttBxHygMOuqK9yMyXvoKDqITCr0xJsJcnLua3UW
VsPDVQc+dTM78TEyGf9QJ49XjuYGBuMjqCMyJnwirkdb4qppse1ag53EYYgTKWIR+EPepaYhZ2JZ
N4Xb4iT0k1YoxB/du8twPVykzq0sCwKl89VLKv7qbzQn1lgglxJRLvTrTWzJNFP5PdI+/IgLoCns
x4IMlOHMFbb6UfVq11wBQEK85QBajGQTX5dBjJbksAzvOQJKJVPZfDhOMDCfE1b+QUlYaeU9nss4
S1RSm9VJT8ylUAxa+WHDvHXb0AbwQZhkfd3Mqv1z9NIkb06gCYWxva7lYkvWv48aeO2nJISPaGGb
DHo8w+RoEdxWhefDq5mQq4UDg20g/zp9lQGD3FwKrC9s9Wa+F1x8/qqizulHaSYSPsG5K/mp7QDG
TwKim66dgYI4JXINwc2HYLO/VxNVjNFbtbXlZpqpNtortQRw9i7QLvPvB0tEbtNQ6nIJ7HLkXekM
TCTkKpjlxr9LxMgmXQm5x692Rh+XUeU8qAQDADY8QgMFkaiTpxDC+HUe/43oWfh7b1kyrpLkRs7k
gTWlFxb/kYxSLd7LCfVVLTJl3BamFKkB5gNRWQ/ffxLzy6EmABP8hW50T9x9O2ELXByiOeBvo1RU
r4vWI/2b3zsopWAehpT85TdRExKyJ2AVGS7v1gnNt/Qv83Kbk6KHDhxQ2Z0dMUQhQ6ck4BIcxn1a
UgNHS2hthJ/Q+27QDLfpJXpYqpPLE5+a+0OrebNFF/KD371YMJc3GPwVlUF+/qT3XarXt1tBK0ct
LA79aarkS3GC78xCcjJJrwSF09Tx7R5YkyNj5y7nMhO3RAUBa/JQyI1B1p4T0dehFFSXGno4nqdv
vMyjxOcF6tgTeYdceSVRLBDhP9YTat8KNyusDRPsQ7Q8RImsQgl59D3K6pzDUmdF53aASueBLALl
ISjyLuI+oSb+MlYv202b9GQ3PMgnStM5fbI5/PGdh5e19kNYgkGcvKwrH/zRRtGylu4JGWZe4NRf
rgvZiBPRrsrPR9cpRn+CciIbDIpJDREJbAEyHotOxYxQ7L5yLjL4xLda78S1f2TTazab5JQL0Jac
u+A8VwvdzN9qr/UQQVshHw3JJyt4A8Ld0j8LZsLdA262FS2+sIH7uUCfX8MGxW05sJr8tPU1DVBi
WuHTvIJSCtGXP199EVWSzCfEBk2zLmUKZcZ0KRfRWVebhynxMXyXrQRt7I9vlj7LqUAUAJsh3IIE
cd677zJVRSWjzowOeQVm4vIAcXapxzDq9HaFMYnRLXij1QRSecPfWL4QkY3dss1259VcAtQ40nBd
PSXzE1BdL+IzqEwbCymQ6+SNHIfzIsNiyvEEDW/qtOA8bpBDIK6z2tC0AgCc6dKb3hYQJZ8J9Z27
Kz/K5Rtg4/G2o0KUAHOWudC4QAKMZHAOoL2/RqT4pi77le1ewzSBLMsiCaEL/nrwfozDgrjX/rq9
x6ZsDcbcnR3SJ94ZharMQvrqoFHK73wO7kSFxJtYaNMAD/xBTq4Sh//lV85Bm23FJVn0jiQqCr8f
Qyx2JSPxbtiV61BJiMdE4YIZjmy1zwZzu4pb7sCwRk5BLrU3uTrs0R7iAOnCmvPiEoO7sCmA7iuB
AKXVrSZFedIlne7/VMmZoA/f26xYE9RIuNUcY7/eDqEnDTrpN7qliybjhW6leuCYAKk1LDnquSnz
Mx7x4T+H1RSfcfj4BAEMCUYDogwIG3SMUtusqdvZYxu8FVlta9Uzt+eDmGIXz0C2F1hUVPAmb0w5
+2l/BhgjNErxdhb4U8fnLvnPlFTspcUJ1YGiZeXHgySnDy4p/mYW4peeF16V8g6+WK/YBV/JqU+q
XwjdTYBLVf0TRnUnX45DivnodeH4cQfxCDb77hGMUIWAOpaTcYvFhJKm3hjEdlHrW2ZLK9qzxEfi
GTrtG+OHeB2An+c9qAjncEoYfLrKiGYGl3Tp6AyWOBOQmLtd5oCtACp2f4NTUXCi4vl9Hs03IIBy
VC5T2nzp/2swjzzr+9SLIpfj+Dd/AgIPBu+625QBru0ZF+hY3Jj7aULUL1Wnyz1Rjz6Tt4hyN0CK
cWskG5Ub8Ob3LGulkvlnFJ2/L/uBJQobArjbF5xlParfQx0gQODSE+d9PDnK7HxaPXmIHK+bsgfV
LtmwAC7bLqHC4/t0LVrzzyc1BPV1Bl75rKHFVDCFCBwcoiDrNc6ZcrYRsewkgTQqzs/+UgPJgncD
oGTAIcVlc6vnSgAyPafbp3bmhQ/dQ3OlyT15BRITJhtkxUugg96TkK8jYEK7t8Vydp8SWwb4h+TW
63qbLqwOBy/8ih8K8ASqB9UFF4TqOIhsPatqWm+u8LvyW0PGtAGskCG5WKddadnUPfrtjPKulyZw
2uATNXGk3rJMIrkpxLWyeQEKj0P7oHhEXin7CPuupj+Ps8NAz+f+b3xn6rKrYsJaoMMGnb9zVRHT
D8Zm4Psif+Rx7smAI30XdfVOP4aWusexDvz4gpG4wpERoVvHR1hhBvGP0oriwkKbTyDEOEj6uKTO
X8MV0dF2P0LNAB5wPcWhFmiGWzlNdCgz+0CTcHIZhVS795YKTVZXTc0g2XE0K+ilOvisjiiSslYV
2Gkl201jHevYHC/GJFtl2GI6zLeT2ggM2oza0NMxxCNHpJaD5braZ+wk4GLIXFBLotqedw8N3pPq
zqL1/NryHfC9cLJGcvl15OIaxUKbAbeGqY1nUv9xXgAECHI5oBqjeSAMytbOJxRW/G1HHuYuPBq6
XXm5OH2YSoOFMJI2RMfgYuHwz+jD9haHlXTPOg6aV6rBhgTm9IvFnfLG9A3Idi04t7JtGrDGBhi4
Dcb6QRhidzNdroV3aPFCaKcpct8dhLkn0ToWNGYvgj0UHPKHuiatZacbAw4IJ6geuxyOcNiku/0y
OmjUo4rHmmYcV7JzP6mcSO5WazWosESvd1KIIbfNg0fhUD3B2yIiLJ4UxlDVPwXkCXXUmHiniCmp
BQS545ujb7c6ZJe2FlFlJcAellYHd+jvIluMWQCC4rQXZ6v2NpgyYzyxMYlE7trI9BKwkkEgP4G7
Z9vpUAe4eTAhLt5kKMvRdzNs+NVk0x9Etz8NTU3qCXHUAdaazqpG5fEDAubc6jSoushzPSk0WEM7
2RS2FG4o80T+PN3XeQrRpMicNMoN52bmo5PkOE2yPED3sCwkbGDU51Xmk1oLcR01WCX7WMm1m54X
SMiiMVf5IZDFrJhbY3xruYjOz/YVpPvzbt9bI+O0t2K+9J6UWm5eG64xdWf70GWSCGjYEIqUUSz+
D2yn+/CaMN4k/MnG+TzxdHU2sVAQO37CJ0zf0Hxn0ClirLbP8EjBim8af4Jkv0ydLmafLMBtqUe2
FJiVkdbai7x4arFpxt0ykkETOU1XEgH2QuCv9BgzQtSSSocmXmcW25R8K0kpiXF9D6hVSnpOSERy
gQ3lMwdto21HIj35OOI7RpNEGWK4NShJfrzbAyn+rebZVqEG8KQMTGhcxJuT47VD//s+HTErV65s
V6kN+oh6r9BLsSq6gKxJrHwUnOwG3y3jGjqyTgS9dfcrFM1DtjFnPdtlqX8ShDJ/CN1B/jLfEK0u
T4gpVyLfuRRp2a3lplyhIxaOk8tA76IJdkfThxaVjU+u6ydDIKJIr7/i9f+F9LvPdLtbvM77gAs5
MAOyKJPKR0DJ0f8IXGMb0yunWkPSQFHHJxACBqusQcNLeiFqPqO4LaECVX1FzIFFrrhKP90CFRWc
WIosVGdvS/RrsxYH2367FWNb7+0+dUPw4BEttSWNR9FDi8MG8kI3VT9JocNq32BpWDD0iQ5BSluZ
qAh27xwffXLnFshordv/TTst97UH042JOnAoYxXDN8K6t77JlkxNJPaGrzEcOjABov3wNQBP4tAd
hF61A8RVfGDMNWMlR0kX+PHgjrZrsozTKWYcGjLQ+Frbwpb7CW7WLylyKJtDMLijlzQ9TNbRC/tg
nMoJZIaiMM7IIImGgwWNypd7z5w7oHQFudbWIpB/dZlF2pHBD7p/m8qX3jC44N2dmynrmY9wVYLT
tPpZ/UBIM7wuTSvcWGY1B+yVkPkuv1Qd+ocIyYsFnriHIkgJKoJMPzRWfzO628HorYq0+e5JwN+Q
GbQ30TqIfATOtx2lPDlkwQqEmh3pkLVzqT3gsyeBTqgvMzwgDebNF35AS0S6iw9vixGhjHLtzIah
SEEmtlDoPdIFy61hPLHUgWlUuyCcW/y/N8+bnx0R9em0l92u46CYVA9pjEmCB/a3dhyyQO7kUhbH
btomD41MupnoozHIWgarhObs2Iwi3iAESlqPeDvlQ/v4DtJiEDBMvWPOBlL/l5Cvxpa160GiCVNG
lpYAMqMh/UPQuHLSQH15SFfbcrfDnAe4Z2BHBCELEnP7axY9Ox+8lKpcJcWLAFbZgb66f7rsqsRr
nIfYwBuu2rA4yzV6VlcsfuBZPKuRBjUwdh89zwQyCkD707ti6Ldp8F7z2mSHla0A4GDloJNxQ4qs
vglA35Ifso2tyXpjAU7KgWdWg+np3Fgnlc3QKepJZxec9vSyPpdahNiRBHqdmMdj03m4xu4H+ODK
UUSHbed6R1nmcRjsjcJNVYv04Xg6O5u30rREZa9sxjem/OQTkTxXMCSlY2GRoo4IiswPRUU0eDh4
M+MKVy7jewL0ra3/5sr9t0N3O5DjMuwwM6TfppGgr01J/m/5cyPmDMr+bVDRBmDTaAQsjIH5MlpB
eImkMNaOs7Y7fIgKMMNO8+SoC5Wl+fjwx4Bta8pI2TuyUsO10EjDpYAUdj5FV79u4eLH53XdBwwV
3pMjjtFdQ++KZjpILVRF1jWpZ01MW74XmEfF6uHsyl7v9KKWPzN+Fahve4I9vB4h7Sdvf5h1z6GX
n86Mk61bVyYzMC7W4yhaEQoHV9tQwWR+fD69FKLB/eUr+MypdMPCJeoSnlZFJ+9VvTTDNeVTsLnU
pf4yMu9acAaSE2CEJU8geLpmotAQ9OUm+DYnnZP/12gkIegsj4MPkdTBUcVS1p3cDUqQB9sFwqkh
IFyKj1Cy7fqOcJ1W75fYfmnRbkFKjo/cblfGyqMi21tJK7i48K1QlL9baKCiBpjCyu5S7PmGVJ6v
Nlzy+qn0yKECalQXHI/xXoIlU7hZtWapligBqsIs3/81SChJLdnVvwH5aIoAyQK+kF0GuDq5LbSM
RaKCdHFmcxoNrr/AYCqmFZyxA0EadIt6/VuU89wdZklG55urC4gppyRe9pIPRpiT90V+FTV1alUZ
Hq/EUAEnHBdAt1GB3gqL/30XilpFUwkbOV+GmrxgSzUwCgQJFAllS3coujygMqGHuxQ8BrjP/0af
rFyvaLkjZ1ikmEU0st4l8Dp90GqiopLMT5pFJelD/gxOHmVvgEVjsKghhMAAULS1J8SU+tc1NkQ+
fzQKOOGA+JRxs1/Jp0k5PDPQYy10YHDCdnh4qrj2sst+79XCJXw4byUq7Gb2EHcVoguT4vhlUtfc
ggq3Bm6NsXevme1tfRsumr9Qxo/oC5LGw59jPdro9LtW2pE6XF8jaSnDFWjjoXyMoDMmPl1EYDF6
PggJTIDWvA5TYU1DwwHdI+ozY8y9+3OnyMaBIwRmGeCpRZ/GHhvy7al5+/E805SCYZUgiG5C4LDm
uxt6/M0AM2mP1CaMA+RceDRRVBT4XrvRxVDGZsx1n368qIsZrJ9+7iPd4h2tBh+nSrJX5Zh02t0c
xtlJ4yzxxtTHVlRrSh1uXtXsnSR0aPcro41w480WiPghtRmW2Sut5H8qJxyMDB/0nsfmNNF7IEXi
GX3ISKWb0j3k+QWPumP0yrYzHCFj6xZLOA14JofEoJPp+ahR9MiMaFhAWqXC43edaftL3yz1iEbj
3Zo2d16bLIoOCo6FlT3S/D+IaGvD3qwCwc4uqn4+GI/QQ3xehQaInr4fpfTIHnwr1U4D5/mkqAD1
u4A4O5LxQY12O2tmC9V/ToCOz2yVHVFBJbT5IFCep05QHGrQYqS8VwUjSLvqf35r137O2Ba+XfUs
Vtoe9QjkpcpMNXAenq9JJffc2pivSK+EyRnat+R3zkjJ5TrXcjMT9bKsLG2LlVq56vLIYFPhD3Kb
SHn2omadmS4ZKdztXu5d3CoEXrHsfjP9AGj01RRZiHLl72GNPBNTrq5OiRkeTYeGATJt0s1y6fp8
qRc2wrZweYCoNPmXt3x1RzVekPJZHwpLwsdGpgORQ0dUJMiRWzueUwKnsIYG/up74RzZQKy4npBu
GzzV7Lr+0US1WGnos7AqMqgDjonhpgmBPzzcqGmD87ZgDGGVjHsPFGaUeDYQjvmCER1oi7Sg+ILX
NByeHutlq3uwO83pZO9yRRrBvwaN1r/c90DLPB+kVJwRUNYWE2pDptzFEqzSosPa1WoqvaJDzo1K
3qQOVqtSuxHUol4+7CbM6xqmoy73NNP5ifyKshm5hEXVYBTY2LHqwV7/CoYvZD1tMiLDat1DLzAM
3CcryJzlIIskMWba/f1ffnEvxkJBrImYNSqljtr4oUGFLYaTSK37bwdBxAo7d0WXWfYRqcvtd6PD
yW2yFuUOJ6wjajpvt8X0/sqcA1wHr1/0wl1tRkIvam30zxKnL1WvgVVhllBoRfdWWj6wZs7PvJzZ
3FLeVh93sO1D4BuZntCySC/fqKM2OgYa2Kr2c4q3q8RIbb1tMLhKgJkqAjKWX//Dz4mWdr1l+Dph
ElHrLp8+RTuywoBhy2vN1+sGtvk9mBdO8B/Q0L9+zoFBnlkWLk+UOQul0zPUARYYFBRDywJVv9Mq
UVSMQzE0yazWzOZCC6F7Eiu+xBXD+K6s5fw6PGSC7NMIfo00SglNStTuwL2zBq1nNbFJtKgysQF4
9e3flYLyBRQywn8XOg3C2oMCy/EkcyjFpUpBfkXU062c87U/gHthnktidfKSbNmxHtBmUyCdNC4Z
OQnq+gme8vMbLZzDB8eE2G7nha9lQiX5cffaDQ00BIgyfPNr6Gs0q+iP5Yrm8ToYkSv650tgnYvA
m2cWaq7u0vXbVrlvoirqP0CCXK3At656frmQgZXG9yvt/qaViEZv7I4TQ3rv+U/SWD/VGYXiLYWd
Yqn0bmsLyQ97z2R9mecdAB/2u2JjARA3v9OKMERYVkWE5Wts91AlY1OuGiyZvh1NO76OqtRkQevh
aZhxHm7S6PS1z05ll9LjYFc54JUV/X71vNFrkXzecD0kpQYWeay4/085Sq2tZW5KSRpAe8mRU1ql
e/9WkKmXq+M6iDwj67EKz4UKNsSASmhvYFgkuyC+ENGPGo2H0/0Pe+v6LKLRf/xCmQOXM3Pms7p4
srmUiLJ0x7gVJ+PaJ3ivvBLhWklLXOGULAj5O4XiM6FmL6k/WpJdnL5RA3VPzdxDdjqKTDxoZPy6
WKT7iNIDezIRxp66dn9DFvihNfm2O7vSM+SYOHjTiHrIe9OIbpvneuEVw0UFyT74lBHmPGteudLT
9SN+dMQAkFgBlmKTvseJayuqXqKYV/DpaGyZYsLRZz3MDLfaVz6IN7+XvTzQPi5L7l2RykhoGRmG
Kh59Hjs3qfQ343pYC1sxrji3Y/8dh9VZf/+bMT3VrR/06NldUxoVBYTZJt8zJ24K8+WlBksQWCuE
xWeC1ay4CxXgt6YYRKp2hFUmuaRIaCsJYKF70XgFc4rDO3kgnp1gmongykDkqSKSVK3glATuOhRS
peNaxlbS92uuVowSQGOX0HTm4TYFmxS7mPAc9JHs96v9O26N4sO5qgPetjb+SIISTemSB9m1HPlD
vTMaVZbZzuNxB9WH3q7I8zUvPh6YtrkdZtuYlQPwJcnRd6p4YOaHtuLlxwsNq1jQedtxzb8rWsse
9Ab9o7GHyVYLb+7xPuevrEwEdPFYo8fyPzwQBdHzD6Vlc5zWfVskaP2zshZ/ciI0Ieq6RJDeDRHw
CC52htuAy5RU3PtJkrf4v7ZGgp1aRCJGN8p1PEzrcigDlnqEnPEk0565bU8IVcFP3tGw472sPInM
zvkNtwTcgO5HnqOR6Ojmjn52FXmscep7ukKfhJvLnxEg6tyYAPb1InCP6A88tFe7d64+tt+9gjXD
aSfYwq7oSkOM0vfcK/FcJXkvmEzQvDWtUldXBtOHEHIaVVaXJl4tjcDvPWUCSeRO1s9jnCBiOtzg
Q1QeBqZCJsvEKH2ElrsO9Dc8beGuF7JEB6u44YAxIgi6mWXtcwrQtnWNqilpmx/dyARxPmqRi8+F
Oy4CZp8nTvoC8p5f334WsV97ayqIPwCIFemIuWCWEHjbwUEZV74tzKmhZF2ATPJ1xMV1NkHD+zAj
H8aB32ajy8fC1djxmDd96iAI9xHrgvs+yb95/0xJcU3Y+qvQxRMGOhVUIzQuY9Rrv9moLtxJNAld
sFu8TaTtLrgtiebyywSxMPAm/xftosPjuFwEJ7T2+j7hsCij/749ixGMvUAM4cK4sLChhRgPgj4t
zPd5yvEPf0/xdrh2meF2AcSR4V19B3PB1XNX9HRVsiYJbOZS2hBkjUi1GNrRfq5tHH/w1MmBz3b8
4VfnHd/A/BkKghI1ItlEZRFiWvH96IaAFunZjrzCa3x3NL66HWUOGc4V0Sc2SY7pfBOpmivKTOVg
YehjwhmIgrOa8pY2jKe/XlUvo5pBcoEEdu+Kor9mEUMu89EUeLUfhQQkr5a48m/0pQ0EFRAtLG2o
6GxnBttxltZ/5u7TeQtnz8vrCQLK+6+e9u8aUd6I62vFusIFnyIRVgfbrdK6Q8NNenmRtPrimz72
tvAp8dvdFZRHUxtdsAVwAeM7CzH7zmS9rW/GW6QdPflwGL1Fpk9axUoByX3fYAE/q2qtiV7LILTF
US6Ycojof/m1mFi5cmXON3zuiPYnyWmHtNwpqlA5tRqx50yNSLicSX1Qs2AWIZ7Gi7s5Mh5SEBH6
CCyc1FnFhQMk/Vpp5SI2EU7vOEbIPFaNjOfiY7zRqzcL67XxE3KIFKn1rHpJtrAiPblOJJCObl4j
v1Dw90skbiKm0yRuTafH+ww7RSFJsZfwwYLPn1PtQokesGUFetWdj/feNEjTgmSzSIeITVeDa/4t
Gu+5fqn0OfEfnzY+ZFqSqBUXSxMvUpXY59dKYSGy8C015ZyS5OpIUxmKKnPCqjvB3ZrkLby+9FWU
73kxbfyp/tqWwESdFey/CAQzIhHNTlgrHYt2T/BekPjCeb3284NaPX+yeefJYsgUfEsq/1Dh56q5
T7AiCbFypXY/Y11o6H5kRahOh3ojwOac1LCvaK0HzhFSeiWlFIzpi6ejx1p4CAooORVtCxWtMHLf
locLmYlZsOTvbKGauLI1SyUBf6rZr7Q9uFB+uK/RABkpj6EBydMrOYQrDUIastHGxm3gRnJl6ISs
Wack3Bbzxbsbc8WklUTTuwzb32mGzDDXM4cKIoQitzLVlzg5CgttROuwHItroMePhvDeLPrbh8A0
HMZiqPx7ztH3jJLJ2ClcDFw4MldehOYLBUAnTqSVzM1l+fBHGCgvMc0bMjyzBtgNW5aZT0Xi8yT/
f76BVc4ps8YUKe2XphEaZD15Cr6MahVc6hRAPL8oC/i1RE5RWKcjp+sBWZUI1JZyUvw7boo5L1bW
+zaB1MyRpu/QqxIqkIfgeb82dddEe1xhVfGAy9hdVXaguiUlXqMqJhDgftEKkrZu+zsDEYfxn95F
IACcKKKkI/fpRnSZ2wLsDTPYPyHU/sJwWvT9hjkc4WmSeVdm9wddAMSWO2ANbUxA50iUD8mdcEls
ud+/EOYQh01bdsFmqGfR84UZ5FWFawRdX9YrHHO3gzFxzwiJDlDaf3qc01de64lg6dcbI+vMYSCe
AqLaqYw8P+iVq0zYCWAWCTHjR7j8UHNuQdScQjZoyE1JTmEki4FcHXbfo/53idgC1kWVw1A89dop
ILdcF8VVvB2m2Y1iKLEKI9gpRnSktdik/Q4/Yu795PhrtL35IoBO5QZ2KXJuDabWsMY5SRXWOZy8
H9Igu3paac89lC98kRhni6o1TbV9XkD1UN0ujh9JTq1VKs5ipdEwqinap9zQ7tvGZxqLFCxvsUCx
vanlBEwET7IHKmIQX7rNAumjTRdfJ0mJI0xJc5MmvV6zJtBmxq+bZSfyW7/nO/Ac+O+qy53v6XO2
3mmMRUvavu5olXL0jbvxMqe1Tsvf+aOccoywkIFyosT0g7UivAeYwMmP5FgA9DuuMV8dVorzDQVp
34PeiE6ScHEAGXyyaFLF7YL6I2VOpTThhkGpx9TQCITxWhL2POsPPP5CQmpcGLGTEPcomOPRXHBr
0mGLliGJSwqVB+TR65U4B2QpwKlNZD+W8Vp9VIu7W7iXEfxLXYtuvONb2VqWXRhS+pYBS3/70rdP
65fizJ6F3dvy0tkr3FvsQdeU7QeLSj6hH1IZVbWB4mE7l9y+eEWS2trL+l6h95j/QR4lMcDUoxFJ
zD8KLtGapOC8Wtk8tDk/t838GZ7u3gCvXGjy6xo5iD6n/inabbyWyhRryuBTr6B5xFIfBqnjJlHi
qUdfRjaIW0Fyxfc84mDNl7IcF7BbIuBMssnFnTAbrA5fdPjY8s7EXrAII0P0e06d7rXfxy3LL06Q
Q073REZD03NTKFHF6XIjQh9+10NdN1sAQAt68zxI90fg69kAaTt51K+Fb1fHzmk70ZuuG6WxQo21
F/gNJDx9Kkqyphuembyf1P3NrnacG9lLc+ckwg3o1nVBQDZA/hlz6NZHpeybH8hKK5O/0nNED+BZ
nEDYWVgWUrKK7/55iDcW5H2SakqN+mRJ/Kd7vFj22njRlNwQrI3iuXgue1kJNhTv1slHrTYI7lt5
b7DAtrpU3G86jBQTbWcJ0ydm8+uqYliadwAkQAD7f06Rpkp/6t7rQlZV5YXBz1b3XpzgVuaFlg8K
q/3fmycDsAZmhSSoZUJsSFXD838UcpaoHR+MaXsEWut4ipdcuWjR1cE2AHqhQ7QxuCrB6NOdgXqT
2mW43/m/rnmkiMZpiSZ+IyHwB3v/lwE6TJ3Cl5IkWdMrnwHwUwPlKgcXXM57X7p3ma7ScBYsEWrf
GmV/LzNO3DZhFpcZQp+ffEWd/Ki7nkoKbpInAZQSHodQx7GGnLqxfOiQZ4fBm0fmoxPCNXkp9RSF
QUN56lQS95CABEQ0h/yY0zY2Emn1g5VF83VXsnzM1l9sarF1AGIr9qSSdekqeHTe52K0A9EhMRcy
IK89cHVheZs0NBBChhx72ZB8h1yhTvq8UIibrJc7ONiVgM6ZI9kExt+yXtEoXK4H+UPHsZdPVgH/
eNCSdxWGTJ5SFQiPArvw5Cn0VwRJiQR4BxY4ZkdNzFBEzjAv16kkQFJ5mRykLFn3nIdzjxccaFwq
yE5HtGjzqElNSYgmzqxojElftDxzArFgsXwEI7oeiz/0Yh2+rtdl5I1zixXkQA+LzLQ44K+kVwzl
3L3QtU59i+9AvqbeRU0J3p+HqXGAYrnBfYdsFNOyetd1qZNr9Hfok2/0LGXL8jeKmvI/BcDtuk7R
M2WNncdju3at9i5w+8pxb/QyeOsWczE8+X0pOdmT4BMtGJN9ppwOiz24S7A5UwBSyOmIjNTYbb7h
9ipxZyAZOAcqL2OD5apH84aj0ehc5Zs5rPX5FmL9Ruluhk3eyi4MgHYqJkjoJmAMjo6oT3vZzAxG
4lwIS5qrQ32mEhrHfPuGMveItA6JFRtRN/0BYJJGwwg75tWHdqEB9Cx6l1zOJE/Na6szi6brX34z
7Lapvqor1hC4m4F6D58qimoQLRBjp4/zhpitRTM3SsrE8h4rNb63oiYtCfqeOwYGCuK5DSRE2xVG
d23bRgrnfR6vZo9+jZT1nczsTchjMkXtlXy6KMqaJoJ4adygh6JdNA6vJL98lASUPVLKTgdPY3AY
yrpuq90PYxbYGlBaSk53CSqwwDP6dVgZTaJDSdaIde17vFIJbZwCbAzSt1bP9D61RruVSkrQ+qSc
yjJc2bGE/LcJrg68wqxAFyAemm9EGOL4wTX6JGJnYYhQKYm46L1jhHV44iOxdxPqff2KG4dNSZzD
Oz+CzdKd/lCM3fkCVZx7QrN2jLNZNKWVbUSxT5oIw4vSgBUrANHVJ15wK1ICsNjtDZxySAmfqit6
2pC7QJKIm2gBT48OGBO+V6iSHB1bOMkibd/ZAXP6Uy8TAJNTk9CxDJysDyZmFe6HUC96g79JXZg6
9dyOfhk/TGtUECzBIjCYJG3fhJTQp6kxfLWCftTmZGFjW5xfasIoLzdx9UCr2q8Q0W18s76MGX44
5rrscp8PK4qL7wCTnz4YuE12WDuZ7yDviuboRyRp42pM5lKEim28Q5pSdchaf7qtA1XmE6AvFzk8
u1ULXXM0xjRwHUCOT6uPRVcj4Fv/Farm5B0YQb0aoh1xF1po5jaT2m0hui+nFFCs1jOvnvr7w6X+
chfYTO5ZQ8ijUMhtP/uicWRNqsIN4fEy4JiRgpgyhtlDyJnnikXfbTigs/ti7YZkJBBNlCNrpbaF
S2iaLv0dDf3kIpB6vQHmZlh/udBtC5dfUpRJKDiwaFZgQ9G4sb1qn0t3R5Qi+YXIXrTxETbH5MWQ
nrhctxJ9lwoFKyCDAjmczOATzr/k/UzR7vUrVM5ChJMeUKGSGjTLPBlA1f2JjY0ngoD3i/mBqxS0
GsA4oqPsHO0A3IiMDSLfk46BtMzH15KngAiBnz/nklBUN6tsBAtQyPnKTTTaPNLImXPpVLEVCvuW
9uiBaKMqOu+/28z4euO1uSMrkN/Lyj77IpfH7PiQW5gw+Y4AGM+rnE0kTEGx6lZNKHVmEz5b25II
gzyrOw2bMQfaWoEHfttRP4f1OChsyhdcFuJq1VViQ7ye9SzIH0J0tNsxBBer8f2oo1Zr2IoOcOc2
1DDl8m8+tSZBtVjSHO3Uwo+Rp2NuwYn0eEt5Rv4AZIYEM6S9kB8EewqQP3Z5clFwhTjBlwfm2B/o
fbq2ydSQszkEgMHGJyacKQyW9avJwtQA8qWLRPaPVn+ojnsg3zz+coxr/snz9nojQst4lXtxOV4C
mUzT0xst96V0HWE3kBE0nFsxIHnr3p6mRZ/K3qi+tJZnfz8btiHOy+IYe6P/j9NGM3KFYZeWleZu
j5JYcKJHnasY8s2MhI1PRKNeQeITaADNXPhECRl66UwJZ4yNIGJ1iWL7u7hcPECNF4cJSBnTDu+U
4hKqbqhnnohzPsfHEWDHKfsNMheNQZvKCi0h9U4lkmum+rT9ter8ni6owbUW6H1vjPWfgJGdO3mz
+zZ12r7wmmaoutjm0BRygI8iA8EPDtC2xT8BtQayqZtFpWresNUQFDIg6+3YWitgedPur4PFe2zG
YY9tSH0Bar0v8sAPXrq3rjbkQbhloFQqz2iwsmv0+jKP3mb5cW2lxh9fENfr7KputwE2G3HeHuaJ
1b/0+MmKNlJb2CbMK0+pg2zw75Sj1Q0AjoH2k2Lx6op+pzCpLdRNEVVvfPEB8nLDLXWroAeadlrW
ZzbB+1Vw1GrdUpin7huQATvoInKhElmTh/IopPNGCKM0kCnqamEOSZvqExBSN2SSZfRZCtFMqzio
rr3AxIHNtOx1LrF0a3HFXNSHC9YhuitMszm+PMHTdTnkLSUTP35mXKQCNnHqesaIQ/GjxVo7m+ER
o7CdrpI+mNzbXpk+K/zBBTLk6ANXG/WY4PD/KXwzvrRENfpGk+raM6Zzkf1TRxPK0Q+5FqaR7fwC
c7yE0KQE0ZuBnS4Y+JqtTvH/E/G6KsXSjJhtaweRN4i4A9F2q8C0nVncejlZcYNUmr0DdPefOQ8b
SDar/w4hUd6TzHJ8PaHyyLzv+y9KX19T2TjeDyTgzMxjEPg/rUIxfutWsQCktyvVyx4qAFWlfleF
XziDclV87hkcjE0EbCV6VNusImaSCvaWcAf54MmwBxxckF+aGSbdFTcnd4+Yt1oUC0/3g9dOVQiQ
7f1srgQDahpjGQ4MTj6FEVVyOIb8yEXh4mw8o7t33sWC3pglK3XnsQu7+NRORCBW9wSkCjxnPAy6
ydaUmUDrrumoW0jMj1sVWIcjpmKeDH6IrHN0d3sODtXZLFHDx2qXjJrQJG86jueaij/KRKKl3Yno
yZrmQRR1SR4FMtFND+kaJEv4yZVFhFfBeDbcbPgQa4YCHKCyEW44g2E/wgvBrEJ4Dpy6btv/JbT3
DpnHsCO7MhSfLrC2FsLtU4ay7cuNi+1CmakdOB91qKy8qinFBHETLA9SZyeOqjU7/IP+ER4Yq6P0
9HT1viWUQ7hBgcDFcdRyMjP+EbSlP6mwbRgy1z2qMUSIVW/DiEX4Cwz9qPi3E3+YQi+0ptkGcBDH
rJA7tRkFy1kvnNQJgZvrJ+RQZwboVBDcIvJV5WEt1dM2jo648APjO6Xwi6YWvvOwbOQntzrdNVOo
vDDWH+22FnOE38/g9rYGkF4QpGsQsdw+hy4c7TWgGr5U1csrogwPSmp1yjK8c9/CYbYT5Xme+0Q5
XJiew9mYFauLH3Mvv0JrkKd6GBA9P7tXlTPY1nhmLlkladH/5WZ7GII/e6b+KemvvRJ1j+e+We08
LlWfGgDDhNaleFuLqyKNxo0ImIW4PQhRYKLip5y3RsxIBSoy4YLUvvszlikebFN60bYAa1/e+CQd
+LP/vVMZWjRgaw2iIyneTFSCG7EFPw+wnO8UIxYTMVro6s/Bxczaqc12ZJRbN8TUAXsQ12Xzocid
Uyc8qjf8J0HQ9eNj4sa/w9QFtqD0vMygB+msAAF5d6tFsigLsHjv7L+uGY3JELOtjePToVp4aoEX
0O8po6nMBBG1XqV6ws083yczM+L+rJuFzeIfdmkqtdV+9+2HvFvYa+0hvs9xhqxZrObWTUdvlA2P
4UvcOE/1kme/Xq4FsmAB5WzixQimGW9fpgLrAR3h0QJtdzETTeDTofnGTlpund1uoNe7QEjUjHfA
ZwzeKfMzYpqIzFIudbT5aCXE1HvW+S+QF0q6PUK/Ua3uVpML1P2Hy2411hjlhpchhHkaSuxtZG4w
9gkXZwzDKKiQSnzKmJouDEtQ0KdaQjOHPG1FFj82532/JX5s9EDm5WGeMIFgo+/4NZhYCKghAcTu
4dlQd+X4EZGhFIsKT8PdPSkDG8333U2EhHLIiQV+t9KenzSOvgNit2h0yapC4tqBmHu42kaHS82F
HJLgJzJQhCwTmW4aLgpbqjhvq9GM8/SW1gPS1v8vbBrvceYEDLHHSH9uBfrvHjxnfeLGkpNQR4A5
USL4Ql1uy/eYGfKP4wUHXPJTqS7aASplFYBTQOYKQvvEWzYGm5XHrZzEdO0ENYSmHvKT76zbbmu2
tFCSrJpkqMj/ThEWZIbthlztf9ExvKhxRSs76/fZZbsEjYYq14EJ9wiWzfu02ZBo42l2DekppH3r
GJDWuDE9WcpkOVIyu0Uzpu+mnS01RxU+hlkE2rZZQCZ+F6gZakyqi/mMPhhwAmLCHzuzPivPG81o
eLP3uT+Z8IR2KpQeccLzwXuI3bTQFxZaN6S4I39TF5lN8BT5/+TM67XQCrG8mpUazqUNXpxEVG7e
XqsOsW0SNk3p0IKQUwIXT/rj3Ql+4qMrW48Lm9nbJPvCuEaThMz1zTVV5QWrrqyr4wvqQvCtCZXF
wVun9pBEtOmce6sGG6i3oXU15wb9utGtevrOHM78Bta0eNDumtAQ8W4tqpS/KAP97UXqdHKao9n2
g8WNT7nkaV/wQFQKzxVZeOmlV6pcMbdcHvI01CEIbPsPA3TVgdXNSi5zgWQO/orT5+B4Mse5NCPD
/8JFWTbBXT7Wxgz1oGLttrcABtKBhcNVy12it5ON/+oBb6caVfnDeuW5EUvfXNl7tKFaXP6VcAhb
SuVBsHfMaXNV7ZeV2+LOFpvVg+CempMNz1ERSNb42Xkf2ySxmtNjjMLpFXsdhxHOibyiRrfAHVI3
CLAV4RlbwwK+IvUGBMMAsodgh2TXFcyLTNSssuUqsxVqiuFeLu8yuhtQQGOcJEFk+LYRb83pAzMr
EUSC9NwWb1qkyQlx3VO8ojzjAZOnDZRmweif10HnKJOAm5948TtOZvLoPodWRkz2V7ELj5wXY022
m5sg2WXnulkWx8yisv61r8k8MjkFCp7Tw5ZjBRGbx3riShgD42NpuYa3+WTFOsDBuolGpr2aEyJb
TJd3JxcqkB6/ph2EAaZ3y5nslpTvVMklSlzzkhp5Yfeqby0LaqULiA/XQYhr43fDTo1xykNDVFR4
SVc4mNQFxMRdyjVlD5ytk8C/wRhuitvoZ5OlhGCf+8JS32tjas5sRkKbVXjsCUg5sNcRs6m1Dvil
F832oV8Vg5iZgQb41pqfhF64VlrRGH7rEMYQN6N+YwHPDE4Zr2CYm1llPVQfP9bHqMqHDQT1VKiy
CbrLmYk+Hi6HnjWY7dGyjZRNOE/ai98P7f5gJJ4EBLVsSZ55EmIDNenOOw+eUVGjqyf3lG7cqKLN
tHk7Kw0xgqqc5bZdSlcLUd/H/QqRf3/PqD045VcR6QAeh6NxnDPSBqxZLZKGP1wk0zeGxSQYVS4E
NWl9Jx+56jgBFvbpcFQEUBkbtHro1GvZf3EQc+LxR1c3gVDZYHFZyZsF10oIVggJZ9H1Xc/pUqWH
ltxt9EervOrkWpRcjWmMWuX9JWwLs/Zpzuv4kBgZScVcmPY5XbdddGLDHEofRXtKwI2mWvK139Fr
RT+Z15wGqWOq3gy5hcysj94rzu9oGAtgy4UW0gykLwkoq1hlMvSArvO9XhIII59bz6mf6kCVIqiq
72Z6nh1/ygYKyogzCsHGn1mxyDn8GQ4HF9+gTIjVZIX9rXcVM2f1hTY6JrOh5/kUeU4QhpKra0wM
kVLr/Bz/rT9TrNjZ+pLPAT4b9n4LjwPG/u4IfSDMIBldT7fwUMoYm/X/bus1HRmLlvmp0CYxATmM
L68OqofVlwvzolMpa8YDXW0+r50d/UiPkNEyAviFR098smG+nqs5Ic35Co6UKqbyFTQOoKxDmuX9
n4BTQnrntL8sqwGw9TYhIyP6ofTxXNyMaE1E9zl/BRjorbKwr4sdNVsPwNz5ObhaYVEbOheiU3TB
23tCBP8LxvXSNM598ZQPoGEManZdHPU86/SrlrBFPLCLtaPEIjrDfJ2ZRf4jZyWISnQ50KvUSjDv
gkW3N1BtYt4H4ZwHWQ59wF/6Ey7rv7X+UgiA3p/XjX5kNyhpvoWAJmoGCRZo9O5TaE+Ef+BwISqI
OBfG/ItjIHUKMtWKYDGpPMF8K6sjHy8GT/dyBNzsk3mMVPw945DnHvvAIeiVbbPmUGmJXrZc1W8d
gzRzsNytNhvzn6lgbDQNP1zKU2YrE/n3fhlKu3j5rnJxfMTdhvgMKpl+7bXwiCCK5eAci0hL+KYN
lbXBRmFNh+iMoXOe3GIKa8gxI8GFuNy0mgc/Qc2YqgPvxG+UP64wPR5L+BwBixB4OA9ZlBPZAxxq
kjBdnCPpzHlhYsfEE2BvEpU6yWQEaTAtdvBOdUyQwVVw0dqKNyNy7NU+t4Mxju0LiBm/N+d0dTKJ
oPq5Ce6aZK31gizqQExAeH9IyHz32KDv7Bss9tfEYicoMaZoC2jKBSvvHs84bU6trxE2oamLvu4z
seKitTjw4e1Jc08shQdZnkMFz/GApaUvdbU1V7bD2I/nOXaOGf7bq14WgBXVd4W9vSY2KESFFegD
BIqEo7PGyejwjJeFKv063c/2ZCbmEQ3KoxqXBgPtt9zRjfSPRcyWGo/CoijPEfFymuur859qhdE/
V7BkvTay35lqGkU6OeDKncrhu8yTFWgXesGzMKh9qr7vov8hqrM9IFA8DX8ThlYP2KGzze/zLfDQ
1QcgZgCfp7gSSrmy9qtJKfW4p5WWFkww8SXWY+EcPQzOEamFU79yj1gWNXKjhvp1rrYwQOXOptI2
SuQaUPfFT50wXeLEFQ5i0wv4YzuOaK2wXwwntpr7IV/apqDCBuKHpWivMAzVVMT1kG3hvOo+q+kk
AlyM581DvsaTGCf3j9O7wlz8waFRLSHhxBKbkBFlptPmxZ/F343RM5Ae1g7uxlPIZ3ixgXIFLVS9
Hlj6OrDCtCbprP/IPVxIA4AdvNWQWoU+VwUKsGkdj5BMohPuwEIS6mQQpKeIF6pg+kb3LoCeLsdu
vzb8Fz/P097YOfCq2cSTd6AssMf50LtSwJ+3frT8D8wjnlCG9VYmFQRUoU7dHJZgPFMn9VFn+1Ry
v+kehb4vfypZiIjsRuRfVt/xzXGdnmufenc2P4cL54ZkXsVHjrWHO3kRMBzqplz7nb7U9gqlFr+w
Llj42UBBgXIARTJLvQlICH35y0B6EtnSPR1MTU/VGQa8LUlVlcFuoDAFc3FrN0W/vcEEW2pFJkB0
8TYxJxU+lxXNa8XXnZJ1bsPY4K6d/laGElovfXthdXnWrCju14BmaGr6A9B/d88tgfmxYEPAgs+E
3ug+MzhvrZ1aiZS0drna7oJEVYvbvZ83s0Vkv5qrqbRdc7GQR5CVdu163oy6dd896vlzrBNgg8mh
mT4f37EZOCkiVJorQmkgbSq+NuYBKcVngVQS472r5D0wTz8nN8D8khCicibe+QQV40EcbOEoEnSi
yIV/8omXD+3SVLCztC8N3Z8qzlAD1CcXdJIsd4apHk/WjtQ+17qIcVYsi5v4CXnN2/8ww2cukJBN
9PK2O1aq466do/AHF7jWqkGUVWJoDNc8LNoajC/uxeDzrx0JfFGpgYGEXmaIB2+hWbADU+hiy1MY
RsHP+k/nn5ylATc2peyyXu+t9rUy60fpqaWy4ZyrLSgYg19/xeGC/gJwePDsEHSkx9iU0CE48tXf
TxVE1qy0/pDfzhz0zeh/E1kxjRoz5ggvA9hM61gANLBgx66TKj9wjyabLRypH5e7O19BP+l/olrA
OeMb4R0yL0YO0XWD+eN43sj7ChJ4KqIGB0tOLVK6D/Q4oheWpYTLXCFnVpsCrCm2GS2TY00pKi1A
UmRK4I9gxEMRW+K5Inepa/5DwORGolHh9JPp16U9ljz23zdf7AF+GmERCS8AwrO/OErUQja85RQ6
fNp4qWmex/Q/FFK3gHi8M37NwetoIt/wBtinMCnJGke8KlkgzeLDZ9fmbFO+tzHAXoOf5hsQX/3i
YMZlxVx3mCjDzpsi819sOonvd4UVQWHORPhPgqc2u6TF6ahDadu7XV2LdFpRgsZU/PobGixSTBsr
V3e2MPV9/9U8ohdxU02vv78Zju9dcUkDfmS1AoouPY6b5G2+DC1WS+sy8Ka+Hd7ppOpN6cC/aXiL
ZiQSUprylCKRGC1kySJJPievfEMSq8VRx7nr1TxN5TBAhBneZQKVWWrUc0UfLX8ltS9iJH6dZogc
vP5i3B6B/1FItRODF6OudokbHx3TddQ1JQmUTPsxuKjFEPUiou97TvaiYCvbUKVIGmSDISOtlHL4
KLOnIR/RvCJdsX1TQCMwM8/anOdBRXS6mnB6357EabsK3Et/ubECAfSapxY0mxffQhuxmRDif99q
Q3Pg+50pmxRO3P2OrnsHM+oIXYS51ccokOH+ov0WdT8gsaCMqFviflvgT3k6TZjoviRVgl/09fwd
uf1xOK5EcUvkM+UmY4Cluhm/Ur9ubTvo+zjlZeyjUuJeYeQCBWsKvknrQ2ud5ym8IXIprJJhdhVw
gw9nFSFzf6Co+qclk+PgVGf5TUiYj2dMUClst47XWldLHt3FaaUI6HVc/7KhLLwJzEExQEACrB2j
qMeHxXJD5Viwc5LwQ74dsPGcfK1sUXqUdMJBsRux/z6uNxQfxpIfe8WPo+s0x6PKRISz7HTPM0dH
q3BmmJ0w5SfcZp+xN92DTpRJyf4CRCUHDM+faOHSxzBJfdbQgmVT17kgr9+eZUkA+gsH7lO60KYl
W5IblfyEU9PRPLua0bUI38QUoVzfv5qJrNFXT3w5aO7xePKWdfTvcxejIIg8h2vzYT8VowxwFB6Y
U8YtyhhgsECNQL3LkxVusJrx474G+b6r/BqDlid73YhbMbRnb5vB7s8SWufG0FFMJaFZvKcbqupC
Zu39WuXb1zShaexhKNXnaAX1Sz+4oD7fImLJT62UWg/bPYV2tygPQZ2Vf01htuIfn7oAxBLzrD0H
xkTvuYDquqoAsyAphrNQUNUIm/JY/RH/lbENyMy9HEnd76yqYLf+nNe8OcT4PW48L+GcBMz9iVGv
h0dgCTYc6xF0ooZLSiZiFaDbXigbe+b78z6I07tWdZcaChSRUkRTyZoSynS8lpSllD7bPavmGrXT
V5nwf9jGbWAcd8UfmFWRqJ3rT8MAV2NRfiMQd0Mrg9vy/YmGlDDmPO/EjjWgVv1pQOorgj7K/lYR
zbrQcV+7fubbMfQ1CuGmUwLBneLthyq+UXwgvnWDGcRoghaOnFwf/iO7qZ3Fz/n2LqBqbJKlFrGc
AO2vAsH51W+drqnDOX1s5Lnfoxfm9euD3dVTdN2qKMiehcZgUoxah8FVGttYyJJf43VDBioEXGqZ
aV/5EmT1DlQpEG0BjudjmIIrcAel3HPHWw/y76Nj48PoHQXilTsU2Xe7y5vXfKiUw8kHveqIURop
lIgJAa5btME8gp3IJlH2eI5qyvDxRF3qdxldRttkNKgEBqn4yJ5tthd+Ih2n0Bl6sYPpNHRcNH4d
p2vHtB9voO0zDe58IC91Lj4eDR+eaFVuBPuLqs91FbBBRL1abcPHnPt+3VwoQwV4cdrm7Sby/gLa
DspRJIQsgqCQRoZZOI1ssHYr6cFkm89s764wfs7EawZJXoHjuB/6AjrYdeDg5gZBszIiEHQaFJNI
126lZrq6krfjZRrvSK0PiGfq2DrZjewuPBejwttXW7G+9F0e/hOMe/G+8M1QM2On7Vr+On9H03N7
wyYqAOX7ahcveiDBYYsz1zVc2BEKm5TXnOQiRiiQ/anQvmPR1aqneiWXMEm7Q3I/U5Q/dwm72Ynq
HbawQ1EivdE5eM02gPlf5kAyDPYMzvaDMzrznWSCWMG+2MN8qa+lm/f1EB9WTdE94IH7Z7cRa/rF
GdIdhDrgW5fnHexflLBZDzzc1/L5VEIgBJzSmEl87Aw5x6p7WscdQApb+Ty95ch2M4KpO1W5IcpY
j0dt0d54YEOvmKs/Wwo3gObYEUy8nmYaG4CY/DV590ddokEHSV/X57WZOGtedL8u1PH+Z4AT1+T+
BFi/0Ocl2/2Ph3W00Q6faMgcBg2y9RRr8Ct5gRPeUrlyFo19xTvy/pNfdWPEnmhvQyp5xhjFNxS8
4j0oKe7Ts3nITL7wnzyEMELBftuX02oLTM4/Ot+T9+aLqcBFf/G+XF8F7h63bg5ZpE5PgQEbOvct
EXMpqpRQpp3uW3GcvNDYUYRL7/4XMSABy4WyNG20lxgkGHvZrwyHKAVj+d2m0/okOKhY9nmdpv6n
IOfI71lyiBv96xABxyJOUx8HOiYK7r4VMZkNebuEyDAczvHo0sVvjTK4T/UTXbRvO7kW7JPw6gfk
kpGscvCJEwKLV63l8BC+yh4E+UmuIDYChrC8AmtBgmh5+IPgcr7gCe/9q4DgIkd2dUA2Bhwgmctk
EY0/PoN3vf8xJkGkZjiiPF0M/uwyhikDMImlMQNn5fUkjaNtcluW4Rn8cI9sIGRtOydX8uIANHij
l4B/lmUQRq7ElOiju8vanN1MTWHPrxc8RKpMq780C6oGnCXAj++SOvyXjcvt4sDauGmtMpDSj7hT
K3sjl5jMZl7DkfoOAwZjlmZUTcyqAU39lAaGnDECtaFQ8xOsDxD6ckUuhrww1f3kJ6czzCzLvsAt
M7TcXCQBwUQ6nz1nir3VDgQGhDrLPgqadMdO6Vu9oGQ0XU1nohmoa03osT263pVhs9ybdDZZFNTQ
MsrqcDOC8ZcbHvSi7OoIIfMwFsyu5c/N1zBd0qt0kIzXSTG1cjwNHarkxci1kebXSJQc1s2LNEo4
yQT0R0pFhKCxY+bzRKElilY/Wfek8q8sSh8k6QM5dxQmgBznA/rROVhEH0BcyX61pJAoQRWogA8G
zh6ShyhAYm9aXO18gXFGxizuvD7vQda2ANufN+yevvqyXeeNdMmdzxxzm7o+S+s+KQbDV15NdSB/
9gr71bC5GaJiwgvgvYZ1pZxqlsc4Hic7e+ow/V83Tec3RAHMXdvoNnwyzRlK+FCBdPU08awR7eks
+FYrX6PnTkuCNUFEiXjjHchqxlF8BA1YWiLcq59mrmQLnPZ2jtPqnD5BlXr8PXZMd7ueIuMwbAw3
ldbyg/AvNpEEo9D8CibLP5LPXNvQlhKc5zFD21FNQo5py2fmV7uAZLXRPl3C/OjfPR0vaHo5DAXw
xbE1KxU43AcBHtxSH6jgcRdJQgFmvafG70Hu/AvRZypwzYc1bebcGCf0rynffYKpptk+Dx2oZBGx
LxlrA3rFSiwOsoGImZ03EihgtFzUg4/NpVh0XB4Se9CWZqpyOeXMNaE2nA4nrbm0yBDfvYsZ9tz2
Fl4Dxutq0NIAoOsxfE87qwf4lUBTVdlMhZjfKqhn3yZnGjclEkiw2HfsXUBsjLfkbOPA0qKdyAN9
9ccQYZywawO1+A1sRisNR73O5FGJH9IqcZ24L8HaA0uRwrJK75cz9htHw5MiBKpTjT47685O0RNB
gDf5yqyMjNRjN+wKBxBAewAmnvqgGP4rBth+Q21kic9GwmTPggwQeTHeBI/O0QbuholVIqNF4bY6
a83M6ngxcj4lQz3gIKtKZqfrRyyBsyWSglMXS+P0lk8+B3xC5g/v2VkI77AyKw0Qzx8ZQRNQp2QP
61m05hKkNbMF5NTa9Z0Jh9e0oHAfBDRP9NLpHhBS4xGGZUs05mmpX9bGOUHd+ydO85XZ9OmgXPBP
G0HpyiWW+xPwt9PuGZWZTCo1ZbHPCAEdEoUKiesmReN9ahuCjTGy5cehxQWUKpEx9medWhl3yu67
uR2VoYD/huaqT+hCBCpv7Hfi/nOEdLWnCUEO2pBPLll2jMTSDWoexMjKBbH1TUSpiDo8gXcxG6Qq
Zqs1NpZQRdnKlqAgRueVBVP4hueXa7S0t1UrbgDCgB8MoLHDu/v+SGWv+i05ATVKa1xyWyXv7T77
7caQ9RI5FfoKacl6mmmKS5a0IquEe9zQJo4c8ypRpR/Wi4jZyg5+AXbYBjtyRIJujY549c6CQq5+
FBYYfGpKKb4G2iiCo6OHBp4I2hOJlf+bLeTruok43LoIgHg+zer1gzlng/471VmEU5jRRrOKomgR
e69egCuLO5cWWF8NY4gVWZAlSDtZnJi44MM9HsjIzdO5Ifv2xnDrJKNHiJaDu6PvyT6JDlxOJ5JG
EDh2i9/ovY9Rm/j0/RVKLyKENutAlMm0b6nJxOKr/cNTM1Nm7/TKUUx6AbzT5OjxAEbVNJ3lvnks
57wHsD7U5yWmsM4kVHmkFtujcwPGcCz5LHFrgM11Mm2Gmdp6/KMcdyU1BYMJwJdRTeMNmSoU4eXh
Ic8bcENfkLbtgH6jxhokfCCPn+u2lJ4bsL4qP8gccU95Dm00n/1D7cpSVE7YUSUEJdOgzh1J9w1s
/6ITqjc4+YVmHyMZ3UVAmSLdjv4SHDKYqzjUyrwkxFLcbBYk/a51Cfh+h498EmJwXbEt3wf85c5N
b+TTmFKfZLFaj5e3nh6ysqtgkE8Rx+zioXT5/S341plWddCUNxkcpb4Uz0mIR251e0DYbcmPBiyF
nGZRRV2eWL9fRNP3aGuoLaaORAPjDuAUbfwfxFnKjTc8Yd54+ANuMfSxf2/+FueFpwDXMF9rwrRK
VLjDufH2bsL5qWeL9C/1nGJw9anIpHvC343wzeZjmImXCAq7j9m9noysgS2V1CuBKiUUxCiajY9B
r4S+N3PwLaTnvR5UUu/jO2LqYORcE9B76/Utw6rvX+Hfcf12qxpSoYou6HpSDDSESfM6+bJgWRQT
52wQIVl872Da7bJZxp88/Z6N/D2pZ6P2Wj35VHbd89phsIW/A8vNLCibR9xZ0rxJ4XYIBnZDqxBo
UvVIbiwkRNqTLqwRi5KgEwETMnB15Ga+tMtMWGgZka19zzQccdTu/amMXq9VGMfa6by4t6Jxi4hb
eBQDJIx5sNgzLZx0UJ5CJNtwtPbcnlF/hgsfwYMZc+HS2Wb1X4hDkNOuERzPDHwQewJXYC+u3xQ0
1eHLCxuS5JLNTwQi9Vf9j4BRaE0Tal1oLjSfc0xsyxy+23Cvm2TTrzxU0ppX6cTEhaZ8y0h2c5uu
Ymiza7djg22yu9t22y3Okltp9hVHj09NWZZsrpy3wtm8r6gmIgOiNQzCOdbb3s4iVQnaHmFWVJ2N
mE1Aj/PaTphb/Vn8njXetaD/Q65tB4SX1jYw9x8ZbKt8tGZYMb4+RudbmBr6AYUXKYo1jFXOsaUy
jjYWQOiwX58swN4mVt8VC/3FnooT5UtrT6MEDCMMFh0BfHaVF1qgUzz0FTZ4V7QuW7I+FTL7xE9U
rekEgFSdYPq21KyZcnN4ItI3RR753gAbIzEBB1QBJaOe54/b/st3xRvKBDobYt3nu7EAPHJ48Fzk
RI/pxp53sJWOugFVuZuu6NkRp/HKfKX61cl2NZLRqSu+yedB6iQ6Il5udMjnPWae61o8BHtRxBG7
z+2N44wjlS2WSwNBwFr9XQhgFXNSEmseyQm1+r4u9/Mq4DgS53YNjDn5uexSYLtNZGjprWNyb3QT
MJp5J6X4OiLxe0UJIEuLO8LOkqaCXVpnsdpopLFrgXTFCdAt6pJA2uCR7CLx9zjJuts1JtyazNgR
VwdEgt3ccsKOAgHot4/5GG00hjjvF/1tn1Sru6qhpYw+b3j2efWMcL6J+gUPjchcNFMHn4UEyWRj
Wchc6wJya3MioMw4Og/oeahZDS480nESqojD3isg9Qy/aDrSLlWeYIBg7++c8bquUdvsI/TpU7tn
DkiQKW+uCVZApalKn/5PPCBBP4AxcH++oif+Nj4jw0+4jqHMJOvbIhSLtZptwCVXU7k/p7+mNUUp
22hy2fpXcrwedDNpbDV4nhnpCFXjgL04LZoA+ir4ojPGgSKoWWqct4D6hiKg+HE0aLZUUb2gGjSo
KIwv+mRFOs5e+rmbL3hg7SLpw9dLcuNQVvI4e8YDvhVkCGsJEhSVutK+Nwwr816AvEAzyj8vB8S4
3PRlyQFQ7kZJtAfTZicNWW3n1cxyH/636zlXEX7UsF9ikPacv+oEk9KvM0mky56XMzpXI+/8VY5g
xE8HX15OutwEInyAcQ+I3x7nqiiJFnxE2K7nLmDY1fQPIkPhq5mrNG/1dpUcMD0NJ9IKKAiMSzcS
fFiaGMLGflWGH+c16y2LVJg8cgjBT+tF2zuQndJFu+BOdo1JCGUlrih3EyluCGC3eUWWHAxc4GTi
ajs3+HQPTQuWDDp3Wu6Mo6r6hMtqh+rLDzhB6ErYNnNhrtbSFN1/yKT9BX6Tq+rQ3DyErCn/7FUz
C2V7AaZlq4vItwKTQpDrHt36IA/BadNWQYMb0jj16kkrR8RpOyeZLgWFjMARChOgwAqPmukgLfKw
DqyB/DZkBGE+3iQnk7JY+7RT5QfJ4AV5+jyvuE5LCtYE+aGBz8/+eVHPr3rx5WserpkIZvGMiTNc
6zhAcXxpXZLAnAte9MnU0w/7Vt/neV4yTbq1khxSwFjrFbBQEQ2yILSO3MaDeRWarRCrP9b59HjR
DUqlVs1gnqBT1qHKUnMBZwi5eG4RuqTniOvZzoV5oLEQJrfuSSWUEcjXmtlhOmc0E0iMpjNT7LOE
hysB/nbWMpq8Lk0sRejE/qDc1DteZqe3hIfUI36GpnVNef2Gx0S0uoq4cy45Ex0JAa9BPDHrekLy
8D+Wh+Kmzss8HotOoEZWBzebW4aK1xcv7emxQzvimK5wX1aOJ6pncV4oxbmIOwLR4acByKzon/P0
EiF1IM42GC+pMwCRyoimQk0QSWLBsg2coXPhBwpPDivktTaaCVrgCmMFxoJw/HyYIYfFTJHGjlYc
Vv5P9l3OQ1JvIoheZgMKs4016SIQeHsw++wRlsbkIh14/1V8sbfESSlKJ5cW8/veX2cBdW2FD6++
+P24a0miiXgXpRbJ8xyKUKM+gdW7Oeqo5H9BO/QVA3mJY54S8zswNOfIC1YwR6tjv88VbbMq2mrv
QRcVxXRxsfdY6lLPP3s0lzQCFnhHo0T+NBBDvB+CERx7ILnhCVQnnb78D+3R5BFzmMkxfC7Iwo6d
v0V6zsi8Rr4b6pbNTbWVZUwd00o+1uAcjWJHlHT9hAv+fqiynGbGBf97QbUP9X/D7ZSDizCUSweY
RDHLhmJxpbf6LnWNoDOyAeIfek3o7U8HgXwFbiN6NI/UINJ9JBBePP7p7WWJyL5iJx6YV7hIlflZ
N3SnB/il9xFbbA5ib/Z6dFhKpOc8zFExADFvZDZ/fCfiutG8WO2CAPW5mnw5CeqbM0F74U3+5BI4
EStJKcCtTGJNJcX2n2XjC+bpJQcTXVIGRCfrKq5WJys+wPnPT9Z9NO7qzHqUN4NJ5Kklk+7sg53C
55dRHOqul9OQwLReWCNYUapfHxajVu2m6V0R8weMayojhoIa2CkYY68a9GK+pq1rp6LKPsOLap44
YJJdvgahHinSgOYARzXX4ZTdmvP2nJJC3kg5soP/T6KK/2pkTvno+5i1+O7imMwOp+6/gOm7YWr4
lQkOCzdGI7C/m5aVgxHXWqDOGUk+vCLQ9+E7PUrlMGSn2IXp3Px3L4/yYP6fLE4AQCt0VQHY6WuQ
+bc1p+G74BgusXQBY9Nqgt+iZMn4QcNowAzJhWMIsxyNPcYoM6JkjIglipclHZG1pfhogPsCH8xK
7z4zjOYHFQgtu7vTaBnclkGk/JkzVcdOfzh1/UywR1jVifOSxpMExuwIkx8Zhtsz7czzEjEDlHqH
6BkAGxfbzNSIxLxM4mbYT23wzsXpqGhY6+c+mPn9VkpNoBl6O0CeaO/SO34K4d8P+q8jrEve9bAw
bP5RyW8Srv86NQlR3+PIkxDyMl7AjovLd4o9iRRosAuXAB4zmdFC+NQhOLOdCS+U4gsrcwbVxqGU
hMjZi6yV0WLMh+3iCAWpPCbNhVFOtZmBOq43wY9l3zuUzoDNX87HTpe0UGNpFsTDDS//ocL5ovM5
f1tmlum/bws9DDb22y6/oUq86T8PbiW4iwazdwLOCeoVJgckoLBvDBI5nxokxTn7CNY9lsZAvFJX
QahjdND/STNYZ2Vmc/DRe8/feh+7jd66zGeSTZNqhOlwcW9wyY8P1nUcbpG6WMPwIPRpoy9C/XoJ
tIfCTYO+f4fuCGBZR3xdw1sbtGidKITQTPE38Uj4eSLJQrPvAGfmD3CCuC5ft7xgGiHYG/gzHtn8
kSzmPs5fS7GCM9MRxhfOS+NPPmL8EMwRQlYDTxP0j7FCSwprgxlbHMItsCGcNHPGtUGnzsfhjtf3
QBwc+oSgUBPssvV3G2sw6aIAtOZKB2b7RS2Vx4CjmJxpRluXFSO5Fmz2JW3cRo5C9k58SIJFkY15
BH64DDvZk4auqjV7b9s/yGjfSPjaiDU9c+hi/JhYo3XdYp77P+OVAb0hZ35Vfhj1906WlqIXxYuv
cDZKFygQqvGyn9Jsrhgx7fzTjlpkwACnHCJkhdExsTrm4oG/iw6i6c8Ed8EG7s7KouewtndcSuPn
b7PCvbJqhS8Wioxq0OKhY3+nmoVR8PmsQZvCWtq/dknK7JOG0qYWtce7RIQBXQzPvuH3SqxoH9xB
gmy7svuBf6MmMErPD7NhuLDmFPyAU8Itdi8LHXogIefv+4F619OIkg2w9v3f8Me+hlCwrVcxKCcV
6tV/+LKZLYrkokZkUQod5CfGieZFbRcv1A7BjDyNRa/nhx9b4TsAXZRD5ZESOc6nZDAqjmk5KUyH
Ia/fzp/Fq7/ogL0xfVdxUXO896S3MqLclQ6NH08zr8Hp7sm93tsFmyiqXKXWkzodwWjyrjUT4lB5
jYPNsJajcJfsDyvLBqXYIxjgJsC8hk4xluWFMgotFpQ7reBka9517fPifDxU39NuwGiwZ3lGQpli
10nV8g5xF7DvJQysu4H/0VX17AZUmdB643h2J8pxjthWfpUtaGMbAZg4Eoxu8pEygOe+eM7WiRVz
dIRPMcqUNYtqQqXR7kHs6/RCdJWCWwzjqjBJTb/SkEKlum1T1bSt7XGWYgxqsLSYlOc9soH4BQj2
wYyRVJZAarmr0VO+a3rHANqiLvia0Ar4W4eaN+OQj9SveNp8TNLFn0Jec/mxN1red4clR4j6LSCX
5QnZgXAF7vLohb2wJpRKSqp/0j+SBHiirK3k7MQ77PUumH1PhR7ZuV7T1bwJjz7DCqs5jsBvJTai
0zVQgtVhcZ1m8YULFbLPtZ3OyXDvpYmLQZ7pHts0Xly33V/gbQAtz2vZqoBLVGsuTiWWA79aE1X5
6jEt5tCsAAtrN60bsGRJjy3pGGc37JKIBEexHmusB+WcNFLaP8A2jSHZprd6F1mi+5qJYOACWJNT
/7d6NqV0g94goeOGziq8S00ZUh9ggBS3iNg4hQf99EbASQTKQYUdCyyNIMTp0nrfO2ewGhSu0iSJ
uy8RBupdbEhRZ03SDOfiF51w3MjxXsieJa2ADKVgf+jQR4a4mpfeFxxlH5lNDeNgsCgihvPkv207
UT0g8lKhMgjN4VLRjW9I73yvgGfluVKFuEkpGMLL6K/8hskyx9rG5EZjfc2wNenZX6djca0Yq1cw
5DbupfYUCvzUQuCzoS1ofcsPOhJDkog+EbxnnmRdCiM492zWYDyRynH9bRlcVq8P9OyL2pinKcg4
VWl1n7ruo1HEFvBUb9Q0JYBhAZm5Ahw5w4mDJIR/uEvy/7Sf4DBYD4hGvn5FiH65f0YQHmyOPR6/
YFslDLt54nDUbf5c+ZWCxd3e1I/vAD3BlYpECpj6zJUwjwB1VB/gmkDV+rijyPGBB6WqHjfibFt5
JN/GGfVjJOzTO2rNB34Em9SmXO8lG7tg+Xdz3he7Nf6TGDaH7YLIQ9/Ooim8iXjJF8bken/cTniT
IUBDUBjZDAqyeboDG7hE1YX8jcxGKV3x0++d4cfm9LEH5YFeix91ys81T652YHkwxjRtR5sqkZ/u
hSAy5C2QhcDIqbUYPSUN0KtMksbN737jes0D/DpSt65uFjTt9H4kY00qCqLK9QmIHTgjwm95WuQ3
SVhmMoLFAjL7LC+K2wPOiwN7v6RIpKVla/VlFzJT1vmmpQlvzrmZg9eLoA19SyiVXbJxC5DzM4Qj
UN9WPn3eqBZqVNZzeCpN0kwuZ/BFvLEoEb7tKNfSxV23JEg2U/CSySFBbsJUaFuTWDsKHFx4DLcz
MzEDHKU3cVx5LDNr+Z30pcKPM5ydpn7hXuCrfjmI/Tuo86ZjKU7sk/jKCwZ3tOesZQ7rQbbKWBOU
q96SElBJh8EFNRN8mXXfbAoWH1SKlgy2/8h+rvLm33AFyCz7oQNnJo9vCSa29iZXTLy+bm04lHRe
apzyZBMQFHZc7AEjWHFwBXgJ7ou4u1VwGwXhwqbNgzyU0IU8syzSOBGOezmi6YAiUwzA9tzn6kFk
q1RCWRfRjUr46WW0yLPxcFDPxVl9zFY9Qld0hItsHduV02NW/Er67J948SYUJynug62nmuSFNO2q
p3HEzGu4+kVWN96mO7i3uu0pqA6KypyvHLk/n0uR5nOLQGnTgqvRdqSJ1nGzd7pF2kf4kdC88psF
WlFw3bPeDLLNAZ6qcykA/7xBqaWNdJt8tl/QZuqqFlI+KK/0mVdCXPxt3F/M1fjfY6i0lr1Evrno
/Lg0ZjyV6N+bm+NTAPrwznc+Q4n7xvn4gsEVekFL3HTSC4sYyppUXZ9FLyP4o1BE68IzfCpUmYJ+
EWdV+4JZ8p+I9ieLDT9EpuXJzovsFBOWqg/CzpfMCWVBNfJxRrh03Qodv46mcgh+jAzzXQ3d4W6O
eZBfmYBgAWRydkkPwIFW6X9vVL2p7y3uYQLWkbDq23HwgzpTz6bGWN5xEg97UVec0ZB77r1kCwps
YNVXmBX0DUBFGVoKojWglVUF3M6X+iSIVVCwk8gHzUFIg2jwphITjU97sNnDSoQPnbWK8Tujviny
/rU5XlNpeMq6cSCX+on3/B2SFJfeeY7oGxr/Bq4BRT8yrFrxSxMwCNDJFxHjizu1ZIRAGeQ3+vxo
rgV2eB85WA4ZynXkH6y4UD2HtF4fPR0zj52KYjONjqKS9HThgp6abtD8clgEAtDvGME0bG68dlSt
PMrhsP6SFRBzNdTJ5An2t9ab1eB9NZtuGvmFvka6tgEULHGSwq5S+GJQkw7AzqnxnW43KGMhMPjd
3TzAUtkMoNfmjqEjl5Nh/dkkHNtSRVt+kdLZffs+pyDgU7VjHhoDky4kA6+RmH+8VdjG7c/Ctqv8
YFouWHSVar4krgWs5LwxezBvaJR8rXJpdnuDmGUhIp0wEvCbXMBPjOWRiKMytOz1MbScwUb4xHfy
V9TRbTzd+PH7n8fGlxxYJm/YG8W+WppZiyvlyR++oEYxQZa3WE+ywOAYgAQfT9guMoiINarhA4Ft
s9mGn19dEQiHfKkyb1VyLVIB72HSmvCJ/9pEwip5ibL99rIWvanSSp/8P9N11DDSwf79kAHp5u4V
wmNFQGddoLF3oVUIN+cPJot3cpkIhDThlyv/vnCZtv/Ep0+Ky2VAhqhkPfYYhLU5NGGU6mu855Ab
RJWD50tgo8B8fpzcMVYpRafexuuRIv1YjiyFstQl3+S/81HqQfTehGuwMuWYibAtiqELyLlK2ZC5
w1xlG5UU/Gz8v09Te/KEqu+baBqPyg/s5Xs8XqWRmcEcBKmodX/YW9uLGfw2QcdzY0WidmWMflHK
Ox44GJnKGrscRFSdUcYJhUm+iXN3Q3a213+avtlD+MMf2+mzSgWmg/KLHUp/z5W0M+Sr2ymmTLOA
BYOn2RE179SCLzLOniZtkHF77DDJv8dM6veTUYTiBtVmVjAejd3u07RwAoJ68QL/LD0PTFgl2bwV
+l8O78TU2vFfNMKOZg6GOM/r6mXxFXC9fptxuflikrjtBWh3T3lRgWQUTaaaDWMLIqFov+/wUfxL
uRXoDt0blgPcWDqY0mBVgecrBLBKBGwy+0JH0bfST1eLZnNNjLNlqtE3ayVaRCHvo6LVlFRB+fom
XL4ZkH/hQE3Rx5MJSC+3+lRRc8VIDrQJTiRTF5Z7FRuLjD1Y+MYn1cmMQUzcPofJRPfDT1mDANxx
KNix3Q7n+dGoe8WpXQHOHEwIj/8KgR4S/gCmEmrieCSc0sxRpF4QFEs3c58Qzxgp97eG+YkBT06l
6CVnMTP+nh/jpxvfAYzvtQDSuK+LKbqiRAgR4z0wZ5uPutiOMBCV8kbKXyZG82hD/qLyiwj8tE3P
sDiJ5UnG1LeOyOR9FY6lUPTkNPFkKrbPlN5SeXkd5g4Ss4jfcBOoBUh24OIHvKmJnsCGYqo9RkSo
L70lJJZhMztGC7U7pXBpU6FSxAWjZr7nS+yavufa4wDWoRIidFFerJxfOEOk6Gq9PaD9NJOw9jiP
X8YtxbqAIwgj3EDcqeW5JTcEdjaZKh/grMdqfCnWVEjVmQtw6QwkfNDwRbOPnpLxEkoMD3sw+8ot
WJOuuC7jQv0N+mP2Becdy1w/NF3Xmo2zy7UjT6wfJhNYgxyPc9vdNcRiLhjylr8m9tjYrc9fdKYm
YbzoB3nU1QJoSlxjTg9YlewdWeOxxbYpw31c8qPJ2Wb3xtZirAp4S/g0EmrIdxGUYVHaiZICRbyP
VRbm026Dy8aTAKpTKvlGDdjXJa4Y4rUoRPtdxgnZfrpmSQnK8nAmPwqg8vv3v+2RE/8RGFoPQy0q
u8B+mV29ZvH1Jiyb627B4idy6zIjsBp+WawCMtGJr9edEzpukTFELyKaHgWFVMni8pMQPWV3uLng
Mi2yRgj4G9c2hKLPU48dmUIlsPxMZIc/VJ+feD8sAPfDysifetATjh/9jdMYbSnaKOHhIzRRlfwg
CePxYbsPtl8mmFpK1sxE5Rmrg49wOdgBhPJwhw58XPjjU9J99WvijRbq7HxtefYMBzZHJ/pG/N8I
05PnhY7N7UlANndLOzbOfYj4LQrNCcR++IcDWMl09m4aAua1W71Ba6LYlxFwhOoKp1nLJTeAgr79
JqjkDIEy9qsvUlJeivRpfE1pFWpDAZXq0ZWE/hsuXcGZ7LlnVncfCktTWHxkObxo2DpzCvmitXVa
ILDvr8ZPxE5w9clCLyjq/XYWA3ZJXP1UN4hn7MeJPEZVK3WmhYQFscPy3D2fmIHb0GLyXlQgatWO
578KEb3aDPmXS/sE4ufwlGTJd28r2bhUJkY5et5CwjoeSB7AOSvlnyghZfocY3xOgIraOhAW0Bh5
Liqa0If9+fpVZMlFARGeWshtPw9W97pVTXc4/Iv2tigcub3ACzySPgI18xRIW2KP43kq5xiz0+08
h7xcFEAmnfWLbGi9+3Y8s/DND3n65MR0gOx0ISBjEm+5kfkArDrKUPp6OWhtDIV+ikQjknjJoY6R
LA1NQweqn0cUV7TmJfcXYT8kNIEtyeEbn9eI1B1JNc15qZCprZbDnN532L4WEdNqkSsOurYdJnwM
EWqm/sIPv6Z+ImpM3wotB9JZYbuAiPTmmzBNWyG+0tFlDK2zLSPTcIA5H6Zuel/nGT1DZHkQuykP
xtA12v8hyrBBhVeaHlrRndHwaHSbn5e0d7xo/C1F0mr4RUU4WFHkuY3JMqeBIgVsSP2xlUrvl5H8
ukISW9bVRbyFUKxA4GcJA7PVKMOmlg2t4zZiFbWstrel8zU2ty85LQzoFSvdBRTp1ouqcT44wSR+
K1XBXLXk4Racq7N4OOlDkdI1FSuNEL5UFfxmiIZ9MBKHpe9eIvzbm2RRa+ds4jgwymNIxVBMGN+L
yvvJ3CQhY50pXWZQXwI3YIvWh79V1HvRWgUWE8qhCstpCNMehbYFEQRo0temwSp+MPnT1fehZoFc
pJ2Z70SvGrQTskY2kGGD/XfuNNk01kQOHWUNMgiCSNCwIiJNcV/wOtMsGiKZT0CdU7GClzkpOuO5
j9/thVZVbLdNVxwo4Uu7l7csJKWQ01oyx0iaggoneIJNMf7fqY29OidZuKD68Ay7gCjQQVhjGMA9
mptgJ2OldnlVapEAXL4Nw00nns41Qlwiadp6JZnv7BG+sFFUiQ++aIXrObh6N2+LF7Aensbh6REM
dB2r15bhCtJvOWXtPNvAM/aQoc9+bvTUE6z2Mw6snUfd0HQUK7VKk6Zk3h7zKqEvOsSrlev50DBo
y47vnGpDD6CrZqP0njpMC0W6vVX/ReLA6tlWsucF9lovdPe52PjW9IokzLVEdjA9L0NkmkEmMtw2
6OnsqWjCmqC478xRvwMp7hAws7isaP1rQR176j4uJDpzxvwUxHbfP6b15Bf3t2+uk1mmloICp/tz
ZdJQLGkF5BZX0E/yKw6BOXa8nQtg/EYsESNjeedf4CIqRSxrs6KbRM0lOeJGK0GeHdsLgOtF4upe
SRbOFEpgb9z2Lu62mMwAFnZJeFSjR/89q+YW0s3SsA1bf208AZgNDh2RBuppkhreEs75PjQHWu4F
1gLJlv+VuFdmN4ZZ1VO7Cgj9YrbkVkMO38kOpJi1buNzcLEFIVWNfIFlqEMmpbP5b09nV7ku517o
zWkcljIxD26PFm9JNIK6m7gFpiOk1XumGHlvTnO3EQLXhR3eSOIE0YCFXSec0Cey7Y1eD2aI7udy
OaGTtxUVI1n5Kc/r8LNez0P9gfjBQ6qsH3SGj8HvASaeOsZr4/A5SzWmXkM2PShkeci12c1vR5GM
yCd57rpW0lJmt3lKgMK8vShIGCU96+RFpUUJqs41hmvtRmb4XDdvga+IX21dSdOLb4cl+3nEi+rh
wmEHb0PpjArJCx/mLAyN83VK11lF0KtMRwC/eJMHL2yiZ8cts8rd/rPItafshXJbzIXnoyU23wwK
pk9qCORbaDDlkdsh56F7m0BeWcJfZpysx6AhOLswdgo52CdIk8MPHrxdiy2yBdox1RU3ztICnv7x
e8l1HJB84Xuo9sLJdNJ5jusi1dCwsgDtPPZHk8O7mj3HeK2jsR1ODhExnQ7UaKEiRze+GYF8L6I0
oThoenzq6f4GO5NjFukVeeU83PvUc7TqDGjd31Efd9wizhZTpuJ4g1zrAd4hl6yVJ1mFnV0FqUvE
55Dli/V59gYMtP3NygbklicqlIiQxJwbXnWYOq4tGYU66Q1y4G+NcRv5Ss1hbMU2f+6cpOyWwzU6
RtAVhV5HiavbKcrBNOEK0ZsREvIcANbdJrim3VjCCVdApwfy17Wv5lH6IGJoeAFheiJCIQfataRS
2L9KcnbNc96pm/v76cjhsg/Khlbd49o/bqimZg9UFo+qlGYk1YNZfxq1M08OVpvqqD4VUzgUCKA2
iT5teRllB2iqxn37P84LtqvxlbfdHcDgueYTW/xtF4zElGoVF8O+SRzDQkuHRDQhi2fU8W0sxqPv
tgQuJCiPYbvF93UtLLHDXyXWO09ndHL8nfIPuDcdDQ5G8s4XtbDXlgZfw71BaFMrbSL3AikKwRLf
wKLUbIZK44Lx9a+t1h+W430hcjqJEeEaH/x3ORz4tYBiOjBoyyq6k0+Bd0CcgrWQ66LAXV5Nbytt
dGsaUEkB1KNnBCCXVXwoQerFEFP0Xr9DMZANmNMHcyRFuJDmKwrKJYM5j/7QhmSIpylQ1UIngDEZ
3P60uSM5ywNgdlnHa8BZV50wnbu3PdHi1yTsDRNL3+FFlwvgemf3fcq35euxOc7vAYVIDq9LFeDO
gj6dFjCyIqVPWH82ZhnaH/vCZNVCrbKH0ZdhjFXm0lC5cmOf1EFMHZJevu2gFWWKKOKhgR170U1x
10GZTMGYzdMl4bJF0LAvlrk9RJFWovT/aCk+GfYuwSgcs/0qE1oQEjhR7FXaX+vey96zdMBtxtGe
Y8zhheuI3HhRTtZ6JJdZ5Uc5hGInaA6gw+JwY6UwovdLNnjx9bT2HedFCg/9ah6csthSU/jXNDvx
cVmhh5v5gbCkssicxCZMDmBoDWc1BwSG40JbnSNwiSnfXgoGIiInv9o7kS33m/iJkX7PG/6YrMrH
OwErjSDn6MLJQmA6g3xNf5dhHZjAe8pKLz5t9vHcfyCR8639ny7vcIfkLGEbVEfJ1O7bTy/HHuHQ
9XsyA/JUjgUXL5lIqBxd40soBE1AhZerEhFHLRZl00OXTzKFZoNG4CsXeZntM4UEX2j9IGZD3Pie
yl2Ln8/UhrjCu/Kbmez884+8Zkgtu3X/aHVGO0tI4r64gQwFKaCxI5quWE3edgmD20axYRJZOS0V
CmBfKpeFh7uALBa9n2T2CO7vTd4CFV6N47sUF4bf/rr+1VvWIPnbOsLsVYckwB1jI3YYMSXOCF4F
YOEBg2o1vNav3o9IVO46+rkxukOUUZmmmmlWEvqlDNV6eXq4dd7ymg30bgsX+pV7RMmcsx5rkZ+b
1ldiEq7gJQj5U6x//LmEE9Q6vtDccs6pULG9TPjN51C9mbo6C2yWrV52p2HWfCSkak6qyiPuK03X
fCXvex6rfwSubqwDfhKJc+Lh9luxW9eV/PcrEQP1tlZe+8uGPdNqX1my9K0CsY2uMB1zq6lr5PsU
idLumka/IaxYxdKH14CEGQlJUhlpxmkTraWDnNMB7V+5AWYTPlc9fxrYDW0Qim94FdTI2XC/YrLH
QVmLK8CG/iNU3TLNt1No+4OzyXSMZD4Vo3e6yFmcTzmDnxQhvC3sXCSuEwdOILYbJVpxxg6FxFXD
VcSyAypZgZWYKC8jd1uhh5DSXAUT4bh4aAJ/weVTOODNthcoCz36x0HgL3PVlnA31w6VyJOWZ6c5
HfccCQ2Yv0ENRp3NU8JPwhNqM4Ow7fZEn6zm1Z98tyrbrXpJXd6VkCMd4X/rhlfJIRvWkehNcLhp
IbqcjXU214zrLBCIu6DdA39xc5lIYHyNMczFOwl6eoqE4OonBUfh+ePFzK08ully8jExDtJnwAdn
bCY629A3fnzCPL8iZcAIm2qovg/1hkq2sxhHDJViovIrYIJ820XH+6CF8BhFM0SPzeQNAqRLCQMu
26h4mTu1O7scFfHuZDQYR667a9TlYeO3ZIbUCJUgd2DBZHHYoevHK7mhJtBgL3t96ZKkYnjRYNop
Q4KJ4Ag2Slnj84GP3iK/N7xkH+JuQKmsklXDff+0EanR+GEhQ+jYucIJVu9tyt4m8ZdcAqMuEBCy
TbzbQ4jUIRfvBeAFc5FlT1Tia3AKN7Gs63y2tMNSyK07LL078/HpRlXIDBIcKHXMjd5qQ8sVeVEN
3zVDniAg0mbAThbWmyuFsC1oNeyEWnR5++MYsnCagymMdEjA9bDouRkFtTJSvXIY/o6TSJ5S7Gy3
ieGql4t1yeYA2K5ImE6j7S831TjY+LFNm1KpNY6U5h9Ii1iy184PTyMYoiWXO0IszNFA/XI9mwvf
sAHjVxtQt/8WH6TfrDmx2+Ppgx4WNiPIE13lw7fKP027XdSFJSqGwp4Kn3N97Mvn4pkPsc+GIqNL
/0ml2iWUYHNtMEnzYXpsA6JIXB8N0O/dBIhkYi/WJ+5VV6jFgK9igY/jl/1OFAz9z/VFr3KiYoLe
reMiL5Wiq0rFQfieeBOGsoHv/pz6FC4SLCL3OMcaMA/+w/FST0HUsGbezmOmMjC20GOHk2g63TFh
orRK+zTFEVeyhA5b5Iqkv5zEBWyLoKVItTfgc3Ldu0fY3FaeTNnHLQ+Z0RR6Pw6L1iQiDdQdHElW
jnaIvQxedgJWXizrPzVNxxYpIUiYbFapcu5cyAflR3JhwOsWqVyIoYUEQkJP5qDoZAhh4/Re2CWD
9E0RYIbJZ2OnDH7aStp8s7gfqz28BWRrAe0w3ZYuTLmnQUvaVg9rJYH+VJbUsBDRRzNlvefZKyqC
jEMbj7DxBGbTo/6u2/2kDB750JDh2mP99oRg15oKnJVvXu9+oi5dZ7nanQl/+OZGi/zrrZkPpx54
A6aH0IjHYEAgHFre/O5WuvwUBsrrg1vA9dbhUcpiJx5LFpLZS++vySwO/v83opKPdlY+fuPwRJ0/
o2lFWGw2pekPh0TvbKG4+4NgJ0mXf+MwxcWhMtWyluLz9QDLli56iN+QBb1Tnov/ozX1MLHTvjuw
GRf1jzM3JV8xT7mbrIk/OoH1ffPGgBHWHaHmHI+t3UazY1fu5qzfsTZTF/eTRoiGg3kz5/S9+4NM
zTEwJmuHLT3+sD4235VWKeZSOgXenv/joP1AIk3OQV1Ge4oSVVungdJfhxvDflJhX5vKF4ooitrF
RNPDj1JyFSp+AMLxx8aML1dLuAFphpbgQwMGAjl0QO2M706+tc6gA9ZtcJ0lMlZWALPHP2Wb/rBW
Skg7fDEpTAX3ViH4t7b3nIG+ZXB5ZFkwa1EMjREdpKm/oeZEqZRH7hzF+SmMr7CAxPzG1Wd+psLd
rpHdyrBKMKHrM/yofr3swW7I6p5FXeOaO3Ut67g+f0Kc57ZMKVezen/jX+5Vq0Q1mM4D4MZCz0/L
kqOwFLy1vdE9MtQXzlMfhwGqBw8lNjlfhPuuDTmNln3UE/3Vg0wYaEaT41Qoa2E/u+Lu10QDZrzJ
xcAxsqpxG920wepQjkVTesgtQR1T9GVLzns0Xm+K0AH7+xqef/vBPsEWV4DA4MIgnhlREQAvcprt
dNC0h/X2/rkPcYqCZBxDTBrewm/ku9on1xXxhG28oSv8rdE9nkVad09YllSxy4Hjrj0Wl5fEK4ag
EwZAmPt3ddyIoV1k46CWZMrjHjfNxE8dYWSB/ieSw+iQlNaxVzy2IcsY/o/1PfEjkoUbYsAZdcHN
O5qN9mc3crvW9RatME5m77WU84GJx/EyYjSCbWhObCGPUTLAo3LcWJyD3Qeu7eS4bc1h2eDgN92h
ba/WcXMbEcb575xHIpxa7qg0V5824n+dEQ5zL2pXpt3vGt46DoLkKuyuuox0Ks4coC9IPqDZDFXE
cTHHiE7RvGXsTUK7D2ifGnEbDfUqLN3U+op4NxAMIf4JibZ1EkL7Y86d7qjTySsJoScEmtZiEWbU
mTcZz7QEcl4pYwe4W8Ih3+8zN60IbwmGURRikN96TQ5wy8Lu42WDvYx0iUGJwtIoNqqX+lU7mwGj
YaCMp+R3jjgEXEpyXlD7xGC9w+h5vPru6WvQQgII7jjiL0Je8TxKS/vYAANysFeA2vvTduS8sHEz
xdPZKg5BPPpK6IdeDvTKGdgDIZ1cZO3ycpDSk8q4O0imz2AUfhhB3+ZGqd18JWFGruaZH1R8yKPw
XJ8vqVUH/ukXzrJwG9vUTV7Y2rEWmElpWlVQFrpfyhuKlNIOhFQCzkGA/jmX5CZntyoEYrblcfXe
Hteg9qGgT9HNSTUX+0200eWGtgaToG38e/DFth85l2NxvwGEjYhUu3Zs2MZ0/0GkceKIrU5HK8o6
99MGr30DvO2Htums2CDrOZeocB/hUhdgAX3+xdhF1mw6qbFvLzmTAhWVmZNM0kAraPxL5o9Patyb
6NWFbGbCSdH/+qMUv71FbgSP8U4+1qvCh8/fzQwm/F1PLvZZWWlvHXPmqCYFfddaSSg6NWOkYaRw
D/YxrCI8EAtyGvIVe8nLf5W9iDZvHBIl1delIelW6f7XTNY1NWShmy8zlYGpzjrXQnZF0exGI4N6
kg6ysd6LgA2NvuPZ5HAva/gkhXwMvXcsT/3hS5XFJh9dKTU2rvOso/QwcFWwqeVxlS47A6Vg/XCl
VOalex00qQaNd6zm0+87X1yjDVpIg4121Xv+yxnnyX40MsJHBtAFEQxU9tX4MYJyPSPHkMy84WoB
/vog/HaTMiFCCjth420wlxvoNftjl+lp+76CV4k+VfP6piF4CIYlXp+hOgb6zaBwL0eC2PZEXLCe
OZ+kC6HhhR0QLdkTzwcfV3DoTGF1RVQCZjikVNU8cCvAzZxdrQoCbATGhopNHwcyFY+6PVErame3
QVmTOlo9/H0MTw5EyUmO4VtBJQslXjUxan1Jmvaogz9sIyPK4VheUN8WuRpNUCxyUV9a53f4DiY6
krUSBBnmaACrBiB24H8CVizd31cQegnFtcKtXrkv2dxAjgX4zxeU+ZXAID6ZctNcJjnc5ShdPi8T
he/6Hk9a1tjC3brMVhjRiwajuhcxfg0FVLTtQHxVU90mLBndy2Rpd2tiYfGVBMPF4uO/NfEMBacV
MJlrGgIyf4WZiiRpUB/x8xe0W4MbNbLu+fkdxKRAoy7faSZF8WnZbrHRpOYiN6mOyM9SempRZmjF
x2RhnkvmCRSZh7KG/AqO3wWIZbSI+dS1zgYw5SGY4bq4jIWRzQ92J3Q/XksBdTOeAzZH8EQjk8q1
VNNZi9YHgGCppP9XJ+HqGHjm5sdIieVSa8jQVaf+R1/ViCyWN52ptKpOP0u0SQmhO4nxSe/Sc5OF
KA+pQw2/BtcQcrJ9IQ/DwtshbwV1nOU1ZD1+X3QjlGgJwseMiVNoCEfWSiJ90wJmy2K+9i5BY7yF
CRmfi71nL33T9PVip/NWcC4h3qkAp08XKyi2Nhl7Gr/AkhyUiONKe++DkArgsCUoQWQYjVa3U0Eu
F1uQ6YStdAllvFGgt5SdgwkQXuXomwsZUtxHQGWG/RAlAdazNIC2sNYW/UQId8G0BImHV9ZuyxZ3
P8AUcP/XdHgKPlFj+JDCLpFFCJI1yps8j2pGUro3SYoh+/KyYo8D4XpW92PU441FT1KXvEZTffXD
hFaTD8iu4wlIvlcgBzUKf+vNzuN94jdmGYkS4BcA9/eS672AKC2xaL62l2xhjVsewHOdg/4fIZ2I
Ha9kcB+pE5Eq8w/LvVl8axII1F9KXxpQiY1Nlv5/2sDP7KLZdE9f8U1ltzvgCNOSpNx2Ppdf4alp
cUj49DLC7A6orEqjZZlPhTwprEB8VFQRw5jBvy3xRKkJUTfLwg3gJZu/Y/3sFeSUk2sWhOF+IEBB
eCwdApuRJj+medCIKblm6bEaKgOH1taLumVHSqCk4uSVMpXcOCw1hGwhFYifg1uIwfLiWF+frgw6
ndHNjEhDj9OtL9JhYsoAY3UQisv1FDUt7I3xel/nJbws5w0dTrAJY38PF10AdZkEfcsR5scjl8Ot
j6ZfQvzIYjqFU7qf0q/E1Etb6GGasUxTkhplUyLOFFdRXcNm0oUpeLMiL+CCStL868o1b7MzWliJ
yv8Ci3GnQH1N8kFs8c2gKvLLmMMZ6Z9adR7KjNEN72a5GBzepkcpfR1NXccIz3Ea3tOsPHu4Hplg
+HWomMP2ew2Zi9QznQfPAhRV0ERHYMxeqBZSb2Pif/mhF2KYEWf+v8pUwrbF5CcPuki8956zBkrJ
ytRiGzUCBhnN69y3tlhv6FGDUmoKGq7Kw4egkayoFGk1QkMejDnduR+lE5nwyAAqSi05S5pGMWSA
4jlGWiT9+HW71DXlrjJeQtk3rTwvhRvBEy44dyISkl8UIkvPISnOjXFEd+xpgXpU+P7f+/hm9/X6
I2Th8Pn6uNTAj183aQ53y58DG7gF/Y0AXy3GRpmGy72epzFfd/9SS6RGTBuHnUgiSeB83pgrQNqv
LhV1kzsFDcFr6PUAUPDxIylls33IVQQyQ3vha5FvV5tWgMdCTJCikcJ5pK8wb5ZTBdZs8KhHOLwj
i9BW1/K+sz5RKOp1bn+0jn1KdIxeSw1P7X3gfDsuuvx2gN7vnjIt9a+GEOV20ZpCc5g9iYxF5pA5
YrlWb3k7ZZornsIgJtA1eLBtGTAtkWze5p5+SKAuy1D793Yy17l7bFwzxanGSQzLrc6NLiNGZ0+A
249moyUUPRhG+njXwi81kd97xBG3TOIzZJp9/qA4GpLOgcuozCSsJCpnkjUPlCOxobKQpHabSwqt
SPpdoRWkL76TnoUh+gA7UN2FO6Nw9kXliC5YWZeYBfZJnWUsvqk+nZES5ZhE9DIboBeDkzacT/3O
EnFu3amX0wc7lwQbqBvTbxm4aJfS8wDLTwRU/VCoHD5LhlgpIUW4tZb6jnmTu4NW/Z/MHckK6tZR
4EeO+gYVa3EpFS9KmAF5CXVz5B0OPhuAD8EpmT0OvOZ/113R6XRSf7jK2LJG8E+/03EX8QEzRMH1
2u3vphver/BL5owrClaL0pVRhjuvtW4w+9oIUocdq+4+shODQBE1YJewy8i1PZ5Tw0pP3jjWz7hV
x3Tjz/1TreETzMVMBhSrrZJ5UrsuGcI7rxOqGrzqWS8s5Ge8UnxkpKK2npOIMKFGaXKWo7ZCQRr2
baNpLS7BKqur9rRhBQA8jUR2HjshkZ4gpWmniL+MhzJIH09lVKY0F6s7un0u7iaWavXEIxElZY0C
MHLspFuztHyods75vHwGEy5FV+cdHy5lgdZOm5YOqqeTTHvXXJTCPhFHlhFyfk0t5cOecjgQPU2d
PqggdlssXJEtTZVgkegU1o6E/42URnnuNSLvTBZMyUtFXmYkgo5dUq5QZiugD9uz0Aib24XXS4Pv
zfvfj+BTjjhlPZjhV9dDbTyfVbdLGltD/hjT0NkUb15kmJVRZrrZlwIxbzAigKke63OYsroNaDH/
lDpSNwGDRB8LRlIV5G4IBzUP0FoMPfwQXmDUZBocYxEQPxcJdO1CMvZTcGTG92U3EKxcykaA7B3z
L+N7Dre9mh+LgyQdGWKLEjr5cW+775mOJLdwrKcD1ZnaDCExW0Y9XuqImfA45MQ+vF8ixH4Z6AL1
u/48EyyVRnvATOONJRkG/0jcqmudajWs9WO6baBvHUVuOJp6wsGiV4/XNvV9ZjvasByijlqJ0Dl2
XZpsqM30Cb9/RA2r9nLmLfO3ukz6W0tAf0/tGHGW47qNzWfycsS0stKaAo7qDtWn5rmRJeCf2EHo
sfIKxmaNTE8Nk+0BUuxxD8Oej2EKXo9G+VZsgcWtoookSOmJKu9fMZU0kGgZxoR42IWxXyUQBhjb
CUZsvBc6/Vn2a3WTEI/f3qkXlLPNaEvvRrd2Kwfl+dB/mac5c39FKh2r5jNU7yxDSil6ZWY4A+Ok
26gS0/F2dmQcnfczVAkKooZFqR1J5pibKdHLkEUCSr+PrKLNQrQk3VQuMIGlSNUplobhgUPxmQ2c
BkbV6UV8jgNoCsIbdaqFaIIRUaw95h9YBuxwBDobR0nEd+brs13hVMKsbael0dFWHTQngs32TEKh
/W59QLbmGANhn5edkA59oN5MBZJp44RLlmW2d9RqPL6DWEcuhHr9GCJGNiBL4JPoSHBirOC1ST+k
f/x9Uh8Uw8RVdkxEaG3iVQXWWUgCHrW6WRCUIGe9yJ8r02hN2p2DVwT273nFx6ZZSvafdkhfhvy4
eQaUh7ZWhHhBEHFL+Ta1aIvxOW9npsA+iKUjT6RyOPuyezoU2xqBx6FNnSG0FOn/s0lXrT4SVa+r
p5wM1pXhjE4mkCQx0mvnuN0e2VmCNP24D9r+ynz35yurNgGD8dYSV0xC4SscCtthqHc0l/9kDwM+
4JpN7mU1S4ptiVvuOV+L1YAPw88CaxlsMr2L6PjURvaO8JGlxjyDydKOIALQXMEtVoo3Bge2F7T5
aUnoLMZFskxWOf5iNBjEUjEknH3ThBb7b83fJNlcFLwjXn2wCbtutmhujUePHQJ0NIr8U7Ugk4ur
+yQx5pouw9uoOC7h62fiEqQ0ZKND8DjiYxcDZaChEfowBNalCiMAWZVRf4b4LIOt8I8MEWfBYEcO
jMEKJwlufkcYYbAFONxf4ehPl/jLJVP6zKIHBqYFeYE4fzRcmPT/D1bwDJSVjcuB0k48uWcf/tfm
YdPAoKdPfbPr/NwO266iOwAP8CJ3YDrPJjo78V58DCCHMAIQh+g3lY3fTmg62llcuu6zm5p0UK7F
taRZ5kBPPTXJrLpHu73gpIrStYBuIBYp6aGdS3o7QQe95s13vJMR881gRTSpfKefAsf5B7Xlo3rz
TsFkAXQT7Yzy5XmykFsMAb0M6Aw7B5LhIQA+sobaxy868EokD/pWNRW9riWOHBPZC0VKF7Irp59P
uxfH9xy801dDdO6nDeSavhSujVXrShEW62xLNe56KcmdnDYKBP5SBk4m0Ql/NIhjoPbiphHSP9VI
epg44R9qJptVwcU4Qq5/pgVuMQJ0PMIAo1Q1ztqKFQXFDMGDdrG2+S6PbmF2nX9wBqutgGgThnnw
VxqjWtjhmJD0yTm6kiWgBIUigcJR8iAeDu6fDPbmDFYN4wld/zJ1O+0m18nGEumA/z7p8h/KK2N5
jminE4n0HilbcuOOLWd2/UhtFuPiemkLpdetutSltg7cyLZFQLbtZuUAN3knFj30wW+/Rpt3NF//
EC86mTMWHzygyejFChOtWxwHWXN5RwmAdjSax00oRw2xg9pOxkzx15PbtRu51gORno3ZVvVaNbcL
zxCcBDZNDQr05U+mHvPMpgcFPhBjCprk7izs0CawtWDIHoDCQXSKWVSX6okssM5zC+h9CHXFRqlB
e4KxIDIzDAHwLYfTNo+MbblN+ulv55tXbDf9FDwP8qFPqF5ZfpA9GSUmfiZYE+hCAfp1rKvoQDJs
QwPndaYRE16XHSAfoXiYq6qVCdYg8s01IyYlQS/Nw9aeHuV1DzBmt6QFuslG2YCm1LwcJ5Us6N4A
Kh8trKwVdH0xPxIb1Mz5n2qZUxlbqNuZnVOvbN2T/h7FDUE2Fx+MHcnqalxwcIPJyN+IjHmfOqjn
oLtDE0s+Ruz4YIOvkoF5mLwU0PRRXNC2lbPrL80zo70hV2lwg4c2QSDftTjMqDlbTsFqTk/9Vi0h
RqV88Urjo607WmAIBfOGAV519uM3HQ3AXQyPngEAHIa1hGR69kkr2sgMZ818MBglF9XIwO365uzE
7RilPAs2nCodRluaLavACQtncHZmVCHCSB+vVVoXvq0BXyEkx/Axtxcb59WOORi79wSVKv/V/RH9
QMkQT/LqqtYNtHs0m02tPEtwGh35ZVnQ+m0h9g7gwAbDyBN4yn3Loyq9ApC2cwhH4+QeOt4Ag4L9
xCYIDsT48zqOWZEK2HsZdVqPzRQ3ijP6NX9R0T4j0h6g17uG101MCUO3kxiHQp+7qvd+M2d7jGyF
7hl1BjtTF7HxOBIN5/3v0oHvqPaKufVuDLr0e8Z3C40eeZUSKq4iG1CuPGQV8fGJcEPP8IcrGtrM
J1eBvWFgKA+M/PlwTXCDuQCj2fht+zmhE2G0OXrkOLLbbG4zocfsCOTtNtPYHBS1MuFWonWzWv3x
XCeG68RmUlxCkxEPw/vGI6q1pIDRIQKyRP4apOcrxmXWUHYY9qw7JKf3aVnZeLf/PT4YJdBSVYFX
VxUTfZoTwSFjL3AAIK5cS9gHbfMqn/mKo3YBMpDoaeAJDZewVF0LRB9dFsYopeJjZjpMwHrmTqNL
+T9u3yvc5kjeG/l1bo9ug4BvbRa98TIuHa2hLDKZr+/Koc0xAMljJCUYET3PF/rc2/LUSsUGyARJ
P0s01lrKbcDo0ASe921gSZumFPE46T4zwBIo4PPyKc+oFy9i0qvL/Jnt4gGkVRMUH6wQ76Y7EJSS
5XHhlBJWhM2bkajeAIv02RD/uMym/vcxUDrWJO/AO2175sunxgCH0Ztp/nqRaYEVYPldR+Vs6pfg
GBRgnqVGIJtEsJevCoDhObhk9tXJXZSS4zHxIwmL9PR7Fs1LsGkofTnKE2/NswK5K/a1G8hjGVMA
aN/SZvcDO5q//KWnOIQgIBIwg0KA63ZjzuxWdDmAVLiqZ1haxkMdXYpe/KfYmmmdBo0y5KliLC6m
vSaAoVODm10vgQL+7QX6+qJhRqEabZXXHLlqdCMLIf86FQhSQ1p8yrHgeAtUp9D+rQlEpHijCc3q
3GcPwxPzYalwhmd8o5gqy+9nLllymXCOu3W+xhz7BFkB+OaIHeyTSk5FfGBXFziE6qiQboEcxF7M
dc+R0LNDwtdrSo4V1zdm7jQzU8SrqVx/WqOm1xtwzDpqDWgKw2qRSV8z3rIOMrmbHCrlASD8GnCl
H2QcK7HD/PMqh7As7El1rOtJ9sKf/1OK6DfsQt1G2rwlV/JUilw7r2IVcl8C/Yc6qKNpl2t6fHFN
OmfFEPPfnvTm+Gu9rpFqfDGBzwtJ8tq9RdC3yXVxW8YmmMQy8skJ+PE3Q/S3n6woW7uN4Qxkd57l
s4yEdHlT7HHHp4nFOkvTFd/8fFTq8Eg3Tjn0oDn+hvJfwGjFLs7vTMZZ0wEe7eYAj3Tlnl3MmQCN
IW1scKyfjieMBQFxOsovl2oXH66W/VBgQkiYN1C0gn7U9EamM/upHRpvefHar43d4AiwewvSotYE
32vZ7VRD1YLcPXXeA/OsnhyloRH6NM7J27+Ck7AlgiTfIfrA+OE2C32yatc0AMewKD5xiQH2FLp7
wRnqt+jhWSz4qKZ3jO7P1Enfc069vppQ4dFb0xbSGzXr8aFFN0Wx6RMCwTYObbe5DFGXoo/T6ivN
wTve88U9f4vpSIASyngvRCAvWTzqgHRpqu/100EqOgMqr0Fd4ecUqPfboHGam1ilkTpY1sSus+bL
diCdVRbRHD9ICzPvObCspIktWiIrhv7xzA+CvEYv/hLkQbCDPCsel2wbGJiYVEQzndjL49JfUILd
QxduBmPlm4U5uExG+BMGmmejzDPD+KY5zlA87eK4cFVUlKSGBU54Udmg+8+31waXc4U6fH7rBd2i
2Kj6C4JVhnXt1R9z0rkJiM9Pr41QyjzbbcwMKYQPpSKxXEMkBXXIwqVM7ZwO+9kZlMIRRZCvE7Ls
UCbWsgrNm0RHlAFfJ3AT5K/MvwJClwg+9qO7jCSraqpoios45R+FF1A67GT5/bKPIXNEsLsWl2p2
GS4LEDcsS6BZVYAeSIokP/AN+Gx8oqDf+IeP1enUasbmqUdjv9OLSWuLqjesfCaCrbh+sjPNLFYn
N8TgcJ44ropdpt1wIT7sD/Lwp5K4VQBplg9teqin+ZZbCx7Zd+QI+KCfFKN5l9guIgdVGD/1dWWA
4rj4DoJHiIB8dV3Jcfr1Zmmt3S8lS58qXdrb0c8vTY76MP3jIOCBEIjM6igjfA5h/IoVXttnDZFo
8wEXmx3gcu1iCgLj837VlGzYTadM5TeAbU3//suGKjO2Xa9a/eThtQy0j9Uq8TMrRfA/gzqrcOL7
zbnYagTQm7zNu+iM31x6XtPONMyTqvpW3DA3+o7sAv7T5Oznwcbmj9H6rK4Lz9SAd8w/wG0x76bi
uj2aYT2Wab1oMxwKDAEL2DcZYGYPkTTDLbQkeqlVlik2L7kTCznuBVFrl/zBcOdMfMCTV7v6Xt2U
z8kSinmrLou+n47rI/zuBovM5klrUWQmVQZDtIl5sKxUFiUrJEEJP4OFp9atE6wK7854YmNTo8S7
kTKVch86XepvrAJ8ymj9xveTHN5X1X4bGD3ANh8qRYdtLosPy4kCBpZCQm7ytHecKADPavD2SAdC
t5EUrDh2o0LjAlamKwXRGVxzIUJGIMPQ4pLBiekP96eRmweNNp05EVXKnLwq64+Dc7knoWN8+J6Z
TpmDDq8A5dFBubaGLSeOrBScMV7vwZoxacmMxlYoAFLeA7dfoBXdtemk1b/dvjRhJnIKMIorvLYY
j4Xnjq2PJ+k2zxCORY3Z5pjhLHXSO6kMG2/z504GfdRbHFzGXaIjBDJI1sdv7uhrmOVplfKak2LO
dnzu9TC2nX1NmZrv78uy/AcXZgZqMoDkll/gI7FLj4/Iicauoa4800ldjbW28/vwU2TpU3C6U+1H
87M4Q/qQGDoQrIcf/SxjFMOZchAIbr1onK6Y/uPsqwEe4nwHYf095gjF/ziMd3tgdQw6R+TqqGdQ
3pVxGXwcmBpFPz9OqqQSQI5Yae6p3wxx/jNFtbaXxPRYY69J1y4745tKBFZxDP9fidLvY4ZVEXL8
AYpuXtcduvcFBwvFmiCaMAVdLejVEyapHj3EDNF9pfN3h+cmp0k7o4s/z9mI5Ogo1ULWUyco/7I1
rPalGimIV0K36IQPPXq6U0HfhkBZuaPIQwTldylOljBD1IPRz+/HV45eNK/kpygN3Xf9eZCB5WfC
8//zLHyluviynsTUK6EXsNYkwzmXEswiLF3+tJiefGBp6yTERUUJ0LVZc7wMzFhIxhXhuxbBUxSW
upK6blP/s8J29KMXYwnlzznHaErBfC/im7rPNvacFiyNj9CWeA6SYycw2S+6HFaRIME374cYjL5t
I1DXXLp5kn0t5imQU86jOYJ5SfoWgf9GV1PeVY/z8yjqoMGMGLso2IshVjxJR8nK/4jH8IdyTwww
55AxeXQqAHLHPvzgmWU3yS+jiA6o3G0RpLHTNOAOHK8NHjilm8l4QoPazoJTJzAKqGYz0ILhH3+g
CuQmAtBb6/Psi+tBEVKZ3eQ43gGb+n0kV/gTl0nS3z+pOND7T5vJtuAQlsgowEOtRLdeP/WsH90q
OqCI3d4hrtB0QlzFmfCHePkvf0P1bGRHbukzmprXqvu7BNZkXKdSIHq9WZ7DFUcx9avzNxXgGdse
YS+ITIDatyEKWsPruZM362W1ZAzaMz/iWPa1DZaKGGUuzOfXcrlqk4MvVDYSFCzVOWy7lZMMdkIl
z4wuixdh13DDa/k9vBAlAEBx3ZVc/Xv4dSCB1olCydOyYvRZJgUtH0/VJpawng/dRyHW9UCbElDh
xBvpdkHT8TMkj2T+YvJKONKXxwxd721xheOXuWHjJp8WKbd32VI/fDsTBZHrKjUSAiuPLMV+Tnxp
WMmi6fz1CJX3Jk1B7isi6iToWZeKQ01eCmtSKGiint3dLbYJXGZcCx8N/WXCQxJzu5bYwhhz4uNY
z086WFFeQX7tcD1SDo2DDdMbfhdQaAvUwiBtIBx6fjaQG6WCWQBW+IEgTSl2A7Q7mTlF9AKM/do2
u0nT1ZNXUwuFFiTzSpYY4h5lojcMYepss2xOAcxeQLzeqHUeZYCwzhJDpHl42+o68fcry9JE/zmw
JEmtN3eHzooChBGXtLGQejLazP39yIjkDtbPErD75Ib/gDSldO7jJEZJGrw6Ss0hVbKDxJRXe0MP
mZy8qv1nesR1C3jYho9t3ph4Pctf1iktQBR2DlH/5BXeIEuT7qt+yAiCltAFxklnsxUUuX4ZbyOv
ce8xVT63x50uxKhPOKKNTjqudXqiQ5K7Epze3VSG/Y79dUuOL4fuU46Q18rQ0nmcPppNlFe+wo2l
/mtFEG6kc0r7681Hr//etS3XsOLQWHE2OAMqMqHveT3a/+ZoWPde3sKNUVOhYOYPJkVdLIfEQs9o
uk0PFVQDbR0N4tFmo2BRiKcCFOAdFCEBlghNVvW9NCdgB5QWbA0qioaeg+LOooZlxGP3x9pdg4pO
HaCHf6XnNGC8hTgM8TBPzdSedE+LOlSCFlpbW10B2z9HsNW/0NyAR+A6OBMoqdrjHJzCCou/Ss81
NpAJiFA7X1gpuf6fGCz7UISSCPWegsi7cUU3xvJ/13OWwneAQyYyCBvh00WTjKzMLKBpJI108/6P
RXnwdUOGUNcK1GLRMzGixjpofPCxl1cIJGdl3TFTYNKW1mApOtm5w0sjVCU0MLON8eFlHLchXDnx
iPltGy/INQ98cGaLwFSx3FGJjkbCMFtlNGLkReH8e7QMbrDqOBWZXHip5UL5j4l6nlRhBjrMaDix
PokIer6UlBVatJpEhW2P3bTzJtvYU9VKyEtGiKLJQFkF+i1xrnS40Hh2i/GLwBqI/4cjNXM0Pc8a
Lrr6FNIb0WcvnUKQb2saNy1kTo/Fa+4PnEkTetJiH6jPuahoi0XGHrKQ4IFyWwa3hif+hNe0Yniq
rGe6v7UoeLvQlicDkiyLbASDj7LRGF6kn1Ss8jZa0YrzCyYBfzXyalKbIWtDeiCfnvIHW/2zQfHU
biFmnAtDTvYzL7vLwwGNTc64telDxLknI7FZSNG54Fk5b+OKObtrqV0bVRLXsB/UKiFFyaU6B/xj
/ze4z4yWVPiC4Kry8QrSrRQ6ju95EJ7X+BHdi3qgpUV84EjQ/zf2bN/fkg/Ub3PzWIJeDTZghi/6
aeLsdHPSZYudApOQWKreE3A1fL+yvXX/BCD8KIuPP5g5KGXkAm6+kNzXVWswdR7KXVlwTPJvklax
cD0llEXrbaQjr1Jasmt92zldVET7CxkXQkpSjj5sr0ShskWf/374kBkOVvr7KPNEpdi5Lzljb2uR
KCYjDYin2O9gOgbXuEcoSOEem/0Qd8rYBRqRjsphrzOjhlw8u/FXKGYVyHBiGO8Qlql4xG7RXuYc
OJUYdIHgoVkCrq8iEN76dIeyBVb4w1w+EvMJAj2cPsgYDW4Vq836tCuweUXbgTrc86ycuPPnbFWc
iZp5ixruTEWntspI5lxdu4KSe5llxDX4V3XlfQTogveDEu1huogA7+oVoTaW8O3sfSDC1K9b3u9i
wmEJhwZEm0/hMqBUhxaBgdX46kxo+mq5rcYKT30KhgOUz9420X9sYU5dk4/eAy67ckNzrgOZJV5S
B5OfiSEikV1i+1NSmi13IvQfRN0+MVB6y0urgPsFoWGnjQAfUdIKTiOHELHN8Bwy10Ja0LhJ7dnW
9526iXLUJORFtiXkKfNCKy04BZ0l/wx0hkdrYHrGKXVSm1LezGLgvm0NCXpEPCymN7bgPvzeUsGp
KjhW5hQPySTDCa58uODcn9U1Piku/mzh4wlVEz1z7VWM8LNncQiOWqZ5gLRX2qDuMV4lvDS1iFim
p00yScOmvmB7f46XuojlNZZC16XC28oFbfW1rCEaPONQaB4+ovl6D2aInvFuLeYzct/v1nL6RIGQ
DDsXZuckDRPzE79/ryqhFI4oxEdcqPyttkhWAQVEtJSkYDR5yzvL7INg2/T5mC+TjqZt5PFkMVck
v6kIRSk5A2YztLPPkO8uol0r+BYBkdK4FlJIy6PgsdkcfxSW29RIZ7r5mr00FwcyJog4XlFjvmd+
7CsFk6jhrc2XfpIlmknX1dtCociXOeoDDHMhTx3RSOezXXZLnQgJJS9Ak2l0jAVL9fOyPcti9h06
YaCQya8uXBapKR4tQUSic1wH038kS4Fm4U42k6Xvo+sCR3MITfL8lgGrNhPAgzv9NQS+uY6L4Jsl
VdbxE6O625g8X4ckoy5sNh5od/z0EfMJ7OHQF7lSYdarRkNezbWPKm8v9jY0ubuDqsL0OXR3zyaz
wBJ4ouQ3k2ulkw5WGNRDFS9r3FHLpcjHW6A4bklg5xM/gXYxr8qu/YueAnXUt9KD4azxXN/4eI3G
btcvSF32vHro+UPphKpuY0hX0w9SJXtsQIvUAHDrV2BuzqskdQpi9eSlgKDPVGczxm9jItFrXfZo
DQHKDLyYasuURiQRra50FuBL34WoSuGzPTkdkKt5S6mGhTG0++DFWRVKqeQjVYNsWYKmt7qiIklG
LA5cImUsHPOO1seeg5RtF7ynHQPGC3MWyHLpL9rnoRbzYZRaXXbv3AEzO3MfrbKnwhvfdbTBH52o
b7NWDApH6KzdDibUM0bSOHdkffP4exo1jhvsV6WMmB/Xi5qDja0Q+ByYYijDQ6zwK8TeYWpJukP9
Ds2CUGKGpeHLhvBOZlisy6sr6baJ+HS/Btisucb1yi8YZ9r5mXnlzFQpCtbxiFOHbStipF6VpeOW
GMYw4+xtcqUdTaEpdc89RY5NSSps8+/LmfKkoFkviAVHB0whnl0Rt9X1C6KLCKe3pezQxDgjwnBk
4d+72h0ZCFcYH6MNU3+xxW1VIaHvGJ/ULsskhK+dFv0wKzzPw6tP7XoP5q2ijcU97J6zUaiZPAnP
CtfMbU3BEu4Ri2MHPrmEdo9jcAZ6HUm10Dv0vAJwYmOMzXr3G0YpfWT+3ApSGCISgRQLAEtvK+yT
yyX95DZgtVBPhFwKnQ+Nua9NSjg/07Pti4dwBDz8QgQw3jJ5PuaHBIplcHtJkJIAOmps8E/0TxoK
rnLcrPS5KrZu8gEq7fYxAAcBLTv9/DZ2kEs08ShWcetCoNVrJMspmWrwz/oD4FgRdpfgDFDn9Jpw
/b5PZvnJaAzatziqkrRP2xXfMwUTUgx+zBSZP8nl4vhzQstvP2x1RD2a80OH+hqG59B5+fPRPadb
5gXSxqghExw4/XWxSsnADqGFM0QIpjJLWCZSySQMJrL1aSMIQyVDG+lLy/IKvoJicKZPgpa5ppd1
kMmQuBTpNnT+EqBCyr9XIgzDd+STkj2wDrNpfXIjLG/bVBzRkYoSDMw5qrrtVoquMnVipPGwZ9av
z39xJPo9IMd6c7NnkOa7ZChyC3W2oMITbSU4vL1w2Uf086N/J2ic2PVoHEDL6Hp0pUZKZ1SpoZSr
Hn5WtF1KJsl8H2417CevTpx4q/sPCQ/qMz5soNFRXnbCJD0diyuKKm/Wwtx1iJkNhf2RaKDt9KkW
dUC8lTGrxftQMMcO4uuKEw2n9ylJ6g03471RrqtgoDjld1jfXloFRyrhYQZRnFrUoNEnOwVvJh0M
WsGwew7qMfd3706Cgy8mLCmTHTFgBiD2ug2lqvqcHRA9TYbWGcqpNwdYzthhq5qgFEFjP6o/3IG1
Po/a0RwQNzLwsj+xjNqOX8PuH2aIzghC1ntmnlVwZ+IR4ckekJMw/eENVKksXtqqzhk3lAzhitia
w1bxIsxTWiVv9hf3eWdMBHAkS2NtJ+4Y2H7OtzOejnVXZkCLQ4qSmKnPq9Vs4phdIKpF/A1vwqSE
k/iEu7hYb8OsYq3Is5S1Q5zJ5OiWHh5Lenpxo7bR3hIel7T8EuutBtGzt9JlxbIaALXoFTt0radP
AlgEKO9naKi8G6aTYqSOVpy8G3jabLrEtmTmsDFH8ORNCAahukd055DNSyzpXDS+4UZptW8KICRW
Hc1naexLZ2O4aoE8KIfrS0LYZV5ZCrzAqQAEnnVGEdJQ/KLiioxQ/mG3CkqHZmignSihhNCiG7BM
KK0esYLPqc8y8BzXSWXR83VxPXOFR7mlLjLNgiCPBQDUD5W/KjY4+Tb+aciHVJedlu6fW0LXiB7v
UathSoMGXxxuM5hfIij/uOWOiQ9lWJHpKVd5bbpRxBKo8HBP98CNEA+n9n1sRFKIita0KprjZMHr
z6hgyUJ+m5zeR4L/yJVZ8ikA/xskJHbSu4JVhKZzoVGVeScbKI7i5YAqsChhdDtX037mQDuXtfmP
0pFQCIGJ22ElCOmQLnkBl8rX8WZUKXvDKh7bTkCw+/Mt2+pmEQx43L4Lj4MmnQ8qtoIGdC59gCsR
ew4mLZxFRgA19EJ+HMBCS9hCKErNPCUR28hxuE2jqci4fAr2LjmzrpqmRHZwgRSoIF+rlBMlevgx
3C8QWpXDjGcTLFaWNAlO2TKyf28bbL1VNipRjYw4Zp+VIbv5U/WvTJ7qftALsRbOajQ0uJI0qcBL
TTf9Tjmj8c2aeaLjrg4F/m6rKYyB8JqDEm5jh3r0b/BEeP2KvfJpycz3gjlLZffSJXU3xMEGFC89
em8S4GCGapsNfPPo3Xf9VtncKeRsEJZcEIuG4Lh6jDnVhshrzDTaN/OMjCwwxPkC59/l95RC6BDm
va/ypXITteJR5jEcW9DgrA6jc7jHNp9p8AKJexXP6xTzLjTdNiNouRCbPgnl8eUAOpJp1HQlRwqy
ucrRfCUYqZdLkR9fPlPuH6hsni3IX1QqqnWtjhO2z4GeLY2A41O//fZD4Hpa7NVBQ1h28psQS0vS
WIMDEjNkSl9hQJOSqzeBnc4LpKOhjHKqkt9xwalE4C6uV93kalevIYn6m1mNts0lkHKxX6rYwWVI
0Z71dsEvZHE8+iRrhJD9hHUBPeDBeTgynDo4vfhvece7IVanQ17gXdTCkasu8fT937ERMOluH92y
bGA3SS2YM1R9s4WbA4ew4u9tX68JmbqdVT78e0b+bwhV0uK2fuqSxI/MRzwB5lGXTxVFqMZlOAmV
Dx8V+wdQlieCwblpGpjqDGKkRH34q+HfPMv1dzed4N5fUo16g4i4rnKdEB6UQD14zRK7rX2BbMRn
MLU61tk0aGSIkbRF2ukt5p60MjJy1l3ebWFOGbfA9Z/0JHII6V/i0H76Ezdw759ZdrzRsQnYXWRO
/n8oHcGm342RyLawsGr1ehoQIRQ2r4P/1Tg48AIQ5/GMh81hVi6hVRcFf8ovltoKltZpiCBL9tn9
JduanzAo/gcoWN5ITxBsLxCOaN7FxHsOUAt94zcAKKig0WZqEPKyRqcybzcj9HZ5/Mr1oLENan0c
WS3UKAaZKnMfPRn/q+iZQb9utjA/5mUmn3uXIqY0ydzVECpNQgxBwSZETNzzqbSerZn3NpMhjLY0
HqI/WJFeZ86CtPc3yjynjaPuez2xw70BNRJlgzPxZMYSMJajPIHWP4F3AGQkGuCRQ7s501jgleo7
lMa8GxK6R+uEgpEWWDPzmwtR+eXhalT+eL6eTmEx19tbvU4/+PHvmW57E9dpi9AbXQJ38nqTE33/
K4zSXGbeVdJkcycGjuvKuY8JvpINx2aaiwY/t2QWqpr5DKcIXGWbK4JImeTlO2L46I/im7ARXIi6
w/pzxZ16Bm65zD9sGp9Iu6ClwhsEIGqgV0TmLvFNd6xfS3MempC/MiOuHocLu4c72p5V9RoS3mDe
6/lkOXFDy6pnsbpwnLRv9/sBoHYhFJthM8Khx3VISoJ5kAE7tvOFKjunmmmWu2Uw+xYSEnFNvIlt
Iqksb1ts5j6aI+KJ35Q+Dsrsua+NYRhXSS+VovwAoPNacvN0u5gqIqopaAXO7dDIvxtkgiuMUVuS
UqTucT2w2td3qLx8WZYfatTFPR7H+sEiTo1/2FbhkvHFfg1hPZ74Syyv24JCdzw3o9/WzDoJoNX7
WElIw2IDc8RDYw43WpAc8LxQSanIxLngRsse2ovxaoW5241i4T8qCgTndJcjzr4P+//972wScmD0
j7FPeJ5GCjQCwe5NznCvhW+lXKpSEAFXSZUdOIqo3cajxONBaFcWjrkLYZUIWXhOKSbvb/EgE3hg
Wyc5/OPKq0gtgUGyIsiCX5f3IHqX51VBhV+BdLINL4GPsQF3SIL0MfUF22zkizcckzTupqvCnBXU
AyOkB9lIT7b+q+KC6L0J2pkpLHUqPAlSeiYOMwu4HPL37ShyNsC/WQGm5uMiyRNwO1BNqHju3wLd
NFHxIZP9gnVU57vgrJGL3EGWi9CO5AqWaGxLz+kSNJ7EX7/mGmeNAaWJEfESkhwOEMmECv8bnBpj
PUHehBjouQffEmkTdgi8gT6Hj21Re9sgAfVw5YyzplIK3+JkJpktUQxvcqGK7cYcO7e0+G9KrPLV
Kkg03Ly2/q8+/cyWXP9feVEPVv1SRHtgSXEqLjxXdmazsdscltI27wPeLISR+O1/YB/wAcg31fto
VcCpEXMmGI7NVhOTijj38RSbrIeOrT3fl+55AHe0TDUqddQSYjP09IGGhzl3Jv6sKzdBVCZrUu9a
Du9jPiW7oHC1riWpGOQBVFpkpoMKg31U4J6/A6zsSNsmEhv9zK1srKPNNdjsMaadM02ybthtBE1P
DuK9HkVp5Z+mm4xYMEpIly3ZTtDCFGZDLHEGyKfetb3x0YpgUEXZ8aBShPiwmQ/511KiBO8uqM7C
1+LTcjXZCn3P9ibtdU1Epjc9nc1kNrb7uhc/EtfaHjKO0v6GBHTVfAX2UNNUrwDvSyVBiXUGf813
X9WhW9OK1pwceNq45jR/Zf/Qx4qoPfL+iXMBmIfQseVV+toVTfiipti6sICwvAWyFxeG4GVvnnt1
t9O9HbIIqGYwkFbpX5RDxkqzhjDdvoD/aE+fvUqDGU31ISkQFEdRlmdRfZ5JBZxuOuugxuuRjBZe
v4naPsh4lUKC2WhvNT87aEAJD+Kq3xKCNEo+JV5AFQtR2tvwZ6FtMWNF1gvdbCYjT+VjTqhP9JDO
0mTj5QGJvbBW+3lcOERRIdEDvfdjP2antrcNRi0SHKK9buFyeiciCblGEkdtrbx4vt03Zn59u233
PWq2Zccxa6oSad3m3quwjI8lWf31k18ETdcdHxognscWMoTKSOynTZmCsnkR9l0u222OgjbnRDfm
GI2nQ05UdDbU7mG+YUW4W7xMHTgdH0CKP/ibTOmCf1ofJoWulvbIvgj3IZ3+JptCQGMZ32cu6Jmp
b+6/ryLrLM6iHql+zATX7vPdIbyUa5iXJv9qqG3+ljhfQSdIi+qdjco7lOADpWcsyDExh6q71tKW
xSpZnelzhDqEiArAWRu7pfIWTDPsFsO4kKXv2dhcXulsXZCyiB89tJz1s0XUbJvrlDIqcAi3rQJs
p6rxhyrVdstV0iB+50tp0/rPx60rSCizypineFExTHBHHLLE8j5XUqhnCXU1ZhTweGBjYOcqh/3q
Lgb0pmV+zc54QmQlGmUTFBXRln+9vdeFQESSA/c6HNxR6mdSfE++100JcPEayvy1A7el56C5Psvu
hnXXTNau8D7OUdCc0SqB+Jya6ra3t6SUe2xVwq6TFPLpSFCnf8VIoP7QLtBC/w33btjYzTLoN+ZX
8FcbyySX0NhRG6HriEZ4zsKZ1xueBCLz0JwBsVXMnO/lvBDFV6WUAXC3mZ7JykJe95xp+BfqPzJZ
T2i7mSCqMr0Jo3OWbSJQkaKbjty83yl3CigKONDyrmBEmxtzqnPQKoG+lue5g/petHQIqqlqFxrx
lJwN3HUrE3SJyXAmKy6FjNHfDGvnf697CC5t87VpQTPlTejX+/lEqzsecpin/7jclRkOJ3jM8kta
Yz1UxsAoXBGVFDRrpTE2TtzuAO1oUI1WLfLVVzkUifjWMzKwmXy/gA6I7jC3/jo6YZOn1MEWvBqy
QMfNBZpyHkPN0Jg8Xzk7TCxGmL5qXNubCtyisIkA6KxZwFw9HBBfezCatfqjJ9PSXTuNEaxZC2YD
n4r6ZiU7KjPTfUSOljEXGHitjhSxtUvJfgyqLQQ4ahsYTFLaw0qw+xnPU7R7OIntuq4qeYfv/x/L
P51KXA69JvYjBy4yaSypHUTtqpTum6H7mKuhVRxRNw4KvC9/WSoUyEaWG0FWNLd30dkTUkb2V1Gg
rOo5YfUEDj8yQX6zoEot2Hpa4w9Hj0c/JltdXNIlZ+5dk6KA2HcmH9znHwM90QfF4PuUM5CdoF2c
rq7HRkbcAn+f+w3IyEL8p6CXEQLxShZU3MbK7ldfKLkRqPrC5WlV6hYuC3L3ptjJz84U4tlMZ2vN
L6hnEA7Pq052aEDB4lJfZl3z6ffdxAI9s+NdF0Z/EUXZBQS3zjO/lcwoJqmmJxuzmvhVs9+mIsAg
gzaUWixltbebIyhZLi89FjzJ0BlXWUUdpr3aOY94uZ0Spq2tgUZhzUHPP0DyDaZzLgqOXoQGl6Wc
Zd6xQNUxZvl/RO9gr/qaSjrJ9iLIdSqdXv31X73ES7hVe5xJ/M01IYWbUd4+4/Msj3aMElVnU31t
7/KeTspqUlVyuDNLFzmudG1VGAxzJ7zxszHzYQ852pSm0KEZKAcD2ey97zqxm8Qu/Ji8VBLDmNyu
6aXaMT20jY0+iSssoVdPak8gLpl+wenvvHcF/B9g01lBmg6Z7B8sdsUOIpn3ZSK+2/ZqcVu2DsCl
JnTy6LFyYC5DUIFs2wthJDzpC9PrP2Zyjd5Se/ltBkRrrIQnr8lM8BAPH3tbeCKpKKKJC9Qyyb0T
yBlk7Nbk5HajfDZnMnORKMGgSMaCiwGeT2ipmWircIGGIa7hoCW8yYjx7pPaZx0DeYwKAXfs4oTP
LUOsOdCjBMy8GpREWM9l2RGBlM/m1GPoRvZjSHUUUMf6mvOOH+jS0gkK1UtikZY8tfjCaB/50W88
H9AGQydIuyCKq70Yjafr9ZFeQZu9MRg6Gh4Kckwk9al3kWNN1qZ57Mx9OqKxBn9GbFgMFou9JKf4
uCKAMMvXL3qHc0LKrO6+9VttNWvvKJtZXZXWrddDG39xNrydSKKnjpYfAT5f/ve4I3hZctd46Yxi
5iHa6+00efZFNpeM+lIDQMcfAuScWTMrUDglX9ChD4FG6YoXuOB7/5mI2fq/dW4E+JpBqfBuNIpP
7rvATEQIC7YOMgF1bvNoVx3WWm15XB55IItvpEhFRLw1ZEys4Hgpz6DE20pBkOnh1h96kQHiwSN9
h60J2SYfp8Jzcu6UXpZnzYjd6fMQ4pB+cT1asGvMFII2u0tHnbOSh/Hsj4QPJgKbyI5JQ9e3J51T
AkwSq/kWtCUCQ7lMmnXzSQzIHVcM+/2INVq3CqjOGwi3JxHBymjuYXKZ8qw/QwifsnrJCkEkut+5
AG1mXoonHUzLKhS4ogVBF+VSEh7SZg7lpWUXYWBfV/VXfguah+/ZEMvtT0ph4DquDay4Dv6gAPhL
BJ1CdGzff5JONtd9d5dLSmCKtwK0xYXL3i/WUHfalGxhcgt67krbbtjeHXTFd2zxE/6t8ZDyokOU
N6e4c1PGmD2qrfrE64MafhC5JHqwTArKdDdbJzLQ2E/IjrwQYkLMpOxX54vNEtCsBu6Qd11sDoKp
e1kY8NTXCCq04oFxYyBwDy9JrnFpw4ho9v3VAy4nzd9krS7D3njSYasWRxM1a3yVRybWMw9usgUn
boANjvKWetaTtEy2G03rc9QmSe2rdg39rU5OuiEdAC7AJEa5e7pnYCm/rykouzD479YDR95D3lqB
5ti0JA2A2QEux+JhSYtQ9glqrDerZ8T7DvN3ojsbLBSruu7Oo+dn8x8u7W4JEPJI6St5jU4V4F8g
8InOniOVcoxR/VqbvYHJ3bn6luRISByGyO3aMqcfSickstDH+d0PSdL9r18us+zvSHWM680Xrfao
WGz+NuoyFDYyh1O5NyzwlOvjAyT8maOKoPYqx2t5mED1UAYrEPO3Oe2RppeAWBKs5et+drpB8edK
tI5Xr2eZ23TdQJPYTj4kmcERJNS4MiZ1ilATfngmxK5HThi+FGe28x7uCF1o9eIglVbK2DzXIAR4
OKUHeXRq5CBoo+RrWWoRih9ShwQ3wQBMCowhgw5BJyb/P57YYtZ8brt+CzICOTpPS4M/OQ2vEI51
4nv2dso/DHIfF7g4YOvdWc0YNHKKNN/VDJqKd1HAO7Kl65zWkq0o8ZqKCrZPXPqUOipK67DIyB8K
JDNGiN0Dz6La26KO67PudIfrhcD3Skj0SOwlRB2kXLeBtz42/pSPNe+wZg2kFResVJVLzYQCx1vj
/YDFki009L3h0L+ipmu6O1ecwa0tL4yg+iCZywuLoDH3b1VIQlirP5KNjSRW/gpACPQycUG5/LcK
bwXsrs9ZDw0wggpA4dwSC1eEX+oMcPKu2EpZ44Q3jPAGrQ/3GJAJUyHZBdCW0naMa0n0gdJxPfYR
4yY0TTXJVq2gNHiJa4ob+m4srCCi8QLgJv+de38FL3vny8uENmJLhaebxd4DhFBR6YgiZlSvflwp
ZocyyK1b8QxlN6Hw0hXwt0uTGdnUdJhWZEGU2GXGnGMpOfJqjBVH2yD2cq2y53GT840Wi88HLxdj
4NuTnfRldAO+3tq4qwbEHqnZH2f6Z/Go+DXOOCDfu/1iF2ED5KwEK0LHciuUpFdceRBEKcH9erFP
TOM35P7tIkCgPv1PR5GIzhE0FLOniv7MSFbOJUgLhlOGp4BU+nW95qgLXUIeCnuPrjlq9ciP/PYq
ZPoIIKpM1X1PoMu/RgS+eVkIc3lMoLHQRwmUf2bQ5bAgWP6Y1mr6eFZ6jM1ZCSW67VVsBb4Ez/Ad
73pbMWT5EnHB3zExYceBjtdKwulEXeCuqr3rMa+5X4OkC7ZZbCWJDJmMj9G24LJq/UBxKQT3Xyli
aTEMztUHB0O9ujHJvhQ8+wVNJcxAhbg0ZqRoCxHtyl2M+F7ZyOMlOo8LfROJGDZHjBowjg7ONzeU
xLCLEaNVUj8wteeFrd2rrEIP4Ubeq8S1p2PQM+Sy1/FX+rMEpajAjl5sCdhzQY2KlN8+f+BzRBmO
O4lJW/YInfNX/qdhaoosp3MJAHR3at0t0D+yLrAVYfTAKbuklcv92fJvd6ItttpU+ji0jL6/9PHk
OM5yVCfGDvw41sP/La3QEEPlD6UkoYKAOzKuKfIhJg9tOzObpRIu/4EOm0nxC38E27KDf3r8P0iY
R/vJVfdO+jpsstAMV/8+XuSKsy+BPDY9+vDUQxIJXXvV1bLOHt8/kGw0xUzGfp8+0w2YXCEU836n
l3U/ifpsqs05KQNjRAjOtdSnnaq9R29WZSV5xli5C9f75Ag01qWuHhOU6khtMjmlQqWeTuploKua
rnmriGqz6s8ptlxR6UtN4uPdYUvGuh/hQ0Xk5bRdXZK/PSuNRzWxw6dSJtXHLJpJ/wfkXoVmr6nB
lve9EW8Rmm4nJA5ahoewi5eP4U5eLV0sDag8y+t/Yy6EWRJIgT4DFwAH9ZWWm+ER1meLUWQFRxuG
PTDBEg6+Sd4I65DJ5bkUSQaaUO7/VauSEmGvKFq6Ete6ZOSxIdLQAr/mtXKNO/H0z6pDipgH+Ms0
L3xDjjCWkj/zzhoGSmdMZMbUZbGAfoAJWXkZP0d78IZbnu0j5qzBBst87eynKmE5GGcNGLB25LXl
SKuN6wiZ4xyMV4f57BOkxFBhQWKQzrmtG3LUNIeXTKrDzPlhiWbyjbqYzssfv7+L8fuZJkGPEtzP
p+e1eP4OPyCc8k8wacQ2KQeUtpIKVwPFdF9liMRdvIsX9kRezxtvKUfP4INELKbFmdDlHtkJ2noh
WlK8xVC3ODS3NSN0oO3eZ9Xn7ACwc3YLsccVuGcSuXhsh4vje6EOVAcVw7lalYKBg95BRaxqbJzk
FmskJNcP0cag7LgOBgH3rH9zPyTKU1wdkKVr8JP63v/gNPAwPFEUR8KI9fTR9h33263nx6XvLy5X
/5UNARF1hftYreKb9mnwz2Rayi7ejdcVDYDkP1GW5s4t1YmvY6sOYfaeQ7SP3qEIXFSBzihkcIch
FTUAUtD8Xrv3kA88KSv3dVpXQIKhpKQTVyLvBn8tdP1IgsAe+QCHkd3JxzKoRFu9r/KWd1vX+KWi
pGaITAHRHJ4HxddGKdALH34jHMbiqBZpyRdGbvhRxwc6zC3jByTJFOg41HziLlpw181YKs/pshg1
b9WzNgL7uHrnVZyI75O20lIRc5HZY1HtghU/BveH2jqQEdLpVzNZWTXlKoIAfBiVjXu9CizQNtbN
9cKzxpQdYGIMAKzadZyGd3xRPnTKjwIx0zm0ucC0ESQr0sC9fdfopzxzw63WyKut5OaXqdbjITNT
iBKlQltfhhStyWGjC/8j/IoN2e4InBt72Ok/UFewom4vt9FvvbIDMYcI88iFl1pl7OfFzelkJrBi
ISMtofu+DnCQele6MXWLEmvCkMYPmOnJ2lD5Nn0fZ1TxRKteC0KywxV5EXQAGZF/n/O0H5wbbQQq
0BTkltqRq8pPrGSO1iEklvUHqtm1ccH3NpRL+OtADCxv3knr6hHYTBQqSLEeeXToU42dARq5DUZY
UZqp//8HFNZQpXThFfIMs/x/lEe1o5Nb3uyUIToBhryE7itE2Zk7tikbjg373Ma/Aw44J66pwAKq
4Pc4dfINKeFPdsTHIM/gv0eXAX+eMDx7yX262yRBAr2CO/rQBWJaX+3xsmAineWHj1+0QSVb0Mvj
pRrFMgCqVyCPViUuQboktIBbFJd4l33M2J42x+6hA465BUciEZYwvpAYRrKvCY+DavrJOArcp8Nt
VoS0q79+zKe2ygiQvjxW2o1iwdnCRipbK+2DsRRoAnKIjAOOZYx/kwOUm5k8DmSo8VOD/o5EuFLQ
q5TGEI99da2ZuTI/jZ01WEvZuvhMEtoiY8SBCbc/W5xByEW5xyfoMSf0MDrnNae7voIBgOK0ueV4
5+BHxkTnJ6kZMH5Oil16Co5SjnkX1uBL3dwtdcHKUF6m67BpxTwSPhnHQiuU+isFlgZgDQxLmtgF
Q/WjqIWqG5EfwbyySY+EsxrJ7975HPeXL70ghbmPNMHFAqQsaYzCzG8M5uGdswnnxe94KGyFjn9Z
OjEtjhOsDTaWPYmBZy/5JNGvaY2hN/e1qW4iHZKRuvj1sqa7iU0rCkzjHAwNQVpFvV3KygC60E/Z
plCEP36OFPCduuuXsfQq+5IBvtvlDjtFBc2vlpZGZOZLQaGTq+ZxUzx3pjuDlTxjXfFiwpC76T6A
jBzOqyTLpUPw5JCBopltn/SxjHaVXs0M4B84Bpp0sGNBR/M7jwEF1fWloJMQ+3jejZuzPSEIYE8s
eo0GCYP70ViSfW+crBo3cY7XuXahd7SpGm7JT0wMm11ysz7/5uHiT5b/YpS0jNd/iRL55wvdQPjl
Pc/6Aqu8JnKK1A1rLED2clNBwx3y8H0+tDgbRlW+k+NbMNykhVqptLAJbVYchJc6ne93Ys/2xMjC
3GV6WcoUDVui5GkmDIJvfLdoliCEmqiIyZbRtOXc6ggcN0HaXXvKI6K1gHCU1ybEnJ7jnHVQeFjt
6ue53Bci7+1oV+Y+YycdFfh5UAN4koig2kERNsaxWgwlaCufGrTupXXqKUOV29GOSOUsERfbGQhy
GJ7f+Bl23yqRX2vG2uEY7bhboH5jM/tRYCASD2fC/F2w48AiUVhHpT0B2kDNkQGgNtAQ8AsQt5u3
X0tLtPQJs2ItjlROxQ/4rSE7SYht0hibwsfafPyBb2kvCrhedPVB3rEEOUWj6W3j8X24ajYgZV+f
NsmvE2P3BKqa79ivmkU1rTXvat/UAcSJ9vvImyNWG9XXMBQ6Bf8pizxw2hHHCZA9vbYY6Ks5ktrb
iSeDdX7mmZuN40UR5z3Qw17L8eWlFKHMn2KDiQAqFd9rbCRcxiR4yvE2zli5F4g89tIR7ixWwip1
QgE9LU9R5zdVdz4vfHDzEwSBIgAbfeEaBiUEMZdHLncCpLFWAF9P+OOfdbFexk1tlH5Dxm2ET4QA
ekj8G22SzzcT3eF66+EQPwIEhjKMIENd40U4OE6tLajzrFQ8EQeF5Acc22bOQuLiSkxfcOwYaT8S
IQPctyK1eMqgwcp7bZOrlN+iEaedCCT69zGmUVSPpNEA45E9yR8+DwJnjvxXVd252EVJCkkVWaM3
NzkcN0PcyIWiDLY9k2966PBm4jUgmIBQMqTqJXvxhVSWNgGzQK5E3d/yHjPS3CrINCO4Up9NqIoL
9qZ9CmZNMc2GNFpaAehB5azj/ntsrxY5tEQL/NpYAdLiDxOxcXvBYiHlh8PjnO2efwIXjucXd3Q/
gOkoFWL+W4Wvwq4C7D+G3R2zJd2YLFxqdFPBxPgwDoP011jMBLM5hjHLIwQfBUggKpt6DUfCj+r1
9mZUtGskQq33l7Rq4PjNOVOS4t8+rIAZzzvUJNfkve2DBFSHqPJBVwAnsurRPDT+9hVYBhoGE/Re
YWxJ2kN8W6ynRJMgYehZOyn6x94i5bXtN+AQpUHFhmBzXvcAmRvmvZ6i6gL4V26L9dxjVKCANayA
EFMmz+OIMH3jZdraec/cd+ThFfQXeuQNQhZFPU8qzhNQplAI0+mZ2nJbxJRvO8OwixdGtCKpuuqE
SSn4hxCprjCcg0y/dBrInqzFcy41fOp//vIRviTJcHVyK5fnM23gYtCUrNnjM43KQJaVvMtjn6KC
XU5a49UfJi5U8GuvVuOi2iKgJ8Csv8ebU39qSKE6S9gtiLHaAjaLuI/2Ud3pL7LylaWfmr+2lIbG
TO3z09bNZ6NPP4nPe/+tyuNRcRcUgr4C5VrLtlBkifD8nvCuO3aD+j7YgiE3IPe4dvbVqFAWNogs
U/3M4sopux98ftzCjIRVXK/WcYf2qwcfgavpUkWsHeP2nnbftx6TZoU0YJLRSAXC0hpLf5vAatQ5
V5egaMGtQIrDzNJrKxGnGGiDK/lu/UYpWO73/XuQ1K5Nwmt9kTVgDc/mPhP+jIWm1/uezz+pMFWx
PVMW//lVh4DCfFIIqdNOMZ2iRsd731JH8U5xD5aDhiDZcgD5zIYBPiayWIvAfpkrFVORf80V/B2S
+Bb+ONKYhYxmWwgOHX8UE/0leJRelf2D1DmDm4+WzK6w7bbZzWMLbk1LEDZCCN4sdRMAmxHtxbEq
b3vX7eg4r8VItVD/8oBuz9sgNRvqhOZ+CY7/na4cNrSQ49k4mdh2MqwrAYrKRIFxT+mSSWUdx4bv
7L7XFDhoOiSgmfRrlGMI5+w68AvT7CqxJghR64wrHLKwok7Kn5dmD3ccoTbKMkN0cZYNFEzrxRA+
cqlox0MSIkLJHuHwUmcz384h+qdQW/dIWT6DcGuAMnIbpod8W2n6DeHdu7kls8E1EcDL69E+4xuC
/kKkNh6pFDR3Sds6j1EKiRQSiAElArfTbyI0SIUJmAMxQgHsUiYUqUq30uuf5Sc54T58VRCTcSy8
CtvtjBi8gMkdE5i7cmhC5tUzUGHRnUf/GwRIZf1GUKHb4T4eUD9+jVJcz3NY7YTu3NnXhRLlD57W
6+uMBfNbp63eClu9h4Ev69B6mb+jCzxgTSXx+cDIND4Q8O7e/xETIHHRKMCwQD75/zEEJg/PUfBo
cDI2/uDMeTnTzj4cn+ioXN+uU+YZN8AHRkN56LOVVndJnldhDGJPvCnKJQPZLntWXIhUTsImSNv0
DlAQKlvGjjVUAuKkybIj9LYV9AgV9lGMFfaHh3HVYE9hqDx1l3jVhv7c29LfhCdDvl0GqFfeoA+5
s9eIUgseybdmjbTkIMs766EFozGFZZtPsFYOH+QH5EYxXguHpVmc/TSanxCRKrto5PUNQAW51/nZ
gZTiop+7tUXqJ47bPE3hRqIjc/23iRCEE63eed0+EQg99KL8MSg51dPb4y8Ly1lzlsvKfOkoXd4G
WOAequpLiTHfDQLEQrXGAAsNhUuj3cArci8EbE7zFo15M5ONyWOZE+sVvsBk71j2sUJyWe+yVohL
ZkpzNUsq4TRIEVciG8NFzqsyypCemIs3OTriCf1DVlIwtuUkfz/5xpi3kFEP/gzS/tnv0ITYIxTJ
mG/OoWaNYI/3A6H6zvBTEIdGZGD0+kuvnXNkeQJd/Ow26Cnr0x6LfGkLIkI5/aT7rxIizLoac1Eq
E0xsT5Yq2xhvlSEqvXmpTghnP/a0tAocqFnDIuDAJnmi51dqdDronlgmw+50H8CeVkVetioIg0EN
Uq/OqHHRZuhLpcl1BY8fKdJKDMRbjnCKS6RBPHiWH5KJyGIIZ3BHLsK6FEhyoMq3ncMDtnKUjwhj
LdiJjdzVXLJ579CNBZwdQkEzhqnE36azwa8RcCArxGNau7vXLRjXVPqLphW6P6dnSeVXEA7Zulqm
oxItTbNvgMIbxWFCV8kDd3ZeZDH8xVn9ZGwP8Zo7yuw6U1WHR+99I1OlBNfAmkCRDxk7hdEiolTD
TZf/q0riq75GO/ctCAA5QL6eRJHxMC+UnHGrQ3T+4AX2RnWaticbT8JSQ8rxkJZHfz/KV3GHGtxp
cEd5St+I5r/V8mFxo8QH9JFmHpXIEVjLCE7cgPQrscgWw83en8ocQUQNqdTbA9Sfz3PDS6grf0en
cGgVvt7wrTH+lLX0JhHoQwfPON8iKyBGs5jQM0UQbNUwZx0/ZtrzUasVNsB/J3jQyMUOXE8AVo5j
bAidjDp0bO5HD7UWab7u1AodJDcvMwbQd0iEktsTb0YJoxmOc7iY0VuVgTZ+LBNFAIJjpEcR0KS5
EUzMISKY1Tmj4MSeXOXBuqNee7i4xy/4OTG+bHwzJqsVbtdDJYpa1nha/mrIgLbanWKmK7Vue7b0
F03cY9JGfmC0r7QiEaOEUNPO1K7myEnCCScUG7mzmi2Fet8WjdpYinwhyOqEqhi13AuOZp36hf2T
uU4i3pMxqQToniip+b+POpXPzWvrJRbWjHl0HXZUUVzoMFNHvKuBNJdxIeUmeNCClAXmSuz7o8dn
G3gJ0x9eHuIAE2DCnehFafP+c+qVdSokew365r6ZLA+uOq1qGcyOoZ+RaW3EMi9kSizEwUyZz04k
LcSG6cTNykmqdQodHNY5SVzIl7ZxTzAQqNBIDMy/l8wzR+02zVxXEP1vJ586TNrD52/VXEq0mI2n
ZAN5veIt9hLtndzMj6i6b7ZkKz/FZgJ8ZqGBe9nz/5W3Z5Li4tguAqO+jhatjmuNl8Z3fKRNgkfM
9PUd5r2okCXVJ+zk/lhFRkEc0xwXWkLlrl92RmqdbimqS1j8EGb0eSfT7/b56ZjjLba8DJBKcqNI
hBkR6oug/2sWvvyJplzOwlwpwRWjVnO3VZKjbWJGFUYjZfW49XCcO5Jai2op0Xgb16KBUpIGaI06
8ZfYyYoqsCS+TLqUDJBpNFKMzNXcz4SkBa1LL5BN0qhO+pb6j2VBC5VzA03zRwTIDYpFL0Xi161k
i33Bb72I0JfUqXxJAWSumJSoDMbkGLH7PgFo7BrrYD8NAFbRNPJAByIXUxnkh9onIExRTkBbcPDn
MlQ2vjFYzxKrmVteyIRgqcARcs5trcbXreMS3l+wcmMHpG8vmD+xCFAjV4Xnaplc6WJ0VNpfi3Ob
XTyvYmVMr5FMyRXtoHK9HuEuFa/q66QhQ+jCZQ6hIVrhwXUJf9DB/92/PUAzhgPEfedUTg7do5Wa
Givlhqb5bchCd4pts1gQ5oAxbQfKJbxzCiz7N0Tko4RrtsyNMVx7TeAr9mKcgEyGp+DAbhT/MkxG
4lmBu40O9iqWGAQuV6Q609Vj17eT0Ue3OOmqdZcIWwJz2HIGrUIihuXUWWrFKDDCIcVnBmLiVYAz
HtjkhZ11RbL6bF87QEoexPMq01UpOtvmRBScS+TIOlXbnXuFczEotN2Tvb1p9HAQxDTUyBaxG7Wr
EqxwD2WqBGFQcij3+EaiZCkl8VqKmNZjOHQSyoEzYutkYXuuupm7favsljRba37YYaXZ9FjFsA2b
kDbviDERCtpF++P2rgA2Q/XnBRwuhUmWDcZOveujFCqkzZmOFu4LsQnFhkJtTAkw9F94O4HqM8nB
8YTXsPdtO9lCoqLuvPFnzM0PoHTtfirpQ3+zPrw/P4h/aa6BIRjFiiGqQkT8JiLWTj928xSj4Im6
axzXS2IfwdoC0Gv5WIZJr73KfwvDVGuI7t0XHKPRnmQQXJOIkFN0/1RMII6C2AZuY3b2KFKJAeVg
GDaykUyPnJoCBI3ZP6EMBUjy3FD0gQm8gbTmKX1kTyoc0wqIBEldr/g5jNvYUG7PLEUgcUWYgE2k
ZDRIATGPTj9JN75XWOwI991Oicsn80DPnTGDzeVlGeMBmPH9Qmelg7mjyg87YsCJZhW1sXzL1SRe
stEw5tze++8aEgaxk7Ke7xO4+vzFVJY6AJj27ZoWwoN8BVlUykFIMWhZI6S76iEXTUKHEjkMx0p7
tVeMOBhQwouvsSOTInNuiYVRM7uUla62VyPAN9nAuUGpLXl+LHCrS1RxStfc/kagMQCyVwCfW4zP
9ySHiHzCtzA5Xu0AvTsVQwyhblSPOpd+7S9bhZUppBCqIKOjggTrvVEVxDIQPU6lricIbtcb6u4A
vyyz+fWGAf67d/RjdAZfu4CDTluiabRvIw55yuzghpaTHm6lHlg7B7o3s/YsE3x9wYyyvFmh+HYo
crJfyB97xE9WsE4xgbuEBeai25zvmTlVNRWTbarTLVOq3YmYap5fSNzi7aJ+cleGqH2yEc4bDMdd
WY0Csmc215TpAgVaY55U4isDVi1dMluLI7H4juM9KgarvLi3Au6j8gFmuvxr/9Vn2wJgJySDCJ/V
e0g7hOvTZFEuMmmwou5BLdVuj25Ccn8LSkU87vpeQ+XUYK0cI2147hc2WhH7b/hZBtsTjkyO5iz/
ObV7FSKdhmkb6ZtyM+hXEyjxI9nhCsmANKMwgHuomqWD+xVrLDhfOysLWZaUomboTtlcidWgcOsC
MyL6ZzF9/dMz9tAuT3z7viw/q2oAm6ozcl/oeWFUvyI+IODmoFJYaq4JQSc3fOLMR0LDM2jNOfL4
QHzHgOikglbZKzXFk9D2es3RdFQDTW++XStv/6GdT+XoZDGLLf8szDpp+PzBY0tFiMUc8TMuEkBH
sxsZPeJiRvKHTXfFbpfdyJUuPo0PZkPs5ZZUPJa5STf2Qj6FJCdn7WK7J0/SSycDbtuisKFB2t39
/5w1bb4phzDvpM9hUgopQUsWxAoKZyqP/9WNdsIb6eZrnw73GR6VGT/iqvxlnDGW9MBrujzl/dPo
OFOieOAk1ly0RLGZUhIZzTsHPKWp6YDgjBXip11XkXkTM25iTPfB8LN2aM8a4va19PN6z7BvsH2q
08vdGiExAfJvvUOBnWBNs7p9izVGv7J/2LO8X6yRUGyZiI9YM8Kp+X9Q2JLYWTILYBQEx+KkNjfD
SGzvUp8tu0WL2ollqqq1wC9OEqEi3+0qWlWVM5BURhtTFbkmf9sB21Zx5d1fCu+6UmoGD0LQzuki
NyfNa+c5XIv5oZJLPGxhlfRbA8cf2b7YDzUhF8NZcArzKDHSiBWGKxCwkG7q/SR80nY571XOSOSp
bxAiHhV47j/Je3/j+dicGqFwAACAS7cxkhiCGW7++pLTUNw+k788AGxE8F2VL6AEp2Jb2KmYZt1o
Rz0726e32cEwWA6eHkxWsmUxkuIHF7Qwkn+td1lJ9PdQ90yVWac5E3i4sgFsV6iEIrvXyA3W61sy
y4GVVcJU0R1FQtI7E2yKxddHZwJgrEokjDuwPvGh6UWoj2FugYP3hmTrlylQNR1ae+d9/92X9mug
pm0wzuqb1O0AN7h6E9MGzrSBm8VNvUsN1L5mc6lY4sOcv7MXywkpzwD5scvpiaTmnyMlWVZRpidG
FKHiqDvBVDS0967QtCj6F2tLy793eATHR6UsgCyyt4w/mTx2MyUhMhz81YuTzNpnwd8H5rfhxU5k
C5NW1uCjJLZVJzAci0cvhL3xFXA6ODxah3xH4cpxZRj8YyDri5uAI9ZRSbrau4sI6zIdrC7EC+KM
3EQn5Dd1SxdrnYs6i5rdSM3vB9MaCZXwm8RZlstrwHvMvw59yhi0pUheC+rO+WE1MlU64aWtt7nB
5oB37mV5STvrtDgv0WU4WETfY1OV2iechxxAsqUVt5cc1PeOXS1trjOQ6KNZLdDU+uBwdW54KsKn
c0ANpjzAxbpiXYlBoRHYzKabp/po/9dHAUZRIbPCqu3aE8eUQyZ2jOKCosCpXq6cUwjuEEglTc8+
aKsTcNnzAJB88gT3rg5Ddh4Yz07XrMECOl5Af0C61yVhaDOMv68/Hnvh1LEL5YBZV+BLO3ATwQK0
rzi8fFkIhWKs5tCd18euuU1kAJlOrl+y1c58suxqriwfrAU0my9p+UM5TrH+BlS37gqNRd3OBDev
OnKkrAdZLHVvBjpITOzBxGVPD6fT+0iMR7NDxI9BzsSg2/eTLB3jwI6E+2ae6lSbMI5q8ZvgapE+
sV/d8KPzym7wv698MzxjoFE1vQo/VQoH4tROAk3PX3EENyHN8cH6Lvp64Rm5rxbUGm/3ghrBqOIX
k/7DSBSeo03tHLg4Z9I/ZWwIFfB4w7K+MXZEkTK81V6PMFKJAoVIVIfQhTF0NwpxQeSRinA4AIyD
Y1hBYM+sRVmpe9fzMGSiIhRwGBqcDtlD/Oe3/Jj1Ru7gOTrIHug9R2aeWU3cwAxpJUZ3CfV15WCd
ZNnRaeFMWJc9aM9XfvOJgCuVuW5E3Ssww2VC77kKI6AqB++yDv0dbURlKDh37Yy3iwyZ+shZQ4Pr
hKLD8j6cF+L7O7R1XBm8PC+DdcndEIFhs30zBsLvuRQ1Y82N3fFD6oU44Vh+hXOADQUK2ZdAWdRd
LW7OFUr9X8T/L/qUE5QaUV7WnevYtzDYm9N5dwdDKvKUaECKDK/yjgxxZ7iTbtrELSFI3QrmN86k
F5IRNljwM8IxbEYKJrUwjXH4prODbhNJVlIpfAgI5KW1M/olML5I4jsX5QdmmKbplAvzfwkLetEp
najfzPovY2F43aI6sMvpIW5H5Fx00S19CQMqEJBCiiYCVSFN8q61e1uYdXzoj5mnqeg4S+v5jqYc
DxCjbWT6Jm4e1WCCbBHTj4t1h6XkiYJCjXtIuv9FqI94iFHBC0SJUpJF22hwME4CxNC0pFNpOwCF
v829RJ/59wNwK0RAYKC1ELlIIXQADaxLzwxQncVzBmOpwllvbK8AYIVbbaYESbdydodJwD2b4NnR
M8tcjaVpZdhlOcyQ7mlDnau1B3N5f0Nxbti3Vo3OcFJxL27A/Vmp1noW1FYzvGfd/4i7I7i0QkXj
hGA3FuVkCLrs+Nd5CY0HCySJ/8YlKX0T5zep+NXeQMzDkDPltp49hiHj8v/NePjpgxRS+XmN5+Z5
EsUPNfQf0GT0mNGMHks3bllrzXHd/f2xJL+KToWjpIp/AZKSkSid6XRMQp4cJ/4DInc0fK/TAZug
d+W2KsICmNOujbU2CMNSC8WVNk08/WJkqtrEeGwgJ1S6i6vTVhdH89PzmDagIt9vsKGEPUd7qK+o
JKd+Fc0S5z8H1ncL4Z0jULUjJKzX+VNG/ZOqfQkCxPZ22RFFf50LgE8Ryu5b2+Hk1G3UfQLyHxIk
heY6dRLCLo+uHw1kMxDJ0PDPaVvUkBf4KRqTbMSU2tamUffU706imRZ4kq4BAYd+eHCEpdNhhltv
boYe4LAyfbQyppKkW3VALdeH1hWIVLkr9W9V4Zg+VJr7OBiBiLi+Z9ItUOLk6+lVLyPe0wJQV9Ao
CWA1PfLc+BHdZqOdfEd0dufK1zuKVHveP53XUze2y29SpGFKZ0pDky5J0rIu6md81FJ9tg9fyVAG
SAudDAnHh9Y3IFqxzMQBGPkBRFs2CJfXsLaIufpyWdUdhAsx3eyIzyzVD/pKL4WAPsMK2SDOPEOO
kKBtYTEjmiRDnWFF7BaNiYp4YChZt0be9G640olLZ+TJqnMSsmrleVVT2J5p6NuEU3CNhr0VZa/Y
4FnRz0PeCQ8gIWYoj5tOGbvUMcLnCiVzvFC7Rfd+UUzt9txtnpz5debHDZCTBcJAJC4sDYtTfZq4
GpsX0TQln8EDwa5n2oj3Gs4ru956ZhNyevNc7q+leUONeWqacC4JTQ7GRKZomIExC2T3uaZKrNiM
1xXLiOLkvBVTgvHbeeucx2BiUg89fx0J4FMOMqJSmx2uGF9Z3qA7juBzGGDE4UE5EovhZUtpOtc7
u7juTEKLKvOQCupL06jh3eGCD0WsuwxlmTwFvs1Z6a07R2ae8JP5qrsCvUiclVFqfnQOGpGKp7k/
m/yCYzugGUNexzzG3B7tIQXGHTN6SWE1eDztU7OXXqHDRgcdktL/zfeQqg5XCFKFjJo0RmB0wdeQ
40a1kEZzuqBGs78x1RFVPAmnbE+HRFv5Qf0PPTiwS/q7OPkKskmu9rd1tcCrOqsocpJbesginKEI
38Qonw4qG/NxCRiWjoQb+YzhfxTETdTw5TgP0P7+ZuSWOdJ7po2iMwbUS6vpC6Hm1x+VI5bU78YJ
KKst/+n4hKhxh9JqLcwIRqwksfunJsAHQy6NpBMsVAvUjUY/dlz4F0O3TpHZDYZJNjsAdrl9tf8j
HfVn9pBQh99SQ/qaBDGunJExfh6UXmaaOxPom6kiniOhf+jWqe32Yrh0Wpwjl+t4E2CsHQV2MrMq
69+kvJvTDIXKjdShBnjGfie0TixX1xEYezPLXrpcYT/uIaq2SqInorZd7lT2dbSAex3JacGl8521
fjiwHQhyGRegj+rK5IehGVI8rTyKVZHK9FlhDQReAHw4ploKN3hcQgMciapnloUVpnQQgwv9NAel
RgRKh8gbckiEw8AV/N/tFIk5n9H+ImOYiEV8u95ZpNJ7SHm2s/O7LOdLmX/ZJokKIDWPHPdd5Ej9
MXF00hySLyXK7WDaa5cwcwjo1MA+0O40m6v5QQjICTqYng/6jckb5RTWVUqr4E6HKw06lSVh0Ryt
q+lYocGOodSFg6Z3NYgITJzUFwDDqIu/ylNaU0DQBwgTjDbqKdjxjmA/908T6m9hQYeJrAILca1j
se87ktT9CUb5BARAUoLUmGW+eXhvIHnWIM2IzSnU4EhGmpLQsvKRRvahdBu02y4LDugOBH979Edt
Nrs8u8Wf3AwTUCtC0wxTYcNhLc9rsgIwF72/rlxuwsBgAm8FxGwNsCclp5DELvuAlH2Otl6r4DbG
axCy8vYX6itgrBaiqeosyzqWb4pjsszp127k7VY+8n1XZ14NssAx6eF9jnUUf5kLbpdg24Ppa+Bt
4GV4fB+MyB6xE2mQPeOsuWN+Rh+Va/F1hNDZ8H1oU+EtoDQFj8HPHnqIreT49R7+0xuedWdOsaSU
gogw+LRo4q86OYGxIUOr+9EFH1LKgJAgSJ/F9f8p1YsPmeniivzEcYTeF+sG3Yhi8Uqm33+KZNLa
QLXK1YRp/gBUFoHSJU5AeTMeu/E+wpxC7yL4Y3Bd2EbZ1cPDCMDgjCFVl4QBE+8DkJ1DOeHFB7mE
8qncGLk9jyBy7L2MQE1Dq2NB89N4tzojLploJ8KvahceRQG+Vxs4RbtlM4e18d2wj1BaS79u/SU6
Bqx4BH4XHnltZvbRGnC97rj7i0eVwPqpGI1VpZkyEnzsqhzoQAsLOOEJ+Hel/7WtjyjHyTFInVdM
kTRyhngxMdLzbDJ8FW4sGLkjYIYcsa75++v9uwfxi2dKZCpmeS3zkbGJFxAqvg4nvEtQUdEty8oN
HCWfgPZAaA86TrZVqLEOwktaMmYo3n78zwJdXUc2tnupG1cm/zE9hpJw0t7pOCsI1sNHDKvElaJL
KbLnClG6zwepoG4ESky0F+cEUaIisBAMxNbTxe3Rnq6Q9gkwYtwYyIsE4/qhOc71YjY682RjiD3b
QHyT205hLD0GEqnZJIKXSjBk6GWT6vLmJKzaUGUwEDWSu97Ugk0N8R4GrmBMoy6r0zbhz6kcOSnt
O3toXatrzrVbfxCTpPXBALKlMdMbx860thPUehZHNwTDTCj9aaa+OddBdL94IGF5c/x42mdJMwG/
d099dDlSH3Jjd6kgkhMDGwsW5Py91ba5hkD4FPywerVqQWEsHodhplQnZwS/MIL2ksbf2/FqHlyp
XlADXy8oh0F/TMs0Z4dnXwYTKBryzgEOybPYn/xtkV8vPVNZ0+mbtNtRr489QNwQIKYmhgoEHrxA
+8vhhWFaGEpitFfv0ZlwFfwE2eAjT6RaFr5MEQGAjgGlo+6pIPj6QPZxDDHeqpPFcs4jelsL665o
Kgx7F1rrKYcR12dGJbh7V1DIY0U0UuFyrTgTWVvYXowTli/BNlGkqkQGM/b1v6SSF1nJR3IHJWqI
6+8lj4ZxpJwu4QAK1AqNQoS0jgWERj5RTQHOkbysT3l6aHJmKNoAEO04D3l7U0oz3Lf7dsWYsEUO
8/Kbb7tH9MftZVra3rOmwBq+JFTX58wuY5tIScP633kcTSO4HaSt6NcvFlZ9buUyhWRmqVHGI3/2
7U1NSUqZGTCFgVsOtjHDhkLffm14u+SqpUzcprQrRSkEGxFeMCui2oX8vpZchDedNajdDwiNU34w
lad1UIK9MuFmreWM8o49GhNKnjrkEaWq1+HoXr/GaR4VwYd7UKCkG64hOK8D2hIKPAP9tDGsBC75
AXLi8fEhC+7yjQKbjjKKOQIv/VCR9r8VFMyRja/WvBp1uaq1i0zJ+Q0+GjroQC0YjSDZ5/vBTucy
8vDtk3eKivEhLxHge0Ce+v6545mSW1AqJx0ctwRt4/ELwjxajE/WNfnIXwyEP02VFFbYlh6H5iKN
lcfEAMAYwMuPAduiGIWUm3HExRY5Uhk4plT1cAsdj6Wvf58RVdu4cVP9h0lZLu/46EDC+TB0Rf46
fQ/i6UE99frHx6zNnYfpQkvX3w0b10IzdgMXVhvHZyiTbCdHRCREEKxqxFloYBLjwV8Chg8rINu0
EAx8Wy+xWCDGnd9s5yFvBSmcDUNulrAHUiZsaMSI1xAuZxLpv4Ipwsd8RJP9My77AXGBBG9ySzgj
zEZ8FGlV6QhRSBmBQsGQgACW7P8WmEBkWuLcQn+8WehGtKpkb4J9rjQ+969XgiuY0j/9IQbRPgFo
XDMB4rZM+Zr99RxRyrMmlg52lm/ITIzppH5szOyY8wPs7J92xJOBgaUx7V8BpA9h9Iqbkw0fdMM0
hsrygFF1/4yMod00ugoSEbUvcD//3/I6PjLa+SQQG0JvCWcyovM765J5j4SmYLF9LMb+5JnJeOKr
LBx1Cf/9OKuAsyGJhJp+u2IXMmyf5KAtiBtKXJucu5ZoY9pzM+ecQ0k3J1s3vNOd0yY9Jd6m01H+
84RqGG28wWMiu1dnXs4IoeJeuWJxhVfadTvZUi9X9uYe64mjitYg16E1I/OQVsxDNDPTFPanKeej
LI45uhRNTVBMZX8vNYCIGWJYDs6ctk2ZU7nOW3pG4M3OMRisql2PJFwIC3/8EK1bEai4UwT09J7j
+1+7IK57ukHXGMCAvQCB/M+qJcyCltl7GFuX1gF+m0N0SZe9ByrvwCl1Y4mU0EDwaJUuWp7PlS3w
rkrB8K7HqZsgFl3XerzJTrVdP4WnfJdTbooGD2jPZsbJSbzqR3THTOt37i9h887Pr9sUZIjTbyuu
V4lAvK38NcTp+FCwwdQMQFm/nam73p7n+cGJ1UnGHrLBaF/t3ZIXpjrwyEXDSNFaYQo/BbcdO+xg
gPhO+r8rJqr3ut65KqhgTpR6jX/M/2HzBDHVzncq7kI1PcS2B2ccJN0gF5CgZeFes39Nq+Jt9Bbx
XKnffVCvlh5iGfVr8+CYEWsU1waJVS62uftqM+RupFVIIb9szH1d9kiCTeFev2jIDhawL9n8tiK2
M11+QMQw8mddd6ne+IBJ+If1axAYyOewaA5kIoHo1WZj6uJ0wgYiXAf0c83UkH4EcOiffsEGzE0Z
Rrru0FU/3tXtPmTMVHnPKg6irNiXhg5Ooeuochv4XuODU3hL/N5WP59hTxeUYcvbsa7kI7GJVDdd
bjK/KkEFI8ps9V9v+gIyfbFwk8QFIeb7BAg9ixJCFiU0+lanmuQG5nL+8v3viG5GeodTcdgVZV6Q
7EPQIFK0NBTWjG1iaKWxdpRpsKnRajDt99/cSQMQD0ZPcJeO2c+0nHGCUl20t0uN3tsVA45yS8xs
T/ZOoM8p18Kxc1rgqJzdrXnQk1SOh+cejObVmxwjrWl+mYaVaCoP+xi4g8wCJfCTf+CXfdOQa1gO
ZMlmUq5XdWfYzZVtvqmAcc+o5A4HX5DHYPDvlRAKPLvL1EsOlq33mLN6rC1Kg48M/JYQnfPxQeBe
BWmgAXA+7zAoVTuaUbHbwpoGnfzNcmBUF4pj35PwbLsZ/1yVMnGLz0xrrtmwnF3o0MoZx1YlWVu9
0N9/lW82kI/h9BCUhlG+KvFnydXBkoppl/kCOCcKzFc8/zP7Xf0L6zCTyO42XC0VQ41a3SNBFus5
5k3cNgEAsBh5y8BMVabf3woFySIA6CFKWkZl71Y36ni7Q52aR87rjV0a8aQs1cMKOqs2Px6GduS5
H4r5Ovuhy5W4vKv9JAfNDupm1o3nwKlYVSgk2ulZ8Yb3bvElbXIbdcuSQHckrp9M0BS5O6YhUTdH
GNRef+PSDzNUSlcLpDPkGC7/hND6fBeax9sEWmnwkVa9R40OXO6uqQ3zV/o6TtSMcRE0rawC28y0
g9TjtgSYv/RWiyoHuUMp5zl5C4CjCTeJbKxpQeb+HArW+KMkBjC6xrkUzN1dFmj9J/u+xMGzZKYW
cGVgUNvfb9OlmVa11PIN49nqiuD8kQnB4Xlw4rixljliBCBcVZpk6ZiyAt47BtTNFUKqVVINv0X9
yxoKi/4unws/daNh0sQ5AfWjIk46PjuxZRdrpwZlPmXJ8ePiJLKBRX/b7at4/C3cOPqcyoEo43Yb
R+r8QxgdQABVdphaQh+/XWLj607ZeyugnYeM/nVjczZjO123H093QzZ5H41P5nI5286WMEKqUmNx
zbwmYe/R6aNLMjguHLFMWjL97XgZyZhTJfuhLhj5jqYWuAnBA/JB881m+f7zs+k1oFMkJe0vZPi7
dqMqWTu2uASIpUzSr8dSW5aaAHv2pvxUYJ/+AaHDpIqiURHKjZPY03Wok+/Gziexmy9qCOWGABZ9
ZEEoJ6jAUb7o2+imr3XkC0/AAJxZMb41p46Jn09VrOe1xQfVbhg3+FxdxyhqBrE7iMdQH/zvwuhW
tCB452GK8fjhAeXQWHrud0XZ83oi0jtho9ieJwgus21PeEyQTt7GexKyp7KuWJ2Vk4wbjtIJFejC
t1R3EvVJ97Ul8w7khCwmDv2zET52qbZBe9BPgQofmMMR61my30d9l5WNtWYhDk4aqthWTDllxM+N
RrSoCFyb0ozyhZY92+N5kbF3TS+NW+WEVBzlgnW8+Kqd3Yf/fu2aE0iYDM7IaVuIJzpZm0bbYoQ7
5wRgJIuMIO6DWX2f6qc07MXeojMNfedGatO1AHDfj4a9Ng6wXdnoNNcnBjQoLhYuisCe09RojOth
B7Sdzi3KAJ/moMAupA6wuCneafR3HyoUNmWr9p9K3Mv6Mwdqcxd/3TvjjMOvsaBjOk+vr7HYUO50
a6J3/VOvS+xKa7tV6H0ve3CCvgyeMM41w7g0dONP+knQE/oaZC7AOLQsR5nc8Chp/V+TTDZsyiRX
kMR93glPogyySiJhOVoZKPTp5griu6YsDmVFVjmiP3LMw3r3ecSmWnJnYbnICy6qy21k9SqBL3MW
61PN3fjLCgC2UKsVFmdVhPX0pB5wFdHu/MiElfV93ii94jx+LhkpG88isIOe0Dk3Yp/Vc1uOBgM9
k22g8OGsVupZoJPSMFDB72+0O+UisA2xDHR6XGfmMdzp7sDpsoyHOqBeiSaWNtBV/mRc5gYruOlD
gmbri91S1fsT5BubxXP1ZI2OOZVgd1rSVrjlTfbCbJ2alLoJ5Eg71gtg2aZWPYQPatt4yJ/K+WXa
1JUY3+EbcNYfSwykSLpPT9HB3qP1bd0/A+p/jBYMPwDlUvFkfil8FID9N9JVh0XTneHtOFqPtDE5
3Lb0uZsJ9T8MvVv4o9V1+7ef41plDZxCni32Liy9AKG50oFmQI1i3OrHw9IDcddVC8+ohIdrVax8
PtJtMwyk1uzfFUS6sd8O4ZE9yuwAMiS1UVfodEEdritS59k50ACUPBQfvN6nw3wn1z4ojJyR850e
fq98ytphlbXrNU6T7YdM035ak13/2pU+E7/Pxtz3gTU/XbFIxeWpFkrW5NHwA2JCRSQC0iWI/Zbq
/zrw7aPmxI60X6QLJyllYso1RGMc0kwf1bUNAA8HhXAvRK6L9OJ9ImzSAVhgr7yAJrea0m+2buTe
qs4AedSJt7/ZA4yCctPb8DJWt/ElRNtrYGBFyE9bGWD0S+4aw9uk7rH7i9CMyx7wePazxb561Wdw
Uk0ctEbOlnRXDUClwAA45WRXCgztd3A5MNNNhMVFF4eR2ZCK6SSRaxE2ciibPbTn+h9H/77aoz9K
/ngzJsPtns2LxxbPot0HhEu+v1y2jtnxGDDN7RCixN8cCoCN52ODU6dfzK0128p4ILHISgqXocJ7
OIlMq/pcLTV1YAuzkDlWNpG2cKWINJBewhnjJJabYecz+bPlT26mm/PesUdrRET1425nOeMkmZ5B
K4llLRSXTsGU5ZlV9WEsbeg3ECS7zc+RuRvzJjhqNGBhVVyqeSv+FgEVRo/jJ6SRAnxOyeZ2Xa/J
yERRN5IkBl5AguRsV5oqpq+bXGPzAFFxxkAIqSIRW+UpHH4nGaSPnV+dPaylerRhEugES4AWil/3
wxpWSXb/quaH0a1EKRxx96upODfV/OvzX+r52FfZIbLNBfR9UV7zmqk1gcyCEpK25oOrhx6afDGf
c1ggnsVsxwFbv4R8P9aDwCQxeY2Ab9mKHWDUdixHumIpXe3z74niRTIvxYVWUBDgDqfm+PR3kbF8
RltXBkGsQHsIrYrOiTGTOOvzAjHGJ9xXZiqZSSn/TUqkMyCzQ3JlPQvJb85nCOExhMPVQvJoLr7i
4Gr/cASqECUQFT+HkxycdhmOcaQPn/e9TuEAXJyERcfdOePz1JBf6ZF6fJVXsX5nY7ric948nGb6
oYjTjjIGsPd8ii50GVSmiD86BG91M4VnDsrzmwgo2hej8X+t8sQ33nekf6ZXw6GeSyc6pgmyp1NW
MFBuyvXXqZAVf2H8T+1tnQWK02Nck2SIVfPHxJkkB2Ux6fNXYgC1nlAHA/0JAfFmoAzvPks6NREb
60+828XNuyy+0mUKSh7IEVrSyBhP9Vns0L1PRF3jQMetgZ3IUG7g9laAUw4vSTlenpPovq+UhjBg
kjaGbh+6dBIZ3XQmq4g+nKawPHIDbkLwVRVO1svaPwcNcYBFYqzGZ2T69LlrpEiQxVyalJRGgCkn
MUe7/9AB7WBIj8ceczrq8Jf/ojduLkOAcYqlhUSuOJkvRr5Du1BJj7HDiJ3x7hyaYu8UOh+MR61U
s/VHZ7H7XsUOKkYHjtUe5xVcSTxT6Ix0FwrDkXoprinu+hRrTwBZydB1jP9gJacF35gBy7ihSA7q
zf2arnn0MOY+LDeCGH25D2n2ivPxekAWCSRE8YZ2tpvd5Gzt1q08ODLe0C//0oHwR159IJ/VTMEN
BcebU6ovH/Lip6jPy0pHh2qDgI7O7q3ApNrjfejd8/EvHxjjpgiYFQCN00GRiEopOWvIn8I75FTf
LQN2V261VnMXI95UghE7tADD7NH9p5huGTkKfwoHCS3W3imQqaba6e+RLeA5KSPAS88XWx/SktYc
ycsBYR1JBWedycMKQ42Gy67sL8Qic3u3cWgQEKBmu2aB/yDXmYstVK8X0b8Qxe4pcUVd46UXVFUw
CPuphbKCRCpGOkqACZQZcwBrdJCsJGawAwKCgVOGujdRqiP+wPq0fSk6PkMaIpOizzZMsUGrPmP0
FwP+HNXEQFu/uPlS5ZddX+jqpO9d0hKo4Zuyz09LA/BkiHSkMXZyA59sbbv3D6AxiytpLG4bI4AD
vDIXKjNWOy5W1U3vMpT7ejbm4CzCjnsvhCOJ5bFDyHLWsBMXLD7BmgvF+KYySlb031yH+b3tYtN+
ESVKTRElYLqp9uAykLlcM0ggoqgr16w4xFpFgqVkx7IRgymDiI4/as9mNVSMz3jhQaCjF6K80xtM
+/x+4xeMAXyzF22FDTP4nCdKAjXt3Bm989PUF+JGEI9ZBx8K0MXEKn815AU1sbrPZjtmLwV2nc6R
l3jSn4DseR6vPskmql9SFuds1LxDyynEwtRwjJ8q8xNlIT/kDJRao3sr6jGqU+uV+fM89pIDiO22
Vuq4ZPssWxxGqW0eWuqyd3exdB9qrWTjfw4IKq3K253NAfxA8mIMwvm4BBRa7aq3OcSpg14uy58e
f6hawqWu2qpsy5fwfNAWAYYZMwbLBfuErogyvh0uswdXyNdN9ex2Wl8PKiJTTJzbowZfT+1wwBGz
wvE5k7+oOG53wCvwcELMd7okVB4GAUGDn2xLplrI863utj4rwvQbobE46iUDmSSbzFKy3Ft8bEGd
QXTH4KrLg0HzzvFcf2qQ8EdsOpaa7crk22QDpLcAjtn/Ep3S54JpdGOfWBok3K5iyFOuCItyWFs2
Eg8fvJxk/IS6RB2zdyUjabmyODglznSycvCqfDJm3yqqRG1TlBHngM16DEE3TGjujumyFzGsNpnu
ZV1//FrGcxooALzsdxntPojxrK6laoYx6VkzpnxdR3RZ2nsMiCrtoK2GIshWWElwmvjo0q7P26ql
SqCudUoZVa53vYiFuPVCMFMSwU95HC2GC37sChxrWLmaa2qwGM3CxG1iqNDo5T1XgpsXOlqraQt8
SwFA/TB50PymNUTG8QtVNLG+rP/ekzvJ+ulJYnUNGlgHwpwuav6O3PdyZRyHtWKXrLYN1UiwNvfM
IX7WrSE8MhOl2w9A26vK6RwCkEK3SmZGKbr/ric6c+DhXNIeUsnWssPCeemhr/3dm7qMPSgBHApX
LFtr/TIowyaqgE51HLJ09UQA45GKyKrU0i3ywOd+7Oplhd6p6uwBXw8yQzuyMuT+FB0kdvYukHDb
Jt6/rhIg83FtIyvMttpjI1KTsbHI0DXqW70bWujhw9hhu9Ax+BEw1zABvumhvcs2ULIrZsfPe1zC
LIQXFQtY7+sMFUIryVL7qSE6DMt5yiL3QS+e7RNfh0fV7Uh/sOHUVg1zywkVKxmjZpZDnmoXUyad
XefIomGcr1ePnd8kqFFrrESCM4CyJz6zrskj0e8bbPDb8hfkiauFLvosdiKrXVlM7pqZqiELbe0s
9gFxznrOAMVtZicKkCkO47XLKbOxBKtfPL2qQa5cQOxCKuIkXvPT7qNpWn2TGxyvcv2z1mmKK94a
zY2hlmtsweq9/walHSRDB970UOR2uTe7NSseuIq5JsApv//sTqzTna/yv9f+MfudoAf1ufLLjQzv
FbrV/7P4gwIOO0HWIL3ZsWbC1bjCLjNYcw+OD5L/AE21Nn0i/4FwOOFjBuUZAXzlCTz6EX1K1KHp
RwI/H91TxuZI0g6g8mBCG6SVs8iaSlIXOWFzlXJDJHTwsy1oMoBqxb1icarpdWUFCEJ3IiflyXm2
rIpC1IBUDgQi7BX/PKyHAUnQQSRXfIB+tudow3nDxXkE4tYakTRzKEJI2lCJjTQvlxxzWgGk6D+P
EOehdiny12ajdK9QWks9BWE0JSAycIIkSH74xa6g4IPhDDdiPVrqfD5NEPJG7FaDWk5SfjjScO6Q
3/NQDP/+ew3fLoJiaLZRcm4mzepr9SQ2pGUzANIpkYfK8ixSUDLvT22Xbkq1YOIAUV0SgQ7UKso4
oLpLD+/WENGmM3gttklb9/+uioiMs49HgLeQPxfC863Lg6pA+cOGJDrQCMpl7t6CdOHFB0hEAnyx
bKjzA266J3kTPrna5sDFKIEfwHsagl7FR7VATPZUZn38Uoz/TPYfUkwiM1/JU8+nJqsDo+DvRtIm
N4LYob9/79/fm3oiqlRzd5d7QFUrQXRce7zgn7AteJxVX/KT5NcJavoU1pvBf8p7Yjy8HYMQjE4L
T0Ww2ReSlY5eLzDjfp0JyNrbPhADqR69kFbuSLo6YxKmoGs5sQ+he00BAN7HxgAs/aFhHxW5BZFz
uqNVqHjLpv5UE//JlKQ5d5dlgLKQbft+GrSiHzUaNqKDU7v5qmuWSCXW3Kdz4TgI1KajTdMNByHy
P4eXALfevk3XPEcO4chNuNL0l4imXMu2Th/4vcnyynzsetUKHBZte5qvXb1JZb8P6tL0csTie1Ag
MiERW6joFWaUs19VxN0jYV26Y+w4Z2/dxuBKtkT46D0DmNpWY2EhSchAsHyT1O92C1Yz2Llk1Dk0
yZhv6QkRX2UAX23/rmPwzZFFSG4X08qiBJry8JYmI+LK7ltAdFord6oJ3aTjMSzPZ1F+BJwOOWFT
JMrnRIE6l4xvELnsNZa4AJqJqwLRZ+E5Gnb2liaGbcHtW9/bjpY7vesgRgKwT6Ys3PSwKk3hpUN1
z7H1UwDBftI+unM1H2h8Pyj3Opo17gAn54t7S27Du2K92EG2FE64K3+HPNVrhC5pREvGLY/9Uap7
RYRRpGUPXHFDTQojanGgveXGLDH5yeBw8YSJH9rBZRWHEpuvQ/PRCC+rQPZc96UoU7p/sDjlWIh5
oSFM6Ngl78KWdJHJSMrbdmHWb5TG/l4A30PJqscM66yAVi8/eMIfsGOwh8FgwpiYfCwLAK4Rbepi
HE9bDg/iY1zQ0PJAAwg+Lqwg/zQxPTGXvb46vLOqAmkkKxXuxN1BG/0QJnKXjMGKzp4X8FxAj7ON
41Mi8TaQOuuM5xgrvGLaouXLFj0gogNU7e1TYfNHFWj1DUX51rdz21DLE0uI8qiMUHsqgahWRTla
88yRV2AYp+HZDUQ0fVA7vkKwa16KWyvzTYJf5F/OI2W3htKUvd5rFViPLFLKIutZEdi1cSurj5Si
U2UWP2iGaEcHu9P2Mk7pB/mFLX6SQ9CchKaKVuxc8C+F3X+DhFqQATeV1pHzVssVuxhjeZMW6P7U
LnZ/H+gicijBPV4LMnz3+JFCdmwM5fdNXFyodppPlyUfTYZm7s6iW/a6zI2WmfrgDW8ZHgDJPtMz
jEqGapCd1oxSoqQgLOIJiHPwzk98pY0YJvDQJmcHxFQttmvhSdk/uiA7CeQ5+al69uFI9L9M7zIR
MU2cLX4K7Mp2LwxQmTbilkZdIEJ9x3zmiBJY7QGkS4+yk2BcBSpqNE6No+/ajd63EatVsfYUSUKU
ugcRc4Hq+kCdHwd7MP9ijt9p+RPDYG7aPyTFpeUVN8joEan1+f+FLcMC+04m8CsUynl1LhwTLs0z
n0o/UuWaf8GrT1JxHDPr2dVRJK6xK7PidYaDj2S5LgZCHlUWndzDORcT0tM1Xqe4pd47Upx04PPn
C+5yl+KdbG+GasY2+Di4O/HvYYNfPfWjEilvIu5jnVmRxe3yZ+n5+yv7PyxeXiuUh17z3TjXvKxs
0WM7y7au86PknFCjdccLbh0Sz9VzmBho6hQKN+YzCxpKhttM5So6bPor8+KUfjgg0hs/ECd0PYl0
ZFtPtrfcodzW1CXcJZ7K3JDzBFJBiaEHUI3lnMJZpz/PivVdHYKS5bHJCC7he3Ud3bHQB1yMRMM6
zVjy0hdTtsEEd1PSYmfUKe9qVowPdxrIf/8nYgVhsYCNhOGiNMfPKXB5uaKmnnqHgg8QyHIkg/cb
xBbdAJaP05xmpplU4cwlFN0ED82MidE7pDLRDnVYbbKG6+yUAhy0RbAeEkBTsbnCIZ44w3vj4rpx
zQU19Ro3NuxCuxNwrFLHuoAd7ZyKziJlAn5ym2f6ts+cQ1LVx0Tfyikia12gsul7W7ebOVKGTYFX
mPL0DEyMo5KDZevS+tkpQJQvezmWSGoZkDP4HPINRGzXLdAN57C7ZRH38y5/leJnhL/UCZc8/utE
D/dscQ90/fUBlmSTGMNplwwBAeiD7cIG3CF6L1PtIunHTm2UVvLDPzc1AW8Opcysv7Wl8NaMoVzI
O00EvE3mQjIMKo0Wxy7glP4pniJXfzgd7EnXNrIvr17ZZ1Lh/cus724y7EQV3PZsNxyGSQKfAE9N
AJ8v1jSkAsEmsTDU8ijXOSbSHjpXvdpSDigiAgawfxJVTx0ywOxJ7XjcT1acS6JoftHC4QZE4Y0U
/5808MfkS6von5NmigcoC5fz8oUy15lJkBMIZUtCfBrtWCNeE5HR8Ivtc80qswTm9ELH5yPCaaTh
aNakdMr05aeqclvMeOgp/6ENioge9b0zDcjTM0RNHWfEm2+UoFHnyQfSXuQOCOd9eLHaopRq0PVG
BO/eFPay1jXiX69KXAe0ybx0Mh1P88f6QVDAp3urfmGGDMzuRe1hv20JY5DGu9Ib0jIyTqvqgnEH
v0SCxRcbxMgiCgW0N4xX0m4Rq8prSY/+h8EG6Pd7rduvUy4OioRvUQhhqhno/e1vL2wG4MD8awTu
koAdv8qlXxqIVHEnkpx9jYN3YkPCXWaW5plb71IpnRWQLOG1TMGkiEEH9doRFhrK58lKyh0kr1Cc
xzx+6W8Rw0/mxCLxam2DRHYsFwjQeyftb+bQKZZ+2iidfHv7V8birl4LSq0W5dpvmM6fJofbn/qc
MvQVNUdk9RpjqCFwIrBgqPRUBCbJZ/oD/EcCN2OutLEH1ydh8exd9p3MrQeU5fklQwBWyCv+X879
KNzzc0vjT9MbcYsOvEj3DOdXmybjAIl/jcZ5KTpAogxulSzmpDeJ70wT3AuK/43ehbWCvA+boTDD
IwdzWrcdYlWc0y/6+bEKnqWPGZO8koM4IQK4wyWSKXlHudQb8oK6H0C7t9JgxWyHDklsWbdA7+X+
/zzB1EMpNKGdAhUi3sMMrcgvA06dDvkSsrwt4NadgUY1+ghny/gC2apgTI238qeDk4aMWZ8TBei7
Pl9R95HPVIfEoSY+NLpxuiAHrZMtiBb4I0xDOhTolvNAROW8m7ffzPq4ZHxgwBYONg7IHUDUaKhI
JKbq1iJmLPXLUytSN1qP3dCBEtDWYmv8KR8HlhPET1o3832ZIQrV6gz+ZfL3hEE6poSWSsZPYVGv
dw0qd/Ys33Se7GRUs+jHGe2uEaLfFCzbKWYV3Z3lvZ2BOokZp+85LOrdEgXU+l8uooHcMDlmD78S
7HYdFL89xNdzA+WT7tT4OyyWGEDVUSyuPp34XEPn8A89r2ha3k7VZDf5j+OtAVrlWb9paO0EKj83
G1ZmkOBcvzKlMNzUzMGQ4Win1kDpZ6WctvDdNNhpWs/r7ykkwOAJjitvMjkQk+b/ymxs21BXG7B6
9XGYzZrl52qualuWsSl+RujVlxy6udUPudHFq0HbOXaAsPHXZ/DwTpjo++tBM336vane5JPqa7bW
VYurkTt5FmOArM21vd42i+gqPwPSufhZLiBuuk0e0G0Dblgrk0yzVuDSEiKY4LHrb4gyg/csgTWK
2q4xiUpgd9wyGbXy51CI2E/cqlDVorM+5mpKbon6rl2trdV7JHWXMVOXC4+aq2GnJ6EpczErDcwt
pBeU4DweiHIvyEs98cAwGm8tSrPbJxNOPR/lqrImXNEJtlrS/W8SMsbyP2vDDQEttrdr4QBTDR0h
JH2p4L+ozz3oYSXGIChQU7oyt1Dip/YBm4ZOpJPcd1SJ/WzcjqTb0bv+U76myJMjqso23Rl1mLDn
mnf4yV5Nd9Dn7UiBPyfjRZWe/wEeBB808kFJuiwCcItRWtWgoMxouxF6qU+gVbNPGzJclVj2dRF3
hi1pGkDuMhc8ijYSsM2gxpWRZH8iqwgDntqscWKheL93dW1EIOC2A1e3LDWCtRqPmW+OV5hSld5v
QOg/cD8y7nrrCKtYV14QkFl+A0EZ19etZGaAkuPIquOl1AnnkNVU33xcLNStUR4pcH2Uodg2HVlZ
Ecils+GC5Shpr5YNgfSVRrRcioOWqK1Iknh3H/joI2lQjEafL3yMmnmrZ1iZwzx3jXnY+RwhAwMV
MQsojgbTvxXjGICaNsL59AnRkVy7L/YsoLpdbOIgYavD3t0cSGysVAQutfWDwzsJ8OEmsDBYkMd5
0UlSSCXuntAl/zsaBBYAxUutbRkqHRjC5j9kEXQ/HsBixtGRFCMeWWM+VyeDs9wZ+SVBk266TobS
hI7qZPuH98UougnKXi3I9SuEersSb6TuFd2Q2J6Hq/t/ULFFvXbTN8BuoZVA+w3swhXXTBv+IOt5
Y3HT2MxhVi917hSWL91qj22WcAPD8COSCsYpCL3LGksU1OnI1nkXClxrOLmrZhcVQc+ephHoQH+J
Vyatdk0qvpxKX7Z79S0AQMz10V8cse/ek/ExuADM+noIXcGl3+DgaFzYWzSXTDDbf9d4rq47sw1w
kVdKt/nKo4JxnKSM5Bf5+dQYvkbZE0sqbRltH7ll5Hlb2+gbESDavFjLWeeDhSIkQU+dbebRoXf0
F1PVccTGk+iiY0a5FV0FXXK/M04LAukFi7xBsyLLow+NwWMnChta3oURZjK13xbsUeh+p5vXnK97
Hk0dW92rebtPYu2H5/c/oAU66LYaVqtKSQiK9ka/lZ7A9o/eVtHTh2Q4D4gH5pmJ13KmLN71a1I4
uvf2k883Up913at82pM4n1m5vCHnwHI0VqPFVzZ0rhPZlbnCuE4UzCSEP2TZ5BOELtDCjwXPD0Lq
xO6Jkd4H9td5rnNoQ6MPl74Q7OQCElqPu9h8h2wE9QrsEVxr06Fkbhnkw/anEYyJ0GYuEqDVggI5
+p4YNRp6M2nsD+++eYn1Ug9j56VkhzQvuckefyGplN23VePLIS3dzKwJjO7tmE5CwEERoWDYFcJQ
fj7nIbjyL2fkGQQrWrZk8MeXMfKTI8KT6MGeBjphYPps675mkYO0mwNCnHl/uUEoA2JJLd0ghj2x
52DyXEBjCo/w5uUZYZb6+OfqL3zHGAYVTT/ff1cLoJXyzF0EG+hFWvHDWZQYnJMJQLqCsOq2Q7GU
iD1o7HIL/aIHtjJ8PeGf5HmBu+1/gFucgUOa5igmwPOwdt4VaKG0nJDFbYlEaVEyDOYTOSOFntoP
X56221JDo71Sog4bopxN4mzuwLN0T4stfdD5rhQtzSwfOE8sSt3patyFUwr8EdTVCbTSZZdDvUwc
hGfPM6T7rMXC3WriL2HvYZIcCkH6KB1XNfREVt9dxeLdWTrQ5NTy9gP/RUsquvdAPGowVVOl0VVT
D29ytnActCdVvqt+BksgcV0PbybTSQAQ3DrQD2iGc5vFNGPz4Y3fN5grKvGy9LRZsAWjvGv5Qmtc
MzaXNNcfr0IeosJ/0w19dBZ7C/LFl3cjgVTwvQbLXOtGSEyflUlbjw+0y2hAmVptNbqc+6z25fb8
brJLQka7naaZkYsKCXDDDbgBYpzIlCI5UYpbjJBau/Do0x5ZtzFKZXhJIFTJSscPdctD4pF9PwJV
KRht+n6aBpyT5pqSsOIjti3eFpv7vbuo019DGtpaj2Hozur5itHG3h6FVNEv+z3UW4gDGCSCnWln
UTAueECcaXOWWtJemXqJ+izdVUhSgWyg5sZvBBPuYsSWrF7RkQGBfv40I6TnEaGKWqRRubz7RT93
Og79GB2ozd91NcLVltni4QJTmNvWPRVorke9IHlCAkEm1+33Vl8Jz8VhY8XJXlnzu9660CmzXyiZ
FptprI0u/L6Y3HmVDLzAcGQwf34za+EeewUHuGlKJ/6cglpc9p8oCPyoUVUHEpg9bKRKpKtTppVJ
iiAxN2gXWvzgfUYPCcAw8AW8nh/J/oDROUqpPKxyc9nleteUhGB0O/Lpy+OhV11MijN5Xsv9fVox
yHMX9CtEN077/xZO7W1negl9rqCgr5bCxSpvXjqXYe1MxmBL4PH6S6GkVR8IgJPs0DZ/KlFkDF6D
bE68ahN6X/m5VdnjCjUqDuDQ6tJ427itvhsOqCyVqls67kryR9jLA2WTib4oaH9/9Lg1oODMJlpF
O5fsqpHuSqrCvvG2w8lezpjoWV+P1iRRMkuGy8dn/vPj8NE9xpUoeIVCdnaBI1mkt7fB2CNBgABH
AmLwuxwibmgZq3u2fWNgxRZQSUBfRaybDrjfhZxTVq4kcC4/Xf0vlr1wmCcCQ0VOSQCpvb37EO6y
lUVKlZLe3hKiOTg321itrh3cubzcH1gLmwAMiHiQYSPaF8627Xk/Ye2blM+UvGZXoQ52JzzAcxwq
Hg3dB1jBta9IuZSdvp8l/48HcnwNJ+UoE3vpgXOQhdgfEFvMgu3t+8w9BFi8r8SsKYVQIwDY3khP
GC8t1tRPhiQV5xV79HExgSYWUShFsRhlvPSv4279uJdDkQnYAT+9/GQJKc+DjGlAUFjrtsS1Zbzc
wUToAeBJPyseGZct8974MLRhdgQWNvJ1ZHoPm1kPGVUyED0ptSZT9MVXjduQMzmTdPwizxhsqu4f
YFJRE/cik3GbV4aLOwUmudo26rD3lI2bwd1R+a7gSiirdVbE9jGTvX/my4uwwS7V76ThQ+M5bLfC
N+nr/Bq6snGv0X/V5LCEDSOcqvkwazFLZzbnOun6d84hPfYjm1R9AB7gGEqEGIgNT9/gpnrvOL7T
rc/zdCjKlFrwKrjkD4LHCrxd/v88yGSSXC/y1pueLJ5cKPK9UeNzwaXZGV4NGTWt/ChloaHS3nA2
4zsrlJJP9aLuPP6cvyBXde0L1gmISDRRLm0ZxSFUZaCOZAiMpVs4LBP5PTLVqpGL9Nl2+jfO/LTR
1cnIpZDvXL7dqllqhQnBducX+UNMnIjX7g5+JrECfLyeP/oe/Wm4dm7LnNdl+OfXrK73Jlz+C8iF
bZAZrHdmETGka9FM+fju/tx5r1/c//WAlmtW44zvguwSDbI3DlyE/a73ZjHGadJcoSIPEqTxYnFW
Qy7pebMbXTFK5kJIQifuSigrGItaAjufCjF/7zFiYL9m4WZrA6fVuYcY+17YRdTf9ryoil3h30Dt
qMHLEtJRAni5Q3+uko/Xp7mkDg6luORF1ggxP7IM97YPFgFfq75hnbVDPTeVqtk1NPl7K0QezMrd
dGgbCsO3adqXm391FEFtm6IHMMGinZeBBr6wiSTG+L6J0F1Sls8EXEBTXuYydXWAE+GkYnfJCp/O
Rl2QtEX11xXqNLBGQo4L1iFtkEPpT6La0Rt1sxDd1IOuaXLY8QADMMslTC9OZQKySqY7k7rJGkST
E83fUqVvvRNYk2O0TxCvRizTvhQiZ3sry5kSQR4eIprdEEzJ1sg8uqXIRCkS8q7OmHROqqriKptn
xqTAWNWIceNpBie6rfED4JG0PQe9gL7McOX7UZDIY/5XThsAeZET3ja4icdx0C398aUs/4/Qemf2
YKMbZuWRunijfGf7wP5jxfGjFAWwVmloH0VKPUsVjZdYlc/lGtW9sjuyvwudFSGh3eFf8NUy2hKy
ONzMo+3JO9y8jAGnNYEZR4o0V526By6Ye64MyVpBgdvEASl6FmBT4kOMZdYrrlkPNOD6PxIfpfK4
S9X0dVgqrhu6kEMpfV8MlGR/Qs9kbiCDBeAewHqocgL9w73FSsOjD1lmQnZnvJ3p0yRt0HQ8pue3
KTFqojQGGsS5UuaXJhpEERzVRw82uERfXfzwf5l2ZuQkBMegWb/7bOtDfursnqtMnYHK6YUrVe8p
qcEny4uwNhJABkxAlvPYYLJqZqFQEGKNq4W53KIBeTubIhVYDhZOUqLmcyW0wajmayogFXWgFGjA
vERsJCOA78Lz5jDzcqk7qyv6mwHlRHSw6q1278zd4vwP/HV9zb4z5zfo7ety4oI/jHfGov71LQB1
s+OUdgOsU4/Dut0rXKhI33NnXj4QhqlTpD1tm76m+JjtMkOrxiU6N6I8Y2ClIqgl0wIH4jwvTM9B
TZ/JmZwQjcRNXHHgurmvgsf68Mz6YtL8tk5XD804xCiT8Cf9k5AbuRiQt7E4HKGqjPszTA55N+oo
MyxtBpyr8zz4tO+dsUC3ugpuZQgM8wCbXeZvA1tFN8HYf5sFiguQv4z3HEWWksFeL+nhnp+sZrxI
RR7x/wQkU5fvX6UeKAHZTnpfAT63xWso6vWRRc3p/BPx/hMqQB4Fnbng0qle8DwLuvPQ9t31oSsV
g0vzw+oCVYgBHjsNC8vbsOXi0e9hsMmBo2AKPlHViXTjwBR0z+Qpg9rx71z65IoXuIAd4S00SoA1
TqihVQudM8C5u2aDQ/wiA8K/XtLlYVS2S/HEYNI6d5h7Zsb+TsEGrz/hpQWW4u1xz8+b5gbkKsgM
hRpRChCXjznzt1cp2DSa5mMZHojITNpJMC3FwbQUoy5S0XsdfL03DyqboMO8D1lvbWn5LBAOe8V2
mYbVRIUnN8slr2YPAZSOkeMF2K1+zC1ugK+bnxgWMBwZsgwsr0W8cR0yctdw96jMBKiQnFZIsWlX
yHyTrGZbPJne8mICwYD23TJtk/3e3YlwWvpGWxISePPCUsWUyQolq71z357wMBxb70LzxAz6hc2g
0du3YleWLTlXDhyZKxy69Mc51xSeDxE0BY0i9g3eDIrf0idvHWnHD4hqDAJJjbeisxm8z1Jb2zvy
zK21Ogky3o4Ic2AA8FVL8oiHN2VzTlRcbVI05OwxMdzs4+799m6vgKP87wpRa8UEUSH3eccC4vI3
OVIVy3C/kJJOByyjMmiDCgKG8IjDl2VKxkOOmV0048Kxt6MmAfE0gIM9bASvPr5AscjX80Ww33zg
xmlaWC+TAng8IuJ3XwFUzxSSvMZmljziUY+qv0FTKMW/b5+96TfxcXWr8K2UuP1Ga/68J2taQPo/
iwCj6YHVFDRtdQ7rIy77Qdx92tZHox1slulizJZrVhDnY07onQCULHlDEfQ9GXzAtxzDcY4pa2f3
k5d+v14J4vd73fQevw8EnpXJs5lHvvQv86vSTevsrFNxrIj6QADu7Bi7hO+6Qm1CyXoloOUQWaRq
M3aRFqb0K5L9mtxbGKGe8t3TidXxFvmAZADMj/7qCM9A9th2Nm6IzW/clkylF4WSQc7buTzkmhPp
EPPDhNKm/cCWaB5T4NKyVMK1PM7/4oK5YyxfoxOTXAGLKyonqHrvWF5eD1AOOFJNCk/KN6TMvwXx
fa9FukugnXFvTrKkcERfLM24dQ+rbpGHLV7+WLl4PzgvLfa/9i4kleboQG9q2Dd+zKLqj2C0+Yw+
j658dngMo2Q6ksV1hufsRAx/xbDUw+5nVezNNtso4bBF9FH5wfWIGRdu+ghwfNxNHU0rwzoO3UYm
U10gCLKrcP16BSXYYji0RFAZ8p1PcAfq9KSj99aeMQXpAGe0BUgLw3083wz5o0bV2TmCnvq9olo6
faCrcCX2Z1XSwGZhFhbTONRXiIhzfhihYoWX79V0kkf+6ikZiRZ8U4ZbZUCPmGQAd8heVXfn9Hsh
SA17LKrwwBKy1REr86fxiGkD/soGmCQLNuE8nC19A9xarY+3ZD4wQIUVotaSDiWSRlMFPY/BpfoS
5dKrVDeMV7hhwIsfFKVz4mkJhUzNQdDyH5d7KwI9ks9I0dCqtjKp0M7QFZqMn1YQrsvyZWhzusPE
QYtk1LFaj6+0oMZtP4oR+NVrIRx9BCpNnyfg7q3hwmhjxiqacIX1keJ1QoMMsrwE3y6qMHlPRD/d
M0YDqi9/4GMBru2xXRBYabcMn9Am7plspXCC1abcOZXO2gmzFl7UJEC2g53uu3dR9HlTVQ6aDYM8
WjB3wCbve6YYIcCr4LGoNxNzWmiQkqIM3Lrqdr6aswjpBWBkuWvP1VqBwvCjalsx/FSqLlZL6LPR
2uTtU+sLaIejXT/rgD/7UsYLytgcKMIZvm6tNt5fPuf8zfhwApoDSsgujen6/zVDrmdrkAcAdrAd
EUC2RKbgk2mVr/YBrk21QNB1T4dh3k5aIArXnoF818iZFeGTLm1dEVvwT2NF7XAHet4ZbkRCh5Yb
k1VCr1zwwwPc20DqSp4etF6y/5g5UGzylzNPswEqj+UMpIduzQb5iy6/kF96Od9DYCgd2dXoKeZf
2AuycKsDpmeOVF7xVQAo34pyvm45VB+iTz2qKzAEf4Uj8TFw0y5esAP70PjaSmzOnme9i0MKbtQd
KsiWiDctGMfYvIJFjVFGsr/0Ls8dvrefCgnfJUrhYtTpRvZr1jD6uka2gavfu/LsmHu99hbynjWF
c9z6xNZhdEqw9g0IKmOp9Ki8pWnMpc5PNmZJFcX11ncM/8CiT/dg/FeXgpW1MY9K1ASMcwOj6khK
Qe8YS8a1PyJ6EdRp8V4x7tjkv2IGlBGOaHl26W9/lS3La+nHjt5n438ZZcNs+qcG1oRKZDbDC3js
ZAZ7TOtRXfOCf2BSHA3aDGpt3FBVIxahXbhK4XsA8jD9a04Pn7JUfBUn1e6L6Er01H4zIZvkrw7u
i54ndtn2J+snsC3lfcNQpnjteqcV/0jnhgbxgXhQtjghcEDdquwyC4DDh0SRNakIZRhnvcy+RO40
1nHTydFLFk7bI0ehU3D81OpaYt6kQUIKaVaEQ0WfXDavw2B8ttBVv4Am9hdI6lP6QxChTd2/ZRZe
TeU5rJvDgZt6vv35BNmcYwzd7wqJ3fY4KEYTXSUaxiyAWP/w28eGMEo/4+lJII9LrIjXqCYroZ7J
W2cC5ufpu9PY4ughLhuQhSt85jSWLu0s5y0yDC9MLjyF/sLJyo8DQSQK3p+RCavFKYrCQs6wm32Q
ar0wTBeaTe4zIgmimD9y1lZLWgKQ5FKoLVGUsyeYpnO5l2vrkWWm+Qe/Ef0f3b/NlKFwLosx1g8f
KzJmalILwvRZ+scEBzaHqPSomCyoaocnnouhqycGCdHPfl5ZCkmQpgKCV60aRHDTRXIn4I7qaH+S
iphjolMDoBUyyAzAb0fa4io+9mci2oUniTuKKbTv3qWnUwcmHw+yEHoKTNyG/NW8ALW3c0W+30QS
32Txocz0llJwDD8r6I/8xOhwSnGrSZS1v2tdbUL9Woy3bZCBEov8Fm5X82dMqRzWc5Fy/MGNaR1E
WKaNgAqFMLbrvVbpXn7EQMtGX04+DhYCbXyTFDvNCFa2kiXBxo0ZW3mBhnxHIAskHBpIj0/G6EHD
+Y633FAWxycN8Hze8wOmRB9YcmtmCfIFrngU9eqKMh/cr9D0FRNR3eZ/bX9gdlhemgGgO9oluHuX
c/kK4dGHNJGIquFqTvEAD4n7mkHBFKeNwi2a9ntvE/d+7LGAZaYCuaFN2K+Wj2ln/BtJ0Dp6pbC7
9GRXpEA7D8e3FwNn4jwvyTe8pshWNpisKIYG4bep8nwpzSAKz3ZwpSdXVIc3H0DpYo9GOGZHUw7g
ie/+MvEr+SLQmmkBZBCOmqztYi3w9bXTfqTfaw9oy/yFzaZzmYZdFI+Fw1SdTuTK2UfH7o+SgCTV
bnzP7js1WqJYTAvFLeQJJBlHaq1Mp9bmz8LUjDcP3NIVobbzc9xwJYbC+DwZM/D88LKrnq1MbcsV
T3YQvTiChNLet4nz5FvlVZdVdO13OFAj7QrTwQzYXwnMnHB+JDJGyi+6/4hcf3PRuzVkH0KByt44
0z5r1te0m8DH/G/QjCEVpODHucdLvICF75674BYMnVxMG4XWqcXqekztIjW/NNCaAR4G85WUSNiD
CCViUhiPEdbje/CiLy3zMOJgsd9v+gW4g+X6tCR3CGh1u960gc2QyND3ul6eLNFWGx7vrak6sHEi
oEjSfPjNZJ/8xLKaRNzQ23XjF0MWs2HGCzTYp1uRm3tIDl5VjbURH3sRGIOiCMKmWMy2TFnHDfmU
R45kGVlV+jdnhv0M67aURY73H2frQ1r/5oLzkN8f7+a3dkZGV0u1Gy0ICFZhIt7LOAspmxZ+dnV4
y80V3INTpcoRvbH28bIvNwtRUlz65cgr14H6QvH9QwGSqte608WzkleXaTDKzLymWrG2NRZX0JvV
2Uky5DmuyiQxP0cuHF+DPNYtBfJsyoBu+NGMRK6yowThIwTCt8V5QQzHSQvStt+36UI2s6ZR9gGX
6DPT6XfKSiAg+5A4ditUDACqJ2blL2XF6uBIzsgtZrVCfLqyZVyrBtNZCs8Ks1qpFEBm14aT6uu5
HwKkpyqpMFoeUuX8YZnOTBIzy9MxqletkO/8S2871eB1iXZ0oN7Mchb9TFYP3E2ummAB3jyiJ6YS
N22E9+16jVUvaRt0F+QVq5/7RETc9tbycn+yzqHZzbh6cEokQG0nrHwp8GzIMGfBin523vgiLgAN
GjEDgHPLsXOPagtnyOnJjsATV8WvrvlOQ8F+LxjizG78TTNED3r0ttTf1qpW+PphZZCm7D4IWbhb
O7Z+8unrt3WPqhM/6ko2+GjYGGtO4PuFQ0rFA+4sgkjwfHd8Ymhc0onmCodBliVv43dpgUmRhN7k
ax3y0JtOxjBdALdCaZi3AMjZyUGUfZ9Dz9D3DJ99OLlSFqoen0E753ABIM5ntJpmfIAY4eSoEW3z
I/M71VJUaGe+uVBF/6hvXcYop/M8ytp6Xrh8wTtB0dytB8/nn/2lGwLh/qk2Q6CqYgW1QS2om2da
QdtXVmlvJmqjCiEMtrQD/vDm7dtSQLwj0QxY0ij5p8BU9oXzRs4qHwYSZ+k25+Av5X90aNsPbXvw
rkK0WhuNfkAbSuzrClw5chJT3W2uyYOfS+6CXKSjQ5zcXsW8e0IplptLLBgzALojzaPKRWDa51Xb
wAgWnD+wDT8W56XwAssEFkYyzq2dkUzhr9/pvzWb8PUBp5G4RtXtZNFz2c2wZewLkmwm6htbkQGf
r7La+0z5hspUXHVFkr48zv2dzaXE2qHyJT5mP9jMUs1cWXpOWTD86bjjA45lyhA8BxPIr0D+1BR+
i/eAUm29w2TwhviovCfx1sg6wTLrwhb8Avec6e9KAznwqWjsgeatEIkPw9/C5ckxxCZwkc5ULMVt
8xiySzxbGKIHbRMg484cYimt8ozSJZp7vOtQKY7Hx7GJJy6jA7l3jtKme3n/uXu3Ti+tgyfclomM
xE1cLI0IBXxK3exNwJarfFqOoCNAjR/ebOQf5/DaP6Zb+8tNcMb8sQM0Ab7PUK1SwoNPw0n0Wa0L
hcPm0Au2aSnadL1429CVvTQLNV5vpr2sCz1nk/bmIYSBhSt1xHapLxR9Rc5bgSDFpHEhJYrZFDym
FAF1kx0MFo1J4CO/cNcbP4M5+vZ+Dx8Y9yhly1ieXKGz0HXMTuSEDrN+B5k+8H9X2VLhTlxLQMG8
EYlRlcmMfuJVyHitvC5u+WZp0Eck4WifWz4jpdBQwyUGcEiNw3hcaz4SrxJQC13Xapk15OdGOAI6
OpPthWbrCQqisiTijUY8vT1teDq9Ss/8fYNTDB5tXtN39Rd/o4yCJke5SkVSzxk4BJCnzJvJEzUW
puHpFfTc9uP+czVFxVriuWNDph3+XU60f+4F0uh5yqGcsPQC6kiyy5TPtkvl//aAnkCSlZyOoFhL
WP/wPBms0hqOsDwLA9iyiilEd5rticn/EVIp7DroSs8NvAPGNqpC9CYPdvU+3vpGePzwGQaGimMc
Zz415pDNl5bbLqxhgHD8zWrGB8ExXtwURDMLvzBUVmlO91TR98ELUk1bqshd2Dg0Hk3cBzKzJAOv
ZA/hpUhY2RsDSDgBZy6AvT0IbPt5gb/6eGLM2AsHEVZM7C22EUZhCcywyNW6EM7Sdcwulm0fiCzS
I7Bbq+SQUJ7EUCpgP3+R9y51/s5JaHrLV/aCP6iCIV0iUe+mgfRk973wcPk1/eAGS3fzb3kDv908
xZqlHE5lebRSn8ppa3gqSpIkIXQgGZwBpYync8ni5gXxH73rxLP23ALf4v5+u4jatcZRjUVoPNHE
Q76tOkZHb4WeC6iJi65Wfoh20Skwp8yLyTEJHcY+6bPwrMDLg2IZNeDmWQoz3vtDch6crg26va5I
Blp5Aw/4wMApAZqTGTD3z1Ceym6d/y+72PJZ/gwvHFHzyzCNuXFZyF/OMzkMUvfLO7MGdR3hkACU
SJwolvtColhmMuPPI7XSKqbzgfuhj+WgxvIRW9LsUDgnPeS7ugDXba7XZbdqrShJ9EG99aQQFH0/
VdtBwTS4w7lK2JYqP44cV8BIkOJCcFk7cDI1xZFHAnaT/JwgA+V9yAUSdyIUYZAMd6Aaosfa3ChD
YChpj/AtI6flStw89M3gJubMSEvWy0/zl4948KR1SF6tHQHGI66ogoMMACdjerwL4V8Na+OQk67o
daa+8m1F3tHk6c/h0D6YWI78fbqAQKHrl2QKP1XiIs186oTR+LXfA7bq9gAeg1URMPLwBkblS6sD
HoRvbcvnOUOeRgohpy8yKt2n10NiNTIRokw2nQ0qwuwGzxzoIUUr9oB3G8I0p9pgcNp2ZfeSJJz9
QlJJwYYFXV29P1egtc/3tt+yyOxjHZcqQ2P7ixnz8dqM0GTMqnoHHtK7bOl/BN0zw8Gf4uYCQ14P
x2n4Lf9lJLNX7VVc+Shtj7ATZRUwkLU9OaKmYik/yjdTDlugExvo1lmazUkk4WABY8T9TtstMIhf
p9AGjN4ORRf2/IWliEkue4OHxGRkYWi/Eq1F1JtEbgY0W5tUnj48SUtKdM5scFRLa+RIg8UG7IND
k+6F3SioCQbU69pX/tC4u6anMd9/UXSH1hrpu3egFdN81mwo8YUprVcSAjBef1HPL7rS189c/fzQ
O8TOaKPStmOm15LLB25Z05B3mED+AV/pkzEb2Nr/g7kfR2Jj9F3fGQL+OrMgvYZl0iZfyoKEQdjX
ifDbF5hOPX6XtROgcaUpBWhLqefYIH/jk1uBj9Nvae4BktpY3F6wcjDubNJ067fJGTCDncLgWi0Q
L5POkpfFD9j1Hf8KmSvqQRemaba0/rYLvMejrbb0u8FZl0m+BPgq4Pxbh1ZDYM9GQ3KQA8O0T4xz
VKsZbQ2kE5dqjrrGnja9b1qNKG+pHss0fj4clmB9I5lH3+zFivLHux12V+aesSwoUUgL90LS8Wh5
QZas/qUFvfAWCFzYd2jIePjfKUeKzZNssBszVfHRVZgQvdeB16gBTHpGjTAaRe9MSrML7rnsckGQ
2Hcx9+ofK7GzWDMcor8qcA0/pdEN7J4UNqOQ/7OgXy8FMrcekQrwEHXOINULOxNw1QGOqyhwd4OD
iYCZKyevbiiUN0PyxAVpZOjVTExJa5+njf+5v+Fq1e4xZe1YqbqRDS5Imh+Nnpb70jfbX04B6se/
S+y9n/yDAdDblUb+/TcGuiuu8QP5Rdq/4jucvGaFT+7NR4milxRCsKp7jMmgnfala9tHuvvotK02
mUJgLaZzsgHVva59OqMuCNA1KLSn/D7JLsV1+leqFKG9r3Ifa1RCq8TX79VWVG3ji5H6773k1O1I
sb5w/mVvT7f5BEv3h4YUBmS6oXyqoDZngehHhschU208JcdxbUFe/KN4JmQh2vFXvUzBY3s1orpD
Ih3lNRFkcxURggcvLCLq9KSeSoMfrqZLkH0xLS7W1cCgh52sxjsz88SXxBT0OMzN8O7QeEI8rye5
zy/4FeLMQBpsHadaBiT7uVHbY0P3UNEIZD6jex1suSr67C3o3nX00hXBdKGeV7aIcr9jGV8e6kr7
JUQfnjXG6n7heObU4p5h23u+gyXULqNlT4RkJ0kzpyctpMnu6aqfBhXWzyb38m91W7hBHjQyJ/Ej
KtBJWrO0Dh9bnQ3ScYcmxcAwDBOKNbTzIevXIlDWDO9gZR3qAxyIDvMCF/DnpfIHsl6LKft9kC23
4vzoGztGKRg4jh6UL50tUP5ekpiqpkM2YXKVZt4TQJH/w6Po5XnOi3Skj9waP450qEv9pvPOcR47
JCMNqcsxDD+viYDr82HEW86guRDVMMIHVekOpqROFblAmw3jaBPlK7CsnSGpOY5Au6RYky+KCwCL
03DR21UpvOPeV7tKVJ0wz2PWch0SOU1TJtWiJl1Rf5oqtPFYHKae0Y5bpDxdRoq4WwWmuPb18Fam
Nmm0KzHuF1wSbSJ0rJksYzuj7ijarvW6F9czYdWSXbuJg46uGAetOClyMjw3L0QyC4dldSRCl6El
8waL6Ypg+jYT4Fqcmf7Vf05B6HkqtQCNpG2HlQy1GyIKSJSXEgk9Tg87GKn/qmNLgx9km2FSx5V1
hY1DgUWB3Jp7A9L5Jw1WciDWVrKJz6RpCswwOtVD0SbuvQmhk3KT5zjf9H8tfgUHDsHthgj7qESx
W2oLdqGq1Q/erogWkj2VDeTV0ieVNWUq3RjFr+PZbpSIygYnVA5Ho4/IJs4Y7NzVEWgTAZG+esQF
wD3SrRSVhl5KzNocDNGoPw40lZsWL1890x2tP6XnxngioJsbGXrfDn8mo7cool/73cLREtB2zU2d
ueuh/KA9EsOckv2/r0CBw7mW3JAyGs2zIKs859BL+ytCVqvhPKNaFp7YUaOZ05B9BqbOPr6mQFHJ
Kc678NuOpk6ZnkvJTVLqI5RPMsN/2rgU/tPThdCSfTGm19vRecb9u9C1zlkd2BB9WR+66T8CFW46
jST2jOR+mYRGmkYamr9foMm4VLlgxtquribJDe+zsnhtrR11G2/g0cS9ACko6V1WS/sRgfhorQfz
B5PwXMEUyqmKNbBCgbEn8udFQouEC1EcfGkjw2kYSOtF+3LWhzX9MMEN/JncU4GhOA0Tcyuyto4G
Soc5eP1IeaIoLX/a7cnMneo1lCkNndsKgAgdOYgTjixPF0HWZo8ei7WEvmIegJWFx25+bK4F1RKH
8Jt17NwSkO2CohiLeVfV74REWfNYZeJrbyJBW0dfy3dWjPwcH8g2OgkDUyw3snowtJY1zq9YfvW4
UkF6XNzCF0kzP/Va21EiPX2IrxtZsAHHAnmFhK9Si88aPqNsJgJgPBeymShk859MFMADtA139Iub
nHTfIMs9kknZ3PAsrS7KDnLEbr7zBo7jLHca1dBEZugWT9lr0IsIdd90Gd20dWKHzpVtWimkzKlr
Nx4Mre4Br33DXqpTQkdz5czbix4ItaDumqakzj8VzVXqFVzn9VkNY23i/t4q4qJvitjueWMn31Ap
utpw8XDxd+PYH41VBWzUVhaiR9eHl3JPKf8bp/h9Mwd0h2e/aVGJe256bdmAgU0eoJYnIdoSal94
LvLo2fYz323oJKLVVM5KuQPyLkatS77MQ9Mm+Y4U+8OocVeo1xmVmwRg6IIWIHDL+kAJK/FxXk44
nVvZhBSQ3NjtCE7zt7//126+h1uyyji+5vD0+bZzV5TaqASH8symQMEgSfWv1N37bW/+fqqM2kia
oMZtAbvwuHTc0XoHSIXvYMCOgCYB2dFRtXQ+6uFm56py3LLgV43oivLtbC7org/UjW5kPJ6RaxkG
BsuKGwVZ+dfRrN3vfd0HhiXYFT7oERUyVjVZADSY7SCSiT0VLvrjJA7XMMcXXVcB/5O7e8FHdE22
L45o2TOno4Te2/oQjZmkTFY9PUs/cREEkvn28RdayrGZXk9wIeQwnZxRjZkb9n+EFeNvd6LyFMQA
UgA3yy83NB81H8TUKB7tTy2DMMeO0FqyUjUisnO/lCmGGhY7TKbnpblLpRUT1aUB26phGeJBc8Ar
2RaeWBnQZE0BSrKwahQOyrAYUEO5uweLjc6fXxE41mG7fRVsj/bdhnIq4OzRBLVg4wtg6xguaNjj
MH2D+I5/R70J2ggkd7xpCDlqbToqrs5Rm06siPJp8nXka+HpE/IVE0EOXQh8NJhecFloe8ZZ/iGB
rqNGzyqYF0aeYLsEp8UMlU742X3+ZWG2YPy0bOAhyq3zWXlPD4LsFwZmV5wjl/EA3ZmkEMCnsnvo
g/OrrUiLuh0/Al+afkEEsoaOl/rxKM8RIDSml9fEgveoqI6p1k3xjJkhIaiTSgzEhLXexBKwoxUM
9+7DJOsvmDhTnYM+xkV4W3PkztICNZxNgmEnq5up2pq3AbAaUjOaU36GWNy0uEU559G4d60btmaY
meL55lsijmShVTkupT8sYQ+QcGxH75yYVZq92ggkV+yUt3/UgqaFtw6fZ36m39zehjmDXzSj7eSo
H5vHdUh/oUpNIFZAtpxOX7TPCMGXMLTx8unQ9Do8CHBUTCvSgZuE/VeXDr6WVi3gYKdCAQJ3BoYh
hW+PiCMLb4Qn9pT12Gfgnale1hkKg/TWv7nS/mCwABy9hEfOymafmDfsDNEm0V21Gn0ZXvsy6NAO
tjqxh2RuAN2mo/Lwltade0Dehuz1ATcpv41+9NnooPRq+YG/ORoyRgUNfjErMLBhbGZ9pkKYgVvl
TjahXx/wsIHb+jJEmM+t7zL0yq6MfGOInzWiY1ziaKAZkOHsebvMFN2gqXZ+vipvzZSbkwrs8IDL
Z6Mtn0CYt4MUC5EQlY6RI27ET1aCOysr1CTmROjyiSy0EhVGqD9S2ZghO6WG+MjliClrZxxShdmQ
oVF1C7c5/TRDHByfSBIOrLE5G+pKHkRALAb+/XEudr6XpWnynxEbvEs8TyZVMbArKMwnht67eiEo
+VbO5bqF+S1ILHm6DcRiiuCHCR3obimFR8kRJ7+uQbooMjulFHb768/8OlfmsKcw55gAB5m8EKpI
OjONovyCBBSVUS5jhOhBdSh3y7Br7ODaVftrIL4vxEdH4FOwdlPbaE7zDUkLrjnqDIWdbcRUSEPg
TaYALZspKZ2lP/RQ8NnKv5OjjDNCOz4phEkrAMvzRPYb+mGiugkQwk2UQzX27NoMIIPbUprGBY9Z
TFRkouTc3EbVQoqgmydoee9XqgK0Ep5x0Nv6+EtSyjjgWDEZyJpOXac/78KrvawpN/1oR72e+R96
UFwH1PE/gP1IcjzzgXPn+9pZA9Qb/odWkxBl+onUA3xgb5sFD+cyOyiZ+2y5OR8dkSJK9nXVE7z/
svVRrqEJDMDddML75YwOvnkJiIM+jlyf1rBlN3MDPD2iyRQl7RaZNRJQpbyyqRBbPOfhbFxBdjtt
0Y7nxbjHhK6UzUKfeZX0zSZRW654cGHMNR/ZyIwo/kIRJt7z9t0bevwvoZ911pkEefPTOSFujnKS
cFpXCaUXPLsmXgke4OZpoWPsDGrBljHAByWeQYfJh53xDJS8V0oLqwKUC72Hr2AuU68UzuJDPRzl
yigZoCx6YeLk/neyVHjKjoqElSglfraW89fEg1VRYU6WLPcDosgsjMu33GnoEzlz/fuV3r+a92yh
kwI1xS17c+hT8uINxzeOi1McJwyG9K+ipp7fPvjiWpOO8+Uzn7lifx+4JZyCwO6v9J1/GSkT7hhN
VOlZihtK4kIIcxPbexuKLvJdIAaLTIo1mWMenn6xlBZX10IAk/4t8FIrCabtmxLKBP7oacvBM/WF
YvGfcCnxW2bbcGm0rAlauxihh7MPNq3+rr8QpA6VHI9pZ/81COA1vKQF2Fh08+WawglrkyWrK6Dg
/aoduDG3WRWEuIt9BboHilQpiARwzB5O//HtlLQ7/JEfzcJb6+dIrsGYAf0zGYexuDZJvb+jUaS+
FgD9bexsgEX7bPKI41jHrGye9aP0H8+R1BwslHUMIlD1eafr/cmO6WYEbzRMkQPkahSWu+H+EQv4
7UfjFct7FoaEE6z+mJs8X6vMjg/DH4jySNnShJGKQIJIAJKuPOj0FL8D45xqbVDq7fdK6kzetvJr
Ze7a7rzYtDbXWgKSfGra4s/XUrJHN4NmmPu4TyQCTzZpcSAPz+/ebQXvyZ70zkji347QKrT3UraM
uvtgJyy3Wk/rMyksunIK+lghrPIGnnBzBgn/d+0XBg/FcdJchgLtdEyBrUzUI3mUYrgA5yt5yTc7
zUbevTMrUA4GPH8u1MIUNuR3izqLtBora1NAJ0TvwgX7F3c0lKuaZkDcysxlKFn21xl3jAbMnQKj
F3WyoQ/gE0bZxG7uYhbCeRMnQqCP3K6j2byguoP/JwQ6taJD6KZuIGJPg1qobF/d2fj0fQwwCNbq
6PZ9zLOW6dDWeXiYJ3k7oWSIDcmoS1anz1+E9ZUICWE30vb3ySDf6kcfSOU9GSjw1mA1WLCw67Bs
ajcSM7aRd1I3bm8t4oWKDep+6g+w8hWcT9kRnM+J4wTIBJrCHQ/JkyCtPXi8m0MJ0DiQjmnNSQ/Y
2lmyuwExwNqQeDT8cyCyN2iABbtdifX1azUWgWLwUM/R8VO7u5bL5B7XpCLtPNE+O5Tut/I8jYYH
wl++nDRyC5f1V3YY3t9wiBEdfIHXNfxmQ6gIJ8wfUWjKWa2ha02asqfFs+OrOY/Y1+pvGNMEWJzL
NCclM07P305B6uWTgKmjZvSGCYJZBHAnNH49vBNzQ6xs/W4B6PKbtR73LTPiNr6MBQS4urNl9Xps
TGjzlYdEOxQx3hkPjZkpNYMmJA9yVeWbLMSf1bKawy2DdhcB3xj05Cs9CmEWW9YhT67GvqiqNaLP
UKXb+DIcmtkgPxnoMV0G8UX/NLE2WBbiKzHkU2DFMyI1N08Gr+zQ9T/yQ4FYk92u7k1zhry5VZa+
QGUHF1zoYV4r0JqVYXjX8GIQ1DtjTtiwxUuIrywXLGOEtEx/I+2kPzZ2BsfcQyPzOWWc3yE34v2j
EAwbqEHN3cFnAZJC2neM14NNwqzP7d1pEcI0LOhCV3avxEU5rvVkHviv/NiEUVCnhXYRL6g8ui5A
1xaGXwqrzAInLS/gpveYoXFHWyNIycGAbwXWPPyokHhJFUGqRBbemdaU0fGcWKkggTlx5HVSFw0l
iYR6qVQj7z3B+uUCn2wh7G3j/1DjRULjRWyw+WXdDcD0YJkZNhkUbx5ncJLbdoC0aHiU41ZIEbGo
AEF9KVuuyqlda5TyVCh9KEzte5IZWLNelINCu3j66oMFjjU03oXGMuHX7MxomBmQjXl98qDfTBDl
fWavVNkloeGgjgleUCngNvVe5SX/h5gtTtcdvLECML+vnBO5ghC5nWj3rbqLeQO5mvs8kcizZQSC
1dBjnQNa4hPENfQnlBeFFt/JDfwEa7P8wYhIz72WEWP4YWqBE5B6Ym23/lBoi5iqx/QMcCZiSLqW
FHjSJE2RYFEbvJAHkzMn889fo4sNs/jbae6TDkHwsdxbUm+rA75tgbv9mD/VBLRgtruNmOnj94EA
aids7Q+J1/e7L/IrJC7mzURO9jxcysk2BUt5C26x1HcD3qPFjSrMog2xa50bnSYmB3Cr3N6k598O
cyK4MMm2AQx2qf/Dqfil0n7KSVgpqhGWvFXvlZMCnn/mnf1zB+hbdDK+G5pW5/xHGtnQwpdvRcTc
79uSavx0sg/Dl3uHrIJwz3sdla4uGhmcmqZNNNfugc+mPYQYm03T2auOsyUg3j+cVJjdEiiyT4Ru
IrjtXeOFim08lQemMuuxGoddtl/g8ZJQTXAnxTBDuXtwy3t/ZLJ0iMoJiEvtZTJ0MDV3yfALf0is
3FvxDYKvnfpEkOtCmQmI5odUUVnTv9hPxx7l43gECcw4VAd9hnKFG+e2676/pMPc+sRrLnuNDosJ
4no+CxDQlKSYM7P0DOP0n8WRohBvnbac9DLg9upHUdZKve/C3mDqeofgnSQp/jNtblk/KscOck+G
8LOrDo9Ve7vMy6t8fgrg9oMs75xV+Ekzs0h0/CCGMw5YB1cvGC3fxNoxQSM9Y/t1USn9vm3TCy6I
OEN0AP+WxOOysbXnP9GO+OAuPuejTdUHaovpirBidCGUVuWdIQAXULmGF6gh4PsjrA4C8jqjDxjO
Q4VBGP4kB+AjfMhAleYRf2kB/QONlfk1f91KVH5Hfkv6IIZH/5xLCppHmONAEVMyXdYcqxM05/tA
YzXrMxPQe2So3R0tFTiKF0q8RMuuAZYAeslA9gRF+e3gzB0K/CEm7pCunAmHmlCznNBbrIaj4lhl
5bMFRf4qeDazZxi0/Qjkv+h0u0sUZ4HcjriEhnLL8Bu9YMTN6b4dMxBuHJjDs6ndmUn6msCwED/2
Ly/9Ef7N7Au1lmA4lkTp5BJy58CidyUMoOfivMxydEd6BNYuosMm1+ChPhts33Lxwoh4pZqqOJ7w
B36LWobNCVQWzPIqbSYLqNqPEAugW2Y2s5RhLYJyykE+BntDa+BrPTgwOw/DJnzx0Sd+LQoDIX/5
KvRpAa+vuTtid0ZjUlJ0jg/ARgh8dmMl2xB3Uk149AZGJjGEIcqhLQ08Aoy+mQE0Ei6GIFlVDAXy
jpHxFtMnQ3LbGbL35x3PJ4WvDAm4k65OtzTZYBDh23kxg0tb0KRN6xe7rmRxEGlpcV5ucJT3Aqgx
DToXrckfVvmY40WkLkwahjmwyRi+CXV12z++v5kL67iOljXWzy0+T/ATQNOLvi7o3Snnbk6sIMpW
oXrAC6B9AAXU1vZiARQgiSDAusTZcEgk0Lhry3PvhzFhpF1dNjzMExR7pXB9xiS6rTuic8cB8RhB
Ro5M8khG030jK9pr9F87HSrU8FYmhA62uLlBz+Khui8dF6fDW10bAfem5zkyH3MbjdWyBAWYCfwT
UyzqAZq4BwcJVq/fSB+cLa996NncBF/YBBwEPyDUjDbYn32CW9mB8PGm8eIpB4mGAmghoQRcg13C
TfbO6NwZXiJLBbM0LYpynPogdkTbmmn5NL1YZjsP+TVuAwOqalNBtqx147M2ZPcybKs7dN9FvBcG
PzrDaE5rUM9TnjP/NNQEOPOkTTlvRbX/0lc+ermmBZX0G8A5gI0k7piOJrVKnBttKSmf/Pmf04aG
gvE0rJhbqR6p94DuixyILanQ2vcY4gMiyGCEf2fUPx1BcWsU++rGQUPWUrUg0XQaDWs8dBgSUnR5
MBnTlokZjsX7wIqqPq+AhIFgkTqLZUnKU5SlHdQRTaD1MTrGNL649D1pJl9k9kcAD5jXcPc5YhSq
7gEwK2qKdOGcRt6nlpuB5Onq/EM+HfWM+rM8EJ++jnBFEaxThNIPIWhsrlG04jWWhSMvNSU6QZWk
gI9/aTz6nzwy/OVi35x9JOfQdhzBSKyyMKJ7KO1/jf5NUkoH/hj9Kgx59OJWt8KZsXCHok9O7lPk
7JzKpM70ObHy4Ishnd+Dfoce5cu0/uVvaKbSTX1dCLE96N4maHVzhwbxr7430Nrd4n2rH5a8O4ba
barfmmmp3pYppD7IvIJ0TnD7YneX/LQbXgzNYR7GPCnkia8C63PsIIfKQDu1TVcEZ6LICMhCEk84
xY4fi+/XcONb6SbQH9DAxDPy9zvcWVy0/kmYKmP7cjnpUaK+vMHrXn6LzJh/xM1EjVu3H32Q3LfQ
KXQTqmAlSb+lITJYVH6WNu1J1vW/WQNPGvBdw/8S0LbY9yNJeUnFZw/Hvt5q2XbK6q5xjXKUY0JI
TPdioQIii8iZcI4EVCExaST4l3PLNmXS5+n0rsxZOd0HUbFI4FqQW6NxQSjtFJ1p355ZdEXjUjmn
K2i6/qRn+2ZUlhbrpfGVr14A4+JC5zJ66+R8w/+kyReg8RVKcEhZmHHZtIFX/8SYDs7XK5/2m1VJ
JSmyLVsB0YpBHLSuAm8TxQkh8ySWQBbYCDh3DaRygW4W9+MT3jrZeXKJzIjQ7Miuvv8S+zdAQdEQ
YHa5u37QVbHk14s++GqfG93FgGp7ewvf8GSTlMHDRJEDqhKFTFRTlj93aSBKEK/PgFxwC4WKxgjq
/BEqZcU7RD4ALA1hSxsKeOYZgIgrUzVV+rNw+A4qUUybUmkqwHhzV/mXZ7DkYitggOfXggbCUFNy
/Ib7g7jmcvoSD+aXyKgS0AZX3GbBA341bZhsd25MfA3xwR+1hdhpVnzc/zenjULsRy5ej4MewHee
tDamEaK+G7NPh0EyxOtGOro1TM1XKPoRfNwhUMdlaKoslEaDBa9dPuzmMOAdxBB2LmyF1oVysuzk
RbHe+VzFj8+xuht/3Y9q7c7hQa8w8s8pGQE2FWY0u3ufFqKX8OJHRwWTAdrHy/lESLSxsXtgC0YR
J5j9j1f8gbySjWkWHHLXGdSBf3PKTy3qkZBsV4L+RfhYw00sfSoabPtiEr5ZMq/Yp9bLqDcQkCYt
not+sOV9UuUdkyOXDcljRvssrlz5WHeUyNSoBY2+dgbdE2Qu3uyyFZp1fe6LGXr5Hvor408lb9Pe
g0/TAwlEJXafPPHH70i5vPUkpOiZXzoJZ+y9lbYoDN/9DcITZN3O/XGf70yMuevW1Nni+RR4tdMY
lw5rjymtrw3RkoYvihqC0kizOO44WV2U0WK89rdXL4L4Iz7BMhN10Xb5I3d+9yS7JKk44TnLFlna
eNhgFQ8HpczRgfdnxS3errzhgj9EAvqod6+9kbLvT56ELfrx0MKAC8IgmpDjDiGtblVlR1upCuDj
Oq5FazPJry5K0h4MD76z/M9plDx0KXSAWs57sh+YF9OlXav+cMDxtLz9Moa/DUFzMLNak3BTRbVH
OsLygMapyqqBmKYt48cFQL9RZ7WTYIRQMngjVtTqObAkElegV/sRZ88+Tk0+7ANrtZbra+mAErwM
t7VvK7x1mS//2fjQT89BgKlEvxThz7nGWuNlB7Wlpzq/NqLK0CkBiPdNq13j/agd1dDZDedS6ffQ
YELkCfJXv2C3HGyf6AjlmAdx4Mogk8fyuj4GqGpeVji8Qb3+4yDUNjIGYwi6ju4mIGH34ZPGNaQi
PIKQhaWwxTfu2fEZtc66ZyASmFKZkUjxBE1zpGOUKEoVzUkV2QOwp9RzLE46NwIoATw7//ROTvok
z7NTIkWoioNXFOjsrzMWhJygEKwn6/7w4hgQCe6M8SmawtI2+6/O7vgBuI+ovYy4/jHRTWjm0oRc
nYdm07gIXkR4WFEbzx7gOdTFtFgg8x5/RLTUcG50aNtZOOqb3bvoTUMttIW+daFLEptum6FodYwj
jQe3k5V+YvGG/h9yUoJo/S/qqjWIGlez5whBk27vP+MMYVrTrZXzLNh7sUAVODtKltdz966ihyD5
JUgAPnTYmiPxhWUO8TEXj0zKrU9gV6kTRSXqKt2ma8YZmuG60KA/+/WJAzQiRNL+EDJ2EXjKf0Jn
/0ePt0coFj1YR4IOWlzc/bQH5bj1gW+9Ysa3oYeuqjSi6XS8pC/fMnIfu5++KEEZdDvLyTHzxp2v
GImRBQkKKu0ANC3sVANLzjK0GQrPG4+OfQDs0DFjF+Qc4b/KEM5vDt0/d1wb7D75S6sgbpiEsivS
6vpmnRwz8tY50ybobAVoYGlkD71t9D9gEjuxN1EE7AvPJrh07/ajlZNu1ohypo1jF1kNXwFQDVDr
j3oihYwkccqsKudUNEJW9GD0US3YddyOp0tGKCpt6nVc2oGkROG7wB1H3fqmHSSMBePM0HsGmo84
37qxqsMiAIKr8ARr6ar1zjia+exspB9TmLBGYyUxuRF4vT/UaJq+CCJxK3SDZEnyGTLJQ/0IZedJ
axDK8FU+gAC2Q1B51vZnU0Fjvh0YzfFRPr29LWg8IhJJW47E3YErVpZeJkpLWdsrpikAuoikXQua
P7RAH4gRHzdBy0WZHxKuzt3toj6yV5My0iSTchAGvRvmjqXE0HvNT2fhJDSJd4tp2TpoVu080YCt
qr/xqUMyTo6TsDMrLFbmzRXUynzOLO6LQx56LCWzQpb7zHY+4Zhkvk49BEeu19G1BNJNWnkzDwtp
GBuuoTeWEvSMfpg7ZVF+idzEAdIgexOllVxs205/hDcU11eVgeVw3Z7mbw3E+qft+bR+KiURjR1j
YDRDhpOz7hn1w34BVrB1hjb/N1Xys9dscSdCLOv1j/8KBXqxTBNdLZ/pChJTKNKHy+TljYvfRIN3
kG5w8t6+5dCQmehp8mBZvYwY2U8jzoXVH0qRpzDQ4hnf8AZ95TMnXyHkCeWvF1+skbaZluM7Ea8K
DEcLklCSfJlg4JxqTmXEk0m8QjwckUuRV1BIZsKdvT2c5D6vMWicmjwy7/TM+0Y5istua+RydTs1
dO+9qFJNw8Nms9U1Fu7nct1vtSjHEhRXNeQRY7IoA43YvU8UppNoeY/53i6i3CiA5oSDmDZAB5/d
BgoGzQBu04OKcF/AFV7UGC5A7AfJi+E5LP1j8414qNGz1BUTha9LZBLAOciG9wp9rF9+PCk0bQER
zl9RNgy+rzQEbFGRPJrZRisgVxVWVR7c6JR11HrLfGi2/rZ8iTLr+ESRd4VJchD55Zh1zWXpQMBi
RCroB2skX6q1ynxJOsqxgP6pmKQU9Z7Lvxa80WUjv5GMQdUfBVbyiNAPvuJM7KLi9Vyo5YckGQ7J
8kiGVj5C1+BxkUNBTARn+LkOPVUZKEG7pSe+YuORtFQ2SLJvZktCSD7e5ygU7BjWAbTAZzCKORnv
6VMt5ktPRYK/G+e9+6vlHICxPOLN4O94K2kvtDPJcx6z1I7IUFsT1Og0hdaxdfoVX5cbj5GVP+wu
CvRTkSbioCHbmHicbjnJU1rdeWXrMEaBbi78iq3kMeI3adYdiADnqgHyClbtEsUByJaOXjyQNJnk
2f/iiXg+EU3yWUexESfGskSDEfnTP5kVTHE8535/Ed+gSt+YI3wVx0GG+x1hbPcGFn/tNtcGs6rW
VZ2z3OtRDNIABAMLwulDKNi3wS5vDLN+pGPfUrlsfsiA1HI+gD3dsOlkd2QJQnc/yZnco7IanB1E
jffFBKsnQdQzZoaF8k0DhkvcR7bnbUBVz/FtykD3cWJ83MzMBn4YBjUx/PnCraLLdZ/uI/AJtId+
5ziUq7BcYdl2XChgmbyCwxR/NU6wM+lvzXsRIjpUJJDSiXKdZlisktilMg7B9PFm0wlOreZkSm9g
hmg2nr03hKdVmVbjmfDfIsNiRTF+U4fzcf9sOYOCk23AA44NWUV4Zln74HuzLOe6+HR9lUgwziy8
QZog+MrZsDYvkfnQN87i9vGa4CtSuJA4QE6B5HkRVnTAQFBwohnM+Wue7soBs9XEWwGIDTSEAC9x
WVq+2Vrfsrp9+ZjczUhQifNGLf8ScTiaQWixCt+8s8b99BPQFesRq1D6c9tUI/SH8FULiT+7Jd7m
7QANdwNSfXIN4bWgKFOpzMqajgMSoMM8cHrGGd+PU/LWyl39un8QB4yCPOgdqQrrnSAfT0jhAhkK
8eTJ3FyQeOfSmwBZCtZN13MTW91UZz8pewn+c2p/kkTHYwuGjuOucLKxEUAX1+J+oTk7SzYQfCTK
m1RzMLW8O5e7B2WFyhe+q8KBWO0Ua6zIy72xyFDa99g4gGHVWLMZhJI7CVF5SuImVtnmSXOczK4I
ivz8FzArVLiRHqa847dsnj4A2u8q10Av4pb6kaWx3V/S8ZId6ndKLtKtWug/w2qrg+EDcagxIUMK
5KtVo5OlvCriwIylKQw0IJgCc0DjEKFGjxMf0r8V7gL6FTLnnnNSlNM99hJEbDLZDJ+BQ4fMWE7c
w7//d6fcWG3moWAIopVtGnXi5favyqeYFvbxQy8N/T/XvXjmYSx6KGCiSO8xWKQub83QVwuzqNvc
2fCaKa+jYLyTumXh/sln+sLBT0jy0N787u909cZjFuk4npdXoU8mFYU+09wjQM4ZY0pd4Y7fikal
GnjaxkJHQP8eDt0gehl+vAzLzG8iHzOzZPGJUdHkHHkUDY2Crg10d4/n4F+oqOzkNZT91Po7NmGa
pYvn7ZHMB8S3WtuLz/9QzNq+C+I2ATRTv1I0VLZFksP4l6S8zB4d5Nc/yTrxTaqe/bN9T5jFomPQ
mFpvj2j43paMuaRX2+u5n6sDhXfFSffe0i8AD+/d4baOPvovIj0oKvz7dM2nFiLXDPXVkh1ygv3l
ZGSaaylQabTDQWzdMlxVUpdm8UW84B8k2JPrNwoRmepn+CwFYZu5+vByWKiQUSm7z2H8DyeVOUtP
JffZ8YqM3RdA8Q2TstI9d3WD64rlgjZPAepBp4eNSt8RRM8OIAtoXnHav37dbkRouy+goPq6PZFV
1D4ujWBbeml7XWgPuzKZbv7VXBXNLdT91FIHUPEwGLEVDLWqhSO0BeTIuAty+xNs1RbM9ACpDty3
GpRNWftrSaBXM/2uV98pCh7QkXtMgm2zZhaw0waqwsyBxMBYDh9kejXeoZh9QPKshJdazHeFULx8
dnQeKGUTdOg1cPgZ6yPAAM2za+IeSpJAwjfRd3IdIffex+i7ARZtyz9HZgwVgLZOFz37IlSHTBrK
49L5VxKO2B2XuWD/FN2EK0EhjFOmGoCskJ8xxMEqRPzO0EEgqagALdZiMIn47IICwNTFzqmsE26s
I5WWIXrhV2p78xRwLuaJP7lH7GcQUP498EeK/1zZuXoCgOq7lbwYs303QNEcKN0ip/YtF1D+PYYW
wisAUM+qwF/2fdrDdAkWASqc5quz6gA1OL0MLBOd4A9Q6aQ5JGZo+cUzmWCoSFAQNmlrQu/RLqsA
KIPmHSqKZ/vcvRm971xFZxbWBwZI6s5OH6KwWJCs/4eUQsL+bRwppSlpH0DFklsqaDmSc6EqDTDI
rcXztMOoSs/tuuRS9aRnKjeJ73Lyq44MxgVBykXlrUSFYKd0KoVbCIgDsqGyopLw9j+di6/7t9Vo
dFFJsgCRDuo8+H6487jStxWRa6uSabs+HiATXaOv8rPv3G9BuoQcMfg0rlWwL3B0DK12kMjbfkJ6
AVdnCCkDpiCymoWlPHkdw/doWP5aTC0pDHxSz9C2eBbd+gxdwNwdUzSbahEKmb88xafPTK39XZlm
g8nTMxB4a0EJ54fZPdlr17JaZlrcKvQHpXy1ZNXikvwA3Jp7gtbZOs33jlAPCUYl/gF3xkemBIJ3
nn3HGWp0HhSwUDWXdVGL3OEizb3WsThgjWLNVuv2e3ONoODcpFUxe/6DcCVVRcg9aVPwcf+jnfva
L7N+oabNFMYFUwsWy6Svj6fBbCl27uJsH/P0pswOZ22CAfwOszqRYxym8PlRyvHAOBNoUwpsX5fx
BELdAbKKnjc8OtWjrplZdpM5QWT0hapCeUmNUs+EJyUkS7YiPH0oWBOuggOZa1/1RF9J2nghv2Ho
h/0jWtqpN4nmDDRulbE4hmbCVFopc+s6IL1r8qjZPo/atwTKwkjIt/+sELd1zU2Rf3MgLBDQSyqw
qCm2Z3P3VCKS70Yg06x8v6IM5E6m0d7YQsO76T+ocT0HkLMpNha7st3sbbda0mXmEFKxnY9OAouo
ZfCPWEknVc+ZzKgZCT6TJPfOtUnN693yEnRRGAYid2w8uEdBLLU8FCVoATKcCoQVEm75XybpijVL
5kiVJEX9VI8bAiJ4q6hG26VxbOpltO5vYX/roAsY8dmTdCAuyUF1wtPS6lpyGi2AgNODukdV6n+k
V+vQBDKVxrG16OOiUSyexGMeZCTGJsErJPtQGChcr4PfMSPIrc/Lc3p7RDl0Vfxuy+VdLruazjNB
KSCQGZwHQnDaBE7Z9GgmnENmTnKwW5CbTLPrHQEQdogJXUy5p7gMrdMppYhIaCk/BanugjZioaHt
37oF8yx8j4U3aVMQ1C/Ho4C+eOvOrwsRyBkgtpKSuH0RNNboBNbr1NRGCaHGD4AHYUfQyY/cTvvx
4VgKEaxitTm2OdwKUJB/3HJLt9+Byq/lPASER7LwssDjpSK9i3Gb6K1NaCr6/F35BjXm0dBUW52d
NB2IQRHmXVlHFLJrhj2kVx/yFSbY+Mpdi0cckVfjnqBkRIfObTMroAqOy387c9zJ226uW9J96eTN
aUyovgbaEI1bjspL+kSmJCbAOQhuzcoOimJ1JRgryTGutTUfz6N7LPTi9wQilmwMXGv60nims6ct
CBT7CdC0QBLZlsyRlxS74Xsdj3R/sWTiUde3o2APqkY7M6YSx9TSZUbTamZdZ8cC3sUl7eLfqMOI
6Q/FAhgu5Tauf1QFOpKxj8nhPJ3WkoCEYky83jJGhU7OJ9gFNyneHIb+8II79U+7xcGBM9bMlN9/
G3kHLgNv7wDMfkkltX5dK/lx7W4FfaAnqwnr8TqDsbveFpxIS2rr7MeFSINm8lIVzuxCrGHZvaF/
lov8Opympmr2yRMZBBGjZWOp8r6J5QPIIfLW/cGlP2O31WnN8ZVJkwNQmFV3sva8F4S2IDnUYQmJ
LyJwjPXBdFQJqFKFSQD2iEmC7J2SHofBLA6SGon5FEZFxtas2HmGaBxqmQ8Y0+0O8JBjV2MdptR4
7iaas0IfwalgTgaQ1cGr2ZsnsOGvPbFvvMouxtGnrrFt1OOr2Vcc2TcMSq1HH8lYdfxGoa35reAY
5jDGxxAdE9hsqQCqSG2cLCaLKzDInSAEsiVrJP8cs5VXPYnaX072ASZrEf0YeTH5WekU18wVs5Nc
qYaYvtMvDT2Nb4UUuvguXazf8CxcfbyoLA3SPbU5qQmtbQvL1LoR6mAqBpt4RVoa2aKt7CLYtamk
R/qbDbFCdvn4DQ3vH0ZYah/jsCTNu8kx4vzkO4/rb+sVfARpJ2alhGZj82bx5NZwVwScPaoEUqGC
BsMkOMuHVV4xEl4JlMAzDfMlJaQ43al2pJDtuMqpMDQzhjt5nPiy9uoeRkA2i8p9b4rTKMZpZ3t4
dIBXaCX2wNPtBGrVVIKof3XzaO78ZbbsV3wdv8KNQKmRTdzCfoUFw7zGin+P6OOwZ4Fv7Txc2lcC
0XqTzOWC0M4HfXgHgR98gmFguqzCnmP7DMZuT5wArVSDLXMDibL9rhyiPjmarbgV2h1XP95mvi7t
6n7yV7ossedHKCF30nYIM4be1u5Anr+3SGtERtIHseVm60JpMkjhgIS3bagH+fv0XJxU9kocEBAF
WLWUl0zcnzDm60cqwx8t/htDDCB6n5apUW1Msea7w176wNWEiLEkr132SIbEmZ+5C6KMFIzTQ4mE
GODRN7/GTxoLq0kyee3xH+7dyTHS4LRB82q4AXRNQz7sOD9VfBILxlpfs79OVdKhjqZegROGkk2E
c7fj/fCmdMAlVdTmwmSFf+22lnUFYVwV791Wq+JDFyTumCki4Xn3M04f+HO3DnqmKn5kVcoOzpbZ
lgwTEgCjBEbcknd85+CbEfvVTqrKSUt17DkptPIJEgCAOei1LFmWC8ZcnADdQj6ZKVe4qYX6ZLWI
hAT53nDLB7d+GJYVMU71OakNjbeZ2oq7DmDow1HGc+eTZRGzyNg6QTSNfU+4sQCxXqg+9EQ+qxLU
CHBtYHiTqwF31p5ZLi4xnrf29Fos3BfrSYP91eHDJMNoPJPZwQ7jpfKdq9ItlJRokhW7g2XOvs9e
beQFyn4KmKnyq+tegHQ5+vIrl08P3Ay4f3x7shF4gIxeDrIJY6SOWLlNKnsZ9x4DRVhw31uSRB+d
4qTewmr4KMmxnU0gqEJ4qnaF0SzPw1zUs33Hvep3uKWd1sOqgfUxbxo9peldViygmvlmtl8gH2g2
vryWcBESPeTOeDfI/byg1BdNHaLhatCtCkan4LCsj8AGukXGpQzt+WuOew5k5KUWIy3S8Hh2miiO
7Rob6EcPqD2Uqw4lt/iMPDMQkWy4NVvg+vp8wOGZxI8iRPhRSOuWm8Bb3WXBatHruT4q2p+N+Yb0
q7sShXXvggJVcBPmUdSV9yuiNtLFFwsA8/JuaDnqT+i2P/pAQX0RzkQOBirRgdIvPWb9G0zDsYtA
3tqyyZvp9zaMHtjJyFcPjav9o5K7ukPyhsxLKiZuoQyMeKpJVK8u/TUtUzbJzfw0HV21KRdaE5Uz
XrA+uK5Wg0o67jenUXT7nY5Ir+nsOflp3moU1ZQoI+ZMm3EEy6L0HEpDzc4BK7uC4ANS3jJEQ0gC
juyseR5E6x0QmgRTGyUsJ28ACTtmDa7I3tSXtAya7cZTE3R9M0Y16kqUUC4yY1Y1C5nNbZltleD/
4n5mJ2JyxlsUe8TbysaJt1dlFQGtMves5idZf9cKkbHwjarEwJx0ydYZVlYQwCK3ufpaxddZVL7U
209UJANKiuXqhevbrUWEJPVdrE6X1iZly4YDUfUQTybUgLo3UXWwMj7Eg/EkJFAoYuyuyHRP0XGA
EZT1pe/kPv0LpggQlTttVJL2A0JELeeX/Vu7IPWkQ0pgSH0r8/N3WHiNb/SiiblA7N1MNxy+EfED
OX4//FEEVsfkGD6BhCIG759OkLGCUg03OyKO7qFJ1Ok46knCfMfowVjETvN4tbhiEJpgKp0ADK3z
G8mYX0R547yRLCiJF0c91aBBoc/btJlipY/JaoMB1Vy/BEN3RQNfCntZ5Pf2hoWKApAJbLXMcr4U
//p1+BNfH1ac7FH/2cOrR6/8DfPwtC74qjXF2KAT7KtSC/bwDkLa7aAIcJwKq77nnH8oXnlUJqkA
/IyrEy4gjqDaQFKz8jsf1zr1/QbBX2CWaA2cU396ADgB339TRmsjXWK2Zj0jG0UjzsfRYxpChB8j
JsHdLqMWnUAU9OZb2Ong+4RpSHEAUBwEoaa+jTnnG3e4p4jFNsGPI47DGNuBZT5S3ZW3VpESvUP3
SaUd4I5wUdUmuzzb04JrejAlgFrI6YKck+XlsSoXqPzX0wRrU72nXeYRPIl1LxiUKKVJ+TvpOEj5
qz1xEGFZGvbmIny704Rx2oOJDJfoXDzvSuJ1QXophhHnNmFvUh17/ZuOLP62BmEqX/Kuzy7WN0F2
ZFID4OpD6MVW4HnCTGt+9pyisaidyX1H/TF+DKx04OaIq6idR9YOZr0EYC0q9Gk/ZD2063yZMwIN
FOvo6F1e1BNF4D3PjhlhTybqhkrnTJ2aAXRGnw2HnVBMhM3oDYPj7JlNXXAJGzqlj0iU3/jRZRs4
VurVC650y9cGqcX1TNsabcmCTJboL0H2RFdFTw24EI8ZxctOgNsTfuiUsM+hYNX16uExnhRtepGn
2RHSuKJR+sjpZ6HRtOQ++rwyMuTJguP2Z1IFyup/eMvzAN+w5FqpmOpcgDTdoaUq/CjqFIHMTLtB
dn70YvSeoXYcr/ckKqi4q1h16D7BNVWYinJaVV1YP82c7NyXlGygj8iY+lTyQTzr2LHY2H7HQioz
z6MSP57LOAaRwnVnW3X0FR8gmUwCAsEjCbazm/jujGydTnVkwlP63IOsEiN7sLwkDylWKuzu/Lly
pW55hakQH57anIg/jogTTEHgrTOjkbKj6kvVR1MOrfZ1e9ifun8VHu80YbzmqWmXiktVVxUdd0/Z
2tjMoMHAjvsWzO6RzIwkGHF0pK1nnyBCEJt6Sj6SkYJZaT0Egk/8BalQqAtxKeNA5bPG8K0+M59q
zbWtLTl04q/C2i0MWctXYNVFSVVVljn/MgE8XkQafU99bhqo/NIxzIjNqO73iA2vLIRbrOIzauAr
6JeX0jeE7Cd7610kPdbYC29MmySTjNiYg6dqE8deeH1D3qQS3oeoO6wwF1SJnb/Ke4Eotawd7KDL
HzwKMy9kOcjkifaPgP7bg7J/zCMKdKUYqbSNp8ad91LyxDj2A1r2xQmnORMjplsRx3rBKx2xhuio
uX1gNYSiNm6L93OJ8bgPgmGoh+3OC7OpckjQAEjoXvipQpj/wfI6G6zOgCcZ7HEo3AoohP5aKocv
z/pC1EhlBBBEyCffHf9WWbbXfgwmBF2dyc2MTlrqcNOCne3aFjNd2f2pvKqJLjCfPxy6TqchpMbY
Vcb66OYM5JDgySoK//G/fHSOVTTjRJysiQpOamR9l1uNT+MOTCHD8NhgXQ6o74jsaDWJtEvviE4o
GunPX7WKG0gmM7sgYHLXjjAmNjjQScB0KBjll9k663ooAAp0rkLV2EY4uSibzxBFVGGtpssxZEDg
TXW2Hz/p8IhSa7+u8u+YVIWpQEqOO3XaKqIWPpC/VbrnhXYyFr43PQWESMg/4tVcRCRUPM6mwKBX
WOd8UlqeJTlnJeBfm1gpK0aqMHjx/IGzdEdwbaIj8omneyB6ml6h2ELYueZWRgo2MzFFWTBd2LcS
HKewL6T/MVUfLyKF/+1r63RMNCS+jt/bBMKPR7tHJ6CB1JLJ9xNzHWPpE73DnrituDAWArXApn7P
XacmBVJmYR0COJZ2Y+0LbyvtEpva2Fv6cA4kY1aE0IOLttyUKLnkignXjgRTw+FT5D79fJWVdRzA
l4JdGS01W02Wy8icuTAuMfBg3foiVCn+du+LYZU+UJtymWdQcl9ZLZNzDO3x+U06iIffOmV/qI7N
2hNNL3+RDoiM61mjC6pnLXrdj3IJ7AhS6tN+X2sdz16L7Y7bc3eFet3lWy6TPZx2dPMVpV6x/fe1
ZKYI/r2ZwAkl29dM31C8UVNQRuQVj+pRacDuo2tnnMvbYVXkRLomNEZwKbK+O+PnGZx7cqKAly/7
qmeb9ggCglC6ydYjK3AG/PyOT6U8Rk3eG4kWVJYatYMe0pVPtHVXfpdEibQ7lkOXr21iMJKS6kxt
svGpqab0ResDwZ4xP9m9H4XTvwAW5hhl4xoTnUe3ryed6TD5TKyxsjJzQD5MfSdjHfns/WRxCV7o
jFHWR8h3QFE9KZp7elZ7Xs3vM3TYRlSN4fw/E3UFuAtDesbQjqX1xyCkhBxEYrrxtrk63jp95fNE
vLl5N5r3o9QsZXt537oPvU5Sc0E7hLREWeR0N9+rqAejYmeBJGktY2qGYHOhB0MAfczfS1CNi2qA
/BxEJhEhK/KOv0UAZweADlrsXLlPxugQjZBGZ/5aO/Jhi/ldZUUHNGJO2DHCJMM7JmCX0+LDHhgN
WTKkDLJdmQRxmahaDrnP/BdZ6hDOeZbQ6wYWmiuR1XqG4rl+U+ziYlF08WLKzEcXTeEixpE8j9wE
Zh2tuA6pHSAIEODwkke/Uv1MqN7jpStZJVQwDKFs+AFasCBijC7udnY6k/ukhX9tXLz9HNoIO9nF
8DxkbZVnn76N4T9Z9J93J5VcH+JFtOFwVnGLAMR33CLZfWC4llTPkcNLVuAFqzG/JQrqAzrTtbAV
AryOggWen2BrhB85bQzi7KCdrTQOpYXcGVqnYcpuLfaYBJaJAKkLhvzKLtB/9hCq381Me5xYz3xH
Cp45pYFcXA3hT7WbySBdSdKbdOP0DnP8bV+XKymU/Jt1xtSWmmZl6hbcNH7YathY4RfvbGi7wFJP
3xIwzkuVDV2nstpixXPDZSnqh4D5GI2CPceQOpI1Ri4tb17uyFvKTJqSVTOi26wULbn9emR6j9wL
ZCf8uFr6oqI9QhRm3vtqHyCZyZlEUFbsnaCzWOAKaYYu/yGX4vOiN2/S/brWocESQeM+HvSeuz7j
3Gi9suH3m+QLTvG2zaWPLyxlJbt0cwIQU9dk8yexG1aFcw4BeFTGo45xHRHq1rKfTvCnSaEFpYwi
iv3z1+YFwxhdWEqrS6oqxojY6EoAfhVM52SK971VNkvHJ5t3Ms+zn7DihhQx5Iw7L0X6VDkGs5M7
ITPP3e8lntF0dWVXs6zGXk/MrWBykRmerxPVM6/uLXUILyJv86GB0k6FO54bxvjHCUyMxXMfrcM7
FTakm0GerzvDVTtDS7xwL5WMmnq4BLX3ph91DL1hfeowWsGNVKz11BuEq9uXvF7Ghx9rx5nQkhB2
Liv9YJR36u6URVkkPYYCyHJiQTbCs2SOSaUfwa3mARwvUEgDOfbXGoM3IJwsKGu5LgqvGE3PDUPE
bUQHWPGYHajpUxOeGDKp8RBO8NiWdaHB6qEALsxva7bOTU67OJF3ZOkNkrJ59ymUaOrn6c1uCgbo
pee17vt/Zcyp5Uj9UkzT2pretQotI4EbIBSa8995fsTPEsF9fi1J4RDCDa7TkRkVkWY22PQ0Oz5l
jabgqKt+EAxqATGWtMSbr/zoiO5bli+m+e+5JHlwehFyw+OHiGNwcJQl1Fupwu27j272ai8TLqVz
0PXatZw3aH6koAgBngRE0hT8TEvTGQUHIJAIXGVZPH+QqS6sndT17hTcS4RasZIGKz0v2xvwOpbc
M/1Ualbl2p1wdTK/yafHFT45znN55sVDOBux7jiTqbX2wI4C9eT1RtPRU0INKiRk84zxt5TifnyJ
gwT/bsYZTz6YFWJhIUhP3D/bYrgqJsslBgWGxSSBOZrBhO1nCz8j5XfsnzU3oV3ahjYmJ88QJhaA
E4TaqEwE8HhXF657pqolC5BEXEr4qeXZx/nES8yZNX39ew8plBnN7MYeMde/wb2e94c1u5B+Ir7j
eVO9hcvK4LpYB/w5ataDaru2GyIWbzr/zGrjpofifa4+7QfOf8eTqIi2S7s/+Fhs0FtxB/qww15H
xEEQBVYBWP8Gr2aUkfx1vkro85cG+/KOyldcG+cFZpY+P5fd2dG8UOZGxeBPBdKS2awFxWgPM3te
earlUts8gwj1VhzEcm0X2NvV8cmLNAnJN68iKUTEzm9JlYp6b9YUN132vQjIW2XVHWJa1U7eivpk
vCv6vAQfY9p8l1pLgrcboV4uavtoDao5GjqKGjEEyGEz1LO3Bh7uy2KgbvXoSv4ZxjquYamDTbqX
O3T9epRatDOwlKdT3KsDzvDkt8GrCn2MnriUo9dXrgEcH8ielLlfQQTzJovW7QgBlPEqA8suYCwO
cucPDTFB2Wa7mQFZW5ZIHhiGFwc0BoUQpDocMMqsg9+aEe1XWAN5IY7R7Yh2pp4lQGmqEc3kmdsO
vd0EwFsyov6aPggzTEwLPaX8lbK6H1XiP90I2tj+8jRmwIFwGF9dQqn/CIiGZQQLNihRChDv7MYV
xBqPi36eFUGf9vlAifnH1L4Eq/TQp76CujHpN4ZXhiQN1yRAUWVC/l5URcUUYZmDtDd+mf6789Pv
WqCY5ZnMzQlemGEg5Mazna8Cbimqsudfh2yzTOZzfeY74dlipgOy1/6ibBr6ySLSXzpKRAJA89H9
SaMQLhpHvAOYBPa9FSYXMapxMXRTLoSaaZaZbuDqlFZnUXKdPoPqiZWkQsD4EPtIxVXIVvqVBAzy
e7fNG+tFktWkSbJsKb548v42k7QG05Dn08efBvT1e0DRzih5LhBZczj7rJiC7wdUwEhpSlGWSOA7
ZSCOTxkzXzsjvAKHWiOUefddQWqPiaUr25MLLUE8nec/+SwFnkUJxgbjhVETLj7zvxKYcx4HhKl+
dSTnciKk4oiyjO8jcIptXPEiAgVOW8gdbYizCw4NXUsL/GS3Ef4bheAAFMmGeCqigIl+gerPJXlR
XuTPq9dz+srPeKNfzAfZI3iD/g2350Lo/qW7r7jgqZDbGAejgvFzK553YEf4MmfO0g1Ncyucn2tr
rVVsPlR9GPofcCJY3BPVgt284bakEN1EjSeY+AISmxApjGIjEAwyZflYz8f0QZHxBNYPJFyzL5zV
AGbgC7J8qwwBuS2doS+/XBxC4C2uYfKcb2lknFTM73Oe2+2DB8/jZ7AevdMOH7gzbOjOtR98RE2i
msza0RQXGuOnf+GIA7DKSx1qPWC3TwO5VdYUdtQz68wTBywdwdVYNTMnO6jS/uNnV8+p7al8DRm7
48vVxs59eic2wBJMmMMJGhUNdo/PBlL3bO+4SqLq7mQlMXSyulmVJKumDkEFHmv06tDlHQVK7ZAP
/0Qw1Ecw3D2htmHssikAkqCtZRxwpGqca7crtfSN+IzErECr/yjsrB+sIQSNIX4om+ghR/0uXmnd
qizHX4ACa5fqzp3/u8t1lRal4BtM4LV/loJ6cEDuw+rjSWNUXwAuL9rlQEnADYC5DRGYm6sgL8dV
gLCKFutymsm3hZG7/4NGUzikunZj3++G+mTeB3JkbnK2PbwPFooUqv7I0yyVATBkPimw7kHZbGZg
vPRTdsEt6tBROQOBuqrziiHw0bCcISuFUuMjec2xPQqRit1yNh+JD+E4OH/OnR6rUMMmevixHBRd
qPr3ewk4Ijflif/BQQIOBQ4gNQJaZsttOGUniOBShguG3TBDtb1dXG8xXK5SWiB9HgdRxx40BK+Y
rY0KtQYbCjnmu4P5+v0UQcMPbmie9dfwxKjGUaA5MYOx9+82ncpcNPWYOlr3pPRXL0BVj9VAKKJT
fkI60BT9EiRgNnEwcTbasJyP4UREtIk/TrZiXDiS9PWA4o8FOOTdZpoWpLpPVVtwqZJ+2LMwiQuo
Pe9Tf77yov/pwuxiGbjgGqW8oZK++g3QFQE27yG2RA3MN+wozzplM8Il6WSEQt9E1DAmft/vxHH7
cBjrTgY0DlRSy+pxRBgLaDZgpiMsALEeegZ8wNQb28a1F15G2ZHGlsezEy4dHOuIcnD9O2EUmaax
2zSNKFYsDea5GHPJPA/bicKKYNEAxDln0XzYKeGoVBBo3DQ2+Na5EGcfJc3ei4Nb22FrnJ36e2If
O5OPC7yoB3lUAEEzVpOAR4PGoOH3vVBbdvVO64+yvGSaOmMPUtJnSd81EOdcwQC+a/hqmfGIbNGK
G74rSseVaDebc+zmSnZEvKonHmFh32iscs32k3i0qZEO2pzGF+m2AScpIwHxzMV85f7MzpME0s7U
Ue2Igx3ZFmAvqZ/mRt+eKOLT6ZfuW8YsizmfCsnawCqo/c/25Z0OHWahCf/nyOCHu+bty/1GFCU9
gbO6dWibSxX6NPEdohDtwvsp1F5n3YUxsiFBMdrNcK8dOzlaX5j50rofVsrndFMcNmCwlaUYNV+w
6/jDzAFtyIquIZeHQAdHzW4JucXvPmZMCliSL8LZDMSn9Bz5AKLGsYK0p4edyHIOjCY8NEyXpTvq
az1KYCp11uUnvVSz2Dd7vbHdGgZb6xEnbGgT4sioktwYJgeJggS6jVReET+ZUlq6Oj9R0PalQaXR
5x6Obdm7Y82YuALNFXspVICz9lqAyyKS+FZ63Z9iTURWS9kcvkdq+dlVlMRWWsWWjRSM4q9mFmJu
3e/yiTr7Qzi4xl64eA0262c807AU3kLBnnqR/rigEd7mGX1SHt5h5IkWljy+5EgC8BouOLItxU7V
Osbt1yAjSjnF81zuVs9+VgAJMJYsoW8Cxx4vGie9bv4yu48O8PXbtWg4iF4Vz559N0Bdw0PolGP6
SadalVE+DIt+ZJzRhMsZe8JqScJ4lInNhlv3LoAHiYz142TWJVgqcZBlvi/qxa+l+53Jd/TULuz8
mXjobvhqWs3XQceCeT40JSvutAWIMdXZbKAHOEoceRvt17JBTWrVRLBmPFxUT37p1ByGCokedAWA
kJCWwMFZ7G7/D6sB6rca/tdP3Xrcb2GBfPa6RS18/7LLB2je2wv5IpYcLctpwinyNlpqNxfPrhS7
0J/mk+lwbfwmi0PV9LeRwBTtBIYUNsaKJ2V2V+3GNH57o5j1C60YDNs14i7I2Xk5vxGfZZqyxVJP
Y6rLlSEP1uM5Kq+wbnS5iTpzljYXjGXVpUU9XkCJyfIf1DCJc/7u3urqm+cPJQ3C3alGCL/2Yk78
T0/o1dRK7Mf5l1EF8xX6LIqHMFyIXISRpwe+Od15Sw2b7la4Yk/XJpzyCZpchugTTZHdsou15d0d
guNaGL6OuZp40+oHhspKY9xfQI7niJX8rvlnxH46YQrViOWsiPstUNFbMR59oCfpOkAl14Omwv+k
PmLgc+3FZy4CBYY7R17xQ9op/GOwPhZ6boFqefoNg5q+PKIdScENN3IcEfctN3yJSwXsl5HT6Zfi
rRbPgyWU03VaNu97uheM2vDMSIoTKbEf+YBIgg8ld+VeqWKSn/RBbKdAIuk+LZSGBZbwqQqicKsi
LRL1Ev3Z8uClu+mJ+zepbGQE50eDAriFN3U6arXSD8KnV44KSLupPZ3zdK31Z6Idn8ePKYboNUgA
HMxXEabBHNBt/tWTNNSjPsr7wmP4U8uN7q5YchEYNYiLCtWI+5iui0B1mB57Zh6dJ4Gw9ekGfDqL
4iBP9lb/Vd/k6uNv7fe5RgInXqq9sJfqVpFVwfmu3uwoae9ERuW57zQ4bn+NFVi49C8+LK77Exqj
fZf03t1MH9VI0U/gQ6nzdoDc38AVpDuZf0GgUBoMOeUJwWqQRROuIlooegzwgVLWWchreeth4YFf
teQOauzyWvywA6gZ5CBk4zeRa3erF40/ukSxcDCc0CPlJmnI17YrYP4oQIDGn/qITjMyGIUlTUNz
osmKdxDdupRfvLftiw1eQs0NzD1H5SZ31TsM3WiufJq1cWxAGXpnMWayXTZTjvu6KyuQmX64lP7L
843GRJSHtEkLDTbn8O2XOyPUDr+edp5GuGcey7Qx0kQ0OCsa4mFc/U5QI2FM5rnQamvt8+LrpMBW
njQK+VZmMxEOk+pzcmae/c8tasu5qu/EFaUZL2mUqFcinoAGgWDNyE+o+zrJ1jKkp9oLaem0IiZK
G8vncALBb4LXEz5YsWCPtsDTMI9CmI6/u5L6SnuKxbIklf0zF/QsBETHty5+G2sP27h/jyqNwGhG
TOWL2tnGpG2wXnVlZRX4jdEZOGVB/W4+r+n/AWNTceQtLULjePi20J8FR/Cs7WUXPkEu7HlA0kb5
pvULg0a9087L7Ph/BK2S4eISdFtzCc+peBLIcvgInNdSWPWNW/fqDuQSENtWWgMp6TUQItXg2bL/
YWA1WRuzGTSLENTMLK4AH/t0UTyI7/3Znp49Abdt7qy1cQKVa5toDALddxcch3HSCoXKCWcLzltN
XN82MyRf4KqdjiFCdltHdDjzXf0dmBF0QRT7T2osfplm36l5eGMVmKrHIlCzf3MoFWEjKPf76yKg
odFHZlofLKWd8A0BN8F+z5Dx/JeH4lr0NUlyOMJaJ2IP/fzzx0dP+O30V0aHQ2DRK10ItWBgRJ9w
m9XcBETycQFCswvtyYA89XmfGyJBkg4LkO0JDwHHx4DqT+RzZSW6cQo5GPfCYk7UQvZ6OwNLpnz3
RhCDjHeDn9JZ8MnV1ZDRpuWbNbgFU+USelTV6RqNilOLxPzHnJ8JB/mxb4mMs4yaKedRdTgd2mG8
LSrAx7qDDfyAZczoGqzftN+RA10QVgWFs/usC1GlKlVUal9S5H2rpkyqx+gwvofVAX/pEe4WnGD9
lsngBHGlDyzuML9KoXb7JoBSnWykNqY9S+SVDhubZxJ3zmcYZ9SL1EECPgWEkR+ZvuXeTppCYmsK
eUTwypY4Bb8NlKeNoeINLm/apePXeKFijZyQVbxRxmbvS9DFkj/WQ5ZGykNBvKHTBCFz4H/mpAmH
eHoXnjPEkuaY/8A5JSWYpMzU7Sp4vZyueOFmgZHeGFosXRjZGWTZ6ycIKxerjjmSF7AzlJGQ0xWm
ymtwDWiPisnSFZynK23KQH0qDR7S+XjAnIpEXLwGa/EwPi5lv0FxqDBwK/D+73XQKQchp8jXW4HV
OoTcJHMkHhUpbcBWT9iKHhwAvRq7EB+uH5vyvw4hV99gu1tF6MUuuk+YOBiKx9rJ0HzxQAVcYxE2
YJbm5yOValD8+im9EhPweX+W86c4tCqlAduMRibUv6bHUXx0ne5X1lrA+i3cz01d9k3BpZuR6lNI
5ghaLiw3zHR99PkPu7ghl7YqIUyK0EUTpZQJG+Yu+UKtK8bT+kIPZEAs78fKhvzpkcOIkcnkYWTt
YzsUWbbAS/ZGViriwlMFGR0mHwSfBhcmHadOBIKx9x1xodVbaZiXUqBKFE6CJpFmdlgGkCSroLqR
yALviZqUACat4HzIy9MJkZivgasSuBj3hBQyjUVqfNXGKr6xG00gcY0GiItWwl4k+KPjoqrlXEYV
NJjC/ZeALNssK8LrgzyPaL/y7RQUkroVICiOncQfwwP1Z2eFe77OchJAVXD2lFTW7BaIherdxCty
vagyz2Fx9xleRbZPD2KLpcinDZY167FnLl744FW/P2BLv0ZsR/wv0n/CTVED3OHtIx2T9ueYueSL
J1iLgoWt63fQoOYRDkAn1tTRxOaNuSgsgyPkau49raMb5y34GrcIqH0pY8BvFq6qU7F7l8qtWEn1
5z/guq76b3f5/5YIeNX7TffYXe4ixI7EF/DP04+cB0jQls5O+bapZ78pQ8dXcp8FTmiBUgU+cn1y
M1BsYvxUbBVDWi2MzjgSKlBKoJCVVR6uZQNKGbLP8dQnNHr/c7x6EqSdapp6i0BCvLZaorYzJnt4
uMWOtKYyDPhRHER6UpAS0/s0/RFGDisgkY38KoS5AopaFjcTGvmJ/JeH1oQnplUO4yxfIVU51ScT
vEeO/EOi/bKkNoI/87p/0KL3v1rMHwpTdsHRF8Cb0OP7wXtPSdWtrszpsCgHOPR/digBAtWHbC8G
UWMcYAJf7Y80jLKwBcYfMnBOsVmJqQ1poQg7o7MFnK8ZfMWGypdUG+l41sTh4EauR81azdyGN98J
Wmr6TzMAdDxe3SjuBUHCrprNf/An3+yjLLpsHbqYt1cMicwloa7JOEOZocZqOKHhr5ZgjHwh3A17
0x1abwTToHVNmiOx8rzOmjNK7I5KGnSlZ/2NEdUSoyyeLo+VA9CtB1dHzRAiW2FC7ckGmlac4OrS
Jrk4grW0CeFpMNQSQpuB3TxdY/VnIt43/ABee2LfmcBqWNa3M0GaQ1OxUTjQ6GCw9mHxTcxZ5lwd
1zzQz7gJwo/EKRyqDhwsN03XuNWGBJzxrkW1aefxAnU5wtvgOKP2VH+ITrJC7m3G0PFb14qX4NBn
Y6z6tP4MGArgwDays+xRZCXXhXDseOIyCT4IcHeGCb9mqURmoQgqWVl3uBoVVSD6XfwVbcEPwth1
jnv+kTr1B8d5WUUNyN8NBv5McRQ7aU3763KV2qBYcKXkU74kEfa1LgTQiUbbIGN759UYa66r/wOq
Kh+pE8TnzZXNsp58rm1q5l6MoGe8rdcC8fac43fP+B9CXBkoSurj666ipPSbl0XKlTlq1iZjikhN
KvPt5+IcOWycfDQX29eGEObWKbFGi1V/oh7bkS4CbvLIUc/w/0HR9v11bKEfheg1FY//0KgKqoqI
uqulHvVE0IhpQbLnLdsitpqCbU2pRM/j/elhC2uUnRvjUGGVfLlf0LXZ9wIYuV0624QUYDF8fxtD
Ia68Q5dwCuU6necr2F7QQ/1WggBGUi2oQQefVJbCnUHF8AlsUvNB/DpEsG3InX8/lgDwwF/kQjuE
nmztKt4GgbTvu4uqu+36lkC/Z6JBbUZi3uB90ZOu3DHOFTX6mb0ofCPU5i18ssQC64FBKfPmkzzH
vpB3DkTLn68quTDXmKOSFeP/CFGc+bMMWQtHNWOee6d8sD3QmuaI6faz9TZR27Myag4SmoAipDks
zM2AMnAeGysMRrl3m7Hbs8+sgVoqG7yBtX7vDm5mu9d6aIO9iUPSxpSomVZKUPDelEMQRA0wdWnz
33394BID7ClZUrKlPeZl2JR2N0jMKRAkde02lKjyffo8Qwgb4aye3nn7hJFCzUo3aLRbYFuAbl5k
GbLXbR5gMyXMP8BUcHq8JnBadHPx69txBFGFRhxAOqDd6NFrICwieSdNmV7Ydau/NtFtIdqqbvCM
XwVj+qqr6aRBcf3bCdK7hLi/1yBWbRCZ6QQudwLl514dtRzJzDhaAPUjthCZ4jpIRdVbAXvLWUqm
i5IHVwJseY41KUVb+6vz+ACkEVyTXfnvbNWnAjYxsZNT4Q8JnBYPXAwhr++6KASKgWTI5g1BfDDz
q5CgwauLQ4TeVbwt6+qcAEFwJLZ8xhz/HqQFaSk1VAiVuTSkgvFpXi4qei/PQp7/LLpOYO68PhF5
BNG54cGtaL+xETqN8hoGelIrfuhMmYE/LfO4fVMkaVbZHaiBfrccifaxMBFMhCR7VrstzGonDzLL
k7c9/Ejv4Gq390gnSuoAVNz9iGuSw1P2Mr7wjIow5zYZw1TD7Lw3x1/EUPAvEKRegnsHnKHI9ex3
J8rxA+jao9qoqlxc132fgh1D0iYcUokDNtcSF4DCv0md1VH9qvchCA28713qcTxrpHaf1ELH3OIv
/4oQw+p2Kz7B2aJLHmLjE+xlWNI9EJP9NTjmSdHxQopq2JQBq0w8g7lhGzzJnaSRruPq7yyllA1P
tKBC87gLKMMdpx7Q3pYQQK/DfVU7ClvJXexNNtPX8je4O1yU7iH8QZTrIklP9d9NIttKNoYTtiJs
MDlpQmXuDGpu0VUDQfTO0grAl7yNkUM/NBpDwzyfaEI3bTB4J7xuoq5vDbKXYbByu73MzA00yGPf
4xNhlCDQhf+TDeclC0II+OYGZdGOoJlc5HiuSr75LyzYNeEJIomoCcBrti2mu44Qfw0Tr2arXrUW
XOK/ZiTz7CPTzsfgfs4zRMHiGgfrr1kLh9svXxgxBYLvGk3MHIPhsgpbJ1UbOfBmACH17v1UI9D2
4JBDtlBVpwtJy6Mk+nC19AlG9SCArMTnM/utHP+gV9S7zRe2jPe+s4srv6/9S7Ge5wt62gvX3XGI
Lod2JiG3RQSTZ0FMr3RN1tZF5BEsGTTob7ItAUkqstARU2ZEl2uMkOUIwWLvl7XWvY+n8zM+mSKT
5wVObKqqHHpEsfhRj582j3rf7rXqiCx6J4+P7DLjDdytNjkUd09w1IH12cv1QWN6rHjz2zAmrXzL
GEpf7/6D1VJnOh3N+EYJ96C+hTf4dzVbKA8bs6Fq2d+/QA7oJdRTDzMDTLGJp6ehashz+ezsgR92
WF7NKWCYa1CrDrsNWx2FKA2DslYjh4Suvd8VsH3fC4vC+EmRGgeGpRPMCUb29AmISMcDmNEUSZO/
NYwEbyvgMLg7cRyvZAUj4dfOR+DZEnB4Tslp6RbQf9IcCLJLKfVbhx3jiRPBk72roJv8FMBp6O5m
ycvuLPbEy0ohhtW4/xA0BptJ7ksDxF9i+M6tJxa9XvyXL0Xlr7y6zY01oGeUMKlL+ets9yvcY8lz
pb1H6W3TZh0J0ucoxB8s2m4i0GnwItAzESfXMa7EcrgWw81desPmiu4prb4oXeJ7yrVn16fvnrvn
lsRQfxEhfMqGk6wckCU6jHpiuy6wCh81RcxMsRnA6oRXQHg8rlxNkT4cC+MLgT8pLKLvALc3pS6C
zl+bizPKMEfHUtvtFuzon/HFwWK66uYtYRylEp/BOAo/JRGiTURK/LjTSlxvR0hK3yU7OvbmJR6J
qN6lsSVTbY0gbtaq5FtHF6ARNs2th7PJQ4FLfmbseWfin2v7Hv6+iQkTnG6DnrIgnk9lbS1ETHdN
ZI8YDnGItnPuZTKZyFT4zOdxm3jgkKUQJwuxtjr7ZppYmQ1rO8lzI6tcdsRERxZlESUFOlzNfrya
hJUiF3gwunSVIzetSKtipr68K+A1oQHZfZpNvIKLj+yB1hMTzJ7lUR9kXbYDaVqhANlDYmWvrCoZ
OaI13ngi15XceDjALAZ9n2E4Bb/rJpEN9ORuw6uX2UmAi9DEwpUc5VJdzK24lwnmGDDd5qYsLvB/
WEOQVy7ak8HY4zu6G9KLoIL05jKrpRqk8Ysu5PlWw7vkesOiHeyLS34MAIRzXJ15qUtHeuJSK1dX
k2OzLxuSZ4W4MVpSAcUDWZ2Ssu29vvEOI+KInJFl5ivrx0DFaUW3Jlv+FtHGectQop0ZXNVhG2v2
+pGFCNBBYkM507M7t1LSE5eU7QMpa5/Whd2+eAwS2KAE2OHOupxOQVGyicRfUYmoVfkINC2+ZY3/
MfSo0msiO8iHfHXpC9jIrEw1o3e6YkT8rG6b3d1tw6z7kuXZSGrpXh0f+zwquku4Tk0bbZV3rvIW
569pKvixTPUPFWXtJm8F2WTWPl5mzL/rHZseTrFPUgPwHS43WzD1paClrLavdvNEdZFuv1YJ/LjO
MFodpGT2aCDkiHB7YkrAEELtyMcsyC6rF7X4iAcuvJIfxhozX3EkWAP+pjUfdo1QfHZskbyLoEwV
9B0Yy5/i7IdnM3JkJXXooLuyTFO0yfTv+IH5fPPtchjDpspdoNrUbzFvnb8vdaX1/9b7VvlSkW2h
27/DRm4CuTRb+5Ozjo8p0hMCIzgNVq3pbf3kOW37+N/kw688gbwlG6di77d/giKKhvko5XfPrPYn
NQzVZy0rlwyTXDcg4zDNEU1k/Nh3bufncMsvy4hNzUBZLrXR4Qt0REDxCXJ3X7J7xW0eZ7PBuVg1
ih1MjFyspu77TEicsNI/ZVhnf/1tMRoSpjhpINReCtiMLsWY3+JWWyRhoZxyy7bobjar3wSZgNTw
n5nyY/1Qv+8TLqwTeu8Dg2gKkB2saUtTkKycRnM/3QgbNc/Lun71KS+Vmlqh+XpJdDqV8DSEBM8d
RP64irPxS55+g2me+tUfwTUxJTj+2lO9nYHAmP7Nz9uK646O+HXlLbpZbBheW6eFBE3bWPLMlySu
gAXbuC4CBXg4f4GHzuFUQ6RTb3I4XXOH7ewyL/R/WjdSZSr5XgsYv+2SWWyopCjwKtQMzcuLVhPN
CjkvG6vP3gLgp/zYthiWhqhO7OTMtG82Ah3pPnl5oAVT2/wSA+ozrAy49GWylD5berqfyajeMAAO
gc1zod47gw+MRjVUR8N7MddNzQwaewpSSIr0JjLKmGuYMNvWfPDyajgLrg95m7nO11mcHWG4ITlV
sXPNUS2+D6ER6HOH/r1QnEeZNdvMcx/ii6YKMJ2ddCoH7n5oju+JgHXU45qAgEgUXeQkyGi0cK5l
0P5DjyZmEoqcxfgfhZzfpnLVbVrdkxHJZRbndRPhfl1L/n+Yi1eVpiGcOLMOACCgjtYD/xQe7PwR
HsmyJwLjrRQnbVhhPtdT1cTQs6igzQcd01Iq7AS8cQzFUoF+IQs1mRdyPeNx5XKK1KlaghwpBWSb
yv+LUcaPE+iN2X0VtQsC+QntAgnBhOhNuqebWXXubZ28E/PPGuZNPAzG1MywxDbuimPRAvHQYLjx
5lhOIaAlMIcnr6wHp2LBfzFssEyGcA9pNpBj6e0k341cqEXTUnGexyiyVk5vGOQNCsB0kBS+nerC
WbMVn7peq6g+lScZ2ZgOivDLOF1oBzB3NxlMvPDT0QFdqw+RHOUS+ggB/AQSxo2NOUzHZBDBcX9Z
GIE75qXR4dNO4lhzyTX5sDHgSeRslBPH/ErRTPH3lZI2b510BRKeVAt9/uMOCIruCNSJO3TkzohC
JFQfSd6GgD1J8rG6epzNNZ89tUuc1ulfOSV96z9mhebxqR0vPdk/3ZmbGt0tPIC2zJfrRDmoulMM
svPmpnWW3YxAj/tzVqhslFAuJ5P+N6SkEkyFBJ8SPpTowgul05BrOwxOV3X6PoRPzP0/XP+Uq+S8
jsEgZnjfbYRsmzNGbEwqSiDEB5kbL687oNS59ipdgWRi/zjkWuibY+Nw29uENefNdkx+HQY/Y3+A
7knZe5ehqUSS9kExFcMAzapw2Dcl8vCaO0s70ntfLEbvbc9BbRBlU/xgR3uampmWXHbhCw0Jk1Wh
if4XDNo87eTevQjA05Wb9dxCVMTSt0Ur9ADkypH0/mLQO7U0H6+NdtB3bwk6w6/adPBuOrPQ0ttc
mIUC/Rfv4OxWA3bHtnBLF7yYI66d0uaSmRCJrfMewrlO3O3AFPTsdKy3T6lzNay0a1VAL7+HzxLc
kyQoOmQW7LumSkyjdm14V+iQWl2fsIjMGPI4SFVeXYXC7a8yA27JLyXNJZGZkLfoV3HzZGYpxBBP
DNWN/jrOgZjv54aQ1JqgK/q2VwK5Quas8Yp/OmkbLLCZ1KjBqmo3gyS6piUAX0YbCZMw50AFe/w+
II3F5vyaVKDMHpBs8OhDgio8K8Bd6r124xjog55FTaam22r8pNAtE3aetFuoewZjOyQMoI2zO2UH
0hThqGL75vgno815Rer/SeTjib3RLZwlePpJ4a/MNVHpCIXrn2+YjLTSQjvQAvccJ5GtJ4Ijunex
J0NRCQbcxJ+0bnVDNFAvjAwAya+33z5q3dkiIZDRDlVm5a0NM3LwpuG5W8pMViOZ50kYJ1Ne908x
39aJcb2d9pFIBvyaohc2i2ENKpWPJb2qzjoyXNBM+Wlfqa9L+4cEEtnWndyueEt1ErAbUJfAEqDW
C6do0V5DlXCVuSoL5aUF+LrdslV+5in7JSHIb+sJjbBczgYYgqju6er8BQr+NoTe1okos1BG782U
fnGj5Jsl+N1cc6SD8AONOJzJoWTxx2YUApZNM8KSI79fJIsUQTwOtv1CVjAIhFvTtn1sy+3YdoKw
9XgzYoBVEGTeKKerQxyAeuXvltiyxvnqenQgzteALYxJnNEMoLjSup/OVHLnXWpzx4w85w1duw7H
oay9cejif2QOoBAjCcnVysLZiQoTrQl5wQF/UJXOraY2lBDshxQN0EhyIEyiGNfRFSiEv8exBdeD
tFO4lKA5inpeutA2VL1YUoCCyC1KJlzKctgOWP6RhLXJqxxXWu0QO1hwv1Nnwh/p1a2Nr9phAN76
AMPyxQWyw89EIpOVRh8yp87JoW8Of6AJGh7+kg/LlXSUT7YZrV6O4UPzEOxihvUTtpytlX4O39Kq
xvV9ciBJj1nAYzCrlM9UX2jbKMdxoRTmpLMRPktnNBnmTUzuhEEYuBbz9cdjb2Syz+SMSFaVHhtx
5Lf162F4RauNJKnRSAbkujF0xo1cS4VwxJr7ua4vgCYqSBUINvFWyu3M+Pk9Krg8GlwFcHyqPQA9
24Df4H4rdUGiYRdc83CuKGzqNOpc7Gyf4OWcg1qHk3ky/JRzRrOi4ZD/bSgUxmlfcogMhgb98ckg
cXXD/uxbjc4jr+LyEk17gNwMW2oyYstjiiHcXq7QjAx6BbZfFKRFmlTcv/zPhFZLsO2EZnQg6rGT
eAUUBu/ZBDzwWUF8FabuZjeNKYWZklZHVwUGSgCzxwIn9MmWHT2nmNsG5hxAkRk3467faKKms9It
+gSHVDngnzLo5HFGrSHjrxE/Z72n7sORRKI2Hmwx2muhLz1q7XN1gZoNVQdUf+yfu6HJnn98MiPf
prJAj7/B/y9wdE4PzeCTtZd/ZW5kedHCS9b/J7Ntr3I/CpjkNeFs2z3Ib+aZqPRRVNl9SUKMCxXT
qf+t8b3auQ9oJQMBInSn3E6iGTKXox8/Ty3+egvQ1otDSu7HNnS/aRex0GM23R2iF0V1W8Z8Lgfk
CfrIHJv5qshIg7eMHGYYLbp7zXnT2USdFvBoiumiB1jwIkd8nMbsUyWjK0vOIYz7Q/Si7DltgfhQ
IwA4hnbt53R4cwP+c/6w21V2vCjGrER5uWmdkkY40/keEJKBuPI4vmP9DOos0RBjyvCXO9ccKB+3
/I/zuRW8xSZqDPHwdscQNaPgao2Azcde3DV03TvY5TuIRB4sJeXzFVUoXweD9COFan7rglB56c3d
lNMUmzKrGWnMtGOh7vqcM+qBNqjgz2J098Co3Hm+ryGMhPgAkF75nrsqcj4eD7F+lxHb6Kurc8xl
tA/4chHJCovjSJf4RjZM9FNjLqhfcj8k6lBI6x8C0tRk9QzuVBkccMW10BhFlrAOdBK+qoiClPDE
/B+rqjLWpTGQ1JqrLBlTgisCj1te61yO0TgJdetyK8fW94R9sk5dc9nMVlLyDGvP3QBUTQT9kFvy
wAqnlTeXOQrehs6z4GJA3atse2dL0W5EkwhuaErBSYQHCIVzOFJfjunLaElCmc2V3lVw1uGfhicO
XxCpLdSa2+zfyQYP5JYPHy/Mp/ipFsL9hazXzAhnhTsWudfkJipPQjw5k7SJWuHRCVvEdaIcU8Ej
ukFZlMnXowdBwmEfMoTcceVO+XR3fvknB4fHFG8J0znoJMY2lNslfduJ50/tqkNdIwZHECxRYvz+
To5T8QDe98+jwoMpY/f2k7BGbKiWhrPlhkLN/00opP/uwGLmONU2NcLQEHkgXN+LanEyJYV8g2Ct
OVwmoz+z2Bp+r+X3q5eOcMqsk3jg0/m+vFF9y7O3WMNwpiE5N6DrbkWvE7jzeWY7Lhr/BruR8bcR
LfEMjRke2fSBtMOTxriBsqUXQqyZezbcGR289LGnEFfGmdBd2HcMaA7i51fXOquUioE1qKRNNNXO
KVciJqtvpX2Dk2tEK0TrY5IJVBG+xwH+76H95UbdoMjSFkOxZ/Px5L0ENFP7v7i815HENLrIPYH+
UYlhOlQhb02x3P5VOu4n+TD1SpCwgJc4n8JTzicrptekwki4Zhun2atmLbvR66aayI0OZOa4u9/t
eOpQtWNcRvBefNbxtwRTAXXtPJu/mmqoZc8InW76QTspjoueygSoNfR/2/7ZpFcgV7C2KIlOvL1x
7mnR3/Fr5Aael9xFX59knHuzOeyOrpfJhuWNZ/UgdwjbpqcGJjawIcYBPCV2TrNIpIRKRWgHMy7u
mjK13iK+6/FjKXvgCRM7MzCuQ7jk8FkgnHQfALsro0AVIAEh7P+xFxQlsTNN2qUB3NjIHMvu32fU
5MAlEF/CUqJ/jSP/Q8dqcHXdAcwMMMzOGENqYRx2gEOVI9c/fU0dRSOy6W0SI+3EMteG3ndTUKcw
1gQrqnbKMpODYknloU1LkIA2qsmJoC2PuuhtTcmqX5n6YO9GBk/oCcY9vrgfCIPR5xir1EZ7FdZ7
q20NIQa3EMdJ02bBtpEKPH/GoqUm7Y6skBmUZOMTHjzr0mT8KfRBZVgaawjq5zQeJmrtnuV4NNPb
7zUGW1GYB3I4Ce1D8XnYeVP8EHP/6d2mlQ2BBK5r9xXzXxPRwH4DnFpC1GSabPXRIfCUC1Dn/DlV
jou0g2Ln6Pms8r+KqmgOvJHL4y18vrDjvFTX0MwmZkN2+l4Xq5osXwFHV8i+mEcY6CA1Plz9drhr
LABCnGe+8AIdjYA64FOZc7WNy8Yeqk5s6leSjlWi10BcbmbqZdSh6PaYqoz2JZDg2IpYCyurSY5o
DBWjElCeVaBnCeaPgW3ApmT9N/0pBXBdlIuoqzs5bvdTeecfHhMS6vqPNnRxbCwqb9I0DZr3SVp7
drsbpX4BcehKubhgrqjezwFODICOBJZtXJ5ok3zKRCvaM1i0ovcoAfpwPWQwlWihzJlB+ytzNo9R
hNdFmQwp8Mmv2cuA0CPWvKI0qKBYI4yCoPUFCYl+BgGvs1fUBYZNDwc59S09F/SsQFvY161FdQ+7
E+zRjdhlRTGLwgK3vI8+x2LOQqUfXil7CB6UStRv6vvk1mk+MSc4xP/0pyPMBeZW+YpxBeHfTANQ
6C85SXR3RGVnBtbX4ngpj2x1fSPDVR5tI2E/9QGoIRISWBlrVN7NLOw9UnOJHwVgMn40e7eb641h
1B6B/5rQjRlH98TpxIAoDkV/zsooxDmZnLVpPEOJCS/iuDV2OaI0krdCN7PGdc26e0JZpo34z+5O
Fivku7VigFBU0TktASUL6lo3egQLx1IoaSv8e98rsE8yI3k4pXxo5Vaf6znMbsBZo7lUPSRZNTxk
8wLS/4YsX3CDau1QJfuuokNS6vT3MFJiUyxrWKesRx9PPjDKM0+u49rOeBxIfqZwq/eN0kN8RwkE
DkDqC+yvw9n3LaFvDD7qLKNTSwJiW3BeuA5yq6yXW/Dd8RgMZ3t4flL8/3YnAEhTgalgp6vM8Qk6
NXfKqc5Pn9/OzYQDn5fSWnzNGQ5bKyasNwfsjaX1nhASZUOkyz0JPcXaU/coJuon4/BRA/WWVDmD
bWtpIbwVqhWPg8FtFQeCGx+7AkPy43wGgQDMtfDRHxgOXqXhJ5rIBPPy5tYJnRVxR9LGN+JkrD5s
1HaXLY7O18BJiVftkZ3MwdaselOLxd3eGgBURRiS7g3KNYxnjgFPNJAchZxEoQQOJMOf4f5BVAwx
SakOazVH4P/bfJDHJsFpknNwR7BdxQp4TL+SikKL9JbNrDtrZd/EhWAy9SRapVnK0o34R4K1084J
S/fc27FZkxSXUNITZl/3kG6xK79hx7gsmd2QdWGgAWniZQNkV+hG44foE3gseadoUPBtqaFQBNqH
fZnn2z73NYiq8MSq4V3YW0IMH9Y9yO8G81rm0wPBR+7lnhRk7NM3ZMGW1WRW/ph+a0S9nT0EYd/I
JL6W5omxwj6aeN5lssZUp0tM1I3R0ujzbig+NG1hTCQ/i2f8MSOX+CDCCt4iPD1lp2OlAEiJfp/M
UHyYW3e74+vcbZyewYrzctXBq6o8JHqPzJUxZZkoNBrJDhHlHjDgprIHZV+Igs/yRMjD0MupTndr
NMBBQlqeri8IRRrPTPxL8w69M/qKSl8Qlho0pemKdSjbQG9DoU5Vgz2GzB8z90UJE9E/lX96E/gu
gKWR8bL7gewfquNIhNXQxOBrIYr7c+hox4VvhGxpNPTUxa4l2Qk4oTuBM9vOPN7w2mG5r5c/RruW
748SdAsI4qbthI+UM7ZXKjq6+7718uHTxn2+xAZHBO9AaCo0QowQmWnbS8pLVx/XjA04A/cHDB6D
15n8xF6PYhnNqy75/Tl3R8SzJtYipHB+VptDj+Q459FnoQWDuFVs9ivBfO+EvCF74Gz6SPOJuF2S
IVhOy47uM2p4khOJGgeXP1/WCzolK1QwB7TtvAfWckQSfMn5cHUDtfi27tTMmxx3JMGhmJ8m9Fmx
3j20eL3CrNKCKRxCuHG6tINvDocEh1WV+F3Xb0PTfA8hK9y5yUiLXYHtMHbqBK8hLGBBj8/vRWNR
lncse2AxBaoew/p4WNVa2EqzCYNgThVB4qW+Ojihb2I8pMcOb0cBq7Y9fOcdpQxTb1YDhfCl3QPv
MN6B4h4gWlI3PAU4ogmoDu3Ab+mgSZ/NvSc/7H5880gwzyltvVVBAukKp6PGpuft7sKsqtgClYRD
/msZCge4wOMav0bnsWOkhMNjRzuTiHEJgHI6hP99YLw2HWDSJbdOs2eGpwh9YpdXFDUyleQrA2Dv
Vp+y7Wwr4gycGrVZqehkqEL9oXukkY6NOxeiBjnFu1XvRx78S2rhcwseIAFrFg/cGaxPdMLh3RSk
HBUO4pGGOBPSxhFX3hVw5dR/Mp5ram5rrgrbkT7tyBjMGdYH3RG/UYVXLx8j4JA/E5cK2Mp5P/Nm
990JqpiZ65voSeQ5tijCJTWrP+Ki273CgwQpVs+6NTqEwsuLIYLk36AIS3itUpJ/DFbvZLbvdOWB
+5eEQ2aLKmUyNK/RBmx50mNLoQ1DRf/PBVG4TpDyZROLJ4ZhJDpwK7Ty8ey+0C0syt0oje1NuWHV
Jhgs5kp5sKlPXYBAihJTw5WB2JjiulkwGkkCWr9vHmHiLBm2cTdcCqr1cUqyi/RrX5P0eoA2id51
hVH3eBhiztNnwnnnZAFoYU6WAaNkFgqUZgAcLof2104uSVvgtslL9bpHuK4cztTM4r3MymDgT2j0
8+1aKYaZD8XUIKaLPLn7gg0kLONaXoiqSv9FK27atbqlDs2E4jonGo2bN5PVOfIl31K2/tVs0fPT
uf4zOXqJ6J5O6bO70pc8vI+N/IfpSlfyG+X2P6BwTGMM+31OUJ4Y+a6nyEE+tMviZJjWQzreAsZh
THxE0m0t6j2m5ubUV2vchi8VSQFPSVD2UgEM3zvVEGECq2+NakB3+x8qyADoU8SVKRqYBSl+j8mb
+Shsgx1hn5rSdCxA2r3gJLxBVWNeF6MhG5XVlnHv0cQigr3pBIsN3kMSDsZItNxCuRpOydwy74Vx
1e+IvCswUSFXIZ6PtC78A/vW4lPlE1fmyD1NlyOynELp8KuHq0519HqncfeNBgxDcDSbvp8gNbHl
ql9dIWSr1xHQX40E2t7mQJMFHdOKleM78W6ZmEDdU4o5pd7K8ePC+EWbNAi5U31O9nxBZC3NUD9N
mtAJsMaCOKutRh4pvhjy6P1wnJ61lmi0UuDqn+hrTPlm+5E4/35h5N3cJtKUcnAzXzfOFlt/s3mt
KIo0z7RblebOv4OtoUJMkQ70Zm/tTyT+JaE2bknTrQrF/+t3bwKZM0HuzjBeioab6kalSDAQnE2x
D/4CzHL9NiklBe3PSzx8OyU177ycDKvnAgONXMkY1P0Nj4ByJ/ojwTwp7VK//rk4UJTz8U4vvSDJ
cBiOjCEyhCXAfX7YYN2OoCjM6dW3IsHc9deWKZqxVecZUtDRsrIrZtInvPb4w4zjTAx9ZVRq0Sy+
IZr10mmyoh7hKFjRPh/HGL23xl85sVbzV7TNWcp27c2vbp0LPJh2K6JYIWAuPInkY0yGT2iuU22G
lbNI47KRqY2q1IZJzToZR23kkzs780PgdmTHhQe++Qz5AVOVMpNkcNbBe4Ub6gibxTdigIbH1lWc
W/PObAHCIQCsK9xl9zpFhhXI14O9+r9R7bxptjaKHICGmoourt6KLNwZH6EnoSGW+fo6nGoIxzxM
VfVB50DWxHqSzuyZngYB//SzEVvAXdYMpnVR3OCPc2k/JLzEKfubnv5MPx0ddzXW+kvOBIyjo27o
3kRwK2B+RzkKdX7euw2503Q4RM8ALJ4srWBZ6AI6T4gyCQ4JLPJZliBtumeRzwNpaLLoPGMzcV64
Pni8Ajmq7/kWnS7SpTZ2AFy7abIXzcH/O41kSZ2yM4oxDt2K5vC6iv42TJJ4oo8jx1iFEqn8axsf
UNWPJes+e0FNJ9ODnbBAyh190Oa4o0xwW705BgEldgAjezi3K+V5Rn2zb1XeIFiGJsvj1blYMuWC
ywa+Z5v4aXkRCus15C7L9mP/9n6OPRmJ0ZrqUDRdJGMLC0PidUrySxGFHEbpImueL+cpdD8DnCnv
FSTiwZrajylZb2Ml1kdRp0Jg+B6QWudMXC8XMed/1u1w2E0IHKQeIX4CvSbXNCXLS5hDUvM4RIaW
oSSkYJ+qQqKoFE7jG1KEf61Uds+PZiJTFSsdGAHJnUMmpbpDai9w6Ax2QGUv5PPSQ4vWTXbjGgPG
zjea8ktNSQ2vrH2JGf0D3ssyp6524ptIAGHXrF4ZlADGR7tFlqgA1SCNn5pQ5BV/mI+af1l4W42J
PaDRzt+Qe1tcKH8ZpXQRpVSvkvOyZF1IVk6najwMIEz7pxUk9tYFnl9jNIOSkb03q1un6bsZqmyp
1sysQpPT1O0tk1uRhmAzoJCDu/uu3KVADSkdZ6xBk0+nZR16U760aQxC082AQnak8c13o8twl5aL
3yhWvElBUE1SmT4ri/nJIgWBG8hdTF2Hf6BDt1CSQ0/YcOJixjm1sc3TNr4QQZoWLQEBH6ZoxQs0
VwZCLM5EiP4lnCqKfgunf34xvhdLVHQYjJLyfOF2Y4KGNdHAK+L7DdccCSUek7hrsz4MaufJIwXG
s66O5mCwiMuQb5KOOw376RsRQItjGTamcuyv+ew4ltup2HCPEEtgpeUw73NbEu4kPwcm4qCvNgVO
z1A71j38fBY1m1JMXP19r7tPs7Kp7bTK1RAYc2mL2Izg7EFFO2CSfpfAhpWt7modtaCIYkr5+KZt
Cr1eqjQk+mupozT9jt80MujByOMIvHPVv2odfuoXjFyV9fDpm+82BcvP8WzDQ032FYwe4kZNfVT/
fen7sPXrYgev6oHko5Wfgnuc1C6m6s0Sh+eXU40g0nX28eHOuMEN8TftGUTLIT/lhwb810XWljBa
M+07XEAxecxkrJKNf52tBdx8eoMhIF+dBz1O3fz4d0r5D/qKzwRnpC3n6LuVvuOf+cczS86h3aYb
YWGpmBBe4NPMrsZ3roK8W794pDQU4Ng4vihMKbG6DVxAEYimJhjXsXwdy3KMWWlWMpO7qss9ZEu9
sXtnSYqeaLYS/sn21TUCRZq+CB/k3cXV5KYgfgWc3crxYqPOnsoGmCVGPGe96zEdZU0VQvNo+9fc
/YyczROxZ+DfX58ajCAFYCxxkeSM6hh1JUvUXkVzs6gfPc8yBp1ESMm2jjMzFEfWGPZSe+UczMoh
w6dOR4o6M1IZ27KTdIiyo1d+qeKV9pVi2mSYZQn0Qac2J9c7IdSmPFDXOhwhvbv1e6UEAjth5ZsP
WEO1ojS64k8x4Ht5riiCDPAR8jYbiR0gUPEqWpW22TGlpOtFl3rUmcMfSqVRrNXdcBNlMV+1Xl23
gsdbKD28UjC3SxexFt3qVSwUcuV0BgBuhz+44NZL/+APO2DjckZiEwUebY9TA3Y7PlT5rSXrhlrS
MTA0G8xjuLLEbkh3LkLMLnA04smWCGerz1jZRly/+ZfssF8OJ/zfbKq2y0ZvoLVSOEJwmQIxjVah
Rf+G7qmQcnYit01QbMIBv9sDUK5aYeBFDQqImu/DeoCqLuFN4L0ErfCtM67kakCWU4bQHHPeY8/W
0wvzdP/zCiBi/Y+zak/fJIdldHxJffCu+AeJEr3TjuHXiEBQh6sWklR2FoDrri2OpjMk4NxgU8i1
VZfvQlwNfUl+BxNzeZ5b7zj28AHnT1kilO54Cg8xCqTsw4RNkAna7UmGzqduNefyxTAuVHkv0bjM
a5Y2QgMBN2knUJdfyleJ1KQOcS/mfmdixR0BvQ6EfOBvaGix9DU628kYtNm4SUAGfSvEKPawWQA4
361H2muT6fUBEJJfB2a/sNRvmUGg9NbDIQ7JpRR1gHgfrzkMgvz85XCiZNmyyMhltzjM/eYwWHgI
mqtlQ1p7EAdlajbp+mS8QPI0t+XISy9zn0UieocWTU2Tkj0sncMfgLBWeIg1eRspz/xcOUmKAVSV
7fI4NUlSoFI1qiqbCEa6qEyW0nwzIWEvFNPtIXw3+sjjU54ESdDKtvKNdCdxKVioecHmc+iE/KFG
4S0gY4eoX4y95uobpj/644lcGlD9rUDXoGwrS6iErXeuM6qcrKvQUR7wxnfi/ygg0w40JUsz6DHt
VKGaLMhcjADKd5xatVcO7951+jvA8kof0JDseMwVrJ22YtU8NF/XsUjs5f5N2SY4zNKH2OXbRfQ6
rhmpY5k5a6PLpsyN8SWW21lDb/4zWPeb97j83GZGget460QPMVsquPBvA7mTaK8KZg9+hoUMEagw
cwat0/M6evqhqcJng+LdnacNOeW9mQZW8FTnN75J8p6Sb39xamV41EV24XEAwoWuLpwJAixv7aqt
hn2TRqxC05+bCtZlcVMeG5o0FLrtACW8K/TtX9fmdUG41KOjIWNY8tO5EGqTew0lmukbRBk8I8pD
Q9+aBE8dutOaHtLZ3iD3CIeT8IyWDobzbacHxpQqrj91XaXVdaWjw8yfH69WSHunoc2ZYp8n16Qp
i0Ilg/Qox5lhCccGkgRtrBFWTbYe6KeuVWRfm+Dk/SGhkH9tPmYv2scO/mH/yZTJlyRO6zYHY+uR
CC/vJR+OaZwuR+NZ22OgB+AYUMRTfHiOYvRUc4N3e3bC6NhYuhYn9OtMgu5k9mMW4S7dcdKob3sD
I3pdi9oq6s2KZACrtrygyeqowuCVWaITSa5feZ+M7NaLHU2PUPR1dR124gmY+C/tn3ckqvmUryQ8
Q1s8bTCZ+Um4Lh91WKKEkXEvx8uqdYWNwXTmlx9EUJNWtyFXTTcXXbCB6/k4RvGRSPkEuHHnRS0Z
uo7cXVspa285wuPJOF/JavphwgtISPXBS1D54ia9vA0wH97MGV821+dwrtmKPlUsccnfe2QO01np
NO2BJAL173FAodEZUUCnQn7AD2tWM6GZvEg0Ji5M+O1yGQiazzYfvIB990pkABapCwBAx9+co6UC
/QOWDIpXoWNdVzltDqTc+bn4So0qSLidkng/ZL89v67OaDyM3a2Odlz+WvpoRP48TSS4R7N/YFMk
DjS2jaqBHXy31ZJRK3qai3RRA3fX9hyFtGWAB1VSWMjqrZEAqwRU4S7jAGcYUSoBuJhMV+LfiXQo
sCTffIWvcWeOqNL5PJSQe8rcybc+FeN8ChEBhOHko8ZLyQfyi3Lm/i5SCGTvwb9DHqCGn/fznE9P
GhU9/js2ktqCt25lYOTugUUrPgpVzfAhDpohCDfx871EhxJrav+YMZOp0ZIQZ+iE2MBnqWTBGyRF
Kex5sCutRnzCwxWtfTkcg306+L+moRLXOP5ngvX9p37cD8tV5ymLPp2ffq/+xefNTtyt+nQVoYqI
j39aWO+EvrFWI+6rW7AHfO9FrHyTPHVOnW5upeFfcuuKoTncx0/4o+aqY7Kps3tWNEfpVU2r7sN3
OWzeQ3X3PDHTyWiaFxzHxyxfS9rqg1SqYbtmsAWnA94M3evu/Jo0ShZnZC5fDV+e8r0J00/JiDZG
9w57WmHZ2bIdfBMhC84pIH7+yNYWbAC7PTjKHAnf5qjcodffei10X/hJsIP2lrNipsNDmg0riJtf
IJ40nhxI1U5WFAwQpL9ZxWKTdZoGu7ZhfbfKII8x4ZZUS3+2tNMdOBiC+ArbrBt09xBmSuGvYXVp
dC9OTazcP1WA/JzsvWEixzeb2d+Cp5SNtgrQVpXf0Ju9T4m9U6/L2EjhZT8VKWn8kj70gTMQ5F/h
qdgiFLlNIKYci3ZICVq1idDHMJZrhP5p85Ne2UhhNY0nMAWT2caoRe9diEOsUWWOVvjN4grcWVe5
kGGeUZ4xQu39JkLL662d3Mv7XiA/btMTwVP2+rhjckMxCowZ9u+YmdLL5miA4F+a5w3q8Hht41Li
Gvjn6FKPESwg6WbkIQnvGHacFMoo2c08LWb9Syf4mOIvZ37zAbe/x3xsuBX03tNvGuCeCS18mkFI
xy1HzyY4b9dGPfr4yNdgQ/zNds9Zt+LNfVCO0TOQIwuTbI3YBeL3HyhBvWoGAxG4Wk6aTB1h/AIn
Gm695teFdTCXPG2rFCZNAjS8FZJxMxwYUaVUX/AZZa+76DFgVTyCMHHf5fIimnEdhiCCTSw6iWoP
sjhH80zB5OMbHciE1oc35LX3WusjP9p0NvrjE/M2djR6DZ9wfhP3LDa873MdFjw/+1COJ2NIfbD6
wS+3jhKq6cM517csGzKkXiCu9omTCLXs1eZ2EYD9QvHV8i6t+oqTa0k/QthrNh7PYvHqQ+YSMbtI
M2J0q1g9OZp9hfpcbdatzanqcWW/50fHjou4udVB29GKO8dIamCSK918AgseEwhtkVvEUfH9L77y
fXA1+FPEbbwbeSgmNAD8n8Na7hfP1yk8sb/Xy01NNJc+8IN1Kgy0Oi8LNMMZBkiZBUQc8e2LKKRd
gyAh2A0oBkPLUIaOa5TmLFwecbPZRHyFGuQYB++JTQOp7TFqg5Jyrng3ML15YyqPOnHSeJr+UhoN
Vefmh2r88OyeGdVZ8j7nzIFfswE87XeKjlamkw1bMQrvEXnBOmQmv8bNjIsxYrXTxX/5mgDtmjsR
IbBHbj8D15YOcuzUbZnuUJzrr2ePuxKMZwNxq+WhZ4ALe6/QnWg3cRGI541CaPU9LF6MfWm+juwd
U2NEjiNIUesr0YVvuhFjH1XSX48CMXZU4r8xeQX66cg4XOSsvtcqhCy8h8mTM0KcVKBJPDEccvUs
y70fdQmmFbGSmLcH/TgvOqTCCDv+dklEEwKDKd4ePgDkLws/8lFS87cLbkQjOmQ2MsgL1guuAmLP
vEOVQoWpWOlG4AWRlczg4wuhsl+zwynRNqLRHxPpkaJ7VmYnyeo7B1aqGtJB3FNjwny6PScl85Hv
sea/Sat+9DqObBFCWudNZS5IlXA9QhvoRv2s9fd4JqgKUDEu8ALc7ptfPWFjFxApRkJPZNFCRVo0
QQFQ9ImZtNQuLAhEpcMWPlTfYrlpEf11qEfA1TSefe7BJY0aipaFel0uts97wSIXUEB6fiz0pz1w
SpYaHn1IZLm15GsDEsra9HhBGPlN7fgZ8FFSbXc3iASglwp+uQwLF7OR8ChJQyIVzDlS2awGizMJ
ZZDJljXmZX1BOFhyDC1oday/+CXfB0apY1Gjca1OMYaWB28VJjFh74ir5RMG2h35AFDpJ1mggifX
MgAv0mPgmrSBr3m7XfvJUsi5H55n6uw0fCxCGqQC6PYyGKsmf3ABGfz88ivGuP9me8OtA14+eQ1o
3HxXdyt0UVt3N8+8DeWNxI99DGH3MReLGsoMZ+9NcdOPhPx35pFmijqwUMgTRT2GElJYiogljKFv
YD7jD8YK/KgwovCOR1X4VPHXBCnjyQ/33twKOmAEqKjuYzZ6SoAnhEnC2FNyAN5qtZkSiegf2AsV
3nxNO4G3i3EbXhpOyzOaU23JEGKa358n+59V9JOmgyjs98lwRdEzoYx/m41gNL8hfyReCyUFP5yx
p9SMTtGRxQTjV+XfX3VTyeKfJs5Evo/60vLEBeExvLsvpm/0xh+fp7vRdG1J4EFY4eiTrEkua9ON
5RhY2h+Z//gKTlinwhic050jt2oFJoJsoCJtRTsUOr+AJTj1/pL2ncgUhSQNOpLYQxHl7S3kKinz
O5gWQXh/3w3s2MN2Su8uqBJ4uK4AV7DS09LKmHgvMUvKREW2JHoGQJUgXRSDRP1pzTLO04/h17pN
1wRLo0OQRhotHzZWJFXh8mWDcf5SZkvG6OQlu0I9ti9iATWRn6KG9OH/KLZDVgq05feeQ4xHkvTg
mI88vMltBBPSICMK0GBc/m+tFctkNPWZhRB/Oz29kBB/e0Cj+tzwpE6vBVFFctOqf9vgINHN753E
RSET4KE47hPN+zvCsbXRjqGJjmmqkVg3gT5jQAQDggyXVEkWLf3iWFtlzfAZa+oYtBAenD4EQhHr
GUchbFKCtMZLou06tD2xrGOCIfN/t9stEhsgYf8pMj6oO5iwGMc0Pm4NCzyR3d+Dbq919alFdvhc
Si9LyKPL0RkzrEDHriN3sKtFWzoSAZ54+LKfQA58twax7c9yc6R30OO+x5JXtnweW1V/vgSt+WWK
b2aJm4SUP4H20EAxYzPBPCL5R+s3BuLlLfI8ObsXUSez7lxspXNGRWL4HG5WMljp9XjuBxz4n4c+
is6N02cugcCiuausHzpSOHW5BQFVpKRhPwsN4r4PnrP3M2RhRsLulxT9MQwRsZkXazvSgcCgsYOU
fKmFWm6SbsGmgKMa7nqZt2MDKesHvRq0uj4vukRDLjgSCdaqlFlJ0HdwrIX4r/7JZH7RV5taegqm
MSAYkbC0idczT5fS80lPYobtobR40P0NEn5Scc6PBKCESU6b7JNQoDuRT184d7y7mJrWEov0R9Us
VUvnK2O1FA+qOCSvsDlZn9Dv+1xrQfnRxrUV8a9cWSFMSJLrS9+aGWNzOPBgRdVwycgq0t7eNcrG
UgaeN2q31SKNrlbDVRabcrAkEAFL+7ioIVrogtJLoJpNPha53oZz5+QoNvQq/qqp/TXi36RR03XB
Nyac6GT8xwI7qZ7xc8W9JDimK85x1L5QCnnhGqCsHbDXMR1FHnWk0LxrT2hFBnvISw9aKCkPKVS9
4j1IRXSi0yE35afz1yNLjHJ3uhIUj/la2VwOTzR2rzcJuG/KxNniP51UduRsdeJg+jyu/KQZgVnw
rxk/zXZct8ES7rWVUiq5VWSLJgfqjWqdaJGxGWrMmjuO9HWDltB48k72GCurBvErz3eZbnahhsVW
uzHIOcB3Sps+WbIJaa3rD44G8WX7/gw2OyJBmBx4NOZLdjHzKOIMaN6EYZxuQx+P7AJQXa3exb02
Ftn150M1REevJ2X0Cjk9jLvV+D7mscRC+NbJBuHcZ1lsIN5K6aQhtcpJmrS8sK8/s6raR7OdRBWd
tu6RtlEe49iUEMA0QlaeVlRGmN71FCxCYsMc0FJ48poKW1slCOuzjh/D2EC86KnpHkhlyvimhSu6
xT6IseGvH7JEwX6cPMwA8KZcxjWumPYeDUSQsAPaQpzG+V328Y/r1RyUofpzewt6n8mABO8asDQW
zVmJsIoHSReIUckHdKjCURJdcuQEot+DsaE7RBrIXFsq4wAUZcIhm98oF9LPY40Vw3Xzc0JNpu2Y
TORC9KR27hfyIDM5s4b5yzhs7c3ZOy66djmK4Pn01tDzJRQ6Ou6nVCxPgyIPYRrsxdDEdWSf+8pX
mtYG2FVXHAvEqrqaQxJtCYOlSSYWEi3gS18aYDNaIKgW9XY0ESYf8j9M+OmBRcwlDt1LCnFoIyFi
aK3Jk3Fv5BEVOxILsei4jFpekMELHquI6brLyj67oMsOXcmqEc3a/qHTYc1opGHKjcNSnLaT1mbK
qym59y/eUOalpTK0P5zOk8ce8A+Bq6KZtvYS/QWHPbxCZsat1iqLiOFWPub7jI8lE8YOmsc8PYk8
kFge3CLgIKdHwrvRWF712BeCeaZItDLwgMeRUZvyJ3UOfnZ7cgO+9vN4MIeTWRdR399Ff6TbbOQH
0zdn1xCsRWSDug8IsF2dmYkB9V013XW82llJzVuL2NxrpqUKH21Fcg4x7JReLkLc3BIRgQDktdC3
RqFKx00UOiGZKa3lXeAgc5QdjouhcwIKWZ1qMGtQ1Dfz0BpHW5wf1CGuqxEs+wvVo5TbRLgxUrnP
9zPcBHI5Ep4AvCOgfDW6VUb1VKhChtXgYFd2312jvM15hVmBedOfm8qZGdOqoDD6PrB47VpiXRZj
lVTa4P81niK+NAHE+jbWQM4ZiZ+IupSkMDfnbMtFxFTrV/EPSwk21160ZA/8cv9YMtPkW6F1flZg
XxwYtEUB9hZgKLeJMGuORyHjg6z+m7Ov4TgO2HMLiPtQjzeq344XjQU42NkPqVKR7JYS2RRJuIWq
OArJS9z6TSpI8equTA5M7p1qkajPduMNJI7HXbKzDHhDAB0fiwPM877JHabb5lXAcCMKzdtFQWbk
2h5Mtw9Ut0gpu2iYVcg8ql3l5PXNommSnmffY02xHxxqBz0JcTbT1USKcWI2hdFtNitjbVALD21Q
Rrh4Kc1RYu4U/TgKcEM3f1Sb/AnbTK5+bXOE8UjCpUikegjPOO6oBQMg5v0mO3ea/95T9ejbUfZE
oUskPpVqAnJvKBC7X+EdRHv8YFZhopovUeUTJB6A1j3MyEKLT+f6dvo23uxJL6hiJ3A5ZpUJ0AVE
OSGqU74gAJYkm7IYZJEn46kzSxsveac4TEWLEABelfIzjw8bmLT+a/ntJEry3I3Ua6aNRfGEXnRd
U6VUfUi8UB1PRkvUVGWANmXhPBNtafHgetTuYDbOftD+QKV1aAbsGg/LT7MCWXhFpvdXo/eP1bN1
mMia/LjELncSkswp2B9sEoADTOLo+dWLNMrGgbxnfwrI7DhF+rTxGpgwYxMVRnJzQHQwr8i3GAcp
T09aFX/xyePBGeRXyT8YDYY7v22hlj/DiiAIH8pLnmItvtZFAtqXweooggXGxN8rxdleOyCMKY8i
2Fjr3AM9rKL1rUjzIUezfbDtO6ZPpW3u3XFtD4ve7ClNHotPhWvqN1nJyhDkhfnJ8LWdzzlgw8ma
1Vc16WSu0hwQUWNEG+WbNpyWi1rUsfqL3f37NjLwTF12pnVX/wIX8Nj5rSAQEvXkf2cYc2CYLpuu
LGriq+wqCF+JHPhIlqBNch11sq10BUoyJqAZBBw04CnaAp+YmawlrcfLZ9s/rwC5J3BJW8UkceYF
RtXtJkHawO0MzAQdi6o0D/ogEC1eKEO32jQSNK7D/MHXQKehT+QkIQjbEedj6s6p0Th5zaHS88XF
zds0WvWTP8xhk8n4YR3eo3MWpkjBpRBNabu1W4a9tH1qWn4AP3xX8CjZqWcgo6PvqB+uGh42gQLM
Gg8xTFoTTZneL5ji7NCa4Vtq4N2gldSr4di4/TsMOk5ppvf/nbYwmKdwTHYMLvQOzaphAN6TLcA4
K2UhC+KW3uH2DSlFP7cbm+ShCfxvkINWLYtvRynrNObjDDp43+iW/bIgv8iF4PZWuJpu8XrnSR6+
+pxCRUlTwVlvVG3e0pNF7ZH37+yhI+wiOFgj1zda9bjFrmkW9aaNJROAtuArFQLjS+gEsOuyA1in
woE0xmHTy+CB6HrDPWVkiGZKLRaTK5f+hfIlOnC9yL1ZAnTtRAG1A8TQWRtZx4+8WuMDZ3PBRraS
Jmdk3A4ZPpNXfh1C3RhxX6HSkpk5y60FLiG2KpfNl6QB3dlCZpMFYmtMpF+k/EdkjCmoIL7JUwDg
X4gEjxITvJdK5Tu7gKW1IEFdW5zYc8pN2w5f1oHnu1kS3sAgCONVUtSa3Rn5HllLtypfIQyGemNK
RXJ8VQzNuKqgD8bGtsEY0BYzDN+ZA6zP5/9+8eJ43qlPzlculmae9heYCrHbnMM+xPJ/YIZKuU/i
4pKbhSNbs/APvu+i2SyxjLAJ6yOzLF8QrGsi7nGM5uBms6RJiS+eCWcp5/Z+jzkkaQMYwJqrS2B7
lR6gKPzA/sNh40elYtt/AkLyEN5nte0dM+6iibS2vW5DelTKDYndhLaN/Knkq1GmGNYfS09kKMzC
Dc9oGwCi8vajdhnOD2A4/RJXpxkbBXbcpWKw6e9/yfZ151a4mJQlTe44aE1StEhJQeIb5GIJxVUe
i7TZE8Uh/7yt73vE4+GPmaVpg7Tekh/RYYRfxP0WsbxH9He7F7anV4HxUWIG3APS6Z/RbAXHgTKH
Nz9lzeCg67uRwwNXqQQOEsHuPgpEogrrlCU03wwzpPbTlraatWuHq3bHFx+DZNJY01kqCj2GLuwp
P7w4HYdh9i6B/yVzToLmc3ZeD6FbfkBatLKa6N8Nf23uMxma2nYQZO5NJ3wN+wUyWySiNqW+0Ixx
VU6wPYDdxIW/P8HwMk+MTShMl1Gg7O4FDSOWFBTnV6r78K33PN06pjPXno4BrqrBIS8IIxa5t1Sf
hMi9kZbaXt0g8LQLn8wOR44WHLnE+gGPvP9TwwY7Hoh1XFZFbkuBXD9zD2q5RzXuOvZKZZUcBtNl
r+O4ebAxM1KOE8t7Ov4QNxdUqeBsMgwD5KNNtJF0T8W9R7kbo363x45A2WsXSYayknAOjQcOCs1d
OpHVbJzhDg2ZiHX9M1vXB4ApAe2XKsF1sXEKijpvOVtncerTMToOdjlG4FO1cdxBJWteYelqhDwQ
SX8iXHC4AhFAFLwzCzJw246hAFuPfmDw/oHLMOa9rVIcToUo3dGbN4bLPiR2aPBIbWlq2eFDdWc1
CkJAuQH9PV4atJnJmhiPI20GdwcLXyosI2zhTpZ5PmkFgeLGnQwHBBuzpZxupazvqmlI0mtYJKSi
kfm9tIUmHyvDaP5jcZ1zPkwn1Zx0i8aJ/ICKKMS+yNViwKMBXlnLVzvEB/L5GzhD7V9UHJ756X64
Lu+3OIhcdSStk6yA7jUNnpPKnffC6vf5aAI9uu8cOOnl7AqORdmL49Yirw4sPrOsvoGHvB4fTCv1
HH6JkyFMvjlZag2RoYWLThalXKr6TaLxTlH6HLPhR4w7fueX0+Wo13ESfX8U71iEvoCr2qwOtCkG
XUvC+MuzNp9xkES/zGgEeqJ+9RXqnZVEt/oDFgYmiTE9cLB2Ad6UHdsIH9jNomHGFFafZr0dqnTV
GN4Kbab+gkzzYwWFNaVIMO8OUevnuf+NA8PDrjPx+HUohICCoH/MS/Zb19plhEl66h8EhSBLyVUi
Ng5qxJlJwGhsNfPRW629rgMLvOfy1lAt0yNbYYaRGQ63WOW2QAGWwsHS90axU4Ulb2y7qLIt//zZ
PoqEWzeyDRXuoL8jGZGCrVv9Lc0IrNASYNMSwfmZp4F7XiE4/oJmf/hpdU/cHfSBQoqGnlV5KGJX
DNW8GEdgDtj84XB4mA5ziMS6YA9LdUK5QDfOQpKeeOYOMJPXzWqfvNM9EcWAHbE3YaTO2pybX6PU
KfEHS+fO6asjQtDRB3AQR9g5174dCv7CKAb5M6BD0zX1p6txOGNxoxEfNBycg4mVTH+c12LAhm6H
H7gE3TjSG7QllIN4GyNruYbElZNEOrHFuNALO9ddpi/xYSgKSZjLklfk9rLQEIaUq35xgcpaNBcV
NFEXi6uupETuvl6JZ0bbIZwkvHvYMFzj8mC+xJ7XdUYEFkMTNJnkhQBhfYsM84gU2WuRFfKkIRe1
jBtVISkaciYN3reOTYM6YaOzEcUtzYST1T1AoPvFHsvd6HAAUmtghK7p5zYIHCvLAGrmUGTJ8LVr
n5bQI4N1FY8S7S3kthc87crmzEXmItmcSeO3sX1k8x3ya/A5Fw+MpiJeXQ6fSIv3UL2bjDqwRC2Z
hO2R8uFxdfhNmGkQHjY5IXqiGn3+Df0L35CruhhhRdJ9k3plUFNIq3KOfWxCKYcgEs3dgHCpjd02
Z/lQ4JQ13r4dFtqUErxdjGhBsU1A6A/rSmwSTgYLrWKrqG4K9gPARhCHud0Wi2Ld1bTtUPiZcVlt
M5xsy8htFg4AILbLKAEE3szkeYCX77wqeJg0fyQTCkDZC4HyUODCBs3O9796I6hXWGb7E227oUMG
RcpUi58WNerLOxvd3VPeyRlQigCKf3ytw1UfJk6EdJuP+smsgMmC33nCMHXnxBsJaTEPtB2bRuAA
q7AkxnbAgTaNaRJAV3JUuHO80kuBneyk02RMXzQFGKSt0cad9v3UfNo+xjpqI6Sh9ExPa4ULt/nc
tT2JCe4mI7mQB/duNeSIamEHeS7oDjsVErq/Wf1GpM0NCdKNeb9hnf2b0PlrEf0GZGqNdDsmm5CT
TZ87Wn5F1JwK1zyqUxxwXkHV9K7qyqHSFAzbJSAOhQJ5e2eT3hcCq+km/nPAliIezDu4KRt3GleP
GVm8Lje2Y+oXQB9GZRuZsuCA2mZgPTck54Wk3WfGJLfxN06NEQBgBf1FQavPJkngJTF/7AxFUjmu
ogQ79gBCYxOIWen79AIvGzwDdD1PK5rqk/EeJcQeFjMsgDyIOplhKuFYl2LdGfUGxfukeTJPD/Jn
lbvgc5T3SpjUdYGtekk93Z9uBksB4qNJaKLAkRdGZx+ev5h/WBJZDbdZgFlSx5JfN9Yp2ZMb1J8R
A0v0hbrVvY/HBtE7+4uv4v47UHNm7kY9nHxWYsKvorA8ylqhEqKSIp74NYHKVtfLF4UJadmW65jU
w4z+GeL+/y3ynt0nmx4B5zZbbS/yBMm2R0WID9TXiwVkA/luO/ALDFVFK3xQu0iZhyawl0UmZm5H
MJXu+7ZawjxE7ks8C5a/qaLrndpyGYu+R8tjLJxrlP57YPtiV0KY9V5u+qSCLx0j8tozzbW+GCU8
ReWawv/NZGnGPIetmvJ0/0UAblD/8JvbOkaWuzZ+B/ILD8QlgqLsU/HbZFaNgFfTEADDnqy7qpMJ
cnA0M7HH1UvoSSDGub8fbO7bRXKZuCROjeqx+Jwir8FaTYXG7APSAkIO9nzlrod0KDCxPRGzqUst
7XY+MYkFtvxraWs5noJ11HjmUJguiXBuoHLNsk4eckLnyx2/o27kpS6t7be+Ixlu12kTmByU7Xwk
0LkYlDXjhzOMj4enQONGgT43zN87MJsQK+D7AHSYTP0QGWuAPtwJn9gfc6qsNp532KBD5fahQlFR
Wkf4JNqjXMFctJUAmG8ZmfrDDcmeXlthwKFtYA+uLmQPEdrLa2vbW9s/RAxTdB0TEOOAt/gn66cg
2aKUqYUCxKAttrkOoE1RZibYtXvRgoz4XDM7yB26ez8DbXk/wDVlvQ8LZCX6xALx2mqjoRJ0HHUR
zIb7cGzuLn8tv9JEjLppekjnldH3IX8g+NLV+7uHdnVzwmIHCbAX/6pxo4p5qwvtpnZvU2APDrwM
1oktnOLCow/JDJAeGDYAYcKdr4yyJ8U7PNpvGDKG/0mE6VofHWyuOqoDYafyAFHcuvOPLSxguAv6
7GqnFfiDCcNdg7TVH78TrtZDYOg8Eu/x0NWdZmwY7T5ObQo6MZqz9+bnioHeLI/41zmJIGqhnyR8
USNAPh/RwLOg5A86jI7haD60K4koOTRPdmFhfg6J0DfHHFk1JhOEQt7T1wuaz4czlIv6rAuHUx1+
8rXGwPo4Oe8wo3nfUBg16futYbz2n98lmcrOhj2Ysc/ePMjMu0dbJgIA9pVx54AHA/CVr17g6wu+
PLCrDpX7uxiATcsE5i6hNxfrfIEB9lAi+QvtWE/66VtRpypzjD9wLUrYDp7LjAdb5j61BB5klVPW
IX83sjH7Kg92Qr5k2ir8yk4hqAu/buvbPdY7v/6W4crFeI3HXVRp5ySfvhLlG+IB/bQofPjnipGU
xCWllq6H4H7y9efsc99b0th5nbQuHU5t6WcA0Hqg5DCPRbDanj6at1pOEeDwURg3WlKOA5wStkE1
wM3OqNHZqwI/8VQuFwQHP2LfkXP2afNJpe2CO4FD+3SYvs1gv6idA2gdiRnO/EVvHdSg+3dnTr9O
KZtxoqbIzSO97V2ikvde6YRVyv4XAX6snv/0n75q2hCmUwuv2E+gBQMT2IeAJiI9g9gFpvXOOq8t
CG4o+UILVJFvjU5DgbhQAHzdBOXQfGemT+2dyQrqNhIq7Sj4eGNadlvhbbWL0h+84ltv/71qf6NU
LEnvYHDy4vRaF8gdxvX9GB54e79ztodPJ/qZ4Mt3kysULmr002UBRsJHUYJ1zZY/6KIpmRnP5WO4
Ue81le3f1lLFZHBmY4QjpIVEepfwxj5q1ITYVabRsq6AFBfy0AK9a/x+faRUlXHE6oRed5Chmlm5
XoXEdC5z6K22Djlat0+8YvGu2JKseZdZ3RiQAGa32/KgbKu2ptVPvOBjB+hZQIUV3AArsvYWh6S4
gVMGB8UObiJDgELD+BmKgtatsDJkOkUMOuYkDVMRAbavthxZSC9TbbzzJGbcJE58KP84E4a2Anz0
NhD25t+Iu1X8tJ1qKKxcQr/57e8pKVZ5MlYPrPnXB1xrdFBy7k2z/+xvsWYF3LRPHg1J8Oo8Ruob
DlLXzXMpNg0GaXzAjMm5s3FmV/jRVgre7km8FR3/uH0XKSO28BkZC7vu5O6NPFfeOZbsG1joQ2cG
7b1jP0X0aw3p+tNqsbBncRl5GosQALDx+6DrYIA+pi7vUDbP8Nb/dIMocAhNisOMP+d1esO5UU6/
etxGSLN7oaAhEwhTVvuLPuWwiQKeoosjn3fKse6EMx6NXEr9yIu2GPU4UWLrzlamoMFpPmVrDvLd
xwxlY1yoeZNwbOSrwPFXC5uUXl0E5Cxgn7K/AxEnQhom83f6+Gvr5WcWDDETpyl76h+NRXt319Cu
mW8fSwij+6AFwiGIpUgrkax0EglNjgOaIpzcw8hYN9h5VW/78B0CrOdGKJ63HLyDTP1jW+H7WC+6
qZs4mR/X46/VVwpG8Y9QG5qQgrIMF0BCcsODDVg3eT/v/6hSJ66p4tzfj8qj2eUPQgfMWxYtWCnS
p6QBWoDcwH6aBrAwwncK5GlotmmC9JsFW6+0p0jWJnhZTjGwv5EtiF0qj2a5ATYEdvl481n1K9YB
h7fUXQ8Vlu8O6nDdrIWYGXD1BYWBxQozd9hcaddtbfd8RYz5Lgs5lYrf26OndHZwDhGUe7fuIACV
2169YH7vBpuX7pRGof+aBMksfJGaX251X8/iMkr8cRc60aycqlirpUTWqRGel271SGD9c0O69qeT
cYFOVRR2TbzkqnjNS0pyi/h5yBmMcNbm/TCXkX6UkHR+GBJzD6m9Fwiua4wVn9+HriXGicv5pc6x
JZz9XU6BIfCcWfHnZiK54+Vcmp8nMv9DhJxrbALSPxXp3suoWFNZqf84jP2LpXPunc9uJFecLgX0
zpMQUb1EVr8nORZJZXlNDIB6K1+6wKpWg7mdA6dEFN5nV02ph7R3j6PxPwuBpk5AqAAR4Vkpiy1H
9uH4ExDa0Keg001XNynrp1/QrbqHPwA50ROLCV1ij9Pui+a0RvPIjXVdkvo4wkNdow/3kubQvkKe
p+TFRE/UBN1KsvHhmP3LB8PjTtYczQDIhrrQ/lHMk6Ed4mStm5ffxyZEbPdHt6H1xy2Je0Jujnqt
WmqFnBVbUiXXTja3rWCvHaPlMTD89yAeZJ16e/b7zIzzqt0exbmo28hiRDye/fKmlxFpFHKtXZ9w
O4tT+YPVrOhyQVWfwpN2urhfAuEiGbEf7N6py6za13loJcavPkD/0fGlAt5ItYImgm9X1iW8koNa
sKDwbhiFI5U0yesRDZRxoG49GUxTphv6GzeU4uXIefrJ/EbqPAfgMDZ6uhE+dV+JyauPHBkTynut
fMfbQrfrp4Os8+lwR9XWUDAtVZ8EF1+NKF84uaF78SieAGAv3H9THtOuI3awiXb1SVJ5XPVqJmDf
5OYGBjhbsnkEgTQSEpsC7kJ3qN1WnDJEPOc0gUWNfrb8qpmE4zfLB57E+ONZKf5ds9gOce3+wDPJ
DWv0RXgRCauUhgzAKhOVPMx2eI6Cm06OFrfj177mbQe3wI5olBaBf/eDWzHxekhDDxQLDR/QxqNi
t2tpya42Rvz/NIXffwEeV3ibgUYye0CvFIkiHBaBpraHYlnkOLv9Csq7CEHq3ma18TMAfYbRhZ7m
Caipxn2uRSRV8jMbjN8KSHrws/YuHJwrMyxtFJcUFEEsfso2v/KCKj45XkRKiEiRfdb/4veGveH4
ZhzaBz4CLKjvv8He0mLkh+HPHmrOUdcqhceqwearFOm6wShgrn4Lbdl4EVKVsI1TMfxbqZD1wc0H
/lag89C4uaiyJzqz7n44reYt+VASc2NhhAi9in6oUQj8GDNUUcQH3XHn1/yGMZMRo5UGouZj+UKg
m7e4ZsJFRghC1mMFbRe0XrBg9qdA2+pB9Hfh5YAUrxMerxbpjaKOFbwJR3YmMowe39gZgUMD0C1s
gWlhsLLx49L1jwCpmhC7+3s7ozBOn1asCbiFoW+NY9hOsktAylPRVD8JDJMylzXOJAe5CONc923w
v0I5B+k3mkgahgux9ducVKDVD8BI4cHbd6di/T910kqjCLJt0TtIxJGLAy/1k0zL12l5ZbGXfGqu
tuzGL4DnzxZWm1VHr72G6exJOE3ehai0e6iRHacA5VUHwsm3eNXr2vj0YjPERTVHwWvrwB9oSiMh
nfaIEXJcyTvwK9ZIY674uL9TrceunLxMYAyzKhNI4NVgWGOtmOZpcQhKv4fg3ntHhdgvtkXbCuN0
Nrm8mqunin9EZXrfGUG/7Q8kS8X1XBO8DAE4zuHgQgAxTtfPatp0Q+zOkOUxAEQ53ORKuA8t0aIH
/kRe4s11/HXFSaqqpdxQLnDxYMTkxZAmG5ePqPDBR+8NZEpx1khVElV0g1PJHxsrBACS6oCp2wYi
A0xMcQFkgNLau13C2u/u4FScSRYQos++Cpb19J5IG+dP+9Huirm8uqy7qdnD5hYACHthnEWks2UG
UNC/XFdv980H+N7Rf/WaDxPPCdMQst0v2k0aXezpWlqlWjfSBHXIlR+HjWXJAzu/r8bUBDkXjE8W
rxOAWjkiHeM7rtXaC0MZXb+S61OUv+AaiTnDr+foHrhE0BzIfHE7Ujxit0kaW2vpKbv/2yON8enB
NnvyUjIX/t1rDEnD/b61YKq+Q9g+eWWFNmbybjMl+wtr491nyMMFQ+iwtL8Jy8IkFYKmCSMVY51M
8CcHIjRW40oomtv1tCxgRER5pZBObIwv02AjbSL0HILoaUPRk6K67uQaROQKd73FfilhhMTOYyNe
NWddWm7MVrkqpLCX02XGsOThP2t/gQ/geryu638Cj0dP1zVfc+l9cxCmsP30PUebrHaOc3rhHGHy
tth7OAC3aKUS2aSrfpe1Y90IhPKGiqfaie5DcfDH+X0CIy0XpbK3ArFXUJFrbRX4X52p1sAe6Von
gWOMe9OMVmQjA/y+dOgKmXrQPg+3+AdubHG05hz8RopVgnh831Z7oCKrS+YGu+Ul8QY=
`pragma protect end_protected

// 
