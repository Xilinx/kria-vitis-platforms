/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dD6sJjMckNM/hk590wWgo7QyLBP7qvuv1GnV/mfQB0w/i/pvS4BJcnppdBuizaQbHZTE85H6pboO
mTjEC8kS1yUyaRKX4KpOmRsaXVL7/iV6Mc+EyHoad/3cx2lAwTCRu6nptqi96Q/dtiPbQirlE0cr
bj2VslWvQXYp7agPImHpkldpbIx4OKKY49/lmZgzjQmz1uAl0Vpqn03TZsorFhKrWNa1NL2PWEvy
H6r6Q2NnxwJibsxIu7/DaDQZ9tx7P3Ox5rT/+t7OV/sWKJMNsqkendhSkyxMCR6Z1Ip9YxyEItGS
Bld1ucslP9zp60t9CzMGZcj/WZZ+ve1NzjV/uw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="NlHs8opBWv2KH1hFnLsdY2EH/Cy8LVzvJ0P9w8zUaYI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
jOrE4515xgbASXSOIDgmJnravK3jfrplQ6x4Zodant/sP97TKimxpnTq9eVAEOxNchu30O/OTWnc
TYbcoSQBrZ3uEjHIcZQlEl+sZi5Uvz0JyEEl//lenxZSkCK/Gl2+hYnn4DHxRsYfNM+GqY7/wl3N
qYdqQ7io7QDklF5murIIK+hRBouZ4jOKNSRWC4fbiDoi4aOuguI9h8msyVrBaVtr4QfZ5BVL6Vdh
U6hQkYiXVm7gghZK1C5quOgXlR5Wr/vXCKacnPo+ovNSyt4OT8PWElAj3FzM2Dok9WcGUBfEAB15
fwW8UKJs8PMRGB+ZrnSIVDdUv35XSiGWO0NU5/GWby3LPIiYpmjKDs5xo/C8UwJ1SMEpk6FvNiLP
uiWDmFT28bhUeRx9+BKGGTdFeA7Uvaji8HxchEz5tHnxu7LCSqPR2EvS97Z2P/lcXQiqW8gqvch+
8fjzax0jxEuXsN4wCfN4nUjh0P4Hra8d+sUa0/SMMj+auKWPl4C9ZE41OzCEOm2T16scnBISMqlB
CR0fcxTdeck1lKJwfG5Vrj1fX91+xT6bmZY5QoXJoQLOgktLu9MMU93X1PTc+S7Bb9YNgwN6f5Zx
gnUT3KotSoI7M0PhoKJcZGsMYcNzBl57Gzn9tx2L50esmmquidKIOIw1cnjak3n+k27XarFS8Cxu
keZMll5PmgxUavfRxeUHK+NnH8S7rpxqoTPVhhRrwrkxbVK7x2ustz16qe36+ucUXY8KWOGMOVhN
jibjN5ee1rByK3lOdcPG0SGOY9vJmvKt0rOqr2LK0D/0zrgpVm7790vTS0hspCuklI+LquhxCwY+
t4l03dP2AR1h3xjF9E0CJVIJSiPd4QniYML+B9lgj70FabwHxvAI9hrAlWNL/WLYQU2SlqOygUZQ
HCrUzOn/VvgujBkSKzJGE/2KS+WmQbiXUeOh7TQ8tDjOkSug9NhDXS79q03Q7o5Lsm0EG27oOBgF
P0sFUVZIQwbkK9Kd2lR/vGbss/NjrM3NminTQET9/45D+RRS25a7eDLtUFNSYOsmWRAokfzDz+XD
FoNEbfBQERTg+WJkdb4VXodGsqSEXrXbimSC7DOOI6dh8S7ssTIZQ0HpFxlHeycS35jTVixOmtlS
7ZBqmQWpayGERU8Fn2/RSlRLGK6LypGRRMOlp1leKbIAFg5ZFIntVV1Qu17HOgd2q/7vHFvTPFgE
f7JfjPf1KqVncpSqv6BLgYLYJrt+0uqdR7choqxF9cEr6HYM9GGu5DcRnlxUcl5DbgKXyQ2rs3h2
kLSL2x/KbX55FNnOMxAqcs2civWeD0x9Vgrdj08P3n3D8RjY/EpWdb3EBaNYp3NseVMEmNT1cVYe
MjpvTrLZzhn60n8mG3MidqXK5WGLkAt2cngs3wBQsymHfHJmAhoiOdpwtKW8tz36RqCuJcFpgVEL
ue0jiYI=
`pragma protect end_protected

// 
