/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
bc4WnAkqx6dlMsl5fn3cAprcqqxHUHgVY/ImIQQum+cRAB7ouhGGGf7iFZf77q22uZ5IUqV83Quw
Hyk2hoLyHV1tsHXgJxRTk+FG0z8kNO9UiseME5aOM/+f1fcoxpdwoF5Nb9O6O9ouJZW/9wU+cOBn
deDxs8Fe2cl/gc7w+7aUoFn4WojygKnIaeby9NCvgShnH90A/5GxWomjUdPAdBRy04fmF471qpG3
rcDSX8G6arFIKQEh5UwVCLxQIuBK6e0cztUh2ocE1tgu0ybaWCTYOjp5wNkYHxW0TxCBiXthO/Y0
21pIqRWTmcspQgDYTjUBBMfo4xnplJBqhrkXZQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="ASJKkguRF7cNZtn0GfYOwaRh6RbIlcvsA1oAuucVfb8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56960)
`pragma protect data_block
Xy3DKr6jQ6T4G9Vc1bujRkO+/BQLnXYt4gYVs4GLtaZXt7vJdy1Ebz0iEgFIiuY4/ooAZBpf5fKs
sMlJuAgrHBoumUVbGnH3rBUVrurCXVLVE/7OEMP9cS56P6Vhi2ddB2hJxme5iHvIxovkhfnbQVwC
/Fw6RH/1pnEcyYpfHpkbtMzFUzwNgClP5GyqqETPmslUJ1CszSvQKOXzpXFiG1xozGuQH2FRR1FW
kdjB2X+vXzx56MXTtX9cnNaeWI36HGgm5lz+gACGlSN8qncowbPk3fUhQjMQYTV2yUjwZAXOMkyU
lLeWWJ6OqgGkxoKYO+P39XUjJJmZ65sehSpb4GBSyQqnqcqQ59wxI7Z4l9NB6oCIsX0M6t2J2jIL
ptbH37/T3VgkRCjv2itNyhiQCvp+VecXIxmMlEqvJd9S0Bi1iPC8gVAPAZCTvEbgmMLiugjOh5HV
Ijz4JhiepFawes+nPsnj+7+7F5AkUTzZn/kUgMYPa5E6fw8a/nW4G2qIn4sZYA2legiTiFZjbA49
BDtb3Cqy584dSZB4HXjYxaFgD9P6tCofJIIqm5YnW8VmHk0eypW9us8TPf8tXJjQ2BNdTPsmn8jH
g+Rnrb/yZ85Aj2dCXbMu3+hQAMgK3q6ivxJ/H8Rf7KdUTIHOlSjjyfg6DLerobZt7S/GvZBDqw1B
62WEsD+vPVBSU8gUEZFRHKUl30zPhz13m2OTsvwGXcGBVhyKPDDsd0phaCI8vI5ibYGQdRz218rJ
Sep/IwpLEBbngUu1pJFrlDMDUPZMzfvjGMpG45TSeiNh5zdsWCnpZkRsMTJawOTUw02XrXIcKYmx
ScOEqS+ACQpgADYPyv8V8MHzSGiQl3KZa90kzkSMwmb1oeuN0KFvYPTgPWZseUuAEue5TBWm9G6/
6YxyjHqB+KbWbNoMuFaVXG7NwggJAyV9Ciyt8VQjEK8mkcgcLC92MzSFx+yuvdfKjymUP6OcZJZ4
BBGnRHNAycrwlI+YvNJ5eI9kxRqdjpy2ZL+MAQ27mpEmlapJVi0C+L8Duw4kBp/8H5ZH8ORQXSJz
Ab3Cz8qdW3vSUG6QpD/zpvJz++ijIp3WW4sbISznodWjVnqCt56Q6vywjFkcNCZYMm1Pj6ctAuit
WvdfoS8QhhIZ5ojFK5LFf61GNjR7lopNNdG/EpBjeA2SA6schz80fs3q0e8iQ3bHBEhXbjQbMMjN
ZQ1aWXk9NX5fPEVpO4SKiIqne4Mgnph9nfgVzh9N1jxNZpzYmzuInN2hlzToxGMUU3FZkVSyJ90A
MkCUxzH/5ZjT5yCNGw6YQX4K1F167mizQbtDuyDC1p1824lusUO0GVOK2QgW5bdlYaMxQUmUpick
x25hQiz0GHS57Zn282iLoVgi2Um2oKFQ6FfNiISUrBx80WWq0OXtH1Fj6qOaeawwd/y0BmBXDXlI
sCufo5ViYNZTblD0DDsTshcKqja93OGmGSXPrMTpfZIo7cc8o026SV/JCbqLM7M3EWJou6z1kpyN
JjPUpzZ24BgzqGdsxt88oCGUw4hBdw/jttAP8jtziEjvE8QTfjCKx8yam7pV+pnCo7QxiWyEoEGp
rBlUbDREfAS7Yx17zKlS/OLeQXTDDzAtN41Vf7SkMwS2Iasw8Pro/arSm2lwmijLZ3/8P1rRE251
ejLPzaEkP9ntfANNo/OpB5JZp00wsX/IiA/fB6I7+Mxo0njO+nMYWZimcoJYHvvkeaEYNVatvW7y
Pwno4xgXj4OBfyZ69KdwT9ZHns8ob3K8XJLNiCkHYzwYSxtIsTh4zKq/LJa201qvwaxKjL7TX8NN
d1Dmzq2tvG6yNpkGtYNz46JKN2Vz/XA9Ne4YMf0ojdFj+x6BaXRZhmHKYE8cUnQCvdy1MzLr54Nf
NLPZAIkphYNQVVfM0A7Y4DZ0QzkGTiWojaH+boJHjRT6JCgYHsSvu76EfQi/9FuvyLZGuBy9qknR
ZfQ5JKjM9FrCo5ojjK0Csacp9JWPYG6BgkK4uo+fbkBtpu1nlh2ccNwNS+TT+Jef9fuIOnB58Xrz
T/Fnh17OexPVIiXhh6pGzBFtj4plximK3aHK8eTf2nUmWwqh29GSs66mPdDdMKZPixKw/ybsfCIb
GopLGsSzH8e2Ofg73Bs6XYybjyP/+IDrhbaMJt55VWpZiJPX1AJ7C73OO/I2alMgJNCbzcUb2BcM
k3fbRWUq10mJPt8ZlgXJG905hmllBUAQZxdMHd5mwdkDdlbXDJT5S/RtBjwaRGD9W0l4Co9reMAF
FrHGWgoMApDHyF9kM9VMexHCYG3ASkEmGzd/w9fWNw60uTvvRMtwoJTi9wEMEEaGkoJGZb3tOg19
qEsE/xoH3rGSAkR3V1dY2Cf+zsqPkuJQGRkbYkWR/eErmgyKyOnMQFot3G7aawYIu2889BwGr6pI
0OXTXMru9+lvMAd9ClfTOr9fJMRghuRoLyZp6I13ZNNMSyvAPeF8+s1lpSffgmC7vzV4rhhm5Aj/
Zs842Cg8z0dmBEAr4g17D/8zS6zb527X3ml5WVqhZJF3yJ37+F5c2SIuqTQo8KMpvA+ufbGuF2Ap
nPR8lD/ITxJHvj2nHPNFC8PXlz7yBtaNRpRX0gmmiXxtmzLqA95dKbY0X2vEnR1/iCtOPbECB+u8
J6OVO8LB72ieZLAb+loS7TWMnoORqQJ/Zf3uP6t+X8Z54Jk+K7+kJqCqGn3kqJgzUjCY5KxyC4vD
DYqNjleeX/A1KVSP6si9LGbjuQi7rqyBUHCJKFsUYkOX3Eat0Yp2DIFacUMBa4XubF6XAiEWVl+4
lpPEDlodGYODN+4X5OFIFV9lv4xUY3EBr20Fk5FG1Bi6s2m8Ky7QjQtkbsLJYvQFOgO8JrMhl/GR
frtqDdgjubVrj9jUPDb3YlUBb0612dnzE5awcfCTOuSnnokByub2KvGonfkb8M6gMSmgUprUeaV0
Arx89FpkNdAPThhm7ro2F8ce5paW8M7sCibzoqYWwUPJQx6EwrapQunohNdqd0LyUA1JNugpKH3R
Z2UjA+rYWFV9+tGlxrR05LVwJ9RobSp2DPWQe+fN/RWFhBPRXh/ha6OjMM0ojlLHGg+/EBBvUtt1
l8nbU/oAWE/QKDmWmkqzJGpSu0WYn+q+/OjtmwoFXkaOOT4ShZjc2ALfkLGG0oGQI4qMYpgUUmKJ
UeXYJzmbwo8Kj6r3B2coQVuCl5LCoxuMDEc3fstXOKr3QnAIZ1ozh2SCWkUmoe0dU1WM62OWOmPR
IMUIfEUGthy/YD7ev4zYEPXCMQCUT+ZX3eGWV5NSaA1oGk8kZezVQcV2gSJG5WcNKH6ILjoRXF9S
IjdU0oGFLqMp27UHUradEV+m1BovZm1gaXYZduyI7AYefdKeh7JDKCAJRPV1D9Q/M31Fzkjtm3EU
9uXWdhaXDASSILmOe1wzz7NyQYvCWEiSNnyfVywPor0O8o+8kk/wOZNpYBrcvpTxoCttTbPcdls5
gUSu3L4WgW6ETdjQEyBGI7CRoPvwYnqxv+r+ZQpzbRI9oINnHD1SkeduSIs0I1VhkzEzyWFg11DP
e9zNms0q5JPX4Qx6AcwW7f2c2LUhxQ5FYVYc4gMTS5zvHBSHrEwm0doXJCa6Ep6y4+Niim6TMSaf
1AjuH9elQ9Hv7RGU3FDRHJigw2dgXMEgmURMzkoiIvCScJ+IL19RvEKvMKk1A+NImWh2op8Y0lBx
hrMI9/ESQY8db17HiOzGN+kGhk8Dg64MmlglQjT/5EzMPqQfMM0q8XHc/41WAvDume1cBDJjN+GL
PT0wrUuDlXw9TdYTzigAiCj+PjfPlg3RCiIPiivjwRlaKN/uTkuY5HQapqU9lsR3pd3rvveY9041
l3XQpsZWH9xEd84XSiP1PPLNZcnwJlP4/+J7tcOipoVW5ltnWP/JizrGl0qh5k5KHydBKl4trqFi
yqqpNxUvSyEEzmcZq+AgCJOHw0E28N9V2A4Phuq7a+lZi6eDERAVHsgQxZuNeH3hIZ89zIrK5Odw
jiF82C61GPkkj6tabIjT8GmBT2tJf6BBAnHQvLriGC/KFwSnKQ4uVcwBwDOldp3GiRjR9KOT9+vw
QtEyOuJjSQzcM4lMgzCigP98lhzdxb6ItoI12W4i5O/mgJ6IlsUpzGG8b6bHnXNcrEMyHuYRe9dD
XIzdFUi6+J4Fq6jvYRi79Q/rbAQldR8uMYGS7Y3mS40EvlwH6BUH1FAHgK9B+HS7CXJXZxKa821/
90251Hy9eTbjl8upiZ3U5fU6O3JGZgw31oC9fBCqMkLsSiXlADbRSTdieV7DZRJvQOeh+7rhX8NJ
4G40VIOkEKEcUsU87HYnUQskeSQrv9KASS9RiiIMHkVIanduJTG3M0svNQsCy7GATIPf9lRbsm1j
v4FMprxqobjvpHLzKUUH3q5PqYjNU0qbeJ7qh1td31kXdqdLJv/iz8ggmE8dAX5pxPn9v2llw004
2Jo30G4wDbDyynaUdf0Dj6TKrlz9VObcq2SUTOv9DDtNjfE/raDcGeRVoZvgkE+H3RCRhnbQxJi8
vNklJKBtzvJa3jAcpDVH/KWEWBvEsB2wvH8/zYMGtDylk56QIHNoz9QqVqa/rPPa0Is3QD2kIcvQ
D0rstBgFagy/YwlH4Qh7ikz9bLvbP4wQneBMeNTwWf2a8JfErjD0aofO5QwsuMWFL6piWzGfO8om
Im223O3okSQuznVnL8KHXZu6djlqREOcYernhfnz1Fwr3Uy+9e1eLNB8SE1euYoYLYBrVmE/SZk7
AyU8ELo0oa6HSqcUTxGAY4NtkWA8qgAj42dMngPgWTx4yPrFFzMr1rkbklT1fTJEBvTlLfFNy7gF
3gVlBwBVJlMhfu/3OST8nTgRkZgF8PWya/HnXHIb2WtK2Ny9nrpSAcqmb6L6u9rI/5b7jsvCaKw7
QPXkq6qqq4MLYb/V2LI2DyuxFfxWtcPA55o/TInglo9uDAlXJrcvpAHzG6dWzp0KIQurQtHEaQ0l
/AleclSeh9tDXGJYA+d/OYUmACcRSnAiX8S6A03v9sZGu7ZqF9IxREIPSbdcysiwbD1h8hUDcH3b
l4vwG7FnRkDHTS8eHCTaPJbAiKKKBSp0gLeKgFvwArY6EZGjztyJcL6nmc9VFmeY8kMP5QgKo1ei
2tBKIWHBv+V8QbZLhrTx3Kn7awsOKAYDPeSI8HHMlLsWMlBzQWv8tdzXBGIqR2UjnVmirgQHKZej
Tfo8pUMGTQl+bH5lvrHxsxnps3h2lU6a1PfF37DkskKlFEk293k1+5Du3yXdCIC6QtSvyvLlExzM
nRo9jeVOjXJkwBcY26uL/WnO2NIjwIZhXlApdOxKrR8YRmZicNAzBBtwB9vbJi6iRGcp/wZ2eTPW
w6LhRtwBdfKcEJRh7r+Dq8eMuUza8VcRZUEDuwRdVpjsy/1lLMGqs419AvHG2nyfxwf/NAlmixu2
fGx3eS0ZYWkOR5dY1EAcnInZrheyK+w4Aorh2KiUbFbVHCwjOHlln6yfsm3GQPb9bs9iWm80EtWR
yi5nm0vFJ3i9hC7BTIkqTH7dOd4POeTo2lSh27tveEy+GoGuXurRIclDxKQKBwikGZaL8BGFPhbL
KGlSgQNdFCs/T/gVmW5qhbxetkKaLkpXyfNZQDZMHpT3uRBQ61jcfmPR+KfMCl2JX4BJT6FD13vr
UbBaAToVbEYfRNsOrU5rlktxQQ5MyA4HqZE7r8xduuVDFbjgHCbi+Aar0ahNGVEyZigOcOpPRkXo
C0IkQez1NYwUb65BBQ7mcmcFQ0ZkeUsIZU46rZFuo5z7UFtgrNvJG21Wl2VRQy+Awsa/hAlhy9QD
nl/brDI0fFg2BQoF+qS5J3xWnwWDUuIdnhue/9C2JxK6QEvk9xc3t66Bw6a4nyvtyGhdFErur1Uj
Fdw4mCYGLSjApyCrTLEdVRYZUsqxQ8qde3m1WimjFcLPUbXp83FY1Cce87Om5YtiFg8Ei+w4y5TJ
7POrwrqxYLX4fqEX1ZM0SM9d7K5DISPEfNmZ9p4qEO4Y1lx8Xh4FRdpnE1b1lIwJSTLa4ttfGCIU
L7J1nM4fC8qzP9xW9WFE5ur0OD++3xMMwA1x4DK4a+VcLm40sixgI/PTSgShCH8CiTmx72cuYHaE
hBhrjHJ3gmQzId9aL84vfpCTI3hg52R8E6G0zv3wtGLjXQvMWAXAfN0a3bD2QiAhcA41F9jeggs6
5Zi+THZkKc1KD1KgzJkxuZVPQPc4QpLvDBAhIz1XdbvceU7eJ0cwQLXyNzbxFtr0gAfNUIfqHspd
u8WHn3KssAbtystMG1XmJG4onkUriPPfdXj+xLOYtsrBFiRCRa0xoL+q26/PYRNhgrkQDcTN02Zo
MRrf8pjY0jhJUCQNwpYfLAgY8dmUaRwHrFD36OMRc/W1XOlLMs14jednVPQ7to1yMKyAet3fOO4C
SB3NpWt2YY3tyyByef1nn9cNw/qBKL1exTTKogrL01mgQSirg6wgRv3D4h1QBj/RcY2SwtQpUhPH
mL7mwt9y6t93EhlKK+IT484rb1qQ0yX8YDs7kuPsas04XbtBbz2VQo6U/E5k2N0Blb4Aa38B9RTR
3kaXa4ZmIlnLH05eJYLan+c6tsSVcBxzOoOnjG9AMF9NfvXPGj+cTPDxb8fvGIQwRZOhDnavlOrd
IxsfJXw4KFxhrHzkWpnM8CMzdkmai33iSYW46N8Ev5h1hIb6M+Ey2mXlmVbvt6UDZzQOQY6rEkTx
zmo/ozu5njfBpf8B8txr44VWslGctuf8hkl3pw4JjLX+gdiyfarFR05YcbQtMdeWNQsyF4AJFv2I
80KSYXKPAjCmyt990tKJq2Pj5pdpMz8Ri2ULVlMSJZuaULTVVpj1BAj0od5Wf0LL9wT2+5WfMMEk
v45zEITjDfv7MO2Q5cwgqi+HkEcCookZYwuFxIisICG0rwckpTPwrcD2Y5/p9wlRM4wOsDps85IL
0cRNwOXCYvhdtJTr3nBc81LZL2hDk7TM1stkr+X5VQTuaD7UE86UpwSCL6ggcQUzSnxC2GeSB/Kh
/kaQhlxWvMmJHNyEmZWqQeBT+VYNeHC0+iVavd09Rmc3FZwkbojLNkAxtFdtdPHA1NcypvJAHuvv
KEYcNGMFEz28nU8kBV3v6w7rhl/3Yif7h4Jvn2Yifdd+wpU6hZGiD83vKqsn9d3ZEtemZDSv+xzA
NgRjlYeGXHJAqfmGM5v+iFvEwsQB5qxAwrtXwQ2Vnqj2P4oyUKajaLs8twya2m/OTJdSV+5LVMAv
un68gbtSr0aoF7YX4J+irfotS5+qNEFEyHiicJ2Cb7/CJWlnsjlS5Sazr9kthuEADN4bX8KzLu+k
h8MNELKXH6dVx7Dk9TW4oFOw52fiCqJhTzidK/bUkAsVe4twqmP91hKGsOJ5EbTUqYVgtJhU1tGB
6p/Z/EdaakSgxWNJqRuwde7zDgxqrLVWgbFu/4Jt8RsipozPwzwi5cwp/6p3o90EC1wLS5Q7fr2f
lD0CgYP643MVEySm+nWwcujf/i053LEv/YZcSyFeDsU8edxk4TpvH55Kf88/yG+7ePaLXjcCDN9A
w7rtQHslzyT5Hd0AxlXwJeoxjn2Birzt5OuJb9uij57TSRnULM0Z2gbLQ/0f77YmVI2BoBKp8xhm
52y7RqZNDLxROng2lnaBljQ0qD1N5xPr8AZDBZT99xMCIm5jZCXKD6YpS8T6Ob3hn27zcRH1EbvJ
v1Hcw2QDw07pAih7HZF5VdF/APzr89NzPSWCCnBtNNsXORdHBwcu5eA2stKrjl9BEolhCN/w6vjp
DzXL+nLHhfQbu3DSbXuSnvj8aVpx3ob0IXkf4xRQERDV9hOlMzov2xyWMilIVATkpAX+cy3fRk1x
4Qhx1LzLmopPXoMzTtMZ4LEesM97fUmL8k/lFQ2W79fREqQyGiRUMy+ByP5xNbv0S3oD2Gap1MUz
zYxLmkjnwqnzPWpuoLx5CQ/c7tmcCtwOTCsBtDObsYIijJPPv7zjZ6FtxzYUaoUacZH4sC22phEX
p1lSrxilPR7ciTQr317/0U/FZB2jxpjys3fz7yZYz3V/KskeAviSU6+Q9kiXpKdB2Lk4ncPyXqDk
bo0bVLdvJ8bksAxky4YF3oa1if6jSN62m5pSCBHSAk4NbehhcQZrFiM9Vo1HfZj5sPbeaj4V/DPw
tIbqUKbzADRbgPdj0OjGkbVOrePY+GDdiJNpOMTWOI9CgGiDQm+acwUH4yAAI09VYbSs7IN4UBJM
y9nOkkZ0KTrYr7A+cSLq0xPcCFT+4ica+c4EeK27f5jBErIvx7V8r9wO0XKny/WEy3+KFdIvEqUn
ccri7V+s4ThlVPhHB7BeXDgVrcWzZyeJm6se7KVwPX0uGAHBUSmIRFKQin3ntaFFNdCo+6BzxBrw
M2Qup23UvrCAhv90KmSdIwunRWRBQvOOi+F6EopM8eElW8t3rfWQnFlFep1ET3VPQrDF2ytHLgZX
j3pWIn9TZdNnKL+ni2DtoOJgjOiS2s90R+JRZx8JwVWE//UFbwoE5X47ZXhbg0LUBY/+QphWjXS1
UP6rhMunvwzIK2CDue+56MRziaUiBIAlyFWtfcSaDWrLGlpaWXTPCNOCiGVqkHyfhoQiW+i9i9gT
tXV4olFRwDgh8rmf/lifrhDkBH1aLYypl53U+0qBYat76QQjt+MkEFl4SaUqSd4Xvv+2s+9TtPhw
PRYY9XFOiImacCw58StIFC5K8CcohGrUJAA8WJyTuis5A6DYIjydbJR8OZV7mW+x7I4L8d0/A+KK
jpFKjJUbLFXFa6v4gEtnLnNwgVmJLIotV7QtME5ePEOgUpZ7oLvs+uA1/05pjVcFwtZ0n3KSG9y/
hVo/Pp5MUuQHqs0MvurmWVCW2oLwUDlKyBngza5mHhujiDrXHT1MDRI4MjMSRkEPgLP8JT+oVmqM
/6sAKMuRtk2NhhnEi0Z+6B3W52vYwZNzbCHg4YrHWa/xwF6902VS/fapWfwZiHvjs4MjnLgcWjxm
3qvBILFOnk7J3uxyXIECm4rCM/n68aRECsS8zjbaCt05A7ZOFHpSYK1O0s20z1HixHDl09ndqOXh
S3TK+sab062YiXeaiCbU6V7OGHIw5wpvI2T5x87FUA4heKu5HJEa+aeLqwm8nyw/owX7QHB0loRY
asq4O7CLEM72ppKBTaa6A+9bYwdpaqrQe7UclR7VeHHBCXZTF5SU+F/wRxY7ePmttbRrVF2D0aIu
Ca1T1R2B/0WoHKDPUEbkCHKjdLydMgY2dXQbjWc2qoWeVd6c3798BfQSnAGY70vAZfQonXQJSd6a
PjNngjjsVCIpaHobwtF/l040UOW+qLVTt7+8l5ZGFOI5vbcxM6WCUpOwb050Meev1YyuMrB+vh4k
TbDLcTATeKyL5uJuGzNamG4jG+3MTF3tNzQNqacPM9V8IDVOU5cL7EtfPZKVR+saj/beqfr9ybIT
KD/oVih/wbVWuzaIB2gbUnjKpztzdNvpLqWB4oY2Team1lYgzGcUUrPPi8MYVu53f1vIpeym1QEL
BxlBzGEPC54YdMxvJFopjW0Cuw5MtHayOYVgho0HkQR26Pz71TrUxeqmxwZPZfi7qyrbEULDkfb2
AkYMKUB5f1Bkep/jd2i0qu0lLq0DtssrllHXVXnxpiHYeUERMW9udQKdyo9YzGdoFPtLO58PTz7y
9UthRfrCqsmnVxksnkSCCO0JJ7+gMUaGQW/J+CnKUXaHJw6ABs7L7VYpvlm71Z3pSuYRfyEOaqKm
Gn5rSqDt+Cczhones5209o+NeakE6bmWgnOgnFNYQl2A/y1H2oNBra18DQKZS5YooF8eWrvJhQ51
nRr/26aZBEBwQP8+H7ooRpKGH6i9bkg3UYcajCeQykeHOxDz3h8T6qJafpg1lh99y4Yd3TFzUUkH
BbTgMoGK9/Cuby9fOZ4B0YMUmfdHc0TN3P42RYQ2Jkiim9YKmROaPJ+nmp407d+Vc5XOYRNhyoNt
E1jTXwIGWaO0C0aFBx9eHBORnwzw8uxp0FDPvttTkmDq8+xzSLRJQwbrYSqf3uANSEjrJobPu6Eu
NUpb9xhKhmov1OT6cpj3qzT0QHBfFiP328vL+FFGIcAKD+3ulT04PGxBIU96fsINRRlZIYStgQ51
0wDWQ0Mb3Tjd+a98HweOKrjA1rMcvqkoRyvEefCVMHwBpYRJLtcOP37Ev3xKjbq7MkNDamirUnQQ
amsvUCufE2Ng9DLZGIiEwHr/lx76MVfzeYkNMwOJqoG7M9W+zyRqDy7OSPtnNNAAkApPl1y53hBT
eJg/PX6Gf9kDEehmcoYJRw1UmG9zhfLgNp/0OYsBADr+m9wHV8i44vFH6SuDPVcmzvgZHWivy+Dk
Wo0E0yxxCf3L7GTUsR+x8NBz70gtvqfBroMNnC4HdO7zzvjFK7Z/bX69f14QQt8prsxcyq2mwwYJ
pBrtT2HI1phPPTGAWXtQnXyIkmbBO7kjbYc4L09JAYMu0qHJtwSDoJ52rehzHLJsQM05Sz1YQkpI
2T5eMLqTKiEIRz6xY3Lw6Qto0JSuDbgywAPLgv5FOeRH7xlhNllm+sLVFWz94BVr5bG6DekuG5t5
kKRRg0nVyreHrc6ox8ZPad14oQqt5YtBlvMfxWe1HU/2Qj2wnBRcImU5bT5JPY0bf6xmOW5Fhjp5
MnAHdEHFfCfBGWuHUM1+UW4XrY1GZ3KdpMJDoez9d7azft9nZDiBgUREbZK+qkFtI4iAfxLE0gK5
Otl+Ejpa9vY6T/J38A6cgvhvqgtfcMRu++yfngUj7MDRTslHlNdVM4ihrKZNxbl5+G+Hg2Ga1wxm
/qXDVWTNyjtOkx2R/AGNflaESNNfzi+1xy/9yVty+Y50LtT7j1aaRR2y7YVLTqRajytcCKOBsR7p
hNr0IuSwWapRE0OC8KsNA5K+q4l3VJ4/J/ZuuJTjZCctkZDp/FsZwJTTBa0DZtzfk0rPXiuJyR4U
pGGrOqJakGcGz+WUM0oJTs3l8DjYOxUr3KJzzOLW5tjUvcoFJBPlavsTGINr2YvID0PVDTbiXVok
TGGaORmLq//s8wfklxB/oJrgbt1tlh8MoQufIoi9QecHVAA7kA5U0HQ/zhMLnNROjK6jNNAxS+YO
7JP4Ur1yQLPCi9sYNQ6dvZolTvIZMNwokwS2mVqp/26/W1MSc+q8g55WVGEcSpixBoA5gjP9x30b
IXpaF63ii+zUxHf+2zGEablQ2qUVXBfrpJAZZap+hvQFLVaaw13exJXMBPjnNf0fKKyrW2EFkIOw
kY3o1mP/SQeVwIJBoKbA8qefblFI6vr1NIrUcR68UbvME7GucknyTmJ0OUUnoB4MyfFXk+qCth5G
5sB7+cKmAAkjvmGf+GnW9UTzmlYinwFdC7bI+zDNq3hVbqF6Bz76wsFSAUuW9vkMtJcUPuGG68tT
C79lLxoDzh8vMwu3j7kP+NZ2l2BhgT5ch6v5m4MpPwQ3xm8KbdCvG0Ibp90xzN6ugQQOQXtkXTc1
lrdOD/UWW+BXdKMWZsS/FM3bZC/CD41IFREWc2dvBS3K+M6msYIfAcPN5o9WhzRZHKkodd4NsnZJ
7eofmtaEZwHda4ULIzy7/TcgV1NcF/Ot6jnz6wuJAnNS1B457mmLNg0OuDw+1SMpwaaW2nZ85Hpg
nTZlH6iaV/m1QdeJrXs2F6HQgSsMwomasZw8H7gkthl8FbGDrtkMsU9gQ2nCcpMoqnKJHigMc2Bk
NZcQxGyi6NIc7jm3zAVIzJJ/e5TwFalbcqCeJLNtutWzCdx9b/zdYRI+bulPtUQJaOKpyZWU3viK
F1l7DLm3Tqfw7w5YU6t+kDo3fnOGNH6JVPoXaUDnddgmZJsgaQAOQTOttzAC5VLl/aiTNw16hcvR
XHxeXIg75I6lcgr8LRhtpJJoGTGab+Lm5PA3BEaRS3PYAFVEBS4Uym+PPZwRjhromRALfnLNA2Oy
VZafIaMFtGX3pFCyya+PUS0RCx9G35112RvUZjlIkwdFZEFBBnJapJPURxBEI6aJoLQqwxfhD8X2
VXZdZ2Z1h4rgWvJHQ53QL/gtZFaEznBM48RfooK4sJOllNTzSVz79zzVs2KAvtHV2UXVy9MTVZku
lXIQIFRFxo7t0TNuFovWcFsQIKWpx9L3VX6UeiRFzwZ3CRevhhUcR36IJrrdW5ORrNBSzUGWGtCj
8oVDqat5Tv/MTmIqW0gbnVNY7cQcJTiWXC++owB6nKPvd8lWYXiuBiituYRechl8voP+89c6F+rS
XKmBkdU839v36M7K8U3t5OXeHvl1ccGnjMh8a4g8rl8WXGPo1H4xdgO8O+qKx3Czr/yRg3Tz0s72
0P1Z6LW3N1kmcMgaT3LobsJkSGmAqAQWH55SMWCOq1MDAp7cewhXtMy7pHr1+FuQo/iUaJyw+xcK
Vt2XpUhV1ZwLfSDa25pLTHDxFPNdIhEBcR+PjTmP+8Pg3IdziuMmfkqSYJDKfHIoD9pobVKOQKfk
tc+r5aNeTUQHpFrTWDe8AFCt54si3rzFd0kBSbfnZlp0OTpLw9qwXwpyxj/wmfKzgfnZn16LiACZ
gFWB6hzid4SsBv9O/yxyRNQfnCb12dIkDPwN/LLQ10Ifz4IOu2oHi+qRxK9uZA0EE6mdczpICBwR
IXeFnVjohR/MoZ0gTNE0BYcjHXhdn5tcwNCMYKXDMlEAOjOs3g0BYemJk8tglNLAgUG2k+GtgZn0
LwLy8NZPe6z6gu3Dke+RnQ6i9AUvaqJJEpNTKwpkya1/s1hqOwpLbwT4WEJR4avVVa5uQlCYTAad
hQmlxwaaJ4rsYiMPmsZSdDeqnHzY6888RElJuxAr4qFefFbzhdue1ADPoY0RS68pDqvt8FLjfDXh
CyAwtqgvyYUhwcnzCjXEMYKEgrcAlaqfR1BhRwJHr6grhaJ6Iu0FWpd4pDHba8/bCSyExslBTln6
G6BJhlfANyUvHIRhSKuj8CS5Ngxg2fpci2u/vXfvIcaz3UeexqXDSmciZ9qJ7B7A6ARgi//fd2NW
Gj7SE/cydbZrb5hIN0US24xfevn2J+uXkxHZy6+xOs55/ZMkGDn9mkd0gD4LTmqo6f/EgvFNE+4V
2EkEX+uQthW0Ke4Sfk4GZfd/psLW34yY4f8CxXEIq3Kvs1qsjyxbGZTKQxwSfQyVV5ti4szqYKT3
IdGrnwkV6f5Gntl4HGbon8ki6CjoLC7xsYojBAsrwpv3kcVAaobvFhBPKFj+NIxnyv4XiJs0NY7g
Q3a/6hAzB/A4V8rSehZXqN2KlL+IZBpjvoCFcJKWoHWII3IQga6DDfqtIf79Z1rqu6a2OtdxG9Ez
e8ibKAv5gpiB78IDzRNDa2XL1BvTf3e8axUCjd4hpcuMF3tJBMoHK540Ew5e+9ac0Demcc5n7Jzh
uUoodODBBzbYOvNAoSy53bEke8ZXzkCnqDHSqRp+QPTSJW7RSEgikwqqvJ4TAdRB0Kel7lXT03z1
i0u+gaAbEodT5lAhwRNWWyE0a1jPregCVg5gA24Cf+gbJ1q+4N+WKVjYL6t2CqKALq03CrrdeSF8
hJvbvT83TZ1G8EFhzXgJSsDFoH9HwzxlHthN/cKifrdjMAggOMVTLFiNszMZzj+hDHHayOQiL8Mg
d1YEKdvGyV0bw/L8yr9KBYKoU1VKyA5s4NX42HU8dmt7PJWcBCmBt3seELaQR+G0FqnzsFpyNGgi
ldvKTInNdZnPkKCV9a5HBu4OUEN0jVzgF/Snh6N2DSbC1JWL+lNx/iUVHhYSPTJzP0KC3O+kI22F
Q4ACHVRVofwNkrulwMP0MEB9X0/lY+AKVu1TEjFN9vpor9+xgnMKEIeWs/+PfFwYxkwC2vshkLaf
R2AGppIape9eOohKrjcjRBHGF0zzjAH6wblkjvKthgUkZ0w4Mai+zz8gOetF/xvhBld1Zfo38wPt
ehSmF/2YuYZahs5LeEAI+TIqt7BI6RsB0tr1Lgmlu/iQyjhz3mwmNSMa9Kwb752ofKRzYuzLi3ym
BIwdO9oU33SS7bvu9AAD7uWkyGxtGyL8ZDHMDHKqPlFJXeqoZsYKe4YZCTatYJgp24Ll3GgF2PCf
r/N+NaoemaGeQFzkLFoVIoIQspxpQbrFYsg9X/NAPKWsy7ob49AcTT0xgBOSMPSvP/6kRjrvtzaq
zXN1OwIIRR/WkaFsNwLPSK2aQafAa+1qmYAM2WteWtPqHHZgvdVj7KjJNPavj4fLy7sD9qVXDeSY
RPhPBmy09/Tb2KkrsMjLZbKKCvxKFaAqBT806hvvJmYI3rr9Gx/8seJR438+PS7UAxRprL/q4Zwc
kOM4ce3Ogxa6K5ikKxQB875dgYbbwOChrWdXilR6rsV7S2jleLzOZaaugO+4Iu9wHWtqZFC5/nT7
ixJqzBqMQGclMHjAtujjaPYbt1psgglBLTpQoj3ozWVEOtPi3JasT1M1YbJRni7Gm1+5BKtSGFfY
fITE6mtyNMESymv+bF/AyaXA/2xfTXz15YLIMdul3AKAM000JChNE3SVTMJ6vq4oPGNE6ACG10mM
Va9u7VLPF+NiXYfMlb5oS/0xenM8zazJ5DnaYqfxyWFVpEnT6hNAGKC8BWM0qJ7xzCtqJLWjZz9i
JYAjz4KxGw506/gQDGvBpQE2UhXP5PNAgJOfcTdOPxLx+YPrDCUoWbYoP1c1C+rb4aOLAID98ice
KFoCJBFaO1w0LeZS9MKaddZFeezm5p4xLO0ketMr2jRY0aZpltCgBKrO46KU2L1vd+lkcLEY5anl
dGzq748akrv8wS5qC0ca3UgXw46TO1ZEVtbZzMexu07PnBeHZOtUnD/X63RDiwuzWzUeHd2mh2Px
bW2qGx4tJ7tX66dYJbhGXPXALsEcAr6JD5SmomGXhO1t6dltoAx10cBopPMb352s1jw5aBGOF6UA
tUG44MHBMCGfoyfXkhpHQz/BkEO5q/mHfwT9kkbFfKc1ra6VMDr9WRow1Gs4iuL93bIMT8b116AW
aqXoGpXbry/e4bV/MxUJ8JhD/mprWs+CE8AK/RGCc28RKETsCQdQNTImwylMVGPMhJ17nCiKe1qr
/zQTUKxzl+dVXOizQj3zWXKdKjQeM8jRuAXWE5idhObE4d7fx9EFW/RfuhTrkG4Ab8TUeK8s7+d5
fEF7ga8STlD+vXHgDP/7PWOG4raahtDAdXdb3NLfyk0WhBacraMayi2ZRoVM/2pXU+aYnToCeGyN
LIJpvhKwfifQWPQe2FSXwlR4wph8TIVTsZkSuSogTZ9pB/wAh2MWF7Q+FQ+K58Zn2YsPgphrDYOC
JoSRkJMZcyEmb1g6hFiv814oD6m/xrtWPe/G6YBHHGbKe4O6gBjVIewCrxKfqb1aanPUO++10oCJ
ktLHqIc17cZHDl8kew0akMAA+qlAFOUrSDXrhzXHj2HCDN6GGFns76odIpvaaBc6YFzDUySazuTX
7FDhtjmNNyyg2k3VoPpdvdMHeS8Y77mVoPWvC+1GILOivM9AOTrwkVXDH9ScNYB+dsP2kjnSyEFS
wx1niSmtI439agtC01NcDtOkeGTSQDhroS0Q40UyK7iCAHV4k+ON4jXbhRkj5bjEaJI8C6BX25sa
LdC7MI3o9n5jUtbF5FNlvB20lnuUSQZx8sv5niY6Bx/xFub8fSUsvCrSS/RqIFzYgYNAdkvvF+hd
jVKoBG2jO3JNLaDMo9m/N2UfwWv3wXEn8M3KLaYHNLM+165xMSmmHIpRVyNWyR4F8YE6hNFmibgr
UqaH104icIgs3MSbVRsjYTzeq4uSkEeDOSTq9tDAMVJba1YwebdSijemrSaNvNoUU88BTZLGrxNW
stP2VUR/Ahovm3NIIxPZ05KyBxjIEZwB19+GEIfkgrbOfpt7VPwuUibPydn9J8xfWnZ5MB93BXHl
hijSJHlrzNG63FpFudjLlGPzvSZs4sReIM724i5Hhu7+N7OARNMJF/cuNnfRammKKO+UCEqIC5s4
hUoAUK2Y+BLm52JsV4iadfCk37kkZNjfigJJVZDSiB20WhcEIddIru/fQghT3/5ftPzgTtorLsl/
eqmxj0BZMWjQ1VYVRzJi69Hg/tDfPPHsjKRJ/RBu52uVAPWYyCt42HIUGtufxePcJbNaieJflUhv
/gjuBCXwlbnkiiymm8SMG9eggr86bGg3e+J1UdJ7N9wys7rebDr2eLCMWxCSi9fQI7valHrJAIze
r5tvKr5aIcjExyFJRHJKmyj+A305O0f1PT+1DFLG5N+9V5IlGQtUC7sGmo7I8apSASaFt1Gr8GqB
gdMU1ZuqehPL5at1YfUK5oLOPISQF5YtDqPpbdGAuSNeih+6r2FXfxXuvqTWmqYpbL4ZahnAbDcu
iPZ55Oav60Xg8rkn4hJNd8TP2eATa3VqKVV3Dei5kh0Xr/g01CDS28hC5MUG9iNGs5PkRvMs8/Eg
R2tB2YI1H7ATxm7XLzgYIiNCNpSU2m9CHZ1b6PaWlVn0zqVbzVcwpFpfX8SjOUzLjyR3aL/omi6z
bpmNLKfoc36ApmKbDH0WYoFm3AN1xlpLc6m2iKsbr9TAtJlXkzVOXRyDIeBvs8zvSmMgPE2sP+KH
q+vqbUZcwb8jxw51uqWSZYivopPZfgUd2zpnsfIyZBCq/HETmLzoSXXuu6fqLmdHGaDg7tqlbEBS
bnxUt2oc9C6Ff97Q9p7zDtWoxjRefHQZZUt3sTAZFkzxDXqebHG9u666DqjW3Xpdeg+JczVGr+9y
qs6tC4jQCzBWXBa0xp2lBptYHxw9UwLGWYmii6dZuouUxfS074Yj1dxfYEm4Ad63jdqX8FVYvjib
TkZ3SW6S4XWvbg4mjKD7b9FuNiKVYItz4x2R2NUxaYCvDKqvBcXngNAjZO1yaxQbh9aJdc2h0nW3
PkpEfGDmSAV0VflN+fStpIKzmH3NrJ0RLJTlBZdDrj6IT4hf4qIAwF2ycfBwygMlaR6c28RDS4TX
8fkIeXzb1gzeYS1RWpyknCIbqlOGcUR0twtWRpbarSKwJJYf4bgzpF69V4WOytYR+DtIaAuhy+09
uWsCIFUjuzGpTIYvy7Xcp25885IRQFPxkLudm4853qHGhTzM2R3ypbiiRz5lDOLtWWv2S0kGAne4
becJIrVu+t7se+oSKocYIOBzQ/4TSGc20TCzDPg33kCaOXuAqMkBU+MKlLUhFs5dH2txlKQAXq48
znvQxPMDWbJmH7UtmUM4UCAgyeXt5Jo/8x/5ZRFXrKaXMbOnzkheUQuVijDn2WZZLzVS505ZxhWj
x9rsC0FpGaT/jf7+2X+u8i5GZmuazUltXRsgEtIdrB2VacNdtZKEN7uVN6XRAl54Y11jZbh6EkEk
bp3b4gW9BnURTvWGxVUNoJj0bumMk1//rP6x9WoYS3uvKsfjeySG66yevjj2+Pf7N1AVEEfVFVF0
RUKIXnhngoo0E6W2fFwHJhy/wV8F3x8n6Nmn7Zryl71QAjbTzRK55dImpQKud1FLoWlrrRzVcKel
/YjVHORXCUZ7VzRhgP466mK5HhRNzhgZ3IBDITcFYcg2hbv072d64z7B8iP+/fHJZwbtvOduAzDI
M9Gp1eZHy2/b8/9KN2CTVI2al4sOTa0H0T2FlnpKc0cVt+1mYcURJ74EmZsuDmRdDDIaPMzgccy8
OH0KfOuqISF0TiNElQ1FuyG8pd4WXj1gJG6vmJ4ni9ttcbxEGFN0jxdvsj4LAyrXJQhRbhS/LleI
ga2mOELgxGOVWzWm7RJ+HLy91izNFTh752ZL3WjOIS+8FluKwDpyPDL8Eirulg6K62Q8nkALUxrq
FquQH2BApsuhGz8JVvdDGUGioFM3CtouJdj/7ugwK0+RINdEnUaDvjYydjCf42K7fmf8lVT21SwK
ehOT7Uhmd8tPdMQrObV/qoM63l5FFzXibwSFE42wzMibfmwLEY39esYLXPPdEoFmPM8gqXFTV40s
2ZN+1oqUXs2owyh8gHxlwX9C5HQWCT0ezE4BeoLe6cgtPFd/tLcMqlCTrlexSICWHCUCGseDanxS
3vDBmXMs1NCQtWBQKa7tXTKgVgd+2XdCKI6MA+EySI4nOAO1LsCeIJn/JcDK0CjIhznloDL8rOLu
b8TpUSujsWIQNdrr7OI9hsq5kAk4zI14xR499pdRJe3xQjUIlMazTYqCZ/EJIioZoRRbVUVLa3gy
vt01LUUN/XSDjm0KeIOMh3+G0e4z+LDEMhBipkYRDsorCwfWVUZY7Y30eYonFEokcDM6kckAbg/x
Hfe45h+SnerZqwsOYFm08YfdiYTWUiU8FU9igBsmojElxiBzyc95ZJaeHtrSpEZ8J+vlLricdnxU
/pwrOHrUXNvQvbLxwed1vARsEkVmzFosjcKBGR7PF4SvnsXL4ZV3shVeLmmAlxVxT1rgfwRwNbA8
q5FqUpM2L1kBOy4jIvxG0zDNAKJ4Eg+dUPjlozWbDNmWgtrRAXb7TbxWh/pl81VNivamdeN/6S21
Fwx2XJEaCwagBRtwaZ/4eJNaUphuUkK+0H50PbSM3NmTS7+j/3JoGluyloG1D1F5UQbzEmdCMILs
du1FcL4hSftGffMPJVEgiWFs/9A80YxE1ZYt7ccO7RoZA+PdETfQUhwwHicRbRaLi98wx3WXgMD1
zg+1SC1PyEXdy+R+A3GS5SyM/eFhEae/ZegaRqsQhZeShKcv9enTD7unWJNsu59saPWxW3+TCL8e
AUsMVPSvOw1jMDFNHJod6760e8ERJcgu3bPcanVz2Xbk+YsKpxIxmU8KllH0MMLITxDstnL7Jqs4
6DOsr/JN5samvYTNkBeVyTg4Uex/zNn/2ZFw72ajwdvbZMhAYK80qVMZslKlViXBYvJdvWi88h6p
n+jcOD5+WTbN6uD6VS0xuPLHMGzibMhZXKUso6P/VteXLYoxKJugnLZprLMj3IAouTchOoTslF/u
Rb1Wsjpl3XRjkIvrctQRGkXAoctL0D30zJTy8C56I9J/ZeFN8hP6WyA5Bda8+vEOsMNSipwbdlYU
0gRBKpXi0kUWtVYpOvPSy/4SJgqurq0VAbAjT7feCQaM6Esh/EoDBrI0LXjFc60nIzjMhr4kP8gT
SomXSpL0q8qEmAWiuQyYRxtduaJCpPrNMV/bGbIkJe6NhnDE1LLARWmfJoZJglrxoqk7AMoiV1Tq
1pjRmOgOcS8NNiquRQcN5x83p5x8PTXCcDjYSZuzs/oS7Da9lDHRRlon+Io1M6xyMfwkUCA0xacH
Abzi2Uyx5mDkCXgAVq2y03zVgWaG8ymb1gh+iE+h00lFE6xbgUFUUuINxmpsYCfqJXCydsFl2k9e
mDWZ7BgBvDCcxTgEOWsvvMkSlReNU6rs6uF9zKZyRLW5MUsn6BgXerlga2FY2vTAO+SASIZPZdTv
Plq2Y9GWIug6jcQcBIjZ/ibGM42PqFIv63Y2eK3jxQSjZPnQbtb8JHV9GduGwr2Y/3iuo4Z1nLkG
0wPZyvc4flkv5QZKm5QiOCuzrV4c5Id2Jo3adT9ZBQD+q013tnz/u3bOQBRNNeGkqG+oBK9aO93d
kU0/iqr4jxj8iUAySqvvIrlcPb4mqkxiEkJVIUf6+BcwBRdCuFrPRofc9OF3jLNceqlRCxw/Uj4E
sV2VVrgb2pZybWzlRcvNvSERB/l90FLrlmOq8I63ZtZbQnociU4RZMhH5Oh++IcipV/Fx/vhQQsR
tYYtXbKvtEye3ZsVpZm+SpNBuU5uJ4GWltK3TA+xycBjFgEga4t7zRpwU9LuNkB6kI2LZc/9yHaR
kilvRxaqk4Xu2fmP/B6A8zH5teWKZLfZDcEXoZPNtFL+xhUJ4T+AaBPJ/EOFp7QNg2YmxghYSyv1
yXWukIK6fLEmr6Q15+lOx5mtC2mtZXDzamj6K7mgLJmhuQV11A6eBBgEUYrlJTSJLwxkHHwLaahA
bnYBdOSawV3tR0xi0HxveqdcpAgnG2wHe7rzS34ZmADJ5bI9Pf1aZW+xnLm9oN2d4Ai5022UxFO7
or2S2Ms3Wtv1Hgq0ssm9ZeP9UCRiMq1PNcJMoOT6MXtfp+br7kAI3knZrFdxgFKG7vIf/jeRqqod
5zPeC9QHLPFLt4r074S9OHnu5F5oiAn93MlI8hg/p0AHz0oUpDiCyIk+uhVmuHO5Cc0Gpvrt01mm
QDtfEF/0ET4uWCfeKfbESbS4wIGtdpUIJCK+aMKhTcYI3+xC+EkBpUrc8B2vQCg3wgmiHUr2N+Es
rAblfiI4yV1ZdzXK3W9xOSBOsuFjUbeJxtUPHx5c5AZGhGNtkVgxVZS2OQ0hAIpU28MUpsr/vpYh
CVUQ75pZtu1kFv3mnTeu9Yqq49ou940b55jOYUmfm2+yZ6Weu2m8rDRAyHSjxHLo1llsK6H21lVW
/Rn9HlTv5ZAeyGrLBIKsn5Rg0eHvICljM0wtORfDEqvVY7UF05a0yupMTjn8LE8rGfJS9+FUTnaX
iAFMmxuGdcpwQyw0L90pbGXrQ2Mi8fLJnCIcTG92VElec0lXjYkLyFELRUuGgm3SmJEIGDnqHeiD
FFBLSjjHwka5H5Na/bIKZs323OwHWe2i4+VFixJFo9eNKnJw/qm4svuKOJif+e++qwhAedLWiDhW
SapAC0a7kBAepMQJK7Tz8Mqy3oZCaP/3BdxwFEgndBYaUfV2mR9fBOzt6ho8dqLCjLrAU6l+nCp3
KOLE0mtS+SVRrd5EPgSrH7MkUrTAeChpoxIw5pQ1UC5WDHe8FQmM6cjdb4ZQZfNOrAqyY3FPAY4t
FAAlinzq26DdzuvQr3repWtxZ14ZBingIswQ+psX+8DomuA9RTKA5iyF0X4NiS6HeLgAsaJ8+K33
wXtvLKDtJCqTevzg3za817eYoll5vLpqJvQWmxr7V2q6Z4bx+S23p1/k0bzlBJOuaWhidKVPzy+Y
VMIJSFjwBMlOubTA/WojB6VkhC/D4zYJ+fPsrN477RfKzMeePc5Ew5kMF/PMzK4VQw0ycxgxgEde
j+T+5I+45GAislzLjGnOcIDk4ueviCs9vhZhpIxiXAetLbanFswmsKn7gXAEJZKCDmEhTNISbEYZ
V0VfTnRDdEkLuKrWOh3oUW7LkPm7xx6tU/EdM7eNu2ymwfVk8lxrbONvUuPgJs7V2Ad1HJUtgMu4
RRi8p4yBfR4M8E2bOLn3XZNOcc2sKSW8cdT7/uj41q6RrJspV755EUKDFld9yh/pN07s8KsafMkI
tKkO5BltPIvut3EokI6ic16htFzTM2e4P/MOUR3Ao0w9v2R05Mm8/LPd8YY8scpymiq0wzRjcPus
xGAZotAjXLNzVMNcemlJXUx03GrxDEo0KAsSjFiNLM2+fzxcqtRq25z1L7MKdCNEGJ1lVDRrQbSf
ZtOU0whbD4MNsGNidoeA7vgDmDy1y3GBcZFl9RA3D3uPl6B4Nlcr3tzXd4wABnecpC1G8D2nvho6
jPSvyAQTdjX/fhIgfZVfuAMcXuiZBFskUP74eyOYEd1qFZabGnaVLS5+jcoaTiiyVuJ1zecLNrrR
/2IlfBrE0sklPGpdM0LVq/lUKKOkjICEVWDVhehmVcXhwFSOhY3P5sS9NRUNMPRzMOIUCtOKyHsa
eVVSs1ZIJ+tQVvC8oFhdE7NcMFsFHsX6Dlr4MGxQbmY/nzkCJnufx/9oScUf8wXSJ4cxY7dvSn6u
dMyAj7nzCQXF8PD35e5OeRsQ9u/7LYsVQQJGQXJ6wxpB+Ux9toILLHNXQrYESyBDzz+Lw+wdu6XD
JmKfpTNCxHEEVZstoRotleb0u6ALXfxVzKD3DRVzlcSsmlEmukYYiiUXsrcVwIdoaPGo3B0Xn03Z
vOeO0u6owI1GEQmoGkSXtSjvoOQo4q6xbKs6I8Uq8ypbXd/gI8RJc2qaAwhQ8G8/TQILHH1R6wcb
BxK/R2ILnpgayVEwGO3WdAXpkY6xgWW0AvJf44hwLSVZR80fX55bQXXiC5ZQPCoXpcSH1/yokJmC
5zarOM5zUDxlBnt18GEmtLboiWr0igMP9kvWYUvsf382z7szzohZJYD6rb72BEhySQXDs99RAptC
4PsdF3LbsvtPtDLqILH207kCjev0qEtOSR8dUljYLy2u4I2NUMeM5DntQ7Qf96fvF82il0vwq1Fw
u48kgwpCPIRPmLwAkK4TXHwk57+g0meE+v9wBXsmtPJuclbMCmQWr0ak6s1CC2Uiia/s1Loyu4f0
uD0QqzEn6TI/aRiwn/ROVThwjeZ31e5nkBMPzZkgtMWNVTlkZHuyjUBrB4KErUAM5I6C7BQt62YJ
6JbdS5eim9b7ilW6n8m0U1XsQ4uqNQNcCk2PtwS9UT52/5QiS0/b8XgDMQIqWS3AjSFa/SQQnLCe
8qIs7hGWgEQc21XDUWuenxBA3C/PMda+ZbJSPvxiEB/PAqrjlC25ouSjDuprlHl2VZYWN8VEv00a
RxFqGwJu/QXWsEWNxWsdlB6vpkOu3qMBXc9KVHEsFv+buomurUhfG4fMUlFQHswV9F2CQHfRqi4M
0jE3hog3prFCvRMSlSh7nqaNBYaLW16dFvQRAQo97fCvJm2RLLw9ufIZ9kcUOCvK6xl0x5Tv/LEG
ShXM8OKcOob+n8hsq8iKdM4qlaivC6d9zFeKAAoADJdXAwwjhWnOim6AY3VWLkz04j1mh3hfERul
wCNQZ6qKwyUuGDzJv7rkaia+yJFJFMm9N/n1Hm2b3S4MH1PCudf62zoyrjVshZwgswvynH3loNFB
UKw+zKMX+KBJf/TCkQbreaxYfmqpQPObooSHCFhDhhE5mjnGFqZA90ywKyLeRLn2wJW3ZB58Y2Ss
7uMMGRSJHkO+UinS7iNQCuzwi6tgM+NZMiqccS27Ld8EBS8mhDrHABUFANtld6CwAR3FVtTOENvX
19x6FYqPtxHAjOxbVn4WUXN/FyU3x7ErHNi1gL3Vlb8EBQkL962K+Zt1L7pIK+wBrH6bO4yIZ+13
tM9QTfLtWNZJKMxyuc1imNOuci/Kn5M9bSFreS6fZggt9Fpt6WHapNkHwpY49iOUA1RbsxPQytOZ
Qf+Ivq6yC866k1rbWVwRRoBmU0IOrvio6KA4CRIysHoZI0vHqOy65tqenf1Xboe6SHvXGKCasEz5
qRA6ttzzc+5YzP3UgvV7rs2G7d8qI/8MtnDfHbcG6DmLHGj8wnJFYv0J5choukEzsLRm1/NWPGb+
FtU1mXnQ2cWbrxqboBFyogQ/ZCwIRduFjkZFzxXr7mrFnpuID2EW6uUEE/cwb0bjNewcJRBOFAv9
XAhROGpCRyiXsc4xwldl92Oj1zE48O7w4bY/zW+0lhjaM1/5XP8dsANBugUNV0ykhblsOceEz0/M
y4jbtLbRSzHlMfMtjLSwiu6J8Cwo9hKy/gMvy/ADGTqnpuwoooNSHqK14YQiLmq6tBUzxfk/xZFu
G8Es1mbFTYchYcCCXoLqUU0jhzGcQ2GXFrQNPw0oS8VDKj0KHVQf79vtYBQ5oQKOimHBIxbPlsy5
Z2saNVnC4Yg/ZMlpVMLC2D2Uso/dEI8buv6JNhc/MC1woJ9sFteASeA1GWGxA4Y4yxuRWeJuUJNk
d8YsvZF5YiYduiD/12wUP0eILUPEU6Ncp4hvJfmXn/f/0tFxzF2F41CQYxm17DGRG1s4xTv/+8ml
aDgLkLDK6pNuyY34dEglj9h+Z4Q9B3GVCKQPFAenoQBCexG2nl6Az51qq7yvObWOPE6KO/JiqLDS
vhjj9VKrL0qHCyPgshGsN3NkTV4qKd1hvFeuhsWZFILanLiC1IrOvt459h90qu+PYmamYzE1qh+n
9D55MX7J+vkmsZjteLGWYt2zN3IbGNkh1p1By2Scl/uCMRPoRUH1GuRuTvEFCjtIRTJu6gc7KZ+z
/aLrN+3mqoLT6t2tjY3IOjT4LgYV6rsWbsLcg3Y4K/rr+Bp99LFBkeRYh0295oJ85qlyA0O7pb0P
XGH8B1hbMXk3YCig3jdOcvuQe4Y5F3jrNwzoIyM8md3MrtpJyl8w3D42KkVsLFaRXzqdd9q31qlg
Uoj9Jjit/ZFvQpbeIt16Vc4w7V1uBnFLyJXBDbtom+36LVmaZCwY6Md8DtWCZDnTRF+iEHxAJHHB
xvV9hjCR6SDYU1qzBcr7xLOtKmpBdqgsv1he8boCi6kTDOyfH+KlnpTPw2d/FSzdVmaOpHC9zMgk
heXKlpjY1g5jalO4o4Y0WwR6VOvzQww2EcH3ULeb6p6e6Zork2J64taADTwKCxJ9Ksnh16nusgCz
eBp+wgSVXQEz/0mkHm0MRlPI+nMFYHo6LrpQ+4wbyGihv6KLfgBxPhce81Zy/0pQitv/m66oje36
7f7sfwVk3CmOfvOAogrjLWs76aMnG3lwesORH3sdzp3gTZknMEhLRjH1tmFVQHTavkH/w6smrFF4
R8IEz/52BI11f78zFsZT2qJ7+pLOJh3WDjC2ddq/MxbXLSrAHXXMtGVB2ggKQjOlzUTm5d6TRsEh
z30wT4Ks+HgtJT8W5b1X1X8cmiRP0lGCGvqzzs6/EpDgOFjkULvdXuT7XXEpICJs1PgyBzk/g9rp
1utWN5B43/3KZp5kNsP60Zj9Oqa8XCFEwA9eM/07xdQPdwi1rzfDql8oLclarowiBLBQoSivAu3W
Y6PzuSl8Z8BILTmUOInTMYnplTYLK/CJPav4QVE7fEJZ6xoDhnwzFSUyU8tVoJhxl366HNkEuMvJ
V2oMnJLAAF/LwhYsFt8ei1uI+1d36flpyz5fR59XaB2cdqhhe3yGHWpJ1KkuEFItDHXVCQWegzm9
UJYIxUqkcpo4Q/eYqWa6878kd+74i/MMbRrzOPJHk5Yigl/z2uxa7tCigWi8q98kKAxRxnB+ayRK
0eVU3BP1hpYZ5csHRExh1hCPBJtKkwNIBXXo9GXpMEZdkbF57JDY/0iZyXMUGpWKp7bb0fGFqSjn
GanJDWlqywEPl2Bje8K4xfuXGCjRfg1RIBg7/k4NlyHkq61QbD5vFtcoIjeNrzU21cjJSM0l7jrB
B7IZbo2MJY7oyeyd0VwCmsoePdFUzRAvRGOJQdHt2Y/YmbIifOQM76ppFSc/pf61tis5DwWJ2qR+
QaSMpxoHOhow0r3ksfL5eP8dzHedkA7WOKkTniIqcuJ6G6/6Vrht3ENxW7iIah0PqskQH7fvQaIr
2/mfCkOx9AbqOBFR5tSZ2PAZIbQViP6Pv/4U4PA6pZjhQ4yqAMZ7YQ7osV7wcggZF47/gWL2MFgc
vBSFq5+5kd8rw8ho8bOBH2bjIYcrgDDq9MaZ2+Q57l6MNjRMw8fk4hSGk5r8Wy5mniuJsOx/tZwP
trqBpZgs8xS1WFXR86h964TVMnVTdY6LkhXXhko0qNkAvRftb6PTrHs/auJWm9rEys0uxa5QC83+
0SfjGsxtWgaFI5QCccmlfvcTV9eulL44GyVzGU1PMb0opWSZDZj/fmpa4twENRpCnCQRRkr3dyzb
Ad5IXUI2pAv5SQOz4XD7P/ngdS19vQiqK92lNq/8ivkPJC1EiIebVR0FNN4jNyW1KDMvGKWWiGj4
937c5WSUJAri9dKJR289gZCWMmy5tetxSdZLiMsN9b4gcJ6djcQ/gJTjKTQFhbIWd2qjvyYJJPav
noi5+ad079WQ5fX2pLHxYLXYdY9lMcXtOobAx6WSgUCu3hNU4Lj4XojLIC4diuOxQU+3HBdALKIZ
RPLtXRrJE+J/GPeCST4mvRD44MhUXtEOOs7moCpoKqG+w3aTSIj3AW2iCSlYR7k/ngFDBMmAiGZG
mjlzPWVaK4odeh95fx8+F6BSdpJa1oGpu+heOZ0zseiT2727zTUUKBPOEWrk7apKQcMXjWde8FyT
EoIh9bW1+6xaZqDHo9sbmFVxZ0QrxKjkuYt7gbrKNp/MYvEe85WjQSP3V7O/Oh+LCZ+E57XD+r/j
1pFH5eyfq7FFDArexEbOyr25YUAesox2TZBdspfh1RGlH6ZJRkwpwNQHPyQE6fLjt1mHqJCrtTpI
trIZd7ZtHJdMGJZUPJe6N8hJC7ix8X5lEUBAxoormdJ0/iSahSppGHwfykDIdhwD7pd8g/JVLN1K
AkIWWaqgDJ7nwTxnRq9LFsLnwals4H1FBg7+qICw/xnfVMTlFvPxaB4cSod3Nc0IjiV7GpH02JjA
vN1ioSuPdU0IGDBt0GQmT5DJOLZ5KTLcLRvt/WYvqBJHK87AuUtcNPLtWW7Xh6It1hMU+wdBE5l8
4UcNheBhvFktqw5iXVN4l0cI/CtHhx3iIP0ilDfWDk5zMM9nscr81x8vbl50BE3A/660QegWl1XG
1WEsauqAcYdmLssDdgtwiSeLIhCwovGsaqhbAwD05FzcIvKmoBRNbEE+w5tIvb5dFY2SXNxXuh0g
/+aDct+KjV8ziwxUZvKo6tXFx3zHuo2uyEjcTMz7R3ICMbB0E1BugmkGbSuaVDMkBMFEvHF32a+I
7Bsel1QvfL5yP6dVDmAcegc8xIUuEdRIhmhyTVJKuWVMW72Bhua0CThcLYgmpcwdDqm9Rz9MOpLv
jy20h8rGI1R/hEfNlD6MAHZNo1w0kI6FLIR/Gmtt7rOd0tbe3ee1NvOCYM+vjZbsxeK9bMTen9D9
5oe81B9z5aA+w7/+N09yPgLy9+JdociyUld8gS3g2XN3k6PIWc8FlEsJHaaaiSfWl2BcwfVvR3o7
3T4o7rOul1WKQu9BubhUpQHbmkNLmLXRLsdeoyAzp9EuMct/y5WtwbdtRStYe+IuM+86htgL3qdt
GAcnJysJtVAALQHs0WKUVAn3RJMf1hVstqw9bNKdXghow4OYGYEgQ+wjw3T+xHJUuux+SzOUy269
8kXKLrGLSW3v/lYfI5uhuaB8OVBANU02vg6G2/+b2QZYwTYPcJwGxSQZPAyosrcyviZ5oSF4wWPn
i0m0/kBV7Nrytng5zCgWzjb80Ai8WM1oqK1qNii10cnuZLJZlgfQ0mAQ9bzGfVFtQFnyYnwRvRSW
tRe1MXpqKHA4+7utYhmJ3SJq+ZePboTEI5cJVJkR6sAyUxq/BnkAPesoGF7+3Oej4bm98dtGPSsb
YSI+VfCQNiblX5mtGTklKzohfAsr6YBydkt5Zdq5GFVsFMgtxBKCQxkUbMzdrBmxq8lUi53INWJf
/3+qGkoxNSXD30Bmsg5HMPbYvL8t8KH8663txK9S1fLTV49Od33HzS/ekBf0L17zpxX06DMtQhQw
vP/jn2/beCAWvQ/xZi03HSVuHNEE1E4oKmeJper802zJNbm9WzakmZ9xyjttIw/uq/m6ed6QQhYi
XjXEP2/51m6PMGe1WzVhKT9BDiU6j8OsVkRtr/cWQRr7DR5o68s14eV2xKU/oUK1kkhU0cNr/dBe
OJYDUB2ucpyl92jZ6LYPx48FIuPMfPT2nZfOySMqxZPjHBy83rC5NofDb0G7y3x/RGuJMJeDHAvP
j5kqtmoMh+fHrn/eMo0Ss55dKISfAWV9TtC4aeqinXiS4BGtxoF6LdiBKdLmh/R/9lqL/9XGzPjE
NvGViAtHs7BJFa14hNp/tA6W9IEq76g3DuHbHRU617j0Qk8pl1nF6cBqQuXXFRfTNQ0Ygb+WXGgl
fUongXFksnoekAeFOh5VXoziWmAPrEFHCIYCWcb4fAAFnG8YfEOYyiff4IT8oY+6oSeV4TbLAOLp
8qCi1I6gNpS+8hmeZJidJEg1Ch/tFFXI+pyynkzTxqIWKqilXnWJ9VjmRB0sqogb8x86KQQ0mri7
aEm4WhOuQWeg1WnbviIT9xkDSwNSshxPjPcQF6SKmSQvNCtU0z/5XLeCVDLbUTSGqob58gkGMRwh
BE/RIkvtWlTifY5I3b1oJAj7feWUHUR2cS2AgQgGco64PJFsSJEwQczfDVvXJaXgqeWd5CObRhVL
twTeUl8ytxLoUao7EzTGBX7Ag0ySqkMaSy5u3tmV9yCL6XR6jr0GEgXRi/B8sdFPEGBK95lwktW7
/OWbR0uTado4anI/UX2BAal4W6jeaXB6SOGhPsDsK7qv9dL5c36qwYokWAc9+6VFASy1q14mtW9C
iWNYPIAHQzkXi3TwGVjCnkvhpaRgZUbM2yIirTTQt7ABcR503MdteJtPKpB05R9hbfsA3XenAgvo
MlQhpY6Fdkkv8tBt89K9N2n2B+rbcM8X9VZR9/z7AF2eG/KFi29t9qKVKCGzcq0LIapjwObn8eA2
EkAklr2mOipudJjt/tWF7CoKjyFNTJ+FFrrH/lNq578NuZeCdYJQhgL6l/TvY6F2/0bYtCya5Jx9
uYWnRLA0eR5IA/feHg8rdGJJPXwBD0qpwNikeBp4+yB19jCvch6L5dF+4rAbvn28BP0ODe2ojfSc
womfrOpnGmiAjw79ITgTG/1ZXbuABRWQSYNa2Jo4uKKNMmLGIxBDJfWro7Dl6zADqHmWxhusTyfv
FHw6ycwxnccMuSjgtTJQ5SIgSHlLBlszX3FajkaANDuC/dAP7jkewxV8sko5fQ+c02orqGkUyMae
J+wnwkZ4BWsFTDwIJB6ET+dASTXr3LXoyt7Ne+RnbGnGARMe7rZZvgIxghGzR3H1jERJPamqc4bf
kQ9YhJYQuDVYTfbe5udZXFQTQ7SKGuvysSTr1TmO4t8HI2vsIDt/Vnj14X66JQC/s76CtX4xRQQs
Qs18kvcCvbhzZd+Ohy4NQjrOwhQWEtM4WjNtGdKTIKvEIU3ZssZhZ1uqkwCBXbNjY3QOj9hCvR6V
Ya74k037ImD9dfw1CgdbzwvcNhWjJ39hZLEX6xOxavYHLYZUFx37h9XhI2XYcIX3K7EhIFx+0/mr
aeXipWd03A0lVkZomjhau7FK9oBVgQ5bRZngVd5dND3VoJMWCRlOjoJCYA4NopCGF7+yGtbg8PqV
5Dfeg+YFS+k74Tgwzcq1+q69FgGqIZjnAUJH2vWRisTEMC/n88VGU8ItQ7C3n7kGUuz0MwB5iFu6
f3w46Q9cTRl0nNn9XmdDMzoLWhM3WR95aKtwhgF9xjxybCfZ8QMH4ZXurHTfDlXENNHM16uSHeJW
wocffgOX0MK9G1yCo+FFlGZIgijPueUE/a/9nUxGNFbKJJpCcCE/IJ9QUzfJN2pMB493gENAtAXm
1jm0SDRjLGb41J+XeAmfJbouDMZ3oscQerXWEwLfrC3E9gWjmE9RDfyykWxWF0Br1sC9DrfBQ5zp
zOsUKs0a/C9hyvh+CtkNYZv3xxks9XP5X3fcBduOFcpUdAg1j4IIN+fFaBBEoMxTbgatZTA6Pk0T
jJqjty1svul/Kqfj6BDk7Iomrf+l4Y3Erq49lMRh7Y4D7DkKZPyTK6/dJNCMDs18kDs8iKncwyd/
JuqeDo4MMh1WmI8/qVPSY/fRrBqJwQJLwo9QradZWiMzishmu1xL4LhXSzF6xZz0K+v3W3k4zPvg
Z5ceYgLif/dqA702t83Qyig0Xu9ei1a36ca4Bx1DQ26B7GU+bnBDnK9BTN+tp52/lr0m3/hTppiI
rTjXJ04I6hwPcV1v6Mq073wFF9+y+QyQRd9ea+QvP6+mSU6vt295t/5QLDKPx5M9Jnr+5uQsIUE0
yTs40xPNj9VyS331Cgjqyv5kuZ8oSMXNA1bxn8egm09NSKFWhUsIUKgfDqW8AKvVjwir09oiblEJ
SJll+EUGLaddoWSg0o510y6Qr6DqcQc837UwgmoA7POsuGgWpXNVFT7lZPk3aaWLScSOWPsfFXpf
WSEc1YFdeJBOBTrBplCvAolCATs3ZRMSroZN2V9ZGiRkIdfNvWr2Vh+SZuOio8ZJvnOdOywYnHkW
Ht0DjrjTiFDLvj5zmIk2vCnazvVNgYBql79u27bPHh0/4h2eMkQkgl/KD32NQNPcdQwU2Nkd+XTD
vTO58Ho4OsVpiX7PjUuA2ywV1LrNL51zeEJrSSRq9MdWPsa7Xjn5PzlpJDCBlRyfj6m96T/+U7K1
65qx18Avm5fGsQjzkqlSR/dUnKAfZYulZ0YxEBhef/yxAIkQzeU4KyJlGdpVMHhZN2XbN9kehR6M
pcMl97DAkGqWRhjAecsx0JsK+GDbHs9J/kf65yAVduEf/FZNyOuTmlC0rx60hVpNJLGfw22HArA/
NCIj8GM6XBQ64wHorreKZDwuDAXE860gDYA4F8wxbTIeFjprVOyPUqnHSwZNEliFg0DAPvePjFbZ
SpTENtNyYwLmMHTswosoEmB/konyNIJ/5v4AFfqVMIFSgvvDTZ3/DeVn4CtDhcmiYcPI2GkjzZY+
IuLncBckOtfVWqN8PYexanFl1dd+sC5U/PZpCm4epA1LH4ZjMN85cfB8eR2YM/CPIaVYwQfPvqtC
q7LhTFiw7anRTGdFYQ6BBSBKtRq7tiClX/V6iOVcgRNRkzmY3T/UlBM0JZ1GqInoEt31bH0ZH5ho
D4RvJXWHxWFXpBRVTK9LluJXmwRvacn19XJsTG3hLhtN6a5xE9npejj+Sgxy3ZdIQ/BaTJPyAmZz
qjBwnB/gY43iBt3fEUPTxz7btGVmpLr0I8NlS1nL6w8HSE9eg7ulaK73YprR+v6bv5CDJWOQHUN4
jk0BD5Kd4FWDsXtE8GSe+A7MrcBSz42xwJ71Y/TtxUUBFPOPrs7mU5mYPWE4klxP25BaL6tPOqCt
PbqMNZKMre8SZh4B2dm2RQcaUTOjHlUvDNbwQ4lDH498ybiND8k148FI+JMMLh1wcQ1JmmzeynRA
LZeTrtP7Gdef4BOUAXPlUraiBbpJ3y4CAiYvJqTVnXWVLxB65mKfkyX/S+Rw/AIiR8ratB2TGu+M
Ducz62X5/3z2H/rQcAdOi2E6J1FstmdgeUJCaOaJ7MdbjFNSsnYVCRpcgfYvrW8MLkj/c8sP0gBh
rSIAjR6szlpd+IrS+63IAC0vSHZs7uGRS1KlSFtxBvqakST81Pl9LMUkfTdsPLWPmCyJiCnN2BU6
qC+OQCfQlYkM7M09M2HTbsJF8PWsZYXVelbp1yWtxJ75QUeBdYeiSOeFNSt4szuPdDwns9A/pnmA
268G7pAsTn0FScy0kqELB/sJkwh4hV2zLZExIT4eXDb0EPaD8xFcP/MsYYrRzwB4zVqy4TfXtP6w
0I8IU/nC3p0ksHU5BxWFvcgRQCfPyDDuaqlTAZCJdcQdifTM3spgYA54nop1/01/wJ/yYX4Vw0m/
weheLkjxgNKqcELTfAjJTqYN6YwNjB0d5pHLwptLVne3+u8EbkYkcOiWDccsWJodgJ2HaQLuzjut
O38ivGQr4iz5+Y9buLPUib5lanDIdlcThNXAgwUNwVFGOJg1kf6bJ5w2GG9lQ5MwT7fMcgbQCzmM
3wmdd/QVH+PW1OSUwUKnKqQOL0IGVF96oLxzojEgIPin1ai/DrNSIeyTLCzylip9a+g/fbcww+6k
VKrCbs+Ioi77wvtey+TjFGDOwLMmQ/b7lVgPrxcZCErnC5TIMxgLk7lNfclUIGQlPDDuFKcEaiDf
+ROQhkp1AlndNIRAbWXI907VWY/kXRV97wf1cfRmiV3sFmIJVfAigiib54jStID54iTLcAuSk31j
1JI63InaUaJvrJKn4BwD1xCXf+kt2aRc06FKSBFj7h8G10Z5RcycZC1jjt3AeoFcWic/8XgIF/us
tXecwGj9Y/3SlHKcJbseUTQI22VQpDCGAIsI3by7yfIiw5IAH/AnQVccm5W02WHstyu8SrWhOVN9
RDm3b7eSxYV7bOlVCyDiIYhwFQUesV/NTnJ+jVHZfD00rfEC52XhBGOtsoDTPvEgdfOkWDZ+hBao
dmrE/HUkjaDmjF4bE2fD0vwp4+4suuHksIqG1GNAVqya6yWAiAQGsNlHOAFwzh/pSlIK82trT1is
XE5TjQAmgqQN2mlzdvBf70+HJZs53WEaPPPh7wvlnNMx4QIMhNQvDHn5FHZpC6RIcT6AmBEZLiMj
dGoXNoC8xBPa9S+ebwVwpMY7OkE6lqrqPSlGwFH7jeb+gaUI3zJqsSHAmAu0n4Pi7yUF630zKsQd
+tctPd9lysPHGepNmqJnaexNqf39yhYJColZBLEddg7cCmuJ8yiv+8uqnUI4pNHAlucwqqXOpNy6
WHhQ3h32ixYDOzaw7gxKm25OVD0YJnANerC712h6l+nu3io9fHJsAmnFVH161hXny2jj7npVwqRR
5Ephqufh8CDnQzC2/OZfaSRC/wy2D9B2lCEfi/PP52GPQriQYK7INYSSOO1/JiuClROySPQO2i6K
tncH87ep7b3w8Nbfoq/KGOWhx9RwMvHbsS3P70k7Qe+y2TrVhb64AYTjWJqvRuviVOJvcnMbGuzm
0wl2WTymg2pPNMTw3o0mv8Q+/7lQ1QeA9AOJKtEDYLxcqCGKCBIRh3EwPQVLrngxmRmsmsuGK6z+
hd95cNyRZ7+9EOZqUq9QonOFb0DQoPzFJRu5uMPdpEO2JHRkSGNTNzjJXaHcFxkrCsdXQf4knPD2
+QCfea0PHmlcv4R4HTgn+KK5WFjV8X+EIP0SDtmeMxUrhXNMDTNMcylNliUYvIynTEJD58olGLvt
LuQgiPuW27RFq0odTpUGTUz7fv0WqaDFjs/yT3uwuUn5b+EKsHZNlVwkll3no4iL9O0JTacc3Yuu
XDcxVGe/WgQaqH7RZvYFudd9x6fMG1KCnp4clk+rkMBLMxeeqTPJcV8k7Sns5nFs8rh0mdWlVPPN
kyOECCJiQRbQL9QYPCK0xia99CbY9G9RH6ivr85oDQ4Xtrj3FlPDUj+/6moNtdVLfuCtGGCdd9/Y
SDGi8Au1IHFV2sz8sLV/DOjSGJYK1nMU1BDTG9B9y8V5MqaSP7Y2a0Ih43sixmAFY81KGEFL3qQr
Sddf+W9eqq5JzOSip5j95gLHvzmJYMY4hbrkv+QHxr42rsGK/UFcotcSYua8IYK7SfFLIjJdgmCa
WJrj8RvwOfvKv6w0N6mOrmk5frrFVXi/pWrBrRI+BPWUCNiWdOgo+PBdy/pylAeaLclb4bAWJjTo
y/h230cCJDhIGREKTrjzBwd0wjusF12V6DidXdQ+fCgU+cTqNEGIjo8PyH96BGqEOHXwRcCNxbj+
gQkxm8JBoLNUcYdMVk+Mk3UMrNMcYR5sDKmsgOuL8DrC810uMbSuVBw0mjeeBV+UnB1AaOWa+g1p
k1P8dVa7nXtwhh0g3xelrOCHJ0lQyN67dWUgTEhb701i1mqb4bXpYaNMEOWBFUQd2qSxIEcANFUT
+h8tZRLs6csJ1TMioceoS8NQJgvf6PBpCFH8rmO0mGEbApmmxwhdMTQKIqHafkZFmj83+O5Fj8QT
tq2r+LoZRxAiv+uLPM+GkQ6klPWWVNz7QMlIsPdPuvrSqFKJgqBHNjceW7I9Ocnbtbnx01Lj3+1L
wSXMxuSWKbUydCZCTOOoQgBHDNQoldanV1Zx/q2sGkkUnk5nKKc52zxS+MV2k2b77MbnrGCtTj5A
mVXgvuBOTfeieU+WggA6Nn5/Ol8HAHSHFRUM6/ekWXvt9CbuWa0zRzLm/x3/31Gv++zkYQL95xTs
E11okwp2pmBoxrwgpEl7LTjnegriTP/Rof7w6UMvFvKXOZ4Z1q4YhaDxc7O/Q/0D+dc8zHC6QnJL
8pvn9gNv3SfmrwuQnU5R7heR2ykHjEFheJnO3Tf8QeCMSdPznMiOeN9dN2cu/CY1xySPNUKCc1sm
HJ6SuaBuOYaZQq36bIsEqGPG1o5pZi8rapzOqr1KZ4jSxvK+9m+Pv/zwficfUY8t24FDmVVrxLDZ
sTtCpSHnwVpy84t2GOSBK/VCBo/kEygS6tR7rb4W8rfzUrzHQgGiLR6Azj2Q0fZKU3AyME25RerH
d3cJhaT9G4HOP6THzkP2xu0b4rH9twLJrFQqVIIrTKkpbk9sWQwCurfgoYW6Z0D3BAPOzFHcNx4T
SC4xM6jND73WAEjzlKRlXZ3pXAilq22bJPCM+UwCf0KuhTA4/6Mp9OKxYu4JRu8IZhPbyXmx3yox
m2UMBXuO3HuzeQ4FAA3ovtaw1QmLAO3lPj+SCiC/BU1qKLAFiyhaO8kOPSg9FdetsXsYzqWSV3IE
Jv/u1DOcNaGQk4D9I/+Z9hdBagQNqw9kGFuTUllyYg5l1cugVSadYPCt1eKFHfr9BAkKM1nMI7WK
YBl8T0qOX6yBm/JFmW73CpgLu3n1WzVhqTqR9m9/PPNfWMNEoTZrbEhs6dlXfWv/WFppRosAkr94
F/kenYTxGJny7+GzoVZBdZ4fBqmoKtmfIsjUpOH2qxXbbhlhQdYU68z8vN/vd65/hjdzzQCitAWJ
Puhtej/XZq6qlZLh9gnzYoJJ+7JJjb5eZg1L14O5aclHMYYfiZcOheZMHZeQ4TPJQsvMmI8RdC+V
9+qruttQImVFNnPe7Ww26of7q93eIxsWLYlap5k/c5pCrvuAC40A8d3NocZkW6tAlwtVghbpZUgN
3xMnlGx/NdFb41wqt9TxJ3IMET6AfdrQUiFCE3WFwXQbEfA6nBXzp9/Y8wfInmMypacAV+o5yYFQ
OqcgKi1rVqebzPPMGjT2chll3Q47aCDo9hVwhTHiAmhklXz56ljGv747VtrBtLLKwaogmxNV5uAH
XShZ96Cd9PX0Y8tVC6GpqwvjAHYpBrP6utVCxcleYR4v/qKh6ImiYNsjZICMlypr4acNHqgq5GAW
YqkJv4Amg4cjm4YZf/Bjy1uxxGrRvia+TCfgtRuxX6WbG35CgG/P64cPpK7aLA7uXhyq0YTK9Jn8
pBGBMYNgtkwfpEtM4ViQhb2PceEca5YE0MxTGnt4T2QPV3I+htS48T+ZOz1TeiTXHXQE9D7YYdyL
GZVFb93xyiI/0yEjepGNByCHMFwIbXNWmfOD/Q9PNJGUDD2RIZDr2dnpfDdoOt18qazrwUL9FJUN
OSv4FbIjirw5wR8Yq02Pjz/SO5D+BVx4ndkXrCmhWAxFnuimVxy5MbasxDakukMxrnGnGjRuOOp3
6ONSNljvRsvyDPVoZD/wPgJ/qadcgWz4ydJhkGjuYlgtBNiru9/uV3V6ffqacaOq8fnxbravYOMF
P9MwpEFwfUwitGUahLw50G7ws3oQsSYPT6p+p5hOmQqW7JJ7+4WCM5Z02zlLhZtYhMcHs1ShslbE
bVQYgdPtHsJAC88GyvVWs3c9+/D0KRHZBMnVl7sXl6yYXQJHIfUkxNZl4miekYRIpSPAyhaTAagf
0xgyXjXKEVWUFxCEVF6KivpiLSs4/8pWCuiPq0g0RO64TI/JWfXTiJksgrMmD5bcK5Bn5gnQY7+/
mlLx9FiGupmVqDz2ZKuEv5ojTM+UGvzt8SlOuWOsbwF93q0Tc/eSxU2bZc74jrXOiIRjvcTDLcUU
uIvzeLyzPMcW1M5CSPDX3AHMwa9HsGEhZ/jr9TWtzusI43IlgGx6SDfIXLuLNjyugqfu2eKxMAMh
TpCunW4vT9A+ODlxqw39/OOORmFk8JExZtweMkK4lYZUSRqgTzHxzuLHgKTR34TYaJIuBZbxL3o5
Ma2ag2NZj6HXaCwOS0Ls0a75AXWkt6HflEyqIcdOMjS5DteSUvY1RHVHZ/Fa61b/E7qJa6gI9ey5
kpCtCTZ4oo4T26SgtMBH97Adw6Qe4JAqZHmzrBEtKcY+s7nVZ0zxIa82HYQ6hki1wQ3x2w0kzIXk
I07XtGS4MY7vaSNuB90Z2bimG3G9yADweJ54ICb7kZoJQql8ToTR/WWE33Oqzct4O9QoqGlJp5MR
pN8OXNKnPk3gmXz8l6Tq4AycDnM/WiNkVhgHltEB9WUpyr8T4J2lxPovva+XxcyuP5GGSxON/269
LFjVteVloEyVVgF1fZNMebu3LXJdB1anc7wtkvg5FBdPt3ul1XG6yj/Hj06pfuk+L7xqhwjdnsOV
NHLCzLt4xEbv8mLW6hOpdg4gEW/no0iPSYTQzozCF0kRuk594ADF7EIJpiXuQycF4pMz3kSYdP4O
s0hdNbG9pbZYefQxHZS+Q9CSWdOpoqD+tx8vX4zH1VwqYwkhk87t2f6RY+Q6EoUpKSzm0efHGoNM
OlWWdVfiz+T4XYHMhywxys4QuA4DcWkWDVgS3m7wbcGS662XEZUFYYZFIP1GFCg/U3lotaOTXddj
w83/uk4xEusyx0Kn0FtwT7Xj1piUvK6TA4E4TvmjWK7Sj0T5KfKrOpHzPfbBs5GUkwTsRmZCFd6U
1i5oXLSk+MAEXEeyiptmlWHgHHt4ittRILJpA0SDrASU4YJ3yZPmE2bHF9TCqpb6p3Oer7mh1Dqs
vAGekg6ElBVJc/QVEMGGfwUOapXIxknvguG1/fwimFDDMzoV6q5rZfgLRoh/hDYpRQK5rlNtN3/e
u/CnLysPhx9dkdmQPUfCZVQ/T9PWiNjpNsYCgL831wOvIAKfFdxT/IdtdI/0jt0lEOzZO1Tzv5d3
Wy1GnFYhojW8JwPMocDgEbO824NlrXl0Er0zkE1HIT/jcJPFy+U5xO6hhrpoEnwqYfvENWgmW9Y2
l+QeNH0f66aN6GdbbqGXueazdVr91R9psL+k6EUmipRlN/opnuQZrzLw0AAX773tkRuGfgBqsiTA
wKaqdKGa35vE1dAke7Omh85bjrPPMXQl6cGPZL8YVDZcvWgQb1QSv4EtqNMbFT0fSaoXyQUxqdlp
XBIC5860zRleXPbylOWqykAkZPvqcqsHHx1xh/dJ/gV+5szotpuC9m9ouzIpSF87Rrq6/fsaztYO
ts8jVmy9ceNpsq7otLOB5oXbbtOtHHqtRtjk4M1q9aTFV2P1vyMC9T4k7P8PrN9Wx3WCOx8QW4u+
u56L9uKFkPMG4wUeCmzVHOGuj19hG8nO3O1vibBI6CW+yNmzBN2dj31yYxjRi57ES5h447+7gSP3
RZutd8mSFDybUWW2e0WEbstX8TBsgKdAGFYemfTzik5yT0eE4dYzbIGipMqVA3haR00V2EMonJ1f
fDnJDod5NogU5TvhoqUfp6WLI+dhJiq7ENeR7bPLhNxTuvOYh26C0cMfl3TEXJLV6xxWlDLRmYZT
lc900ps0Rj2x77CmHgs67M7oLEECuCVfAFX8BeuxACymXFKE1n81nl3oCQcJ9cWxYBmOcyiVGhe1
+yKDImWcOkU0kVq7HPGowL9U+V6C31/lXdZkxkmp5CmKHJGVn4bgKoZ8CqDyMyx0kLB3w36ZCulO
myrYmWjSQ+2rV7SguutEY2lS+oT8hsGGao463CuJ2VlX/iY0u2lO+1ij+PFb+3qosgSCgoONm+2Z
F1N4Lahjt4hMPC57qWEr45aPpFwSoKwN0lVMGeRSpfmcdqCCRILGiA/IT+WDW0mVinEFyJWFXjyk
FtBTisRQg/e1Eg2kzgzeyZjSA4GOGrwwkxKskEw3SRpWnZ2bL5lgxwLin35FymtAWvwgUTNYkDIR
lmTopuwv3hbL/bN33dDg7PX8Lx3vRrIUedySsla5/gz7Jpry5unOAbwHFqM7zxkA0zrMSFsw8Gvu
ZSOeQHIfOx0lPMLk79LBBCnzteSNIIuVmWppeS4GgcACt9B2d9vkIAwvx/f5Di7PvbFQbJ6aeAvb
aDQyeZ05yCeVJcPrTWQTgZPBUbE+YHseF2ccK6FbsOdAIeWuVm5XZCEPwvbJ3qB0uXxyPuiPoyy4
dTS/QG/RZgPUQ9k48lqXxnLyjcpBMl1t8w6oVGoBL1PkirYRD2PY4/RHrH7rYKW5E0FKJZNGp6w0
+kOTg4BjpiO7N3218Xhfdg1OpHdZzfZ7JwhRAiODMDchBCSbL5+4JzlMe8kdYA6b+tiQvgIhL2lc
3Gzb1HB+q8j3oXA/4n6knBCNN4WO4Qv1/y2NfIGRUjqUTHhigh80f+dmy53at1mp4unemYGfdlLx
nnkB5jWc3X9rOu1aZQ4mII4eJ+S3o9834FU3dq39cMUxR0Q16dRzIbtBpgCBt5Cun+zv6Zg2CYrT
9vg5hNfWrS/hxWIvEAMHexVwNB8y+chmwDy4wdI3oiQXD/v9bm/BuR2bmrgoEqFrurpTq5uRsVxB
K2wpDKJHTn+2spcs56MCTEzVbV84Ck6n4vWuLhwaSjyAeH8qrLfM+PYi4N3sufzPxXQAneyMJdI6
VwOnhkt07Km8rwtQlA/9wKvXqEuKd2eJOTptkED/O4VWpiJTBQE7o0SEy0A0XAZ5nTlIU0BiydW9
94vwmOrzYKhMNO/vDbw7kUanU+6mBOI7Zf8i6Y6EIkpxHE3EdG24tNKgb0QEv4bHQigCR8rhdGb8
EYiRPADuCpNS9mLuT+mDxyjv4MeUPGVDc+/mVUScRPb7S+wvoIqiBoYR7PXqgQplFm2/pxXjLjHi
0gJCmTkCrp5oNcdO0Srwy8pOeC7elsYsbGJKFf6nbHoF4pRZPZaprLKP1QkYjSh+dVCstHZQx4rJ
xDPxy85ontuoEDb2BRPSkKgvQbWNxiYf8DoTgmRnzirrqlkisyJmWHxJLy+CCeg0G9YXdYoIh6f4
vUax1tw9saILmF+GOASwHVXSx5/hfMD7FFtetS0cTmrliic9ZaFQwbLTt0CSwqusGeGbsG3c+odd
tWC/MTi/P18f0NZw5yGOTIAQZOiPUlPNIYPgx4G9oiaI1+uy/gVZ6Xe7R55tQ2/1k+PdyotnmEr1
gBd0UiQyhPPs4pwTn2VySQ4w6938uo31Cs5Lt+ucnqDkttcZOadOe4fh41s6kRJvYVyLoBn+Ezas
4Dq6pipKDqQ2sWjO81rAcVi/b5oUMo/HQj/XcpexziFkYkxzwIaZ6V35ib79rrS5XxemnUmMZR1g
uhi38vrXOeCQHDpdmk1UK3wpaG4H80fowMLA4390PfqkSrITKkwNs01i5rOlFode1QQqj18TwXIw
pv6vGuQ4s3/fJ0/74x1SgYfMvNWc3xIjkTMq/5TpTusIEPLKcYOeGuNzkPyl9FvTRsDohHLlJTha
2Xg5auxYDQF4gsEldBVolUxtNBNwM31YJAov3Hh1R42fg0c3QIS5t6F5lL+dJF3GPbT2L+VieiE/
/7GtRchtNn3zJABLi0f0EAObQZyxSD7Wx7X5topaQUlqsZ2DK7LWGj+7u/cmdjgO/yMitHGrQXPk
rL8C1+lS/SS1ZocO7JvNo1saxNY9k0ddMX7a2FTinhhX4wMYtx1Rof//lr1iTFZnJqRboTDbNq+m
pCVS50gZfpW1eJTwcbDba9uRxTkhVF5SRN4O4z9TGBtWdm4bzLMA2mfQ7a3YVlHgy1fYvMDjVsmi
QT3+MGDT6FrUoH1NdxkJ0H0JZqyqcesInniO6wfMo3SFT7WQjvHRWO+RlEt1wlBhuRSTffihmeem
UXxPktkmluGXybxKR/QhbFZrXgjxNoMlAYWZIAUzU+5wa4ZjSQaLkpNgGwV5Zjv9sX61WM82Xglk
q/JQ+4l1avkaPeytIj5jJnYvXujcjt/r5BZavBGeknGeWcLAR0nof3lXWiaNtNSaIVSaQ8zsLnFt
c2Ff5otYFq4FAq8+TOtejDdFxMp2fnCFMn2Iq1xUeqpL12VsTsIweBW3kFRzuD5vImfqzFAk+jpp
OO6i0FcJ0tSsQY7pLJqpKoX1XrRNg0PbhBjMKk7Kz0CfiX0DqEvsV37wIsNsuPqMgBsxE448f+Uu
GQCeLcAPwMqWFi+AUBB7nJbRIgpNb6ZPnyrkmbzjB+6KpqFxzxpXAGO32faoH13i8+qizFR9AGEZ
ERZX2+tP4rQzizh4ydwABWDfmu+1W+e/YSatTaUbhwvQ30s4OGP9GbPis/0lDVAzPIxbEbRrt/Lm
sqgIsp6O990blbl6Jv3APQzkSc5BsgPvsLv0DPJnWNeCo0GD8JcfsacVeu3BTVHmmTy9nQNRIC8q
d/TUJ2i+oHUxyzNnZpyvT+GP5Kk+k/12DpAEvsPbx3nY7h8x4L8qDg4ASErtNxUIXqNA1Tk+5a+e
+uS/DrQgfVqos8WoT4GqtJDY3H7u4eYdPuS33ZAOR/STVWsqxkj7Nfn2q6XWEkn9jeHXBHumhg+i
VJeDV91JflsbS4VkjKSbAEvr5/EsLIucoZWzjivBQvIaQ3MNYim5I3E2s7EH76DINHMS3ZFR5G9v
D4KUSWJ+u2k5lzohnILjae1LKOBLmiMDQccyYtBwA7BRb3ey9AjDYCff/Jy5Bbub8eoHfvZPLA/S
9OiA2xoTP6uVfc55E2RP31Lo+Ky2vRV2c7VzkLXA0fRt9wUz++5BCjJWH+FjiSt0H7pD5mSaWdAD
joN7PEdajtET4tfc4wrltTGi4kt82rnc6sHh/LtM7UrhOujSIXaw45TqUWPbB5J87VqFKrdPXTdO
pEbxQ7LMA53y/gIYAWjf9+/SvTunzrcOcWLXNORaVGqRxZayl66UCFBeWgjew2Qgz/nJpIO1cz3o
ZRqpNiB/5sffzIWG6fOEZ+YPPONx45eBoR3giTEnRiS0AMmrD9tyxLXDilGXSaGn5MUlpX/65kWe
9FTsW/hGl0SZUGKXtXSBV1Fyp6SZKZFSo4STQqY2SaQPOGGmu8ewhmlulB5VCLEWTFSel3ah+V6U
qiaebXDeSXfpx0o1ZVi+D0ycUxcc0H7MBgrVqzXiaSxzMl6DvRRHEgOxapigbLX74PURHLiZ3JvS
fIWmYBuSyviZaQwku3wF0crbBExVfRCV/HKJFFEgMZQ0aqo07EgKQaB3hhSxp3lm6ySVXSPa2cBk
u6AalhkmLj0qa6DdT8tQZYROAPBDPpAGTU7WXKhhn7Iayp/fpd/C+lcqQ0aicqNPCFrXFomxeR0u
n5ooBWx23fxbPCjaskzc3FnPlNTG6QILKMYa/S21s9W7kFnlnXbye4bnL904/uxglDlrWvJjuGtp
sUs2W9eLZTVMyg3lKqAG+r44Xk4Kxp72/H2dxp5y0jJZ/eDqMCtycsKqzZBc136r+ePwg1iqC9va
DhRFO6o8ETBMozjp2/pRYt5C314XawIFZcl+DzmhZ/30BAFx8Wf3iMj6l60SlOKbfmMFhJYLSPL/
ydtOYchCRay1lTqVXeevKCiOVDLV79mc1OZPbArMnhSr0QyZ9gx27yhOThiX5fL1yA12+hCtmapI
f3Bjk/emwW+BiMW0t0SyUfd6wW6+K5unh7HbUXQfSpCLmilCg0HpscU5VOHoNMSdF+qzZ6AHf85N
vd23B6ttHbq2WI4KGttALjeiwecyvXkQ+Jh1Plk4Z1qyajdQE6b81zwrS9AFJoJcYdo5JEUCFHPR
X9uDf8HjaoChL5vwhVbIf0xyXgvJ6semp679m4QQhBpm/+bjyzEa9tGZlh68yq5XohJtiOnqsit1
K+kgFcyIof1Lav/J/F0k4/+vwgNUQERH8I9EprR2ryA4lQq3nnoORhQWRl7nxuBh/RQBCIo8Dvy9
/vray0Hn0kpIIHZ/xFwD0jx0tcPmZzJn62xpw6jxaBwtr0iKfmV9QsEEfdRzu6F3i0w6e2FZoQ+V
eWahz3NjOAiwuVsMSSboST7ZsvV2GnOi5JfVlUzVWexFbX466lg35j3dByWDn0Wfb0yEFK5adqNw
E8eRvJLveAPeSgqtBnuNX8Ed1LfomDQ+0xSGxovpSQ2AJz5YMyK37XvR6Xhd9H0KMaOdW/OMQt2R
T+F1AqX/6hXNl63zp+UYrfQqNTU2Dbzfn02YY5X8km8+sJN8s38wvGPnovjc8XkIU5R4cUUq0qDu
8bgAaW98ScwDParHZzv/h20HKqf9dYJApbbcs4t3+OwXVd+Kj1Cys623vikEmHJ0+IN0eNgRk0CK
3ezPxPsX/x1UBMjIOuLDoAEu6cKRnee5+vH+YLwRQEEyyMp2XyLAGyrC/haOpWrrOtBh4B8lzvYH
39qVd4St+qGMb9Bm19yGwl25hf8Z075Z4zAhxSzFSYNcImbZ/7hE3oV0KXwG08YFZFBd/UOktvzB
VeafisYawyJNYCMXnOAbHU4A23m+GDGqqNQE/Oa1ube9MOzAlNgYZiq1k7I4pRsNgT5BN8+2VhaM
RbSeWYvqvsiPZnjO8tpBqwoFW20BAZTo1H4Nt0jIf8ODyUzv0ZbZ1tB/2sWe4DE/W+e8SPSa1GAo
d+PqqWuea2QjmGO5T+wGipbJKeGH5zoh2bI8ulpfLgWALGhVHAacWqa0qEo02sUClTUr+e30G5D7
W9eBRRuNuTBxRuWJg2iNy5UtTj3RXCDZyawSg9mKX063yxOsqIzT+JGHzKsdKeaib9NCO3m7LCKO
QGDTkrFxmPahXl/Ww+0G9tZ9/yQYseykP5BNSS7J4+9g0hTRpDLfScnw+1UoGGTSPGQHN4FMv/wV
K7nn7kQlDjtEvXS774HRabpBXzWyKETEMTIoB1htfv+qx3SIv8OonQFnxu1qSIZiXifQxYyk9lnv
hv6dczNGNbxuvrIuVnG5vqsIBx68lkZqq+GaSGdrAD3/cKpjf+XAa5c7tSD94NY6B2tuheeZ+rIz
LbU14m+hzF4IPGxvp3WHrJUQIp9ywngEGZNMYiTN7JqR3uv3Bt256tOltr9N+LQxAEfDUUEtSwpq
ThYyQ2fKUe21Crog8eALBYMaLfxbK0b1O8apd6p/ie34hbqX9zrcHvqQA1yiXBH5Ehon3qMCBilU
h574sYoDIT/kcDR3YxWU0cUJgeJvU1SEHQZ+AOD0wQXYn7TwSHb9a+Cq6St29L4CvIK/GzawgBCE
swBnTxCQKQfJ0rwnkGLnLQSlE3zzVREDquuAU7ZUE2E6b1gsAmW1OGlQPidQ3cXMWkoEZuEmo0xk
dVxaKh+XoSKntcTI8CjmBaOA9AzjccywQwxp0sXEkiKCGNn8LF5ONZsqzUgyFCXa2vDC3iBafTha
LNb0prnyRUQTgj7da6uWRvBcBujF6udTF518/teKTY5eS4xADU3mgyISUw1bVF7IkqEbD+PXA3t/
UKblJhTJf+gVeGhQmeCSgQPndspXK0GFDeaavdsy+PpIuu1tkQ+w8KiLXIj1riZApY0ASllhoBDO
O/6ONB8XE4kvP3PQcTJ+uZ0XxM/d4vox8Avt4ojZERXc67EYCb7Ik7bRDiWaiObrRvC28aFrItnM
cqulyILrp7V6Hvyz6oXPh14idA0zhSbIxiQAJpagJj6pcQTPndJWVxJNBe/6CBr62HuhxPpc5/xM
diW65g8nurVNW99db6vdC+3r953kMNDZSUbYGVHtLYzQjqew80D3zIIEe0kSVgAUoOtwdscbhS8e
C7CVkqJwLSrQX7ANP7016zW8hAHkqol/uVlBsWonaW2Pb9xNDtNpT+yfL82Tq9Z5Pyo2eoT4I955
n42FX/NWQSa3bfMBXWmgW7ovuUDRPQQHj0IQi6l/du+JsR7TEsyKS9BuBE+NphLisoSySpcm1USl
xixrcue/AUHXf3Uye2wxiLo4i3ehvrNAfQpdFYdhXHd0uU/Yjhp9rEX8QFykoUsHcVknRTiz1Ptq
ivOguKmqXiIePMZL0mrM54bugkWcB4rsQ7JtBTUCDjsS9kB0Z4ZeJnbJ06HMNLe0xhfc1pN8ct+B
dhPythP0M0uxF8RwEFEP/yhYezZiKB46EQpg3ZJESj9yc0ZcMmKHYNM62Iu4Jx++Ismx0n+5OmwT
Ycjsq3P0gYh+JihUqg+4OcTW5zY0DH3eWjrVn4obq602jG4ohAG4omLcUlb+S72feevmqp2ffrHp
Tq6T/g1E1Dobs/OHbc03FQiQ8k3to+wC6INIqEHCNtWrBw7DPuEyOfcUCc9VwWHSV5e2pQ8vKFvm
W1U2Ryla0FWy5UxaxI5gkCU2uYqecL26OF1/iz7KckN3YHTBFiWYArFXNRPxOfqSZkImeEQn3p3/
l4i6GIeqDKROOEjkiCr/BnKnyExryNFseFEcbl+zFMTi24nou19v1CQ85LpOmpsgI97IOUQWbSnp
OCp4stmwCLpmxPxMvqt4/vtFDX1TnZsCT4NeSKqLU6kc3eFL/qW9zoGP8JNBnSe3s5971Z3YuS/N
g3I16CERMi373vTzhDH9PXxih3nLXTOPLNxCdjdI9lg2+MM0gUtBwwQZM0EGPc0EVH5kXHm5IYK/
g0t0+iu87ZxbEikzMhxbCRoVCspTOoX7fINU2HTW4Ra+IayLNenqFS1DQDjkkqIvDnIpse60QMyE
bIBBwoXr5qerl/NRWtQoX3RfdzoCcbFXNO1U4HkI5WAE8ii8h2L2auHF6sbG+Jx/yUpFcLFoeckw
ZIAqh61SsZPc+hzyiUepvXsGTGLFMtLXuYaDFTivBqmqi74lyJC9tH1o73ktHtst4Xk56vPAQJz9
05v6yAw1e0BSK5AX/vpbhnbYxTOHxvnAJQSkyu9TLIHSK7tSY6ZJrGJVbLUOnyyfG64GimDkAWqH
Lba3kf+c6j0g9KjKBMyPfwTrcoV2wBy8miMsvJVbR36LEO9oLaNh5g7c3QAlL1aJRazzJmTMHgiS
m+tpqS1SGiEBL9nfW+iwfeJ8pBQ7cBNDpdNBcJDSEAFoCw1RljjiYDcUo9jOuoOONleLVy84VXzO
q7pYYx/ZbdrtrRRgAMkn3gUG8QDfK1bVbuo7PsQTj/y8HCxACcpqgH3hgSPMF6Z9u1/Bho2tJYBn
mwTVzoAZMEEoe1Cw8R4W/TiPe1+kqHcKXEcpgTB2dxZ0toP5xCtmv8c66NFVyshCtf2/pzWRXDym
DcKCerm0VLCqsYe5uDEQ+enIaGXtmsuhDCON2DV0vlv7NGSCvf5sKmoHg2H8FO53U1tEGjHqlOA7
JRypQZxThdmJQhQiAqh6+DiZo/loAVYNqxjgq/SYlabBKZPR9EYgLOoKI1x3IOPXUjRH7xBLzmrV
6/eJoEISqKv/T5GAIeVk7vy8QUmMPMZAZbWrCUemL5sQIm7KWYFSWy3JQR3KiIGZRFof0/lskvwI
EvtUxJRO5g63xGuNKIX9judChflGUkyISEgExv/ShfQ6BU18Ne1dlyuJw9YA7ZJPp8EWec+HxjRs
zqo8du+bfg0ZAmCE+0SjL+g5Jttfo3o6R+RiEkmQoJN7adWUNdDDjEa9hkNokr/3YWeWNXxbyaG+
PvGsf+iyWitDVbqjy7b1mDTMfyrwFe6eecZSRMPg/07bjleJjIGpmiOXVkJImDevkxEtPWBGNg/P
Wm0YkBR/PJuq7JQX5SNnkHFUcAvsdsw4qYngsnpO8GZRO6IRvMnljqvN9ntMG8cDPUC4cWRRDd2q
9F5Frrk3A88n29idk6hzOstnhAH2MTgg4t7EDCIEgPFx7HJRKuBTI1xuk5EoG/Q9VdNMepLbT0E+
mR4BYHzh+MbTwrACoC4GGjwmeHArLJBWOuqZ7JW5SwHyr9CYOkxb5MrRI7i0TNcsS9Ofbz4JU/9O
+Lru0Fxv+rV436fMWt07pVhEkNOsEbWI6NVQZCQlhQFZL7A78YbF+N0wiQJHOLxNWzJzpnytnd+D
9tNxBQn4ldglmQ2f4c8E1G61r4TSQxwS+pDgUqQ6MWa0wEOIeAf80OLZKKvix9C5xl80UHEUYqOK
E2JJZ+1pb9rPVapoDsMDbuAViQg60jp4n3br3GXYS98cx8DDd5Tnfx8p/1/7v7Nw5CGcMj7wki/c
yYxskzKQ+Nbn6ugWfBAuNvSS6CswMIC7E3NUZ6qLzI4+W7VTfrP0RQDEKYboe7TGUU7pkoXug6WL
UdiOg848YB1bev5vmKJBftiGRG+qhduPYJ/eyDE9faeCAT+nDICi8seNdBJwyfAu1vMHNEBRYUHc
Q0OXJNwLHUS2dnz09B2QJY3LIRVHK1DR0MP0sSjrYPg0qRokYZPGyaI5vArGnSSn+SGB9fMHyfmp
6QSZGmzjB+Gh9HXk7II0l3iaDphewNQtGNZY3mm+oy62G3MHtmse1v8jVLOdIpHwnwAh8gW1WRfX
TFBS9ah3dzWuC5Gzu5WcGv/WfzGFSJLqQngbF+oq15ue+D9SPWdahn76/AZXXgqBI13fLCtf7Bna
o3Tu1zNa5g4tarMbTqzJYFWx3q+aP31dZPgfnk0kqBgToO1km2rbHngAFNFIsjGXxWeM9sdDa3gF
rpZDZBv3yMJ0VV5Bh9Ucpguer1yQNS25+KcL/GCOZF/9rLakCD9mCEknG90PP+YA5JjUdh8gsCLQ
ddKcLq0eKHB4pkfvNOkw/35GPb1rqVsOL/loIZ2kdFf1x028FMiok6/zmOSTWMeocgXM0x65NURN
a0r4fNbiVMVUYRugmhQ0Ep6GrDBrU67I9i46OPU5P5Ckq3a+qIe/1x6ETfD+m63E0+5QJcw3fx92
gUYHP7rMLe0r1dHQ+dzf+m2N2JjqNKnYkoea/VD0HzgLEYH72Op0ngVjV9tvVdimp1py047FrqVE
IHrPLmb7rUiIC34PoqDmPxLPYmtPVFC7pth61H9D3XFk27yOPaFITAk6Pw/71luiVQMXYci39xoO
u4HJEDhVpydml7iT4nAUBZE6Hx24+PRsRbLujdQGqyyJrCV20Fd9YwM3jJ7z8P15KmJWWSMh0j5f
NHIHrpXZ2fZObf2OvTVBn3z6r0ldLnHl0pBqWQfmD1rqiqdNpTYbSjGJoePab+MSTQrt02Vz+3gQ
clnOvBulbMjcs25I7Rn65wst+V/ra52h+ZyWj0nHwcxuc8DFUdlXMi+Jhd/1R+3qAoAJUMBkfljY
BzVQLKduqDCkkHjxf4U0tvqfL/jSeXwAd5ZMepejF11vHi5SVHJmleMmbYkt1afaa/vbN1BvdOlr
4yEeEFna9bqAm7md6vgVyxHvvdSht7HcVfZ8rjUx29OjitGPWmxZtD2sdllE1zxgIB1MlouyOXmr
N4PWnNPS7197QBefEVJIouFCVVX/y8wvdhz1hE3AfVDCCvnk9JH1uvl3yd8oSXbhmt3tE9/qIhX0
nkpTFLHxRMabIPZ1NOEuFtFwrDXA6ddj0ZeMuUtiPPEolcPDlCxJCelEH2ulLAevwC4Qjih3m+XY
MhxJkVrIL6kT8YKjpJnT4O+ifGO/l45pi03Fv3n3kSpaHqLnzPLVeKAv3aCFso5+rXVblhY2NF7W
CwcP5nDg1HJtDtPxxfswZTRB9RQSRZoa9A+OvyO3AE7aVUrxIZfLnZzGj4nQq9mjvpWXdY5zeqPm
u+Pfq7FQAzaymrqikWJXWlVYyqVVD+lgvCYynGu684JWat0m57+RSDWOzcDJCechVA26MM2Z2mDI
ArSpv63JXVkPbgmc4fsaJy9fURa+53B2R7RnEugWFrUf08h3IobhCOVyNWy2VHO5Lliv6IJ7Zfdg
HwahErMN+lN8BgQ8bvH1HV2sSg31laKIIBtppU3LXqWOL6BJ1tdsPzdVzwV5Pg7sf8Ysiq5i1Dxc
6pK52LeeODdvLifGXloei9bb/Z/iuSJWLQN/LBlYefoVx96tFnTEhaqpmI/zukwTKIw+Mim9iPkg
2oK+iW8ynH+/QWJCbhtoT5FA0h85JzY8WZOGLePkkf2yqRb7StCGhwgazrzR8CuUpOv5Ch/dgCew
xMrFirYVvhwCdjD9RnXTBBOONdBWUKLhj9vpkcuPqaNWnL8vtLBMRxR1XsE8r/8dytHLRQueka+D
Usv+k027rzlpuXIuyiV++ZyLQC/BmcEr8ocY06gA43rqKMPtHjS/7loHl0tmyipK8Nqr82ML0Vcw
PtT57gsyhFi4wZKY3WT4Uv4v1LM7GMjND+AoOUc4y6nr8UrUPHX7l8in732kTVOIq2C5TwCivRTk
sx+9O1VW00Rg4pKEtYNcIaFiHN7FDmET1rSCHC4J9POs20rFR3DPq8UUvz7RR2oqrZzNCXTpt3ox
Ict2TVcE5v4EogzR3vo4LZDFCX59xwMtK54RgsfROqwnjdol0Lbg9YqqYJE1tfLutQY6lYyIQ6BC
JhdIieIoX2kc9e6SuRRzv3hti1efndy46PT5GXNU6eGrnlosJB6OqFJP+fk5IG1i7iAQLa0gsJG3
F+LFFcIhSSnqoZfD+sgzZ++iNUrqnwK2y/F/Ki6oCK4qKxJRpQFCjfiAheOUXRLEKLZoIkp2EJt4
noquIiO3p/yJqh8n7qqC0kAIV3+UjJsnyfpOtUM+lLxp7D7NgSQ8W54aS2abIIa03Ls1XoxxEZIh
c7bHibzbFJpBNrSh9Jt9annIbOD5nMQIdH3RdpAaANJSSHsNPGDHX93VmcgvTiqBqHGnALLnbPV1
f176eNR29aS0geXyN1gxd6It/XF/ZDKKhTY1QfY1Pgn2uh6Jn+G44/z4q1jsSFL2ROctYJjAfHY+
whefw1cMM3o/ehiDVxzET9tXGDGfOCFfZltwJzGfNLEsIZrv9I8Xfg3h1iUekfD9BQnzRC5Z5PIW
ZGTC+2fgDKsPwkXFF1gTfZc9DGzjk6lINbvJbpxP2wKy46sMostSKee/ckChwv9OdJlmvoevCarc
Qln+KQ1xurBS9o0E13F9kLfz5aZZnzjJjTlg+vbCSekWRSbecmu+Uh89ZT1PNXaqWLSuClcuK+/X
bcT6nJy19rHAtmgC/kzTrA90wXNvwnrg4J9xSzYo8deZZeG8LatiYfe0HWuirx2TCg0HdWtl/Whj
ZqWV0Zcim2bTQb031gWp9HN9tQtwDGrXDqqJqlIkx/e6I3inLFdgRYhg7Oh1v3WrpFtpFtBEE0PQ
i4mZImrnmR7jGhRsHn5ve8DKAZKzG5zOjmcCjm4mA+VeZepBq1of71NTXlmDaUIVvVv1U625nFpe
o180wLH5ACUAn0U2ZXEHQ1ahMEIKNT7j6rk2rVnFcNAVCdAeFGXInG1xIqSOi9BSfJ8HT5ey0RhW
+wUuyryJ0yckygxTjiIw3b2IOQCvq3DlCzq3H3tmvuOIURBYQ9dysP0pxd4Kfp+QZruc3rqphfUK
vNmjG5vwz0IJuwXPCpUAuUaw3h7bq5hrgu3YpSwypguDrNMKxgLByjQZZWVad7kII0jHt6C8Ie2c
xFm3r8UiAIknd7AUuxb2yBQBSQ3pQh8WuLn/KEFF46XxHq2qEDnpixB5lEIvFA25mP0x85LQbW1p
SjJcH4gaKVaXwXHncnl9rDVVaSUWK34qMNAuDK1KoKA6kRp11pwMlB2LM5mLm4ImZONutN4ubHr/
FKgNDs+X0egy9mNWtCqiQLYDmXEC4ecODrjgdQNmtwmHCalXCw25U2eXbR+iUCmd1EFWRwxCnv8x
EKmdPUnxh5qseUG8wHfFOCaSWqKD8KKy1VWzmF9q/otHPh2W7wi75w6qsKEjmcXsAMqGMWqtz9XW
5eLzeNlWMxtQrc6JtchXtFsS8NxCTNXodSSWdIzvEtRuOsjshscfwtQjQAepFTN3TWd1CU6zgdhC
HUmgmK+IL90UcVu9oL6Cik7rEtrxDORlslJzi8oPgks1a8PhN8I4nTzvctMW7XbPqjlrzKF+1pw7
k0yfWYzBZZxraxRGoG5HfoCXajU/Vy7PjU3Tg1/0G5vH7lr2P5p4C88mueRphONs2vLzDb21eGwy
Jnvoit12636giD0n3xqzEnVV53h26dWn28U/o6fXEvCM6qfFCCakeExTVac3ytUf7mXP09hgGm1t
LcOhqAhkFCjXUWTjg6wrZw2sIOPWqsmqc27lKPpHim7sYtf6q66A5Ob7rwaOWOEySYmRX0HlLW29
3LaExXsJgXh0TjKpxES3GjtNZ1ereYjplVr0AmVqHtmxMTKOSXUw12jtaBELSnLd+UkciC3MjZj1
fN/V+t8b/KXKlq8izJa30PPAwWpWrZ/PEo4Qr54YE3SLo1fm3WwCGLnVGaa+/Fz7iOblX0gb3arY
zp4wk8GKMPEablKZG3xhaL8FJPsELSTrnQYgs1ShbKuKqvYDlzpKyho9RBndTG+V0OZWpqgmJXvv
mKEOs0KVVbrbPmBTtgOwLcUdq18r9zlegHmv7QGiGuJmsr5rjr4rPl7pcj7gA0CPOAz6210lU1Mq
nE9xN5iRvwQomML5d3HOqNFiuDRRjERR4h4q8cBRy/hTDfoTJr/GgYJJQozh2a5VoOVGPnb1Lng0
PbgkKwmmuoDMLiZJu5nPna8M3EAnMuI5n3tGnwluLsvL4H5g9YztM5/8HgIF/r8H7nriyVJnm0mE
29paDxjXxCOKIactrZiF4NF1NgbAzP8FBnwBppiIraTRstvq+rStM0rXQsdZmnlan6NDKB/SZ4SJ
6CODz8nMImcn/oEtpvzLMc1aWtEfky6C39X7Vl3Ft15ZxFNSNIFVZgSt/IUX4UMvkuts1i93/nKk
GCg4qjgQQUMKT1f/lJe+rYdCwwke9zwCYbhraaaJQkP1VGsv3lhashUE+x7MJks41BOPqrwRU1Xq
+IGcdjy2+fkRkN6ZQxZ6rnyXKmEkg6WHhT96I+3lZimyXzrhuvuYudnFbMuhPqHCZCBCcMzHH2f5
7lnfa7lxvX6OKuMAOlfTEZYyJguD6IQo30ORNreyPMok6OpY82eW2SLNVURDX8st/83WgkaUoed4
we2qbCV5Zo0Nh2OFxPKQADMUo90OSYOKqQabZF2UHQLwSX7Al1Z8GiOqFsLZ2WsoU8melvFP8p6z
Del8JQskpm0cXgYXX9haOAPzoGJ/I6mrv/eLy2UvtIMSHdVTJMNz0IE8nOq5JXKPO1wi3Ci3AWLm
qCW+2nyfo2ctctQaOTe1+NdQ5AUEkGtbuNb50Nvc5R5mNJ/NKiW8ybdmFfNdj/paH5HGY5v10dFW
73/xYYxPo+gw1xeASV36s63eHyKPjqaZQ3Trr6zXMTe+Go4sxj/E/vZl9L/+sAIYRK28LFkGjc1n
ferusInRk0Y7xAfxc0eAvax7MKVSZWceVGsoY8qZNugm76sXVcf/J7V3w/Xy81BBt5ETt6jL6+mR
eUDVyDLyscV8OhjIpJ5JrMnYONU1FjnhnPLT8SIpBtZvNE3Ucu20wETTHl3HL/pLL7twU5EVVMjo
p+ef2lZKZuWJU7SSKuTGY27oWc8GL+3+6wB6Y02AZRWuNyD5stmEyTOhZw6oYqOtI7GAFmUFNnfQ
QHOd9d/U2gG6qmnBdFHNCmODIPK1wQWUuAP11jNGxBmbukCZgNQouQ8BxFueL5SgiQHBNgc74WgY
nZ7myVDonwu60vqkqPEZ7ozhjtw6nHnugC73/rAAfWTU0faKFnkt5yY+9HhL6DpCmQWGuL475rJo
r4aEyWbMCUuKtkvqicpZvSZzmVjd/DNpk9SoXsxHEccECS1EkJlRFcTPslt8jRoVuo/0yVXR44GV
5e0DOG7GiKnj5is0rX5KGPHCEjLh/JcX99RJknvRKbehP6td+uAHJAeetbOLwhp+B4YTBbHjKsf3
6Dot2aINFKh1oTUybByo92U7IPhbdTeij2/z9G5OUZkjvOcge0Fh3DK3q50a1Jqnv94izlPBc6yk
SeEumvXSiloVWX1yuJK9D7IVnuhBlLUp+YLjaXSRiLe6R+qrse99LgeDCWDhpeTMctglDrkuWjjW
LlEIMvfT0soqIOfp2tSLIoBLLnljA8UCoAR5PU4xnbQ08ub3LPeJbldA/0SxEiZjmwh2pJapbHdH
cApMvctUg83f0F+7cY4EwQJ/vFcQz8jBbn9W1Droc5GBO4ksQtMEhhJxb6wDpL6M3e3ASUQfkJsW
7ELbPDLhPyjn27meogI3/O5YuK7kDrXl58VNJcgyhoug+ylIU2afI1eo8YgrpznY99hf8BS+24pc
lr/rP9BVInn7NaP+VCD2ecMUYT/bTaFq/ll9/OVl0xkucErGmtAHaXhCk5+HW7Ax3tOd9/VaXAMR
l9UVs4siJgqyUT9sBxLiFdrCCxO7ljUstHgrYbcHYggEwuD+UsAHFIt3PyBv7HXipILiwFBcnX+H
6/4ouTxhfiYL5eJpdq+ya2FyqdVSFztSVQoxFd/uXwjQQzEzFquiJfltuTUkzzp6GJXvTo2FiV6F
s22IwteXJIVMw7oYmNHjKWXO/jtLMV4r55OWj+xcYcKgP1Orz2qUGsLYLgl2Gae6D1rWFkKrp4pt
K98GDCTWvBELigScjW/R5dRmcAGyjRXgRi8Wl9mke/mLSpFzW4JOHQtaEZtENdIfFyWhZBFxXmWD
qX2dVw1RVjvjKiAopnzWGnBEIh/iaQRlB4HqcQqi5y+nUPsECf4efjpNN0mxyiOgijMMQkWBqGTc
YEv23VCueDdd3WDXEeVmI9cOZfyl2M+LDv+3PIr5V7C7hYcafPIA4tncUOLb9VMW9Y0EXGH9rQDh
M2YMMWSG0NLa8LysRNCOtmo8h4TKVZdRf19vEYIcqEfJGsa5QCR8NbGTSWGt0JuPP7wOYRJUIxxn
RQpHcLn0tErN/EkgUIRLHQwZTpcHV1q6H/GNDgpjiFrMziI54aYAZm91qX9nyR6rUFCWasfHJ10H
1HhPA66d5cn35yfXeDUZmz5+GD5vCe6fXwn4YzPfi2qsVW2VIFhWDwOxrnJaoiXoauTWu9SAsDx2
FE/zNmwv2ODkYHeoS7I3KIja9IEJJSTzUjzO04VoMyMtDRJjscvi8ipI8YofD62J1v8lajb0ghPL
DNm823KhRAeQ/CCWHgq12rGIlxYs/CPfxd9ujKWuewRo74VyTiQ6CGeCNy7o5slILT0TvFLBlcGr
BPdtZa0pz2sqVjPW/lRmgYdNTcg5suV8oDSg/D22E5gk1APhvRgravFvjUv5OMckFnZ8jJEuzjYD
DmJaFQfz26BUO0yPlpI1oxuiFmoU9DQFiyjL1WZ+cBosSHeI0JLIVZfbWzezyzh1vL4C0DGoiFIH
D4ZMN57sUeCkCMqvsSVpZsyhAxEV5ohw4ZkrmhrhjI12hKMXemYd3jYopSIADo0T7ETaBnU/unPI
hV1JKhqI4n6i39MUwnJw84RjFp7GoE+m9SqMYKADxLd4yPRy0S2/YYN4gQgnoadZKLk/HTUtb8eW
F7R4rh5mxh8bLR5ivM3kCimNoRDC8qtxVz6cXehRJE0D1IjKFYN3vmgl4JjfKuJCl5qR3moyFb9C
8quXfIxJeGFDHIQjuDFYvt4I/mujsbu+gWwd/wUYAlyM+RldJr3OYrozxm7wLS7pnOffQSni/HVW
WLChCZ8mliRAz7ayGhaPyWzW/gA9geVhpJxwa9xYCeLhlSyEZOrS5/qD6HYdnEw8DiNT8JsljmqJ
m2BEm/nmeNh5WoetZBzRekqG9eqOvSFeQr0/mNpoOhdreczZaM2Nlq/1PMZGaWuFkUzsYYmqX1rX
WJv3zTzDn+x1wAVgtoypXQBfidmOwuMOqOtcSjTWAul0SBntgmxxqoPoFGmMLTporbSe0tzQq7d+
SfpQiCCKQK24b04x65fwvQAH7omZCk71SoFx+u+Le5MAl4w0zbKC5LQyR2oYtGYmb3pGIpjeRTM2
0KnWd+GrsZiDrDbx0aWk3FkganrF6j/vOk1AtYB1iPjvHfS9Cc16lz7Eci79nOWnPVMRfkwi0CSh
8DeCqMsLYsRhoPhJ2aDylzu6TFytZK5Vc7sut3nrOtVIwxR/M53qnUp26cZKeDH8SUThGUB4f2O6
kzbRV3asZtHJDLEV2bszl9QkQ+bkHx/etWc2Gt3kpDE5t6L0CAdU3c+kvK1YXSzIJYL1lvlfc+qE
8W4ot8d5etJIaCyh5WKjv+N+WxOYhPlHkTxhyayGQIqspdML8+zJkfX6D9AFx2qlEGLLyiDQsdhW
HygdrWU7f0nX63OD3+kHnIXgvnum27EKOJk7fC6WB3wVdHnpgjvZpsq3G7eqd5rULYY3oHm2+GWM
NpO4uxJUpjF/EJVoJrrs9X+dyr3e1ukM2I/Fm/SaRKtOznUmYQcz9Xz4Z184Y79RVLOZ6Xb4Bb93
rewIHjpSgEPDxnJkqHjxoB2XJTjK7G70ku0kKSuRviBTD9to7EqAExTSDMW8qlzBgdeRfvJUqmD/
OFT8tyxdrO6YbleDgaYyBobUTTheB6KbsakyVBf4rUByug9gbNQTeiETxXDNBZ6S3OMlsNs5c4nR
sJOj22YaZDfV6zXqDPuI3WwSnAjqqgSO7/VeRpbYnCkucP/uMqbxMku9ABm6rTvzaFk2WXHj/E4K
QeuvOyNpcuksuK49EvGQSyIh+ckzE3dq0jr0NQAey0gxPf/lwKydOxT8GjaPA1zlIFw4fSz/X2vI
INX0FKTaK0oL7Ck3sjMRu7DAE6c+JmHcaD1qZSsXN2Jqqhx9/umcQDTxneS/OF/WAKL2wKKRsmnm
Zhb2CprneWGZYSxvVJxDOQk+tbQg+xyACh9Qoo6rcq3gmXAKY106ldTypF1ItXj1CUIXhYaMSSQC
4hjtZmDGcQC9F7Fc1Tj0pcKASpLnqAX+cOQAwme0RUvisSvqPMkNmNRIrLR0z9pnoWIyInGQlPpf
+G9csmcEdLI/vlCn13SKnpQ8lZ7Cx1dgZxAVPSVxcBZWJcv8Rl98O+N9hqfjG2wLlXjxylNdz6A0
aXJ0E35wSzicDeqhRrUVlML6+r7dOQOOiaPhVU0qNAkX7jAFp+goqQ/VDoHc6eYbw71p4r0bClsn
u7umS+2fPdYjgnmhmcQU+totK/9JMzeBAOZkfHFxn7xZXcKkLzAnur/LRQi9Ngu7a3SXMIHFZOKy
9nkGyCdsz+HZctLaA9IYXD9jTNLM//oR4ZB3nyLJs/ATmeasLl4LePnCzn4yIATQ+Ipao4gApo/b
0JmIJkzzjIjCZlgflNnViesZxf7aaxEpl80L0e5+V7wElbgSQ+U5aI3SiVgGlpXAX1ubBJxMgIuk
wtfy0ujSdXPepRjI1D80hZUg21SbQDqrhHLHfPQdYY9x7cxEzq+pbAldyd8gc6+IYl5BQ61LixwS
a2wORrRZxE1F71vd8Qg9I4dw3UhrJv2Q/qNvUsjrgRubamoBSuTJ4ZfWdZUq9dPqq9x9dbAAgW7A
m/8cy0kR0RWNL/MbqG1trNP+OemXGP/t6jhZl5YkmDjT91hNOt9i+IyACUJoBggqHNsHKs1nVvA+
BNc5xxIgmyLiLvg48FcB5zCFpX4vYfdcFQaNHhNKd8uUUV1j1u34YLvrWL5G98MTlAz/sS2R0wPp
sPpLdBUQLJ3cs+fuyUIPE6GmA0+Msk+19UYzezOh4LQSzKcjLMbtRDhyXBoZswsJFQr7sCinSzeL
R/ejY6XfR3rV7csn0vtojO77NyySgR4blqvkPWSKerHHrU2uCtnGlz0wjhzHQHEysVOEg9A49XRr
zgFQTDC/4xHKa3ZXjkyfwORYvTqDWgbsAQCmKwt2um/UcDLe7tdbUu8xYg/fpKFMK2ly5w7R0U/T
S+XhBrKPuQpiJAgcuLJQnWlyXu14k8WzRoHTdRFLgLnF9saBrVEhNe0M/RMW9dYwNmAdCB/sD68A
w+PeqGSOadjcY2EIxxpoykz4PQTYMgUSiGp9pFeFe4vo+FXVTf3JmVGXcTCYxGurMzvbStMbXilX
WUC9sZf+0qyBDDsrOYGIjOxrtNYjETQJ+vEZyQb/l31lSp1XO0mQGcj1WxDzVE/QzNYOtLztekoW
pC9SVGubKDtf/aNzP7xxX+VIXA8qoonZcQ50TwrvCw6fG5HqScn9grC6ev9jt63fTd2laa1rJsGr
jHyXOOtJSAZGuM2uBzcXav2Vn0ioSTNqpdTagvn4Xtp6eFqmes78En++jKjZwTLh3hbcnhoouYlw
dNf3nEeJuHqQp7N1cMH3hOXixFBReyw8dirnYuJWcERiDwpvjznN2Ftxi4KiZJsxYt42paAoV/7U
nvdL5h6jF8ESKwzzaqIxUyC3Fda2z+j81CCMwdF0GyoAJK7oZ1LzepqaDMR76c8uFrNBZU1y7KXw
T3LI61xDfvsBfzoW6/zZttRpigyFE3HACib+lPRCeDp+6hvnf+joDF0LDzpFvzzKuoWOoV1S/vvH
4bvc71PjqAkwHMx48LJFlORcLc6JRTa5nkYLUrzJ8aJ8VKAHx5+YJRRn/VXlNOxSGdtRTgmOIvxa
YC66mNrByWCAWroGC6lLxakhuXbHilR6SQHYTpYagqtyorZ0Nx4+BQjh7OE8B4jgV6ojzPrag6Tj
81ZDAK9CYHZy1d2hsiJgNV/HpDlXCqDCuFXkVvi3aFWu2ZjQYe3Q7j8HwSrC+vpOpDwyY5LNbM5X
a5Xt1v9XhLEZz1XgTcwYT9H05q2Yn70vVWOHxCtnAAY25n++OIU8MfEVGF49o3pyZZPytraNNGWS
m3aSqtMIQsIgGw2BxZD9nmQ4GtxvWqtB3+UX/5vbZlIzzNoQRt9RSeiub5yy6uC2fs8ci+DAAxqk
LLXYJW1c6qfSmmNZ+XNMxMyIGAF5mIFdG1VXvqBCoXQoyk1d3m6hNtdScH71BI9LAVgG8U9GYvqF
MiDMJqOOntD54FCgD9GIlt4OHjPwURyFhrrZSzlImkeIGaAFW25dSjeRWPevKRXVuiTy3YmkICyh
QndEhas9SnbzUNxES9Q5QDgRznfCNMhlVXvsWMavdzy9ZXkvCYJZIlaJX6ajfBavIEx3Log+V6Q4
9RY07zii5gq7xl7Q+K/YwtjpWI/tPZkBbaV4ImwwrkQ61EXHYnwC4N49v77JKRVmPyTEPTIt5LSC
ZeNIhdADNZWVahyjjtwllVR3Wq4rs7/QjmHv91TaSrLT8WzXP8/X8aiabxnCSTyoVTpRlSKEYX41
LZorQrFTGVHQtH+dg7c68z/8SkOcPf76zdI8lxWbcAPpylThc10l3t41z07TyhwV/L4/+r+Gu9b6
165v+yIaFeOTSxCar00LQmYMrdu42XYSVqH3evEcIKQF6xkMKRvzMBGUS7la3RhYI87Lk556mmEb
6JrKRnl9YJgk9QBiDI7q6tqEsrV/tgZcSK8qXJQaggQv1V+LRXFEt1OYGQTYxbXY0M3q2PovPp2t
hs7tOuOz6SQ/CacLnWwcrQOpBQBLfeIODXgKLObvHp8OGYTIm9auNMD/s1oFyyID0X0YxX59xYnV
6+qPhWOoyDL+aGZpa6qhhJAtqM2s8gKRIFb9XiGbXxz9+QqISsdr10edZcAP2ib7hMjgm1yHkqYm
dwQzZssqpRcZ0ooJR0wU0LEr3osQViv0xy5ZUcMD6PRXecQbpynDK7kEp60HCRh6Tof5gV7Y7EGv
Nz2s6BAL8sBVTykGvbc9PRyRIFq3OjAVZmNTzPZiE2o3qZNaJPpClFtG3oYKHnCHqce8+W12IatZ
HVOaZDNTtZBkBFnuzRgn8nlPkFh9JSEdpCA96CgW7rRjoF9MeIRidTHF1rrRk0hv67D8qSj+Qy7m
AosCfd9R/Cs7KApFmS5bCYwAa8+3PPsRD0/g8ZiPmCLMHGyTmPGDTgdwuaAn6G6ZOtU300YY26UL
8PzmRfF7RNlVj6JwaThSR6LknP/DiNFQ1gnjwrZ8vFP8uHxzLIK5laKDh7RFLb5IG/afCFStWnYi
++wmCrjPYdRu47ll12QXjS9iXbRemm9GXf4YiAP71fJvOPiPxxqAY+qFTjcUWROCQlPu+ATbvPif
iysygH034R8VJUQ/Y3ov7S9/KIzWvXGPbnS/pHHL7vIozBF3oRjSYXGyufJKgI1qRtwfrs990CzH
Jp74wzmUwdvkU21zoM+jjM1YLf1Tf+VX+QGy8SymgEjY4IT57MS4AXjkHLLZrKyvVaguuld8mWmf
7PIXDKp05ih8cptCsYzXHV+A8omdJ/BT/5MGHSqs00GHleTy69rDvdqrehxsZ2KnQEDAk+6q0rSC
ZkAZbNquXDJRtjGzUbOLHH9DdIq2LEJg4GFtlDGRVDYfVDlWUOAzCux8cZSHzyxeRmWri91RGrHI
C3U0o7X1KyL/Il8jPsAMFet/A84hVMCP1XKqYA4ZqLXsurG5Eml9UdfPFaGtrA6iUi0ohrQFVwmD
LLkErX2YNpLTJj7wflnsJs0Xn/fNGL/DkMUBdBJgDGzEkc6ijBE4LTl3UcZ5SWOmkdbr28VWTpL/
SC2TRpCsj2apVPw9kTL5o2PJCwClvNoqKzCkR2EEjOWSlKOO9+177NwNyIvqeXlMts/s5hFBWsqT
gvPAkk+Fk0x+5Q6/xmQ3UesSpHf6Fry3Gnglq+Nns6K0nQ8hLP4wrlE8mh4Ki/VML4TPghjUZvc2
4Wqhx3j1lt/FVaoFYNEesQ97wb3Ydx4wfO++78S9fQW+buh/GUiQq+rySTJyeYxaMquMVaAJM9ky
lnXS5ZLeQ7Cc73L1IAIgNO/VXgOv7rylcC7Kf0FUH4ZDYUWyUP5xOOpLLN8kNXCIpBFd5q7UraR4
RYxZmzdbQVv2kZLeQSVrACjgU8SWeavAD16p5BUmrfIIMhwzRsR/64Su44rBQVPpv+jbN8TmFq9U
F6Fx0hSxAVys8dfhbhmLANvicUmkZ+SmeJe9Ohn/eOn3cBoSwlKOyx1nvojTHmhAJ77ldaGASj5K
B9j/P8aHjXwt4qZQPRsMZ+X1V+IGIGR8qgiU3CPCtTfnaseDYOb9rnC/FukfNoRU3XYTrL2YDquj
iG6tw1A9GG8jxdjZwZ/ks0MDc0BH2VNM5fwk9Cvs5QWlNgnpmcTToeDbaoiRY4l0iiBWuOS8CjAi
Qa3KzDnkd8NnVkqzESG34kOhhrLrvfP5sKUDEw4SuFZ68z4QI/rtBBHN3YHF5nGPG7snobLoHigb
UMaAJbCeBjzGzZ70u9Aq6Uw5+28Sc7Az+vDT74jVJO1ApUbHLv7wybISqQhO2EQRiHK0grUyTb/o
mLrid8MofG1Pe9L1FXHkROT3GzSP+gFj9PyT+BXdYd4BZTziH1PdrvDnusRspYGxLnaKf/dLmQ15
oiufNAJiwq4I+8rKeApc/8/MBloqX2KjBlzztf/hQb8+vquidSC3OHPupAV7jolln2vEx+bqilhP
/9O8m7z83Sfu42UfZ8BAapEaNypCj22ieuKaeFQbTa9jJkQZ9GplwVR78hj1zqYDGW1MikYo2ekh
Wrh3J8Tk80Vk1epePE/Rt2u31aLPmNqnKOL28JbnFtrsP2tHB6jRJpvXE2wpzCb0pxmFy5Ou96N+
XQfusmPaJMom3TfXNGnd0eviv6Z6/Uwc+pvhG4W+Y0IjZ5AuwOcnXmFxrp7PIBSeB5GoeFwtE2eh
2tga2TTiITGxwBaDU7tR/qanA1ma7knNX3uzZPw7ba3tF3OvW4vXSfdd+fVJLmmJTeP8jCDl6JC2
6Lhh+a2Voxfqdx67FaSzYV4zsxvLYzXmlmIT50x024S4BhL0DEIpcEDOSSm1HjGjC/ye45Jka+5B
dqlL+WBt/287dzAqf3nu7MXAxjjGpc9O00nOBfPEk1oT5f+MEvdArxJpV5NxazXj/CkDi/9JvRFG
sZaMcvZgbJffgFt9L45cJ/7l1MLRRV8eedw1tXpExAUameIYx/1iOdIF/n1B90wuJp3NxQnYCyBy
xldZZl/wUg2ex0lCxE2eeBLEiJFHmwFxqQ34HD+WUE23QoG6VCzuR4PvC/rf/7lrWjSpeUi7Zp9l
bBg1zbkPxkPHNs9trXt15+woVN5hswOgNeRmdh8MtxtBDRIwr3+pmo0xZ8GeIxfMsv9MCr+/Et+5
Rw/WR02FEU1hHuEuFDc1QMxH9qp/PNEQXrFcBV58EEVwZV5lnnGjLBvLAiPmQlCqWEk4GwIvCcNo
UpL03IwGLJ1+5j+YsQv762Jn1keWIsqrDeMfRXiKBGrBI0JL+XSqUr8rnCfIEfrrKQZ4RtAG6yo4
6SPzJJ/uVPm8Sb2R5cmIp99amvHCxvxQI1iJfrvZJBhVpJ04/xmO0IxpiXohqGiroDaWKg/FhbLn
m4+KDXyWzq75xN6ct/7YgGT8GOGDDpSMUTi2Unznb8uZgujXMMAmgQ0pmoF6limjjabJYiw9lOS7
7kwStQrpfPGAKj+owke5RSN0K9aOvc2JUug5WStQ9r8ZbKN2J9a6VYjsW0byOu+B5GAy3+i20mhY
nRq0uDypZ2ZrIyVvucCKroROuGn21zPziDir6XLQ2Abpf71cWsm6wuTwM4tPn2b0xjhS0I2PfRAz
nK8Dg3XFMUYWvVKjKwmcjzA+HxfoZiBYh6/eIG5VEkOyOQhGWpyEXw2uy4RStIPcCR8qYy9IsK4w
XjW+KoGWH4nVBXS+7tkaBB1mABVFQ5M53GOFMB0KXtsKqIc4nIM5n070KIlWd7JEMOd+MSr8+hsl
pY91+ZhoqAz8sOayJENqTzMH5Vpd61WreVdqvCCVlV1rvAQrSYzNERvqjI2HLAnewJMXlXMu2eir
uS97pKQhwvXG5HQwbe7tvqMZw9kt366Pw1CrS7A8bem1nfH83567dY6GsImLPaZKvIZZD/NJSYgz
x7T2Q72YOJPxwanTQBSqDSPcdVkPV4T+LOvIFx5fu6eLG8bRD/JR1UaKFEM3dYu/dko8/hn4W6P8
pr22AP+YXo+EPA8pQvZ6ZLAK5uUAxMUNr8hyx3QqUf39aiF5hjzv+e1s5g2flmhxYfC5JVz4KqWj
UrE0NaYFuUnonmsF7Ir/G4GACxELmoxdZ+spTvS82d2IubiLDaQlhTbuA46vVoXpe3SybJXeHTLR
YcIQNBr9d8iKwJOmOyDM2a/0W4ZWYXu3V+v40lq83RWU60pLc8tv8UTDCV9WohmKHjzs/BmFRlVe
J4uy4Hzo+ALXZx0eY00loJs7GXqk8l/pdTRwfhWP8mLc6FtqeDsfBOf7rJ50K26x8IAhxQcqyfGQ
RilE+zhjJNcQXR6V3P5eYs7APCbtegZdZmQs0aZkQ6U2NcioGNHgN+wLTJZdUKLGy3sb2Mi5IIyq
WFctkrxTm7sjfV8nE2SA0O/16tisoH26G8THNrydwj9+vvVo9O6WDMqbJd8Vw/Qbqd2+YNqPXuop
sj840K4zq3bD9gL1JFoyp+AnIq+5JM/9xjcbxhn1nB7EPzuH0xv+NQ6MS2VvwxLb3P15TbpR+cJ5
2i+eSNvqTxXH1lKyitO1cF4TcDgMZ3lXUBieHTzzr1+oHovBXQY9HuBAeg9E8F0r/ydJmiVs+ct9
YxqJfyesnVOdybsj/96a87ZQvJqoAG1hDYBJ9iLCNBqZqGzevEbi4AqQHDXyY5pMeU44w5j10pIM
CNYbmKzCWeaHuBi6w2T34E6KafX4Y07LtNPcmRSyExtTGqUANaPEnhvBZAfBw+v8jI9pQVndGyae
ahlr2OQjbHP0yWRxbq1jhkP8kZsl8AXSaQsHvqmBH1tGAm38Y7Q+7UBLTD0Qu9JcRsM4NlPDLnje
AJaHqQO64W408XZvPtt9ngA7aNTgg3W94XZziG997KGw27mEI4sfQ+V9NsabgA/nKUQlmse/j+2+
l0h8/wydPrRy6FxG3V/oiPHiBSFWlPmBOSGqOQp2w2KKzlTUqlW7pwIou42dqCf4iIcjD4l/+b9G
g4OyhWVUynJ1bLybIxnwdG4b8mGfDIoKqkcRFrFLOPbIkYfmj9JFH9bldhFk7hadSvnPZLcAMQjt
PyxeutFsw7ZT0W+S26EVCwW6diaWK71w//ArEqGlbTzlAGWRGseAmjD1e8CE8iG+fE/ugifBEWBg
plnhyOIC8EgrQ7j7Fnst2F6Njbe9yAoAG5LoK4h58vZ+bnPP5l07wbJfFelG1C5Q7QK2xsKxjulv
B8Tp6LcjzBEdq2hYoGmTWTMenktzSqdMX/UhSSyMpelIgLGoHF2e5b+YGxXgDvD6ZoDKzoNEKvHp
eD9DmXeif9H/ueorgnHaAGB5Qrd+VDPwA3+ulT6YGoExJ/jlHq9bdDHj21dDY0ZDkXl5dBfearUh
km88caS9AMvVwVntvv33wYuhpPGw0semwKx+H7F8pNfRKibHxVKvvWjzyQDtBiINXjMINCqcSP4A
w/YYGeqh7UAamE5mT10lEwRTwufWJsoq5TYX+dyKa/cIOyt7ZDKXRPq65gufN4YjDSrhusLe74nW
8r1yeiIS3uzgnDvlxOoPE0IJKTGomyHUT22NC4a/FgN+t6Zjsa+sQxvAYycjpD3aKfLrUWyBIvNu
L519vQDzzTXe3mOwLiIlQiSBwtnMBTLvWpHrQmFEhkrRNPeoakbOXZqw249yu+SzRW7XsCTo2Byz
DKxOi6S1c9KenxUxjDPv228zjSWAfW2Bfoc+k7VjanvDkfldxi2XhNO7X8hQjLyZ13gb1x/KwFBr
oYjr0aRvZTWLob0zZS9I+CY/PuLJTgUNjMyF6cPkM8tVUKEbDSL0Ft0faIABK5H76wuorV5BISpI
BgzKM1Fi+f5lbN/y5WZAlsd3THUHYFfr7PyInMGwD07IymNrAcBXSSLbN1arwX8vHpTpHGLNxcTk
7NAeLJYOcINLAhgS3Cig33sXdd0XquhGcVcd+QpOOlzdUw+jtIwRIPOVzt1wkALyrHwSSND/73bG
UYUlvJWNlrcfFKurML8pSHkF6n0clV1zsFts2cTVYzu7pK6UrjBuLxOG3kqeRTxf2aa1oSfPrGuf
Kaw2lW1Kc7K6Aoynv1BAmtLO8PWp/qzu9HxNeFRjZoKKo7hwd1eI1mLLD7UDO8zcxitz8E2N0Ebn
VQ0GKQ9/PyJrWj10tx6KVN+8sBBBOws3jiCx8pUGvhvnXtAoxonR0rGCXJzZmh67rWvo+/AIZqpy
McdxAx77lPiuxW6M860blJatKYsYN2yk5pjFg6w6qo0PRMtXsGO08v+im8nzWMqDi7nJ6HjQu2MI
plctqamfFzbz4Ue94B9xn/6KmjY4DPruI45blE1X8yUDgFuw2R8IP6mLAMYEy5RVD3+hZjvyQWDu
AGzfLiyM4HCKTsHBAnq3GqfUJyO6zogHwDniTJq/ADaWQQ5Wumg6/krCWaZCy5IKFSprEN8NLfHL
dPPyNmRjrGXTZXYzztVwjLJ9WbQA/kzrE7pulweyqypA+p6epSPdMKO5+enFraSjnW+1UZDJ6Tl8
apjl5Y7DniXH7GuuzPtqZ39UVa1Vzs223rg4a5SlVi/azeVOoBzE+/+gCK9AQ6f5gHrFVolJgoa4
01y9uLz29MIttjQ4oS+vwpxbmIN2+j4V72gRa7eda6txXi+Mb1yCYySgFw+vu7HK7o386EsjWOrF
GBEOWu3/A8x3+dUtInwMnnvOxzcyqDbSgtwn6JkKEoKdKo+yLepnOxnN2l34DKlotT6nBYEVuhBt
1AFEZrpzp2HdTlApbAeNHo+A1ZkzHijUW9rQmrQKiGwOm2zlOYPVPbSqzA3rCdGrflfrF9MpD+N4
5BmcEJnSaJoikwC79zNk8OebfzmZrYKwcH+Ay8ZZHrrjlDFLSVgf2XGUxmx3AeQdZUHwNAuoSvTy
17qrcUM7cjmXxBim4ne6+gjl5gBPuIdIh0yFxsaGYvy9gdvgrZlll0sIjN4yORTrqiS0LDb1oBe4
WqUWDEqTLjIzoNG5QQhwVpxqWyRaf2LE9opr+AlYr0t/z63Vma22OJrWHaS4rNvgi88gswVZJRXP
Zncufocjw2QZzpQuxTsvMKuranqrxU5trCJQ+iV1PY70sDbA6NNHHVO+K4V5cKvx5QTtfrIjKqx7
ShsmFLoW0K/ccJhu1KYBTBYpUwZPNRCPmt2RF3PfaMNBJYb0x6zoQQr2DhQIaw0J7BdBuUA7fMgR
xTScuB8gZ6ROvclNRX0g7Vp6e4eAJcKOTBpWw+paNx7HYKBT622IWHBnRoUpbQTWosORqasS9hVr
KkWWfRXvYcL0cKCgseJaidQLq4Q0kLHqzwobHynKBSLA10bewafsYP/JW3PV8ZQlCe2/83yMhGGw
CVHaGDEQynf7P67e9DOhY6Qndxx4rSxtGWyrHMiQz7k/nnMz8Gk0izBr8cwtnSWIoAwkOfUaXmk1
tsMLHLrWBoK8OLPhUub7QYuf9z91d2RUQDXx5knCu+XDZ+/iNjpziYpI+3A2It9e5s8g8BQumfYQ
LnWCN7vYT0SA8rupMy6Ws8RpR1JTxnkXVrQSNJHzEqg0P6Z1qzQq9ePf+vyhq83MTtHW5HS4PFuV
75Yn46LAxhId1ukoVxHMM3y5xUl3TfFuRAPl1YtOHoMlrw4zqFASgzFzYLNMIqKIHJpXwTI505O7
hLKRSaH9LkzEehoyH2CvAfl8zYBAGwT1EjDFJYCa61RLuMvkyPw/cVTOK275q4MtaGI47GnjTP6V
X2EKn0mB5DRn3AlWLjWbh5pomlwPWoGlqUeALf1dmFpf2vk9TsqtnSxWGMaMDuV45ih14qtMVNVs
pccFMkoTTzsztGtFWehJcR+OLMyspQXlx399qkaIvpm+0PfQ1F+Mk8FP5h1ngfq438cSApy3DwKy
/V10qcDXYJV+LBwbDFHCCeSOOt8ee3BeDYTs+hYuBhZasnF5TBTVoLYXLxW+HKxsX+vK7oOk3tQX
cDbECa9hMR3cCgql0K+poqlwiK59weSG6MSWxH4QSe98uIHkBkWztIeCqMuuodVG4HqPoz00aIOw
vD1ha2nwqIdD+K07m8TLcF8UYd83WLpggTUbWBTtqEH33P2CVcIBasg20NUyzLymuMhxSUM3/hK9
+1g8FqU2ThTQ9DJaXZLN+sfHxUvGVbis2CW9Sm1o18C70UBrfszoZ7CWpfzcMOyYbwgrYJFW/Wnb
kikbeZy+ptV0KvgCUZFl4CK5+qInlglyxRlMiwIJ2KmAS8N+w6NaFhMcP16jIxK5YD4m+6VkMta9
va9EydPsTuZCPLs5OxzJ01EvZgau8KVdFEJ4PewwZMYIm4quYr8QUmI41v4sqO1F/BZOMYosJ5qT
zajvc5ZnhsSUM8N+6DfDe8WJ02Kr0tRUe5W8EU3UzrV7NWxGdncqiAuaChq1zGjWr94OIVYIx54v
t6jVme7na5PZNkaPX8R1Z/gFfDXQb+HOe1GOs/J/iMFjth0Lt7/jcEHlorPxPq16FIpkDFUV1XVf
TCfZMYBwl+l7n+3MgJPvjyVRckVUCrvsx2/mFi/nhwM+QhqSQ2fUcf35R48dJA5K+muQC4/0LaAJ
el9Hf+9ETZAlKFeJnXUmFuBYasbHfA1iX9jxkWS3dfHand6pfuf41uDz9AbPATOxz7Y4o3C3n0zP
6bRZZI4K8RX6ikfQdhXw1yrbERnzv7ZKdujWxZAjiBbA36C6mNxqHEY7Bg8wOvyD923DB8WWqwGQ
ePqzDCz3wra09piVYbgJLip+tDB5L8rFXyhUyXeIqYYJDqqBCcJsHU4fq7A8nOJpp7y+oty/AuHi
HkcPPAwmqTVpmDZ3AtwPIKSyT/v1Mtya2G7/VujfBoQCxZ4FAQXnlMHB1E7gasczcf+JFtUEpqpT
FZw32Un32/4sqCyneloQdAVunb+c3hU8x+y+dmmGXBnUrosN/NH+0xA0XPp3dOb8zAT/C5CEBIgK
zIxAxNssOG0C9yMbWaR3ckxBXKT3ReDAj9+2Ovwxcxcw9589mY0BtY26jAZoMHUNY8jCURMNieI1
9ujxV3KE4SjSfw5Ws2roxyRClod0ptP68kogZZI0ZUuQEwJ5hRWao316jOk4tnk8LT43nYtGEV4w
N0e0dU6h37896H4GVTRrVfup00cwdDs2Fo2tEu86ZC2AYE3cGekhlOcaxVF41S1saYoUpz87ch9g
xcUdcIIUrmgJL7R1TScZMRX/Qnw2ZPz9xTYOoCpehXrtx2UHKodvWF6zjdje96q2pQzDpf29KXxI
YYQQMudfv0mHKpmTd56LckK6JaNljFMsRDyaKbBAn3e7hEphRreBRpjOpRtmplu7v2MwK0kHowDW
DYHSTt0DAGxqP1laBbPlbTojt/ilik43uEaCneeW3g+z/a9KbjJhI+N6k3wGBFrqC1oADxyLbdCm
qBKzULpWZpSe7ipyRDh4ABdgNMUAElWeuhmnHFGBMOBb+Aa4XCd+Peli1nZTnfYDRzm6vDKHHFiJ
JO8in5HJS6yTj67aTb6kNsTiB91txarJVSARWlSudOYtjDMvfPRQrFrUmke0Ot33XicT7uJL5AGy
wjAlC88ocqm/ZwGXWPxGtA2QeAf5BTBKnu2JsuId05DuyMqkzq9GPSUNwk9dxbRI6v5kdakrpEQx
4n0klqeRpZXdh9uNaOU0POsLRGwB/eNrr/ta89HeS+tmRZEkosJX9agwoZ6nGtqV6/oIa/9a2zwm
snl6c0e1P9PD49SaNNIhunxmQGB000T3vTOOzcGrn48MXeo6pF/8LG+yr6tFWGcWMdCE2AqSl1k+
BYEVTHDFBx60Gdp/ssqjUn09T2Aoo1+dLs0/1XEFIUuwDafWQRrGiXeuPQ2ZpEuChqJK0MySAnML
UrLYrH2rvCc2vo7NJH9bXBViN4tFRHHLkZI3k20M5+fx5M2LKMZFder7wmxsotME6sPskiXPWt+h
mpqjFcwQ5aF5pxgu8PDpPFp3UGv7wXTp0xKT7IsQl9eBwd/RtjAWlKWjy1eKL6i0cqCRo2dBCZB8
Wqa8TNJvokk6a3aFhaC4IVU0a4YXSO6R22Pk9z8zPD9pjm9I3Y2FIowHnvkUG1mfQ/kzGPzp94vu
KxUjCFD8YTducF3m20t0RKuPGEHusodOq4qnUl0cqLxgWBCpINAQPsrNsI3ofzkNhjhJaIIfe8YB
eQnFJf3Xt6tC4ILIVIVpR4qbkO3656W8bejZoFofqzJZtjKfqqFtpkmJ6/2OkrUZJFEyC1W00fbK
s2Klsh/jrZCctoi4fQzhE2Nfo35xZFOvDcB7j5z7OJqTpYTrCGN2JNEUycTCAd9gtymlVJVLlV0Y
ZNdd2EvO+t8fqOPocqffMmVhHfy1mMmsJB29CEn7ts+GjT8DxMxYzDiuXLtakRLm6Cx+Eo1L7nyf
rUGnMjCPC1yI9ytSZ6r7aUK5D1CWjQo+cOey3AdKiXybZXhfmqQ6XBLQ2SanWNt6DSRpW4arNRGQ
MBxe8OTdeq8afz+fqRtR7LFsP69+Z4PGI42bIedSABLXGmjM/8oO0BmFfJKMeVU4SHFlALz7EvjO
bJnzsMuv9wE3jjMyVKVxKAF2yu9CY5WWXCRQ4KnC3MZMIt7TuQbgVCo5yMD6s6NvGD9yFDiUrQry
jxCYZmpYmLqRCM0Z4ob3gFS2eTYfvIaoJC/JWrvbYmxgOwgauA/VarvZlL2nsJHOGDb5Gd63akBA
fbKcJP2qDvnH4Y2fCvxuXgUCqFXf4o5QaBfCEtVh4buVdxYgSdS+K9dDPmvLCPaXk+MJPzqBQN2K
wH4OEhrk1j2MlPf2j0H/EAkJ53pOGhEuGeMSpM4gjeEjEF79nT2PaUJIzBiEjO5mD2gOr307Ern0
/r6qFE08YErSaH03YJleg1oRJQTCghftGTBLqGiJjGXjLhL2EcZI/IBfNnvtMkR5UP+lYe5/0AFZ
e2EPA+dmHE7FUgNXIdHYjmsmjYFkmNa2J8pHJC775v2xAPUo+1yKsWH8eJVjboB/ULuafnm/Kyrj
3qXD8VaV+Qvdd2qe8JewjqCDgbQ5PsjYQGSCbwA9osq+naAV5lOGcLwYSv90wHH3Zi46yaJMOIxi
s3mFMmc2zZYigvIg6LNK2fL83lWfumeVKazG0V3V9A+5dm5JUQs6g5wFCQMbgzKGm+rM6ZjZ1Iv7
qna6O4kWO1W2E6IFxAqha7FjbKH1BUl58rf5wKK6CU0uHLXOZ8mfVlBk0thK71bMsaKd+5b3GyYe
HpanmL+fjCgo8OGHm9bI9uy4hOICszhcHaQf53XgZirwbypiRtHhJZU7agNiB2joF1vqwORdOkid
Wpb/T331OXGN8f3Vl7tx/2+E+gQRxoKjvFChZD8KL4zApJwfUnBQbYBaktd/LVExPrGrk9xjCIrN
35PALqak3efthwLDNRgb593YhueCd8jRnfbklFj75XjqRitYwVgXhUnjCGI0wMxe5OR1q1PVxkLe
0BIuqazYN5uurgIr4ZgN/ByVDGEWMtmrnyBYnX4wBgCcqr0KXTBhNm8aV4lzgGv3ye9vZ56+FgJ9
vrBvBjipfn0h5Jxtx+xDOlBHP9qNYsOB31YQGQygrEGjoXjCo3oEUwY/T2dkzdnK5WCvNmot10lK
QvZe2tz6ecY/ia6rEdJIuACTL8YBT1WFLB3we73LAdF8GHgIyfxuRO+dfVIMh96ewKwT+ZYU888B
UkWNnTnIL9GpmMKk/+vjdGtBwNWFlUQL731jNSPrf8/WguAy2ErYP16f1LYohYHtXLERuuBRHmym
HPb7Ocx4Q71gLbu7TEr7VkEU5LtPbT8Xdxg8kJsuG8mwo9KltCl5aH+9IXAMd4oZjPQLH3toYHKH
ls+efZMjLV8GQYjasvOLJ97Q0WwKXLF3L9uxdtGWudYcvb5oFcOjzYNe7d74dcB9h0H7wnQTBZJj
j+BSo0oVFSp393xu2H4vhLwdfAozTHYUme71wmH1yL89eTjWtAPnJblQFu2eZJaQEF6IVS7OEMq1
8MPZz+msngkQQ0gcJZVLX/7OSiD+C4qXIBWX/Y8vgYY9jQgR+/b8FEy95R0jIYwJ3mW9NSsTFxfY
ciFRg9aB2Wh+2BMtZlIJBveYGfJhvX3QJLpysqP1hPpwls3RkbLhldX2lOvDMqwF/8XrLvUdNW5i
vd0JQLozgJjZ6U0sUFiJkQX15/qbXylo9EW6tfBlg88CSKvkcg7bcuyA6kt2PF3lw4SdtYJbAIua
XgSP7p+M7b7UP74ahmfPjdO4NphZyWR+PdJmiOAvhLwnMh6sq8M4QN+qehkGmLQf7GlKwNLjSdOO
LlqdIcSeeydAX0S0jOTbTt3Prp2CkFKk2Cw5OdT3s84nDExIDPBS3g+k3PrQ2jE5JjHqr4/1jtyP
rBUfQ0K6oAJKMMfBCJKt8/1jqyQg3E57Av7v4CwtLbLa0RSGNXKZleiSrldWYhfnX9HAaqiDmdRo
B/Qx1r9UWY0RzekOUFJ++6P3oEGG14w5M5Ybpa7/xmPrzctEP7uY7U74R+etXfcNqppHjDteOfzx
2ejxHOQduPFH4MZXtXE+oJQ+sUaVyYzrXdiYFtWAX7JeoPzJuZGB2X9pwMUhjqei42Kt21qto98o
KTDXuk0U8F52djQO0wk9vAxG2wi3oDDaV3HozAYwoZTlxW7cyriceD8t7DfWWq28InHhFMERJR9s
PCf7YQFGXGlJ6wcwNaSo28jokms1CEP9YieveHTuosyNC8Prt+hCFchSU3h8F4liVX1aofEWAEsM
/Ohwnlia4I67fWzi2Byh1Zo0L/ki2DK73es5jfNd9PO40auL2vwGABQc2BRFFjzXehRDm4VzF7dd
AKTJMGCQKnfDgZW8DixPkU38msPSD029deb3PbUP76ju5EFKD2XKrUukbLeaiy8eV6WaC4NEYFVQ
5UCM0ZTyyzWbz5/8iaItXi4/h/FkfHAnBhFIHLF8QORhiISvUvM/LQh/biDFxPHnlKFJI7bvAijh
rDACHLzGEFluRpNE9Idy3/9Sx1FfyUsH1hUFwud1UmEzTUL5Ciq1Y3fO0cQtsPN1g6B3yTvDB+8P
5/OY1cNHxZewBnogExgXwaoRX3Jah8aYeLXFMWmusjyX5Rw+iKst1Z74TnZMyaaqzu8f9pECpnjM
qpMh+Kc32B8SeJJNXcTx/0J0qbNTWxPvdxOQ1EZRENtNj/npf34UPMLsIpb/n01sfVaQvQSIfhhu
gEbVsIoxPr65Vg3SA1upjt6uWs9tHDnjrdAmUcd53VJriHtutu2fum5wgNCuObpsKI8WogJT9mUA
+9e6ikXYwNUrP1verr7NqeUwEFLZVN0FjjdCYNDkX57D2nnQ1f6lOAR1QZexsR5tYwm0lWH89nRJ
65nHEpAd/0NCLmoB3G5m8Ivnyr5kRw4gzihOGRPCrSoHfcp7kU6SiiafsNhgEYKGNBJV9F5vEqZ/
I/D4N7KKGz0JTTwonE0zyaieu2s+CZgw+bPIcAg0imMHiJ5IG9NC0hveoeqeSpSRFMXyeC9xHFgV
scFDbHiqBgnAvv0zEceqWdNi45aZ8eFvnVCz1YvEe01onkGr5I2j1y85IArJRmNR5K0evB2ZaXP8
f489pLpvGzwwsN14IkDT7Wa1Sqn9i99KqPC5NVa1ZNJqR3MM7b6DCJDEPXQhPsLC0+YWBDB++jIK
1Qxdcd+SGprN3/s2w4vgaqphpv55cMfR67TXpSwekFv9qq9ZrcPctdz+eziNMp/AXWwUBuiD6Dkz
2ZWdPJNPazD4C/EXuYTCX07OVg0i5EtpuqVXk/SwNRbtTnbCVrwxS70u7pUK+GNOq2idu5jxYrwG
AOJU6zL1rMfDnhfzxIoEvuKG8CB5GPYQPeFRv2svsRqmPEN/TXian5ukbXvY9am72sMOAbp8yiLZ
iGHzGUEx9Ha6X6OHH+2J6q0f26uZsSWBaZRWvXkqHgASnaL4nwyo40ybu6wto9qltqByQrwcha9C
Kg30VuU99TakvmutPpMY95HIe+GkHx9JUgBGUqnvRCpbRsq5RpbWFcsQM13QLoPKMXdYk7ofKbFZ
+bX9u91X5CNeNgXMTzoHG9obsRmv0QbnoZ1FhRwTkLXFKDlXNeSn1FANwvpyI68oybCidZ3wnd/8
DR+ZFRRsNxBxX07KuIsIpYnGN2yJtSahClbJJRcqW2fwgbMqh5ZpACxPTE0/nHAsBSMl0vpCvJxi
gUlDwbCpMrNDDqm2LQVX7jKJhrbtlMlKOaXlWCmO9Bnvsk2j49TnEveB0T3pna6uxEmss+uxqcT7
bi2IZNatBGbE/gVR+nuPit4PWlPNDsCtJu2O1axEbObUPZ1kGMuTF7ROKO/MRAdMGrPaC74UHiAW
5QW3x/i4wRepLyffj/ySvLiuq4LqYvNc5HxgLTWoFVbSTVTe/I6TGbyvYfNfJZIziNPvH7fkZcl1
BNO08/BHM6wTQUgHAJ4C052DaqWiZTkdliPt9tgnDCFT19wC8AOcratqVYrccY0Sopflac88Su/4
EDGxBJ1YnJ3J0ZugOsom8jfX6ebSwqp6qpo+7yn6IMNoa32a1TU389rT5Ix1di8yC9jMXVE1NfHC
wFGMe7+QucxUuk0HUXJ0a3xbP8JZ8Whbj7w+qCIJOqQwVhC9xg8rICS6iW3nLoz5r7yp/PVhFN6U
WZredE0+J4VTARf2iP1K90eu+gzCnX2LCSugvHtkyLjxiWdDrK4z/Ch29UpOhB5RTDSPEv+USHt/
wsnPwssCp1owqgK8zEI8uMQVoVbHiIOog5CREcPXg/fM1ChWMDSbRP+c+VXcBCxcRY3aiQpVd8/L
tuAx3IAnY3kxcI1Ymeonhv+4tzYC4kih3U+RzYUbl4y39tURvUsvZYxakCuAUDLud2MG9M4+nT8u
14c9Y0osA8uQhn7zPslvZMY3dPXPBoIf2Eg9rKrqwdkc4cd/PQc/KbkS0O23XQcU5BEpThZXWonj
EBwDEmmc8JJzN9iXgU4aihYNER9hi6bAqn/Lji980tv7qXHBX3LvKLB461ZMNMiv2IQtPL1IpneE
2uIR5E5bifb1FYxGrH0qi4pRWExGA/C9W3c7Lh93TItDBECuCHvna/XasZe40xbly3Fvysezbi9B
2Zm6VI1VLfh6sprRsPyTpsBTKuwmt0QQaF2/bpooiWdsQ2O4rRs7PhcyE2bae8og9SEPKz2o2ZlO
QAzjvnPDlHbyfLF53qOc9hVmOVJx0JCK2pnMNF1zfu9wD7cgthQEqssnWknDNZbhPF9A+hbpQQ1s
nh52Civh7xOZKCw1V90jKu285pCkYE0sl3x+KXIxvytQ/rVKJzbQ9AMHCkIM/4vWBCtRJrK3sFWz
IODNxKLwde0P+MqqrBvv3re0qT5O0EhQ53kWdRNevizkcTrzjNVUTS1/7C19RA93mhsL96l1hcch
5EDL6K2/j68KKyiRrlpC5tgPt/1wO3kqX4cviwX3Q1Q9lmG1mAgQ1lCDC70JkZR2O5PVT23phidp
3nPidYB88DkwOf4wo0pp/vQJPMmYmJ9o8jcJWcBKc5D4UwrxE7DsaKT9kXfHFViCtcNAJqfzB06r
Nb024RE4gNvWopriWgDjh2mdTGbPZxoegS048ejJDf9xoHP9DyZonwi954jz9QefsMaYAUNSORu0
0l+0aPg+YQM/fCWKpWAcpBLr5rD5dUgnEsVDPOW+bNEtY9hc2l90QeaLknJT5iph39gMYQNY4avH
VOagEQJ4o53zVsnMGpOwBerwQwyq+iMQ2JNWF6MxwHhV5fh4aweP+0gm/lxYAoHgJypnAtN9HiT/
gqkDjQF1J2pbsuMZGOyZXQ/GN4FOfLnYEycYXsc/E4C4bGK1jE8WVUW39HhXnmuMKmLtP+HAvYlU
/Ghvcm274v4T6Bt/PxMIzSmqdQlHFxuxkm/xsss3Yh4FWBjjr5EVe+jWkYtvzoNaaD4FtKneNotq
FQPyArO2dnHOIcY/XTWv1sCIjYOlhNYBwPtgrXO2Lb3DgEIDzwozSe15eUjhLeuQm9PUKh2oYSNW
hBEZzE+gAsmG15CYVzdh1J1oxe/gYJ8YY4MSVC//hbgt70kiAZfEJbU8M2Sb7Bw3z+eIs93gTw38
4ntY+pTDMcCD3qNvet3YOdXpGUx+CrxCFNoA6qV2igTe4mTRC6SBTT5N2SeDcyxD+YqNvmAuX/5M
U5XMVm5wDD+sJ5E9KZDaqAHPG0cUHuGsKB8++tpwhI/iYVEBoC4shUk47dK51usetT0tFDUs28uA
1dKIQMxVjrfE0qIQvCtWTuhJvRxFoXk4GwPG4vktwbKM4A5u878VNQYE5/TO/mIToRd8WfoE2Hp2
jiCeeOYpyNbQFqUbAvmJ17egpta65q8vmcCweMJFaVf90eL2by+Fss6HjIuE6OzdB6Uwn7nctose
Ot+k/2Z5/uJEK1YzIGzA9cRFwAmvbTSs9nENqtQxfl9yemeCfoC6//vosHqZ14kYDkSg1qu5A+x4
PCbz+CZ7t679rR9iQV/dEih4BbcmOU6z8ruKzSeuoNfQd/TzIwiO9yC+JRrb18TKjdQwaaTb865U
pcJqfE2U1qNKSVjgUwxIrDfJKc5av3phQElezn+DsLQB+1u/CdjJwn6uJrCYvWISbA2p+L/nmIWa
40W2YltAK50lc5LfNrsRDCa3ml4TOWQcmCZt1d63tVjHJgsocvFEhBuJEPAUlyGsFc0r7cw1jhmr
S8TtEkE0TJiIWKvu9yk2vWI6+LgjRtyjnhYd8n03Ef2QvbhyL10GMxa5WxGWRGNQfEuuzIx2RDLw
lmJVLxIaiGTQgtnuIp7RFPtc/xOUP3jz7A9V7moiVFYlWL7MojMWhYufDV3FRgZwpiP5G9TuDO/w
+8jMFUXKRPoVHHYvn68rw7vfcq5LAOcwRLaF8ZHs/2VvkVLdzdC+7J/7dMygT29APb6downJpuCh
np9/D4JeJ57JiBGoEPFghxILhwRGn0T/xSb3ojz857mLcJKbbvEZMOITHgca/oe6XAwFBtGVgfJK
E/ky+PyyzdvdzmxdwsE2OtwhUco9PsDs9RFSdc8mDifzzIisK86l3km0q/uzePtef6lYzRRH0IJI
Sfc87zSP7UGOoBTgsuhG57fTpAxE4cAdaBxd75gt+DSMvH7mfAmm/DIbfKK8KfSWL+pNre7VFIEK
bMgOBp+RfvnjrCYxVaZkZ4XFgu5+UiJ2RjCxb5LPgc08ShEloIJ8ZhjS/r7MRRfqrtO3VSizI/A9
Fsl3GltH5Em+Iz9LpyCxljBCbdaYK52nEk4UeMGh1r93rlW1POqOjf0mlVwNhwz1icnc21Nv7+Rh
4y46At9CyllyNv/G0PeM6YFLRmGl20zmnVfT4h2N9oYgjIq4MOsuOIwef4BvCdUGovEWhU/0tLUi
nOo0CgJmOF6EjeFsJoD8rQXLdu4AVVDW0TO/lDlZ7y/wENmrwhqUP42utmxyGfQ05b1WG5lSWP/9
33C4tqXe+vDMd6iTVTY3Usqb7zmzRQyKer2U8/270lWw01E/trXQK4rN0Cni+cQlSEW/o7x3Ch1h
MdTbRddB3tNO9bhHV7ofX+FEpOsyYe5FHp2zUWiykazmZK9oHQhb6xR4DzXDBfU+hnxWrBUsgmnL
LOkp2yikW3RZ7IcLz+ayYp2xuG5xoJzqFlgsycig1xG2Iz1YSpUFKpWQZFcSPGouNzbBsZklTVR3
r8BLD8oViLIdoD79veFi6jF/je4aScbkynDhMMmxVgT22EdHzjwwBhQKbXL3GqNP+25G5HSZmSlO
ZhEtlCVXNAgzxqvyMtRLj19YW73usOfBgz9p0Ica5lg51WAKRNVFyOziPyMUy2sIX2UEZJ21nQdM
pAEdbgk3Kj7G9/ey15OCHDtuNaVB7JBw8NsY2bGH1An26RVb9uX/phAm30sfW9eWTFdiZJnv8TEz
czspGG439hpFI4ljLK8wKrjpPtriDoSWGOf06Vc3+cEY7gnAllCR5PEFroBwBZyC9J5/iCDEU1gt
2vvmxIs+JuMxL0AReSILFmZuP5mXVmDC9hQDVfTU8oUMO1l0mbdOH5bZwPwHHRGIwscy2Y4xSCjg
z1DzT9hts9xpIU7D7Ev9VzbR1t+JTCVh/KdqoeV/oog8KAuJYun1iZFFXTVH87ah10tdiX8f86UB
fdhnNx3Dk8nZ7c4dtIpJDxB4N+3xBqXrtbjiKbrRK6pM6xiSvWHiG0a+KCWoGKHISipkkmT9H5Zo
Ii6iAr6cbAw0j71OwUSu4ki974fHhoOyC3IkAtzeeomupRqS5te6Yvc9eZuV7TQ3+izlo+KOluy0
w8Li+0l0ieG766WtFMS/JGdfg9H+WtoEYqbBinENJS1NHrJ17OyUYyFyCaWhA7GPDYopEQSrvnRN
romCOJ+/XWseALT7817mS0GNoYjbXXZWlF1FkyuQ3i4q+cQ0FkKXHt2OWu6Gyqk7wQ9Db7sR3POh
7FdvfDprgyPljhr5N7+stNasiS8w3jjafSD4/bVnG8lQmaFH2QJ2qV/bxQ1aOv4lE1K2sXXIFcPP
SpHlvz+X5Z5GtqRbo05wFuKf80oXW4p3XZYg59hj1iLzXoOVsjIeHL0R3hYE9+ZHQQYwgEVPbKa2
b8BiGY1ydkdq+gc7F02DPJltivfpSRLLnDEg8Gk1PTVKyh37XrWH7n8m2DcHkhUqpUiNZpDNexFL
IhnqDizr4fuO0InbjofdEX7NPFsoXPTP5pFp/4EUxhffhjKjgRhl/lqVNUh30f7TLTEeMlUIz97d
OX2gMKQ2W8X2+ZnasVAclD6EmKLCoeNx7y1dtaCFuj3zUiMdx0NeipLvnCsjY3BX0M7kI3RcdGBY
T/lmOMwUFnry7bJMBARFEOjJU+RTCB3lr7I+n2Vk9DN0y/XsxNmNStrqVfm7W85ZH0cB+W9qpsv7
1XsqHZqeUjDQE7UyPLRomnc1ptX1Sukjf0fUAsXT6eWFH4I/PrS/qly+Mz2RDpBBAO0YX3pE3qRx
BVj2mzxBnrXFUBsyaMRFbhyicsn9MdNL3hUWD/Ex+wx1xB2xIz9wJv7giT5ILYTnAo9hcFOUjF0C
yYi58SI/4INV21FGakU2a+HiTiVsCchHDU0xZrj8b2bcz9nfxiRtsuNSztJ8pXjKZscfuEnT1Xsb
g0ECKqJpVdTdZysh51JfgJszQnB/1AjNLF8fSra145sb7SOyQJYqZYAmRtH3k/gPOiBwIheiTBjD
LVqwPTmvtJ8Yj61nbU8Qa5Gfl2WtGjV1PBIMufGwS2ApUL6eJFzbu5dV+z4rGFyQhM5EkjXP2Y0F
mRdq/x89pGadDK0nFHXLiBKhr1o+V8n36WnaZlvtPjJ4tW70O0AkAm6LmCYLecmhdUPH7rZsG1J1
J8Y3q0pjj6MGtzs8KIeVuivqkQOLQjxfks6bq0GyLYUD8PHCrYulA3qPWKdNC3ZSx4KaKyN+AlQ+
6vWkTy5gvXedy97fU2z2s6zSOuVIvlvYjC/HNtdy/UcN5nP4CcjxV0zsXYHBxtYCo9fW2C4nUc2D
/djdK86bgZ0Au5Qkc1CzFdO7lobFS0+e3yk0FoQLy4PcYVHs9mu//GECwYe7W+LJLUAJ3Y5rqEio
cL/qXHtbL8LansuEUTewXi4=
`pragma protect end_protected

// 
