/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
bc4WnAkqx6dlMsl5fn3cAprcqqxHUHgVY/ImIQQum+cRAB7ouhGGGf7iFZf77q22uZ5IUqV83Quw
Hyk2hoLyHV1tsHXgJxRTk+FG0z8kNO9UiseME5aOM/+f1fcoxpdwoF5Nb9O6O9ouJZW/9wU+cOBn
deDxs8Fe2cl/gc7w+7aUoFn4WojygKnIaeby9NCvgShnH90A/5GxWomjUdPAdBRy04fmF471qpG3
rcDSX8G6arFIKQEh5UwVCLxQIuBK6e0cztUh2ocE1tgu0ybaWCTYOjp5wNkYHxW0TxCBiXthO/Y0
21pIqRWTmcspQgDYTjUBBMfo4xnplJBqhrkXZQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="ASJKkguRF7cNZtn0GfYOwaRh6RbIlcvsA1oAuucVfb8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2352)
`pragma protect data_block
Xy3DKr6jQ6T4G9Vc1bujRipQ5Lnfgs9oypvA5FB9A4aN2sNz4/+9uoQkE1Jfn9DvfeJn86scXtK6
FK8P+b4MBLDWDc6g9XYxj2lrCX7ykc+TxA+RrLJI4wERCalb7MpVX682ydWyyEOanE0DNTt1vZLk
px++FiA1i6cQ+XWDQNcjhXhAhw48VC8YSj57qvQK3PcL9jrLgp4iSZf4QvQUisBs3H6flUVyvV2o
Tvtch0FF8kuVw2GpvtNy/o7IFBEay7ZouG/5dNZkodl7Io92fecc+1R0XDKnIJHbVmnOwVnnGdJu
nBtpipM9W+k/Bwy/EqLGYJRvxmIfDlzRGHmhL5a9uYAHuR1Ak+929kZMP70fRMMd7smGHmdNx0wc
plMr5jRVq30/Po8jtkX1j5EnIYEpY3l8gbgsPs2QzebnF49YPXe4UvNt7LcCUaMCCwW6Kw2ZTde4
w9Cd7gcmo42ADdNSKFIwScfX0VXPISWlgsMffh2vr3swneXOKlZNuKpBrviHgN12bLhAEAFAnuMa
cQ/5f7Qt9nGRW61GZIV0W7lg0bflkHm4mJR8tqXpbKmi23mG1rrUU/xek+prB7h3QjMNV5kF+QnP
MePkh6aTnub9jULot/LuK76spcVrfdw7BPHxkV6hb/hSbNlLMKTeeM63Lxn38n/tXoqn4CMZggQk
nwnuL4XphpxzO2yrS8gDm9BfjyYhRPmxC2caj+m4It8XM2pOuMjEeC4H8z8nM9K71DyaXnQuqhXy
6mydqlAYwvLEVcMBibKkfxyziXeXaGJIL5cSxI9nqbbmny/b5GY6Sgv7t72CNPvjLh6kCJkH2ddo
NdY8XY76rtyPmEjkchbE3ucdz0J7PBq0UvNOj/iyzwZKixdW7Qnzch2jVNM6QMSg1opGKOlbgU8g
EdSWw90mGvhaRYoJ/o2wMeFuZbih10udJ48F53ltar0gnzj4AFSyJQn5Dln1R17SdZ3NjNuubwbW
qBflVMdzxgHkYdBWYegJs365E8fpo/Gbg1J9QB8mVAG8zxZHWogZKfi8FJDSCcfH5Qx8lKcEQZHO
zVdmg3ym9aN9NXoU1kTNLt7Th8clwgJTu1rre6dUjjF84YOpMfIVkR4QekVrWJPSX3Nkf9HpoEER
1SbaK/dX5aB+cZlSWLIAG1OfLbq8EcIZjgKpiZkeewtpbskQnu6XuIEWU8WEN1P6wkEqA137exBU
906A7jQL+BAgYX7B6hr/UBL5FLy1CPjYHs9c3khs0ac+KUS5lerqyB4yv/orhddPUeKXYAsr6q14
vSmmtZlsNX1niEN1DRP9wk7khy6DpyXHe3WDNJQCfqC4fsgZbtLNCxxx7zX4miBURvnmhsSauyUj
j00o4t1de5esrz1STtPajgvVsD1mk+3j04azqn3IRcFa4++zfmJTJX7zt7dJhJvA/D2gq0oIVHY+
XpP/aBGfgnHZJwj5z2WlLCylrQQbIlXBumhXTT1xS+22PDcv8zF7iqWmGd8oLIrh+E+EZtCLYoXM
Pz7j2OLp5SFz4POalyGdH8jdfe/PBBPXrtVvTff4kNXPuAUIFXz6+rH/qJsPa5skjWDB8P/pRet9
f7I5M5lQqT2ZDZGKyEA0zPELtmWC0imDSDUAezJuOuH6DMcD3jUyVpJeYl/RgiAZq7X8ZdXdlG/j
TSuUGf+GUI9qaSyzlHUWmaJvrFxNQMQoq7S+7bastCIjHm60LSb3gMK5Yo4p0BP95uQUo9Zeb2qe
tebAjtaQRJxiVofEvl6MkmPlzSyTbwXANi0tCLbhlDSqaM+2bywSHARChURJIxHT3tCzEaJy1EMT
mbU9zPQmpa+mtZHTSr1zPJxDx10cbrN56Bz/mycnu0rM3Nrdt4QFE9nbGhWuMqgyB962gxkhu0Di
fpJYoCA5YVkISEzXkFQdlGwGC475OZ2VIxs1b0e/dvqmjHySHa7I/aca6zfhIbPZ2EN/AdNNKOqh
jlkf3OVYJve/mqo4pdp47ilHtBjZMooI8ADwjkcgh+IlIoSsUayB15uVVEZ2t+gRasFToOjPkV4f
qALjIxcm8Ie1xP5tmlUY5Kl3KpmO28BNWaRAAv4cpLPrXVBCk2MgToavZWlmSvbdWHZUMD5MhUwr
gs6KyFbwZvLIIL+SMuY0wENp1DYBRXzJMvpyin/1099RmU1ekRwNkX5PUQuiDE8g1oBelQ4Kpwx8
Ux9A8FEpo5MvQ9YvexCRXGRKqfpTcO5NT9xyKZc8tbqA0iaAQ/puJnUCQqRv6A23kXJrgk+MJG/J
fpfxaXuhXTuzj4tAkGJfruo4CS+Yj9M3P+Fz2Ezfla4T2+oSuBeZOXsEEmVV/ydcaiiUzFy5JtSY
uZ0b6tcAku65uWZocYJgxQtkmZPU0PzQq8njvz738BWtc3hhIeJf1/CbgusD5JLxH/CMOSlcsdSA
YRciAYmmKZELJTD4d2HeseEI/gDgy2MqdIkAJVzU9wLFylu2w79G3U4HgkDQ1WBLg7PELgP4mgvx
618hjtmHvsvnMUX1Ckniw2RkF+zcU14+Z1Zbfu/Rlt2S+1/pk0JvqIuwqKoI+gn215CvRijuedo8
aDj2hfL8O4vI2S2BdowdAMlj/B2lfq4RD4aJnRt1JHc+LCNFHj0T+Kj/v/CTVnnRRY7lLF8x1NpO
708yEk8u5+qWFhcL3wynxWnnyFPMpzeVx9DWApZ6Z93HMsqLH+FLnCh65v93RILNWIWTdpZnxcaG
k70ERkjpPfX3jerqJLyNGEKRHY2FavSHTI69fTyWUlGKPfZYGp5hrSgQcvuddOLKx4gbMCfFLs1s
OWdlW6I/+uroeZqW3x9oCx0aWcLmpFBGTXNJsacfIZHP+Ik4Tg4JI9nkWwtaa/cZtsT6A9GHhOLs
rznaPE4TTvHwc5nq2SdEbvz2/socWqm2DCDC3X1vDCK1NwYzYreBvcAGXuphjLDfT5GPMuptEiT9
WWfGS42Jea0HrcLOFUlXSv07C6K0GeZ1oUD2WrBluwcve4zu5iQbnLDBvkHpty1XCnI3c1ZFUEFB
GaHfdaYekzGHKaxiyWbqgKUqb+U90icX2y86kpcsReV2Orahb0r6Wdbcz/kMU0u6VAUtV7YHo1Em
uovXLswI7tp2HL/FqwGv
`pragma protect end_protected

// 
