/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
CaihNQWwu+qKJWjcmdIgzgKIXQ8l3vMImmWHnChjYqoa51yMcErBScyiE64YZSDih9WCUqsVfjEZ
HfdPZ9ljuyASaDAJWOBnJBbhrePBDPO5jKkFmPbv80QoBXSWaNMFc5sW0Ulg3lCiE5qq9SVr7IMd
vkFVewJkI9IJKPXIqEiYLMio527A7EkzJrjUXC11BQnTYghbA5n7/6q2WIDOwjQ+BdLZXxGdIUKi
ihIieqBZEgdd6vwETSGv3sSorIwnUPSueC94L800xEEoFQmghwgPGvLA3IEIqt1YNZfrY4rcuvTH
rxE5ve/ar6tMYP0QdSitAf/UOVre3EWtsP+Jcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="IxINXwVvXQ/n7KwTaYrPoEaEACBK27oPy3cRIdl/LOI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
EiGu1ShDtOnFp1/lwt6VhT+Ac16EF9qZs7zPfUtiocXG7NFCRUrZFvQE7QROnM5JeJdM1Z0h/Bws
trvjDLQJcvjMG+ZBB8ZFzh15O5BtbPcrbA2l8stE8ZzNa9TA/441LDhlPlOqSfwWNmUiRZXXMccU
sHe7WR7du0q61ZRV17uJiPmqysYV17ryGX4zYp1sTJ/uTRERepqQjNB6sBfonIBcKQ7qp0lrq610
rZ/NYs5JEZgGDhH/dTOn4VNvuSwidG+w/VhLXGbylYSXlXdc42AppdOEMeGrAcXtj5vr936qk3Ao
42zbSOjgBMtmIldlLiZCmaPkoE796rhVmRP7t+g2dKS7E+MxM93N8tfZ8BEVCkaT5vVE4/11SQNe
rDYYH/qbJMzzwhySy45e2uUajxGeEn0zz//7R+2otpF0VT4YIOrIZ6SFBSugRZsz/MLnAa7iv/t/
LRm/+pua9owggeqWkikof17d+pDWBOiKy0q6QIcgg75f6NkjxmNsHMBQjq2qsDTxfiOmkQuuihL6
/79B/9HiUcjgUAusMxph60LRyfH9mgevRXwIdCymxVxHRCqGu548ILnEM1PDie26mU6friqxyls8
uyIpFpoyqBz12lto0HQ6+yBFRKDqda4KT5EOD1Jlw1q5UdXmQPATplvG22wc8zS8/AV/spM5hOPX
VQPPHy8MpXWfnjZd0CKra006hUKWprQdZOvItz3iln2fS29tAcuqt802SHHrlKJqAmmgntx51GtX
Olwfmzaw3Y2jDjKxtFyg/fo+HSHseyOQ0LZW+KePsHkvJYITc4I1MHcaHD5JKGUjmEu2VA9OOjAE
b7Ce2CAW8ICQJJnP4YBrVM1Y5BjkmgM26UBPo8oED3m4eT8qz1yQX3ptlKx/valQSbMZxt9PRi1Q
21u27si94fZsZ853Jf3YjyN8KFCuGWtnxgkJaHvgtjLmtLdUPTtJ7+8gGmhlZ8RF+xPOl11rdkyz
zPudddePMwb+A+nw/vvM5DfD3+k76I5oai1uVl71AnGl8S7aPjleiiT7v2QNPhx4+WYTvuXrXM0X
v6tY6zdfD/8q9Hzs7OKvlKEQTjmRauY2vO1cpLcF48H3adh25rQGVT7dMQkEge/i0HlirOY40D8j
FdIVj/GV5YAMZBntZ5LFn7Cv8ELRBMMdmbSDzVkf0YXLpMCG16tL/jcnDqx+jhhW1aw0LAR4xt55
VKt9eK4llHmV/bc8twLAO6jY/8D7aseQL+94OWUYHJZNryYgTQ7xzVhCgTnVTXREUnwTZFh3ljWT
l+n/u+jRyC7JBhHGk/84KQTUWMajOnMcRe/uba3tMwfJsKYEiwg87soIRrZFZTnJP3NhOiGPRbUz
72kiO88zMQmVCCmvC5kNNec2XpprmAxrCLhyZs1likL3mHa7vhCU3W6lYL08gH4BzQph1rxEd36F
YbIWkg0=
`pragma protect end_protected

// 
